`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRkcajQVnMQxKjPBaLZIaR7/J7zs
kEF1+54ixDuIyNX+QBxUIanAUk7iqIQDed2hUG0kfoXoL3vuow/GsZ8M3G4iHfWrH7YjpZpxAU7u
+39ASljNjmhxyj7sp43zFjND7KB7yDk1EnS5RQNQKgSwY3fvRC0feceeFHyy9eiKM0+E3KW82xi5
RDh2XoenLekPW3PgKxqpPoG+gCC21CBlAB1jv2k6OVsb0sJjvmBbm0nN4wPphhhkwJPqYyPtdgZc
CE5JzhNsel0O6jCLkBrxuiBOZlErCfgSSrBPgcN45n7QwDnqM8YXjIhK+rKY9SfaZs1mMjBvIXJu
5C1aAMdPPZCuSLqIc8c3INo5AGl7zHLUyS4zLwQssoWbPpGzgg2t/5+9ofd3rTN5pWOYIzdNJUGo
9Hkd8crZi+z3m2YlVBIxNnSNCMKqbXfECXSi6t2dUUJ7MOuLUZwUfX6bq1FMF9Luu25oBj+6QdkD
0fMCayjknP5i5/SOcQA6F5pLVFgcI6Y46urYwn4N77KBQjgBZF/s28/nnrwuZ8jCasHhwrgA6SQr
9svwL9CPjtau1p3G/Ek+6GFpZbFcQeLndmfaLn67fdS4+ojiSkyk6FUKXvXsDJG0qvfTIEnClnUz
xFxQgeQWOdUPgSMP6Q/a4kymClDjhspTVnlSFV9cQWEJ0Jb5U5bwqvrPFsS/OwdB4k4lH0cB7pdU
H6TSJ5MZ4BPK5OgWXlMEwpVbIkcjJKOioNY6iV/QvQVrrgdmaZbw6+T+NtwK11xtgQ4mDY4SD0Lv
sSWshew/3978F386Zux8Bu/u9KsrLu/XjgZxUzfEjF6fDic2sBi8z7NW+9iCLBTurA5CxvsIBYlf
mY3Px8X16lrjbMKZt/pqW34mP4YJ/XEXDBd9Hq0CKvDxQV6Y6/Mq3vVpfhuInYV4PNTTZqcGuXHi
BKHAhD4B55QkToMqLs1hWGIjCS2KqrDhfTtWW5u123Y0liGVjPMvE8Ws3Ao5UrqJ+Cb64cI15rvF
gd9JJtA8i92DsyTzHEGJ9Hy73CfcOZuZcIjBjCPF0AVVR0GNIDEOTtxjv/K3nDlNtfJechxhevjp
xbazTJ45o8dGry80dBugtG1NKPciDAllexH3sMlyI+NTMd7nC+7WpQ1BPw1Kemdqon5w/WTRwCw2
8kY89mB+3+sywOMir/pI375K8tjppPVnAm2ryaCmiatH1VwKe+s6zN1OcoKWdbh8hNHtt3Hx2HQf
ehWduYiPqLwq7fg/EE0av8r8UYGyUvXH+MgLKTKlTP2Z4lPtMVueHIFI1j4+ndl3GMkd9N2e3Ed7
gPAw7/hxBdujktaj6bY8xTLnib3yFj69T+KzkH2aCMobxSdv6B3YofMJ7W91R7sdnc8Yh//FwwL4
yG1jmY/xqip6AipFGrFKxTsgywwPc4krhz1uTBHKWcFNS0nhaocaKfSGlKLxeUH+aT55y7J1EdnH
E8ABGeMKuNPIs3yqzhHRTc889cL8jntcWwKFgPWjMBKC1Yp/aKxSkqHhlyA4MQI0PLqevF1H11u4
P3n2y6jjbQsTCfsHbmuCYFiC9IRpxFPXME2vcKaq2dmDyYD5VPZt/OJNAMd9RzVkInSzonVqsiLj
F2FClOxMxr9UvymGevN7KGvzgYBnZlNNPLTyBddofDkYsqHe9Clnql098h3NM3uolTRnX4K0H8Ew
28XUBfSh9TC5a1YXvtOYLHozU1QHyEWrKXN4m8uWvtyZ8hjZ+1PMMDSwara1X57HtujEHqxlzTTS
S2okC+l1j6e+uvkaB/x0EJzAUfBexUKmL3CctdsiNp5xGQgJEcmRxfW7qbrNDz5RgY4xwIJxy7by
0ReDum9w3Ls/7kSp67x405Nnt0t4DxwKKTWh890C3zLzhB5qLJkzB3EfSE7zm9D6oMTVUafmTVB3
ZVkj+2rbgWbkhAxjLepytjX7ye8ZyYe2hPCEo5oLL+TQLVJ+aGbNZwvbFrq4YmKkZ+DhnJlLJZrl
ST5qlskpu276Lbc9PeB8e/im0lHAzyzQ0cYnClByuKD196TJF3TshBk4CpKb9YYBQbMhvNdWg7HO
6tm4CuT/3f7Rk53PC1zRC+ZzcQg/OcMkpf7PxVeO9ulOy9PWn8XCUVL0LGIZsJGU/DcE1AlWg1Pg
vYwR2uqCIP2kyIaV1+09Q/Wanqt4f5tt7O7hnu4BQhHnuCPR1jOQY42rWDZCPvnAOyjgb/v12cFX
nEmkawp0QpMn5WDJ9k21OckhvLCdnw+EOm79WMSogAYBeMTLIJ4vA4PYxMTa51x/e3vf2Pp55z5o
CQqy2vkkcKh20uQVIfWissWdK/VgQCr+Q73928+0HbKDzIU4IdarYdI+uFmweu3XEKaFecMv6FS9
XzVnS+le7OFqiM8esZr8xPxqZ2o+/poZfPoIVyyQKxkBf4jQ289fcLUn3pNBeQ+dYXv2dbVLrLCg
rFWY7KduVt7TfMmhhl3wJ+WU8c8HN8u66557ANdiLS39W7OUabZN+No0QUG6YB06RWHb6Jy2TXkg
M4aXlXhfDOKG2saG189CM3xeC+sQit2cayddFgnXWkwqE2Erq5AdNXEVvFrifFLH7LeDdpq5jh9k
sbFvcrXuBBuLEUeH5VogaFZ4koH549+xaMji3SlvitA2bwScxHqtouVFDJIB7/ditRqxmxGueOqm
SDSBisZWpTrUPADc1cJNIPZ3jYw9Ek/pWN4b2hpf/slMcHKcMjEjqYdjF1rQWNkY+Un1XqsGkzaF
f3NOiHoJY9Fxisvf/0kdpXNm/4EOahHG8de7HQ7ChFAIiqOFfe5whLDp0jrWNWv+EWHIP4Mzpzxu
Qi4yyg0BFg7+Ho+w5Ii3QN4oF5uIWbm0svMjMTUG4WAUVmL+zd/JAlYHjZW17gIowGCikBz5W/7V
AfT9dH26zjf7DS9k4ozcVPRclT5Lrrmek77hQfI3lG0AZt8MvMPNVNzeqz74bF9m1QexWVe+gt+A
ea6WZFqsNS9p3hLh7F4z1HJBv+LaNm2UshLrc8Mqe9koBhA2cJDbTtAkV4RSBWwBNuJt39/1Eh69
EgVBPDV4ZR5dfoPJqmRV4KbgRMGp2oisOH7zpqd4k25dzi41kqcfADS2YZJ81xR8aG75x52uGrD7
AmnrpvObEZE/fDuh6ufHX9kINH200zEBstTZrPZ/HY7tQ65UAxLt6MoM51acyuSALp+q2bwLvBGY
oj+FCrxiM01oIwsU1ZjbIIe95NTLilseEQrQsqecRatXVOpgN6pIwnq7TkBdiC7VZ5D9db6ejJaB
MI9mtk9+2DI+ynqAJMtZzFnrOA/vQanlIez1Ekth9ZGOAXmkaThofQBLV7LWe6tm5KnnqTehttMX
l9mxbScSMwhP7WzwnVgOZoVhUVaUuAwhCprE5roHFsulNjNHoeGZa9xNkk8H2R8SN/txZTjQO7Q7
mR0LMCZSkVcwsUoVCEtkt2FDNHmYusIF1yg1xALW/2cPL9RRm0W9V+KXdPi6///j54FkTz61RW8T
TUNMOX4Fxl5sLjdhzQLFYQN74zcxzmPkyUTAPP+xKgUgyFBrhpcwrxJEZ947AjOULCz4nYVLAUxT
JC2cGQgsy+wXzSIWQQwcRl1bMOdlzyZStpMofpKikQHaqINmiaiCP/Efge6ua83fGAzDB/OtEbbN
WY08Szzq2hqV3ApIa1ZqBCEZNWvuckIaLLwsoIXnnjk1VuCFZOqueJ0yKjytYuabgsYjfmOkbOZw
nkL0k2t5J3J65XKnd7L8/B1QHC0pSrL+xIewW74q9vJCy9EGNriEk8KoOqAGtaf+58lowfSE0ewA
P5FiPS+m/qYTDttqvUQIQSQP3JSm8eiebsnOqmMOp3G5yZAjQFbXWTmR7RWirWrref6+iw14Szkn
E/LtZx1E1JfqcbKXYWD9CT+9pzlAJyN9AZufJlob3cqTdZhIuzu22vsLHi03S5O4dVeAsy7GXrBA
BBMKE31ZBEj9qPBNrwigTz2avrCvAHSOenhQpzTVhyWeSpOjMD5V44lV/piKUEWEf7KGQPD0CjKE
QWBR5PxpSkuN6qorvlI2ICr/Gqbx3tj8tGCEjJhoDBaY2m7bXAzBGMQdcdakCfSqLNhYVClQAgyO
2fYIY27ms7akwEr/b9uYYO+h8JJznsE/SFzMYEvKCAo3xwJZ3dFBZG4gMobxh52PZPKSSVuq9sNw
zIVSLSFIgU2uZBLVOK/ngS+AAbR2Agg1/y/WIxTXlhOyHteZjOoDKMwyexBxKUrELB8UF33Zlg4M
LO6VhFwyeftT+ri9EQfpzzIeHowAx5lr7oQfOhy5ti3AJ1Wz1Ia88QnaLQ0Q9bIPc/gJwTimmELk
D7azfVqsquCOHNsSVVWirx/WnyFzoVu0v+xjpwvexTJ3z6Be86AbXrPZMWvUMey3q8Qi3bNKkWt0
9IxlCGizOUgfUZlcyqUspEwDPuoWdH95UIN03+mZFNLIRtuGqdP0I320H0Ce7cks9fQ/5soYY0ba
8cbtJk/+49E7rjd93s9zFSSOKfTgQyg55lcF+5HwvsuXzOQZuU0jr/ka6YwmXOwGXU1MNnyJK9zj
ngWY5LAnP/ZuCrfG7WFsUF27YkwzecFtZS1wGK9flaARhPOatMDseXAdwtZOl0yKl0p5GxwbDGXV
MpsSsiJv/RUSi6LgZAsBK1tU6+TWd2MkwJB1elGX8ogewZa1iov+7drHj7ya+RSAwerXZinoKV+Q
pK827f0+uBU/6+VqJXZaslre6Y7o9NhD12PN+UNR2zXb3c3RO7oMyQ65Upqrhz2+wmvnGCw38VTB
wF8eWa+8/pR7db2bJmkZA4eeK7C59a/5y4iMUJomhbYgDBMqSMXESb7x/Ro4JsOkFqx+FbcgDWMy
+gYlXuOMel3Ph8BeastYyFA9fX3OHJm7HANfD+Nn+L1rSNpXUCDeBkOE2QIEGDn/At8LcCzfilpx
n/cPOqy8KZnzLP1neE1JLSERCjBfE9iDoA5QUhV1nncowQCJ0C+LxqDthbNWbYG8dv//DAUY/FUN
1noZIOQ+KBk8FrZYfAqHUiZcpfJv2RBAS8ym/1+eQ3LN4kKwsq+NmMVMDbeEr4pm4RGmucHNRV1j
ler0b5JvxZxbu4nMMZZgkT6kh9uNxmiXfMsiqe82pWnS3P5cYj3eT6oURoYgWy597q9XMT8I3xcT
Ve0X/EVpilboTTwRXVOvvvzXYWk3R9CAGG7BRr9uyxphNmhsotlVvkWdYWcdltwvSfrPn915x+wn
mnSuq6ZI/7EPlTukZQRZFWvajA/YG4ryVzJQaAad27Tj/boPsyJ5qIShk3bZvJf5LkQBfy02d9mS
PamhIEjrJGpC0dLrZ4SW+2xn7dluNWSU/00rUodLzCFri7c8eEO+mOOUNeVbr6FH+6oZunJIF1Fb
Sfaxe8WaZGeXNB8m9j4hrhnR4u+mddhpjTEIajVwdlIisr5EqVhB/ghYsHMfuxr20oRwq2qked6V
fpQtfSwc8bT3QoTsqh0vCqjK9+OewkSKrT3q4iJyZOJpL5sLWloW2I70JrapWI0TuzLF3H7CNWg4
m4SDQ44Q5KjQKr/PFkxBfgFJTy2kMX4jjIUr6mr1eoxof4ZLyQ1q2e7mScvcPkEP3mZJ3LpjKBJj
xxDSkD8MYAFLgu08Dy9RK/cUZ959/6n/OCugArVzK2fCg3iAvVvTKiQdB/d8+zfL5+UbR7Ct37kF
tQfuE7rpUZAz/TNsBHDlkRGoYlljxyOyBG2qTqBcZoXdrgC2phxZUKSJXNP7PX1ET7YbCh73Yw2g
lucypbOPzPcft34FE+GxFq0TJJI5LOPGSBrPM+ej2EeHUiFzdaHFspnezRnT1p+hUBFMnmEC53qK
7Xg0SLm2Gfk8zYMrf5ur8bjVLxn90T5HQWw3EObnVxWbj+FG39uYWvtQ6rBoFmMOqPL+4ANy/NLu
57jK5iWNqa8R5isd/I6DSXrx+txlrAa6YkJesrJ7VbRg1c413zCrJHCiTUUnvKLQ5ah+uphq0xVG
Kf8ACA5z38ZQu2Nbn4tuR1LSDY8OKtDaMJELCCUkR/W0Wnoa9UgvhHTAgE3PsUQT/Ez9J+KknVVa
6osGWNdcQEnSdJCpjMSvN7p/OyBT7mm/Tqfpc5FBWyc1BthI4ahZcgfxjz5TFwKrJ5NBSCt2981m
ddQ7xr8ZE4q47kaIQCe2Hlmpu5BVOgUj+sHJgUjKW4/n3ux3lReyOEwkCICKma0ZPGTkRmOcF0y0
glDOWr0sufD0ughrSnRab0iyO+KrBbXcx0ar4ZCrbwXGiKve6epVbOsTtpwdlmNM5vSotecnqHMc
c/SIGeyN6D9tKXygMFwCjyQjvpTDEvM4M81VNoxyw17ZKY5DpD93YNvBghTXZ5nFUHcF90aKkUWv
bRRQYV9tJN/Zc+26vwyxfNLlcM2A725ResbEnb22dtbtoHcRQ8zjl7BTbD6JIAlT3qhRxpKfYcSI
J5F8jFSsXDGPQ6B+a3+SvN7kNkQp78H2n8rOPLU5O1SdNYfhvCMVtTmQGXjMLTNg1SIigpfWwM40
p8ZgGdZX+24INph1iZitSep8SjN2lsCrGlL4q6NylpBbGuy49upl222iTU5uMw1U0DtPqR7ASJhj
RE5HKnlDBwD5gu+3oZWj6tdg/PsaLmA419v6VjWYl+vbAYgdnEXghUnq6T86/kXDa9KX7gmWHsqZ
aIDOEgoYdETHrCSaB3Mmt3ZtcRvf8yX27BQXfxQQp9LxYqch4Ri/HVMrDUZejdsxWXBQxZsrpqGI
QreOW/syJv4Qld0qCT+8EJq8vDd4/7CBj1w3uqZkcJESiPmRpYD1DnaC5lebhjo7hZi37bu0D7uy
8eraeqDSKlnsbVV2r0T9Z66XoMhyii8oEG8f1E1RZlXrE2W9OgmFvn3AeGsKZ4j+yhTLI+LjQpPU
Qh6dYPdOES4uZwC+F7j/OdebFcB/2hdmFELal41E4ZrnYFDqeMmdBR8DQ5dlusyeKB2MsyOONgnX
hnd0LaDJ1Nx8shmlhTr2T7myuiXL6NQDN3hAz5rRd8P+/Cqz/AdpLpUFHYX8Mhn58UXfVFjJN/Fr
rs0YE2pAesN+i/RnvgIJ/WduPDUU4E9pPMdRD24p5epQI4aSEypshpkwHd/070H7O446XFsUe78Z
5jIwFVT8Pjb5/irK+KArqF4nZ4n0UjyHV+BG6RkNVQH+2PqZyvSJjrY8gyC6HMFt/5U4YMpp96xH
lTAexB4x7AhgWdiUairmlOFJNEdRkBBGCw8prHMa8OSTMD8D9U28Iu/lRfXeV784d/bOS7cKYl5r
3g2Lg77rS6b1G82Z1LVAze5OqV3We8nSHE9tjX/gOxsRYvt/f48+d0ptB+BF7En8CCm3MwZz3S8T
bjKlO1ccicnNvhUyoUvHNv67LPIZdEv1KjwGENyyUY3l/gvlT/xq52s3OAFp2yPM8u86URGfvtLV
+cqf9JFbzuPvbr+2j7CksYZUtbfrHMrI9WkoWsrR5kHIGklUFigCyEQxATjhfRZs0/6U2BUXJJUh
U7rIE7vFcJ5JlLPL5STT6YBi0QR5qDRjk3AuewU/L3OGn2kAh1Ax0bbP/EekvsuPsZeVmP23oowS
x8wDkz7ZCth2ONJiwVwxayxBfItYd/F6siDwrHdxVb9noMs459ZoWia6WisSgFB+RMjdHbiVIyrD
zvterwRyvj6KR284nh4dPLb/6fpBca0ij8arxJdWx+BEuZuZvsBXcIc/076i88YbYaFFMVRoYwqA
VMzrFFswqft65riKz8YwD8etpzc8sX9qvF97Xip6rRRnuU8+XDFynKyLWMvnsWqqETjQp4Mbzwuq
W1jwxFhr7nGyEgHVnzpnJRy9tEy/NDAGNEMFMSU8qklD3Bcr83gswqv583T3fL+iIxrQrGbhjWt7
1X2bRiAwUbwbSAbop/Xl+yvJj8LoYoWSy7gbJuHSD8jtHuyJMh9IUwp9uMcsDVLxG9IbNfR06gPA
u7Z3vJd1bfX4evgdOZNiYJrpCxfg8eoQV2TUkAhqTcr8dOAASBqWmx/etsge3uQOQJtw2ZdCRlmp
ofQUi56wjrCwVsVTlNtj2Uzb1tuBrOedrd1aSvbvXln9qiqdxMLDrKgWdeFY66CMRgBr5jjqJcVh
9eu+xBF8xVqcB9lUsqs8kAmpqvo+ZukJjLO+NanwOjoiZ5zV7dUmnOdQryJVgD+WnAqKZBzf+ag/
q3modzxmL380t9AqLcIRa5lSU3OV6Mwt5A+2coCgiryH+WfgBdTpRX6hUAxgzDTC3wlRgnPFHn3u
gAeoltEN14lKKZIky1WnAv9IEPnSQykBYoF3Afx11QsiMhXCDWtVHS0X7HlJM/0KeN+lYlpmOaXy
B5mMzsbo/s52iYHEPcZx1plmwh2MFBL/Ba9hTDKFyTJIHwHCsCJoXXvdUUZ0TSikhkhthGvKLRag
ab4X+V0HLgIvASIj2VaNXzRx9JoHlDpSeI5RudjOjKziRbWTg9qJwdhVrh7edOB0APaxnU+OejaM
LPrBQGrg+9NkjOG7fFwt7M111x/GqzYO4BzFFgXK7Gnpu8C22uq8bD0EbKb3T62fyfr++ofZeNAL
5j5Ed/77uPqU+BxnUXjQQ2XaWcwtdWxhlZoi5xzakxVQuJACwy862B22p7bTGGN2DjEmN/6PHpIu
zWA6aIDh6s96RCCDF99cBjW0Kg8LPQHQyPCCxXCdfgdw8MN1jP6S6qp6tv7hwwzEWuBP72oQTf8H
ryTFmSe5VRe7GNcXjiVEcin6k/Ey+XSbfVeF/pD3fh4U/jmQ7DefAfOkdBhlKtJlJURPaKVUZCGG
LG7f5Wy3yeXjzklexuj4oQKT2SCHz9l3/5UJ6GnsqElfGqedp2m2iUt8MyS7K3B5KqS+4cGdDKMT
jNbPw6agWpAswRfOtc6t+X33Fw8abo4Fh+YN41Sk583haRiTo4Tst1hGfESMSQYh0E6vFFAtLfi+
FLXY0TPsnmBPX51dB0q3pZkIX76tF03ru91elzISAXqeL9HJv24k+Ky0FEHF/t1yO1YR8nbiIHTi
k7OT4EsVEmXGo6n58E86Uv2niP9Jd7Cs9JPsW8GqtytFiOHgCnmukPRffbzgq768GfJe8Fr9yB+d
aIWfHdkSlu8OhiftJPFsrq6f6bYwcjgn1VCGqUSreArwGvfSuOL+FynCOonGe2P/bVVKfp8OpHYu
BOI6CtoJ6R/jqraDWjkrkq+Gl9gYY868yzrW7Pgx3abD2ZweznFc35eB6JrYQLWhr4sspPa+6ut2
5u/TKleiqOMf1UnJwlhc0PZDbfWq2y1Nkzl7DftbfLiNIL3b2d9S8Y3YwugC5ZmgIlsr0UkqvN9a
CUl3EnjXP0ZNrvX8RGM5kUlW1tD1H3J4hrpHcL76OQ/++hiDxjxWExbSA+QY21wst7ixmQWPL/rD
Y92zOHSKT541Mra6g5iPeokTw4moHx85Ea0zLVztw8XIWkbQw8V980kWScX1Ax6qCmxyIBvpIjmU
dRmP1q1GOIbW7Vlcs8imBEMXSxbunpGew0QqWk8ZrP1xVAMMj67qTb8hD+kJdCbURtaSmNTxfT7b
wCOw0Dt9unCFItB+ywMQ+oUm6YDBgNqdFlIQBU6qJuTmn2ldgCZW0zY5jxyqxHhGhSm4mP/Qg88+
cdY+KZ9CCFCwNGWI7u9tN6AJz3pKuTmVnYunsuIq91vn/uteFzIDaPBHmmEy8gOAJm8WSmSMGM5T
WyzcPJI+lHuKzaV+70iI1eaemXgmN6LKZTaOvnYm1vVLoYh7YYz54Yrj4fU+PTECvoNS2TYliHLP
/hQeh22NuSifb9GhUpRKnxnIbNLbftpBkloeqvTPh7OpEDf2drddToqvUMl0lg3ezbxP/AQnq/BV
mpHI4tfpnMOVvCLccy+BoLibVStjkfIyzJkRCMr+D0T0IqD6oraNSVjEKt3cRSznMKIhZFCK0LhH
GRMtOO6v/mXDhHNNXBHGBqZEix/W9NIlz/XuayhFsbi076+HB7sjDIUBIsDpwiqjDNnNKYcsikHZ
WAWDmyGW8cv+vFXIqMk1E5DhwtcLou9StRy44+cHWz75U/yZ/Zw3LfynOvsh0wtk/xjjTvqL3g+d
9ys7N3pTu/9Fi73Ul3G5TD/fUNJ13z0luTAXFCDebqUvJpsW7r0m4cD71XpBxKEqJGcJRFLYG8AB
RzStuU1HdtGS/Z0+ZoZCjvKmh1iDvmbLujwwmPhTn2206DEAVPllbIA3YgyID89bR7O+W0xmp4tR
GIa0fANcLNanul1FYp8H/DcoQA6tnpBiBjrFpA4efs1OvNcIA43CT+mZt8id9aRMY/H8Hp9ANyc9
Tcr2DXPM6K+C2/Qw7APcU6vM/ZknbJcqlhlNJnWyw94G8NNW2ny+j64h+2jzA4tx7PWvn13vvWIZ
q+EgSjUts7PSV7ThJ4BRglPUQtj2RhtkVkNEvfFqb+hV7vvPq6JCFG8YaWMlF7wz+1Zy1O1D/2E0
HzSPEL8KYbCx+FI9ALYakO240zAp1isAsTKggeQ7jakRrxPeZH/JS1KkTPHb5Gse9G6UDlCTbqoK
ptyYwSleiNsrzEdjDUth10uYDb/0sZi1EV9C/mlObY6xeDx5BwT9vY9wqEehCRkS5eaHTuNgMjSy
Orp54wwN75/IpwP91G9v5nx8T/DK6AHf15TuTNMdjniUO7mTu1F4wmuHI8QrhCHANKFh3odx4iY2
bpYTAiUJGDUV9yq5eSKqat3SCJJ9s8N1YrWwjYPd9xacGBaq9+X721S0K1tEFt4/9WVm5RwTrUKh
90zzPMPAj1Dk37WTWft4GZA0ER1fLT4aPQeXkg6wT3DMzURFtRkAA9e26GA87HJyD3JN94/QD1d+
xcENKPp4jdVRxFXNVBQl43RftWXt8eHIGBsRZ1SyN3UqlBT9kI6BRU4b/JXMtSrRs8EVTMBnZbAw
2DNMwvP9AhdkMrTrX1BLkpBgzLNPasB5o427oA4Dr1JL0nrcCNC20NZgHuH+X6/H8DOMdAQG1iTh
oPWjwslYakEGP/VNih2tUFcjaA/XWJUSq+YQ9y/6feO/iSohoaCcQ3MsNY3K8hPTTKeXBgdAWePn
V/bRpgyNs+ZpyIebdqDujJWJVa5KPAmIKYEsoPL9+mxDwoGKK7DhLTRI0DNTL2tokjUs548NtXkf
g1OoQ9XjpqX7o8VI87pTK/jKSQXUoUZ8tjpbFR94Ruq9EUvgovmx6CRDK2Qhn6pHlxxSB2/S51NZ
tdZTChyQaXbLMc/vQIALQuNGTytx533vkC7k2lv4nfzc6xp55RIDqDB+FzibXW5bZJ1t3YSSt9nk
lxiFWkQlsNu086qFgqU76yNZZ5M1+EuMcZe+tbBPUIgxb4Z+Z9jNwsczExGv009PBMdCOYFiS8xG
ynj075yvBIxvvP4nj0W/LZGdtxqiPC0JMbQlnwYP2e9du42O+EJbkMJcGyj1VkbXT1P/hGsplvod
b5388cPiYS1WilJzVR07WCU2yy5GLpRBUycmG/9LtAzgQ3AKPupPW60BT21c7xonvGeVI75LeeL5
Yss6id7QnfdlFTSPSiJJQ4ocXWgpGPJwtgepB1fuIN17j2kfPLwsLUr+Iz2YZ+WgGbFyaZa0Uo5P
rV/xwXDtmGCMcD2Xq7THdB4VX7vvZdVDz+cD1ESbKrKbxAw6lbV+ahj1oLUyAWfbnoJfpp/xe1Ho
CSX18mLAEmREpFYxcDktS1+THXeLxZaTdMAJChrtscLV6o4kkGQiG/PV/fIRi59LwhryT6HqkApt
l/M9MdzP1qgFztaYSeFkdEDPMOuXVLcrk8EdlsdfpTtFQbZ5qfuAwhGerSX+bgCLAQpx5Aa2GsGK
CDYyx+0W3kSWKqJq3gsZDPTj2A1/pT2pswmb3UK84m0c85yzc+Ce9xR422+33FDPT6I8/iVTq7Fu
WVUcWko5NJffsBRijg9BPRMTIWvw3Niorp/7SSdK7b11bbmbHIWrV2Uch7Z0ULGiJXQTgRuczJiR
qeJYDZKIaXefHULB1mLUIITyOJ3emiGQn8HUqiCl9OvNSPl1t/MmZ8RbMfdM0Epn+Rj3rLYe5hTG
jHVvsZEJwyqpwnr2gA7HS1/XVbLjF61fnNALbUF5emIGBwO/+dQs/Wbhxiv79NUmvO/1LOxwvSv9
jyl21hObF4dghXhtwGgftY8NBns6WnqXU1oo2vJlBgbOOYnk4xFNiybjXknZu+BDe8mzXjJ4rKLo
x1d0ry8/hdw33x1+AQ97P3UnRRe1amL/ezD+aEl8l0aP0uUMWbiotUN6ZAbcnxxbZRxBbHiAUgGm
l4e3AanHjd5qc/ItcjU0J5X3jNr5zT16BDiChTu/Xhs0AbcaaXHd/b8OQ3i1wkgjXVlPxf7Car4y
zy4yziv/3ptVtdaR4/Wrx4WFXfwOpVSVKe2735sLbtOLpa20r6KtToYInFj9tQUYjNEmrTNbW5KW
f9prIK1Tb51pK2N10KRuvVysGqdWTzKQ8supHUoBo1C8PxCYXG224bYh7X8KNXzshSFazIOSVkge
vCo5DElNehiHcC1DZdhTI8C64PGl4rLeiyCb90yp265tTOqOSLv+wdp0elGbWblWQoZdEM1083yr
hK4NqOotbHA37uWNNxqwWliLMaXD075f6ehuyOl5TFUWXEW1B3J+1ERojcuPXufp1lENHc0cU4fB
Yw3FD9JuaeuJpLXMDTcwXvZQVq+flZyG0pumOXaD/1aUjwCRZdq8P9NfTOUkFdsKLQEWucNugnAu
7fBLV4zvE6T3eSVMW9P2O4EmG2PLSfbPx4S9U+ahu5ti7pYDHCLgzmSgQ+eDMHL2KONbf0IOGoF3
gfSp+zz9bx3ZFEB7u9CuZYxJm+DRD0LNyB2SEJ/NHsqI6f1dhIakB3jJaQIeCqUBt2UGsb2nHdgM
5rReXbIyyJAg6f7g4cB4aZtCgCiOMPB6hxX+KVKozvoIdBqpxqUROcVMPhijyuGpZA2m95/o/Y5/
g0IzoY/j3CWR4iViJtRUVaH0POfFJ49g4x7mdUV36M+YMzSr8y7qYLizvu+vRhskPjoH+Wh2ucUm
UQyEzr8hrt8wJdU9p/tAT72tbXl9eVe2clN3A9zICYD0XPKrykan4UL1gF/hm1Y/mlaegQ89AJTy
5ApEVcOl5HGbHahw1GRWKnNJKDvD/mx4EHOpxJK0F8R0y73TSwtHkgi7fAIYwcrfgfuLvKEjasCy
ub+DCPD3AP1LGkfyB/zJaH19IhlY/9vZSslUEK9C/Dcmk5mmiIQII1JUrfPmH3qC6H0Jf3v4psZJ
rFYrt2pDgT1DrWlspKkrU0NpYR4S1J7tQEfmnjQhKXCIpJ2ky9yklH/D5Da0UfVLUs1b6zj4g5s0
dEUZI05RYDk0JM7tKwiUp8OOjIzMzBLNrc/L1Q8TxzWuUVhH91+XC51M1RmrxN4KI949j2opBie3
NOVrb5+/ovwQhtM/xKGofuxrMOtLYTELUEanGJE9jO4YjqYVpQUrsHk3mjlsWzz+Tgv0A3G2wTgh
JbO4zGf7l4n6eiEfRRiOBND3NssfLXwKrc9LGSCbgo2WrXtUy3jrFWZeGTFesRXTdxEP1rtYTqld
gtgeel0rjNgJ3+6zpSlKYK+TQdS8cOJO2HQ3s4NgB0+O5U/CFLwPOJ32IcW45rGF210/szuSMz2n
Ls+SMdtAN9YAwi1Advboy5Bzh5bujnvbT9T6Bfqb2RnUAslEx4LvGr6G/FK56tGpcq6ArAJhCdNr
ixsQZ5HcjrWxAh4TjQFHF6TLcDVrKlcCO4+ZQ6jZPNxszuUt3DlbIuuYGT0FpXzAWaLUVMMtnKH+
0vxfNPFc9fUjj3rDt4OLuyETtq9SvKu7C2KUu+vE2exNl3Ys2j+lDSkdVoKZxxLEyI29WEj2Y6JL
qHz0RCUuL+CwQ/76ntZA38SbRcmPziVxc7h23Mpx+xvjzjjRcMfQrq4ou6fN6nDEAKnB0CZjBn5I
n2dxsvf0B4BMDQGcddzGHQxzN+pQe0jEpI9Di6dx3wrdSSybAeiKo3lqJ/UXNLlVpvETaENLQuqV
FBGejo045n5HeTjmt3I6RsygzkMfsymISII1j2/8uJOUTLreYsk6rmf/3/iTIRQuXRzj9iD6ad04
K5lMS63x5YAhcEQvQ11KsTHv4y4kT0HP2Kf1djMWr9hhZHSvaqhBpx7nJ9yeIJKBbz4znBbjxnxT
LgbgnABcizIXyvhGTWE/aCxzs2YoDuEJvjPDn3UH/OpDsANlL5rMU84TF+hKEazIBtP58Cu23y+G
eAyWCAzoqkxgrrLWlA8Vj8MySBr0idtYFrFYtHzPpcIiDsB61Xa6QxBz+g7i6l5seVfiNcrgqOT9
kl5aHyJWSTPmvpbojKz5JB/gt7aqQ9pqpN0+BLTCSLpmAyamzlTri0HJzXxUJzU65fqShgo3xiOA
73ZDqA2fFpO4/pFRDNWkNA7Ty28wYYjRsdfZ7K+sNKQvnQKbYm7djWvdZ0UY6NwV20LLfvcpXj0s
VPeIp71W+NgPudp04dM9NSVL8li12H3jgtTKJAgijHCXx7qQPUV187Dias1Tm6NUaBNp5EfjzV0n
2y1AeSksZfFU23nIJ6S3luv+yWPDjHMxZozU0+8ZIC2EJdQSlAkYx97OPFpom/9Z4dKJq10QZd6d
IFI1pXbOQmoIGXDHLZPhSvLUl+KPTsd6/fRhMGN+ZRaXnO7R2ZX+nvZ5B5VWfdbDQVWv8I1+nwXO
PaOGbu+AyvDI0OB1sq60vE000fRUvSQaH3paRyVbtMZDbS9f+sfzxH6MWxuz/85ZxTRY6J4PjJkz
Zcwfc7syzhdvREvkiv0RLCA85ywHv2D4YI7WiFXTpmdhDuW9EljmD4FXTJddm4WAvEJu5KlXBAlP
ulzxOxKO2n4ksx2MVQoEcMus/69FksqCruj5J4vYAJtQvHt3f5+GOKNxrtfNwu9aESna7TZddxyc
ldBPu7eTFcuQ/aPfL1Y5xDlURII2g5kUQEjvR1Iw9Cm6elit5fsUiJqgMm33NSqGFrmNMK7Xs6Pf
KgJpgCZIYbNG0CKQtFf4N7g39vX35imvhSLXF4tZbAZordB+zP5M4pMORRFMiLiKBwUPRBirYMPB
9fD2hv+9+vcEUi95XgOyE+TORzqe5J/JW1dt3lJesZBTkpePRSArTQClLWH9COf4AC1eFhiRcQBw
L9kba3I5iOEUZuYCgrGSMM9TuNU6WFEJU6+HQiLDJ977kKYKMl/wSxxWvwU3Zc/QTpwFxCg+wCFR
Nk7S1oYxm3tkR2OL9qvdl2hXXCfyQi+BABWO1/6WQlQZV4IQRJBirAmefdADqC4iiXS77xXu1XJ9
UGnJpy2DMo4zCCieSWP1fMk/iX5mhNALBLfkNs71kWFNvXr26x3aXg3OUJjriqocQmXajrqKxBQ7
bItCXrDtbs4rEXUJcv1AdH4J10dWdqRpkgN6RV2hwKAnX84i1htnTTUF1hmbhZ8wxG9YDAav/klC
AanFfzT3bBcEZhPjkRc1S91MCSRAthBwmSwIcOZQogTISrPUSIZfObGr405YBFtR+nHl2hKwzNRW
8J/Zrh0bwucdgmWjXuM/VpPhOhovxqrp6+ejvyPsGODa4+EwCmtPqrfuAlJOSbFELKYZeyMh1baF
UYd73SN0N5xaDIW6C6uC3YC5j85I4T0ktPSRdQrn2f+0j9tA2eGNf5NO33TTiWWm4Xp16W0h7SlN
y+uOGWkWGb4zNoCaZ+QydkpvlLkT6lijUDW24If8XcZ64SRPQ5W5d+cidsa6XD+ht2/wkOloZQrT
lRmEqvFF7Ry23klwb1QpuzDwpMaRpgAdbDeNzQOa9G0kEOqNTbD3l89FGKKS0ckwgUTip5FC5Jga
aUA1NrtTuhKRAbtUa0yWosyRTHngpT8PSWIbp2HqX8AChg3QXs0zCooqFOYtiMSlv6tDxflOxyje
Y4PvRdU8NsP6GZahp8SwFjbSn2PqlAvlalUlqwOl/OiLkDpRKfoIlqT+az7jj1boQKzlwinfYUaU
320WGU0xZ+Aau3w0GG/e9jMhOagcp7uPO6aqrid6zirZU0vBrhcNgfFgD3txJ/a9ZnhsZ7WL0l4o
KQatzU6sd1bmXiVzsuIvGoIt9OS1eb5NRNd3jdTOHFXu5ZcmFlbQttadFPvLWkt95CayZhxig+Vi
rL13PSuF5Z3eUWXayPRuMaYVotCb+QUWqXQpg7ShhwlgzT8TiA+eLUxMzVaBup3l4DUrdMIfprQy
vk32A7ukPxYgT8AaqHbfCDYFoLcsgvmx7E4YfOjSbsZTPrOsDVg1lRwdAjcpMoKW5cUx0im4om+v
FNdR2HZRsTBEKFd9jfXnfFB07k7gkfUigZxPPqo7K1RPbPcC3UTb6NvIa4oF7nu6v0m2gp+B6ybM
zgufGrAPtXg+aosQ4r1bfl5z0tVPdZ69MluHDYQbfaLrWS+297NasQmXMQsepnuilyoo6/g2nuQT
pFf0uZudavSJotRmFm0Z51viDQNJcNCnSoDfu3tbOQ6W9kwVc4vJ4NgVN15RDOaIitNLmb1PRsBa
SKiN1GSu6s7LLpPew/+NOe54837W9iP+SmdOCVxddZSRAYmIwKQVmLcWSvjpaxfhQksk/AxDPpvS
hHE738OdroRy4Y5bXn22gJIMX86827xjQTIScpeymE1liqMrIHdoq1SPUk8H8egK8cbTiicub+TL
k6EpbxM4gxOwH/H2OWy9AD2zge5K5xHPOsRqxUh2IRlaev68lBuloZNPC/uurNFIRGuWL7qMuHAt
U//ucbrIxGkeAvx8t3GDTId+h5ZIaUncPzG40rjqT+epNBwq5hoWMy/EgyQKu5bK/8jeeyuL7XQT
Q4uNJd5oMsJ0sJL/216DmS0ocDh8eddO/PdydxLqebpvlss6KHCCCXkM7Q8kiGorj5LJTsV0SccJ
fA7mHNQvoK5Sc+S9ePxDTl61ke+BMrx6mgKIxSUjHSHkpfq9yq+iBy/vCAAjhnuB3ODzJLPtTdCR
DSXcQsPxhW8HFZthlMIy7KV6LvCGgLS228l56R5gtm6/s5bnn9RAYvSrBM8gI/ayazs4Chhwoms5
4bB6oeSyOdaiVgxEKm+qWcgMO0e+c0/3xLgoew+RNHdu05TR9/QCnTMHtpKUwW2BX/SrzNRaH2fz
oCt0g2EPdBSz0c1ASUUBpBPn2c/FoaA2volcyGh3q0O/XZYMzMNsnvuDviF3kfKDep5cfNPsRVYq
FmxIciOwAhgo2lT1RLRqF5A9KAJKumfpGtMwzDh5NlIiQs5nTbMRlJS7vlb1eHgOq7pV63xwZzDh
gle9LaFPjvsDRCyINsqkENn2+G4l/hjLKT5UtK20tVACgDPYJOkeu9tquyV7hjGi1zGuXwYTH4mg
6EEXsVbGSUaxWZvGqp+VpmKLb2hWuqL9H3ABKs01Kl0DQQhTeJxdHo60FYJivZe2++nQtdkaKD/r
WSSASQZDIAfQhDZCdXqOhtcg+cM90D40egFW5LK8HhwWwvCRYBAlce0/XTeQJh1bHs9yS3BqIMWl
fy1Kf46x812Wmxy/Sveuq5UMae1aAfO+NNXmLxqqUS0VegXoeT11g5PXECepiM1k0nvrDQlpxdR0
afC7j/Rxh/GI8ZeLLCOFcN0CxiSjv+ivY8Uu9LJ6spmGEJTNY8OuLa7z/a4LYWekiLjEOacrgxBG
QDm06s5Q8foKdZC6wv2CJ3+rjL0F9IcCprnOfnbsSa2NdZPhCdZKbOVWUKCizSLuvZYSqoRCmyne
Ne14f/+X8wcICNS0ZSRAheq8tv0uG7nXdDHcx0OpoDJ7YQUpdg9uK9be3X83+FqZyP2J7231bnTF
5QNUyjgKupnakY+wl12BWYn2FwpvwG1BjHWpZOd+9nFOONUUkpO1ViFRNIKGmS0xam945R7xXRkz
yOvUkqf3v9Fe0v6HflTQtBXVdilhh19ka64dAch/WFrMUI+07ouPxM6nX/f8LtUujSgAdhHOOw3A
cU83YYAVc1ADrPxxiCsDOd0DhdbhMAK6akL+itTZvRht1XhMNu3Z3DmBJOOe9B1mJx54AUaYLPIk
j0WT0WQgZTeABseYG+hLEONE4TMjiga45Yp5Y1OY+G8zCZhaZdwfEoDh/cbPF+zB5Glz1lnkOtXB
hXYdR3QeJfKcAkJcf5+6Mu+iRZwuyQhpet7aUWcqsU7sVndsRN0fUMks59hM311cyTESbCbvhwAg
bYMe6pn9+EcLpfsDC0+pSrJp5PUb3NyGkmYr29EJbDlSJQH9YLf5rN7ZXgqbJfZ840s6+C5xE/dX
hKjStYOvBrjRlusqZq5kL0l8KcwbxNcoKnYwK+gubXDnRRfrbo5HU/sg74hWjXC82BW6Xss007H6
f+MThKOeznABFOWJBAgU4BPmS/VrG6QKKPZ7F1ZSUv9KYIngtKpaK9hr9FQJoNsm3qil8FY1A7ld
dq6TyOJ9Xbw/zyJS6auUM90iKQZJVXE1e/uRUSLoc69nv2I0+eVo/N+7GsSxHvaucymyVg8CzWzG
xG62uvEG81Y5TMcRFEYPV/2nbuXKYfhIaaU0RwQsYELo4tSYMATlKk1iEhJXR1cJqc1iC5cQl/fO
a9Be10HavnJhzSmY2KsZWqH8ktQBzhqqEYNAV8hagSh2up/6JoauWrH5gjLrGDhGmS4dQWVFpSMC
4UoZ/jV31D9BeXMumiNpJnYgleOBFVtT7uPjcVFWVOao4URDWDBv1CV4NiTYE+T/AhdikPI/5fUP
WNEzLf1Fs/YQzFmGQgJZlR9UrSIxBuZch008V1GPssbtqaMsAnHBZ6fo4Sc6Ll57kXyAP7EIYK5d
r1Akc1GL3cwqWUo8ANpO+zxqpTLX5xdHVd0x4fYRHUgweoEew1+o6wbmZf47BIpqAslhl1ulf3yG
Fux5liib5aVM/4DZgE10RwUeN47+Yeu+Gyi3JJ2oSs45K+I1aEUXHykilSbq6Q3SycPb3DE/0wGy
+KxgspLmJpsa3X4TFZQnsJvLFdAme5YXvkVODDMRkDkFy0NDpeEjm8ffRs3OiCfBzFjdTOhKQqbd
HtVnvQCoVLCiDM50K1bf9zoKXwhEaLq2/D3w+p7EZYz55P6K1IPHbYHdnMMVfQEVeUJGFhKl9kh0
cpsQokoL2pYxpvHuY3hpVZQ8Hop5ZLGk9YNs5MF0xlL6PgToqZ144J7Cp/RrsZ72O77JFRhXtafO
CF8sOD1AUcdzcn2D9cfrHtcFpQws1ax4+JWJGwXvrbJYJGzLUtH+VsMDHNiZhkqdbS14uj5k5wNw
xxe75PujBxSOkMFkjZp+iSsqYujYOa4JICP25Pm8ezihnrkf0ovm+CuNC6TPnlI5z1flrXyBlgs9
YOeIXzOC9/p7fWNNBKKSaDSHwwUCCv/4ukQ07ULjXQibmRz2pQaNj4CDGwCaZhGVskx6c5Zby88E
5Q/rHRrETFr09+ZfOTSib58wKo/1fda4BMKdcPfNmEQZpA6jDGTf2SNm5WMZKFJLmqjyG1Zly/bK
cswbeyC8uQk7pnwCjT14ghUfq5ERmbtu1MIRrVnKiTt0F4T96/lBep35t+TOGf/TNA8lyWh78+nL
BwU5fv5qrXTydQJe47jegmowQsFdnCU+70dWWgEIPmbckJdRu4w1nCkQEW2Pt2hMkDk1bqSx1QSo
elGlOzvWRXtaFpohxYoBlacKLkZ8DwObJEtvbBgda6UX8UJZ8wZnPmOsY9Y9d3SdfjcetjcgxOz8
aye2mRLjXgn/mGpun2+smc2z2tu8otfjRAgpUzFRyzQfqWr8o97ONCaS2SL56QrDG5K6sQW7paOJ
U3TND0YL/H0dXtme6/VWqF/vSdrn5u/EYfIiw6+W+lTltmD3RLp/R1MXWeby3RlwfaAa5HaLpW6d
Z37kKjZzVYKdeN3dyrEvLf/Gkai/zcjLTEEQ2YHUT6n+sgB6vWKoX9MDw59tDHp/QH11CjcAjqUq
jly1s5sHNA3UHS9I3RfL/2o4tKT3Ky9S0pu7c2cg0qizrJ7Eyad2hLtLH3UH2j+CkbaaZEiGSDVv
gyhSTVVvqN8+UY1n7PtcjAald3A+c5BwnIVGk+N4mf8giPZ/RvQ9eDHRJSoH0rSUyK2U+Wn+Fsjr
uJYGQGb0oJgTk424hqS2cIpONNQeeN8saRkrP5vGz4DTIBo8Zh1di02hHIjv0pREu9GU8aPLzwgZ
1cK+PypzW8Far22d7Micw2qGGSVU4JHfJUbcmUczpiZmHHq+36SX/7LO6Nz+uyLoxWt/w/isxYw+
XhoUjvxD6PP1XD6tBOkwMgTOCd/zRIEvruV5Vi9bHqoo+oMY0NXZB7THwr/cMwzXu42Po9uWwy6I
fYuhY/GINIgHgrxer3s89Dr7nAe5Y+Ufx4pEYvOK5+JHvLve5Y+egUKVMQsng3h/uI8NwLgOywSA
fRH/j7YqdmuvMT19CIc3nFCj3ig+skq7mScjZPVeu5Caatz9F8tF7PIL3VZSiQAxyI4U8ksLSg5e
79oSSqYMWHIDeAfmWEfF7JbIoBITZf1mac4s/oztS7FZnvebAn883cSktg9epgKiPg+m95Xbr2rY
lSpflB2cbkI04Ff8TTma2JbdSGcJxUVGGRJyZplFO114hw10cuBNIf5pbVkRALGTEL/jRY9hnOUd
NnbDB+fmTAmkOOxLKlHvbxO3em4R8QPHnBWcALqtI7p4piKE8G7cTsQc22QxJ+87mSrtOKaEwJGl
/xYS8yXEzju2INePHBpGqsZzsqlcJ3fQRC7WAF1O4Mg9Qe74H+94gQR9g5arP6Sd2TD6U7lQAV62
i0aYhgUDzKOdmB3kUyE5o6nYYj2ThZcTcJOFD/l6kWAHuoyt3FV7SI8FziABjytaO9iEvz91r7OS
gIxmdrLogc9yIac2zRqviB5BG3BpNEUJZbr4EddYguwn6TJUjt2AFeqoo1w/ceznZtct1vusx28Y
WYYcx5qxfzl1zg32pHDVvTAXxpye2wMYe1aIo0OOEouYYWf1HLdxlnjVChf2aWDFgpwdDXrj4Hx7
Ug8tzltBF7JDsW9NuydNZyRSa3g1Q1QJHIMFSy/3FfR4yELhxJxeydWeChc+T2Fd6cb4DSgmIbhf
ahhZeNHk71JxVtVVQcNPOSZX+BaPMnYoFBO4ggVOuzeLxuva+LbqmZldwzYj5iPnU4/qevUaWWEM
DXd2t/nk6/LPyKwpPW4wL8TdIsB7c8yAr4z+VxOsoeIgMl6kqJUSgrE2sIFTUdqQxZ4H+AqqYRxX
V+ChGSCFUJkIcio+2zGyTLz1BljBFVnSlK0j8cbwF1HsJjvJP3QDCno/Q+nz8opRmEjBsjgkHV27
imTrBg/SvadMvhmT5cLlTSlJtHz4GHxaQSeVRgmMic+IYUsuy0zPkyCogTYDaBwchLKoVUTKnlus
S/TVNeLB2Rmie47g3je+LJRB7UO/KlzvRRAmI95zDjfrkq2MgdFlvso9s3r5FQIkFDkoXuseePP5
1O7YCN4Qy1LP42AAXFFDjbJ6kfIr3hnItkMUQKt3sUzmLh1jPIvBRh4cr14u9OWjLHUGnu4DlH8j
fksPIbaLbsWfPDy38t9dVyQA1ltoYmAf/nK4/1/wWLPC6ZQq1PDTGbCIRFc7h/nE1vlzVwoJtCKQ
Z6bwdpOptNc3PdOnHElrSIfkzcA4F7i+jjE7LBbo+mP7CK2S6bpyWi/+KSmMosiTORbxoEbjO+nK
wYK0ozV6AFtlO1Z7RzLq70be5tTei49urlg4KjaJi7updI20VCzv/hwgRrVs6mDqbb5P5kbgG4Hb
ez8X7HbxmAGSP310QXcs476/G6fVhKYbzSLsTrMYr84NWYIeAedja8SUZawvHGesJjT8jmfu1oMn
fXbDB7CJEjwP7EKXORvgOPFfRj/QBCnzYNvBIpM7O+igUfilBdRL9jG1scsHFv6KatZbQ9UpQeyn
TxrMJN5t7HdTtfssyJrofWRxXsm/LI2CzJDwLtz06UhfEJKqBC3WFKrSEkQv0fp9QeX9gkdkCKRp
ipX0b99dVEcofc8fX2lj0IxFX8Lo6BSl3f7lzIXsy44F/eOARKM9wC1lVfJ5DWyK1o54QyP2lDd9
E4bnwZTD/s9h7bQO0LVNvcyNgi8OhMAmmGgRP9RGAxjT46/NAZkIYwjjYIxmPPqUnZuJau/phUK9
zblfPo7Y128UY3xiX97fXpSURf/17hwcGEpxAA5ehq++3IwqWMHugBV6583+IdxcQ73YPR+YZdgG
A0lQ+k82cwpCKTNJbYdCv1i1lhUsuTRZ6vWaIdxyZ4LVP/XisnN6NSCdkAW5NEFvXOL81e+LXFtp
SnIgfSbldGaPOGDnKoRP6dVfRH5X+xMvex/YVCWbCS13AykgeTgB45m5BQm7WtmOAYXlNPh5x3S4
+t+93imjfEHR7suWjLCkAm1AuW1WbGCjOnhijEbiXe3h34oqDZlKW65DwAOfAIIqF62HJUF2sAlW
zdso5hZK47v0pgPRLXjFosi1aAPygQrB/vyMtupXWZmoS1vEzgGTWDZKSN1XPYHI8GGk2MiHe0Ha
AD4UItVtc1l8cFHmrMLmmCmUYjt8sat9i4Rcm8A6v0x1PAtlEszj9pVvIYvhH8IXQooydCW5pdCh
1DxTNBR0cr8E27v5gQsh39kD2bm7JXBWF388Ovwsg5UnNx3OxvCtlAbbbJJF5hSJyL4xVHja3pvs
0l0f5ziafk9tMkRRhncyxfwFa9LYBmf4x2vnJnofHj4EhyUOupobzO1DJoJhe8dvjlwLooWnJh25
UWWwm8R/ZIhb62+dycT+nw/bvNSqA4lKSBUuRyQkhZ603KEaHl1v9W0CGN8ZBLSGxtqMt8npnTF+
Yspjzd29ejLVwqV9Bi/X3ZNaw+oxWh3QUduUMTR00tjr73HoCCT2cbH9zMKxoClOJLz/CqlQXFcT
LCQa0N6owhUh7RpKntutq/iyXNLlXlZRgobIW8hE58DaJhqpweKEmmQpfY8qEYN8p98Wy0AZclK1
FY8Lvu5d9kbj0Xo1IpgHsKaMBuQ2IpSDAtGPOakizG7OdmGe+8CT/KVLWx6hmQGKj7NRqVTl/geg
xnke4jMQ50XKWqbGBJX01d5OuIzhEHP9BIhs/D+zVGZfvjjklc/Jypun3viuyxYhEki7u3f3nZPo
vsnwvGKNxItKa2Qj0UcSAxNugMgLB4YyDCATPWKkPQQrE75DhNYLs+etaKKeS64I2IaQBBuUmsNU
kvDnDyfRLp+k2bDE4AvbV1Y92JVuxqWItSnai+5eMO+NjCp9o5vwsrmwGyn4f+ydVWR7tKVCA2xT
KpnlxlgQEdnxP2hpp0MxElzoFKArQZJIAL8IwReKHzN31Lz/mmid5z7AJZqXWHvHcrWSF9C4b24W
PgH8gfeaeJKwimHqHUbc+RhHJ4bL08ea/HC6nOAWRij85J4yk9Q5etG9Q1kBcZM7xTWIIZfZSV5r
qL8Cue+7xIuSE5MmUoAlXSUmXJn+gIQkRLVWl3nvk8fp2aZ9zOZNduH4+utsfnVocImsvEUA2pZ+
rTMCSfmVP7JjUgEEdqy8AeJem2QczB9p4AtSH/Qk/1U7ytBX3qinc7BgOATKa1cdxDnL8jD7ngWM
qFYJIVOahUsMEQlIfnZx+adEJAMPwQi12GnANy+dWbQM3Xx5x5+OcHAwmicUf9bJZ88zKwtxYUwf
BWw1Tdy0kcUJvatE6ZKlCnnHkCd4kR8BhO16cRX4l6U1PN6fOKOpIvG18m5dvxdDcYcyJGguGlin
I4o9O5c0sYW1j8mIDM5is2GRYYVrgnAoGmEd5vBMEGNX45itEUTpG4eMU16lB935+oSrv7bImRkx
SK+Gs+3eY4GrqKVZ4Dt1hI5dI0+NPNIuU+n8WLjilabk44ESd+ic3Z3o44TvKjMB5p3d9caDqoMC
R1UpgjTGKewSr1RQGPR9z/tJUgL9Gr0Wgo3fS09Ikn3MfcDT7sFAyiFQku5x6Pziy7yl9cqHxrZf
zb/7UGPT3XaF5YTJwYeN/f+BE5JC3Im/Gc5Rhi8bX0Z6iDnMLeia8eF4LIYFMQ/BXQyhIvkrPZYA
OnAldZXVmQN1clJbbt/dkbzi3KTLTdaLDZF3LEd3t9c0AouzAtNHAs86hLitqJcCe+mey71AciKy
pV32PE+L1INr8IEKnZAff7CtYQeDqLLDCSCuA87ypoi0vjsHrCHHACF9GSqQUSCxDCXvEiCjqwTD
aFKQ0A3m3yxnV+FwQB5bwEN9e7JNN9w+AzY6fJdFzdHA+euc7xz+bNR0k4yFIdqQPV2g84zZ4ktS
RewfHNn8uIDs2MjaYSMV9bZfGKmmpHrQ2Ha38y/K/Hwqu+0/4d9tJ5Rcn9aSetrvHuxX8jBj8eR4
1a9s5MLu1IvzUdf0LdcTzBvo/FnZcx0VbuwlDy29qm4SwzUsVzT0GjLELdmP9rcbyx9Psm463n1b
WSxDpMjNjquzUxns/R5FmeOtWpDybcIjyR0Rb+ztSKE91TL2ivshud4BtIriw8o2ivc9afNAK8o6
R97Q5giet+xWmsgqhqnfcW8RtHRZq3HWYZPShZUsIX0e7UEHd7PxW0gJBSudxXIXF0+jzE5/0mG/
bxS6I7nilMZiw/yYz6BQWchyjac+3FTrnAgjFvcUHEYGmxvC/D5YdZrIDlR5jhWVUKu3zF7jFw2u
BfvGD51qEWDU/64ou3gFpH2LctQRsezAscAv6/ys9GES9t5YSUjsOyuSm0A7goGF03GFH5rc+1/s
lSbtcXN3F/TvQpDKy9pIPuBh+tVJbmVvTqxgazaUHLDHr84JgjB1rXTwhAndfK+h0vXT9iUz/4Hr
tDNgBuh8xBPvyYePC1BfP7LOTuJ/u514uSajHqHBuayJn3AwclVr9NOc9H88DBrQQlfzWCyrp/Bv
HibHbjwe6Ka4CSdNbz9insIKkDnPpP42W5iKAjDEy+BxV6Rkv6dZGTF4kV8ckuGxeFib/HjzTcrE
C26eTi/m0tq9f0SWkIfHxxuKFELH86pw7WdOxxuFNmdJPofnS6iij2iGU2auGQZq8vxeiprvtjMs
wrba7vj342kgZbCtNZzYTdtz+puhwCSDGT+xg3R9iylee/oF2Rm4iSS13jAEYjT8scC2qsrCRtEx
5zAf60+cEm6x9HdGGUduKnYNDQ1yKYxGiIneOu6U6gnJ3aLOiz1mOP1CJdbm4Xdezpduhl3r+VyP
4VKffA1Hk/iRyN1Nput7Z6ORfhZ6SWkXk5zt5hakyOvXrYsed/hVs9XepDyK/ScXqQVbbHy2UAOR
tMwV4o7yjZB+4YWVdcUb0bosQPPVzfAaneNq1np1YCZZ8PkXrNhZH34vX+o1tneHbjdkbS6jHiE1
s8VYlKTw5uL0uLQ3GqVAAryW6EzTakdlvtnqOdIKSAa1R7C1ZIZBVTO5L6C/tZGQC46tcfhOk/xe
VkBqXwSIJborwgllEcaQ+SabVUD5L+e5+/09+TBWiZKImFC3+pqsvMpGID8h1ABP22OoJe9F5LkF
kKU/TdqmO//hjeM9O2ZzFbvhUkotMpWDq1Z96dSiLZMdlJPHFCXTlTXLE1nCUxwnFnw7kEaNoM81
7m73Uzh/2ks6bp5wMNlCc5MaDXG+MqQ6gzstope6pXSAnolV6/bjT3QAonQ0txOEVdIJrcvtcDAp
hJz2Mc2ZLGWktvxzue3wFMfdOyWVlmJAlP2lWEvaui43LV7R748giluzMxWgpCJo8gDdlSyV9XrG
dNm2aLOnYL9e2n8Yz4vm4Kdn4PNpVYujwgusK70UpImsGJ5RJx+Xo06OK1S5O12TYQUWRTZ6b1tW
by5uB/i6HiWjUUe1OHEiwMjbJrZYgn2Wfh4C3jtNYkSfU8eVq8FtndR3ANERV6N+X/+aiJJFk0FB
MAfxNMWOE98v/mKGYKzOFULjRTIIlszr52COs7C+uSRNneIM7D/xYfWor/ru9fpvOGusdX69191A
FSYfDDwAbcNfnynre8IqfYQOaD6voH/qIZWZgQgKMoW+8ALtDOYetWmTyBs7dFXTBRwBX3E3BEpY
bWVrTBBavxh33bGr4nitPyktz9GyIvzcp+nQ4io+hPyncw0U+qny2/wjZCI4D49owL7yEJHUAAb8
UhTbZVUXbuCqT4QsB3NseBz79JjX21prkVIMlOd4EVrbKlietAcGhw4MteeTHv8w7EvOxlLAoM33
95MHMcsHTz4MasdyY6gX/mHmv5NnSoKxECfagZvwld/h1jLBCnsYfASRS/Qu0otuGalnZ/IioQQL
LXty3g7I9ZiXfKaI5ArduIgjfLPcZasX7OeG8smB7LLz6qgmSHQAJ8Do4Xv9FJ0nLEkRn0/hcOxB
lz4xmAcK8kUmErNUi8LQYrXWOTyILfclkfNjYqbO4HJd60BQGF3t76DTsVQL0LMGultC7fbAABy5
tJGxJ1w9KbAJQyTdaNtYYX67KvQWUOQaor80cajVR9bzlHkzusRUDvzrCxCq6C3UxlQvisec6Fdp
W1U5FNEIydDvMWvH3RE2khPDr4h7kRbQqgxnPQxfIyp1wdQCWl7RdAbAJ7+OqB+Ot6ovVkWMMpAl
lUdZL8VT1B44Rq53qDNNE+F5/1J8LP01GDgKxNvjwVgpNSm65o9aQ9zh5BHMJHhSE3uuCixRuHWf
oZqZmNFmPt/Grg0GaZ6qxe5OnjcF/hGPuL1l8IpMZJX0CnE2jPwMZ9TApLbvofzLCT3puaYTlkg/
fTUPp/Rt3XG5YTTWzmsnDbCMKVwZQkvSTPYc/5e1loRYkiT6SYKKRZZ0Sl4suArlVfg0ovkpXG6s
dST1keF3k8NWBcJKuxT8AQWD+wgbvhBRqgJi0a5afw/d1hgBOV1l2+l/TZocDn1O1BmGlvmIS//s
PC0Mc5iTkeemzlH/+4n5nTJSj3Gt2geoEIXUp+1IGMBGki+1M8kse4fnUrgqKcELsAMh1y+4VLOt
LjXxW395j7dp/sHBe6Vefq4oXZPw1Te4LyMLuAiEMj2Z0yz14x3uBEp2vD9eJ3bwoQ5oV1kQ5byY
2UvxIc6NVDo8C0Sm68ABVo4buiAdwxaH//kUIUztbfO9Mmv4k/214TjPxZjaVIe4SdqF0henVZY2
7DpnnRxSYWlcN8pLZPwXMzgGg7TaTzeOmVDTT797p6zyQH/zPeyI8cpJ2XNQp8QtloF3448B79d1
H3HfIlyoYHJ9PdIzJTWw8hqWpi6lbGhiHEKTOMj+2JgW8uUpg8hRwOjZ/CSSjaydwTRyks3m8RHV
G4GRP1Qmj+t1+/ZDsekLPy4od0b8K0JhtItZXzEOBVSMMMcQtjQNiN30EY37jlLfRo+Wp0zfE9d4
MwoXgERGyWE7wNkY3NTS/s9VeH5EklvnnMynvg1CekudP4sL+6prVUIgg8VH/v8BMs9iMS/AJrWS
V08vyqOnvfDzUNgqYjO6mOpZ9mbNujRSJdZiHfHM29uX5ereLUGv6ND2l9qzTE7l6TX+whcB6Gb+
MQf8cdpmCwqG+qAKwjwKRqlRkl7g9CHLAmeezrZr0tLrd9EjLG4Yds9HQL+wVf/cZVAXzukn1PdT
tK7Wnd/mGEIwzQ+fM1le9L6HHGiPOfgkQpk35//DsEIR8LH6iz9GJswrd4/9PEarGueXsaQTUKNP
XCQinbF5bt7Nn+dVu6kLP1Hoyau79CLNv/74HKmnugFuAmjJjeh6ZW8nMep9vIb/ZcyH7CLxMM/N
IGCCg+SN76ULGsGrM/8hsuzY7pJi7OzI1BGExCslYy5VImsni+nhp/EvP41BiojbV0pK8D8X6UaX
WPSndcsr5WBjDsXwioyvvW0vKLs8ylCtUBEhehK1XoifN1sCsutw1Qw0k2HHg4fRxBC25b1RB3nJ
7M6FI69aic950phtpFbxXlFUnY1czYZm58I/6azzDZEjebcex3KD9DO2Nc+WWMDn+moheV+mLP6e
qtEdsERS83M7IJKuB9BObaybSzJFgSe+SlR9UtsubHz8bsDXg6jofR+KN6fqpUlJ1TlUarfu2YBE
zstZXFQdaIt5VsIEVgMB62zb7Ka8lfyBGTkfvT33w+cQb97HAsi1Ub5lfsn3BjQ/VETg2jDwYmbr
aREIcVjRg44Cu9VvXQR3flTYsJr6Xb7UP7/tGK/RXguUJz79XVhz6G8SV3h6p0eJAPYU1DAPF9LT
vZQRWlrnbyevjJXBURTYWTyn5qttLOm7gj/iFsHhiaC2Go7LF135Q++zx6Qs/NWi9Ynj8Dcae+H0
22KyFVEMmfk1Uw4OzETvu6HxoGwiSthKlkxUOsn2e07o2xffoN5LWPc2oIgiq5ZzYEWF+vcYNNpf
F0lUVFD2Hka1Bqpt9vxMHaP83JpmHdjw/34KKaGtsh+UCXmdVI1bD1ssJarXvoFAjHWzLsW0/jJ5
qJa4otfMyhMnRn2dBgmDIzyA2OdNMEFNAcZRsCdeeIn1PGCi5iGiCUoWPz4eexyiFnxgOVD0CIuB
leZ+thN2Ftuo7NeboJNGNOdnEbALrQWSkBL1mec20QGV3AfvayWYLYiwjWesLTmFOzjv7pN7SkuP
l8nFxRXX6GWJmqdJArSrCpoKA+eG1ee9pWR506L6Fqkt9xIomO/56cWx4uM3tkU1anguT41Fbf+x
YbtwzAWxwcmMQsgqOJtOPlmDN2SmeJPeqpVNSx0ls8v4zJDd9TisAGacrMiAKS7vtMc8h7ZNmdwR
1vbmlEPvCpqi/yP+0u4dSztRGPxwDU4JSqHCm4QsJoErgVNzAm5GNunzPQh1cY8rA5GGUKeXi16z
eZUXFXU0vSCS14rl6Wie8GgzlADVxhrO+knX/kyZVS7m/olYyNMIXUIDS4xm/uLjGTxp5YHB/eA8
iBh20Crz+xkaoXGyQhKRYHYRrlBs5YQe0bI9DgYS/C67XDGgBKEbcG3SwUHrDZ9kbseyCQ+H7UTx
A1tnYaO1X3THKCtazi+CORPUbyn8m480e5+NWvI4O/UmZM5ggHCH1cR6k/UFcTUXayNQD/WYpsoh
F7ka5SFxJVnZpR9E4WZBlN1TtuxfO7S4yvvtuXzpgn1+E7WOhxi2un/BzKI5hqr0qOswS8BCFMFN
o2WPFrEmq8U3cP/VN81Y5lBPokzi/vJQwQwF99OKHE7gutRuPuevabeV3B2KWFTZClg8t2kV94uJ
WpUG8gteAOW5Gs3cR0A5OgrysachIW2WDNiw3wfkVWGAVq0lDC4IrK277hy6NKRvUX2AE8BJcVgy
MqG4RwLiJ8r1yUTiRk7ZYG43YzSHInm1HfrfeH+H86SnhIswQI5FuddJsBxfyXEkCqQEKVUqrDFG
TyelVhdwqloc9izkZ4gG4SqRxGGH6yyd7kdDBFLFE/nb90ZKQ3ODCqmXjJQjKN4bwAtB2mvmqOad
J6CTXsCFGcleISIKQjKqvYIRJIh9dyXUO3TnLfyl0ke1W3APYDsyinYTiONOoN+WWL06Z33s1TPs
Hi7y+9A2UsENZPyL1mGMIW39ieSq7llMHIzgZSGmHf5VBuZ4D5oshrAReVxa4CnGfuMtbxPQ/CXv
JsCJ7FsmR26hkh9VLKF6ex6lU448E7gOYonMvpxSq8rFyJGS/RKo6BTL7nUbt7CEip5jQCGB7NS0
SGsMKUMetHxcmpt9itQM03OZBGF63mX9sXU7sn6BE9GltvtDkNOPQ+igMKiQXT+ZIPD/SzV8zjrx
ddMBp6ylaokWykneJBW1i0p7+xo5ftAHwsO6mUUP5YUT7RZRATROYk937HmQFv++1nPtGUqYrPKk
futHAMHh2LiHWM9s9QKQXd3bn92TEmJmb01TP51731wec+YS3zluWjR6K8N0SQFRUfJFbfW+o1lf
4QA/OUx5NA5LXZcP3BLUViqrJ2yJQxM6ewfoSwhefZbPpmLFPfBJd1z7+ML52JYx/I1kI8Cjurk/
pc6FtlI7vlcXF9dKuWo/apGqfL31ReehPUaNVBzNRyio7cNbmOjATihihnirjlA7NQlhI2c6kvPw
AGlXY6S3NzII38DzdyUw4Ie+EvWmPU1q9GYpO9EobngttU3iHNpd6rz+XaVoyfqYPiugU85bg5k7
B3topxPnFTMU1T4YBDfDvyK1pJlDs7TU2aZGTzrbSv7Ug0iLINUzb0pSR18Xagvj7xESSpZfrmwl
d+ov3AgO9Z5A3mbbwxAFsKAcMm0NOOr10/ia4h9+TQAVZQ3lrZfBp+maG1ROeXDxIj6CN9CvWy1c
wNdwAKINCToUgFWXmM2xKIe3oD8VpwY33km0MDdAFGZigevhr2nND3wfCbZqdj/YkRfstLWPNhxJ
DebgkaNKRw7JkT6Q2sj5pgOdGXO5taax/fVM5yIytCQfOpnTXUiRpsog7P10oR5n9LItZOnNXD5M
eKyuIXGudsL5qSMXeNwq1L+krdXkBX+WAP5fPlMDVPRuN+lMNneXz7k2+dUUXbuFsQ0QGZeRIOdE
PAbXZP8L1ed2H3Er3gcASGh5in9ZBy+YaPbJR/lMtXYl9BRjM9BWilHS7mXT8QYE2XkG5i+Rib5l
Y30YTsm/LQgL2Y7LdQZBBIDuxNAJK/mlC9Wp0Sd2VbJRYo6C4RXJ/WWA4eJZwJvelwGrr0kdcRQZ
8R1a+UNGcwQsuZHENmHPo6yA6+AJ4AD0P7uERyL5U9OKyBtErn7RS1CPlNHgtR9Y3X3bWZ/nlyM0
ZWSy+26HPOo/cAw1BfSscg3b0hRE5tQfhva1XRY7PwTSRhDgvxAz/7M43ztuqm6ShX8lVffUKjIn
Y94G1m0oTvutk+wFhiqEwhq7SF3eC4E6SZxrBcoHByKkyReKXitiPkE3LEdiwRp2p3Hd6NglPhud
JJWPaD4tzrvICfirHmsxE7wL/685AzBHkGB9xnF16xOc9eY/ZmMgRQ3x33jDEhM430XOF6ngeI2F
Mcm8DHSIw3WjSnCs/WDey/QyUd5OEbt2Gl5s6F2CDnLYNBwkKd7/T7Xgef+q7Tzc7jxM/owXH/jG
ZbJEKyYcBx/mCq30PomYr2NcoyJyFJrazjaKpbeqm3KhNlKUixfvmmY9ruDBae+yByPiQD4EaAUX
nDKXaZaDHy9LlpRy1GeYskjjAgiHprmtlQjg+3IFlS/4edv/n54KtKUwdq73qHW+NlM11EoO2O2A
KjlRzEY1dbfh31IVXPKCdJVX1fYpZnn7Uz2sNOxiJ0TlPPua/7nP332aCnOT9aihUvqAc6cDuf1D
7VZkgHJ4Xu8UdI0QXgVP1KmCJjM06+ZNJc4+HqX0MBU0ma3Q1Udg9AF7zXsm3uvZsYPL1lWgquSE
2DnwD2kNgbM3ngYUV3ZZnuaMFN5avQvrvFxFNEEPfoNDvUPi/FFPDY3qCWZQtEohh3g+u11RVSkZ
m+EH/FX+JbNIHlCHplAkk42IvHepF+lCCji+hTvOE2+e0XZtB8TiS/k1B72eBt+252Nu9rL/yc6b
JdlIR4Jc0Woi6uG3E7o+S+5YjSnXXPAPiaYe0wLFYJZCNQCqlabjeVqG7YbeYzdaSiOBFCzDAoaZ
u9Rs26Td/9mNoWZYq8Lt2YWjIH8nl6/iBM/8kybGy+PFnpBp6vnHdWHVOzAHtUW4Vf5rEfYnY+Mh
Hyypz+619a8VGnEwjNkYDAMcA06W1R1tPphy/O49Ua3zWENHJX3JIKaKaAtLJZGQgpn2N0p7pMOA
vhdpFV+Odu/FBGvGJ3qv+/wdDVmwfLff4EwVrNHut8fzuXcDCprOL+tBOnsJ8DQle9moMNeE4I2x
bZlArP2SvcLvG/qdDG157zk9fyxs7vXs1Vx2N5P6mTgjtubh8tolaM2ayZnlg2plCP3O/gget8qQ
K6UdIs0SBvk5r5/fv0m/CR4wzuv7sYuxQSOmgrxXe4qGEtPpLk4+g5WiB3Zr1IXIr9Es0Wy6aqKN
/qUfQmEHWE3zMJfbD0X+hBnf9+u4Im1Czxvs9meBiiZclpDJsiebNMqxQQTtSfAVUUZnOXYBAkDC
sQBBo0nBcYhcBu2DzfVKzGj0RN0kPgGpeZcB4hjuUXb56yOQ6BTV5Sm1exuOSV3tPShE1UUCo+TP
UyqJ1HXuv+dt3VrzGCh2fMYJTVPQwpDwS66cZodqoHt/DLOLIL2g89+GQvSUqhDN9DH8kE/pXrw7
s2uRt3LLcKndxBnWHkIsxBthCX/98w6TyqBEDRSoycJmh123HkNVUjMM105CSL0okref3FgkpiFx
S1000oQE4v0EIc2Zp6oL7fZKKU4l2EFo5etun6hoBUAG+1dSDVtB4vXqqhXX4XG0A/O3MX3EW9zW
GetLN6yb3dkY9Y2crvNZlSLjUT/PnHOxxaPZGNG6nX/IWYQ3ZpE5i3iHgnyc9QEymYgQIjs+l0S4
BGWDkrMclzlzWsmwHSQc/91xveEyx6rEk+1t5fXVfPcbgfioXeTIZLjDukM83NDBbJBbc0zxROGQ
3PaMDKG7s8iQ43VL3MElQSLPKSmAzodByIHihaLhCHE+tQjzV7r7IQXF/xw163UpbPpkLRKW+aML
yDYcuS4RZenYVmOsuU6Rn1QdaGlf/7j5qZ8d01popTXadiK16w2CVCFAjVkdkKOCR7nocJMAjsGg
VpKTAgAGiVqBSEbR9XR1byoVTQhHF6k1wENrhTMf7m8sz2IbwZMUx2mMoLdNZXN+Hz4VEaxNj1fk
CzmQVHeWS/ip9+WYlT8cTSJigRgBbMkjSpCiHv+Vz1ypaB107YMT1oou4yheo49NTk8zkVlXcckZ
dueG/JBt+Ss/Zt4SDXz1NB1UGEtLEpXnfICVDXOTUFdbH8Y2XIedgAL/EhgH7Q+n5Vv+t0gL0BiN
Al8DO2eSxKQch/ha7sFKVB7W8sLo2wgBvUaZA+vKbs3O90HoLJDIWKMRcw5VKAfWjZ9Grt4QreI/
47ZLZVwjlD7Sa1p3VboysgO/PzG6Nhtxsu5tjLPZWbYIo9CsK7iYBPikmsi9CDrZPymkHudu4njs
Z9ygvC7AiQ+AmNTwWYivjmqW5FCoOkiMoQAG2tSy1jT6o9gMGQ6P1ledVnPU/pZz68KY1KWSAwzo
nQeWJ232lIOkWXBza0FzdYSHNoVYyHpwSYEEWZktF/FjbJUAVU1FGxvJ5qO1QWvvKGHVrSUD3wkY
foZZZLd3NKOj4xvknoq9Y/u6oIcgjyrEjcE6cczgPeZ3CwVOfMPqvo7Euelrw1l4zWOJuyxhdgLY
CVJsptCjdhBb+03vgqo7UvmNENdYc/PBGUf58Tc5F/GpJ4OunSDRSBzEt8ImWJmioJuKIlR1uWrG
W/E3ZXanGyGZ2PegOcdkvPPg3PTXahFxfaS/o4Qwua/ZoCaXY03w7bgGubB9NDFASLSGzLDpO4AE
gnL3JA/GItOU9JO1B+xcUZFmTrTqoeOXaKJJEDIXRUntAtroghNOMop27f7IadkSYbFMCpEqkSsy
mkRAEjFI+BgIdPii699onP0afmJv4QDTj7A7Ycs71vXtsOYGfvI3OdSxk6TkEbAZAooNucmxAHEg
mE45ZstCGWbAlX4a8be9DYeJtFIZKqaU4HPFE4oUWcswiaJG05qwJyumlVL2TdPvfe38AblT0Cn8
p1y86zCMV6pcoIit3mT53Z0xinu7gTNzKaR22opOm2ehGDVbUCHeb3fONNEQ7hmL23fjlk6dEPHD
Fm52PGZN9GwV5U/v3+MsQZzjlk7fDsIzj0QdILbkj9oyVFIoaSysKgdkr9QKvO0bWtEgc9/L38rH
gIdeq8JHEMQQo55XEBpbIdYbxr0wyGSRrUsM9r1Rulz/sVTpDdcLBcfBSs2PuoNN2IJHqa7to7KW
NGeEeXN8iDwcQjYHK9V9z/vYNxrNI7WJBOZzG8UCGkKinLAR7DIeunKWv+fz7nN7jf33vwN4TPhC
9CBldKCjHG5vg2hh98NuiGv6P1z4Jo6nO+/QaTRiHZqqa5F4raNbxdmVNThVx2jGrSkHtv4eKFlO
jeAeo9HsW/mqQ7jjcBs1tU7OwxLlSrG0m8LebvbX2DwYVp++8SWZdCIGTHEjlMbVOidug/i8Wc9v
xxJR8QsHqiqA10fcqPU6VbD9dENuKl3J2DKMtnkep7+PhTVZeQvrhWnwCARbRdStaSDM8R6ZzF4m
kdnKKtAaXfuL2Yveu0AurvvSqn3PMxIACvO4o1e1Vmbit3QRiiy9vB9A0UNiUTbJTO0e80GxQI5W
ULug0IsSn1SKvHD5bossIXwsAaHinyJQYyiVTJSwgOn03bvFtqTVpPxf9yys9hZ6dHs6Vyfb8V7/
4zUmPwTak46YbAoVlOrshTgGei17aXDVi8tij3CTzulXgHtsO0Q1e0cdt5BRZENjTkbShuAaIIjO
amWVb/u7im3yrf1mH+mBhFtv7hTwQAF3ocIyrH3V1J2a3l2VIPpaC+DRffeyzl/pJ21ccB7bzzx/
SyijSqQ3+LdOI64Oo+G6qhbQ6gMsSdzrJf3isJ0y75NwJfghk1ZSEkyYvuCcgo/ysi8cL4eUwj4o
fBaV2IWNyr6R2Uh8eDSG8tNNQh4F+F3d4EYvWSV/L0PEgq2m2kkReenk8oBS100OvFOmMgJuL2Fx
WFa1+vb0mFQusCVxbOHK6mWSgrhH7i6f4GUc+AGcalmALOvj4bjMyoe9hkAn07e1DZC5zmdbmZV1
n2Qs2hRsND6XZmrc0tAhx9YAifVOIaB/pKi7xU33EhdNA8S4bDC4oBmmnTunPwNuehr+6Blob/13
sOiBiWcYT57RDXW4i+23kOHOEFwpH88VppftiEOu1GWjNBZjMRdduR36NnBR4+CqcCPqlqJ5mumD
w40/9b5csjZ3/9GTz+jjuoWm506l07bywGMSlresww/sLTkOxao9cJ3ZbvMi2iBzU3r56je/Zhk7
7NRUhRXhrBAOanc+wmwlAN4Lqd6yzUfl7qLQ10I//b70+5RS/jzR6F0Y8CDtAkV0+nBdLZ5AmBC1
6nKAFejIkK77zs3ru6Dy/cMTqByupawie43o6ozydFnlmQUSr/QnssjRE3OF5++8XY3KJjfhU6ve
JCRvkKl8l2HzvQJPBH19XSCfDrjam4fNflR+UZr/nMtyOyN+4BLLTFB+TwO38YhhKppkk/gOIGPy
GH6JroZO40mabZj9FpG5NNuu8BVX5M6/KAz5iM9ErFS+0agjDJGydjyBfFlX7vG0v2b+KVJbnB/E
yGfF7nHB4cGXtGKHc7hExFsgVuObydyn6vOFkOj9uE0rJixIV7M+SEZxJLu+LACO67Z4HngPxlN6
iNndYk7dYLyCXUeo5xPvE0DHhUpU7hIDhu1Aj0H8+MrdaLRnMyjsB9KwtKgS+K3GSsreCPchICId
Xfp1wuxVFrzpBDSvCvBQwgTbtKzrmVYmYPXpZgV2FJLZ6kDCK4FbIKIP/sbczycn0zLRssFLlYdt
qPMPSI0fDe47TDgnJa4LMETK6DlFUn6S3f/c3NrhhgJ4ZX2vUxxxOjG5X4j0gtm/sLOaqkD5g/EK
3T2dYO/BmJRNW/lUaleI1U87uc74cWlfO0coGMTklz052IztiUaq5C2Aa/f0x7Wv0rH9X6zHEfcM
AwnOVyxY9Pzg3xSjB/znqpGISwWRwtzPF6LbU2EPcm7Gw30Kw8ZPvn3WAHckk3ddCAuREhfkwS2G
WJxdMwNEaZq/sHaYMaXfxKPUiZsZ22ZU8ZgPazEB0bFXuke49UxuVTFjWL/k1BMaw5l5XyCEt+iu
5n9y0bRwABhacS/74o7Mc9RtySwOcJEB01lbHtcncyWrihEws0SdoO3L7lAzOAO9g3GIB01COth1
yPHwJgbokJsj9Ram3KHn1DPan4WZ/LDhrE9SyavkZVJYi1a3EbcUyGsEuXRDEVca43qGqBa+KoGf
zZZY/IUP/TYjxHOmwazeyBn8xiCrB8N3Nc5Hju1YCH3hd90/ki28CM9SeJfZkd5BCdm5yD0cM4Ed
JLgwphiotA4NAPhM/NWH8ieGww/oeskDpoyddzzAw70+ij8Uhl4B1FsfFIO8wXzA2uqH/xEYBV8h
zSwETTjiYDQDdTWE64t6im5ezvdRhamOp/NGBVcXBjWfN89vqeCwIcteRKHC0oVXAHy1XBom/aYw
zzYQ6Q1in+OWSPWl73OvfXprjLtVC/IJjT+oJaYG4ELU92g2ojHEzXwJZTO8+MFwW7b4hT9MOkHp
/iJj0AZcr688I9M1E/uNrQV2q0BdaySSxoGHPYl5VX0PDyRVkHuF9QM7UVRh3h6emsDe5sicwOEJ
19CJ7phvAy6TuxHGts3FvVhOyaXj6/5LQGWGJwHOTnah4XZzr6T9OMT5eITn3WVZLzAyr/lX7GyI
B298/LKPKWcugxcGkW4E6T0chJnkrC2yzuqKrf9EGUkFq2OGZRVUHcRmnPvlBadqMBVeXZ4WPN4V
hWIgcg6paoHOEktbbh/S6uGyXpoUZL7w8N+REnU9msD6mtyeSFj8OmW7whZS4i9pLpYheH4nUqmG
zfFY1LJcmMV2jdlymhjP37b+BNL/TD6Y8RvLGvDtwoOYqoZYGDh6mWBY69Ld7INrzgZ2Zto4duQU
3OFqojX55fWPhLIFo/R754CvVwyGUD7iv1Blmn921jKeyLpUzxazJsumUxtuK7yFLheDybNkpu3+
qiuvvaNDbQ4O8xvszHZcbC98hMHps5xvUtVdX7v+9o7sieF6o6xEbkfwLTTXZ7ld/lepOhFWXoYs
GZ6qboQsTjjNdbMKlSANnOtDIisHr5ET0H7nKRppm3pDljsFX8LWKAxqc5oLCv74LlBYiv6xMW70
qd3n69aVOh+ZJ4uZF38hCfR2zdbKWLeXNLCB3RLZpbk1lw5oY6PkXO8G/l45M+uXTAmH+OHfuhLj
SvG51oBvF5OmlHtLKm1s8IVfBpD7FRV/kYtFYxNahRBdFhuyyda28illYO4xgSvF/KEDTao35cis
NZyudC/MzDePcFsklwFaGjtNQSR8AwIxzNlSa+QJHh2uI6bmCin3dbOCwbPU2ZW8MExKeOb1ZoPc
lcWs3u4cPwer2dVmE/vbg3HxXJgRoTlUzjakqjiA7MaSDUC6Sb3KIxbJkDh2vqyw2+YN0Fx1xOdR
U6pbweTxd4WQdy6ytal30Dlb9AJAwxaMy/lzHI3YYWjTlZJVLVdC7t4lP2N1ka63YZfRTZXCxEII
T/8D3//HjQB2z5uodPRNilAhOvL+N0OmSu2XIASorXUw81ykCrK6Oq8W9EMWT/XwdbZ+mr8ZQqKq
rcnAsTSKyggB/e69urfpv3gnOelFllQKEcH5+tJ7CcpWdcRxcNeu5cqH4snSjE3tg/bqqfclcloo
CEhyrvwyqrCcA7C+wkp4Q+u1VenN6uodM/oOJsdyRxRNl3uEvYFe8erRSq8XAPNZdmAUO+Og5FbI
e0QArnKGIBEJ7q1P+6mDjQ8zl+Lzk7y6eO9gtA7JwhIqNJuyplt69vcbivWcLe0kw2AeU9Rjzb0K
rPGcDyRUetJc5jy2ZvO9N50M7xy8OBmS0/CNe4/XlKr9J2MT62n9/C1jc1dvl66LmS5nKfs7t6nW
v9CR687c6OoWs83n5OSNe7RyvaA0BaRG88GtbeFfc/0g7pKBVjwv5i8k1moWvgqaO1LZnIf5GVIL
0HZWz8Mfmk4RDtGB+lfwC+X/Nb4P9QauKHXT/+bHLgsDdY71XPunF0sAQUPZA4Mnh4amS+DXD9mW
RWukW68WsCeDCNxDOBFSwf4iMof2G8vzzbq/HRQqOOqs7OvKwb9V4+Dx7ceWNYwstgoVqHA/QhJ6
jfTqdLaJAo6aZ3m9QhXMsTWJUPQq/xpx5Ki67oDS8AtWUlv8w27cxbg5UqJh/I/JfIYxbYLoJB8z
813h9XlTmY8lI+HKBq5+12yC7dZTGrDovhKyl8t4fRst90kCQJnki1klWMZdMO3S6sOyPHpO2q+R
Zc0ixtmhB3C3dQAbOBPk3oVda4M0/89WFj9YjgwlXQ3S36QqcWDxMbPQIzVh6sggHCkF+qS4Ggs6
rGrw0zLw4HrmGegYo0J60zaKHiwD1k7WjBpT1Lt/gulfQQ0X2T6Zkm1YIQSXzTCPNia05TQo8OI7
A+5BdKMysQZ5Tyro6ZhmEqXBsEskUsQEGmon9QJZVmMwvsETbVBF9GbnTNTiGzdQFueFmZSnZGXl
/W666ldWEa8XKQp8rIccI5htdBKa+W7FYlZP0Y5wI7BWRbP17OTT8ZR3MuYJf1gL4sNcfQveqkXY
NlCBzMUVmDpHu+xYUNlQuyPu6SAU1lR6kc4RNMGBVygkSMloGr/agIKca2Put3lCuVgEVLdz6h2b
5awe/NKoiqmV2daKeRRyz9UfU313a4PHfOuBlcIeiTRcwnE8oEJJcOmoDC7FzC9kMi7H0ESvCUOj
iedNPRs/zbtaadaUWRN1CeoJuy/kKTfzrXoukrSRs1OgOPySLzrnW4ma49dRaMOo3UwFp8HaXKYR
3y8O+DEsip7/7lnV6eqwCcZ/XZlWZHy5FF1/3CZmmM7TmAkNFGv0KcWIvFJXYlunn9i22vJSkpTd
aq9kRGe+AlKIBEnsO73vmEo457Q1I2VdGxIib9hQ5ZgKNuyKioRkouGuLlxRooorq9AmQ3+97zyR
ad1ZDOqQ5dVPTwoRR8FNdI78dR9E1odvLXRqOnUeUne0X3ipUdAF6pKXwb0bRH3bavhakrw0tVyr
5f2KHV/G2ykyZ2Q2QjsLiIMInNgbRiKK76YZJA52T2qPefUlkOVf3faEIKYXZBFJz0dJQAWh9zax
gtVoBr9DGOEIbE4AIkJzcWorivHgIauT37UPpuQmD/m65o2XN+TD/lMU4JuIxLFld0O+rNwhzc+E
wE33y16yo8/7crHpdo+/pDTJSNq2L/TDkm3EHtI7iGseVPHFaNV6lcr99kzhExzWOeR04/R9w3ID
6LWT/Nm+32PdeGyXhABb1Ufy8VcqrPDv/AoRxejSnCnXjJH1lupY8Z6xaEEroV9jWH5LcGIziF1B
mpjoLPjkOFiGxBwN6S6b0Cad1QECdJD5AVl0vnrFaE8qbRBaurOxbwOISEmK9BvZXDhZSYCNmudk
5b4ciiMaqtr1lhRKXKc7bla/3H05zEpCjmUA/D/CfY0wklbJS2AAQSe3f/y7Fg68MewARETI58EI
m1F6F/ztkc4wA7RlpnB3IMXPBDE+xHM84JOfe/FX9Qs7nQdbIwSkFBlDWVr5GrIPGYUrCmsZiLgn
mWKuz4vZlDhelZUFaJV6q77QOukkq1FHCceee1XcoYEDk0L2O6himowTuF4YidfIDUNXuAlnucKD
5m+c/2z5OwoPYmtuaMb9d7avx+nfskzyXPnegyDyXn+W5nWmRNPsVQk6OrAeVZ6Q7HHgxlUGRzuw
YyPBvcqj30FfknK/FuVYi8p49MCHioTRBziadWybVIfY0iLNV93hNjg9R5KDSOzvfI3q7Et31kFD
Hz9apO6d9W6vOOO7EjZW209VtRQpGBnh6yh/7FmXPa1UkQO7b0bHQ1PbaOhNOwyr1QerARFCXgGg
yAUqJ/DZYcXhykTfKDEW+CV9hx4Xj372segj0KmIXveteUvSwQPE4bUBJ/qA6ijdSTmiqW610zBX
H7H7H+5nRcWBQSm9+EKvPO3I9QdNO8vdxXNCDj7BPKM3v9fpRu+1q/lKpvutNGrXMPsE3ZOgnfS/
oce3UdCoMjmR1Q/NwhBJEaha9kwh6ch8iaiXzYeyok1EUcljZvjA6VfawALqZPuePZdNnWZGX7+H
+/Tbivx8Ev/Jo88c4AyRxEEG9dXNzXQfqbVYn8XdzOx/vOwpxhXK+67nOMLsPDYJOaRNiA1tDhJu
j8yfWgNJb4B7uoxrVw57dFrj1D0Y4K/IKS7+mveVp/iWKjoMaD6NI1LklXgfy5HUZqK0qBh4WmIu
5Hg38fYidMP+Rah6JXuNbobBtQFa3GO78TfDZ7HtS10fExxVRRk176CN1bF/c/XP166JTd20Bhr3
4Jo9XX+Cc0NL8qLoIrzM4CPLEGtW1Ajmpk+PM4UqTbE77/JnK8nToTGoGheHvo43a0TN7iLqXVJE
2ipgyXUDKX+mLn/PRRm8PNuTZlS+Grx7z8o4w4epaHP1UcdLS4sthw5GpoqFTVwisWzNImBf9v0P
cK9qhli/hvFULSTcDBCdlmTeN9GHN+BMTIWK6/jLqpkC/dOC9/sc8DlNSQlxrAxLQSMLFHr4yiJj
6YqwtdDKryNzc/vpfSYiYEk4Bq1ms9Yf8PjNHg2o5tovmOumRVD0w1gfP5tIAd23Hq0XVzcCwNVV
19IMORRsGz95L7BKsV/cvqg/QUPo3/tkGo5AHnFGI1pyeuaTcoOOVWdVZcI1XdwA2s9bTkfbeEGN
9/7MI7EOIGakzroxHo3xDPBg86Bkfo1+nIS6elSlc6lDxIULZ6B+yk2EZ1BP/ZYyRDRy+/SvEfIO
eou4iuwj+CSRv0s4mWugnIzh3LeukMOmDWsHenvXnB8BrsqAZMd7yIrQPUcAaIfiYCL9dEFYYhRJ
/DbbSS5O5lznwwBKiA+WnDpQcFBKChAmWO7G6oYwQdeQazZZZqQwNtY6Xi2NR/funvN3xw01NHhS
HIinzJGVRsURZFqwxlLHdia5UcUHAMxtM9OtAX/UImeT3eXo3PDQz/rtTor9/ouSvBN0TEiI9+nX
k0Qs042CHRHdPMZd3ZiiFITbxn7j4mE5wYIn88jkHzVJrBA9W8N8+F6XXgjW0mQtgVZiPi22TtlM
9O7OmIiWUpzvIYek0RHaoCl2HvXtttZFBS//a9I16jBa0/yLK5QYaYHpipMvuwH5THJv6N3g1M/u
Ee75eeuVYJVKnhj7AGqn4oNJXb8E7ZOFhZixjWOnzlZEa6QXnW4v3nlWnh9JI0BqZM2cw5CX74cC
G4bp+6P3SP7PRws1J6ENDrBVW5il8aaHs2q/hjz3PJLCASDFvdKjzVi5AHH2pLUUMYR+lotYswdf
98TBECpWKOVSvC2CZD8FL1g6upNlVlSOAjmsPA0WyxuzsnvndYwSbhE4CLR9Z8XyojDRwOf5X+DJ
XESb1CmASpUOQdBSbX1IDJkOiwt/desac5oRFCdOddX8gO6ISWHPSsCfGfduxD2YDlP+gGaPh1OV
3+sIEobHPAsrDqaOi7QhBkaGcUzrh7kPYBV4zG29hqUhjT5TDERDzLQYZ3X1buYZDjHohFq4Amjr
2tw/V33vNe7CnBW1GOCEg5s5dr3hkkKa/XqfQQOtCEV5Dl/1AMzqng4bD9B+8yl/qiJFs+jH6vNB
k9sdB+2vbXof99dGlwfPpyL85Z/3FIUJeB+tKdEe2cjWgTr1Bc9x0ZzdKudrKXw7dugquaj79bOl
i4CoVcr3h20dU2ka/IA7tzNkL1Atn+kF37v2BR0O70p8lI7AKfA4kRl3cyUkm+jaPK6yhOsGI4hO
lKwQTVMH1TNK16kZYXfTnsmon4v6yacuuS7Wwn+e+9g2SjGnesIRuI+EEtIMEWAWgZK3PolfiisF
Wr2zrBzE1tfsHID7Co1WkhTlAypY/txrR4gZczF2Z5z8WDTlgapmK+FDH+nSGaC7CC5QJPyN0luM
a2FYXtMJlY7Y3r3JCsrIGMv8d72UL1YNbqwJhTelaqX/8/IykjHyVnN4l6TvSWL56G7CD+fuj7jZ
Py5Uq9qSz/kuh6EpU2cGCx3jOtZNq4/3XdzNpDHLkoDb9+8rG9B5CdtPAfrMvfpsFK/AVDut+EjF
D8P64AUm8QcumpEAhbOu3lR0AqDMfDlWooriKAmsqP4cOJ1tmDOmZH6ckRnbsy/fExrx5d40aXsz
n3GV7gZkwvw3HFbjcG12QKOQamd5Oeqm5ig4K5hecWlY33OgtaJ+EREUwNPRNqLjXpG304bEHl4k
ejncYq6HeCIbzLDsDE/+vCJF+BuY/2iOxa/4h4p9PEdGva3/HIWMITb5NerbPF24DExP95ntlnr3
ynXi4/em0UbE6lRLy5anzY6XC4mxjauQMnf9leK+HygY1lURJhaIS5dOeSVtHZAHknIPY6tJotjO
DiLcxF9QYV7xF+0WVSyKCi/+lyjurqLT+wI6EyDLPNWGW5E8YsNhV0TgG2verkYRmkMMRXSvu0d/
KBNRi82RgeXdX9R0FiV7lSpfXc6Ec6Kvgtq+h6sMXkCKnCa5ISNNXoMHrgmBHl5xleWwFsMVoeGD
caaVMTkNeVtLVEzxePUzGYAFmTshc1KFoGIDNxifg2G5H/qFWZlGZnNGtnQHxIuTDTpAICdUyecb
NU1gCzy8IRG+3XZC2X4fsxZDidfeDxk4WfBVqpN+gM1T94Wf9sTeJX2WwQYy9BsjGmQYu5qwWJ3l
VWGGH+xjh1xTWm7OE2Jo1gvcEvvXRlKIXB3EAZ9yMt3YrdithBpvZvLEOm98IkL04qPIWwvz6QV9
ztwtxkHfIiWmDMzzIjFFAWnIfjIwRBX5YjmYGDq0keDbjH6nd8WsCvkQvKIhf2haaPOVX1IQYxFn
cplR6g4virhxS8en5LpZAa6vj1hzZVqlinMbaQHUmv3NvrGtmCA+q8yKHtgf2R0qcsyQAuX8qw7p
C7FdtwtT7BWFNfr7ubg0iGImSM6nfeFTbo3UrdvUJPtf99Slbp6aHlMQiwXLZ9LfeKftnxsvQnfd
P2gM35b8cs6PO1TZq3IgZ40c/awdzQULnjLcxnx+pCPtqn4xmPOrYc54JGfVJX1NKnVgKojpUO6V
dZlH8HVmXydsk85yG7TKWD1Io3cfczaX8LPKu5Wlba3o28shVC8UP7duwiDckotU6W9cQxl5aAyb
Darj+NZ4uF0I/FnT5U9UiXtFsiIVtwTJS3PSQWI0sc8Nvf4473izWkMlNmJJ1NojMSJHvseF/pWG
powdGBVUElk/gkRqpPpzot7g/G4FjzeOuaqcszxJf2ua05vKqhT7GgHM/mH3PNtceJPy4sJqQvW/
0LlacdodoaFf5p3Az5B8g1OCrb4r+EgS4REaYDPpzi3vFuU3T7Hs++XP8oL6qmexFleeqtt5SiEp
djmx1wGTuy7Jo8zYlIR4FHBtG9lMZwuXCmO8SWTE47hj3Nn1Eh5b29j9XCQRjC+ItJeMx//QCKT/
7vnL99/v8HSbx05oFZEI1tgsoGqB8aitLS/jXhaXGid9n5/qoaawIIG3QElJ9v/7kcXMrk6k7C/G
shxu5lZLPF1h29Fim1UAjMxDV+CEyrEyjoub1UBxVPPKZVAaMW8Fm2s6dAHTf5hFmwvnQn6Mf9S1
WbdectTdSVvt3HSWejDLDuBscWzMC0IEcY4FYnc6Kz2qS1/GWEiEtHqEIoFhBnATT32rC8OEaOYA
rTVw2MAJBPvdtHpl9VOmkQTCjAuKdpzta4OPT1sc6rnYrBhTv6+7L6Q2fxq5itlrVcaO+enWN9wP
Fu8tklC+ZG4QknWxLpd5il6QzUK2Nwm1fd7eGegLEmvrvaKpzq3m00UxIVdca2QZHZ0WVb10g5vl
EQB4MUB3uDRQJeuAul1RQVMdj9CeoINTrG+eAroqRDmhzfQu11whSy+91ZRvdDmqwLIZh7RsljbO
mvfDEBTSgga71F74NLpd0JAr0J6cG9O3UhCThE9qvI87dRl5GeoPVzfue5uUnQ4zhkiEyMyUlzLf
+/VLV76j4lNVM6jRMPJmoIXMtDW1I8CXYNwkwhMue7VLt5xsW5Ip1FuZNGf268EpGf+jk9Ai65hL
9+5gawkxr7WrEgbs6esG+ua0tTJzW7YXj7s93DMaS/cAuseYyN6p02N81cqWR2X7MrpnjmZ3KtIL
OdaIeZd7Tg4a01ZA7XrzTLaKhLi4Nwxkyj8HuATVSsSY/v/5fiTvo5qLgZ75LchmKs8Dlo25Q0YT
M8d8G5kJBGTmV5rZtpt34GJVTZdI9vaGxYDgDeNUO6eQ1n07c6o8Y7kg8d2oMBGnYCwzOPIPLDNu
wZy1ERDejmh8tUqxirTKhJ8NXkWeIbKp3pvFpDLxTg34h57B6N7tXpp/yAHt3SgWiqFAI3pXfUeE
qgtIIwdr6+UNJSEqPm758EXiNEeLEmcgfZ0E6FpgDxitNC1v+ChfrV8MzWhUJALlCPkrUu+Pjtyu
rs30K8tp6HrH9ssCY6i79xED+21SgKZ1uGFsJN7IrMfHJ3hQdCEm8byx0ztfdcSb71XQDQFyyTIh
CQZNSUVN18xd/0PHgqgr8JgkbCxC6tG9Gy/Sr7evXNYgFYMi9uFtpzreUc5gIZ7qNRQkFT4qcDV+
Kjq5nwWFL0ivRPxradTtzgWYNh/l3aiYQ51FBqQI8GT8eWYHupSBMOp29rjCU0WDBLo3GNU6o4b6
SFvjiOE7X7JlgLJkfwI33F0bPYboVHasP8uuFJaqrg5oYnUofMaloFx8ZzY7hJPiSHSZ0/KNwSeI
ZPCXcmGfHWjGkbcl2pJO3DzzcIaj+ew2DckGqEgB9PENWzIJwAydZOukj6RX6aMb9danPRkr8ofa
NFcClu5vxgZd5NZZyN2prJvu/Oo8Dcv8WRyLe5GIvYlOYrMRgaSDdOZS5+FeLQqB4XW1kT4BRmT+
kdVlY58oY3TBAFri5TvVTo+IhU2zc0pohPHDLN19jSp76NjYC1z32cWMzIBmxnCsMgEFr7z5wyoX
Ifce631xsFtgxGKcdiZsu6SEOh3sItlLIzjFQv/dI3x9qhE8RiJnliPAgR3W0x3fpEREX9NdKvNA
FWej4AF9OilLHeGeTKK/txKCl2qdkBJWYmlM0ZV1a1XMb23faZ53JBD/d6mwtJmNXu/e79rE2aUf
0ShTaXd7x0DdfQqvucJQqHWp4JfwCgcAWFwyonfR8mMy7Pwm6qAvHolXbdT6gAD1xYGk0LUPixTN
oVXbpLco6drORzvi4N/WoZdOqpmYLj5YAwkA8DP+gjCJYpY6GIP56rCvIpeLJZfplZ8RyHxBlYcG
ZpzaCsOIBF2YnwXJMvn8tJk51zqP5wK86e4MROpsD90QPjrVL7N5wIkxWZF8dZ6mcHckp/6rmlgJ
lYRSu/uCano3nSYjazVUVSZftYJrHfOjnj7RGQA1EMX/Zkh/cw6PcNPkBBdfQGy/KJBlqeF9TvDP
5++O50bdwJ5FFOcnxTFns+rSSmydQXEYPlxFEZ13fCeFFa5I755GPHFu+7YaNwzdQZCnIKPvqOcC
kucc5h4CuzdnLPni8ubU+eNb4mJt3oxeEPmZLZUDV08eP1nk7gqU1FPk5sB4SRybM65I+Vlnk2y6
u8EDFF3BqUZV/Lc3RPQqzfK2EY0rFT7b5S4JXfKTGlV+fHNo4HO0sBhLPb3BZEiAx38MDgbe94xK
m1lTLsJwSzj4gpdSAtGPiAcJ1P5Qyw8gwGVVA9EK8oBTnlCkPLMb8YejJjiMWR1svrYgkv/ao6uA
V+m1i2MOc8enqSYhpwmvixpiurmTMXZDF9BmlJP5YQQ2UKo7+5QQ7ewBiIYQGKWYR44UTnz543uV
Ol1/bkBwW3Vet9UwGl4GUc1XqtQ6M6FnEJztnb6kvilJqw2Q5u1HJyd3GFDd4D7157dTEiBD9k3D
ukJY2lZGkWQNH0+0L5OJj/qEdB3fDfoCWvjLnqORO9EBQICRvUy7hDxCkBz8uH9MyHTr250hQ/d4
chkpfM0jWCXm591HQUiQ8gnMSk7i9x+FbYy/Jbvg/f/czvy59TaGhv2g9IfFv4304exH4aYEwv6N
0DIujZirDyJxOLWvPVDdSRYVonQz7uftmRkb/qLm4xn9Wc+ZGozrF2S/5LM4JeSHmzfBn8+w2J6s
TCnzPiEGbQG1KKl0xnZk7Rya/ePHLS7mJjQJ1K6L/4GJKF0tF6t9W80vYcj38GTs4hLUHIA5wYZ2
NTG55aUaqxrcq5YxSX1w9/1nn42yLAZvXsWmPHa/hN+pRDcc59kz2n3PAb9GdT5sRYFzLjvgyaFk
5T8gZGGr+QklsaXgaNNOMTfFUJXdy75v8dJ0y5t27Bwf8jhTjjRYpfh2YMBU44Cvz8i8EVVUe5hi
kHIgFvt4/cIBQgmNo912E+9tV9u3fVWA92sEDNFiCeocBLPi2ACmrmkCiBNFfkMOhq6Kh9XZtf5S
0crUNShTwXVS7rtZ/GCqiGMulMiwcq+Ex5dM+Mz/IRdoWlScPC0ntyqdspzGOzR8as+GJSNK424i
cN+a7pZOXrbDCv1ee6V83FI5b0L/6ScTCnrV1afsGK7cf7wScJsmOyIuD7jkGyS93winrm4JqlQB
dCP+jFmKw2gZgM/gdP6kyNMxA8HAQGmBxp9oEOnKJeqWsFpwd/YwtuOwSs0pB7rYQ4OyTkhXLzNs
3Go0p6nJyJKG6W7+nvlzunSnM7QSrsu6vqVc+fDLm9wHvlMZf8q6mqgIo+N+FXJdAKEd+UZz8dTV
37uF3y4pGZS7zZR1q5fF3UVk2UUEWxERixcqHGcld0iHIzcZHug86OPNYOHOqxV8NUxjvEInLman
3pYWEjhxfxpudpQG6auRexShedCBAkcUKk8m80YV4w60ppLbanp+FpRZVUdNEvIK/HtBmcaKot0K
mF4E1riUtSew7K3rqF4SkIlPq10Hxo4YvRniTIvmLNo5AlVQXGehC3/RamwuEfyTbOGRJTJ2l+Eo
Y1Ze1VTD08xI7D4+aMJoqCtiY+EztXCc6lGcu/X0EMlKb977bqoy3IivXMUJo4jrz0CjWfFzr+tr
1Cn8UfeTP577cdw9upeLV6DuIxsmfEzniy3/dpCyXIl5JLZVvPYbeMMd/05OKbXzKxzTIQfqxvPZ
qAkE8WByPy9DIGmgZQou8+7H0p+Bf7UQoN6sMNFvDqRadR4pklvz17hD46X5gQejmZWMWqNXwHJ0
8RRE1Zpor3tR9rhOGg05IDiYhBJk8oJ9lYxaA/VxtTLDZYqYy5WMzYof6etzTwYO28gc/k8N91uc
6n6Hd8UuNqH/V1Ae2fd1ftPpfCyc+xqK18PHeGmfySf8SYBwsLs7gidp30wG8OzUop2UbTi4mf9Z
plX8YJOwtiqhsIcY6inBv8qnTju0vyMHEfplm9H1AwQxQCzjw0DZK3CZcPLQrIRcEOr0HjgIFBzt
kysKfJRhUbZClMec9dckCxabv+OlBwFHcI8MTDf1np2IrpTGs/YumyDHpsDgjnskjd4U12ARGdQs
jXDAj/8OCuL9OVwhtW7gHpIajOTBqWtFX7zGJtZvkeXY/uyxSMKx+2xtbfYZuKhR7Mb27Ug68eEU
aeGMl8TkeYj8ewCLJYUV/TtlOqo9iTEELGbgdWItZKeAPGA5/uzKOTXx4NX9eLBlVOb1ibd+Sinl
trZ96mQ/SXo1y8UZh68hKMhLmpALOY4UqTGuZEchJusswuJon13NYvZXlTbBm9a1p/YibhYMpkEY
xj4ZbcshYW73F8Kp/e+cct+bMz6JOGHUPFOz99lXjXbG4sAyIONo5cY0rQnFpB0zKD83evyLFs1M
J5Vl/TiRuI0vzTVMqh9ycCskIloXN9IaiMedkL4S3uM/+na0THIWUQvg7qWZkUijhzXnAvspGqxF
Vdgh5ez+jhEY72ZptrOgl+fAS4WJWmLZZ+5gQVeXZjj8Y4bFikfaI3bC5zXuMUR/2AX6LMnsVug5
ZaIz+KBPtGgMkX7/++F+VvMqQi0x1g7yBn4f9li+CabLA1d1HLTGvy19PS9B6igh6Ueo6+dyClka
/ioi4mNUJ+dC2Znvzy8gd4rbeOtwQ1cV8xmf9LH39Iq2uB8GHDyfjEi5HcHenTA6gogREUpF8oJX
mlKDUXxTWbKDpWrFlGSV1YpSoNrkgpZtLG5OU4YgBuczutT2vkGYo+fIXtaavNbrssBT8i+lesWp
bnbMLGxXylLcPR0cKu6LScu/lkMOIhBk+FlM1UPeSEIhKCVCuVNUXXvVLfk0cd5G8fPQfkeOzlz/
lfzMIdGMLIyNKbZQSFyhtSVUwSUkBt0gXf2oVRbHNRl+uSBIuuBrTAq0Z6t6PONQ/Vq1vhRdy8qQ
KLBT804dqy8YkJk8wUpetTrEal1s6eTWsej3HyGD2k47+HspavpyfqhBSs3D0LIErFtIif5XfxxV
E7UoZLvIv7VuPFbpwBNsrezOHQAy/k010hFwg9DJu9arfZL19yidnGRG2q+3qDvV66Jlm6dOYQG1
S2vRcfPSMkg5tvY59PCT6AhUzyYjROt0Vr7n4b57iFC9//hvlC+ZAqH6/sUUcoaNb2LAoe13L/aN
KV/vr1ilsghfYSIB315Ah2UW1/iuHsKpccAQLSzVP5CSRITA6dIiCrwFxkSP4hNrOJOca7XKUS/w
puecG4VPwaXsAG2ifPwPMIptIWXAWzXd2Si2y1MBFQBwU6YF7tvKlsXGit2uPCOxkDuQvXOP/cm+
ualrAMPFizrMsngjwKOc4hgR+E8FEzKffPKK7Xa4Do6lMWXQ7G+N7tzhvOjss2sfwfSMTjlkeZ03
uQvBiaTWlGzhS01CJRE2j0vkasdisioMXrGur1dAAzRzwQEjBH7dozNHzTBO5zSMhKqlG5s9KZq5
zJQX7LIQ0VmrFkMB0/zam222qyGwos5+L1Hu01Yf6QJ3deiN0GUKJPo9loRp2h97fMsj1MlCci6c
t0BWqOMsIPZyFHK5D8wJ3YB7CrY8jE4txvXTFOwv4qbhDmr+f693SepPGglM/06kG4HXYnH2XmR/
iEU9thXtVcedDvPFZ1hmzESwbl+OGqGO90JeAFLVm+7u6GZeh7eohHar5xJT7xFJ8HlXYZI+Ik5c
B5XioSYjtCPDU95bW+5rg4O7izKV8VPrc5DeWe2uDT2SMpxkkIDDRBVS4bBnlivKYlAvNrTmrek1
OiZ7LsXwiTlfnUcEdOsg8NOwjSFcAUu1AH7QZy14RiIZojes6LOpSrm2vzFQ9mlSguK0X61zQYqf
EDkIwVbLtGMT/9uE92JjbdcXh6z4Q3iCuP7MzUPhCZeQBwi4SkoqGYcgo//+XFMFLzsZnM6aDykM
OLwfeSGdLqsTHnyH+N4cfyUA7iH7WC2W0+eBpdcETa9qquB4NvTSlMvovhS5h69bOnJcujJapdOF
2VAYAt7hsAThGqK75zRl4dCzR18AucR+BjKi81sLI4NNrUHkRdSFzv0FXhdji/kAqCMlvpB3d/yr
z5YHdTmQMz4A00RnjC6TgMb35CSOouNTFyqzUVymrS2UZOFVUdw24GKnhpnDfkTkdOapeNq76XfF
pA4uuHvSb0Fejz47HGSr/Gk6Hx2rNKYOixMXT8ggeGhbxTsx69WyNdob6otf1e7qI6AGB2Ciar1X
ZEZpMBpUUi+dFhM8c95Bs4uEGi1/Zcy0DTJzBaYzCd533/vQ+4NNtVQrbGLDKSDEjNL/sMaEOASf
sh0p3l026AObE2G7rvW9YSSFTcruVcyM+YKXgzrudrM3QHdVGEJzit6zd+qqBI1L67zNhdpgMXZ7
qXfTYrfIFK7T3maZKBQ4LW+wzZ0txblvj5g4LzIf7BJLhCt/9nuckZgJQGBxU8RiWgipVu+6t4Kw
ipx1vyUy/m+btJcEJOhLbAbp529ZlLwrDbY8GzjfGLriI2VZRpn073mydK+RiyS3/oInOsMxEo/I
92SbdmtihOq5a9JMTm3b1SrdN+VF7EOsEFealSqAu6mqWFuBQc4TJn0C9NuNJcwWQwy/nVhMZJqV
4uQzGXNYzoOn4sgFcRmgJ8uVCjKoQWoOowYmymG42rSuprIVK0smrzT1ZybLGTpoRU0qglkIBy/B
1+1dPRjlRFl22N27bfmgNLdgIyBJumiYf7F6pW/NzBmgBKpZd1z3qwTG1YHFzq2ZAhNmwPbk7Kyw
s5hdiXyWAccPu7Ahc1nwisiA8FmNbIEab+b6l4lExaWS89RyfBq6UNxAxyfbgjY/HfpyHUlT/v4a
Tksrn80qxxUjwZzuxEyn1qQlFmfWqm5Hw1QBO8RlwaErpKiwfn8H+hNOFKM6k8u3gjtLLsPH/Owp
DO5bVVgD7hn3mog4DSI5CvoVT9pxOXcJT+9p0jEoKFfAYMqq3XktfCtQZjh1PHxPaQzGd3WAW97J
IrJ6Ool0OveF9X855y3MbUxURKjGdqHrDe6pXA3vYQRYlxhtgDHLoLNjEux9vfuNtXy/h9F7gIup
Tm92Sblt93dcxLq1xKlEqPJIrLxES2+gV7WP28Ed4CEJSwvmUSZFU26Kg+nwZPtmTBQn4wrDAOCT
jxthWKI+LViWd5BXkQV2Qe3iiF0OveKkTECdL9MP/R+5vq8ak69+g1Aasnoet8COrD0jlLfP59z9
Gv9S9CAdEGAyjitr2y1h/03wMoYeWt3RcoTImS5uIRfiAJIAFsR1XHFgkxLu/e7nFsUHfmlHONG5
nr8aZwEg+6ZdDUJEPHZfHmPQBxcxIoZrOcGjdHCJU5soEFwF2zWijfEi9rofhN31U/fKITVVRFb2
TOskiEJUiyGPYLKWCq60CQ9FvcXwfYk1X6pGfOwhcOzBrg1AoBPOsPX7aPBzQCe0lCdoDid+D/Yl
TNyXbYQJoYrhHRLZ7FDuhicDf5J9q3aOvKnnUN/e5nuGIt6V6aQSpy+q4QicUfw8xXFc7lsK+lur
7YzHa5gfOcc/6G5gR5zdhtdi1Z58al+ZkmmHvgAr1k8RNg6O7ZxqE1zKSnFLXEpqJU1PHZJtrxDM
FiplbCRfLWIF2mcrEsT31BhP3WUIz0d8g6STrqOGlbo4aVZlFC+e8V1FodhGa6Ri4KlgIMTUTQ+L
45lZzKheliJSEu8P3H58KnoDxnhNBm3X231QGZINSB6ojOHtOq0it9EbCvIJhQsZQdxtGyRAiU6z
bXdDHn4LJXJ6sdqTIGANOPRzlO9Xce5JL+I29R+0DCPrpj/wjpOta8FCFOHRFIyabNg+986FVSKq
MX2SAzq/+ew2C9vtQkn2VLduhAJNhnT5/Is7KQJlggN1lW6pZF25UfWPLP8o3hhsnkdXjupdjr8r
T8SVzFw0PI6/gapqk/L2u/G3GZDAgg942MScZuPrJaJA8mQNg2N0PMsFwxCoU9n6IpIQ3Qk9me2I
WHCGHNIlYbvT504ZTTEXPKvlZ57ybVl4spTvHmgC8wMZuz7iPhvz4Dht8jgLIAMSJPRbaa3ZKGW+
pkfFDzoAwHrMThgJLpofa7+exvNIkHymxiWzuxJ8N/5SZiQ2lRoSsfrwpbpTHSkLmLXC2I95hTQM
EBxkgWWKDUPfnG+oBjEqGD+kOKrfuXLo26/NDUemU9ZtIqa5AVKxT7NSocMlRPaXufj1qJ12+jNM
44M8x2IbqxOi8iZxxwk8mbNOJ3ORmaIXssqFGFNwdjO5Mr0Ki1gKjdEAvOg+gD/dugTFvXFx1E2r
2kIhG+skYg5L7PGaAEqR3ObnBjEdf+cj7Oxw7r9PYjq1MPEosQngeYeInU89iqHV3znZ8rAm1QBG
Wc/4mmjD6j/XkB2aILLfyEMBOsI3CJSmHA9IyMjdwsDkMBEevihB3VUQeGxVeVPjT0dEoo4SehQW
Haw8mUs852zPT+/LMvMIk8XCt5Qj3KAxmVC+ovtmDFGVPeHIfqygoIiyOdGsSJ8R5/e2aJNBGLmY
xFIMzE2BLoa7U9ZIFZ8hQ8/g381zgjfEO+7M1oP83N2T91gSQAHVZsLMBxBNVv9nu3/FacT4/JXh
AtYXzztA4850dIaEY6pq+JZPaICWTNy7EgOwhbJTWZ0L34uB9PMJYv5KBHMDKlFhL3B9IQ3wgtAR
6G64R94BuaQKw6IWmhb28RKtJq2pGqhGFJuf6JKhqsbyElaNO6CdwTYTgwdcBxF1gUCDQ+coIHZx
uLcqgGXOd8We6OzOXaFKZVXvvMV6QmCJaTkAnQknuMbhuA5dFTVcsnybct3CRPEQSUf2CBsD5oTX
qjuBUeGmgaKtw/ynsTUuKcXwP6y6MDhhXeYyh9VaaDHnTX1llcJ9PLEMUN4IdQM0V6VxSN/7iIGD
KhL2noKOWDOB91cBPaHT2oRuRVJ7gXij6EUCkp9IyrdrP6g8B4nDhIOyP1gxUWC/WW0o5NyoOX3A
QncWEc4UcSUnL8K+MBeLJVqnIgnyZmbLETmLr3faJeL+XoF1OaNlmHeFJz1lmqtKIbclFVvkFLkw
5E57ZmHnf5kyz/PDboHw0ALAZFRQpsGNWAf2WnNOgK3y81HXKwS8PdUutex8R90e3t5eqRilYR5m
BqyBqxyEowGKqYdtwAgEcE4wwO2Ft2xjULq8EARdyecfsDzhkaBBoU8U1LNsQm1kfJh4DdzA8q6f
oTXCCcrAUh5qgoCaWpMdd0BTUA1iXVUHwMweER+e1rBWTuk/PnV0XLdSs+2vCHXDmvz188oSN2hI
YqXbBk55x9H8DMNnTWG7V7e1Fn00PVJIXC7Rb1xrC1p1bQPYmfiYbhHxV5vPbmySlFkvnhdmEbru
qTF757pYPOZgXb+s6/jvdWdoKeVoO9zg+CJKz9/NJWxJExM6ib8QfAyEDzplZb5QI8/t0HboaBJJ
oKSDkIHXC3Rd15OCTcFgtlmEkbnTQSDNtFkg1BKIjUmrRtwnFc5q54WM3tzpvg8L6DZz30q4FRxz
N9Du4ycErqcuYXK0bfWTI3oYZll1QimmTn7xXWwy00rkqMOwH8m+7/1UspOZsWTccK285tfyCp4/
1noA+YrEAVO9jBNiG4iK6npH8PjDNjWKkNrUPu5+xd0cmN4g3Z+Wfchi9kDLYcJ5gMckzHKZ3sm/
G57UlJql6Tvf61iNjnW6sTn8Uhef756jYoWX/wpq/WyvFiwVrkh4q3gqu8dk+KOXMy3oJJcNcYVq
IOplWJUUN5fgMmuUt7KOhYrRTGv8y/FRns/eQDcxsZpOzcwS5MXnK0EFNUlojieEbeMFRbxstxuF
Ser9ACssH9qx+5nlUgFDWdDFxhjYQlYi+z27zamZ6O0A7SKeSK9Q+/TKmRw7uGXDx89SeS1VXJBR
3ye0sGOB0cOqH6lS32GwNzRxOycmNi97Vfb/zpxcVSdUz4fWGL4Tc1JSQ4+skh9bUThDa9W4vRnf
K2qzVzknw8sWtLFQeXXr8EDY3ie3iY3T6XTtk6raq+umEWmIvoylnIrYi5qfjPNVVRGJBBtDWNT/
ik2Jn+v7VhNpEoBue2988OBhhVmp+QVbpA3G0hIaV51A7ACY+xs06oICpwQRd5rIFuo73xIlspCk
4xGd37UPrXeEc7GRolMDLZLO/F+eM9UDisHRNZN1j5Twpgt+GNN2ABTimMCVWCpzj3rs/wNsWl8s
J8O90fL48fqsLtnqiZcjV1q7+qckfN3HwUYHUwvxGIM2dU9w7CpZMzZVCeP8pQe8tvD+NjnsZ5X6
3l61DFUhOl29bOB/lKbmD9Vbh0DCwTT1yD4++U7tny5HYDiNUP3fWXta3lbY7/HF5GBy96r8+Vm1
lMpTfudV2Zh71a8+BIKIWwucR0anGe5p0PDtDk/y3BDeWyZoG5Xy6ugmVo3rQj7kXf3Y5k0BCv/Q
3rIVVgAQGP+8yQLCMoL1RM+zJUtN/UZeZJlam0RHxqaMUH2qzx4q0Yn8Vy+dgIG2RK6VZYgFe+wf
mk6dJjmNILG5TWHSnVrLyp36UOs+aDLGzVvfGmBbvXCTDD2ThMAEyGiUBpEMBHl1XYTJ1sxI7rn8
NHubDt2qMgPiO1cxHWzB9zEeEfoMM3lL+DIT242h9kxIGif2NDixh8cHg6duMcWZAU0vZwvofmOq
4csyQ3i38f2wC69EsUXSspa4ZLcAEoakjCmuW/Mo4y9Hjdn75yJ/eaNQ96mYN0iJEp6LOM06o0+a
Y5Y6xyGabIAlAz8cRIw+4NZ1XTCok3W+vBdpyENCfzZn7EOaQkZ/wmHwdlxTbK0yI1fY1ZWjmiLh
6dKfQQYnDZMeqNg0ckZK7/UzOHkZ4h0cnirg6XSjkzbEGSSqcwc64DVGMpZbA7Gk/3C8Pib6l3v8
BDs1VQRQ5mPYOHl5GmHvddJslmgRdY/gSIaX7OV92+iAcdF05asyKaat4LT+L5/UTN8sjjJWHAHk
Akzyr3NBih3kVja+YYaFcMqSBVaMQgLr4M2Kdjd0OQyiNL2W+I965wQT04h2SItz/QmUhfRBFSLB
u5loGYuSSK02HtFAkiGLfe5HbgEQ8HcGL59lNnHrrxxHKaZpwr3dIY6YjIw4eHjBCGWo92JHS79K
V3a+F+S9Bu8SoAvj0lLtx5S7SuEs4Oeibr354JauugumNZIpENTkUDWp7+iNIlwCMjQV9NfgpWHK
buzYspBs0LdLtxwq6zy5utFLldVbRirhYBzh3u0eM7nHv99A3cPYn1ANyMp7hUfNI1M7HquVW0y3
fkCTSyFu3bU8lnibnbD6B25BEBt892FAQbrXu1u5X2oStEKEVEgdfxN95FCMSdIyyH8difuhax4O
vnRZcV97GzKQ0yWQGvrLGsuEaLBzLW6arI2sl0k8SFnOhALXtSMOgRle1n+rUOsEiQ3dkBJmFlgw
cKuiR9Ebk0+B3dIBS++9yyG3N9aj3ByKbdM+FxnUf36Cn2PEiFuPyPecG5AHHLd+o7OfGwks6pBf
tPjGvB6FpUly6aK/Ko43qlnp7HnMD/b3BVtfSQUZkvShEl17OOlVCPOvPsqcTTZB++rzVmUhfZu8
5RE5c73bNdiQl305i2YBMtCGjUw4th5N+Kx0UtBB6HqO0vxmlXWSjs7uMCMoF9wVDuak11vjRXlX
97nwsAo6iqTTBPEnx10M/v9tOeuYqAWWeSkws9L19dXwYo+MgzeViHUu0Sf4MRPEOPlRxBQfRBAJ
C0IB3ZEmxBQQ6fN/eVi1UbTJC7OUWhARsju/f/B/HHfcfYQvxyIZGOBJJwF570DCyjkO/nDRTPrQ
GfVR5UNtMi45oYhDslNk2vdsG8GXey1bnDTEbgSIz3zBC/0NIr2oySGSNmTmJuxeM8DYxIQSp+b8
w4c0UC35QIKnuH1tE+aRWAyojQ34ttc0lMz3A/44n+vJZTVF9huxKpMqUw8PUGwPbUym2q3Im3Ig
eZ342jfebiIBFgrz90hLjtUneuye6ozrJIOpoq6DYAfeSq0X1tpuN0mFnqvIveL6d39X9DV0IiPS
cChqnecdL7L3imuixtw4D9jEeQcVDWdLEs2W8+c0cVNKhybZK45ONLEKxf5bc6AqLhETlYyToVqw
A1BZjJdWveL6ylH2pBkt+PjT92JlT6BUm9lHL8gjM+CnjsdcxcpubxFt72T5xIshRoZ3szeZjAz3
O9sk/U+jOY4VB4xL0VBuXj4bV9Ml43Jz3K2Z1YEw+eMpo6BD17xKHesWcl0JGzzYphxrkuZ0p7Ii
0+lmCDW/XcYRCEwOyZXvpQ5Zvq7jhUzeDjAMSnm8xpQiTKIZHljmaJk4UiR9FMyWtyagHU9VHQEU
UCQT6C51c5i28DU1+ebxS1jMaCoO0xjljx5UyYq+FDlAfiK+Tj23dtevsHNoo6G/CLdhWbIleyj1
KQ+AYRR6vqBX94qUQtIIfG00KyajpIlOorCGhnxMsajp8vH0JJWf1bC2AdQIgSMkQbKY7sAWdw/0
fLS9OxVvE3/TN73SIKsibixOIgXyhErExuTjlbXdC3Oi09akqhv989X1vtAEYpWP6TAkG4CI14n7
fFwR7Mt7coHtPguh1COPPQXeiQNA3m0HtwWwCThmxCDGq/sECrNg7kv2a4oIrT30CmQbPjuJ4hQ6
aO5jo6PI/7JN3ia5pIlL/wG1yMPGiglua3w42W4ogh4EwAhkXUjIMCAOujqsBNCX676lLzc7Dap3
inOOOfNUFbvdSzIiT93J0GIniK8VHsJyv4x/yjo5SGvi6K+JYg9/uoKmsLrwSyruyXmV7820I/gE
+pXfufv1PjOadN2b97lLlukO2XVGbraWlLksUoE0PT0DAqwmVanOlWchRiSM9zvXyjTFLGItU3nK
xoeJm+bM+LvBSnsCaWYSBMXICk3zJaFppc1NoMo2+cP8YLvoZKoipgOTJSuXrc9+SoH0D2XG9vrf
0FBidZdVzco8u3sQ5zoL7JVKDSmHVO82WBnX1jrV0vUHWZ+KqOzMxwNFInyi/FhgKprUlkL3IE/j
Rc5JwYN+9Tiw4S9rRagtvv08qcbVYNm0E03X+X+m6u5wJyJ+yORC//zqZiz25ErXp43ZkS7zjIJr
gOUSj4C+tK9AwYcg3sSzOsl+iSe7pll+8Z8EK6E+lxVG/tde9oUj39eoPSm7WBfhdYW+8qVWbXac
2yw/JlEWRuMjJlHhujIPV1sVXC+I/DE9UTt2YouXiDZmW/yeWB66vpR+rOPYjN9Gc6wyZANO2Wmd
ecUjlVIVU3l96CcyXYP4MkjnFroCU92+SvUjjmsJvKI4tUED7T/jaVjpFsrDtTcuPBfWUVahxvl8
/LABzJTpvNgiUi6clpmSdxIbrJiXFiEOLldFWT4FEdxEsVJcbIuaZMDL7UcUq9RMhqtsOrDIP6XM
/rDZCXco8Kounf/CW0OgtGPJvLDN7nKBfFVSeR7iIdWYALgrSZ7BBm/Tov9DNXLcSz4lnk8ZE6e6
zNKnoBwHwrJtYi5AvpdRU6dBzjsbZMyBD5RZ8cuXASSLLm3RtR2/V0mRSOPu97V6AE1ZAALt075/
WWTetzpEhgpA+dQbUk9f48kcVYJXApLiaWRmYSm+1sRx+1sT34mHVd0mCgw8CWE7oYSOqbYvQUQp
EiB1hQY8N8QpmT/olNRyiNnPbtYzjw5vhkMK259tqlvZR1NcotUECSFOJd/PhfLZVcJFQd83PbWq
/y6U9TWV3xHU7jJH5eRx+yWar/FIdmkgNWDlKKe95WdUK8tdRBhjpPKSPZunkvqDz17tyPFhLWrq
6gi7KqD5O2rc5phc+s6R/a+ttdZ1Q0PKxMryYgf8Dujn+qLWEfLLlrSH3vzyrAxspO18yYuSaIC5
JMrQn805dHqcbh7BYBB55MFtVOEz03PInsoE+0PcZIPsEgh85uE8BhG8fSfx5RlVLdMyxQWBtUKI
0F7OLD0TZveV98AQQwaHBXkNqUPNKgP3gSTxRHFDMTwJH1D/HWW/+TcU//7VXbFQ2R8AKitcxTnG
pmnVkAGn3YiCo2LcHpHnEr14VC6OqTvzi6x3S+aUnyY8K6qFhv/9Od9u1K2c7Wq9kHeA2O/eGUhH
pqWZxOUHSyyELUHTsot9Kzjd5gauRZL2fBdShYdAfNi9mZzMBvHRx5Pv4CmrM9lauwWR/9MaHC03
P8MPizz8y6lRJ9Qpzq15KyuolrNDhHSiIKrZGQD14ur0Uos73e9eNbMS86qDJH4B0VSxG6HrTsco
E3ro87EZ76LhVHJXmQr2nT/FK74zxDXrjGiMqBQ844p4lRb/gsjda8OiJNHqKdo63Ld5Vksjswaj
dANJUujw82Ss0fKFeq4QIhCPa8IJFtqnUiONdxdJl2TJ+FL1/Bho0qaRSKGwT0lmDNaUA0YawC5q
i1fNtYI85wyWqxrYZ6UbzoABUmlwhWs2QGJJjU3cx7RhbyI8lFZmjA2eZT14hkUicyHvCQuC8d9f
o+vVlB8Mykw2gqPFZy2sOO9N2yKQl3tWoA2vw3w9bR3qsZHfznxql5yVRi572X1B88lGn7O0KZqA
xtoRZEpHGNSs5Y7PeLsUg8+Y8aGflci0/hEQUaDCT7sU5RLVyuEntpzJBPuRVP3IlryeFv4UQUDk
ZVhkBEk+fdR/l0VmWpjDenBYUSTFP+RPYRjKkEpW2NHfLI5Ndgs6hAb+VcOwbfj040EzBZsNgGhP
eE1Q/iAuQlaD4iYb4Km9NWJY1lE5AJbj/eZilihWf+KD7cgzbm6pvv82T9HvSoB75Wv31tkNbP7q
eLj635QU84MBYrz1Mgw3Rpe7YAVtSSH1uZo3k0KeFP6Fa8MlJFjPsmT/6Ddcmg/ruDdmVPnAZrZM
jFnhHRAt7WZkE++478o3q1wIhLiTxXuxjUqjPWCM69U5E00lu3Tld7KRAJ9OedafUwHWoBtq7lSX
G6P/KOEnESEcmaFouAtjsKFJVq37sl/rtyhJLZr9MWINydituDHBnmVQ48ScQLNisWJbW5eCPwNU
rixJaP5IL+VfmA+bygWOfgacRS3KOOLr6+df2cyPSoN6hM4joCOhi8thynxMfy04izwC+pn3ENCI
Yb1zq2o+FDS+ySad/Id35YYms7Im5DWV8aLlHB6p1Tt3riJa7ejw3HQ799qkZLZfND6KIKoTta1u
pA9994RGQgZY9dcrGMSWzLCokK9qIXSiHIEup49TZaGjBEoV7dVmdjg0Sr4C/GOLF821BnHTPWC0
Z3E0Koyvn6k4bOkaxDl54fBpuJXBbeK7955NVzYQ5D30lEHOTMEQCGh75nNzXtxji+m4129AWeXn
4aWm6eL+d4fX5A5NbBOj234AnyZ3Axy4lOJoMIWGOLOI+nSrQJdlmyiqz4lx7+F4ktQUgBdyY5FT
G4eaHGR/Y1Uojjphdfig53dFe9giCjkkcOYAdLiPZG92d0GM0gEwKFVakhlYu8YHgg9ny/LGI7ix
LLOlUcPmMIYNOtMeMfz9WYzFAjIBIngN7Sp8IsPdXxDfUrE/rIP7La2x+Lf5+HMQi1SVeMt9jSs5
d6GcJPS2+NI7f2C3HFpGLJuNi/Ax33dILb0cvJ4IbMb878kGFXpjILRFrnwXhKwGzw+IQjgef7i2
EsIAHkGd/hT2WVFr50xG33ZELwpEBgeR7UZTONEmSzJUzp2V7qab3jDflQA6jUKRFRHQMhAwDk4Y
HJxKzdVM3o1j1lnVx0M/WrF06rWIc/yip4/af5KE0NX91mBuRL1HZ+oT+TYep0GkHUXKFqlEhCgV
nza7NQqkAbY1t8v/f4RPA7PLskjzvLWBbw8Fug6LAxo8xd+SRdSZAK/tqnqs3XNJfds6slzTxLeN
Cr++JiZ6xaLg3smIi4TuousbHdrX7CVK5e/4OEnbZmtk/rZZWeTKUaMLMDELKSJXaiPDanhxR16q
6Edb2kqBpKhoC56YCSVyTnyMNIMIb+/tinzeRFv2RH/s5xVg2KoEqNHO9iw2Bm1nsE5+10LJ5jQ+
yXHcZpxdiS6fNBTCKcYQTz1ZIjr4FXrU5elvBi9HOzYX0pWee4bet9z0gGre86LP4/g49WH/IHir
TU0aCuXvg1giZIxtbKB5GCYQQ2KPjhoLZ/FiOccsuDnrW7kVh46QjiWsPwrN0ALOsFQu704zneJQ
anPO7stklqC2h7r0WwbIbM5zoLulms0LgdXfL5bPHmR962t+T5TW+p9XjW/xkuSWpguYV3OwGPvG
r0bEXWP/42AHGMbmtIgb5OGhh84G9/3bxB1deiPKcMYiGI7OlVqwMYEdA+1aRjfAjLmoiWhb+2zv
3hOx9BjlaYeNcjbwisuQI6n31yK7kS/8itn6a8oGPjcdxEG0H5S+bQ/oS/41xPzlJeN/eW6quPH0
rx+QrF9PPs0MGl2OpPBGZK436kubRHOr9xD6cE5vixlSVTmByTqUwxtSwBvxDKuMeBzb9qYYoAoC
B1niwgNih7LHJaiViC5VRfT5oxLpWChqAF9p6JAH17eS4x4efTb/TCjkMKjPcXFTc6GRyMdNEmpC
IpZkFhXr28RbIUp2b+SssCwl4VCQPTEeYom6KyVF/TrDoSRdlJQBEqzPXMxO2va6LJaeWwuLW0uK
8zmGfkLr9yh6gPCFyDyQ+Vvp/NEcVpz5Cpvn3yo7qVQnJJD0FVHHc0x8VGVcBhE1H77AJhnQvAw0
rJ0pYR4U2IZ5vZmgV18DoVTmK7sSxuRw5PeLQsi9GzvmCkIIAvQ91sE3XgWQhV8xyxCelNZKkfPa
AO0/0PdyCynS6tapVMfeRvAxzt3I9/HMlCqi0wHKN+qXbLoGTyzq6DsvcCC4VwLJ7gIZAzYepEcf
3XstGS+1c0UdNmAnDAtGbf2w3ImpBCebTb4d+fpsItDaD1iL1LTRDTYKDmIN2aQcD7WpmYAMmdqz
VvYGauw+eYoCPT8/yyerraEzO+SuREGoOpkPKgDPvjkKiae3ry8/I5HvTRUONpioE1MlgzEgYU/U
lKmgVN9AwUgiC9ej/AgJLVPyLGkVky9JIlba6jLRrccbnyn0FTt7cTBxfw4hEbqhEoojr9MQgZ7H
/Cf8dUJdEH/MXXLAAG7sjsmi31Z2i91N1iUHtHky2snXhaug6wKJyVPcimXEGC9cLj0ZfzJmuUq2
Bh+fNqW1sVnInnmYDa9kCjFjH+yufq/A1Wpr5qpCtSPsT6cTm1eawwFrX72xaAFHaNJxmN4vz91u
EdIGIBddRHB4ZXAsjPJPVzS63gzSXJQ6uPKVJjZkDJhanuXnP0EyXzIOULG86/jewBi8lbHcFQyy
qrlnAzsV30mIcqxH+o4asEKi5zYxWfnloRp/8C5uFiDHH9484DFhAaCnedtTh6phgUa0+uuIQyLV
l5My4lEs1OS94on7ltgPB+KuQqklN44UYLnz6UALGHiCuCaUTFoDbRGX/krE50+KO2PGHP84luD+
/XgzmPlapBkXEkIhz47gao6rkmvMoCglmVrPCI626CtIaCC0etfw2RwsJY17UJ9eTB339ZA9iC35
IlOL6tvcgzh7NcK35iyC58sYT1iauMw6u8pMRclKmjFG7Mg90fxxl4moGUgCvmdRXR5goWA1Z1xH
KSIr5woFJzzVTJzorARHi2RzEgTj0EZ17MInhCu4SgXpiFDj3RBZCX2KUmvgM8q8U0IRniJW9xHY
TRdlG8mVDqmGwmj08g9FLHIAg4+J2Lt2Yoa/Uo2NwakGsRvPXwvuSGlSz0gwbbfLh8j4RjTB+e80
aEkRFGyJsSWc+4mjWfmfDuWb6Gzbg5/8uIXFSC0WNHsnSWCPIq9OvWQITB77XBvAqNJafpKKh3Mj
E1xYMMG9D4s9LzSTROKUd9Lp5ByiPkFyxBBgmF6xCKPrp9neyZEHoJRx0YZlObFCzWHGFRD5iyxd
0MLYGxZzdPzptTbUj82MSs0ZTRZw9VXjwhlhkpfQ6tJ5uXo6XVxw/oPE+i6laj5CtGJCoXdZeuEh
puSqtHtF27c10+y9UaJpi7DWjojZ+MDdaezUA2RI988knOQLZXUA9LizqayNUf8L9W8z8GGnKxna
xMCDIqUJxqN/NCEMYcZ9D5Ivb6jNxUkxIkLk0u5m3syXGcQ1b093FkhV3bqF6QRyqdD0eWOyog99
LuyUsxgs2PqgyloN72Esqf3iyDaxAifABpIK+5MabfZTgG8CXMBnA0HewF0a1gtgazfWQVxFScEv
KL0j/NEWxRs6vN5XSXAWwL4y+hxTWZyW+rTDH9RfMBS3f1O/CMHCIW4jSVQWpa4BBgdfXeXV23/f
Ll7TTi+/eVhywGLbYZ/ks75jtIZ2EoRN+GsQwI167xu7f4+3ZrKqw8JSMSsmlFs3dNqe65sFqhJx
oYEzXcmzeHJ5TVmiN/bECXmzqiBuMS56fSM/LyatNHdreJziRV65sJuS2QTWKkfgA4CQ60gUNaCz
1uMTDlKZdgYMS8NUyjmUKeLS5oG9yG+QkWaO2ekzgZE3fXuAYE1bVbwLa6V4mrqASoEikGwhUWl5
z23t+Com1goX1lbYZF90NymrkvaQPYrQDkoP75lKrqSbGGCqA5iXJdJyoDTpBGygsGqjVcHCVngi
OYJc7hQkuHwFizzYe0MkRmrZs/LBADz/VGbWE8YhBqSW4LP51pUH0N9/zY3HitKS3lcAeYZuMQBN
kPuQeVd9lNSy8lKM37iucANbGhiA84gbrqsq/FEs6RmQsu7cgQVqb7RT2gEAVF3twRtPmknHotmE
b/HXUYu5xzX0bNlzaeS3qslyoczcWdCgvgd/ceUy7jhHLYQS+RP1KRaNduuCajchpClSGg45i51U
83iq3YR/ysedAZkGlVKv6qRpZFQTywDA3DzK7qy+kHSsKLivFUuXZ6S0okv2i86+aOfhgtUMe7Kl
G8+8KMs9CcGpS6kOFvk/3aGQah0UTcL1UkvZEr2nDn+HN4CJ5kw9Kr7yn3oZxjqRCNatH46ET+tX
8sFzwGwFrjpIB7v2xKl0DHCwr6rVAnMIItdAvB0yATwwsYuIx+KyvnkbWjH1JROXcU4g+BsOXr12
r/y43F7mubZrI2GP8T0y51HZ9zuJYXLBBBGFao05setG9pJi0i9JxnYgNTbea7UK4gvETDn7iRUO
huAlvHTKjr/k9b5awEZHsAAHP+TPcu8OMQZgx/DMoSs/ZvxAacxF7YueCyY0dxiR22d+XL8xVeFj
td3VrwjFGHUcjCpifActhSIJrO8pv3KTzo1TI8JBYhs4tUb4tllMiHq3/bWKQE4wsq0bHXNXzkGG
CE4C4mUY1cFnIenP5pXI4/Shb6r9NUiw2eedxs3L5cTnmYuo1Ea1BE9uea/Zs6HEc2SCkZywxDki
jwVxkOMnA3jJ0+rgmZ/Z4ovOtBXmHkgDG5fwIsvkFEOaVOzKqMFlz5qq2hTxnoB89viIiy3Ka1kQ
kxUUidUW9uJ+9dwmSevSa9wc27U0mKXWSh49N9CzKcX7l95leVFGDUd1E595ZtY9glsDzSY0aEy6
i3M9qPPzW0MBLlBk7g2+ETsUXoN5xSUY+vt15bjzMIDuuE3o6cFFJLvG18zDLWlzbENthHji0LLB
jFifllhC8Wq4j3L+NvuvrK6DMIHgt/V7pXPRi9VJLwt6Iy8d9IoDj0IQioSApnqIrQVyRgTGC3xH
47/IolQLSNUInhjjFRdJpG9eWMsX
`pragma protect end_protected
