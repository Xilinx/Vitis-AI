/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 303392)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2k6YATDgJl93TomqNwQrJc8NdbI+vcDjdCMLVmchv38lW8s//oBIOH7o
y1C3258dieGAccHAAyxg2xEdUIp1DS72+Fw/aRrst1Yl5PXhC23Tnb6VqXb8ayOfqz0d/gFDhAnr
UEYSabHC3Q9gjOt804dYgEPhaBbYCGCQ+kyxxl7JVraKg8U84+GtnjTHbGrKhDv7lZralyJh2rQ/
ccOzHRo6VUrZL9ofpTCrPpjMKlJOcNLUwJEhxd00pdFJCYsCSXCj2YsFTcrLp69gT0JK/xMr5PIt
HCXv8Zzhl8krpY+O0nZEinV2aHvZxejb1HAUqq/kpEogadHozDdW5ORKy8bKSZ8DB6YIi535Jeyb
kQDvqeEHzn+8P7Rjhs736Zc13uS/RGyETH6QDL24tegesUX2klAn7GF4eJ1uIB7lH5SbIborfb9j
EWsWaMM4M/nf/Eze94lLn88GU7jac91lDQodUeLZDYdFD4fBFF6kBJoBRjTavkce/K/18YW6Sor7
M5yaXT16tQmI19ZGueMdEcm6iru6HdTy/HoQIXrhK77XPWU13Yr4r/j+NhsPgavr2fRo5ACFIJAX
nrd7mUeGVkUWXoX376NwXBBIdC0C/nldBro4eciILh+tnvtuwk/cylcza8cF9XUh1jDykiCmK/Md
Q1DN0RntBOOAfX0q1U1h6JJ9zJaPnxxz+jXD2WE/52cb2PHFiT3dvrZjJCUpouW8Xg/b5FQurhy2
3hLIDr/iEwueX0uAtkV67JTNwmpRyiPGgVxYirGXz1ttapUbxsQ/UbovWbORa2HrZ+vooKAgwpkB
ZpLWiaklxxtN9Vj1So0kJeioEKAuClRWB5V39HgmVYX4E2HbTphhjD69iX8WlEONAISJCEcuov9N
Lp9csxD5CNP4uz6qvTUAUvfnPxsphOqp/2Q0qaSBHwL5f3Fag9QHscuyAR5L4y0AS9c4+tq+h02+
dS6DDeENyo2DSBilz4nDSI+5gSGOegZ7RdCrdWT5sm+yryg/05JrGKmDFLtQeMHdzI83RfnaUn5j
zjmqKd/h1C+s2vcE61TFFVyexFANfqeJ5ZQw/b7DlusWVzLWNiD6sAU90QhmfKN1yekIcQiVV0EG
MCEa23DRZOhl1FJpSJjXO9FWRkk/rWD0d41mtUa5AlEroMVKYdR6CgOMD/HYwGNLLvzDG7W11K5s
VhBflz4Cc9C0LliyeVQPC4ptAMmvDK7NHBrZch42K/+xJGhSDg/A+xdIMfOvQHjVsAxGlj0p+mGE
OdzaU4yT+X48sSEgf+VHNHHZkzV7HDgY0Piq6fvUPKO1DXk9KBawR2AwWq56jr4lcs14Ml0BaxtK
5VBnVW/2IPsQB2psWVxVlPG3Ah/zfiRt0uMrAH7+VFsB4gFptJ1YK9Atwme5uSIwSbjVlgrnK0cb
h7PcKlSSZ8nKyGGIBn/SnjQ3+KfTzbLKA9E4DegitAn6qo2md4kz2Tt5JpMApnkn5JO6icp9iE/k
/bHvCkudEuGkEBIqd6+8U4AEkyzNKOOkunRkzvEuMXEfgPEkCSDtKi2wo8za44Y9gwL76kmOG/S+
bRRUzzTnFkdVJIMN3O/mOvU+v6vzmsX3RUy+WmakL2o8wK8hfDs2f8gGCJ1kiqH6VuxbUkMX0QvW
vKBPksm5eC+JWosXG2Tfay22KiF3oDQNaqiy9qytRPNlgiWUDDOuN9dp/Afv70h65w5UdaeQeK00
Ztanc0ZtP3r4CpclWJ3pOqoG2FbCsJTgCEnvuux8yU3brzxfRitIwrYL9yh2GCoSvSMVHU9eoAu/
LLGRsuhqLaekifw3DKxEtzBzr7Z8KYZ9HsSo3xKKB2o8unESkkwMVU3LYABbH2+wWnPxQw/j0FmX
fRiuuvH4FnsXGK63nJkbGWJWlqIqfl3RFJe93WhwHMcyBmke989PysZkpooBK9HBXvwR3tI88uCM
20fPcD96yxDZzqK3Pm8o3nFVTYWN49RWSPWxDTWOqaXlBSqhx0GtPCR2iLm3w2gHalt/CUfjFUWI
ulh5gs6uroJDwtmFEGcrX9dsWwMYL7u1A9rBXqniZYDGtC0k6D5FKFivgvbtCBtJv+/ooIjMfb8p
6jYJ7SudEG82y+PmOUWCmKN8a7PCeymRZ4W4XPjbXQGDkEH6l7r09l+ftdPjiC9spwr+G/G1toF8
nhG/v17sgyPZdRQkiAdCPdWycsMs0sEU93tzFTI+PzTrGAIZVVi3uC4X+fBjobPhkFA5yLSzMpMj
xv1bCgDW8mxhpmH7gSIa5YHr+gRU1HVVTAr8daIhwfy3jLqvHe60+7rQ5weSHUozJSM2xs7t82za
GCTLCmXtzkFuwZOZQbtxDy7ETwmKIadSfSuoR5fuIfaCj7O5Zn1OqMGInNc7amuPIMLIlCgCTXvW
dF9HDZJ7sWhyx/P8xe+J7Ozhe+WOyXWq8rR4cCNn2tJbCHX1+Ro57Vohnw4XzQ9yaxek2SRpBILz
BzrrPot0q550gHlM6a0KmNqHsqxfVDvGZNdQ2qjnktXy0JzwUTuN2Axg9iwqxfzF9pVWq+75ul6k
UvXbY16nnGOvJCGFleEVxoZIxfa4MgplgHnzFavRhn/AnAUaLL+dHkbCnL3trIoCSRH4CJIec7F5
CBL7xlfHNyjogVgOMl+cOBkYR/HcI/PVUzUUXvOZzSydwB5Wg4HeivIkYo/FVaCSRqlmb/jsHouR
wkGllmka6urTElLhZsg8lrbNXp4kdrwi+xqUqpGUmAKcjrbuVkmY1UCaMWVv5SPS4jYx86tHGYic
xgQAKuv3ggbvZ80cZAgOJefsDnDuV2CJzXRyeTbBaMKhFNhk89JGTRqxAO5SFmaadCd18JDkJx4p
TSzfds4+HW5pI4Dkq64LcJ1LHuFQZdGio7jr6pY9NRoMjFQqITboX/RnS1q/Jnt2zyninCffJ3Ve
gVg+6dXduflZ9U01/kzcrhwggI/ThGtoyGMtoAfR9iJnO/bQB5ZmoiQdB8PgJetHDZPEXr3csBc4
PwXa1kkikOhDdtN2AEWJ/cPWeiQd7qD88pbZGK1lvIj4u506iHaQM78FKPSbfRgqFeA5OLiAmYYf
EOEebtVcqP1S6oS1DrBNNEgM4ZfOVobZ9QcnXha0qy1TEhIg1B45bxPq8pb+4tjTTGASZnYC9J61
oKCXVgeemNQP4n2/XycCQPObY3OEtuiSqwrkd9aajQIxz2dXSapi3QkyIFVcTtcXtO8lOT8iyoPw
b5Wy0S2kIPlDh9G4+1hiYcBP+3S6eLn2tMLqMhohExFCygleP7N17Y6NmqSy3A8hgEDqYGNp9+6R
nY7xn9XFzZWoX6refe0rxrXzWxzk8wgaftrs64Lqhd2S5cgSqTFj7jk/59a8V4FHFtbifn1Udy2H
neQ8SzjtNFJ1AVrfIKzt0MgX4+O5ugkq61Ekbatw9hozRYqEJvnacFljjFTHNm74HMGB6ijbBtpU
nI2qMC2fVdKG4C8idRYq+oT/bGeebKnf6y0ibi/Wsvqo0TKu1QqKx+oqwISSJyjoGMLVjfAD9dGS
Ucmh1FlAmW1hPj7Pn/PZzRmxXd5D+9xZSfPSsrMbkU3LaM+S6yH55VhwTj6jqzGInNCbyNlMjgpZ
PJCfcamaxMmHw5VhGNXksDTYEEO1lJaLpBE4dWhG2Zj34Wf2sZM8AINc+LpgYHmBSsvIMSedbqPg
JNNBDzD9IFKC0uLpznLKsNfunu/8ErtxTAlb2YbP7+2g6RFDCeHpkkQSwaiMnd96KG6dtCz420CU
MarK9AEmcWZMGeXwjLsZfQMykRR+cK9oA/RI5lnFeLoVAARMfBZJbIElSxnkP7Xl221f43wLKmpH
IKpsi475uU/Juk87WtPHnvCyr0PsZeQrx+p3r2jTQephQzekjuPbj/9FMeXZANsjT3D1M95NvjmA
JkiOb4Geg2a/YWgJBUJcr03MSTgiW1fnG1BRBPZiknZaE8133w6gaG2BE1zQTv91sEp/p7mPOIQc
dJeWavGmU3XzvB/XSqLl8OCFgUHm0vaIrlsR3slFKMDv4EgADbTZWUVLS0h4rWB1FetdD9DmVLbL
EnE2BBfUVXno7ytA/unDOkwjNZzRV+Ksfe1pTYMNuwA6trpZRgtPT66urzC7xlxOjbnmyXWM88PL
xJ5s9wEu0XUSYGWAskcGrpL2gxKqZr2NdGKePYLsKfxdFHPPVC++WBE3FbHMFWh2FrWXFg9znYQb
VfZtdH2OAabI7TxoZMwESKhUKaVm80SlvXt4xKrK2dek3veYY/IwVQXQDeVjluh4kC/Pio26t6wH
UzIlGDAZI0p2fZKctsoj91T8mJXgNR29Ic4NhAO+GOHvpqGLQwaJmAf5XihFzCH5ZGxPTQScCGqI
Gpclsl2bBqccg0BPMD2z78qk1slB+ktuKnrLP7meEg22YISkpqVwURHV3G4yaYYwBQiVjN4sh1Hs
YeypeYJSqzG1s0gKodyw1nv6jV4/jOAaNkN3CON2Gs9vt8vFfxK7D+9tWGkVOK8HCwsixWjF/16c
VuRDQpgja7WHSD4azwOqwzLsEkxFeUTVwe46gY928lHL35hVmEKB/KZ8+/ZDt3fKoBmzAHG9+/l0
OPzeOpNd69Svjrbg9fcVGA4KDZODChz1FGsOAd8ca4cgCoMi9WzDIGSAINVwUwlLKWVc1kVYYrVL
UP4vxGM4CbSBMt4DKblsrc/C4MrQ4gSOOcESdDy+OVC/5SrSLarwy+GrZ5g6GRvpEFLcPV/OU8Wt
pfByXyfMx3ZL6Pi/zyC0nZCYngYm8duPmsTO8hIiG3CmFmdPWeahzWxvAR5ffRTAfXmKBbyhu/MB
teR6pqQobaOex37NW6JLaYSYDax+MtygrjnVNbmo4GMk7miQNEKILlPoGCERYqc1Wakv2wcZ90/o
mvP8TsX/NtRu2q+htndBuPywqjEFZQ7Bc4/ktztQyd6LuzZ4rZMffPGluhBhj8EZx1Bohleym5Qq
eeXQsxHr0i/+7sWP9PRwUa8hxkrLxYQHvdD8pwa5XO+fREvi4+Idmlgn/jSgn3leJjXNA1B2BrpK
KFcxFWB3aIm6nF9qXB1YTushA3uVx23HRs977rIvAgla+3Ymo+tYXEIvjzBCfTCfRwic21bXp9KE
+4tvRnEPRxUnRNOAQOKk1wbelvzIouhLrolFtxPwUjn7YWV/infejN1UY6x9T4WtA+NBjd2S3UWX
ouhib6QdWPM49g8EmMT+0AajVbNYvafgtFuDMoPMU5zhFNn+Hq+TDv26XXMDam6PtnijE9nEHRjo
fRXcX27XISE/EfX8JvSi8vHbp9AqsUbgYYeqanBwThSP/AG8Zt1MG9jtHVI5+fITpmj8jRtq840X
RlESM5w62usayp+KJAAdAM2QSc1XNO2GVSs+2GXdAaaPwCyPmW/ezrbg0tPo+r9QNQLvramurnZs
Va8PLD7DS9PIdY05bAo+ogU63khzMLlb3pCdHTrGDzuJ08PaKE5eko0DexONsXRZ8tyMUApqi8D1
ClRfwO6xUOPy+ayQVQj2KVLibGRz0GWfCSfqRdM/95BksB3Jz+l4QDTUwXzOW2f79m7kWmTpPFR0
DCPuCfA6BScAFlvdAnggwGG79ELz9aBIR0OxNy66JX6asgkt8gcOWfnj0QN4IwJZa6nMggNvQZaO
x7z9iXPA/37+w1OEIh7YqwLBxg7RpSO+53A8DLPwxyvxb0AIk2JTiIKOYP9JIoiJEaN393Csrxef
7rMkx4htzfiz2DBjPCZ0Xuorsx4BvZxXpPvGhn04gQOyz/zVckS5K0eXHRLXS8K1LVITiMLfYTdc
afaMAWgabY//fih0CPhfHlet2FfHxmU/ZcWCDe9oSYwUzvsi04Dea8Hd/bnSuBz5hZeIbqGuYCLl
M/N1Cu79rFzlKnWBX7GOre/rMDZVL2nIIwfKxudJB3ZbTe0Ieriy5TdiaEMbZCYgjX4GWXOfKC7S
FFXafKe4gqOqKH0Si0KdLCU8zwZLbV924S5seApbGGWZm5OBfspzoJ6Q/989Ggx3Z0csqrWk1QcW
wojKlIg+RKY0hzr7FEWSGDq9tVQE1z2dq25CriAZgrZMO6NZqiPDJa9VN4TVGHh02wjICOhm0X2e
/eJIqcZU326M08DTQ+xLfQsIdr383w3IK1L6KhH6sdOx3bRLtl4sSVCa6Cn6RDTzUbOraxs5KcHQ
uYQyycQExEcbKfk7T2cmCucQ6TV1aJNRn/yMQs2JU7+9WTSASvhkHhA7p3AnU3K40qclIopt9qPl
ixwQ/jQDzF6RoNzL2rpR6O6SWnZlWrEY0SIIIZ5Qd4fbZJpF9kanHptf8/+thfvL1yxozr83XbYU
WGmjPIktqschGGTcBuMY+0t5MSuRN1FH3bWKIE2v6QgzAxAHeU2IFwsm8+6Yc5JnHT8BA+NoPN1H
owYvVsYQjmmhcrKyCOEdluyCrsz/2tNYDuKs6LoH84mMgvUywoEBeZPEdSZe8c7B/MHK5rYQE+d/
foNQJ7wYxwfjIiX4oY8a83OwdujJDdHYvL63nR3uU6Kans9amPWZbSJrxr5HHHCLN0RXNLW4MQRy
YAK09qmeqcOUuVETgbxh7I68RQnPLGMsYVzi0I+khhJX9P8qfcbuoN6QDwJux59j4yJdqe1Ojd8u
/BidGe+uF7u+8kjfbn/kSAOzwolSTWCxcJgnAIgDhmURclcSav5ivBrzgWPZ7roQFFI7CT9DdCm+
3ccAVlGtqkfD7z6rj+tH++eQtyrneH8SnoihMZZwpnm0SRjw3eIXtCOGa03oGyl1F31m5iOHsv3u
oKEO/CaJiixL2FDxaDUzaEKJ6jw68ZQQYTSQfqOxDJFGEA0UR37W+QJemF4Ed5dQDoE/AsdM7kg+
wYkJI5kQTiPl1JID/H0fRaUBXQ6rfEcAOacVjUgN8Ng9+ITf3GXaEaUcYpN26dMEAWRE8MQOfVMm
O+wM1fzJg3OZjc6rbpJQxV3SlTXhV6gqUDhPyojSnBVUjx6NxjHDnDXza+TCNBfbbAOfWdT/MJZ/
da8i/ix679y7QZogVAdLbPf0sku7hks4k5sT+M+3fRPN9O2ifmMAzdQIAkhByEqQPqo6vKrCKJy6
HV0SKbynb1jZcU2Gy0Ef3jsmqryhM1na8VUBZTtOZNutVXNeGhN7jFsv57JyqhX++ZEb4ma+XTwe
iFQ8h1FSB1fk3V2shVuUhqmORRxX2E5kcdvSPz3/tmbYmb6hIcUO/4hUCc5evLlJ8PslLVdKbEe1
fMR90u7ZmqI2hl+IszVR1ql0RFv5taXwVsLrk/vPOt1xleL+6lZuq9k08jybEvdN/iwysCgKroqV
pUdAK13ixgnp7/s5MoPxTZjvQdI5kbWT8nO2WbbivXAw50vKSEowTm2RQnlDJF4adcqFaU3rw43e
T7Ds32sD1FQooyr0UqhvxBXkyV90xDnnDVrU2bBSplil5bVfimy6xavjten/FpP0e0t/hb+O6Wrp
nnaJGU72IzrXSDzmCDEDiY5+JSLVM1Pp+jD/oWco61yb0Z879/dbDCRS1n0RRaieSSxwh3eoRwLD
4gMFXTTK3+Y5eYPJZCLF8vKOqvQE1jlNfsulgvhFVdgxZBh7dURxvVsU5YJVp45u3Nob9l+5SnCj
SeqfEHpEsSN83MuF9THUCOx+9+gUrrlnZTvJy9sgVlXP8apjN+kvLrSHZSreXKBRqko+uPemkZYJ
OOVfjBqJvjWxpwXQh/2inze6+3BqrkeqO3hAtBKRN6uJTVPgPEo3FiUgvPUW3ySuF2ezaCqo27k/
dJPoTxj/qrWb6nwigju+O/UuNsGgWvaztxgavIm9bUhmuTC7G+yM15Zhjf6xI5inapj4/5TVoA+/
gYRLbK03UDPSA+z1bKenkWQ19p2c/MIXIr5yxM8knJ4CKVgruHKJFOwTzvETY/ND2VOZQPDqABiN
rUFPYUcXsX48K+3aYzoDDMl4JtU59ZyI5DPjRNfb2Fjsz0cmaIGSzIFVyLU/1OTaQ/gjJ3XUv938
hfpL+h8zO7/vX3rFzkDKy0dwET+lwvHuIl/nLPTjJANxX5Y2LplDXbvgVgiEsJ05UV2EKJlLv91W
3kJBgrh2NiHPLwoQB4N7wZY2JvWMb6WD06Q3zy3Sx12WjY36ccZTYTFdcHK4j3F/1oE0dXKzS+jr
FbkJM0RmrrJQgnFdh25Ro9LVDxiJUzAbpfBlUm9RA7Q7muEeytAYcpWvP0RcPFe7K4Q9DtddutVX
DIpsV+wvH44OCHtN8DqRKbmbWxSzRq8DheyzQhkKY4GvCA0VQQQrmk69Bx/lmbznQLbn69M+pEnf
zY+upwoYbCJdc9vJkmoMHjAXwaGGrBBf73mBCelxOX0p8KR6kuZsxoSN4+lAEAOfbF96G99E9Cm7
lK9VpaQEhWLwEYMzrBWCK1MqHkxvTNBoyFtszFLWMzMIhxSr7rjlq5HFZ6CrZB5BN8TTnxNmTmlQ
ecOXJg0KjicjZX349nccMCDxdQ3avEc0fYNxk3xdkD4NdhLJzwRkVTyIIYID3YbBC/n/Ddfo/IAC
RR1ZPX3vTikowUydL3jWvj7Io+b1Erw9MYVnYPHAleVq2HPld3iAohcjjd1EPIHG4QlKPI1ZDsnQ
u7tUknmxza/g3r5Ns75LKT1gmcZN8inRz5pAwrsoBk536H1YrVjtJuMC2df0fUOYlOBhkTFi0KP7
s8yT9b89zBjUorYPV9b5NJ4iQ3mz/b4F3fqkrFS69wtEVgMNkp3fK4qop0Wyvw+ZyTSGEv+VVhwj
UXetq5wrUkgxjjVQezrUY5RJyBZck0Z4oFnwuSjrfOKErd5GU9W/Mx6f+w9fRYbfa2XBk66fVMSV
kevLcd4p9doCm5wlcLiHxgjKOhh3li5p4hfuDZHVF5kW++485uwe2rodjAGLNuuyX1YfbSoFhpad
OQoovrou6vuJbqn0WWIFFdI/X5noaS6xhY+2larRxX7EK6kSxEaGv0qgC3eRpV6lDXe+ZS50TEEw
28Nyhy20sCNNAaRNXt4IY48hb77sX7TgcVoZZD4vCVTTL8hsJHwuTdzN4LwHUI2tTBpwjFMKkG96
pMx+3AerGwMzQeMdVnwkgyz/J2vbWLQzTcXFklaxsjDXAIzoSxPFAEGpeb7PegTQU7yHM7ptpLd4
B94r1i1wlM46AWPQsJjq2GrZnk+jI1VGp9U2B3UfPbObYwltcIiEpYrVnRn0P4COxY0I3xqPJIM/
SlDVMu78jE/KAGecA9qL2V7aDS6J+VXf3rfAKcW+cg9gt63SxE1eiAhweUriIURRqz60QIQH2grY
iLIBrjee0gzSmLljSTiTJcS/HGm9mAdBGQG0CYUjTP5v4VT7tzrXPn5zgI4U84zsdE5PA0Rnm4s9
dDPl64TRKN35tdappPh2L7PFrwY2hGCi1W1PY4qLluFgozk0ABoq94WfPG3TCCH0p4iFb1KYWSDx
4ZLVdhm4g9O6Opo7GsHsZlSCHiI9LQSfyWqEVjlAjDLaJZuD3wAYCqTURIHVxnMQBExvqGUIjk8l
N9JCLOe4EwZ6lgVQpoS48vNx7fO6SLxASzNWHteY5WkefV/xGOUxreFCcFV5fYaJcu3jqbY9Dpw2
QZDKqw+XYG0/B6GjhvIhX58ncCMyEodeKiC98Jmh0ihifgMZxaVOtv1UvjJMo9GQe03EOp+ZvhZh
qjZSsu5xznxa973BVZWpMFIS9WjrDiMkWvQPl3dfAAQqGTrr+YgPz0hPZUgWj4z1pM28jMjJT0Ja
0XLxK5XZ6495KoxLncomzaoiC7JZvtFhACYO+WOkOl3vb3uNx5lPNPiHSgl1o3c9Cpm/eFNf/Kh1
tWNWUrjf1PL4x73jfRj8kzvIyRsHzZrUAxZ2h7tiMJG5wlduVVyCJKVp5AjEZIjT9VdLSTVKrLvY
BnumPq901MrxOVRv1cm4/oqLIIB9npzU3r9c5JB+J1mR21SVVJHEuQT7RZBNeAI/Busjep1Q87PR
jxqdEU7RrxkBykI6iJhsc90GMbl6xFKHGxApCsZxMCVxdNHf+wY/MGH6YxwOM97kuiRY0RU+g6kh
CRcbV1cp8b7zx+A/PnTAxT6i+BuphqCMno4+wOjd2KsYOGCc5Om+evdFRa3UrqftJGOxeCp4f7/4
O6F/b23mY+FC/n0AkiTYFODPPl29u3Py2Vpp05W7TTVs9uh/n1h3tsfid8AgvzX//LJfo3ecgbwm
Fty5phZ3+DrG+m3wsSLPxj20uNMRNhiwvUafHaLoa4FZKbsbK5Z9wSrZu71uhbmVTH7Xpp8EP0hS
Er1y1Myg/UIyuS6YblNJxxqvQPCS4N4D4fDoofLwIbfeKGGB58pwgat0wcUySXB0Y153GTIakdJP
Vrx4JgGRGg5HeGaOZbD1Y7jdwbTg+UPz1j96IpOIOix3KCKq7qO/DfD8aWurNfchV5PogLiyuFPX
VciePMKuq3mua1UcIk8vZuYCexKWbv4h1VBqKi25hTJnJPOH8GaqKf6s1wYoeB0eryAPeT/LJUrl
n4BlA7Oj9V/N0MuYFNgd0JB78Yfq7cGHJ9DhH3WAs0BHQZrdoDeYOGYEc2DnA32PrCcx2WUQE3SO
7I3Zvhf0bVw0hQm1j/XFj6oMQmhF8bwsxHROK5JbK/a6YXsmDQs0QOJwpAR9n8Ly4pNt0ICfqvNi
hswWgYKGB065iz/lKlcbxj/9E03MXsBnavlKMaVZxIavU1gwlcplJt5PqtmMoYXkq3h/KBsJ8e74
h3KEuo4oLP5spvfiQlTz8YM/AC9VU29tWaRwJH1HTzufF6VbrTDhHRWQlcWazVOIDGcumnjogQ+M
vIoOSzzZKKjY1qXBWFyWKf0iPMVrbX3aCMkrCicenU/vpelPVEDogZNa1eIZCklt5c682AqUVAgr
YWT2Jclf5YvjRWQXAwv+U/AvuK7mSu/ZJkl2jjbheAY1mUTRzRMtWKz4Aap3/66RCPDhTU4YKTFf
xfUaScRZLfIqMyWdf0lqeQemS2LqBYFvt1kjmxiHLwvsp5urpPhDtPCuDFDvMhjglifL86kpsNAr
A6PysrpCI2pGXa0aHuZKMuusDuyu8sh9H7n9wJM0XxxCKgBGa7wwi2C5V5GM3cOAYzHSUn6zAzqF
pZeVb3h07qq+W9O0zvFgnJ2V/oXT1erc7rGWkNDS3A81LzFKjsVsj1mkB0WublPQRt1DNCtNkJbi
7HZRQZKY5BlamMwOZyYu+2/tKihxRBOxqHvRZNq5ePtSLs8A9kxOXKqTwJM+vIHDcQfv8I/qDtKb
+X1SHLgFFWRS7z2toiSQT2poVDiCpL7RGyHNHD1/f5mWrUKXsyIBu6MRHdxDu2nALw6hwey84CKU
Rvc038gFqSZQn8KufwvWi7v3LGosGSfVhVH4Bi6B7B6lPH3zz/7sqYlKYTdhEmW5VpuuSneO7IFP
OviatCZylbEUpsAqTMtOMhuDoG4A4j4x5LEHGdhVTY8Xul38NP/im/Bebt8+ic/zTTQ7AV9EQXFT
eboCOc8q7g2hEeu/qpxgUKcxcz2oLY7Nv75hXLS20R6BxsWhCdNTbr1lCV9J7NTfRNfvKJi29YG+
oeWNZRF/gHZTd5CRIVmS6+IqleIha828eMlWAFIxLoWpHjO9WwvrJ3liHk4eamSd5A/2n5CHXHIG
QkW1BxivitGhuzjxZXkk1hY/Ziv1yUkm+dNpnZ35t1Kf2ETX9jEQtu5kwquw4WizO2XUk6OoRQXS
5NQdLhsBYef1xhrRVJ0jvI1iaFP2pwpxiPGbhPzrZbrCW3Bzrp1thCDFK/pWyNM3Y4fC8finnTNY
MMqcpHN0uvwOTyMrvipRUqYGOHwOPerr/sMaozMT9cH9UdKlVcGYu9tMvk+ZJpQCH3yHMM63Su7F
zZ+rk9E8KYgQR2WrpOPrkdUevOX/It8DUHztgDASFw/iB1cGUNUmCxG8D09vyBYa7CpAD4k7yq9g
UvE1rkpZ0cKwLEvan1lafmr1BooQUcMxYlsmzvPYO4YqBgfJEnF/BR+VWI284Vr7ynVcxW70NLRA
QwlMUkv1YXcEmc/UAFFOlankkL3ONzGPX/KW2e/ZHqyoDUWzf+0vDi/BBlVPsGtVAlV0WyOt0+L4
DUbY2tVZVSOYvZrBw6iIedLNIbExmuxIDECjtax6AKNfwgaOIl4/A6TdQzDK2tmZ4UzYhiZDi/4S
BANSqmRv2axPxNolj1zMciPPlQlCp8xvQDj6dQQGeh4xXU41EQ6tcMyXNs/Xx6yj9m7f13/4vRK4
PgAaEFtTcmO2Y9kbPs2ZnwI10emhmhIZ/ODX4RYWf4+gHZqBh2i/HVr12YwHnLeAD+pqzFQ+wgCJ
+meMNyueEFDjdIVOnOBLEXqoLETD9bsa6hV00iVTUPKLNr8Zbmabl8dYLArEh3y/+5kutIfhf6D1
p8Y2KjevFYlx4YmE6w0FA99AEllDNuyt0luMSDlRP7fpKXKmhH+zFBcQ6CZFLOFrtxTerQvm9eXm
IzKzZutR/6mTXpfGy5y+i+dv+uNF3FCfATZo/HQ/oWKC+INMrM1UQob6/Sw9xFqPEs+5k2wZ6a+Q
tS36Zo+xlFZbnGNTq6HpEOsr+kLmfVFx2mYgVuFI6rhqkWllUiawHPSBunY4a2kzpO35mkZQiQU7
ylHK2EkJKYLd8fb7SnYGOhukyB02HVCnmC6hmz4FDg6oHP2hXsNwm0olDoWegtMt17hJeTcbVusy
bdJfLjcTN+qgaTMCHXqJwHArL/achiBI/KLSintzPzk8Wfgk7L/sGdc9q328iK5WU1gGapuQLp9e
6DuSz+3YMQBQ4TacQV3vqMT8gSoG/N+Zq1OdYaDGc/YFqxFgGyVCZgS7qE6MkqkxjHUbAZAzizTA
kg1pHYkOAJBA1x6P/Pfnm2XAGHvWm9Shozf45qDcGeovFL9RZ3jIHuHKcC4FC3dEgtLz06AN1kDk
D0pPgcSs0cqOiwAGciBwPyr7VHpEqzP2+M34MDcv/8nrEaKc2nWc5NMB3NhTBepJXy2SBmKuwdcI
NVJON2UeU1nbV77MsTDg9f8N9lqMa+ucrj4rOoOy8vlm6OBRC/ykLAjQ1EvCznHBviOoUZTyU6Pe
t6InUS2qKm1UfiSrPnlKMKM8GqAz360Fktz33TrkrnneMzfBdSA+3hvkOnW1bXpPYba7m1RBnbPq
3A4NAjHGNswzqs9AbqlyDx4WhZNbhPsQzYHlaTjV3C97OqqNDfBphY6a/P3ULu7b8mWcBqkmxgP2
w8VMhtQD6vxBIgfdsXvbFaSxJYQVTH4MzEL1EtgV9xzIm21jvJE7qkDIoMEAmtCFR2mp8PoGP0jh
yVB88bAxoQ80Ke2WeJVHf13FO9jDEELVcMzHU3tm5GkG15jTejsTQ1oaROOy5ct3OwnfEp7fGGsH
kOMnrZE6GkVQKuR3rcgAMiBXCz8qgtamAExET98R6mMwtgw0NvxxFSQaGyFybnGTjo2sW8OgCiYR
A5fL57Ef5Ibj/HIool/7bpFFpRbr5QJQnUwv+Ant+goohAV3rzvKzOMlLx2Dna7au8X/R29NbRvQ
gmmIYcY1/AzPAuhCKGDKZ5PkOuicLx+thVkW3NXsGGiD2GY15Nqt5AlmQDcn8jbbmgIvfLv9ThWq
hgg/4pSuPQzHvXfQDItxxDvSJeDoNxbiHO/azIMvLhu/ozK9yNHlecXRypB0k/SA2f/qVxkQtui9
DLjdC/NleAvVSRzkx1UaN+eVSDg3imcm7QDYDOkN/aUG+6PWLmC3cJVK7jUppzs2p1k1KaQDV6RF
jx3G9ny0iVxKe55XcIokN3G+y7+Y2uBaSqKcntfcfjmNAzjOD1rmMhQSFkp8A7ZWV1OheXtifl1N
G6dmKBd8bhmN1L97iFPXKX2Extrq5O26Z1/qXK219J7NvUb/HZtNQdK0MSzO0h30LoiVMyoo0Vpn
Mu/fGgBtCzodC1evZ9yBI9+AUJWdo8Mee3vcEOqe6kTsqXikpH1ayhvV+ZB20IWEbrXFaBJf2is2
WbK/em+PZcrbc6fZbK2ZrwyL8TsRVDKWj1xsXkfeB0EBlUUn0iQh0ev4WboE+7mjedFzw3HOx1jq
X9NsHtPifm63RAFmpgu+dd7L7YG7HbUoUV0C9r/JyOn4lf9uv7UjDb+xH9ZMd5BmJWmJAvpGaH5b
z+EeK3FxklFO8MjIg5/wNqou175Tsu3yay/qe1OLH0rruDt0l2P3rDBf9qkMGy7ESCYbLWGrTQUM
eYsPKxfb4DzpQvnPJeWi8motUNZky380fCW9E/u8vUzqEZuoAedkQPm9GKSMtTgSWXAkTv9sNDne
mc+BtzCHej3EvNqxCK/JIp1RCxnXtU72I9JTTYpucgGAG0m4d9/ek76xeeUOCROVwuFFbDzJryHa
7hXsQQ/Dyq96uxpXWW0J5x58eYJJhfD5AvGtHgPmAWI7/y8uUqNhrHNlM/Zx89Haa3nq7N9KeCDo
/CZy4O1VItCKeklQK4DJO7tOxwXFhhdxLMt2nYFNQXA6CgHjuthBK4QbHidfuAY8FQGosk8zD2Fh
Y9i66WV0TCILUbFz9go+PQXZeY8I6210VU/khKSO51sqBoxXDzUv0jDVDuIWQxKuaUF5SfxTtJ1T
HNh6PgYfPIbx0RbI0Nkex1O0Qez+kLh+5a6A16pUWVf31YRmNi++H7YhXg/wI8GD84idvWphx+/C
tR5cQ0CmW4ZyW4hF3dESq32ME9f3EcqtpzORFagSXeb4yBxlQqr01DiHzz4FN5eH0/qbLgg9aLC2
f6QwVFXVcxsjpEX1d4l3kvLl4GUCYc6a5/jMoVnhaebQUTx3yrKOg7039LIc18cfmQIJ9Fxh0P7h
yUcgIkVezzlPogRiBgurPpDrHTMgX5H81ssmPjhMZZf6EUTQFft39+n2xqZth7sVxqg5xRoTTQ1t
MV/AwhbUpOs5sM+NjMkl+Rg5o3KjBC9OfGaHn+QGqzzbJWNnp/UnioE0ksqaLRk3m8XvHxUXn22N
X7CHXK4M0LCfnEN+pTdDErhgTwSQaliN6yrKRLTBTwNnvDZ6nO/O0s7DXIe6cUQWNRc1aAwYZFo2
N0/PsKV1A6MAfObFiv6LcIp/Eweew2riAOkwvUEZofXJYCOv5+A1uQYylOE9LlPc9TXAJftOOSBB
fh+cAywNkgujPydgD6MkhRGfi6Tq/ZpK+XqOP0/fYJFvw1oJvzXsp37+KvWQ5M9Fr3JmpNj4J+LV
VameSkUf7X7fXG1ZK0V1O47Mh47g6RuO8m9yAnOLztagFb23YJw3Pqoth9nu7d4EdRCYyMvCeuxs
nYb2oNOImFJaWWJVGcPDdRPN1pPqDBdUzOWVx+DOBtZKNiZkjMY5dh87eLdYTXFXgervJeCb0aEw
tpFTxgdP60uJk68Fo6mKFRbLhZNlZRlAD0CQL6HmZwbiZUhUVRWrYON7upOcx8IxYuvvyaHDKfgO
R3UQMErzd7JTAYVb7FOkj7HUBiZ6RZCWbXDHDT8jaJTmKS7ez85B/QklDg0mhy3ze95ojBsgMw4B
tqrKahVSpCC7843ra/fMLuMIPOO97n29O+EsMg3Gva60RBWrc+Kg01VgyhSljn9uWi82yy7i0ohz
cT2YhZ3dRO6xn2IBg4oHibIJSGh+2n6BNETmR2KGR7Nf2FzWx7c+gb4EXqfsAA30Jem6QoFWBsd+
Dm3RugJdVzYnXgfhI98+HKzSIai+FGuaNRqjPOyBFIwJ8XtMBu6Q4JxB7njwac2HAix9sphQ6p8z
GXqK3OQWMHPVYK7jddvWx58WnpG63WBBliTQdyv9vN9WYh4XAm1rv/1Wk5LdklqQdjDv1P+GG+Oo
9ux9+MHeoKOXhGApiymZnlXbh02O62mPW8c9tdSWSYpzA8acGgmOuDGHvvszB2M3XSXed5JKuLEc
A0QJA5GKFLdQneFzIKgM0l8WI1lXQvdJ4lUX9EyPC0Yd+8xhBCScc8Ofcvc/K31Kkg8N7b4II1Nx
/tO6f7s2fes24yHhVo2i9kUGXoVJUt0R/sRqitBKrtG32o6oSlZAQD4o0KfB5wl0vEvnXlXhU3cI
q6nG+8LtgOz2YRSUjHsdSOrQIobXtwBAWwbr7b6E+RmWUcUoc0yHiEm7pXMzxZ5mIQsIgtSI1ui8
3dsZwHmP2FrhX20N30N8VchODbwOZaFj3KgJ7qCGjQ87FzzCZYF/JEOsihBj1ZQr7Efz4C2eik1G
pdkIeioIfaFfylp6PLnB+AOJx3vM/EEVHkphHLfvp4caRXG4F4ca33vNOwOERVEy8eLUZ4kc/ic5
RTQS/4TJVhm3nUxmxw20GChJ1mQTwIxq/pWA40Ff+fFAnAubeIDxid33Cm2uS5katX8xhy7NoK5R
yRLs9SDaiAHTNe4L4KU038ZkvkpSKj25ePGAsTN0ttQdqaME9iiTaIoe6+UgKPashfnfBc8fS7Dj
+G+NRLMy9ZMCxIEKXkifndXfKSiD5sZ/MAH0FBr9DCV12L/A0us7f+vgOt8j29e80yJWm5Qq/wNl
C+QyZI1oy8+Ah4aZKUU28HtCm5OvugQ2NWWU7I25lrmDQOgAGNYqt45bVAMZDykF1YUAPAY4RHGT
zJV+vMP0EYl+VHGOg6NZ5l2p28hekRp/rsTlc31JvuyEDJoLUozD0DsXjUQQye0Z/SWwNE7XK6nN
Y370qWB/N5WjU7sKw23weDqNNVm1Nnvg5NYaoVo4KkiYHkEuBXDVX6SIGY3R0t1DduhEE6q/1HtE
3BOto8h2bEWDBfLFwlhh6YTb+61EPS1iiyFScKW1DdzYZ7IkO976TopblYOqB+sU7ad0lDFRKNAi
AyP/3qI9jBvN5Easka3/jEhZb1mhN+CselFOvXTbIFubvkkkPKxkL0b3Uv3/K6UqrTWyWmPJk9ln
X2wa4kO6lC6DPwNuZEN0Q7AIRvo4LoLSynnbFU21hrZes81vn1fM1AnUFFM31otrrV33ZF8/MAto
x4narkyPc/Broto8gaauf/ZEnEsklfehe2Mjq9j4WBe2wfagxtm9S38YgkAgp2evgHDgj72+bFwK
85uPmuIrx82Nsejft0T7wta2Uk6jyHxqP1W+nBHrgrLHtqKSbrE1qCQhH8ZTsyQb3TM1ATCdclN1
BqZexY21S/V9oOmuMbKPw8rxhqJ1XsVjwGZ+FrF6M3ISK7lwm7s6WB2s1/iA4XXqhqyI2KO+4bxP
e9VQkKyVuPt1GOt0mzwcTl9QiGIMlFqouKyBuH0sfO1tF/YLUDVcU9splxClAP85EzVCsW+hbj0m
NsufztK9SUYQEF/ifU2fSzsMWUUlcx2YOGBZ9jTpvHM9vMh5TYevzsXoFSyIvPrHZFHmmOvKqY4E
YhF7RmxH13DwqH+qliyYjjbch3Z2hNNNpMmvp3a5prhKyMWv62xPhldY80PDJk2Np0A8eDC9MUUV
12MCQGtklqmzYqLbNKOJc9bLLs8QGqNZurpIEm9DhZDaTdvw61NLmKg2ed1sziQAjkhywUHJrDT8
G67RveyuZ/GTz2egQbByFlk5M3Kvd0jRfbtW5G5uFX4EDtHPgNR2o5k9FYhcX0CKrA0ktcIp8Cn+
lMUWEhijhWYAzhAK9MSvGXo7iQrmPGxwMfv7LuOmq70ZrBFg7/g1tSrqu9+PH7A48JOsNpPGr9TB
SGRRqMSQGgatjib6X7b0PaO/BXpwcWdSose2XNnIf2Vk5yOjhELGDpdJLsm2NspKl1VadnVkyXdV
+pSYyBay671/Kms/cz7Seiug0A+lo0cAs8fQxdIpfrEcN3XUovrb5jCkmY6lHVebMhEE7LvRDF6q
82j8ukBTyiTI5S9M6i8rPnojRGVCDQhj+/ygauDExwIM2/vorhqqtXavTe61WL2XSBcSkQzUpSax
VrCydFp51ZOJxhjCOqhjpPJSCy38KR39aM2nOIfhnEvDxsM9sWzJ4CL4mlH8aksG/zDAyXkeLaXM
1MWwlRrPj+mg4jOY7It/wzC0BEGascVuKRylFbzptxo+tHGbU+2EQSvDj+uBT+/Dg/SeeGVEb82Q
wQjWs64PjJwoQWRjUErdwQxuOt5EqbJ5GjGFDX7Wmt+UEUb/jEAHiGk2WlHsO+jSyl9B46xaZJCz
1Ef+UTBwOL83/oqkEHdT/a0CCE567aZZVBbl8z7fL+O5ugwN5+Xrsubz6xPcszMsDfg1W0SwaPQ7
bA07ObsAnhGoR43Ay8SClZnGKolIvHDXpZPFFzNYJgEDWVYDt8IBkUFDwewC0hqqoPWXEkPPNa9O
37vZQLjUS2GI7tj3zr1ZL/Rs7E5H4GOw+3yfw9qocjAyjliuVMPW1jZQ4syT7w0sVkV3W+d1Gkje
LIjksa/p5Bxod+Vo3wq5Ijm/7HZvdLo2Yzx9bDvnRtQCiMOz6HTnBLA2pTW7xeNsjoIzxF2HSJm0
6bkh2y8KdlM7LJBuVzjFsxjj0GRInBy+ocLX5KJG/6noPLBh6pVwEhce519lk9cC02Qqd+fsSJVc
BDpG/azi7VUdnieI7ym3ZnehkBqd7zhsUTZYvMxvehUqDteqXtdyKSMRRep9cwinAe+9T8a89V0P
c334dCy507mtMi5ar2HS52z3dbkmIDCee8W8ks4wMCecQ6L3Hdg9lI1+q9hmvPQrqlTfYoLxQEMe
n0KE7q80gZWLPj/i5EyYA9vnDk93df9kNz7u4jmcln4oOofV70miutDowCk3PxQ3UdxX0k+EG7xT
eqKWs0ar3rigkSSmZUDWKPnvkdV5F62frUhEm2U5RUnEmyCMp1LffTEDoj8ucNepUrqFR9uZ7D5p
uzlvIGUj96nNnsTQDaIZfH3LhBTvp63s1Mp7QAzff27ltitGSwNmJhaENJalA4z7NgTwI0d8Hu02
QmM7sM+4Z8vWYqVS+O7ZNBgEwdAF715j7hgAzSe3UPXyE+zrM7I3fDyWflo5oqR9jfA1s1bZ08Vj
pE5S+R0v0eQqMJBeSBUrmkmnYvk03HkvUvTs7ndIEvXJNGLYXy2Hi/jY5eB5gdil65YGdArFbQkV
1dV97KKrJyk3U9lC0aGijFGesPenubOXOblStDlZQn2f5pWltJF/ARg4OMYIHeuIZ3YISHO3nTYp
DnFINJZJsNpFwN+3IUV52IXOJbnWUEguC10JdoegJfI9Bv93Yk0R3KcsT+XjNHsksP6WjypZDUPd
Yc+e7tYGmQhBpERsLXuUK9phb0z4FB71izBTg7/i+IsK9W67b1cdiSM98/10J90I3AU2NbfS2LhU
d9UbTmznuQkCSARZuCH2P94DilTI1Ohe6cYBX4MxnAkQPvCBxAA1l91zWZWtQtXhf0xLr4Ea6Nqv
QHjTXKi7W31vCMFdqFZzI/7w/ixUcY+vZAVTdedLPRYCNu+X89A5M1BV/7UHBKUo/Bx9boJ6UmlB
lhs2XIfdYxPLJRYnSsBtKxVhkIu0J5RSxBqBpsI8yTccLjo/LuN3C1u88MBeP24Dy6uVExpywdna
5dYDTbC0p9N9nLTC/TRumrl9FDvdjvU/Ap3dgfPTYnWRCASm/ihrZIRA9EIm4pS3bxx9b8pI+vw2
gXyuAss/caKzWDr8ZPNW988lDo3hrudzNb/kBdnjPRlxGkMPrrdVU1II9p3epcKQ765wYyMsP++/
QGWik5WjU51oHI/lErKf0rIwcp6KXIuzbNhEe3QDNulywqufUBthfOIUTca/RV72xTeks14fornf
6QhMgY7Wlx5jSCKxowWZGzOTX8oVWYbmURPzHmve8HMBn1TyAdpNmhXYeJM6K/UZ4EDKBI7GgQ1M
rXYnpFU2Dc7TeCbMeOw+C+a+N9xOs4gPsWXzwO7KFQ69FllFBtW/nYvyI53Tr9oAf2vO+L+ctYCE
zR74q34UxYKiDtFJi57vM3/Azc4ykn0XguuqzWHtl4sBXW1I3jptruxBJAirDRq17IBD6nciidvB
xNSZLsMvv7fhQ2YKhIk3l/SELJ3i8ZR0GwGZ1hDB5zSJtPZvFiZ26NXjDhnh0/USEBh+JjSE8od3
nL/Vhr8klx+tAP1oOY1hVouG8Ekfq5WRTiNPfWuKxUl/N0KmVZ2PgnnnKLAvmQ7sbi9inFMQ7pF8
bR6RFPK97pUgrUtXYgzZfYeFoZjnIEE6o1X7m/UlXPK7xF8BXpU11D9ZsLYlADRl250iS57piyrI
7UxsNrLJ4VuxC1q7639erLRn1du8tbyNDHLFJ8B2u4+UvIJ2kdNy/U8Zn69qbN2n1qkH530dD+dM
a9lTV+bqoGUh0nDXedExD9eb3jFgJSn2/rhJRlRxEtF0S1c1kYk2yE6cPtuvc2uL9Ml4GV7T3+SW
3h5QmXoT9X+p9Kv03wGqH/9lxG/jTQZd9Y4YBZm9tCYl7sOwV0ayouJFUqXQdFt2Kp7sPhu3jkrs
dCnss9bJpTEOMuC1uTgLNAVCFS11ga1PTnRCQK4TLJfx4uzrYGsC0ArxfSrwHrAutfML9z9gdOSi
HQV7PwLS5EJ3BrKbVbBPym7sfgXcYhZFbYGydlDWtetfqkFdq5ufD/r9Ec80XMIVJfksaohGukxO
rWOY/YAYyjDbem6FrUmk4zzecF+3UDVzdGamfT+Z5aSEpqlgLkyuihqBsSPdJFEhO6kNb04LuTsz
L3NQZP3+GHcI4l0VMEom4u66Rl/ZbvuTdi6vx2CltIv1Lepo/0+YEs66/eGFJBCTUhiKWnD3Lm7r
IWhkPKnGBcNp09xhmzNrlZ4duU2hT0UJQAnd/YeQyVJRjuPWJRjSi0CuYL4JAbl3eIq5iKi98osE
aSSEpw7JwCYWB/ku7bVM6ltfQnoNEGFgKzTLiA0jkVMGuw2K8lWZQ4X+75SfMB/DTjxpHGLWd/NR
jcBK0D1rBigcbM4nq0I3fUjv0Y1XuIFnlxkGkyN/KroazoFodnSaYqhkWOj66cg2fKSYL2nhyFPZ
Leo4S+czP1L1mf1sMn/sk/Jn+s3JauYN2+2f2rii201KobsQJ86cdgSbXwUfkwmyOYFX89Vyl9xc
QRwvTwJ6bP52J9ZGGeIov+D7eGfdNcXs+4umjhA4H58XF9HH8mKCP0pDPeghQi1Q30Pz9mzvC8/f
9xNlUcFl65DbUV2xwcTIA3RMjsZog/v5pBjEiLbHGWTlElWYFk8oyYP3w26III2yUU/e4nTGQvXq
XIhAVArSRj+6S94GVZRj+bDML+8Aid+r2cbvapNZR/UQmEW89kMe+eTU9vSiIhheXuKvs65l0VKa
lKSjcj23fN46lCm6zAQV9leBhy6azAPvrM8VwhceI31fDkERqNHlui1nNShLCg02FIds1FqPjVj5
79SxJWeIo2P+wvnlr5zRlG1lsft4G4QKOG22PstudyUxKZ0vBup7RW/O6O29VYeukPggHqRuXfuE
MZMMe8QqBRz62tU1bpTB27FHgHhviHI0ccU8IxFzJhB2u8QyTyxSfRImHWVC6gA5w7+LUbLP0AHl
V72nUseJqDKK2umqWnfIGpy5P2vbyalKCsabcqw4HguKyJ+xBaV3q+oj5Z/0YkkHjotVJkQJVuAg
NxF1uKGxfGcm7+rqeUP5JTGWqBjmsjgEh4Fq0YWV3wHv8Dbo+vEqVLbauDKQysKkdCXGdHbInUWe
AyB6WWQ4Zi9H6XHwXVCzvuZHyuYgNR68opd/qiSKvxwFKQRWq6M4uq9d2xw5EdKgdrdTJi+FyShU
swSDU9zno2Vuklk6SSMEUplxKYwni9Hm6LZ3nG3D3GkU98wik5zuzFSbXMG5sbe4nDLDMidkAEDt
nOnxc/um4fWznXLNmyXf5SaN9xkZouTaHJfTqHZSuVWGxRylR+l7OL2ZqAS1diMe0Bpcpbuf7yUR
9Q3WjBZJBR17VbsTj1uBUnkYGiBGK2l00A+IZEEwlUmvNa+Da3gP23DgG9B8MgnDphNlTLBtBa0M
hkIYsUOimQp3TY+Ktv1Azn5mPtgcHjVhjY7NFicBnKj+ldz1OaHZevelNxJjKHJZcYNWRgILFDO8
C+Jdfi8dDOIZFyHex16HJip6nwPh7SC7cEWMiUXpbuCLltVXTSG+4Z1olNH/mK196jdkegk2pJOP
PEEhZi06F7gz5gDcD41WmuS9VIo0e23VORb5Qh1ECZzErF/K0YvotlzHHLCjr8cyooLJJCjPt+Bs
iDVAp/Y3/b3upoxW7QSIAkWRnJGFZlFXzmJo7l7RPL/dtafzDqv+G3OW4QwmqpUZD0VGeFtyrzKi
h+4KBlYbri1BSL2Tw0TkJvyUVJp/v3lw7Vh7NIYUlGbbmdpTsHeH2XIYuQGD6/z1oyYR1LDzOZxu
WUfr76c1B6Ajp1fRbdAyatXfBCMaJcZRzHlDawy8Hve2/wxD40qaNEC2Bsu+i0AqRm/AQs7aDvPX
0Jl8LL6dFgYopJlf9U4ZCjq95iF44/1yON/0mQxP6irrnqfOPuZZWBag9X/pfVRW4iGDDOApKuMe
v7W59600QPlJhJ0fpyKRyfrunh2jals1YiFIQ4rN9o+ZUpRA2nbIPx+8sdKAnFwBHX2Aln9uM249
jFF2RbbZfVSLJoi322E2lTKKx2JGRBExiXnugfr8b4zpkooN4dUAynPoF3RQBGP9aryJ8LZ8+i7w
L6mXco0xLVxiITUer+2PwK1LGVfeyoxGpYJ25N9xnlSnp8Ho8gK83T9YWP1//nqj51sNUrdiP9Dz
CLjaD5Gu9uJxKHHD8oJgO0jrLtThRr+LOobTsMFSi7csF52Dmji5AhWv8wb6QWBPqngcKCCG8DVR
+CPCiOePtP1PJsjqdmT+i+uLeJBz8kg+v4Ufcxw6F5aVXVTTL+MkG/0Y2cbPWusYw9eAfJBzQLwZ
8gl6PySQeW0AxNrdiB2pdqFf/RPEM4Vcbg5vmkwdlj0I+cwdu5KBvIoMaMNrWJpesDMYbHbqnSYt
x7WqKnWs5RyoAbGIAqsuOInACl0MsiqU3ZK/yO2huA+Y88/G2qGrXz9sqTng8yIQ7udJdnxwX871
V2HdkWeSodqasMnE/jvTUEhgvTZsnjeNoWO/W78e+vB8Igxw0poDSJThocaPpbE2ct3nXotOp84w
yj9ZAtMDUZlgG8n0g12/+EG4Ah5xkmBXFikW0Ku52rrBj0tDWfVVwImGlyjS/sxR/5WS3UoHJWQ0
movZUHbtPeYBOumfRcSRyBFmn/i38YYH5yNiFTVx8Cj4UZ+Ba6+b4+fi+QhkF8ZhklhqN97FPSAa
RZBuODAWi//QNb8awGgIUhKOZSRvGK3kJWO7VFpw7q//uoVbD7NTMrfmnEEAc4Sc4gOJjpNVq+in
CmZMJggT8IgxCzB4+QhxFpwzeVjJqp9t6vrJzsGWeMisJrAZf9amPeuPinwGFvWi93pFvGnhYxCY
XYOSys3Rq4fiYFSozUU3C99ljHocu9L9f1QplQch/p2Y/k+8eZDenbVVzeTjcojov97Y0VKmiUyC
Jka5xR0Cbdm0LXx3ySmTC7Umtqa+kC1e0+cq9KRTrV1PIYw2ZvNIRjjdgVFfAuRSz8Zq3GTbCfke
iG48h/5C5CMoy3XWBDg2w+hFmlErulmhYk2PnDPgI7QUOCjRKiraMn3RT3NVc/7SuLJQqL221nyi
5clPqK2x0SZXsvrsvMHKGSeUyqRYI1UCAx12ueV5E3Z+7pdOq1aWxA2HswU6KF6UiSywKKqujVOm
SJKCTtKxCyVWc3xYQOwBw9OOVYivP//X88eEsAX2Xm8oAFCPUXAsfpW8WoGEKoOtE7ykMYAwJrtw
hGEdC2lkLPcuCpTiK8tbFWP/ccFptLMaSr4Qq8FKUazRAvj7TRIl917I3SdI9NjEnlFOFUA+pkSO
DPa3RpB0GtwF91hfSqI12ZOnMPovC91fVg2WNZmzu3v7gypZDEnxDZLpnqI+a8WZ6BRWrQAOY9WO
TrooMhP1hhpcItbeTQNRU5YhzA5Ghmcrvx72GzGZT78SvqH+OlgAHVQ7ZLpBHtqOzVTp67jOfjXg
DL2VFup4PLIz1wJpKlOiYiH/yoX0IgAsxhQmh6tAYZEmd8QYvvqXdBitT77d/2u62C0d4cJKtnPZ
xmx9QaCu9nB2k9zUhEOC2WI3ISKuKdY9NFzT+kczF1nyJtS11LIBiQ9o9P9KfNO03312mpQXa6F+
UHm5oyxJBuVqMAxUrlK88uxirXf/3Wf7cIqnYWwi+L/Q/XJ5ZnNZ/zzRAw3M88UCQBZTx10+yHLo
owMaxuKlFStY+sG/8NTowNF2j2wEQeyPdFEXC0yFLY15c7MKJDL4s5xy57NjtEJDbrAOWmhSpv1N
eLa3Jni7cPxzQaUMxOXQh85+4cKd1sx3fgd6G8y9CRFEGAVm9A2RgFe2oTvj+DT+2u6XXy+RuVCT
sMus9LDMM/wz1f2tNZOygRUfDOtENzP1nChOh2PnGSchk/xuxO4ojOYnDiaGZnjJrhabBVqddB2L
e0UDhDtYofsJkjhLWQgMOfteQBgS9oJ6ETMMj2WV25vDLcddU5n5ZvmCDVHihd7NW7b4Xyhdbbk7
lLzvf9XYRPrXGEYDFknfFfT9LdvFCS8Bx/hFsnnRBREVzJYp3Ac9xPAkOJv1Wbp6Xvf6FmU0ju0B
dMVkXD21gKp75MPVYP0egUUJj3cwrURSnxQ3eTiacpFokiVzb3PW0yue7E/cUvGvLZFROO8ErjPw
dEutje91/xLjY5TG7o+1E3k8K4cIrjGhk9iBxV9nhyMCz+JaxeW4lqm2uFbTQDkfnvqSPNBYiW4D
GLhz+Jqm6WQ9KDeOzrup4jXJw4uJrS0YnCuMg1IP7NozIT03LenOwRNU9a+TIg9K6NROmyK2FtYg
J9QBE0UKo0lrtbWCCFMUigTYJbXH091ViwxCqMPJWLbhpdmtCfCv9AS2T51nS/q0N9bGgBZf6D0M
tq+DTyvJxkwnoZPzWYFrb3AhHGntwzfhwqiwe9CIiIVmCMzRfkvLAakACP71exqNPlo/is+mt4nl
JuAPWaIjRmpHiWYnqogvhnqbEvGOl5AjFob/xWSa1sXHgia5GIaR6gR0xjPyOPH0EoVLRHDCBeTe
U43/9CzApXkGsPhRpGEa1tvGtX4eWHzu1NjNB+8waS5haVAHNsaONnKUncwBCPf8/SXlCGt9onTI
OG/e3gv//cLjClLwLkCtX2EAqBdhqUDtmBU6paFySk752L/NdfyKoIfSWwJlLCU6Uo5jUr6ersOA
g8A22HZOep1hzNf+BdRNx6Vco1jel/N8uBtJx9ve7BJyfdb0P5Mm4+zSrwyGT0HXMIA8DTzqxn57
kuXqpXAmoLqCiVkJwq56U4QGdVxDe2lR9Nk8Vd3K/nBlWpkezKuYwLemh4KbNXvEANwzMqR6TEGR
i9G9vEZ22GqVc/i2ugXVYi4d3RQvEz/b5HeAZ5FkH9WaJgsq128QrRibM7UUrTM5P0VhRbaXOnHf
eac+BRLqBX5edOAjwTNuxX9X7x6dTCEQj92qJDVHLB8DtZZuTRNe/GV317v9D6D75HTRzNzOW2lZ
Z9SJfd92vR6RlEfinR0qdT4Ek/WT0kCRgf0I76uZtroxBSFUXgM1KYlBZS5NnU8qJYHLgp6H77IT
ey2p6cCECQ7E8Hs9sn9h9f/XHodUFam6WndY3okLicIDIDT9bKWr9WKwv7Ace0cb9fb4fCuboToV
MxY9WVzzE28yl8O1CCGMssyXKCMKUBcEjiyzbXZTc7ENZBdjtO9uo/PAsvsKP1YdbwpADp7OQeYC
gbT/kPAXbhkpi48363NcLsw0LrMZqNPrinUUGgXvgmt7MOrok5cPfw/PFUx8gYJvkSJhR6fko+aV
BvC/tZ2JTuktKTctzM+PvDFPzVgpvX9XPkTrqNK0LuCW2NYg21VvDplf/Uv9WwjoDrqL5LmJ4JWX
BRorvHXP3UW/+2nSNpPmxtrl86q2vJJSqPbLovs+McRl4MJKBexZ6mNFnsE3OSHjBgWjj+BD2wgM
nwb9K0ms6n0WlxC6b2BzVWylnAqE0NB8jboz8tvthYwV7RyiXmcLCbtvNI/rF0INCRnhqn5HpiQ1
ml0IV4EgcBkCLKlOKpsXbAmARQ6LWNXz8cBVfqXmSwuZHTowOrn3v9alJhBam7Tj8e0tPwd+DN/+
L5PnfaXgf26JB+SPK2wRCdZUMzTdKuVilZJ43F1eSEx6Qwa3JuyYZxt6OarxC6KHUrpEA36+mh8V
k2RqypyHlm5oRbyujWz18PL+wB67T2z30aSpobA42kLEaR0oYQO3SYhW1uBdd1ZJ4z1v+I3EEziv
+pRwOazjQuZYJs34UOTw1j/4xrD37inouH1wNmPdgvW/mrDLEAYAxl6czEyvnszke8OktgwBovnK
HRBhBvEA4rqsyKX2fkN2JNfZols1aQMqhaYzyC2VlOIckMeUm5N3HB492KIsKQVl0yWm/fWMOqb9
E5KfI/R+YKZ+cNTPc1zvCee2cLUkAxhY8utffcQOgy2A0m2xDMpBKxJCuB26zv17gPMCmoti5IqL
B0BK9VVPe/eYuAD6FsntEI+cwp7GaN2LSw8urR/NILxdHnedA8UwRJjETzRVe4dWvAS7BVIBXEDf
nXL7SGZ9+F2T20c3ppUqYK1RtHU69y0QOwJtNmAuGiT7MfVd6eQpar3fNq2Se3gQqaCaHdpO12ud
tuIID0kqr9YLVqd3Ef/PYMJXYvbVC461/1esRc71zxma8GDW+bl5WgjaxZp/fiQFMGaRVWppRybG
NblgrfyKf50GwxnXQrWLj9zbn/9d+ktYrwmSDqN3iR2EcF42eBWTF8euCLc1rUOwAcIf/x80kbgo
tTealP9q5mzHTJWNigEAsJJfF11jpA3/U3J68DLpXZ/+Qfsec+n3F7/tRDUASqOy589IAzWhajKs
biYuAqJLBYuKFroMkC+mGhmUArB8XBkCI07CXa92Cb/KiiHLkonotMqVxSYGyZx32ofTTIdgVt+C
VvQ9az/Nyr0uekhFaBjPO3G77DnYbUnr4OuCdjsVvnQy4rQK4xI9PoMfYdKzeLCcElbx3EGHG+8Y
PWqy/ygyklHmgaj4rQslR+esVa18KADinQksPIjqSfMMjzS4sD3QLHc13rdgyVmDLQyUjBXQaSPd
Z4DH+bptPx+Z8ou4vCy3xWEn69emUsuySWuVpJfv/zW9GT1oYNS/CWgojP0pjQU+XuEi9XLe8XiB
Tojw8Nm3TGLYTn8bLUcVQFL54v7jHY4uoon0nqUIpgPJTE7SLZpUX0+jDvCthy0yR6eLwooJYDDN
nYaL0g/qIvmhRoWtuHiCnsiRp5K6cWssIVYRbv3g48UFY9dBcOw6KfjKN4hlc8LJYqwkhfwwVPGT
fCxng1O8oxDIvbxLD/WDzU4e6pfobM+H1JSQWQLv57R3a1VfHFYGpS3/4Sn6MByxZRTpP5iUV5rz
MMKnsp6EsPqVrQo+MYwBR3vyBPmVlND8vtQ22xfLbzeGS9uFPIU/mAvIC/AAmJX8nyV9qicT5EpV
iPSYv6bt7i8aGMzkNIYB9vaMzCtPeeByN4oVJihl/0bMlRynJhFU743N5W43FtOM39KRNvcrD7dz
1Fdh/23ppV0QEWfTpmlXjAYq9OVr/ODxeaB6sfrsMF0tawfoTIGbBL00PhdJ0zflJtBIfm6aoDru
d+W6DUV/8Gr1AqLpyOTMPfiktXsm8lVeAgLjiWU5QO4GhG+xyC2nMlD2xY3EDkupmTnf6K2zufqg
wA1YMtiBTha4l0OYRuTodjLDYpjCWAstMc4S1MWhQtqiPxtk4BSb2vATGS79JWMXmQRDW4/PEIKv
YzP9sNU+R9UO7WDo9g6Jh0X7LJMA6/nXnaZLcnMsEWlI2BKe3WUNV/qnWyMta1ZhTpVlo/1/17IX
K6MVZ37D78gGh0O8KsieHNZGlFTIviYif5XgHlaFIa5dzDybPgcuBAOP0teuXvjQRYWhFYAOggKR
qmIFzrbke6EHca/zyBBlMkNMhBMi91dTzP0zCUq8HOwKPWAqPDn4L0lWmCrrQfdf8Z8gOWx6H6d/
uHKQZoqxcZraguSGl7irq+7An3/mWHcphXygEoduS8+pqP6ZOY2U0qKw2sGQ5NL9I/Kr46uXW2CI
jaj+LsWOXPYoWUJZfgC65B+q+OKngEoSSA/6qfyTcn/5XAnFTi+WF3BJQZbTgmBjKU9hJNLcGFPX
hg/9qcrUZYE3mTT72N8jhtFynrtvR0gyBEMup7MNEyEFCxY2gMCv2qipwhXf9izk/rpLD39iaVDC
gxMNrO8LvYRNBUVdY8fZdteHRgoj7AiY+iQ4+oiDgLOWLEycAI+91rbYFzyGYCNlAgatP1deKQlQ
g2AJnn/+SHAAySxA4jfRtp5u9W6Zh9wNvtcx0s47FYh4+1QfP996413yIVg7JdAjs8wV8CW6XJuB
iNVSbjDnx4UESiu5ePM8kzsERYT/sHkOv6lPNQ5fILDzTjfrKY+ix/uPFby3ppOc5IR76yZtoVJM
FErQNzew7V3cEGA87MY3JxCuR6nYGkJJPhuwXTLHK+Gxd6YuVm0elMZyY8TiUvxtb2128ZJpstnY
y3+ebGitMickWIV/1ZcityD7Y5jdndXJi0kNmXVxQ1eGdfWDrpMUpQ1pr2HsmHX5cYUDRCaofGdH
LQtMJyP5hzwmVUVxE+Gcuw6xDnC9Dze7dWwOkwPTPj1WF6qIufIqm72SgomkNyfR+zT0reH0t9Jg
Y25Za40LfU1czIwDyJtNDfLWyYSbt44mEUs7bBR5zRTvLDDJBrjcrEmzGGSm7kZz75TiJFMYLJ1z
KhDg81s2/f45rzCcwJ+rxYa/o7odinAIUDA6pvcgwzN5K2cpLm/Vyo8Xjf2Q1s4wUO/AP4SkIZqh
x4YXxraMSBsmE0TdreF6wIH/FlBwwc8pqU1Ij+NovH5OV8yzAq2C9P0Ahe2gGlIpvbKKKkg0hPxG
AZbMU5vdd5YLy8eDXP13HrHNsQq2Kh8mkVJLlPRVTz6rIB/kt61FbuK63UUDyS536D2yXOWmej5x
BwXB7YIrCwTQc9+1jEuadGGwN3khqyZF2Z48G1erapglEL7fx+D9rgG7mEtYRf+1cVA7qqYykTuQ
Uqw4kh2ekEnIDc05CYXGyRh7C0Liw6+q9DOHbYCSXA95QNjpcERGwwOTHiMNUQce3686BOWMdpL0
ODUc4NW5B1XsxfeIBJOSsagjAFhhRYeNtg4l6V9fvTFD9FKtCT+KR8DNiRkL82wM6fDyJuF4KoYp
m4HKmZpk2lz9H/KXjILv6lGGa8OlGWqqN4fcIzz8t815xScjIpBVfl7djHPlxge4N6uzAw7UfM0k
dDsuhUmr6RS+akOsR7Lyj89nPesPgq/78tPOhm8zetQfMimlCKjv0G8fyNZeCq/skF/y/qqAbNYR
wfokmWZKi6dHtTQzK+ExwjSQd7beESQUcrDGuKNQ8di4CqA4EQboaRpYg8TLwAwPEqTWseZsSukM
R/wuptBml8aPC77M89cdgqMR9XMTlV4nZXOy2iX2RNdgNDR3P4BpfkMJQUfv6d8rtyl73XxdnxW2
+wu7PtfFqiFxSjNMI+Dut2Zqf1XQtDlM0j63guAWrFbllcKZRNXby6Zaeh/vZnp9IuWMvXzVJywc
HT95wVAEwBUqXmXx8+a9UrSwFeas2rQN8Dxd+0jpXTPqWjQ9eemyykPTRj/mgCd9xDrP7ONV8nr0
+OaZUqB8AO3Mosp9AzuFpDaNXsr+3va0vRPdgFDDzK3M+qLOgGTb4ysU7T2IZWMn58QOtf35QS0M
VfVhD9nWRYd9kZQEo3giU66L1WH7d3BXz6qcBWJhrfNst5tdq19dRTpHF2+jaKu+JmjzNIzGj23B
K75+hKNQsChxEA0i+xmZsyfByrqnmxWcdJ3EV1WErSECWxPHND5M1p4UgjM6aeepMrCtmr5kZn2o
YE4XJWUqDMN1vEBPIqmQ7MYy5zk9R0Ckp5yzfi/y41raQFFnx8lDFaUm8PabVeKfiRJYukBKwgbV
Pc1kTKmnO9YsW2SnpL4J2C5dP1mKnVmC7OMOF78gneOx6yt4BKSt1GLafJmCKt8DaLn0onUS3uTG
U+ZicqMXwAiUMwz2VlT3x7k2Ip9OQgYcdic7lqawR8652Flkcpwk5Ke72U/vmdpDGJRhtmW0Mcww
nako+irEfd3sQX68MiRFyGMzSjjngOPvTDIIgIK1zZfyMk34EnGuI2wftEH92jp8Bx29pIV1Y9cp
CASP0HBVGgzQHaU0ZR5mzxcDyV1R1+BSH7yZPjraUn4t7Q7WOwbFpTXfwA0iY3cqWFXtK9/p9kpq
x5QUJjOa9JexYf+MW1pmkeOlmBeT2MS1DqDJpxpdPBs9bP7MIhPDmIBeuXqssBww0i+Gwm7JLD1o
3NjAZtXmS2H/t6HReeku0RYO04N1xc+2QaugU4bcFS3g/UrtpmPZWH0lc2RLmLyLVXm/nuko5vI9
8H5OsRHGyc6xIoHsL2FaWX2H3PXLDDzTd33xQw5MGL+O1yk+FkfsSc9XEyQcemTY7thp9AuBfqu0
hWeNkSCfTCMGgfiITJOCHy9nn8BaC2fGFx9DiOIZuHiaU/J3jeihNkOdKrkQE55QkhONy2NI0sYn
qGM5kuzv6QSpQZSO4+ykP+HUGV9vCchyYH7XRWoASjck9NibrEIY0g/m57jvAA60kREpyxaao0e1
8799PxU5c0xGYAFx4Baa9+2UBUfKJh6VA7y+jJCmTFHEnLCoTLIqNpduD/ksUunc0alzcmv5C3ML
I0H7nirfKSqBQ5xMF5dpsXPgdU46B2wMNyJdMFSVzex7oKs+yjHgmi/IGGyn/5ediqhaj8GzcWD3
77wV+0IzckySIHp66GvCHryDR/EBsjSeE0Jb5wCjGuGXJCDaeDKJVQrxgiOZPl4Dzuokp/VJlNvo
hRHG1+jj++t82Uyc2YpuEI2NPZddaeMAmnYFDZF9efUgsxWGsM5JbpNnSTnR1XTGa3DoqodnMNAr
LNvsY3w+GGvW47ETz/sX1nZgL0eQVzhRhaeGCQLK6z98aRUkPqq9NVcxUJYsTFN4rzkI+yYK/pBx
tS6HDnGmEYA4Toh3EUjqbBPaC+4twSuowxzI880juYvubTV3LcJseLfxynFi/79yNHdmd7lgTW+y
Nn7JcRjOV59gssQ0Uy83pz+X+koL/nckw+768wyDjkCgQbN2qXlyogTs2Si+JvQfacn/xN/7dXMX
vLjrNg6LSv9c1frg6lhC6M08ydEz24BlomcqqT6vb8vUSgMqBmB99WUw5kOzIxUB7MfTPYeP8CsN
zHpO+tP4rzEgezj+xeIJZg4vuiuEL4+mnJdMYbwkgNLntb+JS8X2HGbxd4lbbNvVDS/kX23CYjz+
FUAE+kjrSFa4gdUg/pLHaY/bOatvlZQtVt2vwhkXGZWJf7g+utpfUf77Q/mpW8uUS5XlhL1hQ+Tg
DGHx1Q4tuApmmKoAorATX23WJ1ycuPpaHwRcKCSd3FClHYNSa8aX7gcbfhaJLKDfu631nGdvmTuG
dIbqK+1MIwisN3AJQk02xOkbPLMkFRpU9jkbGQJW88rV2r1oFhQLs17CTALq4Sat24jtJmniL9Sf
mF4m43F/3YwdkQNQktRiwKAxTuD06rbbsPKfdw1gf8VP0295rh7xf4O5CjikchIE1jKPUltG2L5u
VcQxO+HUEUN2gzBP271c+L0WyfrKUiOddoX7SBppVaTmRGYJaewr8Lk1zNhxucCq+4K1EFVCZZeL
BUdCUQlw5KCBpole612CWOH5FRqsAWuwou1dwabu+PuWt1LAWJxCe/lljZCUJL+wDeQEfuhSi33O
Akb/Dd4UaN/Y/rGzhsJGwDYKKD2GRTpfz8MjzukJDQ5sxnQvlCCtVJ/ab69ctuZXLrRxScvb3TF2
aaKQFluEhy6j6TgdTuZSAIV1zvy47egNyuvD/WjzIAtd9EUUpp0UFeC7tV+gdpdGAF6C99q5DlEh
eIZFbukweaX50WwlBvbg8OhZgDTDJx0Ow37x1KOvtaTyKin/2sI0OLwnZc6wG+EY00VL1YnAlSXF
YH6RiJwaOnCURyPngAU57rqpayk8lg2JCAVZhGAGRDaiEtGIVGxdxU8ZvLXMklP1GJSdTjuD+s8M
raXa6Flef3Fw0edRZnc7cQQCgX4/A9AgHelCB8ieh6dqF4cktjfs91Xe4foqTYQOrwmh58eRVY2z
6cQQRJH1b3XnO+dDwDLz+kE7pIAqID0z/m3MrWFo5NKgoKvIr+kRQ+DZn2gedFhuEobavHCmU0Lk
ImPqJWlXZbpAbKOsskZIAcbfu+hnWQ73JIu8rdkDdCMuSr6MbrHEKnPV8YQHJ5w/eolWJeCM6QH0
i80GClgwZ6gnJ4i5lK+NusPpHnJNA1QeVUedZ83d8pGu8irw0okaRo++zJKQNI2P/M6U4czWVMY/
//TNhLlUMIg2bkjU9sp5wN0O0j1cBTphwrXLLHxeuZol1OljL1cFlNS8WiMsE4ibptSNT+KG4asS
VS7F9Gec5oeq1HYXU67xws41uAUaWZa8jUk0kU5GKcucm2r5LAS+W2tvwbgFF8Woj4ivqTJu1uQe
njUMtxQTx/WiMTxfyP+pwTAUuRqJxatJ6aEyTLHijnjCEMgDOdHVhB8LD8y8Cg7QcNiNeedzXu/Z
DEeQqG4vZ2L6JjUxFlj5ktC5qApErVYgGCU5mBilWQKhR1RANewF+oPkVSabjc6+oiMwfbcCBh5g
B5rX6tFKvjcbht45BS/AG0NXGivvcjieXfxDQAlmvWtyJtg3xzkJNp/73PcriklxSgMZVpbrXF3y
kyZS0d99HstN69FBJIaTTjGqGeESQ5GvxOA28v83VV0q0Gq7SfYni78zeKUzlOGKGYztl6IkeBk/
yoHjggJY6IkKc0IUvI1TGlx5bMNgh2eisyTVDya1CGL5IgByuBw3Z5kOsQsukWCCWAHEJCeuYvsJ
sMQpeyKI3x5IoB1LTFAAa0t2LLldxAH80lMF/+u0QBsH/E+RgVXvDlEPxTj5mDZ3/aFYd6fPyWsf
1/nfkajrSf1GFPRgxQCJzBMmCBe3DKEm6D1jZDz9W03JBXm7FiWNshX0NAxdiKQFtnSYuoRr4sqK
WvZa2/6mnXmc6kLPKYvmQGp2M8cTqWUM2jjV70cS27G3ne8rH4rRgQ+y5ZgMpoJm/CbJpnHXp4GK
hmq5L99ENGRtOcWmdgQBlrEzzup6vRVrssGBfHKnFzZNDwxJzy/KbrIyxNJ3B3wFj9LZUyxAHlwP
GqBQC3gqZrVTOEaEuapH9L2E+nYUuFSFteBa1wWQ+eAu6h6pAxlaonJRCEjqfPG3ozvCSErb2vTb
ssNLGacFT9MDpnU8m/9iYgudROosFtlqm3tycr0PsRSgXcqZ9Fga6FjTdAlwVQuME8t4fIagXYpu
9wLti5iWnxGF3H9FBebuxH/DXtgYgcqcxDs+NxReVKpSWEQNLk8XJSa93dHQYJwztAIV67CzEQ4K
1rJ1r5JF2gWaBC1OYF4tCfOmWDLgeVJSx+zFO+lV5VXPGfYkBIROXZJZJ3HEmjtdgmx8UnnBUjRH
sIXaYLt0n3ngnNwPC9p14JLePwdgZOl3sz+LbD+WmgWtm+Fz4yBtjory3inTkvoCDT+e6PIBT8K6
wOHl+DD+DM1CHe7mKx95wIAPD+hoOAXJ4ADk/ckKV9xQfG4n1TDuz35ba+b1ZHf9JSlUINFMiyYi
SAEO5leDTt3Ri1cPR448owr5LaSu7rBcrhLTknMro3UBfpYSEwZjUsE80TuB1k3oK4RnGpSKTS7v
AYG2DwVXrNp81mGfz1L3IX2ynhUOz9jH9j4FfSCDmcFYaIjjGcpKAH/6s9tKGz9kQRHS2zTmX1HE
oxl+e0egYEhBJsCuQYpyMNX1z1rITxnYA3irEdnq+MsNNu2/j4omASUVtL7o9DfzsH5K7gnzGGK0
AomGs/NvatMprAgQULnXJ7H5E4iJX284fCPNQg5aI19UNKU4B0Y8RXqsyonh38880G41vyKK5Z+T
OrrfJ1qXW06TSUcoFiSJEKRAh4b9DEQglQzHRJTVxkN8W4FXNy+1eA1ehORF3R8xNcvRkQ3h14p+
LFCueZl8ADu7v+9J/v96beCSXvX1fIdEK7fl77VQQqL+aDPz8dp7UvanX9cjxRNBTgbDVlghq2Zm
yWdO6RE3AZpG38yku9ZtzIoXGPKhKJ493chRqutdOGlS4+STj3V4aHtKnnUoRPMW/R9OzTM28FT/
z9dc95RDKkyGwhDolOFMcT+yq1NcziE1wlGS6OhaeXlVPqwReNB7HocrmLkUOhxJtl8KJSkZ8s4y
gYuDCUDkuDmBBfcht/XMl+M5Z6PPB+2wsFzLLUMQJmWyOTi5a95R5vgy92S8324hZ7WOTj/dfFHx
e/gzQiGQ29OFboBngp3tL/iB+42QU5WfeOMwVsweiO+VGqHi9k7WIeFLAbHr/V59D6yZ9MYA7RMp
+bLe5YVwM+cCM8CYo7zu0A0nwRz4VFnpOewBhoyARA2e+XuDXP8ZyActyuHPgbR6qQ0Ljn93ll/u
jlBFLUY30ldu/uqFcaT9uOzSNhZzPfRISmLBSaBqoIWUdl5q3bs/F6v1V1MiazprD5+1i7Sudbdd
/wGzMt5/w1N5G0Hp6GjAR1kujy4yDD0jWCN+oIXZnyWljYd/6VsRiKFgEZP6ykbR8HBHkkYeTOhh
3Bt4grzRrPaAfgcEwu99pHxyLPVQqHNQGrwp/szTuvNapdXYRrk26aQd/hkA5QiZLBh1olUjQhwh
q1aL16qOedPQLaseWXDp4hPoXEcn4jKHfjJ1xpZENIE6VdMrdyFc91qF+d3/7GKlNRvBO+ELa00U
wSuCmuWBu12BVangdhVfg6I5X2FxcwBVAS6/RXsRXIh/SWXqW7YyLxPjfpF1Goqh3famrJ1Io7qf
W8SPkzIz+IxMzPJq6FZ8vZ0YYt6XUa3JOiColOqt/x+K7NfQqtJggffwUp1e2u3+ErLcHns+//p2
TV5DACbfsonZbb1RQfKxxqUYnRv+hW5ggf7tWnnZt0MD3LViM4jvrlAV2klDAhBbXjwYP7nH2JyF
HkLfBaONmK9in9Cw8O584Vj9eggixNwxeBFiFqiHLXfzz9Ka1ud2K5tZ8HqQ58lHkkLqhKEJibzZ
zMellEZUO0NW5645rqO72BRMn9R7ziNFZLY16x51G4Zle+4wxZzAJRTikcrJeh/QZYk+RQJF89H8
prdTLoGfsXsR8Ja6kgNrUEm2qytR5/X5+yIls2KwXrBFxVFg1tb90bBjUyYH/RZQ5NJ2tXOtCugs
g5hwaHaah3EWoaK95snJGDv6SoBxvi+YfstPEylG0CcGzNKpcMKc+jpJmYUpXFjlsP6fzwYc+GOO
VKcEPR9sKsFenBduT7IjlGRgDxIDKc9ZtADHOrE5hJ2y1VNxGQsLH0HVTTHtBZzi7KrJClcQzVAb
zIWbfhydQRqWA2g+zgTEkSzrUibTnDuFEnifAyFBNDbRt9IGg9YjJkDgJzmOFiu90yGjPBr1bIk8
T9QP64fMnc4ZVfW6ATb1rfwyAA9iNvLGp4dTjCHDtSE0i9/tg21f9NnFdyNBQmWVQwelp/Cq2Qji
EnecMddMmPt1BCVSMNhV4aoeUZR2UWcJNs4v38da5fy8fhHAn3myFHBXxwH/f1Fg8eMEtLYTj4hW
05PSpR20IZ+Nu1o55fgPMbGVlF8gp5dHsQgPFwBBjVMIy9i55k0C29bbSnZ0ZZ8+U3fSGaI0FF7q
pKAui5FiAC0VXcN2YKowG4WCvygeLxHkYIGK6O1xaH7c9lWgS6cHS4/NIomhzibDtfAeIXQdWjLa
hPjYecNlquyvi4HVn8XT3FN4R3flCrFZJSUrjUo5J5fIUNxHDBiLJk3n+Yq+7TbF8/xlmdVoxGxv
QLhzy7RqHizkKcjBkyn6JxYI3+WjpZDSczcwNvF+TYj+vRH8ts5K+blss5UXCYU7nRPVVnnD+kKJ
xgyJORBXrQQwM731yEXu1xXu/1OncVd1KiNJpxcsQJXRsNDAhE42d2edwkmRiIEDZiP3A88GTRGP
QjJhnQHhA98Iivy0u0m1LOdXzt3vb8ZtdRksBd5vbQq3WsKDQaF9FpUqkQg6icYZTTcNXDIbnIsj
7+CbFd9CFCPd/mkluVcZB/a/lYYbA6OCCNEqgZqgUhyzlLPzXJux1GYXvnLXEs7bEZSnVi/PSKBJ
cOPQFuhTTJjb722qK8WyxCg6gq+AuCl70nx8Lp5CC7AApOtJqWTSLbnGLqGcRweXhRlMfeM0uzhT
Og3J4OULv3fC0R4swt4zLBwKYZhJOUVJRmptgKL4GSEaJh/dgHqvTvnZrjN70aMc2GzNy1g6eI3I
96KAn3BM/IogNh7XM3iwsxhHh97FTrDYl7Lill3mRxGQRXbuhA+r3DDPzSAm5zbx03OPSzbb/AOG
BnEYYFbKiT+yLHBeTqm1OGWSJPW9ZpRAy4QR5yKE1LxwBIgoY/P2X0tKvXaUECFTupMeuVuI/XgG
5zsr8Rk8qFhT7ciBgqejZaOuFxevMdmZeoS6XrD8X+O0mNB3RX7y7Qe3il3f6/vNogiqssPk/hvB
G+5MFUXqmSMLC7HOv7CP2FZZoN9JbPMNuyQznHSeiQycDvSJjsPWnyZueHgSaoFCX7sLqA8ZYxev
KuNktdFMXhXvv3XCP2xcOc/AZSJJCk8966sDWyE2DEQDKaTUFO+jrKJ2e5g1IJV7uYcT8IpD9sgT
6E1gn1lvAtW8OkMo8/mK6vYffgbIp+EjcDwc/c0NCONFlpENsLHhUG9aYN0pq4so9H+YTuk8Fno8
Ks2hmu3urNOhBbCjs5u1hD+3sY7DrWGI+OYujkNG95e0GUZy67IOgwBbfwGqcFaauVepPUKxLABR
C4bkMihSBJvr2hERGzIgZIiVTpmE96WiYrkQUOfq5lNEQ1qexlkryGeezsKZ/X1nFsJR9O5w5+ow
JTZINKIclWbWJgMf8yqT48X5sAAqlpzNGUFqzGDs3WAWLNLDNgGIEBq4sKFRZRUSFZZNVZrR7OPb
leubHPF4BrJs/lfNrN7HS4inQyJ/GiFtrIlLwAAmbZjK6wBw44e1z7mE+hWZ6nUb1UqZ5R3+0PYC
h28KiayUXQbhOKq58KmQOIaV+2IzupBDtkbTkBd3Bo0tlakGMafql1U0pNB84Hw9RC+Mzk1Zjr8V
UixxrydddHnsOUEdRXQ0E9B6xefe7Ey53ISKHhnRb59eWUoYoT5hpou6AYRyfwkFoWuuLxHy9ar0
m+T/zdMHHeEnFc8PPKRN1Do1H/9qMxGK4yhrfmMQYyjevFXwAivd03ga//njoSVyPjzbhW4ocaLi
9avMRQ3caWvNJ7S9WtCYIxOgZ5ijGbnSKPc+IGpDJp6bWZQYaMF6+HXkTz4k79LJTQDAw3zs2qfa
FkPRAKkOnhlIEXdvwU5CvPBf9ONu2/c4EJhAfHqiO92biHHrN7EjgkUefwGEtzHnYiIYVyYx3Sql
cCYwD02kQAdtvzEhoeRU67KPuWpp41WugXHcSYe0SDKtzjseMjMdOoxwWWjGIZeLpNH4su8i7aTL
Y33DxMCnhibsEEKBgKXEgY0yCMAF/Jp0BNal84hK7bRA+xY92NVT9vf5/+2nIXqYj5hHHVORfwN7
cFOmAyXnGdEZd1ZEvY7xngxGgVelXog5u6ojoSPNo4Hb47NdFNAPKJwUoSzvZ4YRfnR4xe8BQWz5
1p2wmi4YAZqg1p2PTv80ycOAgzRJ9LuSTXVltTJ6YxiqSFrfa9M01fDVLPev7NjuRTCLvhcvMQh2
3O2bBVIX845QxUmXGAW/hOLtLZfl2iRsb/nDBdU2a5T5GaFCYazKM0nH7PkpdyxoIzdlKQPbgbqf
43Ikkm87GAaATyAO8dJYZXZA6V70fXzj7EQYKN3JHQEXrgPlDf4XtwKuNztNkWlo1jZIEPUL+KID
6JQxgOlNo/I9logwtGDHtUf93kBQpROZ8/W9DNVg+1oazk2LAqPRZHb6P/SEeEq3aM3zLe3OgZcz
hkP/J6DmSsZfhbBUXx0wBhMjaDVyIpxpV8y9wopGtneZJidYC7f6Rzyvw0J0yW/MrSG3pQxy1tyv
4ai1hi5Ls8xKj++kTUfe8dWGwL+XK1PglC7Zw1p73HfBqsR87S7fylci8kaZQ8anboP+2UohPHkO
Ruj4xURO4Obs/INOZMboCqP79CS1h2Dl/qt9ElVrggscskATMlCyeJfplLqV0Y5vV6axe26sX7yv
l6Lu4Jg15gTsk6dvRVailQmAxchOUgf8Ej98fjlWGiF9zkom3XNS1TbcGq5YAc/Qr0LHdNaV/rFr
CILq2b4Atnkgxv9Dmq/ccZIYH/i3aaanLvsGSey1a0UCuVRjvkSk9oUhW5wGyRd4CRjCv5xdHLRV
J1n9Um4X2G6JqX8lWS/IGUVJ5BUaR+6OfV5nIjNmSIKo39JmhHB3yYxJ26CbKoCR/7bAxTH0tYEY
b8Nty10Phg5q+V5OoBWCpanIh7bn/dRqOQqjI6XkR29nC/bojAYPd5MW8NVenJ3tJa0Ppd5zR2/U
U98IsiTEk18iVrFaPuSLkl6U+Mckld8Q4fWmko4yughW2xl1aDSk1PEZWOEczuUGGkjJKad6i0k9
H0x4vtDMhWbtKeLoJW5RbqmbLIiSDfQt0mKqL7ZVYLgni/kLsqUFJafFMdv/XOnSi1AwTeWxIk6e
/uQABcOMW9JhxFcu47bkkHe2ScLVlhpmZua3ds/m+8ULsNBx79VhMV1eDYgPzn3pS967MgnmWB45
w5IGDqTqubNRniUWgVVDOwUiU39Nq5pqQMwFESyqPuWgvGa+JPgz0yE04ldO0c7XDLhByhhNJyoD
KGOtbSIiCTsYEpttslXujVP4owXIutQ7C/JpMB3TgqYVhlmjEhOritC3AiJ9Wgu/x7r8TXGiL4cC
dgMwP0leoIm1fnceNNLyBC8foVBFByL360q+/6rxFLB8TpbIcYMocTM4SfeLUdqkvU3Lgkp8P/Ev
YHfsv9S+0I0E4wWu9OaJc9uKTo+iwjnc16ts6E0bP/HWNakkqNQnfsbldqUB+0stOdfaIvgmDFp8
YE+d8cAF6Ow556p9FQcurGLhvT/gAfr/Z1HCt7/bPdIFEYQ4kO/C9eRAzUtl44Lr+DUjB0nbF6wI
3Ye3Ak7PR9OdEqgJUGvvW9FAhzSqVTSmeRn107okiEx1p1EXCnJ9cS6YAC3BOq68jPaWizWZkJC4
MYZYNX1WuZw2hvS2vZa0cSPsV4g8geOAEltYrlhqnY+F/4XKbKzpeWjNS5mnCcMnelE8S6V5R7oz
6EfBk/emKFgjBYDKjh63qn5GyPBVh6NJtN8hxTu5VFJPRVqMiphTYMtDemymM1WbHhThP1dIRMC0
AIP5zUjs+GV9bfRA3PI5nIWB7L5H45lwIFqmyBh5c+CUfis2Ffsaw3gs/Q4ObgwTpK3tS+Lz7VUz
BG+GQXjfIYcYulbgG2scOWl072tbQdlaFyRXllH7kh3s6xfni2h19Jv6kavAYVW5PD1wKEHyiIoV
RZZ/JGC9uKoojtnv3bZmudFcZsCH3xqGoJ8WXnkoCrD9UJXd8c/mL0CrheJK6hOWJcZaEXx7hy+Y
QmXg2Xe/jw3yPACLo1ELr1xEndfQygCTknX+5TzXhBOlZy4uxttyUQ9D6kkpWLn6xv8rxylIlSNf
Bucm6pbgpCy/q0MQZ8J+IrnumEBoMQ+dXVOZMXbzvY9zaF6JdrBIkx4OotqY0q7i7DBIaySI98eR
gi2wYWS458Lcz+CAQ554/JDsUg8dKuXmda5c+N2WJO3rKBxTY6rOQ1ih+b340S+TNZmnnHWo+JuJ
gr14HaR6G04iffboNC84VTYo3xwuNlHuWFjarVSJKwT8HINFaG1ysjXtQanHizNalAFFDnWB4YJz
PzOm94RpdGMPtCB3h/XH0WKfq+73Cua7lCsZvIDhcJ28FG5qkUsxoCwujWuub7LPzi8Pb9lC0TS5
/JVcyKVAClCwAaTf8PjHs1MpSkHoLYOrX5rvF1EiNWqUM3O12AwzjrpOfeQ8kHakx/JUTwXXOo4i
84GQ8YsRzehZZq2ogWiFaU3i0/KE13aCEWaH3UJ5/oI/B3wj7Xj6H4wthqfuYgv6hatfthiJJqpF
fS+QXxhHEiY3wkMIInL91TKs+2uJssrYjS3GXBjZTX9jVvjVmXpYIl5Xb/zUSAJ/V+Jvr6RsMq39
DUKg0mYlEs70xhV5xHGqDUB+sxFiEYez+V6kLrk1iRhEOAtKW8PjcJ+otQlLoZ6pT+ZbyaJnZxcV
KQh6RwuNnl2UpJeIEUnnIRI5NHimWetY8Uv/Utchksb6kI05HmEKiJiwavJt5Q8cOl1i6ZSE6nWx
nr88Z/taowni+lNukc1KTETpBytfBebCUoKV5Ty03/roL5L3wzi5PEdJ7Sj2or+bBr5Ui8Zyklmi
Wt20/SlKw2cNaKUPOHPMaP2vqiHmSj+u4tM3yDGojErECs+7NvnHjH0ucupK8wcf9ql3VvSGguDD
Yf/lfGpSzH6+enbsVWLxJRNgwz1yUThs/MZNutwtqkI1qkCQ0YW45ZvWGof77DohodVbL0EZAsZt
1J0+N7P9J0Q0Vdog/S9iR8z0zddIdvxC/gcGPqEzzQ1x+XJTMvYbizFqeapY0wJfdGwELlyVvgg3
GkwcIKred9J94coFX+5bYK2cCvW4SXMwfL4ZQ97S/F+q2KBksxBM5FYOqJxP/lELt15iPyY09liR
CLX8MyPf4hJYccdp7Xu1HnNU7xcFKGr5wxAXlH2bwzqEl3wbov6pm/fDLZ3cqx3knnPbGHKwNs8N
j06clhh8YeiMnA1SRKpjPzr1wk2FCDPLr9ZRZ1hewnV/G25tRq89yj47Nqtm5aAAIw/wWMl1tdWZ
LidyUoYqwBZ5t037AHHhlumrS/TvNuTphgAkVSYQgutOFiu9E2KCFH02goGNVyWwGd2TImdJnUpm
XSVLwCYqRgMu2tIshHe5PPx7JBvU79j8xeCFS7lE3Os5rY0BsMzFIGHRzrcw454d0T7BN8SLx3CP
eCkpZbvJJpZYzD2eJmnRz4V3elCztv73m12PPPKKAH3o5fLVPazJaNXdz5iWEb3qRbw4bBJZML1l
EchozTmIWUADmagBxjJZ2Fea1rHuEW7Jv4GV1ES9ErPLDQ4GQPEjYmWpCGXrMeYQ2wkvlHQ6RUBe
1bY7PvtD9rTkxQy21TzbzwKcEzu35COa79c8avOJR0h5KmZke0TVQHavCGIjWJfamckMVMfV5vZ2
Mr+mXJQEn3CSqOHy8B4P1fGMhuKJ93aRtQZu5MLKBnL5OuE39agt86YKvyUI3Dv42xPFVONm+w/A
9HO30uH4Hckmt6rq+n5KkC2BesXwi1myK//0JQLDtIwRmgml7VLSt3/zaTap4LUotQ+YHjhP883d
IhmQsLREQQynvqeyVEd0Gd3x5GrIuZzbqcUUmI+3rpf3vAFnbpjWO7px2ecCN3KUIX7nVGTEcIp6
M2zY/WkZVCP+rpqpbywTukTnROfmRRdXeuUeVNXXpYryfAygsP7j6jVZs8zM6nmSDp442BEgpoeX
CFVpvdyvF0ZZq84dizM0Zf5NAEuCr8QpYA6NF5UyNrFSMFwrrLSEEr/A968bfUTmPMneicTdeytG
5UX4kqtk8y8V3NbAPh+ccvUHpALdNKC6JnlS5J2+jpZylYGKTUA+/hr/5ReYE8ybYOriZyE7xZLR
MFpodCMZBePKkDmcZnN4xYX5OnoPHc7uqafOVIMicitTsOkxnW3+5tjgtN5domH4B0Z+U/ysirzR
HBbfurmrzE0fAlNwxBZWclpvV4qKwSD7cd9GYHHTVKq0AD6XDrRfcBH5Mnyr35MZ0ue4dnXAFtOo
5hAgK3Fx70DdjYuZoCpe2R/QBjLH1vNP9ODt2CHirMJ/s9Z2xGshGyNARPUZLhQsnRSfAy+XR21O
s7K2iyWw6aQ17h0U5lCpZMVFfFXNBzsuQGbgUptD+A7kcNGHQsi+chtDJTbdTDqDRDj9UoxoHcne
NW6sw9m+ZMYGRcDkZv0saR6+NR+r+MYi9QdtpyWkG2tCvDQK89UjKIWFWS4W5wSx73aUQ8MpUycn
1tUhXjPwLroZcFuNwFl/bFUnsGytqfB2lyHblNi9yYqQRsYsPy4mlPoXMaJ1ab02EaKBreYD1Tq6
n47De6vBDGK3rcD54901nkNa+5BIw8fEfIJq1S54GW2PpkNVungCaERLysLZrKPdyfxJY1prOzRC
J8pKTNtH4tsI0lkJTCJxStudm8CLTTsvCgVKbaTWmPQtxwa9C94277wu7d1Hw4+jRB+imBUhkiFE
XBcZA7PTw2exVPEVxt7fCM+8RvKOp0OXqPpMxeEPj4vo0Csf7Ulp6QwxK6f2sjxcF/YenMQs12Zc
V8sUfkTHVspQBnKlUuzjEx0+W9BQlQX53rveS4XFSxxAdp//6I8ZwB/PkS3WIMiYIli9vnTERXBD
lmORsKjL5xyiBlTgnS2AXeJz3zNEsEV/+aTNnomIqUt30sA+pw1OpbCuiJ0OICcegsTyrryTLcBA
RNI2QDKX2XhXu/37A2ohbX7wXuBFhZuKLP3dhHjFUiKnG7lT6SF/5u3XD5og89XjU+m43RFThuDF
s5QStfyleIexc/LMxlTfJqRbDenp4EZUYfXR3udoPahVTqgMy/zv7Di9yMGq/JrXFxiD1RHByEg+
MA0T4RvD9+1c712kovJk+Ngi4BAvqtbQYdhuZnX2toRX8AvB/30zHvNqTifO0hkRbOJfo0RiKCkb
KKtoeTtv6+kjEqe9MnzJylIFuqF+oR4W02nEaE25fis7d4eMN9FgJ4XGxdlwZjVdW1An9NIDW89V
y0slP7Og9QcNNZyg8hxTDymkhPRrkShosBM+xSvuQ2oNPhgVMZo5R4p6ukeHy2iYxRJlma03kgew
L88HXcxLzgnBqc13eAGBZuYcVw5Bt801jogmx0M4LuPc0eDAc/hyzn+bocDa6F4jeS0fcABsbLyx
q5GutqBlu6PN0ySjXzcVL2j+VFZDr2gybhKLZpuFn4LboFJPjhZyVRISB9mgCnnxgXAcs5c8AfGT
L2I7powgQBoyu/OcjGO86mDgApc/ZdTzpMya7IEcNqP9gHX0PBSo/lJo3pjOKP2xQH8PHltm5/vR
oEcErk9O0gb4dCrW0ZHZXMoU88LtR46B1EpGGoaBI6PsTYW3vin+cyancSrV+M2WUwdvx9hCYTHd
R6tcQ3RCXs/P5bQXcnyTexeypczuqITG4dZj0Ia5qI1sfOVMmhwOX0oSCTQmiq2bX174Xgp91Wcr
jLTnBQ2YsiDjRJIeuGB0QiCMyDBR7KOMToCK5V/NjS6c1o7p1Cy76SYQGVtjID6M6zYUNl3gn6+v
bl0I1Ot7rnuxCvyghcUQFhMKosRyY1trKiYHrp77UP3/zws4TbP+WkvVP/uSxuRrqpEs+Pv0evSn
s1ck4Fl+FbgGoSHPrXTpUin4XaefkiYsAu+pm3cTHVBKSq60CHpHRAmuk2zzqS5YMeBqXE2yqYQZ
rnioHhYnh78J8TB03ddOuxeadXEHusL5xSBZ6r99tzGY9kki9j3ErSzZkFpoigiF0fohWvCMqmVy
uUPLGbONhfGi9Ks1f/KvxCeXFuYTsz77G7yA4Ox0tXHD2XcyvdRNjZ8GU0V7gzXpoN1GUsBAjj9x
vX9KNQTQm6DT8+mY17vi0TKOCLz2HAT4hU1tYfFA9RjjMrX+luNQ1cMQUWB2jAcLBM8n5pzobIEA
Xqs8W+DIMc9Ns39DlF8Cm2C7pjW++wk4c9KSU4LzNlKHQ+KgvU8ow1IW3tTlxY+gD/ADNBZdxPhI
M5sW4MvmH3Uuuzynfzv4rlE4/m2jyN8grTWUtQk/nk4Mp918h62RpCMLH2mD6r95R/Y77HJiDBDh
LrBr6QuDQ6ISH6Ho8Sv0R8dKDuMfHzUwj7PIklfMTmsV37JSR35jlHCWFQ0+C1S+7Z/pF9eJibqG
cX6cZ1u0nMjD3ygZJ+BVeb81GmmSkDyPQJ5GQEhcDDPFMERHaAZbv8qTnzSQ40Z81pw76A+/PbHg
IeYenSJG+YGVh9aJr5ltN7hwzj2LUwWDumnbEbDXwfS5lcaqxsReXrC8nbPRwvj3VzuXMnl99EMY
HOasDsu2l6MZun78fhMliryTaAgHdNCukYpe2BONAfRu/DZ5QonQ8Dytn5Corwy9wyovKHzdAJdl
KHdD7jhrbQVRhRwHCT5aoiIlNSRbxQLeAV0sdfegwp3ZERMoqJSNduVZFHG6e51zBs2CrwH5zowI
1T5fqAXT1SN5roGSaZFN54qH4gkAumUsFr1ylw5a0grlu1DjBYFeGYwcVqUMl0XPcPHp2Q9K/E+7
CjCMuxWcsgr9hVyhb8pPuei6HpJqQ46QCy48qrA/HDcgrSlJ+RYeA33BOcBhcFvR9Nsp2BtVT/Qg
Ahf4Yy5fiChDT/5SYuRuzDWXAWozCo2o7YVdVas0DvvjyXb424TmO3kxJ1qkmxIDZMWbYqnR4zDf
4jq7vB/66i2XASsi+Aqu3LA9+XDKCio4dZuFbgXCTnMO3Fj+NTXTk3IwqOdpYlSd55cMEwQWGugB
MKgPS/pf7bMCzhZutFe6ym6/mvB+rKfT47+oI9e1EJ96Mo/HdA9QQig99ZDl4iVTSTCHBb4aFIBl
2TuStBn6aEQHWYlth9S/wUIk5fQ5RF13ERVnjCEFnBXZZpObhISpntXGJPJdh/qkCfYrvVBmHKMm
ILJUf0c7x4dubQPC6tIMfYmw0EwEfz/bkCYMEl5JaOlMLE/FBm/pexUel+Qd3s9dxr3bOBNcr2M2
5+y3MEAfjsmOd3JH14cy0EH0scNu3mBZwWU3JuSS9zdphGtRTp9a81guascA/cSDGciy5wEjtI4K
XN4n+ua6TR8wDqNSAlHtTg/5u4oLtNnBiq4NA0WHO2n1Xx3hujYn3UX+xMYTJjm05ROukgDfHI0w
bu9lw4QwiYVPjCTNw38So/5zJ2zAM4pkbE20PY30fGKaYyMJznilPmw4wPbCAAoBMZmeXjhZIj0E
P5u55vRmBwpoaqnaF5xHgTSANtDBFe0kchdF727QFpxWOhUjW/f6xAAhZElVZd+mzNnE6XkoLwM7
jgpkhRmjYFgpVB0fIdTURhFUezFyjPem6PUdqRczj/k7LOz9cvxp+DcdhOfXownFNBgfAhCsLZSW
kP6WKLKE3wlrTqtDRI2tvtr9vh0sRyXP3R6Miu14sJ6T9+Q47wiS9EBFi1bfpU++U9UQXoMcmrx0
wITqPcY1USEmzNDQUPEVWtngzgdmd59oSQ84B4/1ttfmXOUkeQ62XCjJOXYFzUIzgyIpczPdSJ0j
zqRUBqvh8OGfhd/xuGWL/7OCY7d7jpk9pMd3wT9iNSg5/QMFTWbNVp9W5spwBnh9Gco+fo5DVCgP
yIJvldg+ERqFS9VuW15P2IMzf+V8H081rH8ZX2oazj5xdQqLvcezLE1mPyQhSfSiSWnXAnXndPqp
EcANqM1UXfJKT4sqekw1SjBumPJSi36iUf+7LFLAr/odggRWAcMqT8gd6MDFIyBmScSjuTIK1Dbe
dZ9D7t0GnV0XfeuwHX4+9DyvDl0UdEDwnFLPhHD/7o1axllV+0XV4/8oJ0E3PrQhy5VQ/fWn+s3a
lj2Vlb+nPvlQDj2pMrnrEdsVVCT/xPEZAzLWu/p//nNrthyfEBTd2KrFreIt6/fHjLOfJ0OBPrvK
c0gr6eQgOl4m0c5sjOsOidJOxnvw9CsIU+3J6HkkCfcgpus6+/w4yp9aUb+Llkdwh+h7whfOcLA6
hjUDvmjCgCa2pHC8MreOJsunQUO2DEHkOy3+1rJKZko1UDoW22n5+5csF3gCu9C+H1eLoEDV4SA3
lpB1pYcKzfIx7SwOpNdFx+OLHyVh2xP66TYGedrAEoqvF8IIk7GKxApMdlcr4H6Z3HxeaTAuh8nR
Kp8sKBcOPH+xoxLVzHStiIha+IY2Q700sWRQFiKLntBF0AUwQQ91jozH0mvQlcTptqwW/EZVgm3h
qUwgm8Q7wTk5JieofNf8HO5nEQoGo9oUy60QY6XCbUpJScjbkGzZUJ+SqzBew90oh8EXYgPEHQBW
o/D5emthuF61zS4uC8DK2VSS1qj4JnrfyBaIXQHuCzdHUD0dLuXZMZ+9n8JKi8apuJNxYIwebxK8
FjmkrRyuqL88IgvMNGEo3Ybcfvw5pZmJLXY7+s8ufx5sevYwjozLsNx6+hMl2V73Fp0Mr/7yL4P3
9VmCcCRu8lyujpauaTT/ac1hHIIWHCC1G3t1tqepF36tDItjNcWsgR0j6Xhk2uZQ6fEwqjX8Gvef
rZ4jsysLXY5Z86FtHGrknRyK2+9HNqfb7xbef/AjS20CmPx80BZUN3+qUlEb5U+/6fG6vuI9QZWH
WHD0c/5T2DYG6oEA0vYLmKF69QMBwh+VdV34t8I1NXLLiyW/hGpvzTdsXYNLdlXWE2mqYUo3JNRZ
ERry+5Mv2eSSv58XVldGuILxjIQy/b9QIE1voosgxleqlr0ulrB6MRQPdQWCB9R8mjrV+qh0tJ+P
/dfzLQuXlPIb33gQr5GHqJjc79bwiplRbBzHHrDT8QOtHsP6MNnbbO4ihffl16VeHSSdSenZp2TC
poMT42nlu1BocKspiaiPDkkhJY0VUULwXUZpwWeumBGTN5772/enT50KawmxUp0zxxWXIRiNOU0V
4/xovb4/rIx/gMa5hsbxv29Xzjeb6XCiWzZrDCKNbeVO5FqhWYA9TQ3aSwFMENBU2wek1F2dh5Wj
N+r2RJH5lz2STSWRnU1mlXUkKGxEEF0IARAlYPrbrgufF7wckFOaI10O0MXB3n8KfQQDTUAOWNFx
zXdCLpkfP2e+Yn7wRZJlo1250bwL7a/D4SDwUCpRtuv3Nqp6h3M77RUYms6ByTwXP86jZxx/LM9k
jZSdn9C62po+vM1aAOeQsHzVAQpUALN3M6Rkbc5onfR8zZogzd/IYjZDR7vZq/Lkq7IwlqcCywBB
Do6SFS34KqOirnrsa2Bvd81VetWmGCOBmMbTJpKcCbQkegfhaqO3vHvXLdmmzDfQSrNakks2DDhP
k5Yi6GeV4/Kir25Uyhcfbp8g1W83YtMpu0U8dPHZt3cu/s+4RRfUr20V5Xpw/msgtto/KeOYK089
cgl8r5yn1/SC1yLAKILGktemZdlgil47e9mcYKZ8FD7rXlstH1I9gJyHSph/hyfGSzBuJyS+IIt8
pS48jzyEkgB9eU+Y+DzVhaAJzCFw1vPDm+Wx/4XLSnUGdYfOWy4amwB+PcIYXFzavI4QlFuEEUvG
RIq0zRQdF5pZ+FqTj/48lSnfo9L8VuLr63nh2DRJXVZk7pPM9/m0xThvsQBv6Nj3cwGzoVpRSqt+
6yXgx0n6B/pjWL+dKcAU4lYy+ED2pdJDP+NQMAlodl2sSgR22gqNILzWfuiKRWHwx6hoKIhieAzf
WovscJj9eFlkTt79g6KwrpGsZ9uG1QZUhYUxnizWcDI5GO+xGtB6ZuuZi8KPtb1tFkttqSO46a5o
UhoxOl2bb0SCmdqbjs9ewiguNpVAGBJYBX65u1RDrK/SXpmuPQhTqXz/POFZJbgOo52SZKglJjnx
rcL67Vnm94OKpRqlmoHdAW2dyk53d29sPdCxp9f6D3MBEFd5VkXYgfuTNIhB5XfapJbhxBEXgsgH
yuKTBOVeu7Kp7lmYGwXajNp5AezQ+EmZ54OLauVJpPCkN1o3BF/PSgUroTGRWzltid9cu36WHbRM
QcmvBp5I+3UZ/O694fX0F9xRowu3Q9voOBRhGqtomPW0O7Hsz0LmFCy8RWz0MCp1+yWKJCNQfnB2
or1txXEJ15ALwdUM81cWpL3XmTsgw5PqUyoay1wuYuETGQ9RY/W0M2p91P5QgvrwLuM7qzQ0G+6C
gmgZo+t1hszbyFUrX19520p/h3KiOSiTrEhC2Z4qHVI3J/7OguBoP1z3RhJqr1DrIArbqTcHAK7K
wRpTIOuzm13xgO56PYMWs3ALqSI/RuYvYoeplFsHT52cTnqLDwdTCC12FfmAnaGzDnZSmgPKcWdO
PsNs3Mxuw14h3rxK6P297ivBJQtQ77xhwFgBV+newSFheOc0huLS8aChSd3a76tqhwsQp++dwqpP
1jVv84odZn8v1GA9DzBLNB6dU3icd9ZcRXeZlPhA5LmNPEV6cStj9HdZQ4LgoSZ+9wZegS39+XK8
dNU4LiXQreA6ey9WmqHIykAQVKus9DbnBftv5zERv/chlzl5RTkXtJ7wvQeN2lzy1L2pX/+zGx9Y
olZJfEuuEOcwYBC8k09vFfpuWzpUwAp3Ii+BK59x46V0C2VeRXZrkIRpAJiZ72VV+BLjv//TT5kO
cToIe0Dfnz+wzPnPv9HcTTWnMmJhVDVEvFc6YI5LGdBbUuGxOy4dGvLZB7XMNq27CSOOiVApmw+2
Y6tZhZpvLvtsxGtKTx3NrGuZ5V5rHE5ZRrkxkTpCeCyFYIYZznYE5xTgTHBUuShCZR0svwbCdtcT
VwB1NIN0KaAVjlz1mMTovG1g1krvqX7bWlphCAbub1E+XwlnHrcEdbffYf2vzFG6Dy1gqYpnEmaE
N0HP1kAF0/xhnZGTvFNGXcVbDf4ZRRm4zDpYuP2uqmj9LogWm5/albVWISwnZ7X+KRSkGEPJOtg8
lKLmUhxHwiiJsnqQh75pw4zD0UPqKhAJR0SP9Dn2edpUarDbpHqlVdB6bPoVDgkt0VY0PwBBdsVz
NCmazO2ZUUiJvzrbs5yXrkZASQD51ZfNXO50ronN2mHfxrcDfQf5bQE/fe5SWcVAgdRMS0QMjUNN
IQu8yoSa6P1uqZWESHz3tu4Mz9SqLVn7XU4yrZj9GI42eLKXmQUgtLLq9ZGbpLhHjdhC9P9uWTKf
UHZ9z4BEogBc9SZzS800AfL85RuC0tlhRK+rF+yZKNClWEUcY+C8j2DqvFL2aUAG5EUQvSiyb+dh
zxUM5EGrkyJonLEFgAJktouA7UJOTuBdmCpDz67mNxaCUHkOQCC79EmXv4b/wdGSYHCmxmhw/Al9
Y6a49QftIRj6njg4bVPTIRnu11QjZOpODK1dgPwLsqXo+cjnuk+dU2bqQRoD5tLWO7hpPa+4sBM4
oRPSH/iJi25JOUX1YbjEfoFmHhTMLgVubfAUE19BrxPn1UpvsoApdywpMwH0iGC5pn3QsK+9JCYb
U4BpRZ8OL4qzsb8ay5HyptGkADbxnwBogWp9jUJehYiHiGbUUJd/YaeTNCS2wArJnT57KEbwAwcT
dXSH7ohWtVRAdA5TRTNhfstVbW6RskdLIVSdWLmrBsKP4c3l1KsymLyJLgEZyKsR31M+fOAy5bh3
nxuchOhf4OB3lPobFy8qJBJHHyC0mJUFl4/a57UJJvmQghL+qQsAPCnzHP9ukfP/h1kpmxQgFgLW
H6VNjpMGaIPhj9od/gsUV144hebwlG1CTZzyYqOb3W8SjIv3lfz90FOuPtXLHEJsLRdBWRDThZnh
McWbSsvuJCOkiBwmT1n06qgML8VvUuBqcAeK3559JFmzYLhT1v5p6juXNk2lx15RrBFbvu1ECdaG
K8xJ6S08VUHjOUbeBIT9+LnN3TY56hTKfl4RwWrjONP8LfwNrvfsWzVa6naH0LywfHmJvsnECvyB
va+aTTQtZoWF8N6P+H5a8BYsdmpTavYyqB4cFvMAdNzcw4p2B0f3p5gfS+k8Oo4htgqqKCYkapeM
rzkehcY76dgVYtu/DGiRrnj3Ey40ATe5ZiDqCdZdeHnHGkFA+3nQQEF9KQosH37UGp2PIV04OLVD
IBS+nEhqIF5STPykl6CdbevQ+EdugB8oIxIYn1uTJc5X/U3dvZHbDZZlP/spFObJEGo2zBWllf0h
ul17cWRMeim/aYiEistuh4iTiF0WVp+hZ81MIPzUVKYtxpdy9hj4HFNpeq4V2uf4nZ3hKMbpur1P
5SBEbm50VDNcAcEr/3RRwR6JshOZUdOCJUUSSGD3pv/t2CAZVi2/cAtg7d54bPHffrKTHo805Kdk
EOZG4xns0a7G+e2SDSzbKq6RfMVUzmOGCd13P0t8GunwhzhCC0Tix3qxHO/xaY8p4idNpAabCs2X
7yNRvDMi83ogCdYH0N3CyhibrVh9qV2VoWVD79z7Csi8yzf3ta2I+QZmXMf/lTwc+rUsyeIrkynb
YVVQqeTG9rp1iExr5PWuo7B2goPU5CDlk7+gD41nnYLznTk6EdtNi0lE63mBgVHrNc+mr/nAUDbU
QVNkLRF6NKMWGWscQeN7qKBRokkyFqY9AJi4Zb52I5w901t+cK6Gk9Kqh3QlHMhrgCuvZ6/iECrV
bjD2m9FGwNrW67HFxc6X7x1j3ukmoZufXWLoxt21goLF1ldow/1bR/D5xWqLULY5lfDXdnWHtbVp
5K/cdMLEQSeuo7CuptJCRXtCZIueohBkGwVi7EuJ9NNtUNoMb34FEMEGXMhlXc7Q9IVrOum35xy4
qZeZCtY7oErFr1kQzYQfcmX8kypWclmeQH2hd54ZOcsJiEBRqlVRThkTUS5/wm9vUrpfqZjXzeyX
Jsm7KOOIfr9WmQxXqGpwAIXKwZTCIytN6ovm9rGY/aUgU2kXE6NWF8z/ObxRni57I7xgVVY+LHMR
z5wWguIKwzVjSFY4xT89K4BvEj37n422ICXvOy3BRTYtmfRqF1V1yjLFyOKkQPIQSinZqYTLFJ4v
bvFNi3XSPtqBdHkoq67YKi9p8GRvFfjUz23gQDL8Rn7ZJQ3Zd70FT2YpuyaLspnG8e72jp9Bf4mo
jyuuRApq+puUgfgH7y9VN9i/Xy8AleV4j6bi6/7BMX0+2BWXxWGbyx3EijjjUhMM9Jm9HSf+mKgk
JzPyOXnIaYEIWFQUdkjErjt/fvsDrkGslWQQSIGs1uB1jteB5HoxK+EPt4+mvG9kezsbzDz4HsvJ
X4vCKXBk11GvUpbynbI7XGnMn/VYYKthxp7K2C5bwPE3e4Wurf91qMWz40FFYRYr5hFEp89RpH8S
1EkZasBTDfNR1sFEQg5icBjSx9ojSUL2eecOiV0SyiNKh8aslduxciH0+NOG3weegH7N9o0o/Tj+
mucnVWjUhlLvCY+vX5lh0D+chRtsauBUpqnuPUM7S/XRugNtl0WKjLVq7BezEJZsiNGpwd44hJsE
df4KDOaZpHrv4yyhQvlVC4WgZjonbBrO+PJ0BOoKNgmWixB2kDVlQWDNT+lRh+xqtX8OIqBQsmkn
t9GrIz83uVhCcYIe3VQz4ojh2knFcf0IZ0tOms58ynqVD5koZcAba4a1CSEAeHj/y3dROCViJ71B
YqKIsB3uIFZI1pLxqu4oRgnEYGPWRXKK2N3pA6C2OEuo/izmfCn7t/AgxVvEwH3dQEMADapgKApA
pbHGHtQDcfckyfXsOhofbqFE5xrpCcz5wyTlg5twIOAVMcsBYpskmdqewXVVqHNAGzyHVjRhGg/9
qb7ijdrexGEr4auy32WgBRrTnOw0D+pM1uVxdwMQRDf6Rs4Eou0HR8mKl7LeCoj1vSpYWcIKWEwS
20CgUsj2ijCY/i4BauvCjaqcdjFK/g8MJq2dAx8H6GmKglVeO+lCEviwAU8wBtSKC72E6syeU6Jx
OqvtpUJ8o5tt13PCeoiFD0ldF2CTW8K4VfUb+8HUGjx3BxbYUiKJerdRUKi1CnEiNlEQ9OBwHgi1
bCaqCpm53M9fHNn4luLibW5M9CS3xzZ2ZCVI4oU/rS2qidDucouKPisrBe8VrKz+jKA/Yj1yWZ/g
zBvpMb75OOsLcQcv1O8T/I4wV0TKY9aG1AsymqYOfExGvsE6ZyvML9Z3v3vsA32HZei7sd3VZJf0
YaQw2XUArQESy5iI3z7X8Ee8AhCC3spYMpQ9tJ4mS9n5mJoh248ptz2Y3pSil/5lt+zgmI6xM0mJ
r482xSmjZsHQoPQO2VsgfT7iqkNV0T8BzJ1i51hmrsu0oPMUspzl8wE8kg4scUNcPUCK+AOninS+
iB6U+Uu9DDcLU4bJG5gP/Lp5UgdUuOXaIf48EtycZrqreTyBupb1V+5OcXkvglaLgXfw8xeb9UG+
KuU0yQ0y3uZyUcYX8W8bvlR9b0vR00gaMWus9GyaFwiKt8dHgvLmkZRAzWOBPw31kme3H3WEYoU0
/DJXiE3JFuB2xXDkmAtMQTpz8lyXSL5sPz6B6M2gtjsMdoUepzwQi6BKE1S4G4e1irS3slxuquuJ
PCMnj9FCExm4EkHP4SrWTH12QmkhB9JeCJnTTs/tL7oTl0x7Q4kgn0zo5YQhaTVmyb7RCWwpf8u3
qLpYH8FikpSd28Mi2SiXEFANWAHGyiiu9RqWMfeF4BXho0GLhUt2iaH7dat/rZ7udFJFfwDwJ6Ao
wA2Zwtp/35l7W/HwdBBIRMfnik7Q85EoJzRXaa2pKFze+zrGMUuyHJiLFOmlld1waT2GiLevy2Fr
myBB1fBCljHirZA/zJYYVYNXmAfmwsbOZuRoJUpqw49GmuKwKLNVklF3tcpgFB1ZCXbGOtt4NKAL
YCHxKzmhtC7vtYdjabFUxQwBHiGT4Bp55reelPTRcnZg9XvwPqBc7uSTF+qmEacbeCBF2r6qdgq2
HPbsAQ9aelfNflpQkH7oVbixBQBkusAOqECSKOrylHwQaoAkrS5PeW3QORkZObRyf1jnfWkfpENV
HUjBPiLDpQyBxYrJWCLXV4jeJdcrtrXkoXsIPUfmyjFZL0S0OvCjTkUiOPCgbppbCdPtHIYVo41N
q2qeWbe85p2cZHjp4OeXcrNbUSj3tSmS5znv/egGb3uDeqWcbuxmDsUrf9ED0gz0WBnp4N9A96s/
AKzWAedmoVmlhgztYttXCDLI2PFa0Wgsbl+0twWGLMw+OvhXz9LsbaJ+2q5RB91ww8e5Hkp51nCz
QDsxHT42r+NSxAyAAdBPkJqJSBsHkzmaNjFbyXBdWMPdrZVSskI6YxBTvBRq6nheVazwvzHObmsA
M56tpdOOlXctwpTq3EQyR8K47nfYzpZ/1EqCj3UcibVcLGunfQhQ3WT+yYmJCtNw19TDDRz4Vukn
D6y1HoQdpciH12bcSDIU8hDUV/xyzJoDO6HCG02hORePOWHSpg5XkfZsXvIHYO0BtIDcJP2ykJff
jMpEvcyqkXcFyfwXhpZW+bChOTTRwhL+rPSuDQjYkIuEvTqrmF6YV4XIAqXwbnEgiLuo8rOetbcY
59aGZTbaDuuXEzOG/szFp4sWp3REPhoIJ92kKTHvFnbRk0jCRNEbjHCcdvTcLrtet2kzyo+r1Ypd
aX/CuIYMAHgIVONY7T84kvXPUViQNH4EuPFUiEyzdzYd6sfJVddAEBxj11slQkVd/aImofYF0Oip
PKk9DVJGYyfsFMhKDyC9a7xtsnRP1aI/9SvVSd1Hq6ZHDrpXUPOIzuxVQesovl43yQLhM1ii3evn
Bn7ktJPgUx6VEIVyc8Ktb8ETamFZdxdlIh9Uhh9Ro+lC0X+Lmi0J25QKIXxRW86kr5EMivD2bjnq
4IE6gL0QcMF9tQ6pr3uCjSAwqHVnjHihvawuwrsxgSMOYjeSwNp40HMbyAE2uq2PJUkDfeykl6gN
JzWwKurGCwKyNckzHXtMao7FC9k/3MpMiX8Il9ThaBfHqjcc7/7uUHz5FjOWTj5Od9HKwNuT1Po9
MXDwEfsFAo9xhJFNFYlk43622+r34R8drQfZHw73g2THweEILptnW5JWn2FIQjSpMi3dzWvvSzt/
fgXkIqhwtDFAe7r+b2+jkXg0pQb3YkBhdle3tzTULF/MQwsEYI8PMUvaJ5qP7v4OfYPqKkYeaJvy
tqtmtMTYVMW8cHNNnFl2Iavmtr0cDpGMrZnxKQ6aZesvhbH1txnl4ZeN2mi0A1gmonIih08JD/Yf
UL9fEbEkV1nbLSBYRGYX9jCl7T8gredTqOU5FuaAQ9VAUXp3o3RPt4Gvjmb4MT5jF+kx6w38HhL1
aeeAQDi5rpGCE6cz4gYXSXpOgym54VVH4ReUPSrkTtMAiGChCN6l//7j2H18j0YDIMhAsDOPYR64
/NdPA2ublOolEISnO2kTpB5fGDGvmoGXvmefjirsnCDCnOyPqFoWu2Sq6Mm3SnmGVCNgphjiiLqj
rGWdluICj8A9lDwoFMz2nAXEcvSu2VZEdYGZmbZhY57lNRJJ3B5brLGlAn5maMHHbPkoTgKdEXyo
lxT8yOa6b+yTRbd6lLMz11E6NF2IfBupxwBVSOtCJWXOC6mtWJHXloVqmHZ9vrSz3v/kCPvjj6qp
gFp1q+FvkhGR1qcLAaf1MLX5peTbiLKcSvDgcpRyFEh6MaL4HgBAPm4B+ouXRBx+kJBKhcXIUkV/
a6kfL7Miu2WTeSR/qbhrLNx9qVG6sMNj9U+OkMYBrhobVVxfjp9PzrvNYcxnEyAJYIycTQ3Fc5cX
zc3eART+ZOXYnU07kGJhsK+2koLE0pNaTZ0vl0kfmKCgfl1LEKPvkWCc3xqWdm4hBFjXAEpORk10
i6dg9lRuLIUzg4ywmhX7pcPMV7EgDWramSnCbG+fg/Oe1DjeVpZP7EeVXXGFOjkSzdfzgRPdZiHZ
6tKl409LCbuL6CYD3z5464O/G1xvx8skcw5bzhQmwhAOCxzcLWI0YuI1eXk/OBWaXRjfTokK+HpM
blrhPJ0i5fK4Nk3u2PpmbhJ21cRevDNQbtoTc5DF8uCn2wKhV0dZdJYVqxKTTMUvW9z2rGRGrAeY
WQhToSioY7tH85YP1QOqNkaSx+Rjqa7UBwBatiAR7iU0dmj/SWYbXVF0BE3Ddz388zjIu7rcWUjv
6bazfLD+o5rh234jTh0LAUdUG4RoY6mb2lWHa0jDeoo8mr1DcInJcqagU+qlknE5G8iW2JqwH6ua
igaFzmgIu0lvgHxg4PU7ri5W/Cxddkwp/SlDpkL4YD/N3jLGpuf2JcClvnLIzIv3OS5kqi/7a9vw
2a61clKDQSbarmqr5KEWwZ729aqY4h9TiUXtZAFwZpn7DKXwNRIHuJXGfAi0MtdHfsKFonbUcdV/
Ciok7hrlsGkDd3/xlw0SVNRyAAB4ADcMiHTstxVOtuEHOU92vxUXxZTudSYK/0R6DRh9IzSL0g/i
hal5YoS0Bh9bjjEeyHSMe3mHw+GFQ5wa2tlwDQAcN+ELDomTR9SBDDn8VcbSS8hNjJzPNIyJuuCw
jWfUBmeI3KS6bwRS24kQ6Vlp28noOAYV1WlCMxxyc4snstUh3/PGIpRObmLVnRweHgrIhf0dPIyZ
w55Jhw+wameLh5CWtLuZ+BOI/KJu5QXAT7TL5G2XYg0WSH60IvRNAYTUeIaTCh16z+CdlcQAroGc
KioKaZF0tNdvL/xUBG//u3rdXsboMiJpwo6WTIfZnCae57B47XuNYERVPdhxlo6aITPzpYbWO42i
EInDtWVTEEe+iNnYji5oULqwDzIzBmsvG9TT01q65qG50v7xMShefLQEpn18ibZMdkG/brRG59xG
o5HVwtCD7SwTKc4jPFUHmrYLsgqyKmZNCbcU4H/WB9i8yIMKJjjzOnrk7FsPv792Gm3voxF3oymZ
rLGilnC7/3owLQDw3HqO8U8Uiy0edUSWFqPNuDexXGKYlw1+jK+Q6YG/sM+nyoMPAlKRMbDt9/hd
mJGG6+GWMmbDmN9eBFTE6idqKnHldmatbqVf5OxLVfthJNp3nsqAiYF+ltvSAsyBjxAaaBEQ+cns
f32Qhd22RIxTU/E0IBM0n2GBgrf1BMLzmD1tZX4M+fMSHpbTiNy43zuFds24XQZYiI5BbJzY0JUk
0X8WXpywgnwGtDHeR77JyGFV5KvJDEq4b6wnd3QAkjSVc4XNcBo0aQDmnOTk06fGrX0RpRKhvtOE
QLg5dHZ/H2Ebr+1H+njib+YaOmVQYVkHzcgIavUcVf+HtxVQOO9M8K9a5fMdFYw9sBqrgLNB2IXr
umnLXc2Sr27DEN0dVBHIPzwrnwzu7PwkD/w3zQpiUaoX5+1e4aWdHAUWt1DCZ7hfH33mIaxI+OA5
QK+pjlpsF18Yk64FacvrXkeAXt4Q+dPInY6RWVT2LAfmvaNMKtkNvIhHGkFrjHJZutb5AI9Z2fHG
pzMXqu/4NfLXe/8UeYhG1nMtlf/KcZCe2A5LpesVzs4P4mKugiOAwW63wgJhvNSnKP7797IQI8mf
L9/L4Bgh8s8iO7PQJALAtaTdksfS5p2vjq9O2Wh+JME0oLi5in9fLxBotzclzrlhJJsKLebqy7FE
Hir0e8P6trFBLX8HPMTrXTffd0vYsQPZbZyNT46Ysh67Tt1YXGWjv7B4wARO+hTDntFlmPp7Cerb
uVKBooN1c933PmuKoYDdXyQFETqJD/FTfKnTK/ZYTSWk8bgMBRog1cWm68nKK9jJmM+CtIaYemYD
aPJAxhrBJp/ZjxGIU9UF+2/v7xS+jgKt65edP2MHNi9Y04ju4mJq+ylXWc3FIyhRZjGboteYCK2N
H12QLS8djWjYXkjKyx22kXuhI5annBddTMYjhbtBZ7BL9+J2njLEq2vbJas9qAgUew1YiSQqLqAd
crn4PHUp+WIbi4RoeMmwhZtN+1x1ffvrnq14ZQDVJoxYvs8gn79fwFeFPLbijV3mEgShpcMSMbB7
qDb6ay37UhqIbi0RoauYkG1qdt6LbbCu2DxIcUXCz6qJRxps/+L+TiasyXEDbUNOmn9APW0kGNhs
GEK/1D4mVZw+EOlIhWmUhtUWoIoRrxKvmdQBbrR6vWQ3LA1WvkqysnH6niHwppQ/h0h4RHE/YNBL
QRk6qkO9wM+z+9eF5ImU3MaXX0kJfsAPMBgq+NHFBv+Pc+1qUF4ctGKGVtnhxxfwfOL2y+GF7lX3
D5quPaq4AGDxNpdYKQRVI1wscjdQwPMqWZE9DCne9dzThK+Kgfu/wlIvrX/v1FND/jmeatKdHvIU
F0YF7C3ynFTQwBzLT5WOhsHyhPQXggjsJGThYO9T6usWi5LvK6jeABAWMX2j1idzFNGkdnBsbVrW
UPWzN+oxUYfb17jeiRfrr6wqosS/itCTnElljWDj1/AzQgbBEXN0Ddl1j2/a3cToYZEeoQrm18bw
S22hT5G/bdtmp98LRf38yppz7Ro5rYmO9wkH/q62drLA8YXnUGmMmYpD+XateYvQCA4oDv/mXMc/
PM+INIbo8bCRMpDf9ZUp1I4XeUSuyhHklSkD602L/7BJxa07lzic4Zc+MzO+d8H7fjroZQoVDxqN
L2S+kBFUSAlFb77twWDLuLC5Dc3KdMmh9nYMyD3sXGzP2HjTr54F/3wX1LiVxLL4jU+i9ACQEDlx
zCHsV36oqGd2RcqZxTZ8KK5XTHj3FrnBjta0woxiDfFjle/MhSXNQJy+HUYCM1yjj7oIv2/aCxNV
w/MYQZboxgBUbPu6PW4PLbrnXzKar4JASIbjPgoidykFSvsGbsN305tH8cFUf82rCsd1RhpbGV4V
lDjYInqfxyUM9eZLqfJx3/opYVHWm7DEZEtX5meVf5CuXAxEgFyNgAutzMm7Pc67607TSQJ6745M
Q2Vm6K2pMq2Ov+9kPmWJGwaIFJccdnqXYjIGzJUcei0wFFqIRAUVYWlMS9TTbO5pAcwA/+MrIN4r
nnYsvK6drW0T7dGOXd3svSQrB3yDh8w0Fpvq2WOmu+0TEF0BV8HqwOOkeVCNvhN4kaQsM/q/JLcE
3uCoBQDNTzy8V46vikatjoLS9sgJF6C8zLVTB/4B2uPLninnEaGuhlB/usgQoEvKZdGu0npTNeJE
j/kajvGPWUjIGc5nICeJX9p2ZAxMF851EeCF5FHLroq8Ktp9vP0K8PJmFzWB/DtXai75D97tLy25
4lr4kVMzNVOn41q+3BMlbtADHsfjccsTqMIZ2353ozSPpbYp8P0kRQDd2q96VTdEr3dOkIg6jkd3
At2L6txt9PVwD2Sau4K9sE33CMkf3irQAvAVGUYOnaIk2A2TVjd0unXnDh4J7+oHmH1jD6hQ91yI
R2s+tv+JjyUjp58vyRzW8Xx4vgIXEMArJzdZ6/jYzViPemRdbJWnp+6muBh4A7YUtY7tfvlbhSIK
x9RbvcNgXr48l2Mk9P4vEuQZFvL1QNtzQH5+oPk2ZY+MtI/51edGsWDTz+9hlvS2R3lXbyypxTAk
kCbcw0Ievf6Mh3NIOXRnvI3hfGKZ7ocJuoxSmF79b57ENbsfyiJDyuaXQqAzXjjb2fF3ouTOljq7
SWep8xhj2flSqBsE3Pp3ifQbk1y+94Y7i3YCrUa8wvuokbqOrLg7kKZFBKXYz86HWkM2Onk/kdSY
rf1ESiaC/zMBN6o4bngy/SZTpYLS8a2K9Di797PcognmzOnxO4r9IBGN3x1q5wB3TJRyd9lqSsc9
tqBkn8I29g9Vq33aRTpb7UTXze8LdxEI7DvEAiQuIVBIW+a3O/nBByR234QxCo7DuSTM0yBfd6Kv
cfatnAOyQANJRy1gxvFPYGb/LutuW09ts4omohf048UgkQ3j0bPN9whos8yw4pFhy0gtfYjVkK9U
pV2XP6ZlKy5BcikHMiFpn/k5sVJ2e4sFzMKCk+mLZDySOJFqOgmHNpmcH/MMxI6zKRDBHLBB/pr/
Cxw4us3P3lEBJFz8XuG4Xqgla99V5Hpp0UC1gGOHCe6gj2De0bkm/x+9d+j4hM3pUXU8nJkdGcC2
g5wx9LMlqC16pSeGoinSDEFjHfLIFqh+U7YXPuIYBP6BhwULgCWjfuU0OuckXWDLUJgbR5Me4qRB
+U3on6vC3F454mP8yb2diGemltXRIYGmlZZOfSYOCIBO1Bob4zJ3BEtFtIvEXwHBJLr2fGv3Ip+8
HHCv+tYxGgdEJrvtBBYMalDvN+TQzQ0gt6ZYIkDXc6S7tVBHx8s2tt1D7ViU/xDUm86t7SZByAaU
zp1f4USe6u3SAwb9g93YOd+I71Rivemh9MzEcy6XxpVl/pixBDdYiVTjxB5PNX9SbYfMQsoK8cMQ
tdhI0PSUskciYwLye37jOK4aUD6RFSsnF5Bj6+K5YN0my8yGIZv/rLTl8uJ6gOhcS7p03w45HzX/
R/d+P798jM06cIyCj+bAxwkrMDWJlRI7M8JFeJjoRAiiPH/2JkiYIqn/VdirZRZLln8LfDMOPaPm
tN5E1T8DPmFp0jTE34nP+8kkO9cmgxfWwGYr/1yvb/2OX/CAOSKalWlADRsBzB7Sfdiicysb42fy
zhMK/iYT5/24qMWGDCRXL1jzU3YrlyVTjtKLRz4xjN0YVIPMtDSxtrops0saKasL8Q2Gou768lRc
iPlIT8Xh5bPb8XNEcVM25EpF8lXq4brzIcsl+L+htxHJKXglF2xMtReSYWX8jeDTv3IXWLo0B+x3
xBCUyFssGaakSec4JaG2zXSfSRjxjT820+dAjp3csNLHMKnWZpkaQx6ufr1P+fNntZvArvFmNVFZ
zWsHUGYDSrL41aPsPPB/zI5OKm/k07OLU3p39Xaf+G8/ZY7TrfxlqTKDVXrKKeJHKeleLZ0ijEDe
sYNR6Y8Kk0FKg3WojQ9Hr4URBzxuAkYztV/ayRqcPQ9DJ79RuqVfhVLDNuLJ6k3C2UaFga9RZtgQ
sJmd3p4MQYl1fDeAqhkv8Y2WAz8oMZDaq1+DznlCW8gbCdxPOPCxC0UppCN7neAtSpMAybuuCkzk
cdT40GT8g7wQhofWHCSJlmTfaLiF1/ohGYK5AnFZJeNK+7ZGnpwCObZ2vt/gGi14FBB7bxm0NgA1
YD6E2faXNGVlX5njoPZasmn+DLUKyxfYtqWNaGTxLhDIuBjokTgmd42aze+YBRMcPZKIWiXH7Wzt
mGdBN5tYmevmYW1nJHkTHOhgKIHYQkfrcvysmhuS1z8zA4l6fiuzmkPi/0/brXTtB3nzVCLQlyVh
G3WCHEn1Bo1HmMH9F93ffuXbbizarXim1AjFYMJEecio5oyGRdPpTUEFu3E2VKwzwrw3+hIupv3x
uF6dAtGZaAf4lJzScSNuZjO4dwS4h8V0EeAc4m29uqN3s3mPg310o6nJnYpnD3fsR6o/cdEk5lw3
UlzbLmd4moj5udoK+QLPligLDlGtjXfDegbIyM3kRyGDCPvkicfplLrJsYVMqIzTWHkkam1oHrkS
U0WS54pipXYkLBvsPiSk0geLUFxAf3GKHWrUOFj0z6hL/xQCvDZsLejfrrqXKJZ1u+ekeFR8Fj1M
uYluitA0eYrQcQiGmElsGvt41BrwwBVmwOY+2vXRjjuqaYy//E8sFzX9+dCFWJIgfTKHh+ht68gR
9UCIwx9d2BhiAXw3eTws+Sv4meuS2QtvxDDOyCDq3xe/bQzB8u72V8rAO3fNXdWddK+ginuQhMRE
57ki2sjsWdHc71k0VeS8y3j4yEjb64OfJF3Rr1093AcSmtzwmbApIumleZzcouTc4w9QsDAnrb9E
sYrhbGqmG4O6Rz3vcp5H1OzxjRaSiuP4NjGyLTfsSyD7N6D9EAhJzIhFQ60QsqoDP26IT1TGZN56
tgoZ6IYOu96yBa9H07M442h3WEI09sy39h2Wd/vdnruaRFx9Kzj46PpsrtUoRgMX0eHUjxocJ84i
34B9oXGF5aK2RrQaOmVhH7Fh17pdhaJ7Ri5RSMCZbdOUwO+ymo0JsMwo7d8nsC9NK6qWU1YNJR0a
bNdRwN5QERPcgzAt+a/EOy1hzwQAscCErjnupOgCrzi4w3g8v0Wlb5wb9P4FnS8GQgedVcn+1rQp
+tfkvC06hfQF4fIJh6ZZEo+i5V4nj/Ut07TqNct6HirjUsTJtleYTQ4psllmPQNk+8Z26yNyISuj
eYLe8juvBGDHXXFhG3m2pk8S0BedffzwfsJ5k2auDI59GmhcSPQmFy/iEBh66R93GgTymglhx37w
LrGWPAyEw4BAHOijer2BR/Sdh8w+4uq2zCWwcvDLpWuMA46fAEWRJnLmePhVL7QZgkor+XChkkaW
U8DVzcsp5V5MWN1M4Z9C2BWN/DcypVLiaXo65zh2cHmPAGfABu5Erszf6XrTo8LzBgBDHrjxLSQz
FDzfa6erRtOPde96aZqY2avXABThs2xKZoF0UVHk9fcqS1+mvSMhyW2HT4VRxgrkbHPi2bwZjokX
tDFJWEJZnxT2HNY1vU7PTfNC6xMRFtbKM4dVxzWSJEu2829lF7YcZ7W+E/VBzv2jYYK+FwqENJ+p
O1WMgrYDRBPssqyUpmmIc6gq0KLiWpS0d9HXQ/RqkPZL2SMd0RITod1X5zDAGiJXKzIHmlzHIyCq
DlLOLpgmMleXw9yKNmAtnp1Lr/yS8qjG3aTpxkpjWGyaaVsYDL43xJZUKZGdMjToNeEAdqJdfgRN
IY3n+WR7ERoUaQNVZQKQpdtoWOv5jze47lIPN9eD6JRWslX46IKsZKda5HnCNrUHYTQH6bISrltk
mt6GbSua9qsxt3GvQtJlOi+wXDiTRL1sQj/MWsmHXcpEXBd5QvkWI9fdt4VZ/i4NKWBGH7Ge4nQK
8WVrsgSD2EJ1Knne38af8tNSMViLlzp6SXPPxGyp5ZJcHGo1i5TM0ZtnCxtOTVeIBdWs7aUB8ZVb
z4SMgF7hbsspdbENha9I6Nb+W8gNS+ZnHqe6zz9/3MRSezX0iMgga3C97Cn904L+Xbgad0GaGTdc
a1NZQsKxRxgBuJONw3eun/ZWHQUsfja/ESdTsg/+nHvg71T8wdQ7YcviIKkB66k8tm9ipOLCWs5C
V0roKkMJyBwrS6PbZVYEJQzViNeN4LuUrCf14HE8Q3/o177USMLvYcxA1zvjYM+Y0XQBsXge1Lg6
zngLTcYHQt19SgzUQGJMC4TbRihlPNv/9IOiJ91ljpkQ9cVAHAGT5wFkLe2/6sWn1/QyhjRWHirl
dgsrsnpG168I2IHfmQJJ1FWXozNkibLS0X8sENrSCUZpsfAnj0/5yqZlHxb5XnxZWtvspQXPl3AR
yzD2t5ZJMBA+csH7lvw436El6MRGHDIlrv2JEJRzajpJKwmOL3uT55eOnxWSMGzHxIvJEIueJrgN
HfRxK7QaieH3LwSwFfH9xQDwT3Uu7l8F/e4we+6T7/i5RxvXu4GON65qJ/i1jO6xL9/rS8lOiS03
3GQH2Bhh5nA924VoAKU8qOUChMf+nJybi6qJbVuSmun7CESRJbrutv97pAlQWpRTC9hRkrZ1MW+Z
HuvA/xMbnFZSbB3Yv/sgthmVRVvsFhsq8eyIaUKTHKOP/IWO4j4/xpQp+on4pktJ0DS4hz/Zc6uc
qq9treMhTD48FzF5VxB4ciDXU6yRd9A94g8aU7vJu2uKmQof+oJrZTmvgDX+MWiOptxP4lixIO2A
KgQLzQA5nFFG4QVylsa6AvYRLLAdiUIFFS6Zqb7StxkVFsCiMK6QYEN/BX8grs5o4bdqPvpNpbys
v+vK5RU7khBq5nwSa0CS+VQQ0H1zGrQperKEQLxOzKqp5TLYodHlddn1I+3zrJWK4VywW6kjfO+9
Z6H32KZuGfkb0fHTkV56FV2Z0HJzYgJmChlrwkV34i7bPUdqjTQCsqoRrv9yl0QvZ46vnGu8s39o
ktoC1neSP67w2pcD0aRZVigmOLG53BurKcAjxsg44eaHvoR9LMxEk/6RRoiiE9hPTzMt6zKQQ8mK
UDSLY8RrdDF4dt6p3e+PYanSkWHZ7y3Ql/UlZMCqmx96FCEA98rqvEBvHj14z9nGhMBHm7urBBWA
/dhBo/ef2jHFD2pEY0sh6tFptaTlHUA35WsX3ZDeURKLUVYNvQt3RZNcCbA85kpkhrhf0OK1Xos6
lSqEFq64bKn19fqkly/qrp0O+w4sSi4wTkMb9uQgU/cy2rMQNZdo9XlnbBBaSszmxNpyXnHWjq0J
vclTHk/Cv7z0X+of68UPDRXPZE7BBFVBoubiRCjjvLO2hVavuZOhiLMvZNuWBML4pIGoWzyw8tui
XdstapzcE8g0d6Czl6DNhhXBORWLK4aeOoGHnWTjHpP6ERzIRLg+dn3ELTshI8VoEhHtd+F1YYL/
97o9sppFazYP8D/tIkRz+AQ2s1l+Igh2bJAVRuwCS610AH4vn/6dzBz0aiFMzAYZQgwRsd8RqafW
3LyjANWoOsjRThkW7CAHMi1psbCrwHpIgpZeNAk+0xG3TAK2eqYYB1sjegFWfsbS3lwB74luMBkx
k23qOm8NM6EwRNtItkFQfWmDadvqaFNGN3xQhmYFarkYwvC9KNN+qokb9znPsp25bz+OU/jEsojU
V2VK/o0+QIywLFG8smBJDMrDYD9liOc4VCfSA45HQs9N/8tluM5Jpm3PCNqjk/xsZrFNMiVhusK8
Z40rzhbvOS4s/E5UeQLJtM+7OBmWCWMfLRwTexKxiW36NqrQ1mN9hMQRSS9nIWTumjiaKLxyAbvR
mKj21I0kvN+nWWuoKpFPwYdNWJqdFmKlnmQyUa+/JSdykAIYC+oPC9ItiWZ95bV4081EY43gJe4q
1kAGMCe/sg+9VM9g5LCt8msK9EVkFDqleQHPqSPQ3lbGI3WFD1fxUTG4hZdyXoGQ837ilWHWJwRx
kTFRbplOCG4U2Qs4++g2hciVFXVpfEZ08J7+wmjblWMLS6BrgtmkxnGLeUSvYy7/C42z3W7t0kFp
8gCzYFSAzChrMg/iCN/ZUUoPuSCHhZJEdgmLGd5c+qWoLJfcN3BhrWLqubA6ud4ZY1XX22P4IN0+
kwtfxlH0qgIAz9qrOiGB7ldBuKfFQRd6XFDC31eE5Sw7L18jOa4LwmrkkFJQ1I6g1FkQv4aPftXf
HPqd4HQvI84yQyquu1Icnf9CqCTZrg77wbRGdPHgw1krHIn805YKH/Pl3kK4zDpz5tRYBD75Zjnw
P9cpHb+2OgBNcGGGNjgEZix22IIy12OIjCng65UpqNMs69cmLLwMMSpvk8qwV5vvVv1iXFqczB7N
IAa3asUdIfFBGd3Pz8rxv/VcJqcJ0RMQyg9CsPkBRh+bHaDDQz7kWgwx27lbIaeAxZweYr/Iy49j
3detfaJeC4zR6lbDYw8aJWGqDfPM8Cn6iV+CNi+Wz2isk1uRKKuMWzXD2wBHjq8LzEIqNiofLyxm
yrKYZ3pkIBTyWmkvPew+1Y4ZQwKTnQcyBSvxRJTuM9Zmc5YLKuwAAT2pnw4BId/Di6EbY1FA/Ghz
J4gWGuxmxuarFP53rNcuUBTbn9DGEz0vHqPFOZllpV7W2WYoobZ9SUa0/8Z2E681WICvM1HDi4xe
7cx1cv2V8ohO4JOqpV1qBSZqh5ig1NszAsjD4tLup3fofSxPqTcW0i1j/1/Z3ipoP1Gh/DMnuxSb
L0tG7p2c/yvrNQisRVCSvrO1Hx0onPGWBagOlqabdgxg0BvIuYEfbp0XmVWEoX+cLlKJrD9nuryi
Y6u77nUCJU3X6nA1I26UcDA8Kx3NhWiCIGNIaQj29lr6HLJtR+j6jMgtCGD01Uw2M6UldnDVC757
Ios+xxP+ymbHZtUtIUVpGlfhCaJelI0zJu/id/HEmF+7RXe53LrdNHt8zpnSSENWAW4VpaZ9Rigb
8sP+KNUTOvRQXvU+1z5QHaLQyBZQ1ljN+6GtolkM3QfW3XfrPDdq/Sym5OKT16PHlIXKLo1vj6+m
4UdrZwGsRTuF7jxYhqU9COTP0Z2gdzequjaN7OqEBs939u8ZNgQuV1t8diRPznNSiAACCnMiNj39
61MYAMxYQs8cYB8ULNoSF+y62GKMtfQLNVOFx9JOMAB/ylVP9k1zDzbaxjHlBsxC+I7HQKhnQC3K
9XRf/oQl2Y4A75KNp0t55D63slV+3YRzAB4/cESv6kGePvLPaQR6MdoSE3sPJi/D7IbaHwcMNot7
IoDjHWEk/QiJm8OMDhlOwdZpt9E82nhTtoqmxzjrn3m/fU7fYkdZ8VCsJmI0NIIvEiqdc8cdWkQe
80SBY7/LelsA0bngWX1qvY+WTyQ447R9hScWa5018PixcrHS6GZP8YUvF6mqNKHLH+om83Ixitgn
nvg4ZKq5HsNiQpRMXgvPKiU1HnuM08WMPntCbE5Gl7PzIJo0SWqiJUVCKSzNgfSiIheAfqfvv4MQ
JJRLqoo5qQFk/ITchTKe8zPp+F4DIUWVeRX75xByqvmpZHF1UAm0GsKfW6yqb9AFfadJapeuZc6x
iVV5bmOo3FkhiuDJRwbcPBRFl2XJYZQ6Imcw9FLwnWyKPu0haObPIQxee4lttgszoqBb4KRO9oav
giEeiMexTZeiGNrqrzDz8QhdYrXP5OfK1azKELkIHEyEmy8buCXFudgDztKMlyup/EjKt0+yb4Xq
/HtRxHoRsIVu8vziEsuJyTekfSQMdbq9/PwyeyYaC0mZwXIFGNBJGUVPs8LgAgdaa5KodSpindeh
csDWNHN/s20JAeTSP5bRsftbEyNNZkiSPma2cpZuLt/TNpaGzlC1LCitkROx2tuzKWO8LBklSk0m
QuEmVh9Aef0rbm+LRxmD0Zu0crTAa/Kwa48SfXIBZiRmQP06OUL8JU3skDLxAk6p//7n4ikDj+Xl
8u6G4sn3ZQcACSMUApAjZeKhqFuvpY+hzIzleS4DFqgCnmJlH4UnwnnfEPlMu0WbpGaaUn84KEPZ
40+CJwI5Nh/NxLSodP9s7zXU5mvCKa5FOtLoHLKhjFZKm2REv+DdGUtrV9Rb+YQpJPq3aHshDEI0
iyP+hshmwLhu5iCxdx4H+8C+wVWImZGTrxv/3mWD3jP0Isxfrz/HPXHO/6V+RXsDYMFribdAusZY
PONKCZ1U6IU7AfuE/N6avYIrqByInW9y8ST8st58y87nV5F8SwDB6CdrO67DHQHz53lf77zU+oWP
yVD1e0AzvAQPV7f8PmY0Sz5+N17BGu2a9gemfbmCfjEZobSvWd/g9CYHs7Meqn0Jz5tv0vTd6fqI
Z1uGaNj9crkklWiqbLO3lT1hJ76JSZufYNb34rQwFqXrdiabWIPAI8bMYPgXF+2vqODc2JFusiF4
PWtKMPEazJD7CdiLyiXKhztR7d9p/Q/jsn9uht7MKGcUJH0OGp/SpXOyVq6tL7FJbCBHxBEsuf2H
91bqT15MQpF1bFvtz3vOlF9K1YYJRadRSh/H0v8l7K21wqdUIoDcT4an2G48fCVP7coLNieTa2Fr
9xbvuI1y17oKYg7iq8Ny2Q1S8xsrbJKfbwY/3lDbrKuYgs4E3YsuatQ6iohIbUNjQDEsyjLCSc8b
t8cToQaIM59mHuy0bKP9opIIyoESZUq3RhOXh2nqHOopIYSvUcz+dwvtIb1VBRPMIB97Znslz0mH
08VHyJMk1CNdzeGbnbkVAelPnx/6tXhiN4pMiHgaomEHkI/ds+vGFJuHBZimdgSFwedxoe78uPOR
2OsMG6tgUJPJR2LLIv7ibThD+oIRYF+gLxg+e799cW2ppVqyExh8NOKxQ5wrur1tZ6yFGu2eJEIX
ER4Jq5wzmNEWakdRAbGtTxxvk2M3Bk/pL8+kPw4Y1K/SQe/VitMTnUFRXhqI8+Ed8/cSD8SIb3gG
k6P0WjDqtrQvjUqwgCCUROp/Zp7kk+mE/E0aDHaHU8nIw/NGZAE4nre4z0wn2VqRoLrsbbNuNEXt
W2BNX0NnDUndB6xmADyL9dGYrD7zI7X+bduKju9x1egpBbNXbsyhk9OnJiCWgZHQLRjTRkisRUHA
XoJBJLe8wO9D8DAz9WBSt1nlk/PIFJ20nygKLIBBIdwYe566cqvNGO2cfz9ExrYp08RK2K5lTLIp
98wnZV1k/ef48MlYMqij/UV+PYyq9m58kVngJAPhgNkbWKGHqCuIJeyu8IPJT/2a25O7rsYWcPSM
krhL5iuHoTd51ByUVM0bZAXePuUhL9GYuQj38OJhkZfqw9OFngyivAuCCZpMsHJ5JoFos79MZMwy
M8qz6+ykO6o2VAEp7hZB6mRAFyu7x8Y44RRJu8Bia0w5S/ZVt6+1wLTqucotzagvj89T3P3UsdXO
SYfzkRmvU31Zx3I/YwXYec/j6KP0CnKoysjaA1YmVhsdTryeL8OA8m5QNdzsbCAxXQ+XMdSgZPdJ
vplxX2DFrwGMtDwtamiA04rCPAmqd/92/aW15UmCj8LoJ3qz4QLfGuKAvkpYdBZmjL0rKoTxluCh
FZsnx918jyS8o8JzkIV6QfTRcx+x2uTd0J50HVHu5DODJSw5NALQDKPg6oj+luBM0TVTLYyu3HKy
Adwh5W5BySzuOc6HBd7vbKxGFp66+xaUTr4nPLaPf3zOUxr5rDKaZZLR136BevClEuqAswtAtgef
+NPcnJegkVVkhUyH56OuXo6/CCAGqxMCpR3ktfj0y6CV8x2+aAuaTJImW+0LyfLUVujvihCdPG3T
5ZSA8aabPRc+idPskNc71GwsVmjMqSzUN3jzqzh2xafATt6a6NbXxN+0R7y3fRcP6lRN85LbILiN
dXQ0ISjn4o9vVd7o8ib07U4IavcRLEpGkmcYBpwE4Hxxv9f24Pg9+GGpZKd8Hf/d+/Iztd97mJLj
U73xDPfkyh390Xv1P0zMnVffkPcyN9+VrNtgeYo2Ot4ahO7G+y7Go44b76xSvbrMr3jDFCXnKZEh
s7vqvvTp2eymYXrlGpykGCc3mf/f0hyCwQxWtNCv1rSp6qy8EupB4F7+P8iVfiSmawEFz1PQOGJJ
IUhHvsABED7VyYMGXdbtbt17ftOD3Wr7p31gq3wUsHmyL5PLUGjWG2Q90hzsAzUn0R9K3XdR5lT1
nwML0GplXH8Wn82iycTCgrlB3IC2MbATt402FrLDWa+YgkaShI3J9/6pESXj7w/TbyFjCPFQ+9aT
djQ3lVvKWB1YS6airP4hm3JwFHqJbRREX/VPqubEiZJGKgTcQBg3P+/tw5hN6UKn7bS9v74MSx6A
0PtJsKfeIEeZZw7qjuCeIE6ha45M7KtGIFDwjVaZLcvBC3wQ5sBIcA9a7fGBo1brRrh9Y2FYpFUg
lUcQ5IZOmmWyZ2zGiR/7pF+Vhn0sZXCXKz7iBycSoOI3aa4vMjChusud7Ca7iUbZVnF4rSow37E9
+MS4yG/NcERbeXdgWbPzZZ104nvyBDY0iCMowlyvBGd1DKSav70nzd4kOglht43xiOG/CTUUFCGm
pS1ql7kOC7Py8tEMUAR4l82FkAS3pL5hVmsrIKbVACcyUKZcacimtXSWAcGs/5FfzjaQLdGczsZI
cs5ImEhpsDarnPmQBJfpd50uMapM6LtvTFcv2sW6NTyk7wpAy6DIM4vCP2vN8MCBidVc40cPg3By
Mj3I7Hz5LDEtloOQ/sMjnCtcl6LbSo6+Xzyqhm4TMXBSe9qFXtCPbk4vsndGGm4l6uLzlh3F72ri
f/+hbvI5hU9X4mH3320VzGdA07D1JvQH5X/BvwE0DD0FaCixEKiHyTuagHwi0LRjmXJjej0dlDV8
RiLufSzJ5JSGUMqSxCZHMUhIPx2zYMtGV5Iz0Sg3Jmb1WQ/8s6LzhSIJyd5F3fMkaXWAEjxq2MJt
YGPbe9al+pQtRe4wDwbKoW4j9JZXVddcS+5veHl2P8kXIpnrT+p237+4+rcrHog9xiHQtDyC/feM
5joOenwEnzm7TRp7W/hwkza9GkVaOU1i6ZO4qSbB02qfHsYBBsvr++aZyT/kKSiagOxhMi6CBKQU
b3W3yTg9pW+BkCPk8Wp47+TuK9Q6cg1AX6VPfdKg/vEC7o7g6iCqMq1jZbwsqROC7OHVQjQaniSg
gGOu+lKviMTBZvqURSef2ahN6GPOmz855KtVSiwbI1HtuJtjNA3tgRNJdLKr6vhpff7c6nY+A04K
7PwA1Nf4HxTLVU51Izsl+50KlGESZw+EATZaLxmIhpXsiKpOg3mILmnOirVHjIVd0xrZ1BLaYqq7
ynAKF2W7O4Z1YRFA04zCmh+MmhXOoEtoqWEdGK0ULcbM+S/78tMKdvgvEpyA3AiAWzy6+mPD24f0
zt7MvFMD108cX04aCbdYyQ7+XoeE/avBr7fBN7OnR/SSchOnqN9Aej87wwCA0LK8pygzgaojo+EN
8CmlQCYST4sGIhD9ngIRseOoi8IUsFzsLOVMaiFQM21mefaW4KnWmjWbCGvtke7YvhQOUB/076wl
7dfIy4+tNtLSo/3NBMwLWkgfUxpz7kgMeP3O1v0NKdbnXNdy5qCLZfW0TY4FOoMCKtA4nTrKEHFL
9qX3D99/i0a1M5jjAc717qa3E/TU8gPZm+AkWSRqPf9TNTliYXDwC7N7Azg5mrEhZHNQ6Oqi7svh
a1V5UuBzlwjB1xb0eUluEan9flKbdQvXxa23tB1lWoUqqt1d52pb/JIKVGuD0S/TdQinE7O1+HNc
BWLsmBn0mbbI+FjQ6Dk4mkBQ+FlnFpxSj3D1KATbpCIwvvYiTH8CiH3han/io4Tfztn8viLyK/wy
1EO+FP3OnF4XCIdMcD81MvReGAYTsRdXN+/vtvf+PvUKHNoe+Pbe0/hvCz1inAqEmDrZ+31iA7YN
Xy54Sl8vTkvTkfXdGHTdnQQikl0LPlMDW4O8CHEdCFAiGOy8DpEd7gILqp8Xw42h1FFGdI0mIykn
jsQZ9Lf5OSqVE+J9+WunAeJLOdEc1kweYFoj1tRf8g4aWMmIxBNmUD+M3w37RgHoSVKPeqmh5g/a
EHF7B3QZuE9iWXKJz1u0OctYHN8Sraii0azNUIAEqmq3ECgo1xYFtaMGjY5C8Q2aObNDE1SX6gni
9r5Erf1NRZGNyHM3S8YzQ+PGEcZ7KP7HMBVOpOvfFQZyqe0A5zH1MNU66uX5Ekeu+7l94eEkWWtj
vN7+LcCXGnPbp/PLw5CB5+k6eThdVvd+Ovhjbsd28i0QnUnXMyNYFqzdvCgA1I+WqFVddlUvJbY5
DLkL5eZlnLn1jhmwEU1Aa7THVQeVbwlIbTpxR0DkntRqCi+STwMYlQp+hq0zRszvw6FP9f+DxY2V
0YMFjl72fNbG7wkJX3xUJi07dYtr3FGG5wKkRuEagUwMCm9YA6OQYKTMTRoEFh8OKgWdBFT9W/M/
E1mXT+rEEZ9VR1wMnDv66pOCiG5qxSP2RI4Izg+savZII8sfFSVXVsrS1+onBFixGEvC2VJm4fZY
HgzfrkvZ4RfibvgnjSkRGYn2YMUvwsdOqSpyucfKGI2F2aaO6hq8F7rGeBfHyCVoRcpHHGAo3Ov1
2BAPDH1ZARKjplzXKGjnwGUdTjsraqsX+r7HedXthvA6LNMxBPqnDBvgz8xMnq9PDY1UL+03tieW
ybdIB8CzZC5W2WAHTyQ2Lqv0W04VxWUG/HhBHL2VDc4zM5kwb4p+Mh8YR55GPwKt2Kl9cH4Paz3X
NaXv6Nj3egcXycDyxhUCtZ5XKljrf3k/jPFvjTPYDPpKJWF7qDdp4HxJK+paKRw0GEVxD7zFQbTq
QF3puVKrGC9NugpFM3wp8Iv7D2KIWHFUGpwjpPiHr/IxpHQw5uTkF1DZcvK89Ce5MngtHujaGDqA
nM/36YHIVfpyFwhox2sm9ZnpUZq4qHQ+SCdCcObp9BHLVVRmMi3cG3dT8z6ot88QTpojGGa++N/h
PdOLPRUYZjHQM4brqZy+nExFT2KZMQPp+/2XvwPt0jAiunLv5LOfCJpQqFameAEG9j6GoXbKlFcB
NwUxTt6r/sH61PLFHj9JkSDIxCMFv1UTCxYq1NIlAk9dyrTjiN6b0AhapFx/qJmaH8sbLHFz/PKa
QzkwhcSbOGkrV9VQQVPvyesQzHKoo1O2asn5IGS11UL2Htd5GtX+mOHLjUAF/iXbOSbfmkCOmHK9
APctF8SMGwyQnNdR2631pIZeRvN+1b5WcKjHliw5SytuHaJvfbaI+07AFVVWYbWQlNd93ZQPu8gZ
Kota7dgitgwcS04ehW0jRMthfRybozbcGTGMhtLbyzsWxeh5/VyxrQET4gnEDI3Buw8HIYWPH3Tr
qizAFuP12Z6uZ8btDDe8Lgb4VYR5qn5AvW+kuTld31EsVRxacHFw04fCaeyocRERx3LwkyiQvTiP
wi6mCM2w4BxBHlD3H6CZCmk1Q7p+9FhXErmY+gLP6ILmt71lQQD1KfcwT9MJe/mExcuA5hT9fWQ7
UOxLI2McldDav8OkXZ+wyXoqAsqVFAjOEiH/wM12CjEGZzU0zfDUwHItOdtQQD1FNM1yoI0YGCCw
goFoaGCnNiDJFDK6NCDAPKPb926ZZeP6xlGkL0PgVsK4Q4GxTWaZ3yGRIsZi/yzW1r8eBg2/PzER
QALG+Pw2O6Aw4dAwZQj1Bkipi4cDTKf3poyejAuAD7miGMopy9jBM2ML6Ztq0oy9vdoKQS8lE2+5
t3IVVjaXgqOyXcijK3e2th8KvMwh1gCBe6i+C4PTzSXkyp+evO1LDovflnPX+fmLNU0/eqDrYHFs
VCEd4U/A7X8C3rvXLUHRxuU2HNzIGgOHwVMo4M+XWrMZO55IIxTHPrUaGxXaj0sL7xIhELZgYM+g
HJIEkj/IHK1V/hnfS1UGwP2prBA9i2ReUkg9zBZrEGNVgFmSK2XUjbLNi9b6rLXrSe1IEzDi5P39
kqppEegxOzunGPuE618UAE0oS3jV92AB5+U65gNWY6vQO9NdDKVWRpnXeVXst5nElY45As5e1dho
Br/TIEziuIgBfNnSSSyRi6AGYwVFkTO0ijLk3ut4OJE6OXms1eE45q5wZXOGomJT5kpn0GClcn9v
BW+rkjVif/pQ4mqmcwzFLF0+teqCrWgeA0G+laaFJhSqBiI2EhaxpTbTgjbz5FNGj7iih+PKebL4
2o1S1MBryeATrnpFFGEih6znz3Cv51mlWEfwwBUIGwUE0GB6dvGGPHuio8Ws8QgOl2ySLoVWDMb4
dqDrnJLCH60o75O5jpk6nBuaLqzTHfwYHTKsAvu1JsG4vcLYpdgghV4Nxrhz2tFE59hQiE1C7YZy
PjGPcoDpn+KKhIpTa0YvKqTTBTnt9pJCvxTea9sF4c4o5LRw5qEJVSpARUcVDUCWp47z/+U/x5Vo
VMmOYUC5EXZvPpvzZeDzxJqCJcUNK3mjIxPfqGtK+2cD2u2chl1EQnJ0j5EQTzRjdEsNkVncIqGg
MXk+SD9dI+vUnxblpm5OjvRxk2tJUMQcnQGvCjiM49TygHcjJt1HClZKHx3A5AQZsKjZ4dWulNMy
4fqhiP6uAJQhPlGsRpRaG0WeHAJLs4ALC/UgL3zciq7A+WcmBr+ctTLZr+WxRQ7G+e+nHMgEdnwn
5btljoUeaVFQC22mD1WSlaQjZ+jXzBKrFQwq41+X07sMLMGAQs6RAiloyYjnnkpUHBFN1UsMQa3M
MoUvfuv0KdLq2DU6tRB+yhyRm/lM5aYNEGbwfwSK8Rw7R87uco+jl71PDb2hPXuDNkgPaED+oz+l
PZfnmTdZehmmL9gyIW3xzek7HCqgx9ErC6EW1p+gZOPYNpzuDzkFwNNEYrvfiV1WtnYm+rMqCppl
mYlcfCfnIMjHiyv4MwvRLEDlLQXbqtFpr1nfoe8tMrNQ4Vu6GFSirDSSh142HmFKEW+W5zDTkERC
n6aGQMXVL3fVWH5fv8rXL/UoL3k+hwQCvG5foengA4N0a9Bg8WB1/B18AHbMdEwYrZhCu1OvoOT5
Y4kTkkM4UjdsA0tdyg5LH3YjKtDrF0RICm9amPpN4ra2lVUbQjRQ4nEWSNgexm6N26Yjhg4FaFWf
oHs1ajKszYG2tKK7nhTk6bxGQ4qaER9gUakH8MAOq6Auy+lANsdYBchirCG/kOP3A0e0AVkBgWVQ
T7J5Cd5uVy2RSyp5NefQdftSS+8hMV24AX7EIsMxZzJq+R/4U1F+FZP6Qc/nA5ZU1QJJ4dTK/WUX
ZhuiRynGkLQ6vv86XgTyRcNcTKik12bfOZXEPMpYyb6cPXMm4a/8/S3GTnQxRHMLZ/FlS+x+0Qgn
euBfvxo+zprNNEUYFgJR50srbaPhLlGjcMCT1dCFGZjGMaS2DsCJutNGr+zRCkLpSpPH0vUTWIxi
5xVe8wbwfQ1sPy0feVfgplDDX8ymCr4vEQiQ6ZK8IYABnm6gnH8jqupUV3Axk4Vm/wvyuzhPffxI
tLQx6Ai6ASGlzl1ecQ7VyXnMGndzSDIi645AdzloSyXdgPf0VpBwy/O33LbfCbR2/iQu8dbEMEyk
N6qNqgFb043WqVZiYpBlgElvIox78MgwSyZuEHc/SWqZfn520MMD+VxuzuIWRjt20DvVD8rzz2BS
XxoQrkYBy4Loq2vyEeXKUU9tdDFkUBLRDflNAeArtl8QDT/FwbAwXS0emRIFaDd2/OAxekrJ7TJZ
+W5BP9OB6ZQVVZwz8jaqebbv8e8HsLZjHFGQ46uyo2N5+syA1bCEPfTLi7l6H5ffywqx81fG1S3S
3YYS43EDMbwkOTesH64zHZ3sDslyJHmqL8HFDigd79yPTlMAbCnzIyiAfalXjVVLpTEsIDOAWKAZ
Bn9dPeTkIaG8ZDPO+O1dPFf3P9kObn+hsWgqk3jhv9J2fX+p6TP8S4KimDMBkIKZJ4GT7LgYPAGW
t5U+uNE9zo4iH6UAULZuuN+sBBhBQ/2uuxsSJZSGzBPrgzsPt3WoP0xRV59M/QYxX48qwfOVxaCx
fc1jOeIm73Ffagfwj3HhnDBuD/YxQWsfxfVIPEw1vB6g3ACRjPOvwoJ0hWIjMe9ybm2CyeidiUt5
fkQqSkifC08WeMaTijYQxhHwGtmXOG6B3on+08yZYYO0OmBO9pWuK7a9aCZjuy6SMbLvhD6YXCWg
TIacC6dt/jR1H1F5kXKbtvwasy9OO3A2jvEZWdx5mJbfP3zDu1QZnyIc9hbApzh/PwhvShJYeEYr
1HcMlJf3GM/+4/fExRqbMHIlVt06N57EZ0a39Va9QS3pt8Yx7DSoW6iZDVS4+iuU1e3XKxTqSF1+
DoD3DyzAvBxqv/RwNgy7GKt7WoP/lbilZPJwz8gu2VgN78viV8P1VuOlFT46kA128Cw3I4cF4WTv
z7TYFTAFwIiTCEr16LfT6ZGu4N7Y3dR3fjUTNra1Iogz7Zy40F0pVTV+CCrLXmQ78Wpk1aaaB/6K
Im5plqD/2mQYeAZmgviHAT8P9UewZIpKo5H6yh/trOU5DA8XAv2BLTqtGbmJfzrBYRc/3bIEHOjn
A4ot9bOMyUMyBsgvyaFvaVQrik1AziMHJy4wlT+lZFkGdLThCVA8iURHK4yfase34Vm6q627jOEt
Gr9uLnTi+wi67fA2NmCSBtfzPJXvR9u7DprvcEjN95T6kyf9ytrme0R2ylCPncfkaOjf6Vk3xuu2
bihhuif1Uj2su6F7N8BQ76IHb9r2i01X+vpQYJIi2w86oKF/1OFUbtPVzXiQT/qM7LAbnvKyUeVw
s7v/UpjD9zXKLOI0VWkE7nzZU1hDvkFEXYjW54TG82ObQG5CdngMO7BrWVxxTXrvO3uX5hkEKjvq
hymxK/qIhAQVNkSuDlEdcd2M+qog0CxUXhltyBRpNciUZ8XZBUg1bvim01uqjIlaxDACTWMqzgGB
TCU7PUQnle6uemYbElZ0wHT7FAD62Mw/BM9rQatVI9OL+bK2ZOiPCZxU1eusFN/DNwyHyZbRvmqr
vJJ+a9fNtOEOR+P6iltaUhZ45lPamkqRC261fy/khgaYDuMXWI8CfqaNZRzC70FZB6ejxGPiaQ/k
UJy5KK2Fi/KHv7lE/a7DuZ1cp9EUO0HJiDx0xVofpfhSmCp3SFnPxSfukZjxXbPsTEYKrS3MMTVd
zQnlDu7dUL43fQSIqzDUl7i0iAaSjWIQGBnfI5dVpf7MkB/gfxjJbvRhX0pFAzKIlJhHBFG5jVfx
tNJHPipm3ToVq36PafjaVnswJuIpJdAVxPef4n50ailZ4rf2eyYy7sLMedrNrXMifZQQRCEDwTK4
yT0nGlky+OByHBNhhryMDBbR+R2tKLufbAsESkgFEDGxtf2L2KwYE1VCbN4/dcZYdhyF9aoz+y/o
LRtZTWZj26xB+xLe3VjkSZ9AOBYyNOTNN9Ax0vdMOvEP8ynb6VhGrkhEaJUU1adzNeG1OU7D2R+d
148nh73PXnVsO0W3Kferlo9zrSXm9ZbDPAmYZYDTzJbqbPd9Uf68O8RquA3i3fnNwCXmDWt0m3Hm
DazUn/igqqBOrwM2SZprqM3rSRDBA4go3gy5Xd+Hr3mZwTSmVhP6f81hAcgAZI0tL9DkF4xUNa56
jHTCb46f48NnPEWP5swtKtolfdf+Jfj0kUFDb6HaIoOO2UDWvGFew7+iTw9DGU0fJOtu7JC9Rbik
Ym4bbAxv4ONvx14co76qtcSuDBDoAFYLHLunK3z8Euhyt445EtV3e0Ok8jhWntWjBNWsee0gk9iX
9id8lNip/tN55THX5AhWe2dDXIaNNVXB0ahK3mBKh2xB+BlgCNHhgtCK5lrSQkyEyoQz/ne1WWc5
GTME8pINXzAcTlz7PlVLyT7s2aZbRFDPYVToZ/9NEMHCGNngpP/4U7+mExLR3Rddlu61WSwN2Nv/
obz8vJQR5xR/Nv0frIKgQPpcxoBXtM0x577LtFALJLFVx5cOE9oCYTqlkthbt95c7Phwjgpkjrx2
dc9ZJIFxo2N6UCOq6842Uo4KviizgTdUdIbWn2WB8OEOJdOqRxCxtGO7aFyvNGui5SyyHXGx4o0u
Bfgl801Yi2VxXcixIaskcN+BLlUgrOtfjkXKlZn77prQ81LuUdXhov8MvOWOOVYsno8tpbl0D3fx
SH26s0UA4KNT7av78tOl8+64rGic99Qi5YQBuCCABLnS8mTRMNJLW+r4p1w1v8D+sr8NvQcFHCO5
td+Lt2SyolouRBGEHH6gDbglSnoNa/f0Qol/ib2h+gGvMut0z8FMr8gUy3b+oT3Ir2+0IOgQCCCz
co3jP3rmtXTnWLRvpcs+mQHozH82pKT0ZV3wCY0kLu9cFrH1ZxbbU29ZZOree2Vd+okLjy27yKJO
MWQlDBo0ikNbkGCAP9vg4QjJrQ2qMvq0KjvRk1Jd1qkWjcr2eXOC05wH5Xu0WIx6PVC8T07jsjUk
FDI31KJ/3P3IWWK6B4VuwfqT+wJCRw6jgyBG0OQyRbrlTXCmM19wDYG3Ly+Vq4dhpqRgecmNRbjb
38v/8H90MWV69SLY8cnxqcVCBM19UmeUrcR/QOl7ndtrbVkKt61BJq93MdSE/QPBgMFqzfXBAtt+
s5XJHVCgH4sCvr3WIvGo+vSd7cGpMb3iS6AMBpdLTCkX16m6XLy4SwI8Xq4/xYwEHmHjOmo9JvIl
LeOrfnpCD9UnMUQvT3TH9tjPYo66pZMFWDIEoxCGuloGRP7h8QqogqRuvnJ223btCPhPKxI30xtf
x8udLd+Z2XrW4T7h6DIZtiLLyqXeKf+eDdnULNrYAdn6xWA2DLYyazcnj0fJJrIzBBhzc3j5j3XT
lit90Va8m9GAYwyIDTPdVWYA0tmJJDLy8TKSMTXNe8T3ABsh6nrdtr5FLKyWgfxwLtqXGvVAZcyH
QftlULb2g39cg6+mwBDzGtS//d6BcL7Helj06LK8I9YrvdAnc9xOnY/z7sLD1vfq6ee2y4IRa2+V
IJwfOV7nx8G1Z7YUFQ0IW410hudimGtCdIHYnpYp4P5zrKfcu/yscqZCjxPwn/X4F8mqhjOWG/cu
iKnkAtn9exo+gLV95U5wgIAFyG4xtyjlcs/8dYRp7xaIV4A3FsoHHnp7bUaVs0aWvY6YZYBpUK5p
OzPjXR7XXaiPyzghHK+cyM7KYXdWZDmubWkUwQCsa79vkLwmlFgzaMNEda8eyOuQWFtLyimwVLA+
I0U4kr5DkYnWkR228o2ZnNug80v4KyGaQf0+2Ey7QtnAItvFJmzntzohAhLFYLCQcAKOPGjSVgCZ
TgRHkgzxzSBV8jQpPT1rqGd5uhYZcqn/lZacIa8G+pdBv2MbyJGNTRMXhm0RJpaFJ7KNJIPEWFw1
afcK4+WOM+ee4xYzqvEKQp9MVDwMY3wWYVyZQ4qzI2d1P/o9KcySsRgzhDElTofXpxv35P+xfOnR
u6hcOuqus2DoEAyGlY/ewV+INZlwdJc6ayg3RWMsyxZy58rkh5vPhW0+UePPv3A3TVu4ciGU2rds
UwEhMb9ZKKTqIB4wq8o33ZuWRE0MLCgxAErbYlEDY3AwyhIHgTTU9cWBrPnRoo3SKsCR3Qqv+QDB
btcKuIcXwPQutXOT1lbXApaL1bJ5D/hQhEgDFBU0m0FNocKSEsOPw4pMFkvDFCajR1eqbHl3MME4
0sSaOT9cHGh+4hY3xsBnXYFSQdm+JdWwsJAImrYW7MuGADTqrtPCoRkxweNbPisV3VuN8DVVISpq
pP1JFFOwZEDLZva+oVfBfdcgtF2jEilJD60RjA6szZyDYgfHLOEo8nMVQjR6nuV5dFPA4Zl4agW/
jZcVYtCCQEL7nUUlB4YkT9+CiVw1KGQ4QvFf/CEmPoYAQy6u2XAQb4v+dwcei19Ww4HDtyJzz5v8
Aj6H19tBEwkVlX2fSCxCjqicWylUablJyGZFMcitEwzFtphU96h6/df2Zw6HR2lqc395/1EHIjI8
2Frq0CuH0pr926qD7dK+f6Pt0pEw+zSdYThUVgiR+c8pkcM+bPNiO+QRx8jk52GMmXVKRAlyNDwj
VOqeKsjjaf70ChnrglIIyAjykeIEhax2cTmxWt72cC3lqPkgd7yTVeW6X70T+96NEy6/STwof91K
Xk/oL13WXzpAuWyWmnjmxHAS/rG8LSZD8CtcVW3qfuHxX7HGrPhmI2AWtc8QcKHDmz7sc9ZiJgbt
G0whkE/vNPUOR/Xs2F+Is3bVM8RSzEMS+tZb2I2bragF9SdHveZR5jQmmerWUvKgDDA0UIwW5YP4
O8mpu6gUQilcFV4pZxv3iqodsjENpyyy4xEpYIHVK3FK7yv4x6K2vk7Tn1v/+iQVITUIgSK1QG9N
JIF9MFhobakBa/GTgUeJLSF87Qkomz81GRlquPHPwguyfAgfNqFKNZZk3OaXPYoVjB3vvrlAXDTW
z1WsB0Yyga/lHYOqPHWX5FopAKUm6OSzlw35PkEY24X3qAJfWjhbSH0+xyrBsksdORwYA42poAZI
Wo8yiAOn8VLFxu26oVYmqYWHxvFxzxvIViSx4pSxy3wlsbwEeeICcmhGKF3OjgajNQPJH7yS99gi
2L+J7eCXN1/x2T0mFxhke1yrf8hFz6llg/izle1nQX8A3GvU7XmRdjeR1p6AYM6bJqLIWqijEp1A
PWnEcc76lW9Zhp8rvXXnDTA2MzUkQGplU1HZRX4tYkCJ6nV+T1G1HnNHtrMU/cY8y2EeJnJUGL9s
saaprDHaM8vDdNAeAnxWdxn+8PDLLFfIv/1VEZnjG3J71O4EUJwj1AU/7GZqXm/qUWzz8U/W1FJt
ICUMfc/CgMlGLCyQDT+R+Y9ZOekSyEEY+6OOwcuMYsaCY5nkjyO1Q0+M805V7sHRD6F/NkUqOH1e
UoTFAVD+Updp2lCFtkJfWoEuiF3HtJCnu1bx3UdHez9J0pbHOY2QNLArlXF+4yL2lCl7awW9EMTy
9uJuJBRanuXMly2lrjw1RfBBhD2ycqGIg5nvB3QJ8QGnjswlyDycbSYyN/uRtD5m/sSMXLcJ4pAa
hDKuzD2zXUaHY63gNLQ3QoLR4Z4+wYiCMF1E8+PZEtwXC/RxJrZsx0F2/wcyo7l/s+yW9m/qwFrn
CjeR/JBFrmFO/1qbSEmRBzkJL66is9zliBqq6zjJkaVsgG7J6y1QP1hk6SN1iRGD+qNaFmUVRKmV
Iih1tb6RtDyCSkqEk41PtiHv3w2Mr5HO2IEx5Jh4P1U/H6yGEAdkJc8CZmZQewKQYrENCZGa1DJh
1JdjFEjLVHfhE93ifWRyJ2j8WXdW4ZhNnrSTdrL7dMnDC+sZcBFZHeTDWXcwZG9xris7ZLc26OGP
VBdPtFRx5/OQo2uWrsU+EJSL1XpwzS7EYkFJJ6aW1f3aU2lzTBTFR/q0LXYIg6qXqRBUZiysyUdz
Hl7JptV9xkVSrV0BGSbCFIFXUc7G+9rqsEZwupgep/6PbXIjaI5N0lWtCXKF7Cx6nBJ1eTjvDXnP
wKojDfWPAcI9J6ihS11Zzha9ZCVrxGk4BFh9CeDo5wFpLKo9RRuBJ78ompItd1y5LRVUzQLBSY69
UZnZqSlVPiIsDxj07mkBFzdGKWCsfi5krml/VodXyEI3fNkO1VQWUYsQJMYGi7gJT5iDLVAskR2f
kho5qt5q0u86vzCVDePVgd6w2Z1sogeXPvN8IV7/sUC6Bw9SZOoJ9hEq+Uq+f/v/a7J4Jkte9CeT
ee5tGtg+eFuL8ltSnLUsg+DVeYqhc1REhyaEyVdHhEFYbtXik5ihR9mf4L8mhcOlTdWK+CZzBTm5
kPMtqREI1gdy4sahtxSqdI7gchk7zWKdpKuo1vi9eMt/KhZtrpWlPpgpFEBTGFxbQEP8foilyYaf
YfqkZTdZeLR0sPZIr9nL2q93dC08PLu36w9bXiJ/Bj0EKHSH5cfaFw0yRB4L0JrI52/YwS7vqyF7
TO+OB9LLKIO9AhVd4VRd3rW4rHPos2Da6JfN2AZ/xVk2y35wv2q93w82Lmf/Z1bj1T83MPaw5ZlN
bjSrA22Nh3bmnb+TxzIdBt6ZCP44LOKWriGw6f2V1z42i0Mi3tnxcqT8RNlhrAQ+wF/Q/aDns4Er
R6XCa4aJgqfu/U9afT2hs6KD2m3RqiQssy9Y0UkWwDMiniWa6h4ooD/XLASoQusJw9iwN7eqdOi9
IpIeWqDd4ATLhbUe8U/6JVIOcgE94jUmh2yNjA7QgaV0T6EznG1nIasNQftHhXI0pD4fpzNKeB6q
y+Ne1qkRMxLA1TJQuYtf+sDFQ0+ZUNjDEsf7oGYnuHrNzmpkruJjTCp0UwPl8n0Z+ZHd+7VATuk3
2ZD5EaVvyptXbAGWPYDbgdzx4W0NSS8nbl8sU0RCu7S0KoNzIEqZCutoqqnIiXLZvKOXGTtmq3xi
eOx9eZwxgBi/EARpVXcQW9SQJfs/OrWDef0iqDZp6id/bcM4+HdEskqz4pD8PPL1n7DtnwolNLok
ifrs5FTCBKDFeS/8hjG8eMi5xSR1vkgpw1ZBuA0a9QyVvDAATWfu2nMg67IwJk7u2hMRwxXgsKvW
8amiTzUYwm/n+ORJek1ltdjOLKpphYFlE3Xezxnuu8I66XcXXDP2Ye1UfeLveNBSH3fSfDRUca9q
2TngFI0IXW41ZocA6ZcsNxEVSawkD6I/720qkzM67B/RMNLyMH7Kn78UekCQ3K82Lo+qcqnimOjH
BZwMBXa23xPoNK88m/+u0yFnmJ9U3DYqpZ43QadG1n9emec2JuotcBUyaZ89Tg30wJjCNe5GwrSg
ZTSPRaFEzIeVYUoIq+uXjfNQSDHkYJa7JYQgT/mcghGpeIqXf3JJKEhOK2r8ZKJDoIL/OTdU3uyv
0Bdpewgoibpm0L7RYXP4WzoUNhaVrIGwRDj7v9KJGl+XcQkH2bRwxXd4WNLe7XymD/EgssqCQG9M
SXvTmH+kmCUwlVDQxq2lvKtVUo+ctHfOVrIZrZ365aLui4N9LzNsaTbB7PfoFfI/wOocGzv5jtts
51mMWzc1CRgckyVpYM4c5Zj2kSxyUuaRrI7ffcH/x2tR+puPqlaGOWo6Nrli/pu2ej7Zw7sYuxg9
LljxniyYafHjw/exGSoWPsLL6WIXOjra+3I0xEhdjL2hPaIPVKzpPcjTIfBD4huR5jyWjqxN4TR4
Nsw5YZjOpAyqPN8ErhBlEUQVhPbPOEaWJB5b0yNOzknQiZK2VGinAGSmybl/pJakYSgRzLoct0bJ
GBA/Wk9tDiv4peKnZL0Sn6/jI+p5RQgiyGWGdCl+lHgtiyS39UhS8szd5b1tSt1A8UmXNwaCTh5K
UDBOeafUOZos61qWeE8h7MiDP1BrNRSV2T1JhMPMKtFL5b28R1j5N8vMfuw1ItDX/h0sUJg7hgCr
cMnFmIgGwDOEM1JgbTSvW/NZWowXB+lYEZuNdfFEI9GwSgpH67C5y36sz4kNSgl242EJMCbMrks4
rBk2oAIy/8NnX/X03CuOVazlzIHZTgwKZxhKlgbsEYegEF68HtdBsD8gf/VoIAlqmvVagYSTl6oC
G8zdRsi9ZLNDUcaW5ld/lXM76Vu2Ocg1hd+xavVNU/t6mxXPv22J+mzwH5Tbd206eVMij9KJ0Cl4
+RQUhy3shTQfYDmlWcf5A3FRqr25Rw2mxjxtAVJEh189PIpLUJln8PEkKVe1FPbNRms2KWNqYlY+
PRmNlwEm71O+1fvZR/JtK2v5FnuslxazZzl8eSlr0hPh3fbbHb+HoQmZXPXMyCYRT9ySeAY3BgHx
CmiFv7UoS7abDCvC2XExJ/5pd8PGxRx0LFnoI/p6txL0ub5vORv0n+QrvLPgF6SEtIgoOOP4fdhk
Yq8N9lMq8Cg82nGNXlQWWNOqpmWhjqK3RAqZ7hdzCIb88eWTPvYUXWYON1jFya8cTCpFfOAS6JYS
XNxpOIRhq/kjvsN2uQSwToFfa65Ptr3nB+8b90QFyXbvSbkOPGa8ngTJxaPjEtbVYbXH0Ci4CDg1
TQVu2mBDjYEp1Zum0wC7vUQeavD4ob5uJCVkLlqAxENRA3PRJZTEkq5zJsMtWCEVP9f3YtW+Rzrt
SnnnZsi+pPOPH0qMQfBlzeneg6EK8ZTjfs7+NXRtH8L3ROlHMC5WQTefBXhoI+za3XINhhnkdUpQ
hbLkZ0whiddEVl+NTAsmA3vBdCl6q3BqzcxdNlKifrGT6fnW8knWA1LTHXd1k9xpAo5lWzZPX8kx
eHLamP4grizUN7ki/re/oD4hAqAyP4WhVdhsCczZI573NtZ7b9huLK/TFuF8rFGQIl9eHqS2qQy7
x2VW4xGFCwFWKLa6juBX/zcGAU2MHHXbA3dHspMns/iF+/ky7j0HrULTkoKhuNkFaWPBYN7CDheb
F3YreJUD4oKC7jhDk/Ou0wxzjt/0ht36R/n/Pz8Eil+bdoBK94rdAUl+s12zRpLzSb5cFvAT8O0Q
vtxtMxVgDpPEKF5jYk6iNkv51hBWtPHq7IBiAO1Ja10IGcOgZxFIDuHYr9FbXCJm8W6II48No5l2
ZnbYo9pZb7cEo17XqBHEVp6eEpa6wPkNXM1d6d7cmWqQTKxyKiP975LYzGYFQtTke1jA4DlB4pnA
xQpQbGNQVARR1bUq3a3/2BPfubSLFEZjdWvcRKnKwqMwkYyUETtaffiHNYB/QtUvVQjz+30EtLID
GBchcFdpnYwxyH+jhur/mEFJKar2XnidgA3NBHZN3yLGPnAO6WgVZjQ1tKqW47wVKLzsAUkCsOAe
LxdP/4cpVUiUvDXfIdC4IaY3wC9ZwRjGwLa4JdTdvBTtARO1VHI5n8ytZhe4fevuUBznQUM8vBYm
5IFPUOPVPzG5zV6CyC4gCkgt9kigi59rRSv2PjKmktJoTAQhcQdqzEqfeAU+D05cDtckovijhXnI
q53HMLOr9q6vw8BxyPLoZxFcxW9UNIuKsfinpetz922HjDIk8z6OxdB7o9r9OMJyxkudoTrmvlmC
KHTHJ+LhBbOIDXYANWFFxA4l1Pwlu7amo8Tf83KNVXjFWOLrULgF265nWfkqCKadiP1rFiO/VB1l
urU/ihaLbFmZ49wpYIjArniqp8rJForM1Iy6pPl/4Ryp+82f1H2V0z9GVm95kZypupeiCQv2OWfE
XBNjqqFYBPV56+kjmd/iHHaWRte14qJQzruLBoEgaBfwpFD7cNShLCp8EHuaX3THJNfLNn6ckyc5
xW4dvHN8E62I2aNXgZq0E13Ou1ZVzXFNakUZ2/J0UXUEf7WdkXNckXpe258xvsK5K2SsHgSXw9HR
f6E2A4fnNUzSs7lUAwZkIKYnnPIJ+i/Z1wLnr1tUuGjkYyF4skJnN17kkr5/j+dgPSwGpkjDOFR7
By4UzOgzTwWxXw629vIZ08P5/y9LDOagBvqtVmLwVa+SJtHxALDFU13j2/dXIGWPzeLLrxFFZqUI
Er9J9IbUT+tA1TEWc2t7WwPtQvr1uoKM7CSSxafofhWzx0D65wLqWJ2poGZpWFEWq75c2knyhEd7
xAAwP9UDi57p39QIWdiWFpTh9KqJHwI0rJ+1PQE+Zczp+LNxlcmMB3192QB7vBEFLNsNWv192RG8
OdCdHDQWiLXw16ceQF7UM5yhTwd2PhRvu4vEwUF0aKrIzKiUN/dp2n62mGPyNTrWZsfZ1Xt4u44q
SHq5KSxtaa7k78ZyHPXkv/hQab7KvpAjXz9O1Ut+t2dRiiKM5goblEOYVECcnxQyzjKSYhsiMrVJ
TQDepKN7FwQIrhSxsDSD2W2ZUDIqNkh0n+WCLXJAiniGZccwHNLExUL1sljBlmoLzhyj0VpQFy5N
3fx2x6lg7rqM6tk0soYZab6spqwvyQRpC/XU8+ZJ4m5YYeH/hwuclpVfSY++vP4yZ1LxgvMndHNr
1p5gwJ0s4Rr8XwdkL9tLB5LhCJHnCzyGOVVLhZvyU950u6R0STJEGoBjpAco6FXPjFMO6IjxAwRZ
tHBM3EzrOxvJOagYaeXoLkDjqOh+eAHmyePmY4OqwvjzkLuWtyIK9M62SpnZRV5HvCnYJt8WcJBR
r8R8mbTqmNHK7nD5KW7F2zKJyN8j3WL4+1VUFHSTNvS5oJowYEgPPfJl6FdUoIEP/Xh6Cvt3HauA
pCTSA5lQ2zpT6he05C7JwLdENyxOjB3fdRy3A7d8UTvLj/8LQMIDqQwarlsQePsdD+UokLHYkJLP
1CqnUTJtiWo1gY6Auw6CCIPTlBSau/Wao9MYY6Y+BrEJlCRQoL126TYXqPybpor4dhPl6h9xC1oD
PmpRalIJAPJSFZTSY0eVxnUNW/s/b3++5jlNfNBQU/B73SbxcHqhXi7o3LLP7IKR5mTKuC4K6rzL
dDFDK6OFkJuEr0d7DfWZ2A+i0BvB1bXyioDrFSSjCJ9SRJjtdEIZ5ZOS8pB8MddArEuMCjBDeiX/
4rcbzbKv4BnvMQSW8I72F1HT3pUOhzwKrE+3nYu+dlcpjwwQefilIi5ThP971S8uKSyhRjWvkC8A
4d2vsljYhaFHUwzqEHv/z+t7s3wPoQLjTGxrlHgjVjfbuSWCvA86kmdY8scJLeLkJzrApHgKbSsc
hUs+bEZUbsUlcHqpscjik8s5K+1lWO9tS+SHMy70imzF8yYFbmwLdoH9Udkuq3ZdK5WfML/WtQIl
FURy4dIl9ip4YUwvDaMJX7xXo/uE27/TxSO3FzJkCQO3ViWHkLkJojaGy6VBwnZPIl68S71gy+FX
BD/r4efPS/Njn5jr1W/IvAYIGs75lE/xILDwW6dSfWvVhvfmhp26lc7MDQ20KskjPVVHqk7hhiob
rPKZYW7ZslOYU0WAfpZL1T7Zstcf0mNSS4JYGmIySulU7Wtve4V8i3IBnROc9n/j38pxOTCgrGBP
f01nzR49YhZT8qnQXLsfK+X0CfbT/9zRl8jSZQNEykheetJY8slYye9QnD9lmNXvN5LxdvHQT958
fOmoHyIfMDV1Cwm6+63YIIwTxByEZkYvGh+mtOc8Xu/XD8pZxzi7pdFZwkIA1EfpZ3xV5He50duw
HarLTHPzlTPmJa5vbzJK/yBpL6NPOUCypwLbi4EIlnCEw9y2w+QUs1r8hrXJp17in5dQHIFvrHSB
DIk2uO1FOhA45WtHqFRoWlpSeDDzd+OPDfNkHcNDTzoQ9lYrihIjlHm6bHRWIq5Nmc13une44TeL
6c8WZ9Oe11Bx9JTHcBD9pILU5OPCPagfG2vxadNYthap8A+Ay1EIz9gb47AuvAiUAVqlqe8ff0X2
XhQCkKA9Fh0tpGoifKKqV2dvkQu8zgG51GR0yDNN4iAwM3x2LJe6kySs/rXh/lG5y7h37+Dq/iUI
QBQAY3dsSlqkoFBmqVSwAuqtmt3TiWI3j+52XlZGPZSadFHwmilAk07fVrydhcdRGM1mvwBsxCsg
LJk5wj2ronbwwQFv1L2ZsHJeq/RRxRU5z7zWcW1EUoITsArgpBSoNb3soNiZmDczru2oy3zM2erC
smjFRb7Fh6kV2cvUDCO8Nx8SwJnqig5GX0PaCMKdpEGiSMtT4WC8O4toTxkp8xO/UAKccklgvUlx
+fQS1OYCQeIhF4wEIYsYG53/BTgedDRadoPckhWsaIQ4QiADl+Oqxw2x7+l0Z5PN2buIOMIgFxZH
lnkM7O2ZKLILZnfhzjnQgH5wx5vibwlF1GE9ASicQbrM7nLaILOt41hCEnaSxtQ9xtEKre/GAyTu
tcMdn7aStUmMXpy8JRKnIW36sQIGdZjNDcxEugcXbY/fJZOf/0jGRHpX2uwPNo3ff/jRcl4/iQKh
t+Oa3lXB1pCGHWa6VW2CbHNjPEbuiZg7tzFOUlq2ZfDFz43RLZwspbMfHHgDy8QT6q0auEboDhrx
e7VOEI5P8+LT/RlPSCvbhz7t0KgIF/CJJD8fl347M7D2HML2pwhKfdlVzFqvw/hKDIcu3ycagB7k
iVh95Mlox6+Q1Z8sQDz3nu05DpFDM9uSuAZv75OrQC0+im1gPJYwsnpJUH0xMk4UU2tGW5vyG1UI
GzEXc+UFpfsfN8Gt73sdNHctm5XHil6fy1wb0yYsuCvZfsaPlWY0NyrnWPV1ticw+1RFTWIHiB2p
j3R6KvKzncVrpQEoTc0k/JhLqAXrthL0pu6cEwn47gAtCzn/D79y1Z6bbSDq/aCqiRkNN5DW4KJI
5lMufIc3OVIgf3vidPCYhIKCQbs5Sw7KEB1ACc7C81qpof+wMQPhUP+bLIa7EU+paGmXm6yIDWpA
m2rsf1DOh08muJkmlt0bGZj19NOZGjWFJ2z8z3+Yx0+9CN1gikcRztaJQYPKVbTJJMvupQQTwFMu
QJQca6gruqON66ZwNQwhCltelB9QjRVR1bZeHntP9IWU+fIq1K9OQDXIhQdFnl/3eMdeygxxAI2Q
vVsKVRrxw3Fp23GPfQfLcwiU4vaf4BDlrjoUc/TyNO2q0/Bee1ROZxz8ioexMLdTAIK6MaOE5WJp
SvuPuMsMtmeYMXbyWhOQQKFrrEsFCEYaooHX7mWJcDn/15+fKkdKXk+BGAVbhY/RqIyk2X0wl6Nn
z83I+UAYNB5xtUFNpyvbL4OcNwsntqlXeeaCXH+NJGAN/KN61SApzeXhZqiupFwlxfgZXvjN6UIB
VujkwfoPtt3gW3nxx5F/ZF45cofWQfAr2SRAqzr5t/NMZDVfAWVNQVq11nPMcsKkaWnuRsrlZEUh
DPd66m4YBMi6pdyXHmmqkJNYH+ZCscBrngy/9G8xLSs5wZv3xumYcmnUqjTTPN8k0yxMt1rzC0ct
6c4+CJWeh5iDCLrTHsjY7cqNa2T4rfYrtIgWi5Q/1tkJxKIBQYxpCgwn6aJp6tAumIfujxB0MAUc
SPDXj99KpBjs0Uv0xnRi/ic9NljN2XNDbiUPphe15cRdoELOuWSh7pFEcBe31ElHZ44tSK2Zl7nx
U8Xe/UHVPyzQrqVA9DmCqYqsAHhnZeWubsMLRzlp7TksuFCypNJ+fNML/Onwa5wXJiBAo09Vb9zN
GieCqT73doaLmkqE3KzrG1iaBOxN4RKwxvOl6Wc2sNtWv5ZmhsYxqAL/9L7BboW3szbUO/diCSZF
IIuFrw9syJ1IcIJQ5s4P3u+jV/E2uXbSgHuEcoU4SeAVQL+APNPvFWj+Oko2Ynr4/LhmKc5tyXJN
PhUksQW33hXI8DUjJhWsUjirPNa2UlOyKFMKPKATBxEoFrQyKQoltchTdmQ8YWHRAHzfTW5fkAhH
NktqEzvr8U5pdoKrGkfEk2sxOwEpZNwKOvOq72Bn27K0Igt9m115TNmGZUiLf8s0o6JpiziGcPA/
cQ5cN9x+hniiNXvaESRf1U7bpAXAHTZyBxxLjpLaOiCoMc8AdByKvb2kwqMNrqxrzi1gnPMknJ/F
FX5dasvfFqCDtZSUlEUTc81EKbxT39ecDsv/RvnMHGpNT7iekLZSb7PK/SPdYr2RgCEx+nDNn6bl
K0LioD9G3hkCQra516kgs0h2yqk8SkFSefEhFNzhotm5Z40mIC0qLwKYhrcE2vcR+Sqif8ZgYVHW
3CZf0SYhQQK/z7y7csntWfHCGLEtKpWAhywaaZZVKpOWU4VGjK27w1b+XM/7ZxFhpgVmjskmHVK9
5hcobU5Li21jdEVR3AhE5wXUO7Df3ezHytrGOOxjeiSQq+PhDjLMLsT87l3wzfOgBlJ2gdVSHuHZ
wNPOEf+zGALGS5WCEl5teIt5U9llCW49IK7l/DBZWOnMzfkVg6pR+1OeLB7ADb4VrHnvJSVSmNaV
SaXhBxV/aFrtAmjj9qMCyH1NMcbMuOPVWOre+EnaFfAr6bosRnOzOejH45UwgaLjXtuyEbVgocs8
bAkMyIgOSd9j+8Z2mmEBU6T6VVCMZzncHFHCENAfOD3/xpev0/TTVN+Kc4ONc2GX1cX8eTi/iy+U
1QZdTb9tbRrzak5UE+EKsPEEwtkX4W3+HP4r2vIsAmpF09XiopQIlLCcFNY4FF295ODmtJBSUrhV
2Is09dE6eCxVvfrm8AVw+DG/igQ0fb/dgap0KlGNiJMzaxY7hg4Jam7JlIfm2XSDpr92A35227PY
eIPcZl7MEoRx1Z1TnGc6Sld+sCDRkfFjZzIFtT2OrSksWn3v+uJ1h4xUAHmIPC+4hRpZnbH3f8v0
MI+dbgb5NH4D50sGp/Oc7LlLzMtY+TKHRigGgowFqOFnesgN7MXwWyy2cqwpggX3ObT2QlI3P9Jn
mmFYzaYZfDIR7YHMI6qYjeXyRLUtsShHlte63kIy9Gm0bA1VLaqiMjk7OBbFumu1a3ndqdxNBUhJ
l/VTV38JbSlDbI+mY/D/f4zC7sxW9Y8Ta2cdfTsjh4mmC/FrDWZFIQPSO1j1jHVhxHhytRhO6jF2
JrEyKu5FCz7J/6+EP9nitfunMwaSfmlnrJYd3TKpTwpiTQqeQiEw9I3c7r0Q+syUDp8WFO09ZCaE
ZdxEVMSEICKrsIf1Fx2YKQe+eZt0XkKAIc4O24tguuWAq2537lLEuUuZl3poivpr8tcsBtaGdIoq
abnnfRhXdeq/vNQoi9zOPlBbYZkzlAJIO9cVgN1M0pICAULgUpDmI1FBnWZny+EbCO4g9dGhNZjR
EeVUjr1u9d6/987DEZ0f4AvaM1eXvoHn19BnPT2mGK9LykrtmNv6OpV4KU8MOay17rdgdG3QMMAo
qlIID9n/nChr2O4E8S/aFSrBFKV/xMKPqwZus6nLgy0InBMgtO6EGbGVrJClaNQvfj68c7A3AFKb
oEsEk1NKsoTv9A4a6mWUjimRaBsKtrS11CCUym4bFuEmepiPG0VYDKFEZie1cqRi1DQaKppDqf1X
TIq7mPA/xX8F/uUT9nR1dPgFiYWaULEc+2dzp8ZumECWzc8YnIo8v0qBqAHjEx47/O0R7g3mFmPA
lxzL9i5Pd0yCdIefxueV9mMu+lWwE2BeNSapMTlw54rZ49zu4AOBeKRn2Ar+JAJa7eHPJ9gLwEZe
l3r21Esej4rZRcCbRs11Gw5pd58nUMKm/oyxBa92GiPIYZnRwbdsP1popcLQhklITy3DhryLIW1/
grZ5kR+BXyeS1axYms9eTLkTwlyTFGCvnSOFHL2VqTmP6OKJHj5cUFxEWWwCEcq+7jOXe4v198nJ
cJm+wtGpRIGXlU17HRnLURs29cZA199tgs0/yByIuDeiwTpHGdbZenHNjRvKleHxdF3avPk4m6s4
kdTAmAcYQS93LsJZ0uba/rF0IHs/TGWwgfC5dilkjUG1tjCcfiIt1/qMleghV45FHO1d7qSMNnSj
FsTTzCkqbYnbZrSk5c1Q40NRNQ8F8qDZ4Th/G9G0EUTi2D51S1XXlKSuI6jX1OiN7c1rOVvK/N0e
1nbXIA5rtDQiva/BrP+LlUofvI/Moy/lswnRzTslBGX4x32fz8sNpW75Ib0c6Fy2DNixBxdI+8Uv
2Ier4M7jOo5BDVb4CqrxvWqnapnKohbF4MhwcPjJAAEek0dB0HFCULrKYH3JKjc9zx4o9XzvjRXU
CSFYQgIPaHUzjr5O0WrqXLeAAe08ldDz+XgHhb1IEDTkbSn9hekyXW2jiSIARCo+ZGf7TG0ReYf1
baXhf6uKM4d1Q8Oh19KOD0Qgfg3wchuI3T2SgkCDiz/dhPwaa8OPfiAE36K+tFEshIm0k/Z+LTZI
qD+QfBdmw2f3h82iQ7FwkvUUBO1mQEhDBFIpqqW+Y8WlsaNviOAPSDWczfSAuy8QGATvT8QIl/l1
WOQNBiYmoYHSxRR9lMAMA9ojhdXhZ4wzFTU5ji+av1/J9/fGkDYjuP2Y6q1BqQa1LBLg0eBdLac+
PCvN+WycqxLWOrLZh99+TmgHBVUhv5lHyjc8COUeYKD7ryhJdANJaeNG4OcByyfUkXdzLq7bnWoG
MNKm6N5nzJe3zZNWKdBNLXkg9b5dLvJvCJsJ10cElaHZsP2B4MEY1jQQo9mqchASe+BEp95wbsG0
eaYkieR2EnFC3JIKLobezjZcYWiC5KEENLZdQTOmFxbHAaB7saaurO8nkcKM0t7cNsT8nP5uD6mR
ei2LqcsQog9JmidL/xyc5/LD315QSg6j0lniLUdpOfajTGpJ5+N5xqBWxQqTMK1VtyFLTcJhTIwY
GH7x+L3mhkzzJz5v3nWu/di09o5JyZRLnn32dfEX3SmANcMF3brFnHLpFbnIPYzQB0P8cZH/Wqpa
cIKIDO6OuPmz5zwusyXkuV6fqVR9TdTVoS1MwXX75J98fDPTUsZbKgetIch7KKPYgs/Q4Ns5hVeJ
Je8lSJ2pWJ/khl4Nn7ix/JRGrSLFYjMfov+yLt3FOJFkyRQF74K/Uocc75z0F9si3rPifN0QILZp
MjZjQghpLINMrGj3NuwmuRiV/hCTpWH2ndKloYJ52L62fOtN1LnNo10nTN66gaOOKb1lQzPmy2mj
UE2qoHhKMYEYrowZxcADM2YLavoLK3BIG5qB9LH/AcH1UisE4/KApR4DDqYNJFOSSuI7Mm3IzFP3
lX9m9tlCM9JRdCaeOaoskO2pQGbPQvCnzGjmUyPwL8BloTD/5BHtow09oNhMSuLxPNlWO22Y8oIX
WBOeQUvSaJXUcxb+m7vxzTXY7Z5qDQtIhGDfy9hDJWc7VJSoAXvjZLQ9BRy8SpEnvRXv3XDvEZhE
fM/9qMnt/bcR5X9GAE2+A/VCiM3FZRYD0cqHMDkNjFu6IKH7SRyV2Jfeh/KG4dMlsOEwM6Iyo+K5
VcMgNScpunrt6o/EkG3vy1MogZcEhvgloEpXMbkSiXzoy0h94s9EJIMFeKFomjA42KxDVT1MUzkr
p00SyZ8FaM4nBs4QHjrvriO2V15Ew8DUtZNx5OroT4hc4IfWo5houly4jk68Fz5zBc7WnkO/ltKz
0Oy86SKa+hJgDdUJCPlFMUa6Iyr64AENScNsHZRQxFLedHQTbQLi832HLNhvVWwCz0nyoXDqdNKM
YVo/x5ZsXcAyItEcwzAjYmEUjciEbz5U2RYFzUebEgAgWnN+sUr6w8Z12StGQHKfsx0lXwycjZOD
FqfnIuKXP+H0mobXSWOrvgrcysZaKjCUn2PVlEEV3IWzEzYa1kx776cj9ioHehDbkR6Ri4TgwOa5
xhJnsQkcHamg3mcxRnGSIagzcNwM8h52mHuX08w799bSCqIqxEimC2ffcRt9XcVYAKcGYnFBPjSM
P7K8OIR6L+lpeF+pI2sojB1TGe0Z4ZlXB8UomLeJaO7ecyBnqroovbUqytBEn9kCLwtuRpeVtDPh
KK/lL4m0qyaFly7iXSlqvajgpXNLzfr+s+jnFiPW9dmjloJhv6kwobxr0msDSrd+nuYse8aeehb0
NfWZF1PFC+hXQ8ieJ5Q6bkkG1nr9bVktZAsYCMSFZ1+cQHXYmxamPQ0xDdejKRe779qA+VtaqqtJ
d0HaO41qhZElUCu3JpULXmjLOxm1YF1tg/SLOdANRUNQ4orwwPrFLqDKFYv5x1PkSjL/sibmgpBm
gXAn6/NIGYOaJV3FJF+3atd4VqDma+BWP+eQwhIrpZN0m8BvflqkwLWqjmrrVHXSv2QJppa0nxeZ
DjlD+ecI6FjYCX4Cy6cEgePe7es/cxp/7JVYR+ZKVQrplojdgiAvWg8t1N726oHaEMGarp66EORX
sjqUISsQ+GhDkxZxahSLDY2vtIaG4LO2sfK7pUmdSWopVhlOMez19T3DmTSQZVfls0Pahn0fkuza
2o531v7FRMuF7XxHyoxpzq2fJYUR3tywLwFRXjRK1Ay+WILBcYWfJo+4s2vDJ1YdgnYEyj5Qz12b
58+TIHs3gtmNMyPNGCJ4f6CgIDUrP42/N9d7kERYh02+ZAjOSR/tf/eLmEnmOudK0Jf9p3FZQlRz
PLe9F8hQi7xP4tSAEyaO1mFhqJsg7/+6QSktnS6HVMTOVZwXCCHe9FQVEyHjE/XO2WbXTwwA9ogz
CkwVvjNBn3dOTGfTnlXEQAFY62AFhERQnEVsL+fB1HKMH6iDw8PlAkKo7LRwDSao/Oi9RmMvM3u2
TIac8nGTJc1b/YaHj/txHSxVTWDr+AuGZbmQrW95hn4NTTviJzOHf98H6ArUFBMHGmhD9jaOjcu6
lI3iY6Eay93zhrQRCNw/JMmuJbT1uYTWhDIR+osKwm1ascYXdtxYo8SqeyF/QZo4zL5IG0dtfiyZ
D+tJKQu3TYBZsBv0fYW6q5RbEp5axN1iww4O8BK/LGsRWlF5thzn4ruohLwViZzKsRbGCXEgSNJh
oC3Tb2bYNXP4FnHROQsT5eL8jxi+M3Dyd9llqbEwzLt1AnFv7b4gA7zxcikJODuvkhLvK+u97PBI
tktbbd7WTGZMMplmD3rxklKB3Krp1au0Em5jmMEqwAmEUAEexWGIrifb1svRkDIOxwoEbR88RmND
E92o02/KwY6tr0DFnalO9+e6H+CSd1iBOaz9nkmj3I2DxgEBoKvVG7peGPDJ0SPIfDzoJnGTGls0
nn4+BGo0Mt2qQVmBobIAsgIF9MncOVVB8tAlj6A+9CV2xF2bg5iyqIHA2tJ91Vi6b7H/KcIE+33N
DPKrbnLb/heLA3J/qk/5ew6ATqzgZri3eBi+oq13uOhySGzYFpZGs126GDLFYpHkuyfYzFCPuNtz
kQTLBZyZUygVPRcRiYkw0tI2mUkFcm3P5+0zqbvQ5xAnitYkAwqVLNE/AafzAxoihrLs8MnN7xHP
waR4fIVta0BSg1dMeSq6epmj1XJKkoRAry+UORIPBFjngaYO4E8f9WNiCbJ5zpMgeaL9U1M2ferV
YrZPaq4vQY8pgwDg5R5gC76zxQEBpp9CU9Zs9m91Kcs0qCcijJhFLxhCnU2chaSs75B9XOJrS9gX
GgWyPHjKVxd0jnULZoNlygcENDYU9Ycj7tIf/rWw9wY5hVGIJHCfwFC+0KeLLR+gerq0LfxB0QNO
E1hTG6nrLnKi5xR1Q7H8zaPQ2RTN3ynRwyebZBCtcgSTj9ILUZ+EbiQOapNgMN+Oref0n90dkRvy
aH2qQhiKwgR22wmL/sRC8sB1PKa6ca+YOykEy22OzsNo+bAo26KLvBgLV1DWw81kjM9dhRzl9pHj
SLBropH8oin/17Meuwh9iPTRWbI1y2pYJljB6azWiWY3iNHktpB9j6cGxM9NDf2WfcvTHr10guhA
BSmDa2eZn4fxEw9xRdyEbS24JFnh71I4hqWa7MWiRTNBxQ5TSflFm/cLO/FtR4ej6U/3/8apr8d/
hm59qPkJ2l72npSAk+n+R/X4gzdapQfjqPIpgyaP6TEe1B+kWCCEWelrbJLUiuEtIB4HXhHCsy7j
Xx85N3NMW3yMC51seuZCm3GaIHittcQM57eBrPc+zafKAM6qkP4waCHjpdDyjewc+zNPyJ+7lcXR
pkChZ9CFh37KfMxf9Wic6lXsyzReLUefZMe9ZXfgIQtH0VWoYwKZUWBl8x9oDETjOlBRXUAQnTjV
Rg9DOAvNoKTdQIKOErk28vsMPnl+b8DwAwcgFcvkMJU6d/rwxyi02K4MonUE6O11n/rT5D5J+c2t
OVhCNyKMo/h2FXtMpVGDyogLRt68yjxWxdz49oohZG5k4I7Ls9Y+7xCUiTiWSzVQx8kvmhWRMBZB
eRJR+hMaZM3lsHS/IY5ADETm9N6qpE2QAFgsn71M7FIbw1gPL5wyY6nnzagQvPhuBQHt/NQAt6eH
GAx08bnNcIDmlv9KOsPZqU6jUfJ11AWv8Dr17UQ51lrzwt2wq52hHml8Jwjw1yUfCQYjOjx6SWlz
vBU2qymMN4N0PisBBBsaMb18kK2EOvoA0+YrMiGlBeWhahS+Ly3eHlQ+A/u9P5vpQi5ZlxCNGC/r
t9hkLJsdmkBZtSrEr35adflp8sY1m1HG3TYzvUXPbNXrjM8Oh5JbxqIttABrNAKt2J250NMDUu2t
R7KpQslpK5r5fy3kjkJpw3Vc98ZJfLpywvjVQ4P57EFdPzAA5uUILhmErKhvWRWQHYqpCFH6hDcH
l1MAVMfcimR075jAV+qK2eUfpK+Ozj0l/TlAPXXfOXIrEDk6OvVZd6+Q1U+Zk1zrALdw4KYUYfDc
gNA8wxgDLoyfGOypZ+hDROv3erIyQFKCDFEPAAYZ3JpGlJdjQeLmx9kZh2Dj8RqodIWIZcGOujn/
LS4UCLiVeD/8H/O5FxLsLbU/IPCnjx2PODX5ORJqJXDgx+Jpfplq5znIZ3NYK6/BNKmSt2zKaOWV
SIX0bwLOUcnYEsntF6VbT1OkphZzvp/kGglyK4WuV6yDUAok4YFpo3g4HoyoR24zIM0YeaboY2fm
cewAf2azukb/3vm6trTMYJNNoIfsijSiXBCmlkQe2A0eXxCch0/5z+6XJ0NEUVf5at5Vp8mYuY5F
7xUfuCyUIcOqvU9EIN38QGpXn5jLAFq0wDZsuIhayHXgD0ANyUZdcasChb1sCqViikHVXrHgdlwS
qwHSr92XphfgK7Dfm9Ef9un34wYcBb9wQ1jymq9mEeXuhwgxjUhogglAFYQ0OlJ/IzKfAn7GSO2v
ENbasce4azCyapmpOc7om2Gc2OqhwFi6UG8SQHjYjDrZOo3XlYo/QQutsN0i40rxFmJqmhQrqkfp
u+6VAhS7AxaEXiO/s5qXky3y/kFoV+tv7mUL+DwrbVDaC3RaDnblTMm37jDMfjmf+0nck+xj08XR
mave9dIkwos+vDlfsFL44tcNuh4UwwDe9luW5WFFIptIC2U50qIVr1J6lisyYBtOYZIue+cJFQCc
9mk04VoKpl1U3DIbBWr8reAc+0PAAPCVccecAvIeSDWo8uEfZq5DQIQEsrea5O8jA3139Vy6tkna
kvLPzL21HD1B0xZOeft9E2/+NdtvN3aONebS8X8Wpz/WclyL6st9GJh9BGCvXIa8QGCqc86kECVa
VCQpKhJXSk1uLBCN4SXC+cVL+4vLXhMNXG/vb/tm1EKIkK+y8c0nOQm7wfguWnwtHHuPZFgsHPr2
kayGoOv2iTfoW1eZJxBy83xipcpB4Ty1BlsLJ3qRQHGuOyi/teXVK3kP9b06fBBDH8Nsiqpgwshq
dy9xBjWqpvNQVVG/Mchp+iXmVohjbaSwx8gGqE5/mmAUKjPkfEysi3muoTGC43V/pCNhtQEhdgvg
7QnFUQxB49H2VHssKxCFSMqFLLE3CwSdjDxpfGX3/EUcMTEeCY+i75xuHWKaPc7zl8Y4DzPD5le9
oo3mm0ugn3dJ9W2FR6Slw6KEJY2sVfb0QOHHG2lf5LeJ24RKAVGnFF7EBBiB6dR1WMNMr/6o7kp8
9yYk66r9ogkItVm+PqRKbr0YrrpQuDWcGBZCMyTVolOQkLmGnQEET0z/iVg2cFnt/GRnMaKyDm4d
cIJG1fI1nv/hCQPWyxtYr2eNbf05MtrQK7o9sctTk66B28J0F8isQc9ufhMAzYIzD1LcGlNZ02t2
xdSO8LEodGg1VDTfbt++Om1A2J0b1w8Q4Ecr9+bWxnEYMv+s85MPPVV0zR1gYWCzRN9BoJ/TBNLt
1VikJzhb04RUaDTdC3VzLTBoY9pnhrf+0aA8vdSJvfx1upNpBdDbwuEJMiAKGHfnNxjiDgnyJh3Z
4EfXV9l32exwYSCFgHdcAjDAwVLJ5C80gUmxKsTRGGgoUHnVVcFgAFx67ZbPlPvskROfVM/t6zop
4RAJorRfEB+emof7M+pUalSdRAWDR69KzcUwl+KBPt5pOJeFBw0P3HhWPmAj3BMFuxC6i39LRdWq
Uf2dMUgUk4pQ1koeUsDiJj4JTFbJenG/0HpzXT1KlYLaTdmdpiKiBF7hIIIQC9UJJW2Lw/ugQ+r5
uexQ9efqxssaKZTfhioSJJ5aUZzZWNq2YTFPFsW/9VnivP+tMm0VYUqmMMEIA/KAndy6UjGFH3/C
NJavcMeB2a1Rv1U+JZD5KPYwjM8wIXgNnqeRiamf/Qkn3nwu4TfLCmy30DRGJAi4mOMMYIyCo8V1
wbFyXvHtPcgYthCYu+Cl0x3JZP3aOG3fbd8rx4km6GttSgr0JcCkS+ranUvL0WUXBVFMDm0Gn65m
3x432GQpfnG9JOZBEOPVIBbqgv6wJlmUUfiUXRPGhBSsAEHj95yllnnjaHhypaEqunKENJ8jHfHj
+0TmMouXvTq8jGfU605OLi2lyjk2KlWR1RhKthHiFcfvCKPjv6+RxiFCQqdrvkjXjEAaiJoHJG8p
+QA/aZMtcnsl4lPbPTZAcU+gRSQz+vxZVl3/52QSh6/YWxdgiL08mjieRYs6bJX87lwiZfEY84NP
saL/UbdKXueIzTbRKVDEVl1I8GjZj+gTM1hPcqg5MM2IrfwnsoZPcpAKTPWL4uBOund8xHKYYuFF
WUtLjKBAJ/ln1HPQkXLVMNif30y6pVpRQCqstoQDdUReUJU6RSgSIpFfwbb98a0l1P8WLJeiMIll
F0XSoMHtnz5vFFAHOap25SiONHa5XaWSBx8pE/ZPgOT5Ig7Fgz0237DOY3TuDcCHGThj7U+k6dQ5
5rCzY3RtQvyLaPBcDQLl1o3kYFg1nLVd7XKRs8MrZvO0Gw3Wa0QcXmkyAPosot6cV3egY4XuovvD
po5m5VfYohSsCTBqZo7SJ1dxB7wXhVVRwdSK7yPvXpwmupot5uwypjiyG4Tpj+NDF7CnX5Y4cF6J
NLa7vfYyKulYgq0d0md1wUsf9wBK2pXPE2nS64nQaI++wh2Xu3BboJkE5Y1NM6EPUrEy8pXuWb7X
1+YLp92EaEZPlx1Pk6FaRFk020VUXDsmzC/6i7g3plSOn6+b/Xb36LfONuZ+dHWQnpUNQBaT1wkJ
pQyLA4On51cttpBl+r3843p5bdZuVybnrGbq5StstkqOgIepxTAKgtX+LiCRnqZR7PCBoWu7vG7y
q6AwAKQNjO2+DhHw4eekNFLfzfgEJkFFVfxxy9I0iCI6ZTE8NCJS7gsvUyFa1IHtPzdupzYgSpd3
V1Up+/33coxEPGyNmU8HqTnQHPrXoIEXIbMrNEGaQQuttqUq9ONj00QdF0wMecBvWohuToeJgsvZ
QHXiFrA7ZIR1bWpoLsQB+3RSV6Dd7Qa0fOIA+3klocLnAuPbwXT9I9Xl0MyH5jh0Ev3rqbu7fLwv
Sp4544HvrEBs2W0AkbY1d1/ycWPQQos3dO0s5SMAA1H/Fg30PIe874U+o5GiJBSG5YC3IwP3O1Pv
98A9tFYrUz0gM9kZzsopzCPJ9udbS9kAiQjxfLA9PjPa1gXG+nF7F4tZghDSJWSHZ+TBmyZ/flkn
5EzTXFZOyTzrDFvgMp2ctOtxmhrG0r2dWSSCF9Cx2nasaUwMHwtDXLY0sCE7quxmeKeSgjdJs1mh
GKg7Oh1QrUf26MieAp2tCBxOyESamsDWFjlQYPaVaLwauLLBYWt4yeXQ4VPdgvWZDTuOfuXk1Jgz
QLICSt0RURsweRaYrza+LJpbvtNWWbGxBCJsT9+MCkpB7Pn/uwT4tedzxezDIlqEHipMJAdUlbPZ
ds0NevVQMa+4tLBsnFYI2wOf7dDFmiArFYa9hTAXVfvTJyE4FLhEt2FJmtG/TcFYxuc4lC+0L0rV
q/lu1zJ6Bed+0LDoHHiRzrFPl8j0pdYYcI4MQDQv6kufg4ml3oCEI5n/5RseJJgutjQU4wkix/Yi
z8oN0GNBYCAs3FDiajMyYAyXeTw1vOSL5PqlKSDPNPIrG71+4zCGo2YX0x6b5+dIoCrZaK3E5VKz
VNtPF/LzAMBOOzZtsXvwFaRJsKF+OsDBijKG4FeHnW9eBBY7nShASje2Imoszt/ZHSGj71LKKVOk
TF4qctNZis0y3qwM6tWcl0g/+6ADuB4rU6KMEO+oV7h5n4YQ3RBQdOvXL+ya4D7ci7P9E2llB9wK
e4kSntepo7SbZSu2wF6bobHVp+Y747Gz3yVOyh7yLFLBE5J0ChPDouc+PWGgShD1tkWZ4t3WSD0Z
jZTlJNd/6r5xnkTunvxoUeW2F7xiIrCbwb7MMdzCz7kCh7hmmhyoX+6GFFwtEQpmwZGgOdslGzO7
1bxD2VxtsBwMyG5MTFL3lY1Izh0fLg0WUx73U8EAMtc7lBx5j+SFlnGcu/ojRKldWpf2S3itHHzW
V68IiJdN8qagBRbMqEGtG2FF+EFnPKh3exvgecAPvWtpOYv2RL6d0U5NHtj4NPWNydK8FhQ1dkW8
TnUWlQ9g0n9SF40oDn9ujudXxqE5D5DiYVLgSBPeLj6MyiuxIRdYy6tJONtQMRaV/5nL29GwcmP6
GRPUIAxg9Tz8gvs9FweN42mNjfJecdIG0SjnkqnmE62odViYXVu38sw2zx6GSB0o+LcPlM4MHt5X
Uk/HObecoQtCAC38Cgy90yzl/bykXbgvrt/oJipX9gHYgfGiIzUPI0Kiach0Jtlv7bnuzEt2VFGo
/Jb4MZmXOSgKGRF3pyEOrDsTMFL+XPgCrkit/ckaN/xUui9ezrtVaYwTT9wiXVhfo2qIuaCJu0Dt
um0Yw27DlW1MPb0wR7DYF8C/ufaaPkcdEtf6Hkeegic6CdLwpTnfeuVkWzYmGqhk5cb7vAxhAXod
lfpaWMj3GhY2rZxB6cSdhpBHufarpLgSS9C+SKL1XV1q4oFGczNOCS7qONPQsMBKl+wKk948Lr16
K4dvDpQGDVqfbBJ9WLr3TvcO0GU0KFy5ORsg5CR7/qJDw3+N7cXWyQmXCScC6JvzvnwrMkqg19rN
/TELFpJwSxpPeaF5JxG/8EnYxzsmLrpa4MCcBJBNjFmyJUm+T2g+UOAiqKtEQzjWZzrqhpFtht6b
Hy4TgKlzfZuhBrx8z4OkedVmW82uAL33wzqP7Smkfg+Yl2myYqoqHSpgE4dss5prcBFOouWBqbG6
kPCasp1hLkj699knsw6w7Qy44Gn6R7Cv1SXoNfbJykfGC35FqxPQhweL03pPe/ygUHPLwAbh2Op1
gVEo0/9TydoVEaPbYHsHWuSWJCRMFxs34Iw3Sh0mwtNEJt4Hbo1Lq6wUo9tN3y05iE1+FGcx7kqc
AY1iLGAg23t9VaDxA+SmuGkT4MQ6V5IaTIwu1s8OQhbW2kIWh5enL9QgeVMaYtoh0tCyeoq02+if
0uWtFZUtPvaibNMsReMVCNHHJg3EAtWLxdSDpv+2xiyhx3o49OscKaf+/957rtqi6So/J6sKLh+l
Pemohj8ZmIZ8GEPoaFeCkJqUqiT0Xss0xzNqEKx+52u7R3PJ9sTSd8/4QoI+OzJNFhhGjD2AmID7
JpNkxZHR6xeQbBtzCm26j7vM1XvAP7jaw4LfEhgYw3+NupGjtnJNp+Tp18tlt0fVYcTUADcJUTri
rQDlF1e9ElMnUlOcerk8qQJ9t8HFGbcL6aVchuKm4RiUvUdcO5rQKtQU6dklbvazufwaCyNvmCh6
vzhkmIWHkowhTTO2lm6QCgWMweUcLxHjaxEfuyebDI07RkwWyw/C8DXFKMZKYZWv7HEBWhn+9FGx
pGeht/x5QAqwyhE0eH69BnYALaMOjsJ+Tc+RLQx9VERX24jNJMpBBhQymQnmB2KCRYvl6Zllgkci
uSWDCxE49T02SEUBoYQL6DCtt3GjupTzW0kdf0eDsCyOn6iM7ZWH6AFF/tf5RSPlQ62mx3I7AFMM
xM9EYrwnrsRkcvxaKXoixIWR2Mh1un7GN7sKL0J1v0J9ZnlwhxmdzSvZrdvIePp3ZYPKIciMFydk
FTrGv2beXFoU8VG4J85aIdGocOyWXgu1AGOflTvEgcUqmQtWnP7aaTj6GkJ3TPLxwyFb9mlTIhS+
6XSOpxutqtiZyVJnFNKga6pCH/e8p5QhcvVltT7Ba/KVI7Jk31jDCVGZZYVUsPnIjJUcJtGhbfAE
L2Z8Xhhh01xgGAsFb8vKK3mTVaYkJuUKxOxTlugSgh2LKazpI4MPwn9RNzB8vdR5dxJrt4RTS7hF
sFG4BKjGqsjrhu5PRmRFbmrevqBlF84aMFeiyVmuBuLUpD+DicIKl+KncLIhzjHYLrKLRMX6T5IF
wD38/QmcTUjxLY9E1HAFgARaN04PHQzLHkBH2r8yMjCiFpZxILWIGVe9M/3cZvetOH5Ns0/rD6lO
7OXmA0TXqCaKOtc351U9snxOIDZOQyXxZVUkxtHO0j13v4Qf76NNWcSaQjxQABakS45F0+kICpRU
w/vW4JcykKfn8VWpII7iz5sulRjH/YtFe7ohc7frx87UF8m04oC69b+kL2KZ0i0zZed3De6aqJhv
xxX0ujlq4lpPgJwhLJ5N/xrBXfJpPLMsJ4TRRJI3DWIHZPP1n4pzxVj/k1v+53KrJwlg7NKwUUeH
4tU0npp+5Fgjh9igkZPl682cKOpnMCDOo9Bp6dtY1ht5TVOkmZRRuMpHuF/mAaxJMHK35lIIcAE+
cbm4OiA8Gnr8xXwP/G4/v9rnmNl41Itky6k8cBr5aYv9gEfZaHmpN1bW4mCh47UNR58ET5yuxI/x
FVh5Y+sJdchPmzYPbBebFH45+A4YiwSmpaHoE1Vh7G3NtjnzMK04upLNrNAH30ka2hfjO4P5C9RD
yLE2F9vwlNiMU81VXOQ1mbKorqIyRCRhCkaiPvVkKEP2uac7Ub6188NiGWWnJH7x4FUedWQsqwPI
2ZVB/uf9L08voi0Ahd8o40T5xlQsJ371iPF2LtUeo7JfUDsqJHd31V32b0GOHW7UZ78p2BLvyQ6X
OwVglMF3S2EorPp/ZaDm2B7Sz0PBKamjICwK3D0j8eSrJ7LnnSO2D4QS62IXiNi0cY0M12g6p9hf
Y8Fa228zcV/ODzTPTpKRqu6cTund/AVFi4uzyUUuP1IecrLDnolyUY3mXx6HaVcH8TP7tYp7KX8s
SFQIJmWAGk2gdmdgRrV+MYbc6FY8KHnFOj1H1SkoolP/7eHy1eqZEV4GB16JN18AEhpkmBqPe5bg
vMKEq0o7gBy+VU1ewYQo5frfx8lzjCChttCFQrF83GsS3bZUTkIj+5z8EzyVc1hkNbKstTgbZYvG
MtwSp9CqnGWkf4Ib4QtF+ctKyj5EHCHJgNZXq5S5PIK/Qi8DIAEO72eRigT2iKeKz4yWdq1f6TSe
ieZFurFxJjPfcwiTBpyVgUDNguMfSzrD3GIprs+RE3XjPxHyUyBn7U0xL7C6rSsLL0jdU8dqyMyF
06lnpqbXy2j4w0tLsUC2rybT0V1OG3jv0eRwZP3/9NS/NwAyPCjRQz1rgO8iSaf5wnuIDKOISUJE
V6E6aBtD0qk/kDzPNzKJM4Ygo6WKZ6LX9DT59DZcyRqze48zJLuHdeTUa5eJUlqMqB5iF6hCbubP
OSmYhD8baPLGJirxVynad8qMHgbTDKgwpSAseL41cjS7n0E+up2OtgBYHAlcyHIPcD0cyJH7paWB
io/FJJzuhwLI8/nFmJxF6dsRDIxVzjrOhl/KgSyuapKTdvNUwPr5B7oDCG+FRtcghTrCMn8UxBjT
jwIX7hIANrYWGQ2f0qrZpEzXP5Z3F4fWyxg8W0f5E1YS4AMXPQ62hQpoif8/aIVvBynKQAPcF8hg
uRJZNGskhuhAA/ew58feAKvWnLwLq0VhSSqxGBKTHrTYueAibMa1Ij6EvkdAcBR7rebgiALsteIB
yEClDQoItQAAT8iBv2AUhRWemLRvAEuz9L/GNQnk/Vx7oFm6ylnvhsvHbsvVzurHM/3C9kaMDQly
KlDayyfYQ0nWkeKRhstCZkmxC32p1DQQ/LVBiuiTh4Jn+1Jja1MC0uQvaEkKCrYDmNyKbioRdPwr
jcMHTLi+nGEap2oyDaIKpiIBIj25GUVs3zar7Aarf9TezL7ac/OhWNRrdl3gZvIg5T4I2+8dMuxI
d778K/IsGBdC5deaq5Zrl7NZ83MTFfHU7n73T5nrXRyctp06Z3QDUCjisqpag7q7RtCuBFekiSrI
qgXL3/ttlcE4ZwaUNMpmaCAAVdy9psyaj7KP/vOUyh2QTlRyIieljUeiCOIq1VtW/Xeiaa39FXmY
0XrCrkhZTAJU1bbg1hH1XI3uGgQCn0kkGFruuadFcDGE8vHPJXJXQHxAaWk238gqRG9UDYirD48P
Tg8r1vXwyYb1Ej/DlAAQCoFIfwFymeeeTKqCBaXFpZxGAiZiPe+HLn1MP4rkr5D4+ZHTBsCyp6Pg
RCGHbyaH1ZYcXOtPJzKj6v0NtSV3/Dt2H/ewGJuBeQJSoCHIddYNQfEEh3glMjZ+YZ6QqPl3dMmd
eaJITzrZX71TAOqLZanBvDn6PaqoOXXP8beH+C0sRqQkIS4QhxYrduxInUstuw0r5iaBo+WqgJtS
TAXRjMJAQnQF0H3G8ABbNY2b2nfVIc7Jfa3ukasyYb5ZXnJrPaMllUquSFUuOSsrSU0duyvPnmVO
hhHwyEVjx8I7Y/7IOIV7TAlg7WA3PH7xzGKcWNAWl67Dup4vaf96515o8LvZ4LuaEByfKTccKRuP
WE8hH277MCz0C740XAyzOsJtc/+DOAt00rTBXFNz5YuPOWxjAwcOoU7qV0mdrCxy1JmiTF7mb3eq
Sx1RjiuETJBX7YbTfkOJqRnSvjbQzOAFhug5kbntJnzvFYSHzgHyVKIDVRF5cA4NCrijgak/1Xmg
REq0AxMefAtP/wkqx85eiDMuK7oc+NG5PMJBk7+JB88YA7A4JNZsgvEwX2oHUsABXQ5pLexWB4yC
TiVcEJ7X2Jr0QHcmYjRajhW9VNe97HlKJLR7cWGaUsi28Ck/Zev7JD2Tg5wGLy+gTUzG3Zf4LvBs
bSr65lMPrihguqKkJb1kkAgFaO2eTLN6aro9j109Wc67N4JBkotL08+GrcPc1TrY68dHhK0hzZTI
wls10ZkyGlOAibpP9yDNU/e/QLRzOnMMfuwsoK/bBkwUlYk7WqlRiqQXbrvJBCd1SiqEZKy7ChDH
WX6S4WuGWGxtnWSozDaBc/J7QUtJERlm6FJfMK39zqSD+twunlMLCoxyCCY4n7+5kY7J7nTkSUWF
7BKwYfMRJOBeRgjBQh4V2XcYGr8K/td3djDykwz7lKfDgG4wL+lQr1e/NxDBoV2g0IKbfYPTs2Fz
Jnp2nvCv/1hS3zJEVjHXkvY1qJS+OIpNXILXcC9yUecCmE22wsmc+nianBb6/GLdd3+RQH7ZIHHK
BVzYgYXLsqSOVoSsRdIXmcF5lsXRzgIGLnAuQzfyUrohHrbzXiYbWvnfuusYn/N13Y7nqANyz72s
nv68B8KtnQPgWvI2NCZfl8u9lgwjagwmeZu3bhItkQdnZaTl6k/bVWlP1SJmUH7GN67lQJNEoa8c
l2UAAKK+A6mYPWp9QU/+UjTXmisckXhFHG/TYhlT/PH7Im/Po61pOS9/ec1a6GTHO5sRxSEALV2n
gCnDPsTCnzisOsKHxffC+1vVTv9GlytdhG7U2kR21aGfdV9Np6e3xw06sYM3EGaB/h3riG0u/5Eo
CUc7S3xb1gJL7BPlYTJ9+2tgF+bCugDTTSzAvodBUiGWHBDMrQqgrEGPwdDeBQ8uEBf+TTkQFgnU
tW8LjpWvr2425+dPPkZ0TBn01SLaGWghRM5rBVB4PzdLYmPR2587ME5LTSvaCTFEm+mFND3Drp/8
pWClhwm6Vh/yZubsgq86ZJ/SQYAz5jeV3926pb8qrzQD85FTF8SI21vQWFU5SwGrzMDRzMDu6RMm
7irWTRXsz623ChJ58mAEp/nxMUNi4cSjDuv8iAndl/ayuy8G2ukAMaeQD1C2UkEzLP2fHLbGnf/a
wMYVUinobcrSQ7CGJ4+g+n/x1lTlDI2YfcTsUMox/vAaMo/MNv7OiozlLTgbhD3qSNUrV9gVsUHC
4w/3c+BOErsqyhwjQe8jnhAFS29P+6D4HO+tSKTt4h26b4tZAxIYn4gIYMGwGCvYcnXyNMNJ4oWe
4riQr1hk4JdH9/5frgKUuOK+03SebyEhQLBLY5uZeC6sStDkHTTiatRANrn9MxaJ3A71xlNlqH4s
yU+1iNKf7NWbN307btAFkfT0OKWVCc/zJ7PBiDSRmVooUOoBZ+Z8wIcbSFeOGgEs6aA1mP4Ga4Dh
74XKaSAow0iVXnB5xplPyN4wCFgUknHBzZQ2PIY5aM59lNtD57nbZPdpvRmowdn/dhdHef8endjU
tykpwoc7MOoeIkhUZQhuds0mdIRlXPxkKm9ETYPikdet2RKp+KExrR6ee2V5c9y2YJoL1twW3WPw
6XcsN+Q8qQTscPNXh1XKaw+k/Fo84qURotcVDWqAy0pkI8lZCFO2uC/69N8BNKwJ2lfKK7Es9O/Y
ekVppekWpeNgy6QodhatkB4PAQMsZAWbID8aZgmE/u7Zi/WalGSyBCdAfzkB2ZMSY/Zj7WT3Sn2s
4ByXDNvAOD/r5KnCpOGp4Kb/79QVZeOKtTGeTs0eeehCvc9jqjcXCL1og+W7TFXECKdCd6vx5V7k
8ZpK+u6UOf2/OpscG0Ic2k9amaMqOW7Mx0p7jvvJBc4U9xzOk6ggBI4/9xUwkcT2w9N7fDFUgM2N
y+aboHL84uhkqmX7jrSjD5heJ7m7qFms0PoXq8wpgqbMnfcg2Lhrr1iM13T7tPFbb0xLMrxUU023
IRGx+01i3oKIrEAjV+1GT1lMFAjvGEJ4mWjkMq+w5oWL3YKc0bUDuEz8O+umHbAFM/ecx2PgDBAS
hVXA9abD3KfbbrvKo7x28ZlO/T5mJv1GOhvqYkfEnbNtpPCDquGKSuJWop+uSu7NcqRKo2znb5aP
e/P11DKPvs5fZS+3WVg545NPXABKWdwSP/+5SsH0YHPOt35zxEYFM8uBbyURiG9Ii2WsGOf7QPyf
Tvw6iSdzMC1ZroJ1RYLnQFLWVGaUNF1y+AImPrE/KGYHaPcOUWIRc3Xp9m1vDDLO31UJU58cyoJn
ZXoR2DVl5Tp06deZBT4hlXf753LwNqI0cu7TYovuXnMLieryFStkIjUhCfsCNG7vzdYzWwSGtTfm
cYALKiM4nmdWGZL4YKxKILeOZH/ixA6q6Qm8RGuVIQWMJTZhs8NqKHfB3vb/V6jIxn5CDbXVZht2
c2jXPlgo+sqyJKy2NUV+xnT+MoYf3H/PgqR64qaRMA6WfNDTlLzLNSNYUHU/dehsusjvAj0OZfjI
tEif2R0hW086pVV18KK1PBJquhDRgYiLkXyYX31xK0IAZneDleSxI6sYn3ezzGdd5sp+UF5zYHbV
OvVmoHNkVvDxY324rbzsMMEZ2+/W4Hvg+pG8SZLblXnVYebSc+dbJSA463q3i2qkTIjN8o+tDLIw
6FO48Oaxlgq/mvisUVucIjtRD5K2puCCUItrWxm0IRpYBthGkgtAJ1DQjA6PGehnDRAijXVCZj5q
LGI719tpsf5rEbMJ9YjPIxR4e542suU4kV09Xp85leb0RFsjjjg3Swr82GV5gARH2VYOzSRBITm5
pK8ETMpO+4+5B+yc/rZLLrtB9xvgO+Zf1xc9Ymwt7C7VzeRaSQlIHgNbdNlF+mhg+NFDDYIXXPYF
UdHx9B0XoIBpZS6X4EGvtiHIBLJWxj6l56RE295uBkqAfOlzZ3kQ2HQMzzuNhVzdyoLZ/s+hqHTA
yggQqAqh0xGyslMlnobJjQciu8cBHvf6ccxi0GS9BStl3Mh9xgmsgc65qfV8xPgie8zPER9FoXxM
z7JtD7QKHmbQgwIpdtjPLSc5iUneIUdS8HhULP9bHkD9e0VSQWuLfDzl7FJ0jd4Xec/7vsYzAARm
Z219DGB82RcOqFPAkNtl+FhG433jQ5aUmXdI0XwkFN9RQbB2vzEz9x35udagT30yIHuBYmMFJS/P
aEcnMOc9p3gpY7H3GVvU0HjpIdTXEm+aKlIuzOvA2unAE09j7yHF11FewUmKg+yQhIV/exGN32d6
QRyF7MEkzYFLXOSG+WT4N/7opklKUM7i9ssH4XUcdwKAhbM1VF0Li2rObMi0tSA1ka6T7r4XxcXy
hpgq+T5dn2Ee2RxTGTh/09nzvIRE1vHbkDcYqqEfIG2f6nvS341HGnnRHmLADrMnk6OHWJfI/7LV
tuTHudH0EV6ynv+g/0XpTVjUWbjiO/1mYg7kyAxeM+OCJFhjLiBBIUhH3kTPGip6IIViv9oDq0bs
fchRJ6L9fA7QhVgfJddE4fD43/IUZBOR/z99TuWDdsGJx3eG8B4di6F3z4bsy+l/ViVPDFy7R96O
U8HjwL/iy63Tx9KRqaef8dGzc3bKDbZ/yCJXg0THLusPEJHJxTiNK6C6GJt+K/T7Wpy/uROIExRg
ZXrGXTIzZ5/Ywk3eFxEsgScOdQw0i/PPsYMr0jzFt6N+ztlbexQ9sykEdvEM7LEfRLwUdnOCtsj7
JV6py26A61TOpZXhjKaNjNDVJgHytHnmrr1xt89o5mzhtkwx2azdwqgNQ3Nl/lnaLXi+zxTFEyZT
TU3NI+wAQWlgoNVzwYH4cb0avO41Ms2xiSsqBSXyJVXJ9nLfNWltZda2sgJe2jCzl74DELdDzil4
GKWe6PpUnvWkdoh6+Fug22/P+JUP8zgPjOBjZpWL9qHiQM4A/GhXsrAVw9wfmPmwvflz527YLbtJ
HVtPoNytqc3lTqApWB27p+4RprNaZMbD2VglDxaNZg0u4yuYYBbKnJNzkndSQVhemzou19gBWeil
b34HHF2YlpNfvh9zhBkC2iUxzC1vUWC4/ZmcTpPvoc/KGPaUVjvXuGJNERl9ui9STFlVeEG/zn8n
Pzen2EG68N9JtCgMq3x1tbOh1LfuTUJ7vC8YfZXnigWIRx9lhOCfW/rEHeIr+ryWkogD6ddlWuJb
kctI14tTvzTk0XhU+SspQP1l2jtMio10F1KJsPJGJOpFaJA5Xskaogyx9hTcDd6J3HKzwZXUooAP
+OhLPIJ3OQJ4z1k+cJTEBgBMu7rjStxwYZfiwwfdhqu9ztP38EWLVa4JG/NcXZazu5biCBc9DkBY
iCKoU6nRIRD2fEcvo8c7UDZbKmfPuBV/KHOtR/tU2VXHvxFe5EW0jVdjeeMxWabulKgJXVisx0is
kosazjSrdBmwojs/fL2/e/GVaqvo58eDBpc0ciTzrWdOtI4oYd5oHZViaJyl4MNHe+OIuSTR1dp1
2SQXNBIR/CX8XtmErQIiAzbvli+0PMoZLITqDNZ5VPCGprNXGChwipA6Q6e8f7CkVpij/VWD7nJQ
EgnoKglaPGUPKddWgrkqvi7gzxhMiRMmTR3A6IZ/PSOJV0QBPE5QZDGYxkl+n2+oq+Kc2xkVsi1p
yJLRnKZ80gUHp2bhr8ClJRyMM4SW6KuxlDXfCRwWEZMHVl5h6XMaOCy9buEmENaUMGzYEaHoQs2c
h8XN3R/9Cd6JV+agbXoZce0nspnOaf84bWj8pxhpbrvR82VumA2iqUd/uR9r21tHTyh+2HpVHL5/
Sc97NTEa2O/0n8qVLzX+ZxlilGzFcbaoNs71BzyZwWulnL6BRVCANynHZBIFM6+XpXoC/l7LfORn
bDJziRLn7HPrrqMF3DBmbvgGc4UXa8yj316BoU0d07LfxL/AZSDp1MlAMNqLKR9toOc2ffnTUqdn
sVd0tcf7gpeULtQthMQa5Cqrok9cqHN86ojT59IN4HHWDhjrP23prWRyHm0HITVrpmMrqTc+muIC
yToNnGeb7sPk33SO805smj9KBhYMBiWJm9jwCmsLjDoAV304UjgfaEFkAIxdRIP6+ULfVi10Sa3h
nncI22cTfj8W/vzP3UOlWiRM+nEb3p87fFdyuAOvzSNIraOkBScG7+t6Wv+QXBQ3Un3BsMcZR+m7
ujksJxHkHeAsVYfWLWdjjEcK7NTXMfvXi6IJzxRp7lxvEvpqZgiw/1v5p4cq5gWK5yaT0pXFAV57
muBcdKJMtzTl4WtFWB5B+VPkRWM1U9IbYIBFUe7DOq9wMJajZwaIeqyPoBpTrfuYUVeeJbK/hKL5
8DMnS8BVER/yjTWn/gzjWR3mviaOMCQXd0E4mnhMAuFkPvT+5DydYV6kY5EFgwXOy+i/IO9sibj1
puKqyTiJZSCsZIe2AZhl19Hb5fMPzOK6xNuwz6quoGARpkTQda4tuvk6iVCpiq5GCCXXz5vpS7Gt
0TkEgBmeWkfCjohpezXp8c2hl3vuy9OMnTB0e3+14BfwsF74KZWfx6OyAzlnnrrIgaLmx1RetgwL
NOO4VskY9VP7ESfxNm/9k49Wwq57TJmenH7VSD19y5ypwf1KyjD222VQRdgAeLLOq5y5Ef6Q6f1g
UisLacMU6jkmE3VRwD1dKGB0XnIQifVgYDgjbuJ1neDPdxDyaVv0BleN32QpCLil/1XJPQokXvNO
yT/3qaiSG0PkS7il1mTKcjz9nOjNJ8/V7QQDLJbz754ZPh2WlWVFsXPo20kW1UDMKCkVdF6yafvd
pWQWNmr1TFMRjiiI6B5l50l1jhFKVtYkJ/xXTmtlDjrwktDdH1miZ2d5pYajUQHVMd+2oVRDOIgB
AFptYRvJlDinY84bZef0MyVGqvnAn7dTPZ6Q0E+U8LzYhKeOP9vQVAuD+Q0o2m3/d9/nuxQaexNw
AfzNrbFXfxNq1Ks9ARm39JnrD0NDSl/3OtArYmy/oRS12XDz3PDpBQsbPIaWVH0yccgEPBygWCGC
dvWCdqDs0C1bshEQ5+Jxkxv5mPET4GfkaKRJPcx45dlMMg24t+LZ4PvhtNIjCN4dhUU5Bm/dKLpd
sZFVOmJu+f0Hbl7BDsm5C8nbbLcXSc9OpI6Vua+rTuZAYfUYm+hVzlE9MbogDz/2hSL1MlmnFJyg
0KjCBaX9F0afD2oTLIM/8KtGx/7zPOEMbAm06Y4SssrS6stIYHAFacGAZR9lQaVzWo40T2UNdiT4
ZQRtHJnVz0NkNS+JwLRwOwfzI5rm0pCpzi/STqunrnszQieaw7IaQTGnupKDNrgRVQ6Q9uVzD528
8zcXGa2EbPirKBuW7LE61ZZcZiDQy2RHA9vjqn9exV0o84j4UnzqedI+WytVuYsDttwyTXeXJ3eS
0K1Muric7328204hTJST6jxPnbW6wRpXz9f1dcenqzoav4TQNn67BaqE2iF1J7V+NGnM+7JbCPgy
wVlPWP9PBsutGl1ewDdW3Z0hoR/IU5Fy0/LDLSMJRFHbBUj3nOOgD2eVJACDTKShlGdFfzktcgeE
loUQYroif0UyXM0IKEx+lRCk2MCz/IdfY3NloSNVkcP0jxVg21Ay7Syk8KkeM+hHJruuo2bua3r/
mSo/uajCLzy026xY1mzXAapqGpA245B7/WebQ1k1RViFI6acgOhHdcUAuiuOvhX+t4By55NhybG7
sq9GTCx5yVNopKSFF5PPTgm1UazU5kQv30jCQjogvxJFEMZN7PWooOGd2DWV1DxlRh5elz7f8Ann
Rb9HpFHwxJero8t2UfJaDpfT8CZlCGhEsx3qHVDh+pRvlPz6FsyZd4plp1OjzLHldMkUS2rw+k8x
sHmZCulceJO3a6YN0fnNFFNZrEwLS0iodBf7nVi1jQVRr7obky9lfT/ZLHtC26Q/k3VZDhvVrre2
wMOo+Yt5MU5DWz/Z21TzGf8Twqq4k138Va0J5ERdhbRomanNbpstBJO7l7NeBJumSLdRKowWi9uD
hFsuXYFqQleobai1M4a3B/zaOWb3xmVyxHO/C23u3piLdBex7RPZzjxTffr89q7aSwseWkk2moIC
rluOCQ97MF6GEc9UoEzYsi+0xxTQzB+IVxR9Ip6QnvaFVLpB/jkB8M6cSq+zhuv6WZTqKl63QlcP
5RDy9wdQLoJCRTD2jJemqFX/JK9FlxQ+ylm8g/nKS8gavnh5N/hNUXyIjc9M/zBjKv98Ec1yyzJU
aiIfY8zI7hWqtys5zRwCLxAf21y9c1G8SCYUXO4RFcyQRdLujK0pi2ha9zLreDUVVEpPzUT1oluX
+rm6pDG0KJin2yQWQNzhrpmLkv61uQXFGYYiJXtxJEasrEoJGLt/rRpEtzOJOmhaphf+WnCZ/z3a
9AQ+FCF75NbUiWXGC3SNbydegEVcc57vagh9ioYyl9YMhPlmolo5OsATtFq54X7R+eKZvlPVrX4Z
2/nYQeCmFcDG3cFS9777fSv7q7Z8VBXhm4+cKwQnYQvnM0syODb9b3MiiRGgIAZU9TIAi21dAJw7
XdpwbVIEhFLqKvMHheQXIoTZdNTkDm2h8pgFhy8X5085pA72kDEOK3YicqthQy8o9T4OmzpIM8er
wd6BWqDz6yY11VfMrqsqDasgW5AtH1UlaPsphd83OxrfWbDR2QbMBvbFXB259b8DdB8el5fnR4TE
paaOfR0OZvqM/bY21RYCZvnRwD030DmW21CAnz6F6Xy/+Lzoyv1GidDK7g0rGPJvvDaie9bFGjyF
4wkpk38csK7u5r5fOyyUykmSG77OoC0jE/Ap1gueFhufxx12zl3u1NCaTtUkLjJO27n+3t/FFx6t
mETMBEBP600zqumYvGYL66N1fvWJTqaUrPKxFqyGubtnoIUeRFQwFP7b8UDjcwm8C1DqY3tvh382
17hZDuvHgCLbeKBhYCN5Ozq69SgX6ReUPMazyVjIDk0VSbgNvIN9e+8t4cbSZlRFA/u005XwLVRd
gKpnJB6DTZmop0I2Xo2eW2Ia48RtNpQn5NhbTxP3KIT1NN/jel48lKkUnk2YSODUPF3B3rtU69ik
C1qScQrAuX0066hb0ksZKVRJ6sPLwUySrOzX4wcTxfLecR686w892dUUDvJ9PALVtQ43se4TN1OB
8cNyfOeILoatjR33STFrYcbP00YpvBCfnrrPbRyRDHYL8zZh08GMpb1ayuvocCkgnmqPqGepbg9n
YXFE6gS9fE0cVsTbXLeHkblF3GFYijdaX1SxsNghObCrlyNiogjHmbQPxfJoUlZtJkYhtTcOxTJX
IRETqC1yGlMMlpQENxl/76Qh+PbRVt9RSR5Hdxi1h8UpktEbM6Lz2RE63+1IYM4ex4/qiuiSgrei
53AIkXeW+Uo3W+YBwoTdYSo65KmeCv+cbHzaAWsQ9es9ObOJ24UBitNQH7IML5VkJvWJP4VBH33Q
UFCcYlK1hrNh557Cyf53fBCYA0SpcjaXcoNmBBlhwH6o4WRWsvs6WUL5Zr3pf/07/11/uXmuW0yv
XH+I9lkFLpN3z8FlCsVgqOTLDOGuEf/qeS7jDZQOoNhbkdObpVCYrT2tEv7+PqadAh5tbNKOOTix
GcBRbnhNZ90kJUXj88AxtZ1jEDILBzNi2shJSh1oIgJCkemlKux+9ghM+Js2hj56H4F0ntz8qErJ
YJTHq5AL55nep4sPvXdv30jKnHi2M9YjCtMS/s1f3G4xJEgRv6PD0hAqriUR/WGtAvhf5dm8z51A
HhrR1LR3lFgggV63YQdc/OVwv7NtiuV1UWatqoL76NFxlNGS6X73Gfev4LHaKOZTD4B1Cfee2ZLl
AZjsaI4kFxmJr1DwKgiCCheP7stAv3QptH20PhI0OIjqmHnL9P44INLKn77bTNKCZ/sIqZq2/D1d
iZY2QnXt0FrWcElLVGztUIwdaN33sy+glP25yClCLqP+URTgR+YWyH0J5oLMQ1UM9TftUKt6kB0V
6NiD/69kjByzv2n2qbIuO+I1TuAvs17osy7U7FKxYUCcDaMkNpc3bzxiGerdTdi1FPINn/rSR+Si
5Ax1Q/SaDiZv0WKkKaJkWrvpl+jFvOdhPdV7lt8djeY5Xp5iU53aFE7mBWThvOw9hax3hHRAz4MW
FChHkouq8IEsL/KCV5myZnoF8rMrwvtXocm+KeWMYlWwHLrrJbTjXayG5IzXDdbcOQsGODLVYJrp
7a0wkeTNS2B4u/vSoAdQY5CGo1XzpSNdGYx/jgAm/uzlHBnmkhcmmtSvcxY7RiDeu6jqsKqbSBkh
/BL73oviIUybYpanx7yaZAVXA/w3oto/bi2MuO5SqBk3AbbNINnwXg5Hmi6MqMlQcySWPychi+VJ
WN61yCnmyRsFcq45yDnwwClR1AeB2CUk2t4eKR9ke/DtXhlE/6UPQBPKF7p5oa1wPX2HGAFYN0rc
g1czfSn/OBa1nlLftRRFY5wLJLWdg3KubZ8NmzaLR3VvugsMCcvTjuVIHGSKmVrVqGE+IYs1xGBf
pE7TpoizhbkRd4/2nHBG4EApoBmGL9UF2+km63j9HAs3F+MTwT7IVEtmConKmXg90cAX0xF/bXTX
EOr0rEZrwP6lljy92ZSk+mrCi2pyPyg8tCEUa05lNTd3bl2t2RcqICnPT+d5gWqg+ZgGnxpYorIr
+bF7QL2x9E73qpgQrkU9e7qQvylOpC5iu5TnglEwBbf13MY894fuarEDaPsg+qFhra/8jONXfA64
R9aoD9ICRykzhnmsL6QCFc+xRk/fsXtMGTCUQ5IJHlCeazDCSnwisCgedpPuljYzY14dcau7vcZS
y1NFuIZhwBxp+tbLCNRYE1siy+L64FtZ8I4Py9L4lyp/MGUJ7LT7egCK5Fn8jiusSe8JUQmQVqYY
9TVACH5dXsFI2OObPsNn9iBKPiOVC2dJ1pxskZ5d1DceGrCGvdAX6/mdP9PElmMraoXZOBWv5/8C
kIcM/jpnWbDAp6OjgAznarG7yVQws+timboahGRzxjnBHe04GjVxhWRbUK0GtoOLgsNv8A7W53FW
vrh7TMVOK2QQ0TIjJA9+6NaQebpdlKOJD/cLYvISQk+4tZ2o2dr3J0VJNR4TbSyF4NBFwqot1Q5o
ZsLRf3hG6L/bxe+GlTt9PXyJ/fT7LofhsBSuFaAHaBJQ52haImJq1zbXBaHJoQzpGn4HmLbZbNK1
GWHbdqofzrx2m3g+OO9diyc5B5Q+NPmWCOIuohtR4dpeBsVh0n2tdybcJwojNfVv2H+71NsTnDYu
9w6GlJnT4cwLoz7OHvz5T9TkxD/zzS9IFWM0x5Lhvp2HOqToh7X4TO+f98eeHpvijN148R+Wmy+A
9XeGpd4O59rn6bmpHr43g20Q2JD1O0V9mAdbT1C0EbT7Sl6lxaE+dKyBGdbPziZ4PND1HNjLFLJI
get/jK8DcVNzy4OP7VzDvV1L6JQts0DG05FJbCP4CUbIqIENZYj5M3jHb4RZaFWmvP/yrFCB6V6z
MyejQXGKEZWiZpbQ4/stz40p6PU3kzg785K/rmrR5EPBtQhKHmwL9ZZNeKuEVb0CwIow5rb1R3N8
bVkFuI7z1OJVbp0KB0uxUNKz/34P4Qls9Q1mbzFm3UwOX4j5mqDEWKLVnTYyZwDvNNElyCICrO4A
3YczCxaCe5pjQv8V60jvHj2oGapiNzFxpGQMUq5ZMeXjsT/b+BOQ/WD/ODlinw6+u2qafeCGLDbS
IVvC1C+TyzOi8VGr27OTUwxbCbubTcuikwBDd6zzLWvLw91BnPUmOGS8Z8nS9t187tx+73RSSsVb
P9N9IdLH63UAr2M3OstUWcHYhPiHWwe88NtE8WgNZvCXtsbwMap0lHhywVYyTKxHfvm2NTsiDe7m
m3wqZXLG/EEarcUz4O7N3wrwfC5bRmQqscjfcjBOGKYpv3fOCAegbqsuBOylCB89bwv4Z7AgW3D5
nYHsMY2n7uFCMYdgDHxO48WbShH8EP6sWg0+1ra/zYs+QUIKe+GRI1IzCLlQaSbELgHN/8OWV0BR
xdTQp13JeWVMdaJwvnG4C+iMspE+OfWRgH0w2s7bEilxcU5W2c0FBEmLSf4lVkgRD2CE4/g5448h
OgcpwCDIMpN6N75hXvELINCJdtHbHJ9lIKfUktIOVVFcn8tAmhDifYeMSoE4uzSlwDGMT4X4sxBC
PpbZOJoq3m2F+Xvi0gDjQTp95c3GswhO2F96pMcr8p5kkwGacZA1fB6mu5axHKk99bm2lT1ps2Co
X1UYoPVoctasvsldh/If9IQZosKnTxhDYaUXDPv89lY3vBNh8bnliiDgZsYUzJU34ESYLglagege
1Qt6HzPU8G7m8Sdw9emEwScYk+dNwVYQHu+/IzTWsV+k0dyc8i15sECsfl8tTRWDq0AWsMcTfZWk
6T6JhRijpyXZYhs3r59purWYMeP9y2X1Ms0Lr2/3sHjDIp7VRd2NKiHBnGfqzBahlbqExRuQPX69
0OAN7pDVJW/xZLkifDrfUjCtTshbx+PcFsldk1LlHjKJBoamXKWVTeqCkLnAoljtKc4kavnTQG1k
QvLooziM3Onrxf/FOslyFTSGWq5++CUrbDp6flt/4K60GdBDpCCnxSxV2whKNLVd31BAx+iRCLj6
LiZx0p51S497uFYN+q3axibRpMMrWJnj5J38VU4ew9FSn4s2qQIk7FK0v5PCedI0tsojq8VgkYcA
Xj8sVyykJqVw9XgX6ck8ZiaeBbSklYZ1ipWZe1e+Z/Pja8NXagBgVEyw8NWHdIuEys0XHJlEpQwj
KaCStqtXBBozmYh5OQnZsE8SgSiYIjSIJMTQfka58uAjbAZYdea1PT6ItN0V19vxhVbX/z8jMqDX
NEIrYOvl67ZdAlYNUUCMlOxISL+pvofuR0yoAqFhlrc2upwHBlgYUHCelEFZXhmdWZzFY3xFudsY
cxKvG2EShyH3d2uCnS8AWFQA182nVk+1/IOZddXHfG7MOHgPZNrT1sh9YBnb57l2UXVvHFBl95d1
JqvyggBKfjsptGNQheDqlitbRdy3mZD8Tl44KE4Q5A4G9bQm0skUcelwPo8O9nUS/aqQg6MQiMqp
Bhy8VSYga6GPqDSLWAJtc0cp+z2cd/nmkGDP/SOZl5kmFLrba9pxaUABs5p+JlZ1YnfuATXZzLDF
DH/U5rAvb5v4Q4+n0oH6cwTBtyLZZZ5nFA3/S5oGDh7AB2H++VKXGcBK8dk60FRC5zNFt1dr8zDH
4Sd8XuFm1IS5/4mAVLLBfXYQNOFPQymdjHjjC1SZuMqskfMTKMFeJtirfp5lfg2uTc+GIN7Rd2/E
g6V6k+ramd3CqxPq4OHEpe+QUHk3/JCifaw/6yrfKZ1KmW/NEky4rS3RmYmMwJIdO/5+Lcppd2xC
mY5dwg1ZRqC9+T+TmkcD39bmoSvN01ERkpKm28cAHY5r6oczT/Nf9ShtnEwdjemAT6S/OOTQw/ps
EsrVtQOUwA0tX0SdB4u3CXxnuJRFN0Mlu63rRj270deMgos7SG8ibWUpq0Ud8Tq9oAqpS+HaZlrw
nAhlvYi/2fevW4eUT8pQEj59nnzhohjM8q+O2FA+Eguq7Bpizm1UneXJmhMtZ+8Bv1pcYPRbhUsK
ZRwhI+NnWnPmyqlG6VtojKIn6M7wtWzZgEpwEjHxGw2tLLfPm6PD4PqDeWIuftBP2Wx6jUlKIJ/b
6R/sUsGoEkB+JJDf+tb3sc3Mxj7VVZQdg8QBKwYmPk6sySYLbSUYRuauK5MfwE1CyLPwkUAJBzTA
IhorpDIPCuy5wASCI3HiOFXUJtQOdt4pTCB9ssfYECLMr62u3n1yxi1gePDG0wZCFoQnXyaNAR03
+7ZUv5/9s9+hYru8jw1Fm8OXlVmvT6D96VYyPGxhhodUdM82Atg6IMojEjrVGexztdTnT0lWlNNj
Y1jeUja/2zxSLbMVvIS0525oDvyZwkCwVcyVYFvUfs648h+s7/rQ84BAU/46gHuixhPmAnf/Ptj0
ZaaRLhKoucn3Uk8ZdWdJey+5kCQ8Rq8yV/lC1ajq/ZPy8Rek6aSBM6T3qjE1Rcnp8i8rrDNurhFO
F7PEA1xEW5Z+IbQDkp/mtjsYfbmBpeituzTAcDZXE74G+e2bfPeCT5tfK61bQ83hSUE+YNOW+Skg
H/RG9IgGRxvswR6af1o6yvaiFobfkGkkZVI3s92UpwnF5P3GUGuLUkb5qt9nLqN80TCHNtYTL7Ls
s90J8TPykP1u1+QxtJuus5azXKL1fv7zotRwoxrIhixfjVHvbbofmKx346uPKqcmYe4TULH/Afjz
qfZcvRqHcgryNOnJfrwWakSw0wJggjZIcJ1jcqCYrn+wDSpJDwSlVDJP9ftkZ+djvfQi6KUM+ASy
TxUsXpkTCZcg6oNLLqcCIUds37IAWVZAZNL/pJgz/HcdJW8Kolc/Out2jN/4zJD2eolH9LNUQ+af
c00CJdzUEO0HjG8yLMKs7jf90X/rC0wEYFiGjB8zUPdU7suw3n/PI+1Uv/C8+YzP1v59AiQhPZqs
2w+EjJLukwdI+MZSnPTFJD28/1v90s/RBTzzNks9DflAUfgB0GC4vbkkggo92pEpHSCMmQDUXAKn
LVMGRfy1q+s0nsP0eiHqPiBFw+PZQVm6Tx8svwnK7gbltMLHw7vI/metKaoO8abLoIfh7H780+8M
rxZnhN9zXv4zsUwHVo//kb9kwghJ/GkfIbl7qSuqj7qTLJ2UR+zGWAetHG21hNvJDXXJkDy4H0lS
AOBEmGP6Y9nAHgEzkVcJxkW6SVADEgdNIWbaHof8JVZX52gxI6n6Vmv8VdKjZwXEhIiOVXYQ8gZk
k4gz5MEnh+9FAAktWTtKcJLBZNTBtlwFKepYdq4SOXwrqtMGDE/hNHfn/DuGtamsMmYtINR/KPN9
q3/ATg7A+w37G1YalOnSoMIdG44NPVn4gMoKTCGJ9xq5ojWXjz8cdyMTQLWIzofdGztpefNP36eA
h/3iOXClZEfVahHuswYFXNWhy0RQzsmTShNcTrP4obEgbtIqTeW8butT/mbO44b/ocZpoBLHYYZM
VkNuya3n9Xm0LuKRIZaXNSyt1d5BMhPflXJF03XgFcjAzBcNApSBUnX3zXa+iw/eFQsuDbDJsyUD
Kgwej5hRG3eXlJF2d5PFmJQIz9iCm3+v4bkuYi84m4S/Zn85st0X98u9Z8iNY19A56UVSEMXM5uQ
5yfERMtsEr0hUqtOrWf8IIUg+aTzsPsK4q2jWFmRRAjrznZgC2L6vOMpFdZXKjaEsjQu7ovatzhx
XRsgNoJtuDEzzuPbTOLX6rBg9f8McrVRUGHXN6iuM1K2D2p9vy85KXTN0/I58WLskY2kjiY0xcta
Ygki0w8j6iKkK6ei8SCZt59pnN+R7o7mWu/lZH14hoeSQA1TzCsxokvdfbftYC3svighz2P3Ds/D
xjy0ej4ATErs9DL7IJUavjK9d+x3tg3dwcjoAgiySUIC2W0nv2ifPc7WB/7Y6Nwu2OvXghHjcmGr
kYDnzrQZUmog9dSwIG/XVhWo0PsaLlCaMs1p1vkybbJ7vgq/SNEeyBikDUlYd+Eq9IGE7UWJfdMm
3PZST1ZDEr5UVrZEnqIfF/6CU7UVAzih+gBwE9ZLN0n7I3dS7KhmpoiLO4OrmlR+znJ7eho7HBNW
ISafSY6zBlDNn6g9W6IZJG5qTWacO/4YH0Q5w4WB6uVTuYm6bqSn4fniKx3GYPwjIz9oBfD1B2Cb
5GBpGFxi1TFSWC9SmHiLDZ80kHR4dYX9OQ+b+t96ZB5B7qVgsHLLElMTdydHpWQKzlIN5yx7OoCZ
grjlHB4/wV7fOgjwcFfzLBo7A4ApTIBuxc8eIVaxZuXjYzWxCXOclQcDL0i5C5QIyYY9Hss7RxJa
GIl/8WUSnuCq1KtrQ7eZ0vUAYCzoWU7xn/b4WE1sf6AVGCpZOBigJrfsOW0VDZIRc3Iawsc37QbM
LZBg9jL8bDEsfTQHJNnIpqrxaC2roM2pIvnSNb1TwziYLaMVX1J35Q3ftmTuWldt6YJ85Gw0Xw4C
Zy4NGJlo0RVGrtTwYK1z/2zjkKgAvCzcQy0BHspKPbDxw7y722TnVfhExV8NF+Luioc9h7YbtpZ8
B1oDqEBMFGimqCRh4gfBg+JcRNFao40Z5Z7lWhY9KVfPwNb+ELX413CY7GCnumMChLzzDzwROJDV
UyP5dnGajrmU41MJqQOggWmVJdGMFNw28/GxQ4L7AJ3fNBHbU9KaqE+JadEq/ZMmylrLvAMA5Fmt
KBIiIZP9Q+Cwfl5wuHt82SNkeWzBLd/JRsvmka2xXQQqMqG4zmC+GE1zFzLO+zVcIPxZzCFRMTDe
aPrXTrNNY9JOg0GWeJY2GfuIlWd6D3BDVxVomeqGAXJnKGdE/JAginS24WqrHWSNxLa0xOHn6GEp
2Akt5Jm2MbvIo5Vqy4v4/RyaCVXe8HN3k0OcEVJacj7HBo8yIT4SRJ8uJPhE8Y9UGl0QvH4eqf5+
eeGKtx+a5UHgcrVbB7m+OHL5zLvE9njE6SxfkgUGQZzSEO48cbyc4jdtntZYTB8EUtOpdcieXhV4
puX16G06LOCHos0M3S09KiblwYmkQvQJI0XC+WHnQz+SIA7K3w4dguYxVF95/KrTpfR7CqJiH5QQ
X/NrfGUXRAPF1gXoLlv8MZDkMXfkYdZCDrJ8JyxtcT++IiTqaDX5stZJp/9cP+k5uoqIop8ZiL/j
b1gnrlizKfSl9idkb/LsuhkYvfru+OiEH+SlIMkBqbMj/WLjMmYJNZXml8ZL25XA6fFo4B5PkyOG
XMx9IHbx6U7OIohFFq5Eua1S2AV7PVJPkwTCvEJ/4b5DKu5oHNfter/BjIflXnuqCGwhFKEQfGHe
kYbIerkE6lJ5r+Tiku/SOv71HeCVwNYdE2PRMfzlsBrW7nlsneDbIYh07oaVr1Xac8RvnFKWxUg2
h1VqC1Ow7OtM5TPqoFlqRMVCcELLMIkZzvefMcW+eZ0L58/88vrduJ8XCPrdPPdxqJ07eWY8wMrc
CLiGPNxlbWxfVLK491V3B8RaI8WTAkB8U+fLhcqxIp4eGYk+dBqiJp3hxVv51tYMFRBrx8zSDxzz
HKkeLeNM13EnRFlNi9vfr2iJo1uBpkHd7K7uAjzDPjr2Pcq/HicIVb1nujhKBf2lD0UWcKxXRL0N
L7ZpqVOQl1itTgOfSzzcNUFIY2QTUT64nz7CKFXRuP1aoyWdiOTda4r0R2J50pD2/NU0oh/NVjpg
pxmjPk87Il94FNtP7j5feueImCBEvtJgLmJB15qrxbTxUsnGh5/u39RvVBV/teduxjWLHwnCZmiU
39oG9yBYvuzBU3GljFEVCVdB3ChRlpDz1XVa9i7v2uSVz+9d47NFtvF5lZBFNJKLwWhpUsC1GJD6
sTCaW+U4ws9bYOyQ8gdP9YiPs/4kUHaCT/gvVK0D6naVBI2BgV28W2TtoaoaL2G8jfiaNmt2M7ES
CycHqlgPZWcKWH/778byI0kaTPvhkurOV7hQWz4Hki3rR+lwDk7i4buVfrO7ZYUVyrnBfX9PORrK
WMsX5EpH4TwOVATsKJkB9+lGeEODJnpxsqdHiQUDY8xOGyBq0sy2OJ4Q9Ne6VHT6gKwYNC0yl1EY
8aWE15A0uOmNbz8T31qe+JFbyDe2V8D3p7sBkV9GnUq2wOdQiwK1YaC7LeN06GEnGVkVC53Wj+HW
9eZALGpwtJ6DbfOJXQsB9H+4fbS6Dciu1BmsiBBZobOY9FiFEsDldeueJYMtw8HqmyvMNpxBmpt3
RANKtBMr5CiQTpBZPHqvy8OdN/z+MEFgHe0y1SSxMHfinDBxv6A7sHSFcBbUZtO/NelhurRmfC75
f4/LmE6LFxaHvj/QxrtfMTLvCeiOd7NTIMs5ks8JgG6pwpnimacO7R3j4+hcnKhqvElRrSn3zXsd
mcVhHnbUyNcGCaV4rTS6PtytL9XN6Qp6lgBTmt4SnfmN9H9gC76yDIWKEtGy9CyE1ct2iF4Pv4Ff
lsptyKaTUID/8WDQAdHMogiz9xV8bwAg+FDj+yI1t9WJIAZN3lbF7fdZt3+jzObBl/f/Mk0nEO58
9lXFxKERXiiJm0MVwwaAa6HxjaG+/8h/spqGka+ekdDg/nn6mzQslRckHN7Gph47cHtpraG6Xj/M
9ucOt1Bewb/xh0U0qN8PgQ6AbeT+88Ritp8eFCOBRw90tI2ezrNdyHbG8jAF1Hl4xo7t3PG77e0l
Se0TGf3jrD9sEKSU0npH5y+xF+zW0RFt1+C5/NreGC/a0k16QmE50xWEtpGoeb7F+gvX9A6NaQPy
opjmouugAl86+yI+SqXj3CWr+o2KJeHDv5eH6Jfy8rePaYgeLhgrVCXiAvRPnamMrPaIXo+0SJQR
gFAYv+BW8On5Pj1FccY0+c8Tq3uOsUH6+OHmq2Mp2VCWAe0N+9ndIjJCZOjeseIx/NeXcnJckhh6
bmO3fx34vFOnTAjKCxujJBxCY/WoXT8zJQAaWuET9f1pT+IuljWv1G2i5ke56s8eUC3I7S6QaW4H
J6JPqM5lXbp5APUcrzstSURTACeByZsgM33s0YMQP1W+g2YyQ1ryDdhxgFps/vzLti+yZN4kgkIA
aChY2W4ijBcHSXbQ6vmeDm+QANYSe/rJVICZvMvVoWCCahxfV7kLCxXF9OUGb36oe08x0ag4Lujd
YVbAr/EWWp8LO/GDwkB88MR+Y2Kc3XD6ioHZet8wFm66C8Zz5fTV1tZZyfTfRu5BvFbqoLSoLFGo
UM9mhf6Nm90DzMU2eGDf5kSsdl93ct4u6MJ4x7miEnSkLr0sOGZjAz8pCeG4XbB3RwEF/daEjlwc
FpILjMKDJj6yAHEtA4v18jFW1NWk15s1EsqAkJltDHSISXVjEyz3mWaRrs0Abp2qwIsSJvXwEmtd
dTSvPlqGdzvlBSm4cz0wkb2EfPS3XypjZfuSbBAnXF4+sCWWOptBfzOg2Egb+oEwTZMSbIKhRs4E
a9Z1EUOygnJr6b2YE+a9fd3AbvN3t0Z0yqposPPbGgyJhabfJv0IAVs1Cc8Rx5Z6XtLPPGgkMnwM
oUtSByEJwI4xd1GyyQpERYVR4yF2cbHrxlIdwfDMLME+6Ea7k0zOEGMRQ0JiNZv/tKg77iy0lpBm
7+GqvWrxS6CrJ39k0mi51I1JBlVFwoB6uny9TFobbzXmXy7NydqMDlENbphqn2lz+UAnhBdgwhc4
8nlTknD3P1mNsOpx3ot76bqIBUVFpUj73nwRyQUJO3+Fbb2pauCFDpmfrxI8JYQ0Yj4OqpRLxIiH
lP5o/CrMEujraRnccWVnpo+6rHVXAcOHaUdGUac6J6QQaCn2O3RpJh1gar8JzwS4qRnfv3jo4mtP
ly1X4Wr6t6oU/S/y6/UMiPbtUzOvVcUHp8VJsDVtPeBQ02GynCm6IpYSJ8bp8qCvrteBQqS0URoe
Et22w6IsuxhDpGeXM5zpJc1zCtMEwTONDQyDmE4IMJYmRlgxoBpAUghksGemZn7yB6m/AM4RQ0hE
T7Mz1WqvlpRs4BplnoydqpBIe8KrrBLHlWTXGSZ/eBeA6/ZRhltFVMqvZB5deRi3G3CS9G9tSWnT
fqq3KorpNbDCjqKJZOW3/vgj/j2rxJ9ra6j2qW1mrKXYsmortrov6fsJ2Us11DcNdTqVVKL8S75Z
Wskp49mCCQF0b6MtDpzzWzK7TImiLSCRHAhMr+8YOVfZf+DNoR72//PY6usmZN1UZuWfEZOnFtcI
oynDHPBj6tSDrliClmRtk7J0GQJRhCNLHN91Wi/RezD/WRPPx+ot2m3gk4fboOgLk1NvmXRFdI/l
jX25wM9N0nPQIEjOkH5Qyk3ci5WYkP6i/VYUKVtIO0NnKwHplketWRWeX0NIrr0KgI3YrMbh/Z6S
PUTykp2+1nQBKQmHDf3/rrdJAqTK+/wITv2vBj9dYykdNwHCxvh4+ibZDZCw9bBKElU9ijUmJO0h
5VL045v9JRt8w2UuewLRmE38bz4Sgl3KHzFP8nhNsKayUQcbkpVtVFmT3SkffvyYdDBztIdKJNtf
UfwiAX13+fYCdkTwwOE2IJL4RoKv29Li5fO1tdkoRNtSsa2FfnNUrHyw5/reJ7xyQpYgzuG4bjsn
i/26TaviOpzI1+Plf1io8QoXczIwf+D1Akih9wqj/dIi2UbPDSfkgxxT7wxHdH0YiRAxixnlKOGv
Rujgg+JJFTZvrezTpc54RQBlalW1IYA5FYSiRS4Bb2QtfFxC1gAjUfbq2Tyy2nQXVjmCxRUyGDvd
Wv70uTnjq1oTQpnqQcoeMSunHyy0pokELR02VnzDQdrFfnyUtE50OLpRNKlCr1I923Nl7NKV8Ver
95BaijIrkdiAt5XXnw0vcCx3VdIWJqkUuUYe7yABDB0GpF/CgyXYQtD0gkXq4dQa01yKRyXv4uo3
SsdmHIC4gaBj7hj8luAIeDC2KKaJahV408136OgW5s1StLPO8i9uhRj51y9c/yUn8WS6iY3XPVmE
Rual3QnN2WGOrlrW4DRCowuXRaxbOjUfzRxx/DmfcZK3U7oOoUI+2byCyHTJCCZqgi+/CopKMHbQ
bJpHZBTikxODqe3n9SluPmd7oNV/hqLuTAIuGbAt7caBaXhYDwTxP4pFs75xsj1Q2vewOeFtIDbB
a96pZ9xAEi4JmlYzJ7qc9jCaL7NgMoAro+YsHmLYH0/W+T9qBQIqkXH/R5+ruIHgj+mjmMshb6c3
MFEChwDWrOoTkmGGCJ3xUC7TVVJoixXxmCMEI2vAb5WJ4hBQdG9oV5Ozb04rEGFPIN43K4524udO
KrHWumw6kD5XQiSw3YYtenI//E79QUdSPjkXeO2LmPGpuHVgRqldr++Arz/ZE5VPgQpUDS/jnBPR
SyFMF1LqXpY69CZcfQ/Y7I8txIp9yoXQSYQBRO493BSNB9f3RT/flEtTgcFZHgyIsv57TOy9DA8a
Pdm2Ik4iIlXiB3uM6seR0VHB4DvCEFbXM2FnN+9jJJvPDWEYXvixd4p2OhZf1A2lchEH3d2a/tO1
2gus7rXGGLOnwMUAi54iqG/m5GIWFsePI5C1ldVe5iET8qJcjWMOTrPdC/LgScNhNIezLQawN+qC
VUZ8qY9qMthNeyz1L8dFfxxlmklWERGpC48Y61hvhJZElB2wtg+pEvOc7k6ZBRWigQ3ywTWuG84h
dDbSW7e3tih6GfrADsHWSzWB2L+4LdOoMMNOMYuiJ2FAViHjBjY5pdNA0pCZa0OmfOCkHU4RrRoT
7JFm3KIwG/6ikGOHbFR4xC66RD4+tu/tMTdIs+7ZhHRy7L24G0hCfQk7EroO0M7g/EChHffciaAO
TtB7oKtSO+X1/vdKMaSQsOtEPwEGppjsTrFuCcWPVxT5RFb6Bc73NoXTACrz17NrGRVNyU74sTfk
sskHHpx1Kfri+K4TTrajVl35WCnlH1gPTs5LHOG03y0Aa3D+AxpSWOUXcrKh1Ob0Hhk77VHc2hcm
wmH5Xw4g+ZEemhotJMwcG64RsI9NedBcjN9z5ja8OF3Ubcg8Wlxv0QirNUP50L574p1+1opotK5p
tu8qryoZpW9te6E7ObGx/8UEy5uk53UzwDnqDguUW+a93NVWBOLToInNuD/micjsXCp4hdjylDi5
BzM3zigajI/Gf6POw1YH5Q3KsrE/Bd3SF3Y/a3n2WmZwq9gVRiGiM7uQM6HGE8VLkrKVfLsBuzNU
dwrBlW+YePDkenqtCladNFQVl7jm2ku5QBPPHmBPF7J4fRVMIqvoE1xWO2xSjftm55Z/S6836aUA
0aTg2inwU5k6NlkpiVYBQ7Wo1oLSi/YjxJrbcWihvao6iAzETd+9ToEuMHh71ZFV3LzTa0ZSQSWO
SQCQXzYZXK2M9APkBn+SKnG5XZLR58OpBB2dYsb2baJOJd3vwBhiXsl/FUc5qmRmfOwQTIoccUr6
xX8pwrtUt6lHpsun9XCxYQYGFyOQZcQ1/4xGbVhtCUe0Du+ooz/y+k6E172j2ynHAP8BKDtzHCEw
cuC4zOVKKkLdElwoxSpEReeShq8j09tsOUq0xWwLrm3qel1wab5hpOtzTV4XK7ntz/TijQm3eDNU
mz5CcZyl+nNJY1tSy38zoE2dupG6BrW7tufs60HW77t8Nh8Ii3nnUXdhEWyM71sxqeD4HbJUmb+/
AyCx0zY6CiUVC0bzeaWeL1LEtmGBlwH9rcxxo9yBdPPR72qcj/ntbbQaoFOJUZn3c3R0y7FfCDc8
itsw+bmkc7FuTNldnAtPKA0SZjkXCogju+NK3A64f9VcNC7Q3NZOroa6rvYxFRwjj5xQweIFx8Bw
CIZTSLIybXtbAbJ3c5pEpoCVlM2Pe6lQylKwQymKusG71Tf/aPrwYrAaut06GwIOcaC/YZO36mun
xSYFyriYzBdbdjPvlkWOL082zZ2TohDENsFuqvZyondEzt3ZzKbZ6uUsMrOl3JXYmpew2zCHA6W7
oVz9OJfPbw2e78OK7Qxin+A0LpGfM1b35H64Qk1gDpSzBzyq18rERpaNtnpb0R0Zc4rKDhqaM0lo
ZxGs8k3m5Xz6UEEUhWexkFbREo+uhIXnNYjRatzFRUArkQnlcJjB1wKlr2mhxPENv2CM5wPVDOXZ
5dHxFdIcxKGVt1vI0Mzw9mA2/uaB4FEKarngF9a7vdEazhB6m6uFa6NJtvwF3Qe7G2HOUoNJWxwF
KUahQxWCqDYq1X5n1AF2rSNpjRqVe7p+6UavjB8A0/tAm7g93lv4rwN6OcrUKF9ltMsi68jT3t9l
C7uNXqPAs62E6ZAW7tmPl6PW1eEm/nO2LjRUQoBh5VYtdWYCecnKh+uHc5AO6Lyv9zjFAWrdGAfu
By+5NuCSRaTjaPsJ7lLXKmnJdDihZP2MTlzJMLls4jmxQH5ZwIYBNH933Vl7s+y2qKiauOqFpUr5
mZyXu5bfoLAbThYGz3JuKRgWMvEUg+E9Z5hMkAV8XZtdCJmO6Zk4XpZF3cMr+Lcg/Ojzxy3CL1qd
e/c+ymJOCU8ZdwGZl1tYiTiwDaTe+zXj9UwFTcdQ1sAKVBYhre5+A/QKx+tMH8bGTe48GPThtjAf
rVsr6aVJqMTAWhgG38LFGz4wu2sqKBoqhnTuif3Y85wywQgG0bN2Jp0QFJsb7G0rnJ76GfJtb0q1
gankfmaebwRXVk1qo4zLka5giiC1Yt02cGa34atxt3FgcMor4zlJsrGJ185iChi/jNdyyim5TDK6
rtU2n36g50UAQAgcIbFvm+oEkKWZkyNIELCX3SHmPQVRcdV5dYRJjeZNk0pYFfs3aK2fSk2OxNYL
9jjaWkYTskQKxGQiceX/a1pqAkVD3W0PKCQZ5f52F7NwG6fGYz0TYJrsiyoAr8sZK7/LNdJvOEBN
G2gwn//TCWR2Dp+FZk//ujz9gU9Ynk9lQJifGFC1gGKgvDiAvPuQxEs+4ri/pDTkslX8lcML42OM
ahHtPPfBUyfmpl/niLevf6Gu3rzC4KwJOGN8+KGYdgML0wP3bq3/+wiOebnBe8hfkf6+ArezvNG0
pme8SVUQJ+m6oZZNQ1GTcjXY0ZbDdFwI0f/mT/3YnAbi46mRcUFU8KrvPkn6d3bGnoj6LBfOa8WH
tfMk9ABYr+U/6qgME9Ik1np6mWPqxcikA3508InVV44J6Zz4WQXGPELbcGr0hkjAchjqeDKv8aQq
VjtK39KDSTK9AvcdxtS4ZwdsQyYuHkGB7cT3uKJOEV6DhklERqHNC3c9fyjlqt2wKsX0cpRoBZg7
kxBFkGHp0eiTpqNUPvDwQvySw8TXQUDodfwadjotGhJtTzE4/7TxrjuSPhhX7Bsr8FXsUgXgmPZy
m8uXOVLgU7qmvt8+4x5Ez9cAtLIb3H5WrMSOE09HCMMlj1uhD/0Yp6cgtZ3nUSoW5luy8/gxqLNd
I/FuePBaRp0kYukIP0DBDtQKXY1RV/6r6Bxl840sWbsyxqTL0g1wfOCeISQSylYJiuez1oo1cj0y
F1hi2x5W2lnAq/hKev+xlxCyQjcIZG29vhwxyx+eqh27kWkx4oqHDpT1CC+6raqjjMoeZHcuCy/F
omMIZDpd5YsgKZzgp1kggGqAZkvBUn42kstXN92kmceyZM8KJqne0LDcdqhcY6kHNmnvFwxz6465
xLVBFhwkhk5CLHRyyPVCjg2IOkINEqjgHxfOYHHTS6rW37wQlbI2T0qups5KJm2S22YRvpQJtzD5
G2KrZeMwuP7/OTPfG4Y7V5WdlsxgSWLEtriBV39odoG26eoT3TDhBBI2e8eyz18GXGQ8HrTahcp4
GsdxS3l73bmrYI7odcJl7LU+maqu3+pVRyuA0eC2zWrwRoiV4tGcB2YrCZtl2WQzovAyI8tb2dZE
6C31x+RwauA1PNCLmu1KeeyXv2/rQWLYOCGhMJah+xPv6+T3UjBVmX5hHBvUdwKAvGn+vrbqi3/I
0l5MBiKObX64ALKB9XZkD6bfGpkjkb9DVHfHb+7kiuyXug+XjZ9/xuPMmjuQY73qjfg4qEk6tvk3
K82waNdsr7SxsipENQQ3dGR0S+bAtzcGuA8K9SkxKCN43NQDCsxgQUAr+OG4+JxYq5aupPf7nTaj
sMvy6Xk/+/GGFmudb0U56DV7D2Jw4K8upa9W+C7YMTFzABEZKRU5Lxujj5yHzLDUhD0SezYGNgLl
Ab2ewNQwoylS09qvkE3kLXwRiIoAz9unFi36fBMoMBnitRwUA0iiXti4+41CvWrmshCPKyucuCPo
orcH0GNIbu8RFCTEoT6qSkgFyh5UOx+jL7GHg+4csv6rzghPs8xpUW7DRKi9srB9x+RJS9E+sKav
kHMUjXA4v2+uq4BGYjzLFSxUnjuoUt5kDjA0tbcONdEJNMCJL9dpujcOBLHL9Kur0F2IYDM1Cve7
YCgNRIkL6uvCdrwmLGJHMlxonnTgwHyqkdTZPaeTsf/rEaZT2pb77JifKWRGetI+SlQuxjfBGQYY
snmIEVnTQPaJ3oIuLiHjMj2xtOf7N7zkvvhvsB7Wc3v1Y23t5u2gumTA4jdTTgLzmRuDhuvp5suD
Gor95swnZIRyD/N2GhsVovtUNPI01uzGI76B8MSlRz86eJzY5gpv+DfeU1EGyyRoPyojbjuwTKvQ
JdwyrzKbbcFqlObiYuzMjvOdNNvr9mqucIcCmhUuT/ytOmHAmAskm00qq4+uNrkdUHUMOfAz41nI
85xhRlPoYKKR8FgJhHgZmOiXRVyPbWamhZHkRW+/itr9EALLYo8A6KpKExsqxCUE+nWcRV9+Mt1S
whn243HmkidrNvyL48jqt3PtgguS+y0gEAy2PMT7lmyqCZyVKBeq7Q0e/OwCBasKps4AldZIO4B5
vYVHLF3Iq+t1zamyl21gLszxd8VCChZqyENpx9VchVWnGAj0P44lDunVdpFxuUx8Wi5DKaWpqEVZ
Y+BevIAbJR5kyZ4c47+ArOLUztQv61h96U7hw/LA+UC6lD9uVNNyfZ4j7L9kaHJBiIMEtitqyd0M
mRjPPpzCue1POQj8gISVB8cEH9ENLyOdP39K3vn/YR37jM+VOmW9sOqf6L2D1jXes3LTOCHktpuL
GNp1/yGSap/DZeN24AGTMPI6ERm7h3lg3IZOhljsZ6KytwFiGT65AUHCpklTzJaBZ18dr/DPI0qJ
qljsC2UrTCFJc8fnS/ICmtGAanZkp44w3hXftKJ7zKeP1bCOO6zsyy5Qk0iO61+g2REKhD/d3GLm
XHEwZdrDDBNBMGsk6iiOGnjWvrAT3dko3c5dxJM+sLlppPGDp5jIdmAkWfs814DN9qn32CDIyiSj
XRUBKeJbDU/9vfWG2OZF8T1AReU2rN3gB30Hd5j53q0xmIp34figBPdS4Z+Tw+IVpt89GOrsb9oX
X5ER+FThRQaPieJ0jzz9TBA6CUIJ0cy6Nsygg4VXzg2YKi0epmdFdiCeaXVLa5KmGE3ORhye+j6e
AUNz2p6CfZQ+fppC0Ko4Gob1PccOLz7PHecskwlIGytcJ1LCg93aD7eA/dnNvWlTlesjsKIgvXXy
uOdvTTzrsH0AC1FZHv+1hy5Nx7HcUGrhOiaFLOsI6KL1s0vtuLaeD0ywNbrtw07q/99WYF5tHV9O
ckvySnxH/T2WWh1HYSsxUOf5LE3p9ghMdLv1hE9ZfR3RzPDDYfEtR49mliYXYt4LOjRpjJHH5mdu
HK7xb2HdUuc8Bj+dWonvXsYDeS1LBjIXwXKG2CkuC6xOuK4wZPS13aS0GozMYIf+4S/cQoI5z6t1
fkAJ4kddfcAjWv9/kIua8nFTKpB5CijflroSA6mGh1H7O9Fyo0fUDxv/PQcTa7loKM/2EIxav4mF
GZwl/8KSGq9yiMybJdw+4Gp8+e7TFFDUd2bzIUf6Nd3wBNv8Q3s63h6SsUOVSmoNS6IqGiRHbZIj
IWXOWvx1NlhNDzqtBnoBWi0PCuGkdtrzK1GsstewQUuc722fbQi4LV4XauU4Y/XLkEgsZkgex0JV
AJZQHkr/7LepYSO7v/P5WKGrbxPtTMwuXqTO/fTyU8sDAsRcNrBGOSjC5mtQ8PuQbSTNznceZwXy
aNoZUHMzurbJ+mc8I5dt6Yw7d7yc/89SCDmKTogICHWVOx9/bWxbzF2cFG6XP2YqcXIH0EDTDl2Y
5KvOWnNWZ/QiwTJQ4X9bXjOf5vRT5uZbLHlPUMZ+0sVlHlZRLEu/+hrW8Ftkecu+R1gsSKsx5qTC
vpCf9HZpl6XOxtklvgA9Q5fKcb/pDwGoTSXuTOCIOUo+X/6Uy6jjKz+8OMK8wTiTCdGHBTahvEGZ
Vi6LTysYKr8TZ70P6gfgReNR5ARDxJRiZaptykvlixaS3ms9ubsZuoWyegBN0YLVdVdXgKU8Bhu5
5DhNCMaMXOE5g6M3deh9AHX6N/x5vRo1p2GkDmF9mqx+k+6eFYNtR9F7thfnH4yT3YVsMijuwQhY
en9B7ublhyO+Pbc1C4Ouh74e+1c/XJE6qAfnKPSYVsR/55hjv3qDiwPGdsZHJqzU5YaKwiD3qJK+
LImgGN8If0hfP6ZamehdYH52J4mU1sRCDewnGBYCVEd5xNMsNF0qYRIJZ6rnhmeHKeOlLA9vadDu
y62XPTK6hsAqOLTaebZ4MMNJjiutTBM4g0cg4Zqe1wojjkVVhhyNM6eFu3/qwRTuw4Wu4do9VlXF
2T1XTA6ERrdbYmJvXzDr6fzLxZkHb9Zn0gQqPyuMqixbQmFETMCHR2I/fRNb8asF5gRSYBgtrJoi
Gk6ezN9n9GrhplqrBgX2lsE9tmT2GXF+m1goRJ03xGUgPw1mAx6Ke7pQrHLBnTkj3mHga4DohfQd
jvDIIuJbr4n5L6WMP+4uv3i+2wC4YA+UvFF2UZfybMulec/lHdUO8SJJcVHo8Y3U8H3y1BuXgcUY
50cDPg5jFpcjBygcbdv2UMMfAIXG0wgDr1Pbt7d13t1YkzxzSZA4I2HvK6bHHeRB6uC2rL+tSTHg
ZhLYeEq5vRSzo+0OYy3jzZjOFj7IeSAexw1+gT9fItk728Fr2SDb6DEPKRWBhLc3kkLG3DXDtTLK
qW9kKfkYR5At+mRqeZcgbaDriJuRREap7vlgTcUPGQWGD9XWtaQjnhf8CrIEMMxh2MY+eYHW57LC
aT142p6N+FGbI4CBNlO7NfU8l19s8y61EyC7ndbHC27vYhg2p4f8vyhGr178gle88FlsnaKxVWiF
y5TcREyiN06Bfd21T592sMwa4dARgFSvymbXHNjocgDdffClwVwdR3Rnty/SQAQeN1L8AhCPkWHb
dpyACU8PpXuJ5qa0ppRMkIybrOVRXQ/ZDhYegWQK8QfFCogeed3gLfs8eD8A+RQXyoxHtu5aPxxJ
vv4NE+U5ER6SLL0w5LGwNzloWdamNHVCIuudeqUx+DfgQtu3GXbkASQ0lo0FwXC3OEvjvpO5ndcv
QISAmVh9Ogmwj9YDitF7s8CCZail2IHF1UCG/LvZEyJgbpmLAwG5TAuesedK8mk7Jp2BQuWDfLk8
wKuAf7U25+8wrEeCPa1G8rd7eIBnzs37ukojfR5QcyGDjYEmQSRWI4upQ06dDQuB1PSS1V4DBJDk
Fc+9q2wpLuk4ErZrLb160djQeww3ZVXPjMKowB6tgiN3jGEENuVJh55STIh9qSbrKa/1OpkNAPun
8JXN02VwIVu8r308pFuqA9epKvJG3ZtwCbBOt6VsldMzR5AL+Q666QenP3c4SNoDM1BHCSYyM0dI
gFOXnp11BrDi/5VUL665Z/S5LBlC6Lv1gzCZpFeJNuUrjK+HzIcdoxBpuiRumwd/r4R0xaMsOIpM
LYNYwiYYnrejhJi+2jBMINvfMir00xTS+6D2zrxDl04cVCxhvHn8F2sHIco1OZaTuAvT1JSvqDGI
nYC4mcNlALulbX6kif0lDD9yMmIF3fIKKvxfXP8wnJp4AE2fkNAMMl/eoJnuViBawNY+or5YGOCR
G9NxmW1/sc4iy8zSpBvxvsDzZsKXVVS75LoswPiSL/P4G1SZ6YQLn/4H7yfFPyUkiX0BfSUJMBO+
9edUM6ZJlBqoRUen/xsRP8t9sPvHPQpeFMTB+zcj4MrsPv+VjyARdrS37Ia2HER5ad2rsVggI0Eh
buMOxu8oclcyiYXKhu73kig9PjR0fPULB+PQrZqc+nyxTY8GnGG0ZKUFIRCbRGTWbbiKcAl4cHkA
1umwSrUBkz4E2DJQ+/O8UHKSKfpbbBJDXQLseOUgbsPJWjVMjI6/VQpYD/7xOUIo1eOjZe40Bqt4
AEDWRnyeiozTj2RM8r9F1Bn4YIEjuwJ2jsLU+9WYrwVDuWBwwyXM/zNa/kGUOeZhBVPLKjmQ7sdw
HsacUTa/vS06trXQfOguGeGHmksCf1dmERJpoS6NtY3F+YZc7Tr8YuV9dnVKJO9QBZt9Pp9/A4cM
515itv/obaU1gH5i8xJpWjKvy+9P2JV4y3f/QdLahz+cbLESy/ddoq0YLiOGPXZ2p13uRWgToFV5
vsuxEZO5WI3xBURBVITcmbEyKgVo6Ruu5nUZD/CBEQ1S/L8jQqh1bAjp8xyR+ZSjNUTGqO2u1hr9
NHq2uZyDGs3/UKuDBSA7sUp0IZdv6E5uHpvklq//glARYW/FC4qH9dSRa24q7nKCf+WKV+blH4EN
AqCinPtIJYomti73I5UIqbvNre+0rhv83ZqNXZG2teXTzsezNULN9Q9mTWGiRJYvcNtPkrJHFkBj
vjfa2OEM8in1hdMIBnADv5ac9czraBySbECyFmXAfrjfa7EQ4q2/CEATmS3zkrDbh8AAbwohAHfQ
0rELk5o+PgQc3JM6RHdrJHUAcfELdawxhZV2bQqsBrFM4lZVWD5T/mWqQ7OK21vOmWVsDEJ0b8sa
cwmFcBeTdzO3HghOGNm6uxC5RhT918Z6XAfQwLWnPWxEjWS3zAbrluSBalkcWwZ34Tr8r0s6ZhKw
n1HGrazQfAG+CevaMQHomUug5DIjnPRnvwtvE8vSzPyKgFn/pw8IUaYZprhsGG4i7jatW8Mv47R0
DuY1k3RHKd7LiQBJGinH1uX3XxkDCpXTtz2/q+LNz1DmVra3Yfq8d2gMPzbp5o2zoGBLFPd6Hs3L
vIMKdqvBHAj5T0ey0oZoQQtdKpv65kj8jjcvV+cicicuDCAuk2Mfj2ens0FHqG4ulEJ4mQeYgOPC
JHm9jM+154mhfUbQb3c4XiNcvm8dRDmyXs1mU9FaDkXYH9/69S1pGbjuNkLCqx4wJumhY0K/rLZg
krhVlKGYVnsWs89CXa+RJnccWOjeKethm+FZKxceY/NdGb6WqdYsk6gDqz+QfnsMHkIvovrQZ7FT
w2pMndGO9fFUeVnMtb1MSQeq4gUjAv+uforcTDJwv+4TjjTEOuQXeC8uZxhwg9trQNCgSibouHKf
lcDlvNSsAsS0aFr17KXbzs4BIldCRLlHoDhJ1OwNAU0e1H+B7phUsIy2/Mti0WfVO+8ssFaUa1Hk
p02+3wnDuVpkITUgfmsfVQRAM6n2HpIxtWqMtVdjCwMlUQJCPLw7wWDIBFOE3HDhZHhDIsVjco4n
ettSRdYzWUM8s1VtqYqysgVZnOST6pIl7m0+4H1g2ivXzVGRYPiWSE/UIQgAdswAr/fJUePtRjYL
YOfmcObDY0Jj04ASjACwiiMcGisrqDMif3nVla+Ytm6ao74g7gsfNwSg97DTa6MaqWxuCCYYYb5e
NXFcYuKfDw4GZCd501flbO9sEBFzpZ0dT2zvQWfm4hI2HoZ4T3Bpo2y/9SISIU15LxOAufaD/X0x
a95xpcOKLIzye7Ryv2oRQJ+8E6jIUbwKneHrZkpTgAR4xTek3mt+jPsoAebde8dgA9szh8ecujm8
X0S3zMZ6e301pOpXOxxP1mH/ct7JaIR1lVVzF3kAI7CIRodrw8nrSzfkw2Iwz+WpnJomr4mrxIoR
ED2kt2EbA2Sc2dVBGqB4U8r+pDfuzj/MqB9yxfb6fD2Zzvfe8HhyRsIW0rd2FDtEQ2moLB3RRQrf
6Pynd0zwA/fFjFPXqsRtO+xCAJLsWn5ujdaSLLMwGGPewHZHwEcoHOFc7yvkzZY5I23IUKXCIq3E
xWKeSAGAqyWn/fPtFtI6bCkLwk/hTvy9GedFoWfO77u43ytDigu0Rqb6rghwaUtlrILLofhvtf8G
hV82BX+dDbwYthkU2OCKykuRCfls0x6bGdxIT3nFAREgpA3FpVvf7VUZML+qu2cexPYIp2s5IRGu
PKbd2FQdYhe7QpXUASu7+Xidt/zN50PCiZSwn3dPoDd7EWn+Vbuoumgx+q4ALiglYPyYbYvDYVvg
7ydjK/5+c5gf9Dq+lyCqgbS+/PkdaAlmn/KKutcHHYuNcq8fLuILkgENI4a81Lq+84bNKbkFieXc
d9RxyeM7CBAK2cizuIEb3w8PF/GFKZ9oCHV9p1xQg/AWNXfY802TuElBNlw3Uaut3EyAFkN9J+y/
v9f3lb04m/B+YMeTBaeU+o0nYs/idub0beK63OFlL+i2HJ8NqzQh1K2zBUyhriiVx9XvfBxMNJ7G
iwh/Qn2pRMCldbRiFs1B0kq/ThPn7lvpG8BEsOpejhI9KMHbPnruQwJh7Yd7V3VuGVfukpnMeydK
gXb4fGjnWSDpRm4mzbalJRbV9l4O7gReHv6DpKYZ0SK9pHnCJtFp3Z0MxGVZUmkwcuEHYcasqxeq
kdfDvsUwwnMBLPb8OZyYLoaP058Lrlc0XYRKWHYewOrCyy6akJsP7iCG2UIwmCrsn/0C1MdgXVlx
7gemIwbULX23V1tBZQLz6j1APWQlxXJtRH22uVIGTsZnlJ8S5ejvfhrbEkhLUVKypFG2dCHlpQ3w
DS41m2ss4HyhiAKkVWiBJnJSEXQUYvhknCeCuwNpT7V7+51KsNksBsi8lwBAiwZHajq5yNilW6L3
LKjJfFMtQNHAFLO7ICzGmGSl4P27frFSe5nSVk6oUKjuupzFvK557c+4MFpYEg0Gdx9G8kWlSmQp
wX+4pr4Q4sk/5KXfSZT4M1Oa8uZ7l/KTJJKZgf1hObk+McZPENtTJYcb4Cn2YIT//r9SJIY6f5UK
w9l61/CRAdV1azKDP075vIXZs4XqoKYufx/qwLgPJqrSQf34FPQh27Q65AMiv4smY37gQAlUa304
3houB1zjz/ZpaxurSOt3uBIMcLLdiIpfS/t12KwkeWW6qaupQPAFHE5/01nOf50pNQuYTSHnnN+S
nPWyR7XMqNQMNkAEhj/1XfUvbws3DJqJOkMkrQk7f+zppsjzMLYRYtj+/Tzy6jJZZjlNV4JPiT0d
0Iu0ENEJ56AOk9WbX3XyRmrbYJVXlWqqQ4h95MdtiPvthYztV8bQWSYWUVTZkJHJWEmEWuZJJpEt
dI5NYKjZI7VGf1aoaYZOYZcbkj1jGMRMeSr5lgaBveVWUMcZFPO4BfPY6Sj/r/6LAJD/58wSUulr
Jf4RZwVvBbXDzenmRUXaMWPXrLqd6/zZMqvCaKsCQRw3vMhUcHCKzxDJjIiEoMRVDHNsy9foaIon
23DCW30+5ehT5d37cjDdp6qDud7uV2DM8ColuHHIpdnwt34MYJxMLTeCJ/hgDRnnqDY6TgGZsKKx
q8xNbjxPTESem9f5nZvVQSAF63zYJuTmOCjrIxksqUJ2Md32unCThLrEwbrbj8b/xhiBAX5lbbbx
0ZTmfX/Kg4ctlaor0wy1muPCPcH/upK2WVT4P94tVuspTjxDQ1yTDEwNNUgqnFDsMqoAYJDed5K4
ivx/LEmkIKMuHJ9fBtj6TJD0F9pVSfYnrx0Pq7hyfM4Au9JhXPer3PtL8jYp0CxEYhc2mRNhhKMe
/OafBsrEslExsWAm3CvNxkssLygTgdWOSUMsC/mLbqmCB/giGgC5bST6MR9zfhJhujEu3vTphEv4
5/1iPQBV0PY7DEg2ltn0oiEPsAkWic/lbI1FxRwQK8auYKNjoISsD14aPJlSMnf3wUkZv7+5d8X4
VglE1Oky+UpKH4ovpZ0cqXZmWZZz7yM/IMmfupaP9afoInJAViRoHlWqkEsJwypYxzvKZ5GjWJXV
OUYwUHWQaRdQ32bIm2Bd+4IawqCXWgVu3qIpCcv8xchYXIQKlYWMxUuuYe36R34oKWPL/YaIM+x2
wWtk1iGmqGCefWyDMlYpUGmVlOLh+nLroqX1eZkbldQbhczFfrYwIhJXp9EnChwlf6NaNzQSCYh+
gfwzH4eR9xPgKbVdprgSF3fiqAkCTMRGKWgN93ZkiQKshqE3a35I22tQi3BzJ6OV0WjWTksyWVQh
s6RSjRIZTK7rrKefDMGoiRIU7Wq+1cNLmpfNhmZAqor7F7DUpGk8LFI6+4mHaF7iCZeBkHctUF7U
/iywyOMf57o0Nd8iythVjjHsFNx8n9eyBUoNxz6YT4qfMAgNe4LDHR7BiQBth2kzVSI3ENB6CFcb
q+F/hKSrR2q9kfCQnO+edSLZ/RtDsnURtrc0EbrRRAfHNQ0mbcGwmBak/BPTllUv6EzrxtI9fRBv
HIe6uuhE5/SfI8kuPLzUATqFjqQZKsG2s+WSpklGHXM9vtZJP0g3zakQiLreM73lKieIFpU39BNV
ybVE1+eh16ASIREVN+FQAGOn2fC5ljDP/jOdwSixkwzdYXKIRcSlIWxqFSMzqo96w/5c53nC8Si4
rrBLeQlvafmSVjS/Ex661Lji7wLQCJiaaHwna28pKXSPfemti2er19qs3WRWIai6tizzVIsSo5eE
U0bcypIYvrgJf9PJ4o68/Bhu+sg4AH/57TYrlohSS81ouJPRF28PhjHfGJ1wdQGpp6PeowhS4pYd
goNtohyW6YBmhp8TOoKKZyK9+ucBIlJf3D6N0sHDokf0rm6HLyDMl+Bq7k1JlBn2bQ+6x1ctiRLR
1AHayIZscPL/qCbC8ioeeqrOVKik5izcCB+HCitNQR361EFAvTRC2FFvxZN+yOLiqEpM4PVpBGe9
4RvTP3cTZBvKh23/IsElWjI1NqI84vLLd3Shuk+vGyxs68mTJivH4nYCEXGsKWZY8ovBx+2c1WRw
wsOs3yA6W731jlSlkWQFCDIFZvUWMcslHvqezyOKur8AM8rI3/dtX/vlCvcCl6p/8tnqB+cPlr9m
TsHEuX44atzIXxlv/O1l/3RTnGf8slUjliHnMZKonkwJJC9KeQ/kxw28Hpw0ead0OppLtzMvT7MK
UdBjz/WoLVAMCWSyDmp8ZvvojgCslMLLFYm7FkQ1KW5x23qedcVrl1h+rzy43JkPEXPQfKM6F61G
zAH7A0nriYbdT9Y2lA5dGwLYdaYjCrLNWhsex0cXj/Ifhtq13yikJi4Vyrp9zIRKq0G8p3nfW4BT
2u88ISCr7XrJWQRvHEpwwMr1keiJ5TAFMDjGdcl7bmBvR8KQaJyQz0eAoFJhotMKegruQE8PQUtk
9GLZXHBb46QvcUKvHxY4QC4Rkfx9lRtP+yNxjIKeOJFsOTmmvsbJaxfoliB8rt0oqgTW4NW1frBR
6nIQZYfQH4IiPxhOUICE7wGXiZcphlNgKX+2f/K/7PDnllebFoYxCenipYpVmC+CeUC0NjpqhkZ8
rhDTF5JawIEHyq8zmVud2bofdbDHvk+eBkMLR9KxtRv2qra+iavSbVBKY+NQFMWDxNuIw0aKQsFF
cUoCxRGaY3qsAevzw826eCq2VWGgJ204KMw3OEqnWme6yEbDuxfveCn76u+Uql9MGLZDrnvf7x8f
VeB6qUFWbIX+4fn3K930LF44gP2Vsoao+HEnlWtGxtmY4yeBbNi8M1J1D42z0+e+WoYngjoz8xDz
Ittinzq2ocrxkZCH2sGoyqeQdXWFL7DWWC9aBUX0tb00PU7Lh78LcLiYyU8MntOiCE9Savj7vSpJ
ngaqQKR0FOJ4UNJedXJQCfDSg+TovCZcI5ssGwkEdvQFw/1jTMtCXc4JKb3F0+AFkHXJ73WwAVkf
32IdlmMfsBUbupQD+veaVQn4mQBsdXhdWAU5mkuk/zB/H0tVmtqxbKLp2rY3NT5Yt3rO2bRyYDf0
8m0X5RGiZeJ+u2LDxgoMtcI88XosRwN/pMUFCOBgJbmAQ7MoT1MkkYfBx0zQmcgNbfJQ39sApiOx
w3OybRm25Q1wEeGKJpfloVjPkYFuLNhowdQdZFW7qyEDsOw5HDJIYs2ujefPaxnZs9Ep0qsIibid
d5yVNjKV0YNpYQ55CTgxZqNv1mFpL/m+x66q8pugmSO/+SDwgmFZHPajywZ5uNS128up+qhpkw+3
x0lB4H+eaR8GoivWm4bmDO/U7Q/7EW1Yj/N6dTBow+3xL79UsJVVOIX2U4Ez6mtNA3YyUVPV1DyO
vZ66hge+ysbfA1evJSexnPHcfppLPdI7xyRhW6Zh3MS2IODKnfPTDyNgI7h2y494mONGYteDi1Or
Xz4aYuT1MZThUfZuu4brn/KeCGBsbpoVkkQ40ry+seLUWNV+AtwxdxMoAQYs6R5J8zQRTMkTJ8lk
4endm8AL7q86iPtlIbfvncZBrRHlGlA6wUmpyvcAKoZJyf/q2d2dxGVnsOmvZTeISA5ntExX56vn
+XvQ3PofM0/wbZ+DT/bQRN3gV0DubgyhWeqc+lR/tsOjyrrYrDUyl069Zpv5luyYf4rPxbf+16AQ
7dY5tDxpBcLP2XQbqo9lFEsak3rCUfxv8PtxZQS3lOK9diX2vmPszmH+EWnQBYDSMLIbxKIwVso7
pfblPPGiPFXhI4yJot0q4CHoJHFmhz7JmR2tR/tlbBaihl6NZgbYkJyQXeGTm1XYzn+CMl8SDG8w
sjgsKTciQlPe7MbKYRNlpfm1sn6iMtWf1P2+DTUboLJplRgzwLdz0vX/lh/h9JQjwoFx95m/snkn
AOEDiiR/SJUDyZG7kL4GZ7637pPxTKB5NceeEs+NvL7YtqmDVgnio3hTnK/41yvETMXvaqX0mODp
9SQic+kJf5pEjtuRSZkXrcEWysCD2kYwTfoAMnQSnpG9QV5YXEj5D1XX+Baga+n11lz0BfCy5FuP
6sUUPUuKqHAdDiVz9Xf1fDErKXMd+hl1UkiysqechtJZUQMMU/mrmiwa0EvIZQgpKYWmVsB46y/a
OkIRgVrjYMECNd+Js+4JTOJqbyq5Pxa+QMT4BnGBvfmC48ns4fyXgDXKYF9awewyuFQFE/n08cR9
WnA9GDiY7L8VHCQ9U2oaqWxOaJSoQpqlimNHHcP3KTiyKgNcOrpggdn9Cu+R0UMuv8vRuK8aa68o
dMLbe6xHPs3F17PkKwrNQdyQ2fQgwAB1ti7Ykhbs30+jMNS4WbOHRw5bsvofwaG6K3NW6kA+XMz+
t0DdzqgQNNOqzCDhIwYgAH3iBxD6dJlKq/pnn8hJ7uJljlS8CvXDrE8qt8uKJxA6axV1tepCTIuu
rzA26wgqXk+P2XqsEdED4MmQ8xs5xnnrtAqZZU5AIOp5wgyrB+dGP4kL0Zo8UajMpqr57VUNXfOD
esvinS9nQIxAFSl7WR4vt0406wxUGEFR8xGUOy7QV9MIJw71YfjqVV1mtr4v2JH7MVByn5czuYX0
JVzJMmeYrUlDpmCa8IWueP73/ZlrFiBSXVK5DmYl5FC1MIgXF6LCijifBlfa0G09rxCqMA29YIm6
NS9hQQBTWeDrcxcrYrlQYo0Ue45sYno0CO2mI44DqK4IzNpVWJk9foOjGlP2mog7v1WFM5gzVBki
dt0x27dJCWVyxhXPVaqRrusIIi+1BJGGK+20v5xoLEb0v2baQWsfC2TeJ99A88J+tVj6aQbhP4ak
ASWIX/re/MFbjgpHzCYsbedR1sjHoRzqe40wHm3zlWfyS0eBP09l/xWEUHpBerIkM2dARDl4GIUi
lGXpE6Qsej+OmvyVWq9E+8o7RhxOVQXTzBTEbNsYupeXtvdVmEcfqjwZEoFcKiBh8O/zxUTm6SFO
MCkmCIzXt0KEvz+bzR74ECgEh1xy2FAcjqTSlCTd4yf+x2LS43vNdHGagMyPsK/AEsStW+jm1jqn
0WucZyLk3ie7iQXA7VIPtdnzHhXKktBSFHPJNH+30wSJob2eQRymkl2tgnf3tS9xL7+oM7UICy3Z
wP1qDwnPDOjIu46jn5VszoXT7e9wAX7i25JFKMG4l8r0VPUD6rhxSIUIb63U3/VtHSvOc9xh8J3d
xdjcDqbpteHtmTIO9KBh6BPbF9jZwPFS1cN9M+ZIILWT4LXD1vjkj+bWQ2hA6ZFrDdip1SwY7tzu
eDsIAMQeG/oFozBbCL/rpm8HRHGnOtQx4EAgms87lHDQi1/nq9x4wzA9VjAwHb2JsZqT6pC7SBE7
tCua1wd6TkRexYLEB+RcYjpohIntoSLwcv00tCydhv7NXuBCE8iMlBkfokEHP2PuQngNYX5fxbEj
6fjGKcsE9CIw+nPCN/xkkGGYXnMU6vVfwkfdi+nilD1UBPV2tRnB18HN7iy9I/iYVm/HlZMQ+eL/
ThEewuZzYgsZQT/N0LHPrqQO3Ys7/cR9vLIUDKzD1HhuKbbE1LWcBDKZ1+VUBbLKmODW0Fp4D/ql
kqhxQjjSHg62TsANDTdcPEEAFYZlI5gv37yYmt6Ax1XSHwi5Mp6sVTiX5VxTQxFg30T1dfqq8v+R
SnC9VivpxzVJYcQ3yQ2kTflx0zQOeRnQ6YkKznmzi9AWFsXq7cThhtTzHsluQs1aemXduzoNsE1G
ewcIUFW563e/SO+wpnnu3H/24p2ekgZyeJlEKdyntqeAg658/CEynCJViUZP+zICQVWb8Cf7Tg+Q
peUqRw97fWe1wmBCpG7bXhJStRsI1+Wjlsv1VNNWr8keKnx5vBiwiA63WKatKbl6Y9y9RsjyoqbI
f5E9L19/HCmzNh532bU2CaYOwBQvokgmXwf+Cgdn6QxC45XIxJUyP0zgxia0q0VpmIAAE6wHCN4g
dw1IpJo9uqLu+vZUprM5LDay6dZpOSkEZmmGWXmWUmzqQPO8CsGfxTmUT0Yk7vTDpm7XLW4Re4Gz
HYUPAIr0QJwRsjXg/fXB6oeAQ0gCqD53TW9nAHQHrDfudNPRF7kwssCiW+67e5GPrCA/il5Rm2FZ
RBKHElNZvc9keHPMCbyZ5l/H/uC7zmPvffbkvdElOlM0Mpe1rRwKwALGTo4VKvuqkyMQ+U2DrlDg
NNyX0DR9XqIjdatCAVkC0z6UehO7IJoXBAWkCde9R/4/wH2HjEoiryEf8B6VoIybD6wsEgTO5aqw
DMwi9f2DduEMgX+VJEnwTIOKidJ2GiFStkw2bm3iWmsR6bkV9lI4VGDfmHkBoEv9W/WjGBRaFsUk
U27TnWXgWf+vOJyNyKZTd3Lr3YazlgZMP7fjUzsVRr0Q2KDFK/+rFFvJV4XhYxctpTILjaJOd/O6
tLy39LB9mQ3BGmYD8+7jCQMCJ1cajuFIoMZot6+qPVNGM94x0wZix4CUc1CMURuN7P/mFAMA3bni
M+SxAic/8x4ap4WljeL3OMnWvujSUD4c12UbmNT3Rr1VMfb1zXt9K2AvNsYp/CzBS3oWKP4x8AaV
a1OGo4ZP5jaAQj62H8luzUi6CgPsYc7gNRxIfBZZvWqX9VKoPVIHsqlAH2qt/m1782USIOZ9OT/Z
UFKH7qwivG23ye6hYlswhptxcOvQpfiYnVe/nwjv9BCEqgyjUqasBVqAwZEPLC7YK88ijIXmbf0f
r4Z2Mk9IC2CMWcQZuEQyTg/8NhZ08McxCwTsc+9AxT0ohLksac0+M0luNNsBVabCsCDB42oDzbZt
HgDNNNHtMIP8LtwacIoMvFJZrwY1aeBGCFyfKhAyMA0TO3CSMt/6nggSo4JvPh1tD9mIa2SJS0xs
nQKGsCr8HhBWP5o1L4cYb5tf7zXWTV1HaDXsyolq/w9wE47/PGPZs5sPwpdmcpvqWzAeXqHScYUL
bq/EfY5F1kCyhEN+KZoRGcqSLRFB2n1n1xBIhpIf0jf4skJ56oPveUR3gb7n/vr26fAchfgnVjGn
emPyT3CthRLnRSNd/2MbRmTsBy3PEmWiq1sNN5qvcjpPLT1/ryxYZrGex2K++GV3gmay60zrqF3q
wMKJAcSkceC2vZH1VHQblznGyl0LfQNe1rH0h8b+hnF1sgqNAJsDhPdRFyV0zNVzzSPS5B/1qrNN
ttm4HSRatYlzPti/dfA5LZY+RsvVrdCjbBLec0bKbb42hFQPaSkm0hAnWi1JDjQ39N1Sv8LLlRDL
x3JxvfkzMWeNEqDJO6P2/eYpmRdZRZ2YrTGm/gslvLpsVxQAiWmojXw7NhHlfICX0nX3BjbWhbGi
RV3Zzst+ielyzpO5hm3wCJlhtbzFJRIXiqgdV7h77DtbZ7C8OAj1CX6uwB6K4EPQwlcGVB92cbqO
zZZ0B6eSWcSpCqEoKtT9DiUtc0Wc2xE2IEiNrC7dW99cx+iuRgwPa0G7m4nfHUPgEFeI2baWGGr1
z1vZHDjj+HSH3wk82ZYSg+bPlKkty+MVHu+O9zLjYrzBkwGlt8BUg9a2VzmL74A5zXmzN8Dv7JsJ
ubXRmX1KtLNq366ibtf/0n9ZJXt35g7zmDzwhyxHKwc8GT8yvV5FAKyTQR2/VbdA2o276esKG7K1
m2GGcfP/PZgUYdlUvilOQ1vYXumld0lNWlJVN5kLJgB2A/iYGBcfJ9pVDKYT01Vj8qQ3sFzoC6iE
xUuNbE1bqkmT8pq9+WyX30QTJ4fieCITQn3Yi0x2MPvHXS+f6VJyjRXDtXtwZbE7nayke5+dJUz1
ArErIgYv1Tk38wEo4IOXWZvvpsQVpaK1n/8Xi2VMtt6GASTOptq3sXXwBn6f77egV6bJtZ4C2CkO
2IF9xuaIXF90mDpF+xB3I0k34EY1sajhAuLtbvtX/BrGZKynnxXOioVn4KiKtLs98B7QMYlU8MmF
GUG5zTx6+kmaCe02gP5J6lNMfjhCrEyza0LCro3MmMou+U1ltMF55xrN3nFCkkGpFTYwPFLsx2ve
NAa3f1bF8RKRF4oRE/CdD+zV0U7Iaz5KQtBgzvuFJpTr8szRtZP8wkdvVUXcNQ0pboGFuz5cNNlg
wSqtRlvom5IxVhKfFzZsMFG36+g47QW8oquV0jUQnNsvTnR+CR+CveDOdHIbfrAHy/lBgodiDoti
Z6HNG2Z6l8gN/9u30SteKX1QPZeV/Ws28D0yEtxuCMdf0sIuBxGa7+/DiStzh0NT1Gz9V/Yh55Da
S3+UD7hSBl/jGW7XrdM5UC3EcE2Qzk1aAxnvsia6/TwlNCOMp9ZtEwxMh93CVd9GTK+oOQybeE2o
Txji/Sm5UXzzF0x897szX1rg4645PgDgetCfr/sISPtidJOBotOzz1m4+vd7gitm0bhVwT6dav/Z
kELetnaZFeOegW4QmwM5zxH7qmMjxwrbhZKYgZXDgwA9YB10h+nBZI7xN2qfcbY2Bd9ZT6R/paVD
hiQssuYC+JvlSIw+SEDZA8FRXcRnDoMrGcqFstcAdxfzN/pJR2tzWDnGNBhEF2yhp0lOKFKFYrP/
FhyxjXlvEXBoJeWGIJ31tmIev8pZVQFpcNJarTZgGSuYGE7nGqnbviJbYq16YJtigHBJmyVB22Fs
+cJBt7vk3q284wuZHVHOEw9IoJluYa6qaBl2ViI/7+tsmOg/PbcInJWOVGhX/MC83Qro3nGyB0N+
iZlQeTb+1AFS4u44SaxszYqaSCuMKehJztOEOYW1WeCwvId7BlOPUc9CWdDnbh6kwqi7k4oS8bXP
ATCe4VfvLI6HX39SgeQ/DDvgPifk9rRXh1DK7KfjgzeSEirW0j1Fk/RkCL90ZQXvSIORVIdOGzJ/
dvzsS07edxTH4KRRGXtR+X2qz80RSLkHglHxN+vzzZDNeGeevGdawHhQcULWrncCwQAuBtY0nWPF
qhlTwM/c5Pb0tyCbMspF1Tag9WkX5K104D+N25zuFQd62WHCVsafR+hRgK5uLG03YUGQgVCl3TGu
uTJxOrhwWu23E09e2OH6bhcYLpxUeUEQ4YMLbDR706P32odOkldAc6JL0vlkVSzeqPfaMtLc2bvd
Qb2UVZ0D0qkSlzNDOb9m7RHZeI+7anp4Pkr2VYLSQyV92LZ6FEvB+H/HQDS1yks5u+rl9X1k07s1
lD/UmXJd4ARkOdvtxsBJzyhg+8rZ2jmfQsNCz82I2WLEJ9qfOHfYwVAgvuYGM9TtbKu76QelLK19
8QzQHLDqyZ3nllefW6wL/vZRBTqnwRoFoY5dYYGrEIu5kVjBHVvbhXgSezGn37lQll0JCYHDcA7h
qoR8tXECMdE9W7ev+SCgtqq/O5FjVxJyV4h9K+ll7jbhTnN0vFUwdwqqHXctMoRTWUGC9pDAjxty
JBZ5KdxnJE9tG2W5GhW6PYsAbLHWQ0/aDla899ZtXgEIeP4Uwk+0tB1P7WPQDyiIAEbRMLGFbqE5
7A6/v6a4eZk4LomE0dR5aDQcYX0zS7YGk5rkGKk3khz8f07Mg3og62FDWWBj0obBxUe9FdUh4oP8
+/USCijdV/OAZhKiRyTenuEKoofDA8jjnE6fqPMRP6Fn+tg2Cjjm+4Qbi1/OXgYzVrOyaxR0qRND
ZXIzaIyV0eajtwL7CtTkleAaL11fVPthXz2AUfdOH+DJJ3feazLUDzdqJ95XRPWgfBZwgL5L6FD8
GKiQKFnACo+7XUAursKUgwJOOfmHmSTlG+9dWtbTP6YBsNTsbG2M9I28Hcq3cgrSo4aayvx8IBQI
XiBlZvEq0Hdgy1NT8Io7mNxJ2Ih5b5KcKn8E3Ury43Q+ZU/OdSkwp499Ixle+gqjn5zBDgQOkLv2
azci9CJovPat1QRA0VogKCXhzXEz1V2NZ7M4i/C2JL4/gjKHLNyptg6kb9CnGpDbRv/D+xuSIvQ2
LxS7D2vKoTrrlg1HZ5j4uBOvP1ecL7mo5ytAsl3M+68VNcrwFX3IQvbnlTfGpsGN530YbNHGpenF
OZciPhWBwh2bh1bEwx7W32vXK5cw9iOtCN3Bnwg2Zj8vcLylhAu3aZS3BYYF4Q/1m2ltcJpVLh3P
n7cKOIVfzYbEGXqhaQqUSn/A1j0hOhZOZHFZ4Zb6U8iXCdYBRmSB0QWmDpmjGG8FLEUczbZbos3i
hbZYVoNSW3Nr5W8SLyClOQUDPpWsF0t4WgAZSMOUqdxqgkJk+ac1q4zvDw4hje67yE0nxG0R0kPr
NdEUdU3YzlWqsBEqU6GcQsRgpspm9MHKkNL3JolSP7S7Ki5kWBy1rBkuVT8LndM1rr5kD/zDPk8F
NPUuj/FyDuRzTO9MOcw5XO8BvRAdGYTJVM24KBFicZfaDPfsgXm0VmHlX/bi3bumZO5+I2YBzDYS
n7rDvWT+EQTyWksULzyjjAFbHa7ZsE5njEIW+SsIP9ZW+xoGuA+SAGw1CHRDeh6c280Wxv/mixrU
OqJrR6Y+XORsgEWTcQatxBQbDntkKNU2RYD5BXdsF/7KjUne6xXLZoQ58lJoqLsu/CZavCsFYr8z
OWLbTeBnFDFTt1cW0STsXuGvYidUnCF3159v1UHWbR80JqBrWrSug6PUiPz7oFhw/q9gBGE05geG
wVgO96EODBMHoCGT2kdq2QjWx7OBw2AJp7cFxdzxwCbYfXREn+ezhI0JvUbIWehOZ+11XktTfodR
d3NTFDh2F0zkunYd43onQf88CoUCwgv+MpkvtoegxMx8PmJ1sSba1KMIS5S+BFF1pxOArvu2c17e
4QvT5qo2yNA3CUvVJ7RT4u/piV68sPhDgcRXNB92wBICleFZUn/mYbBenqumFbisGrmAFYxmdU63
5Gj4m1h/NzWprig36tztZ9U1w37nwBwd/wM5VLTv2KZfNIrDcGE/QEO112SCU4074h7BYFoa2Qh0
0QOGXVQkPqNPHe7FLkTkPQG45vrja1/ne06DSuKIWdmFA8/5RVvFrcNz7jBUpPD8Q9hvzOu2zPlM
+Fa1jDS2BiMA81nACcsnKUG7iRg/K8LT+qtKy5ws7J5kMSpkG2W50zwH1NxpoE8SjmydwP2rjYbz
S6/PYsZMivoV/cwVBpecSZ2ShjlvLHdtEjW5n2zWdwZpKmTmvbzu74Sxb2yHNGQdvx6l6+r40wCr
8yuiyGHXYL3CnlZ5IC2b0+i1zXoT8eGfG2enevmZXG+QKUxwDhlpMTMZhEr+gFGhM06MiXKYZFRw
ii8UY+UPkPZqG46uOzUO19dLF8Wpj9O19jOWFOFI0XU8c3dpw7QCo5eppMr5m7y++Kzwmq1YIx6v
WhxOB8iTHKatno5xGuvQIUwKHgtg3swpfGY0+asDQyA6sTStJEDRafcivExJVox2rp36viGtQEUP
bwZR6vgMj2XwtI5lzTFkqhS/wuHTbSgTNgrUUL8TgL5gWS7KWdSuyh8tojaqUP7WqqEGaAw16Rlo
/cqT56a2MetBUZ4YnOyb43aQHtX7AtVoLm3yKHT81VOG6865B1JbGAB2SAK65pAeI3zlM2USLVd0
lupsiQmTbrxikop8hDDuZt2b3qpWbVRenOyqMYz0iE715j6VwpE5ek6D8zdDrCyMrK1t+Lm04HbZ
wdU4Kg/rs+WNoaDh3nsFLCal7VJHB0DXJGxevz7zsl8WarPEO5ftn9Xo0jL4Gg3GgxyiUszy2qzu
CoY9jUYY1HSkfxgcoxxGQcZinSC532BuprFY+nMzGI/5gvGAhzwVX87I6W2kALITe3DMRsrmVXM3
CCzM8BPeYJTNWUK240pppK6aSp9DgMxcgnGJ4Z1LKLwKrH8KEwrynmiK4b/w6NwpFXMNyqC1uNCL
Z0wLDiWTCIHlsbqkvVZ/iqz7dovZJloC2ACJTRjUx6JaB/mahBAa47XztayHFZibRDoojpFzbX/Z
YxFVPxUrVI8/1ejnDujlMySHotaWVyamzGJVMaUjLyneNFdCLCTkbTHRnFQMniBhnP0G5oFaXH+E
+8BpPDYUK2SAF7tSZczkRTRwvKW3BuM2RGOdDNor2hoFUbkas6q/KYxdBMfwtxDjuk3CDrXR9tRU
rqH997iq5+hXzI+Ok5CtWzx1m2/ljq5xRLJuEOrB7dWe2AVJLCI8nDCW8nGg+YrH8cAfDQWhxxHV
qZYzi8S4ephqscNoDukcGA/sp77pgnBLB/n5aToTjpXEjgn8cOxSK8T3Y7KVM5G2uhh01RG2Kea3
O0RYMyjaLZ4ah7LPEDNvxPbVyTFCG9EzT7SAgdSinHk3L3mcK+a6G3tKDCxIyWDifZ2o/9h+7bc2
LPHyZ6Y/XIb28eHBbSsJOYpFb3wwbbcRf0NFBhXd70uFwqG8HFIT1cW+ymh1RupW1gEdpvG31Iu3
7FMBK4Iy7Cz8ik3Bb3J4FDi83gHVLtAxkSy7+ja5kRfun9nOIS41J1Yuvr0J20/IGKzOXLaUVEG2
SFj5dC3As0dBTQlWk10PIwisytZrAJlrV5FxFxbZwxa2iEdbkFB5sFHaiG/LeHzdhLr5c9aoTjyh
ioC7fUnPIMQ2cq+1O3in6xoVMsrtfRbfs2mHSWyr0AXzMi8rSASl4mtSBCwdCoYoBDOf2NSxUkd+
6QzFpvmlRt0zezCkaV4YWxra3esTpyH9XieeDsooX1nIxrK1HX3M+uIc2H4qWW7iBIZbIUKFNDpF
b0FSQC6UJz3MiYdwgP/12iAA7qQo7Bcwk4wDg7Sq2ADcUU76PuhnjZHHmaNWXYEBBzhrwTanOv3U
udwjpwTUhfN9zJAGMFlNt3PepKaEbllJ79wZk6+1gnWHD1GaBKbUdgUNOApycomSLqXuwCy6QK8O
ZWBZIl0t2GiNgAxBOqpuQUwIbgYdOxUI2nLgTsFXGGQImWnvPriGPc0plpEbwBs+8glgKttbzREd
vWpuhUW+sGu7zh/ghVWMgcuRkmXR0dHkIwao4dJOsO4bG3YRvdpXXA1YIVqZMcdYuBeNZ2JzpJux
n8LmcfzCX3eyKW3WAgMCThwvvTsvpjhqX7KWD7olsrSJYU7xnJRGkBuk9seKrCIdgR8HNXonnpF6
AW2CjNyAOAimSltrk5+KYHA+CMakykBZS6U3XYn0wquHIlX9dIApeVkbYDVBjJu5qJSuFTUh6VxQ
qk83DtjKXoI6hXAxZus2qDc37jRHlf2v07o5CHAZjgEQEChr5gxlw5IHMTqeDk2FP5uwCynv+puq
WTuzwijDZFOf0rtK67fOxR0TG8CYUX1GUa0TCop72in2HggvpM86PlcQG3HEepwsVyCvIScLcuLc
HRFrnnX3HjBpyVpvuAjUdzrplwJ1tNlC79N0mOSZEiF5mqstvymFpMPmXoy1Q4K8YgjMXEH67tTC
1CXMW5PB4/dBM446NC0rS3QmMuEx0q3hVZZl012LXEQHVRl6ZmCuG2h0e23b98O7vgkkNxBwPXIG
SdEZI3rFchi0E47GHOeBqmXW4/kROiyOEbPYlRW7t4sP2UU5+fiiYT0aMInqJmzUuVsn060NgQHQ
lUOV9frYrupvH46PL/q4E6DNBnMbKOOPIz8ZKVy2v6jxoPwjd89XJAMdv9kX8gZy2L2kdg32OqK2
V2bGqYpSuGYojENVGFmgZxv8qs+vz/AhIfDiqBnEMp+G62nvLs0YUc72h6XxI/QwUnQAwWCPY0nJ
qDcoT9cjWxoSO6D4ycuK+whuUMDS8zTzdDOjV9FVAyAgGA9q7Yp/Z/T3l6dPR9Vymum59tM+bvZN
tb9JdSjI40kPWtKPz9bHFf43zvhyV/ax5zC6px5hlI2ZimWW+z1e/ZgH9Cbf43aE0N5sQSu/SI/7
3j/cPR9jH69jrLXORYxhBO09dKn5pcs9khJ1zdJeZ63MPrxK0jZaXA2cAScibbRFJF+iF2PwFQbv
jxwu+PHtsYz0a0zMHjbK5M6tgrzpdkqa/SPakaEnJ3HMQeLW0naGenWCO4DIddaDl1caI1thJWcP
WC+ltP96jNVsMrPjlCrPpIWr0+IU+5lKEtUvAY6n13LC84zBMTPUFBZNjFoavR/7+t3yRGuoETib
YB+tg+ISrzWx3tSeOqixvOb89Rk700liGYND8IAzavGr/Gt9jM1cpleTwW6q8le0kLbRoXU752h3
M8xM/NnfUNgrzS0IMChA+mDfU1mtZfiFWSqLj/6Xx5oCognnNYsfLv42arHuhf2kkIuNLoAll7XW
mzxIwjlPZmLvLfMrP8AlETafSOBqnnd8xHbRMICx61EjOj/rRsNAGQyqNfmiRvuU+A5m9La3cr0/
7uz2oZfMS6iTXrHOiPgAfcR61RvNtcDTTJciQ8Sbo2iAXdbdjxFnuIyXHsaXoJFpOP+8o0Zfv9XR
aAhfUsOFaDnfWnKn1lUKWtbVSImYBZ8ycxbWs57RAHFFl0Jc/aapQvf3+evoVz41QHq3FkJKTMDk
5Hpv0+A2mqIN93fEamX5dJ+l88q5IBqUu+wjSqSJlgNztWQ4nKDnD3z9qjhrStLHE3FJvlPYDIfE
9ayZFvRJwaiDfJXnBvSGlqfcVO+/xvSxzSvaVBKfI/arvWHGz3w/bIUuY4yN/fwJS0g39hTwHVzc
6kBKzYM9AItjSM5JWmsjtR1OUtWr0le99UlNuFhoMkl2RZnhajElj4bm3FlLaXiV21sE6cUWGHaP
/j6AblRG37XHuuEs0m43yUxpi0E8EpywgTzwsg+f78UXWWeAAo5MDhuZ3IV2TF1IfaGQU8Yn8FfA
lUqFM+E106016Bm1akrOUkDXypLthYphWcF1DcocGv47YpCrH5uJ8ZbPdk4yqH+4mT9B19ykBkyE
7bW091R7dQFThg52b1kUx2RjUrMc3hCNu04H44tFRAo9UwFCl3k9VAqnTzVp0qKjxHyfcglctRrc
yUNHI48j4Eo1cm2AkSXlvb7LdOCd7QNfeTeMJSxMJnE+s4sHtOMaOUIgrbLZs1AeNLBQfzHrwkE5
7LNdtiIyJrdb7kYiMX6cRiwBOhcX4nn7UrXytfcvqysk8sbTehPMpMZX8X3oFB0QSg6I9++vLctD
c+YKyQkzSYn42eGPiUomZx1D0BtXxAZRB8zchWNj6CjrPtgef5XFtHPv8CMVge+/LhEI7VOWv5mV
Jo3wlVh++bn7PJWKdy/NVPBGGC1YgrGE/6VccZoBBr764p/n4pl/eRNTp/BonRYUwXBV6VRmy03v
WVQo3Cy+cDo+GAyjala1Mle3kvDl4HsXOA4Ri9l+Hfy+tA5PVO8Jwf9e5hpTHUHnULn4vZ2HERTr
9DJJ8qRbqQ/As6Ak/olXTZZOU27Lc+Ms1QJK9zVY62S8WiKGprgC3M0XA6J3fJ1NE+VkuCDiiJIq
3AfTJJEKV8muOUt5j3L9Zdv7/SorFVHVUROAtUArHVdyrcOBtM+nygr+DvBh8JuC0AWOZ6JvBVrv
d0Sq9w1Aw96wxvLBbO0CnupHXT/J68lzK2dhE3FATpFvLCgIVBTljr0+hUd3ylwKmYYS6huyestz
fvuJgCMcR4iz0vPUPSNLhWxJY0ATSs2p2nZdjgK6k81YTNJQFsVnRrK7PnQCaqXVo4SXj1MsxuZB
AbQOn/jBXX5BwFMVEpibGAXk7y40KvftUcDpL1w2Y1yzVU8680Ry4bHzvsEQNg2PkL1Ya5Z5CL+J
S+5qInUPKjKdfCiqTnFFLiOiY72/nao3nhh+kzWcCDDE+DkRWmi3XhfsoYppmwtnYuaWLp+hemcP
Y9jgID3AQIOGf+YGkregPrIHsPXq0GKnKOinptx9V4Shf7Dl3y+MPlo5spp1r3gK7sLcgAysSJcf
3TI2t6ynbM2IdnXddu79tzo83AQouOoYtlq2ZgJQtnOefTviXb5UuB+hjfl9rrxd98hPZvmKKiU9
bAGh2eRXq4bbYUTNGD8M9QL8p3ASVo56dn5N2NZAwEeBTk4ePtm+IZ8b723A7TjFanyMzielPAXj
2A1tVjZUFkgCX+oozcaqjmieR2NzbyCmltwVHrIucGrr2sBmzcIDncxLAcY6sWGtS2xqIhzzdx7j
4nU8rTyl8DdLQCtL/Xdv0kVM3x4eAxVKXLwO4bUgYCEQQ/XHP5t7uU5vGI3xKsgWHzDYeeO31kiD
Xzt4k+5Hvcs/rnNin9IgHUes4b0Uz7Ayj9U3O8ROA+/y9+iI3nSw8+0Ryy3SkB0azIPK9V4IRIfS
uWPaKRbvQDJuKfzF03FBCLYN5sehaZ4FGQgBpT4XqKQKwjYXfw/kiYGSSlYMoFwmnG8nQIZjES6W
GFaATcawbQ4dUHdrFt+rpYXnOXHXInnKfqc8WWQb2u/D9GvJqgwuMUCBVSLTyIoyTs+9tASOxO/3
nI42m8GPWAafjx8ZfOrBtPav32tzU2I0+vaPAWw2RDGjLoaLBa81Yr/LnV8CHu5pXK9mYsg/C2sF
lHi+2mxojRqMAHFeU9JWNoJ4lZQU+Px+/DVd0jhpnbsIXhaCKfCao5Ow3XGNUgi8RqLbpsNxr/4/
Wf2xkHMn69CPLoVWD+nwcX+IMlasdsaFU/agkZoCH33b+lXzx3vlkKA0PzpQiLjr315mT/VO+85b
Wv7r2ZTPJ9Zd+PwwHERH7yAjoeHeTYv2mNWJW0WnAZB5qisMlevfUE6/2SAW0IXnL5TGN6JeR6IJ
G6BwR+ZBwtiTFz0JAn+6BLrATB1hXyr2Nz8KlazMT4H/d5fRYKUwwYVJIuK3x0WnKF5CvBCkp1yN
4vsaBxY6uRc8nK/drWO3AaUCqvKMy/bRNFXgx+GeuJxWOey7B3XmLU2zEKRxkPutwno0Ozt2EmfT
iFgC2jwbsT8PnngllLZ7ea8LyU0bO8yNSOmnergS1Is/i5HJQd71BN80heWblYlgHwjsbIo96Cq8
GXrrt8fPHumTEwjeTe0vetI75OzOkQrPMO3lfZrROLRjI8IjwCCn6OexwlZcv+h4/zihqbKbERvK
C6pRZq+TkFa180/OeDG/UTjhh8lkv2ntKQK86gI+jFurbDQ8ZkwSw0lpIZaxwcvt7VKbfKYOSjBY
zdOtpBcrF3MfEbnegy5Iy3BAjstV03OlJ4GPxeMDMmd/UaTxEIzYTnSPWHArYt9dXPHEoSKhei2k
Z1KFw+6C2OU9HJ+osJdgpWvOn6+tAC0WXeWJSrgy0O3I7svEjYyNTxLtC5GuNDXoFtjHqfW97+8i
HsREjPc6/OVp83vbTAEMUTCUiGijBEw2tOTeAPshHK7+bsYSmqVNsXxIK15LkdIDH12cOx5kOZ8W
0EaFiGm4Qxu3x77F2f+uDMn7YbCLUwjor3CE1dy4xEJ9sKFgrKwSu81+Vq67m9Uez1Epfr6Fhigj
K0/px5bznGv/5ne+YH9dUC06dhlGZhafDGD2eq32B2OUIPGlPTnzGT6xT1Uk4AHywSVZggrCK9wx
138haLZX7vAl5nxCm7sUozNz7S3WYyuBg2+yihi2qRHr2NqFv3e74/NWWrZHVnniYnwuxj2nWEYj
hZcmACdmKEC/Ys3AYstPXOs+q9XG7zK7AbcwpgJiIFySOIjxgWx9tEjZzErAddjlHK5ZIjJeF5Cg
M2ivutShvbVGZ+p1X7h+sYGhUpMUXGutA7VsQi1/C0a+lOsgjnsVqxDmu8j/gKiss5esuT8xsp75
uw7LZ0+KCN+m6bm5LiajNYxFKy0426PsQtisljPGQzgCtjdLffJsB9GZfzHcYtX7TYE91Qo+SDM6
AmzpD7QP/fTAdHUKBD5H3aEa0NMy0nkIrHZCG/+po7vi6baG30Bqck53zejLDG6KjNUlK7sY5JlK
5oSisS70pUblpCT1ervpLjZx8GvEDhbmiRM1PH7udFSIT5eR4WQkqqeQzTSPrWGhDybWWQ9Yblz6
NWbZAf/RO/aNtNWZRSASKZ/pGLIMoJ5WFG/nJzYOrwytgeloYpXlv2gEriFnVR0Rjv6J3w22gPk6
2076m+NHYQwFc1B7KQ1kQ7/v9JzUoUd4+ctS0lB9RXUdB+GV9MUV/7+q3PNMbkIfRA/w/rHLa0Xh
4S232V3DMCjhOEsEMRnbfXyH3GDw0svZwzeKfr+NHyefCqVWqSy8yqX4Q3G2LAC/FejG79H3Sa/I
NvyQXHVvfpwKfIXYUhHFynjX067AO/TiGTkSqdFZULUfwKHicxhJzmjmk+z4C/RsMuoBN6jAEU9h
HSgrKFl5QFeKlro+GexycN87Ii7iO1jgtslon2uBBFsM9Py8Zj3L7X3pcKgWC7KEWo66XFIQU7Av
LCwKUPBqdUcQ3/3LQ+bwLtmIEz3yWrYhJI0FlX9UCfcMgPJwh0c6xCaIRfvAOMaak8/kNjDNeZdz
ibA/gEVBJm0o9weM7eWvEwgf9srIsA/08wqfPXYdkU1dTxN324u2SfbdRXmjbkvvIeETr37Ajs10
ttw9lHMx796UeW/JI9oSqOT9+sQ3xMiCjaD0LpBp9ImXbBeagULJ7tpRsVd3ybFtc9+toz63nEfJ
2AMmLvwftSVsJA++HVHL3n4lU7gJ06gufmXk0zyuivLlIzhA8+iInsSiip6jayaD1G82s/Qf1wVc
ZStqgVn05MMxUrn7TJjyXsalJ8sCMEnXEGwL9NqscLQE+1Ys6Z4ghBB1BAX+DFja+5ncXLgIdbYq
fk/ohBO4yFYHoT8xCat32mQub9kDKmjQ9n6aGiENDzLVewwZIeNEAbNucdE2RmhaFg7M6VyI6cGY
2C1UO3wbvvgMgaZ4Hn3ctANzPbykLDgN9SedBTboIzhnd9bWxqWPz0bdiZU2mz5kxwtUxOR8QI33
L0/4she3sxipl/Ll/H+FGOKir4H4C0iDRmPg955wUNWh3wqnGScCroujHqT69XxwW6OPslRMO51f
svmMyItWr6/F0B/ZJcefU899AwWir1wP8QrGSdpUOfDdfOmJA18i+VjmmGn7kez+stCMokRLa+ah
YCkDAUv71+L6GB1sGyzVdKdsZNX+BJAZ/EV08t2/FL5j3MUVvOafh3WtcUrzzEqHffZ0sBMT0erZ
uUHcpHa/rWCdFJNBoWHSS5+DsbRxrkMjhgPiYG3J+yVlxcABW+w/QIADbHlWbowWnbrm99h7NWnw
Xaawyb97GP/t5IysMEVVplTPckajK9ONPGlLrPD1A9fxodaYBAJ9+H/xeG2h92gp35FZ5cmkvbXC
fY7WI0Ycpwvs9nv9OyMCMFon2UqF3lyDeWN64ujbZlDVbHBO1Jnq9NuKRuFZM7gP7kPJ2dn4FqAD
UKI45OYl98brwVYqgemOVrGrGhGzSMABz5Hu/vEnh1pasZQ5Es7laDbFZslM92Jld9gBr1hF5eCe
1HVhxvLY9PTy1uwkpq9D0/MCudvkuYUugNoQpFFqSFh0zTRYVQivCCALsBiXtHCkEG+xvDdJqM0U
tZFo/ZukeCA7P510L1CFO1yYHo98fmBjcunTkzQZcf8yYTaXWyANiIUTiHEwIzqn+Mh+dXCDP5nv
ZjB7xZXv7cLlmyEoFTC+GTKIs+otECmZymucLmUf8IP7u20LB9PzyAd4u9UgKbAtwRCQmf29/zDl
/l0RuXX3QKxQLUtaNiVv/4wevenn55ndfvL/F27X8B2OhSyVfTM16KEPA9eBA0Mny7U0aLYjmtYU
i1nyJjv2fxyoej4OnYcp1EwE8+ufMUBabpAxlT5UVPVlQ160XIkXy2VpkWq4MT0a9HJaLoom1w4J
FIGXZctaEnsQ5d26O1MMcJNZKDQzz6mwMJzvdym3cKLqJ74g8/aqu3CLpPHerLbsP7/jmIr4kpLo
KaTfaaQ/Q1qS+/KNPG8zmyPJc03J0oFhjHXeukOUAPSY2uQQxQyMorKTkVedj1lKSetr6koRAZlS
AdhbDq2/L3Mx3OD9x9zJ2dW6cjAYyLJvtJl4ikgQvtZJmTGVUF3sFtkKKxmyc7RIHIBBShxjA28h
eUEEUs96vl5WIf4LrdmlE2HBkNXBTbc7NhbW2fVv4/GazHCZDLX6MFKQRL4Rs3t5uNYzhDM4ogD5
IN2jaelU2NNVFo7aOdqhkY5wBjSIxECOzE2h0BslJ5HTxTROdHR463TOfPC46fOBxXTrjAepPSTp
hrV2g71dZWT+pYSsQUkeD75HSJHWpX8S1YqCIToKT7KC1dDLyCUpWFznDpnHk/XDd/TPdc9qyK9d
1ri3RSVn75xCu1LRTFTXJZCU8H4AwL0HHNbWy+fEgG1LcLSq4vDIdrMqS6WcxlmfVy+l2eMuO5Wd
OiQMjyhMAN4p0oKBuaPn7Rh6pMA6DO17QatyhzcEuj3G8HKHOmS6GvhklXvjqVaFEdG/PRrjTU2/
EuydJ8niILHs9ABKbmL5MU+vbIsrkV3Kg7NxSsbIdQX4EKFyAQP+frv++2TB94Ldrblvvl1TU9ws
2zkVTS+gxL7yZNKlKZHovm73IhuDB9NY1gmV7bX6VVmAyHXUc/DjOSeUpcOAd2dPHX2hW63ePVmI
0f7R1YuCDtH7oTpOS/Iw8T9iuts93R3rPckgT/5euJk88YwY94S9U2RxzEhilsdMhW8UctdQxBOa
5A03ORXtIUX9EhV+RKElq776JlUDt0I1Yhq2KdI3ocEDaCv0gMeX7pPKlqUj5uR6wYlJ0I7/QQX2
U4lYYvuAZ9NcgcKK4CAWyalJcD1EBJ0fcmMLE6P3Ffhj86wESdx/nqsqbuRHDkd9+48NfrKDWf4o
OzluD712Lnea84SPrmRRGpakcBZK1bS4JZRZozaNr6QKZ1EB41hRkTskofPbVxC9EmGou5U4lSyD
9FJ0S/d91W1vh7pJAK2muFQ4iilKO/Z+V/yNYLLbrW/nKj+xvQkz2JUEy4blRg4d++Xx3bEE4MlB
G9ooRUHP+nRgJaGCEpdoK8gDG37I8oe1yHg1ZGgbze4M6qYAWxYUCe6toSZO7SYMKvIGkiXY/dBA
k+nrjXF5ZKyTGsfW22eEPivopEHujvhouEBkTAr7gwJN1RxjPTW4IIDN++1KZgbnBLaCq2tuKm0s
wDUHdO9LJxw3zvd4N64Q8ZrIJgkQDomZ2fLZFL5SmE4YAYZJ0uDsqlH8eKvZrACjjlZ67NvE+KEv
YuTTPlyYxFAa/UURaB/C7GIMhWF5/9jrLKM/EXS1LJPmUk8x3TY2DFrGid3sZss9i6ACMy4CoKM/
u+E+SdAbLyXtCxHjS8FMQJGwa2MQY7Y8DwAgtcm+/6w/meTpOhISJW7Mi5Wpzqb9xrHBZBHna+E4
MBlO//LVryDJZpzqnDrDijP4o8y1Kh6fNiqGV2ESLgb/RZCi8UPGLnAwhzfEp2kpkuESngNCstSs
9Cq90Dj1xd8FfOgiwob3kbN5vNioxMmyhgz8q6xGgjzc+lqVhblnbRDF6KAY6xK13Zwq80UIlbV6
kwQpxh61Gd79bD0eK26c87fiH1glW99knRGTKEU75ppURp5XO8jSqF9g3z03Y+MuUbs/Jmo5cqhU
gyWRQLJd5qxu4THW48ewzdKHiWGoEOzd7z1vsN9cvWUWHAZOC5YUZgrdXydYLTYExMOe+DJBWu/Y
YnOkjyJta8k4ouuruWkLPPsh7UZTEigdzjmIF1LTR96EX1btN6AHMBYyPs69P6esNNbseYnnogvR
95ZZHeaHQjHenJ53LA/FNw+x3c1lUeDL+mKWXJzR2uVRduDHomIXa4GkczHNGhKaXfURL/+2Kd+Y
pBv31EhtoI0PXeBmZg8JiOZXHbwtJ4hubaqpFIheGSOxNvCKMoX0UUcY9/vsKiTSWFr4qzlA61Z0
1vuyhz9xglpdYpdkxFt5mosvHhFzGmQsB85Z+5EaG8xWl4vs2sl7fF8wFY7QCeTjjWAgoofFuiqy
pNo0gWRDFuggep56cNWv59Uo1KK2SJYgy901RICjZ1pwSXHHrNs0hSM8KfuJ15AKuifEVy7CYmvM
SfAmKb4iOf0DQoBouVE5WYkj5aS3LTQGEh1Voe241mlWgDp9nSJDM/jvmsc8oZDzEsyvmVYkNc/u
DFA2sGNln+PX97hI6LmltI631Iyl2025KbHZABEbLrq9ITmc0uc8vUL5n90U2n+89FLodHJ6nlGf
flqj1bVv0IXj1JnGV8jRfIEcUleHWN0PBxTwGcKKPocvfpSg4xzy03N6/nzg2kzq1TFOlZAzaIAF
86CYbdDt8/wBNQCYFo3CGcpSk3BAZBaIzmBlnu9WMp/i1Qfe+LbruvZLG3ceDlg+MBhp4JQAgj1Z
QgcbXH6UwasXIWLPPRDC1T74Q4/ACzmRCPp2Sgdhh3txwMk/34ejA2KtVYr163h/z+Kq4kLDJtmU
ddJeHQOaYpjTjRfOi2oNZVPyW5kVT11q4m008Dt1gXdlkivGmqrL1VaSgxOdbk1RimllEcCtVSTT
ndMSjVKRMA8+rOWFsbNFht/fM8cf3MBI82mf/jdhAm2PrRzD1PZ0wljZdnufzRvmMGyLfhhfGJjK
Iz9ywJeYSLsUAc2J4w6s3BoxPL/lLXvrBz6xSG9sEpkfiER5DoLgVZrp65ud3fNQ5Ao4ov2NZKjN
/hIlLAGkL/8Qag6xpRSbKmUBJuO6vkgJ+F3fD3IbyNBZ92NaVOT7pknod3BhCG4F/JiFNGWOA1/f
uMlx6r0WEUckO4VSRjtQ644qGD4QwKw5oc37tr3YvVCrzbbQt2cAsVXLaVMy4aE5is+O772iFZKP
TNS+1EB+ZZsvb5X1YKSwqZngsbw20O8IjngB1o4BvXpSRFjLj2fyentQw094EtnwcGHTU9T241qO
SGI5KuQbW/zXvXAcjgG0namAO+gZfcFkOmwyol1TR7OOOtFWMhvuu1QAQnZcD6UUU4o1t/g4kLt2
FZLSYwo9ZobHRAJ5qS8OeGgLsq78BE3dxYWCpbEenFoLmBK/1/s2GKTuejinzD8IgWE9OdZfX19A
nyFznjG+5IYt/5iKBI+iMNuEPxkv0TM+nSGBe8GWcqj7kr3QEzhcg45bDKWCovC9wX3sBisKOn8h
11brXcKbtJjTL5hg09Mph02Lpyxd0oZJE9SfAJ3n08obTveFIUBA9EmVRshO0qWrV+DzsSpZN7cm
8wbGkAeloqBjioytk4TnHXF1u6MdcJk39273IAjMaRWXgmZHUsYyJLFaQQQMOgUJ43s7rqgjYReq
8vbrO5x9g4EDYycRJfBWGZr4xNmwFzheN9gSgLazJJfPZ8mCnYgI2OVnqCX9TkOs08Rd7DOJSWno
pyCGQdhAPoygumhkfDCQaOnPOj6f/HphKP01Uh9wHTjpfIn7bYxz+kEgUglbwWwgYpI1DORNZ5fP
GZDV8VL3Qrycl1mbDM12mvryE8BTxCUee0Wa/hF50e2RtW+S5M+3AUrIhiSH+S7t1QfAviDvc3CT
l+JE0qjRti7sTSyApHJK3c4sUJy0/ZpJvEEXA8uGzGV4jRm4hBo0/LX/g9pme3qM//7S/F7E+0fB
KkE08EFNIV4pw7V4G3Nbn03iMMgoRnGTPhC8M62AMyHJmlZ5MiYTb4aMf5VNfi1XzANJEbRmvuTE
3vClXOPHxdLhYykZk2mBqGbWFj8CKolE5WWYtOM1A01EVDlIhDuPggWL8m1CT3dPUtMbGLqIKihz
fQtqxpaoBPiMg1p+vFr8awRWSPGZLjN3BPLVXhzZxvKFz8nvJUkmbPYXelMd0HG1r/zxvfJMp2qO
ObDqHW9cu3xz39p/aJbdtWZCyDjuv/UAdhgDlN6WiBIsNkidM4K1TRf4EfV2MlQJe+kQqqfsdqHK
crQfElPeHFzVwEsWEthRjRIh7TI4nw7N7sBb2rDNQYWaruN9WcRhbCUWLCTZFPnf8NwrdX5sF4oB
8w8nxAPJJi2d/hhc6q4gPjtkK2r/3hMLlVXfzYqXTL2fmi7Dj3o7Oj2ZoqmHWMeB49mUE6StFIKA
iPMlQ+/pw5PktOk2EsR5XQdemNok/m7X4WAPsGYpBe2AFPpBIrKOdB5nR7YO/pBr/PzpXV3AjX1W
gA5tETLKm8FO1Z0q2VkLwZ9gxeCVZKb+Vy49fP41OBjymKVTGNlPxHAlxBWHQM0Oc8m4sDOQVI9T
aRbB0rnZfbqYJgTtEQ57xo82LCAGyQJDH+cFk2ts1qeBugUUdDsqAONtNIdBqhU5J+00xe646D9I
FFuUfhl7XVPngrjYL65Bj3BefvkBQqrxCbOD89Bdd4xWlO8xrv0p9FxP0hOlx1qs9JfQhMsc5cbY
G4U1rmJNIHrSvBx3Cy4H4IPPaZjf3ZdG2vfPRaShJwmk2+8nZsqlQbcnGu2ghPP2mK3qFdLGLL5o
fUVYrTs3EYjF1u/FTMXB31iOFyg1kwAhmf1Fbhg7rYOkd3l70kTzZoTDhKCEAdWl8GkxqoexbRbU
CFiNe11z0dBwpwFcuwSYJ2ywa+V6es3dl8RQyz7ly6TpIxPwvPDoJVwj9/tBI95lokfJM1SKyvdP
2mHWMPkR41secJwElLEQQzSyrzEvdRB2qhzF9Xz1D+nK9vfevYv0MI6ZGjRqEBfwce1ZprIr2gSD
aMex/SpXXQdkIYJqMQJvWw8Vc3UQ0aHVI5kSu6sHZEXwdRv6iRA/nY3lwORzjUfNUTWA1b6os0nv
TjUxxLj68WWMBpt5n/z8mta1/Fnc5PpyoyF8YKHw+PTZpJ4o9YJ/TkgMkZ/YyfmXZTEeViGS0vRa
FPRfVujo/XF8mDzTLQ3w0Y79AQF3thWv+VW7JN8xmI+UiUypGnouQWRpfTE7DT8Z+WgLxL6yIZ7M
ltoHW+gWUjILtB/YZNoeQSpXUhqgmo0JnY9qyi3bw+dB0nWSP161WKmLgS0xv+Py9x3ZOty7uqr/
jvvbv0bOUUqUp0TIk2OcZwQn6R5CrZnghwgfXikQxjw8zIJT2kvCNXEmpvuEFN9k1D+wQ9sfBqzo
ksSNqQ4T4KFPkdfStdIKLr4Uwb5Nfo/2okmpSRysXNeZZg0bwmQ/qQMaonc3mleMxGoAZ59l+3CE
ycQAxvXSGuyuT1ERs7y3hUH1DM3ihM6c59djpIqEmCmkvank7j4Heitp4qNOHhLdh6tit8M4vIIu
f/mBDUn123yJo5JbDPZlsbArvfdmVrkoTHiPdFwHAN8oG4Fd0+ocwTh4ml8fiPxwWOgKQCajD5i7
Ap6m7t0Mi/6fX3bJ2FZyS6Vh+kuy9byOdsmWEkkNlsI2wp4I2sq68+Nntb4ZRQY8YS3Nr7OTKBx8
Sk9BIqtFY1KDQp5nsLxn+p9PuEoabmwM2ED6x0PNRxejH8GReO93TOYJMfj6R+mBWotBEcL2oOFc
BVZlpVENaC9TKSggToC2LHQ5RdigTgbdhf+OT4mPFqcVsVFHORWlB1anL5EUD7XOGVgbyIrefkrg
mgz8dFdE2FUOCnRf4fBzuZPBJEI0B3ikzeT3g7gDy2hmWJxhzkUEflyYdtlqJ1GEorPXKMIWH+E0
AhyNDoHAptDcY1BZxXTvYSdALWJKbP59fcmczzbzaUiNX+LsZZmTUKRMhoyJyKrkEkG63JUJpzQ2
zaPGd9xm4Z0KWotbGh/1o5E3C369b3hxGca77vU6v1vSBF9mZDODfenHRHjgx7jGyKmsKK8iboel
6BMzdQKvEkRtT7NWR1P1OMjqMEHWILxY2q4nyW9cL57lwBfXkDQXcWbQCafHajUArg6DZWRv64Ku
MmZmk1gRAD85i41jCynl9vw2au4BcYuZVvKiyvLxqeY7/s4jO+CDktR2Qtn/6sp9bGntMUTF0E7j
UO+t1jeqErB2ikDUwnqKuAj2L0Yb6UsPsgXJwrFABWhsDMohGRPRLJXI2+ko+ixH0wQfFjG/aIZj
GUIm/FlMiLQdYxUjZnTNUUxHkA7am6x44I7Gxpoyc5Boctdq6P6QnzGjUxDc8qfi6Iwi5hm9ziJ0
deRSIxohsnqYyjAppCSUc/poWXbwz8Wk//9QrutRvnV4glPBU8ROe2NaZGSekz3MVKv6h6GtnoNt
5j7CGQNOGzy/V8+PwmvprE3FtHY/WmlqM/rGFt+L2cb/A0PjdJbZFVB7AtsFglxR3aY31v/xKPaK
HP3+/IISEhlGgiGnwvweYbQOrKKARgVhIC2Fx0VBCAebiDdMR3pLd/UJQCQmevlVT34IJN5/3lAK
JRHwuM083OLCQG95xEKRc17qlMlEeYYg/B95e/uoERByz43wrtxBjd9Y8kAYXWyPVP8CjxjcF5U5
AFLzTUoBpnFtYCJ7U1oVT5nZSNvyW+3NQrfoCaOdfxdMWuSZg29dS8rSh5EQ7nVP6Au0OGg3eoUF
bf+gCsW4tiNbJY1h4VASuoRxwaXI08309D36TgwKe8xESuPz5lq7i6Ch83+fQoioh7xJbPBYvTay
OrEHfT8pziLOuSlUIoClkw9nJAgoQH9sO7B9I6P6cRteM+fJRPBX6cRfO0NCA7dwI9dh7j5hudJg
FX5qk7Lj/feLtxHHVsP0jMxAa9ztCIwxeeDm+0XH82lB4N5dyTcESgX6bXEwgf18ieH0h9Pi/daa
x8k/LZ1LCJL4/tgm/IxsiKH/V2ed4kbbXVwA06ULzxu9ouiW+P1IAaWktSigdglmtVIi/kDsFCMQ
8Ey5/lUwYmPYW5bPgAQQUpKjqYpfLxsUlGMPcrZHrbnavk690XtwdzCSWimwoQ2AfTugnw5F1Rjj
KFT8Ts8PEMUon4Wh6cgq3lxaUAdWT6Vv6NYOX5MqR6KtN0AbYobsInR247vFpfxjrb9ExcCbJc0T
dycR5xe/KDczWhYEfh3arMtHPwEl5PyFt1TraefFgTujgjpBkxEE9WNDg109d3Ssrs87HYzM6bLo
OwuZoGQXTMukfCU1Jp+HwlCRGOWOQggpXi/4iR30V0zHkdivFV3qstlebCSxTPfjRegRJXc2D5x9
ijg9NwEZ95Nysv5cQqTKf7hcuLbJXNL0tT/VVRph4kl+2MhH4qoRe/YvUUi4/Nf3PIMN/qstwR/W
okT2paQ1QxeKdgZv7J+aR784DKNraDUB0uM0hp3AbJseLSuC9vVLPh95DjEsQ6wKmhi6aexgNb9g
I0JHJ2xRjttVfpNz4lRkRQaZPrSAckcS+jTdmFL+dsPuggjaXYLKT6h8+6I6wMmWYY+2zquGgIvc
E2OddG+K0zzfALmwzDZE48CpJBwVQpZx/pazXBCSRSozeo3atPwBxcZVMdQUDGhpozPYFWvqN8Jq
lCv4z6cxNDdaP/pwOlbssR53f+Qj7aV6otURrK0dbhd1SRPuFuqEZ0uBOLTvGJhfoQzmuClZ9ngI
O/IL9WxHPPr1LN48ui01HN7uMuTuQauWHWANrxEC5Jy1IegqDYOYH5I19sXb6pbkRc8gdecIbfq3
FbFcF8iLrCXp2SZbLRBXxtG0j9eBbnLRk1tjutinDR4+vbfhNbp/WC4d/77hCCBYwMd/fwhxMJqA
ju7So/9Dd/rnK2QEur2JcgWelcni8p9e36/0wteqqBCVWQrRfe8q5sx9agpr4VeFqQr29Xtw4aAd
vKEJyZe+026M27EQtlRB/9nWquLsUbURqUK6glXzONSP4DQg5/N7lZOXN1Hwh/R9tSyOSa58r8fF
IKwC1Y2AYqzjCQvbRBZb7aqczRzV2MFNtWUzjVEOpRmXjAsYyosRL4813lUamHRPEnZDQpeSqDa/
JHXAnUhOyKqTxUm7ShtKzyxGEi1jwzwpKgOztr94gKe2WYS1Efm4iZV+EHLco0fJ/nq7eZlWh5pb
THW3Nu3VttTBxaitJa16TXaKDy9OjYj9xju6KJYxbWOO3jlC+a8A/uz0ID1DUqjroxzDk3mtEbCU
PW/fyXf6Sj9qhmcnNwbijimzun8NThHPdUD1SA/FsoSIdoR8gSWSL6jE5QF3yLPBd44Wt05eWbgP
A5+nWliIYRUpEN++pNBh9xxO/fUFmF+idsREBfQbJXnByzPVr6n0NxqPqBamNNhDdnmrSCkPYMCt
qAODgTCHGV7KFANWCFuDxgXoY6DXynT2ZdC8V7L6GCCzzDWM7lMTynMq4zK9/jneBnXhWfjRw6HK
vOicM4hTFcbU7RrmdtkoibJTverUxPdHUd8CSvPQtEbCBZU3BMYjXh1qwILnN2Dd2r1t7vCbnxfK
Qar33cxhGjezdM8aJvI784zLN++MJ7Wk24/cTKyLYZX0MnFKvK738sulntWwSjzEVanLsH0TAkZd
/Vq8ua04xn1njYHW5wrII6PLjXX5ium9wtYAx2ijEqWFWX4HRy3rCtpZzxISuVZv75TEcfju0Uje
ZSGvrFYtmC2DXk6x8gMjigKM4SsN68NFt/ezdFKHmvESEn5UAZx3f4WdqdvTvcDqiI6HkXxujqBK
3LAn9iVj8TNKF2FqhlQ+Nk0k9hHcz6DZMIWquho4GIMOZ0iChjPldzgLuvYyBgPTvL2h6lFtmXVM
cgeuAGHdFrHOYa3XHIsJRFcZG/B3Jvxzj1YNTDTTPKyXqUDgY22EJ/8o8cpdTlT8uM0UWpqxdAko
NEWkCU3YGRJlfon556UvOAV3ep3delg8/xWdxMHcmwzyZ8F3BmS8cuTyWiTMbYmLZubiu3EPtHbQ
Q3Coq1eTA2HGU8cDAd80e4ru5KafYFlOh5TxuuhqqNFwW/ci6gtsFxDb3fGdv2n4VWD702KAEOBz
kDqsKptQ2dkwamfDz1TVpqhOnvi8hr83Jgm8nNKqn+9YrZMFZN6Tb+/jFceKtH1aLDu+bDYLQnv2
Ebb7OGHAaClhFJGPmtD99pNoAPP/NbzNmu3gKlAEN+Owr1JiwycuWOnsrbbqNgYhHsOkiADzX0+y
qpt2D8AzBdCKYkRtUAMOBdVSI5mtaH9qw5pnyK+EW3kpgkaTALN912YNWU9rupOj98npaN9Ij8M3
h4HItN32m32jFZjnsr1+9ZDiwJzCSAjbBpJ2d90Lr5KxNMi2t6OkWW8JGxL2SPm1z6G3qKQS+XsG
a3ThPauHTSRt2FH+rI4/wt5JE/tdhuhEClG3ne8/YN+v7aoH35erbzhr8R5wpdeKGHanozmaDy8G
JeNL2U8EmUMGOvrwjBb0zMb4NI+oBEhEwKinyEA12M4bLC2odshx6vCQ5p1Dpch6weiOMeaSuIT9
pv9oYNa+BI7/LNhAoi4bAv1qkLx8iiCru0UqCXdqint+ylLUZHxZ7yI+VGGmA6RXeSgSnbRKpe4w
P5J9uCWajEaXnWTA94s+yQN5xx8lpRy/ohsVF8OFgDpK3ODRi6PKsslux5C/87R5NlxenVRbJNJL
hwWv3F4bv7ihU9gdoPSCewVPSjPpQyxzXlEYOIkrfw+5lLT1A3mlzOhAq3qwbrQLPC6z0BNgJuAz
7XJv+eHKMwUKC33SIIb00k5WTNiS7ggAz8d+GVFJyVg13Wm0DI1OIQASNc7lc7aGaTXhKB94YDvB
rG7GJ4kMM9dSARVnjbkxwEENYfzUQU6xEjfyxarO8aDd3pgURkcRHFTqJGUtXAf7wicRczjLYdkI
CdLBHS4Xi7XHRR3iMjVfCkySvgI2eTH7/vySEA5BcTku1cNEibD6j9R2emos9u+LTLN92a7j18f6
3KfOxrWLsOtvEx+2MM6ePRcX0HiD1OXZuipPnK0J8o6BzkbstCxVUrRN396NbUOT24p9ikxFr1Uz
MEErK6AG1OSEC2HOhoBD6iizOgULnMY8gu80fiW4lw+kdCjVq4FscyrbWa9+2ONmb/KIWCjxoCUY
Aww7XdqEv0OftERw5x7ElRiu/9fx6Nef6pwmlLfB2j3zWu9Z1Wbe0y3tAWtmUvRPHVdTLE1QAaRA
IQRvSOcRNNH+XN7ooA0yIxKRvBqqKOh/KF2/mH/iqjWCo5cgTjbVfKVdTp+s/IPh17vZeYBUR/IA
fVpYU295AtwGK7zSOCfFtIS7NGo6ezNeNbHuoRanenaipeLLhh1tJ/pFrTE2JIuxWrnSf6OZ3Iye
DQZ8jBIfWRLBqJTAjfVzMtZF7yGPepT7gkV9cSAPEh5vA1uOiayUJ4bfiPjNsTLZ2//MO6/bwug6
W6pDh+CQnRpqU1IuJQuLgbcjk5/bWS45GBRGHvBKh5kRggCttmDkzKrG4oO19OQC8og3VxBk/ESJ
plTJxh8C/91irqE8XbMSEwBJL8UzD2Y7a4UvBB38jO8rp+ei6Qz0Y0Mq7xjC65UFyG39XO0YBlD6
B3eZEaCTuIUtomMYdPDahNBPaR/I1WAkXicl/y8L9/wvi8RcLBTiZmdxbHRbmED3LV/p4oEiW4ex
CFuRSmHcm2uuJnYvb6MpODg0xN9A1LW7FudNORkYltNfVZn2PkhK927R5Sa/TMJCGDFJiuS11Nie
DRpVJ9WcV0fz0M2M0+8C/ChdfS9kxaiDKBHrU3Rz4H3znARSlsNOjeVKV7lMf9b7dOABEkDtcP6F
t8QC+KRx+vlQXqODHPxd6z5K0X4MoNVDb8rreqnusC+p8zA0wF9bg8le2rKgf/ZOecnWCkQUfNOW
uzGtsxTLEE3inmTFxH6329gakhIZfZ4JbM0eZDju7pxmg78esChGjjuNLYASXZpBEOfn8dBDMPN4
Bs6JqHarBA9Bodh6V1oxMBMi8y0YYmfFVXDymLaPUVGwH3Eqc63G1mdi/i/qZnYu2BLBZ1Isx9sv
LgEas7aGM36eJoy2kJfALBc1a9hnZ7RATkFPosx+Vim1mkIRsyOvGMYu6rQV/ONlPGGw91GpEYAu
tWbnHlROC4rtEExPNhwgmubwmYqaWO3XgVj90IM0QwiBDnvDhUM7Mo7JVwVmIgIpQz/ljvt+L1y3
Qilj1s5cYuaA46dJsaJFs1/43qiYRBcG4wr4lCHZjmwqZKGWTg9QvJicwaogpz8vDd6WTAWaJffB
mBk4ViWZnOa4jGUTBR7evTBSgEPiyX7y1XlwtUvSt8hdZgyuhECfLeURaAPUhPioDlTsQM8uj61g
QVDHVdwpZXeEyvUYT1fCihAOHVHGyh/lCbzIW+K8fEtq5VCqG9xVzJU7LrwLcyKmO0AntxJ6mELe
BYK8JXEYIoQqkH9MIoqV5n/fvh67PzuXvhgj0NXq4X91/UFR91LZuBHJYX0hpZtGkApP+zbH9XXb
uRhuUWpWvskUcfAbSl9LtJ2kghK5UXg3kou6VdGfCwXJOBhhQB/iOByc68R4JYjk069FPj4n9z5U
gZDa4aB7rZow8WlhzETl6t+hpOodR0yu0BLfIsBnm36Uq1nJGJse9EFOIZGIer6kKksqosAygIGf
1oIgGS6RwhmpT3ckunoH25aOn6dG8Yswf/oIcKtHOAzMYxOjIztZXpcN3Y2Lty/SIxohjxNRGT/r
tFYlrtimJgt3oOFVED0ie5u6LwE+mw8E2Zh0hpJJ/FQPsNMCDCHn9SDtjYQMCuQ55BXYqlb2porf
ohHUrzJHRk+ol2R1hqwcMuDuUwV/n968TM8Ssd29tcZYpvB5m1++FfQPcgsGi6mVWHXa+9luKxEa
ok0bjidYw7A38XWYICHMoB2hs277PqwgBAa73i0BOuEqUKspiKEAMlp3bT91F5CEqM6Uu9eKpA91
xGgFChGl2ASEImQDaBtsZLk1QPX/azPZlrWNYZG8x7U1fEgU0k3gAYJEaPwrrO92bFwcEOdLkWIZ
GOB5j6DpO0WRqVyDc46UvG5AUtW0UL1qbJXuylQmvPHPiQEiwPu+hSOo/ZuOV1wdGteRhNLstk4E
k/5mmdxrSG6SKDMo587qwCno1qw0yW32Rkx2gltAs/lldDIFFnBfgz6DublHoyfbzOQxhLu3DzXh
Dq3QacQJ9eDr8Gk2KHUsfJL5Te62cO+wE+p0tPqnXwGQbVuqtkjYokmkUNAN7JgfkwiIDk1ZgpZZ
iho8mNButUWwyH/4LYvwIaRBQ7ThwhT1F/NT+zNPBXqxHEEb4LcyE9xSPvqehzL9S4+DQ8DMM/Ol
z2z++iW1uYtPeklC3CVSTQMJxeVlxzbftSC2tUgiH2/5FYytfb/+BXHPDO2mcQet1CpWaRBXQOod
N+7biUfG/BaOv5JZybT//kokB52MZoAX1M+DqAoTrfLkowlRtFNoKyaSSCpqRIXJYFl/PFxJy5ng
tOEJ8ZLtca8tRjOqn/kbQ6pyQFUflZD9UHq4u3F0kMHasxHH/UASCjkW4TDIfla/CTW9GaAGJery
yn3QTub76mke8TP2zTwYAPaND1sqeleoXQthnKgctugt7sQllRhr3LZykQdxYSbK0awaMl5VNLwD
WgSOo2NfvMciMK70oYZxUXSEdMHFxWY1s2sR4CsxLppsXek0DP/ABUJeouHL108V2KWIvrGX8k1H
/YZZg6JweLCD6QiPHKDEML7r9RTDEInHMDYrBLZGUv4rJc5HdBxkaQ0BrNS70PD0P7BjvR60yFRO
x+6P+/U2Mw4dC//GTXoqupi3V+jQuYVSI6/flmoocuLXLsOiUDJNBNYPMhlMTD3dtq/+iNwMtyXz
hKH0YTvOBsm9mPQqv2Ur6fty6woLJXXJWl2LKRKYrRlGqH7CXk9NJD/VpAiT1fEnbyWkAPcNindT
zGsl9AvLy6OptFoC9Tz5Za6CQNru6VLv8OmPcAPz/JoyLn49YnliL7r0H+uAQxukr9JwDzvw/O1X
A8u1brjU6+zbcxXN4I9g24W2IUdflUdljYnYgfybBsiPUUFlPlu6xrhS0QUh5+txVpS0M90IK/Il
Bwqqa3xLbcqFQOPviXWE9ZEDbodtJJUbKmmyfFHLmdzbIQcNywiFqrT36swhvIl37py7FBh8qj7H
aZHdVSant0WSlyJtLuKEGlgV9w1q1D22jHQMXgrcdv2C8RetI821RXjgi/a9te+Np2RsX1BI1lDO
P0P+t9Jo5e/tBe8Pg8MvaHjpMaqCdJnghVJPwqv3lqaTX3mZIWVuzXT4UcjpRLyUiIF8J6E4lrT1
33u7FlGlfkmX569EqrMf8ml11NQnAqX2jYFRtJW3zuSc7OWsPVCs60DMByF7MP/q3OVIMIWaaj3Y
zfyIyFFLD2VnofC+SdP8vPlHtKAklp4grzQH85h0R//g5yYjOH8fPrsvBamnrXgD5BvCSntN6Nl2
Pp6HTNSHElLBz/yKKWVL2CpXbtcLBEXeUGd08BDzXFtt9EmBl/TENfNlcuN+ElJlgW90y5ntA9mq
b1kAeullC1n6EmrGK7FvfOX01AldUNGis8bU1L5dGURsmCR6+ai7zbbcCQZbfZv4JIyKdrD/7z1W
9hPo00b/FV/kMbPMkt58B47kqIe3mL48qINFMhRWL/vBgcfJgj7LGocxPg9i25iPUTUJC0Z08KFa
G4yL+2NCSqpyOQiu592fPXHJBd4/4x8x1PYqo9ydmCogIJXFvbFq4sDCTYs1BL3Ow8hW6HuCjo57
J/4Xza3yaoTyQq8XwOIQq4myP8wnRnc+LHUO9Wk86YxvxXy1d0zuBjtuxQpnKRup6LAGsVS8XyzS
FEurqykU2NB22rUGKMX7XYw2RFJtIyzcdeY3kEOBO0f4M4CeEDeeCArGOmSUuIZjiM6nRsnm0wmK
irbHu4+1fjPlGpCVBJNR2U42q7b1HNiYxOpr78vuhzY0DVwVYUfNr2SDgRVEAGDBOvTCoTGJBQsa
QjPbXaCc1G7piJ90D9TkYnXBiy5BSz5y99MJmDQrHib42SEXv5yNwKxO/xSGMfrLM7oAg7FD45l8
vewAcGL1ts1cmJWLIXzfczIhtOeyjaVSyRKqMQSvEp25HX8B2XW4kKejHo1+j1UeWmcCyXRWqCv0
DgwSleoVqbrjTPHaT//kuxY1kDshP1+Udj7d03r5Bv21Zhf6+t7Yd2ncEWeWWj3ZRHenOm/2AXAF
tHZ5xUW51BlBbgmj/JcCIyS78lKoHIc/QYe2pT8+JHzukiWQub/qZreUJWHGnUivkE7slXLcx4HH
lx88D9AfJwyaK15iG+Sk3y6rKK/PvIhY18Z2JsMUGowuytw5uOkLcpU7JKRcf1/QOY53/OBhImic
PaI3+U6uYrOtW3M+V1qJMoNx2HrtfBS8Fgw8MzH3FV3TlOAnI8sTkBbbf/m6XTHQpPVTamZ78pyh
NFrcd2h+rFtyLORhcMjbPbjUGd4CYeu3GnxkwK/yDkYVLChLIEh6M+VyYa4OQF1wmoZh2XX5ACZk
EsNzNV9PBoWSTJHCsFlPvHnTU7al8ibhEnzvO8FvgM531XMM9Jr4bpiloVpuL+zX3+NlImj9ipuT
Ar1xYfbYL7XHO/jtir7sFUG2DrohaCZ4Ath/BJRKyWrKzmZQpTVRE/R9xyfd8bQR5h6kCdeiyXn4
cK46EXVGm0G+g5G/8LZEl9CmVddy5St8QiGmjZpdkyrr1YtDrKECzoYbndjPIC+8mRthPZpONUgS
OMN/lT1nvJyxxAbuYE6toF/tLENZMQvcFGGRrywnKL3Wkca+hX0HksYE5fdpps1czMMcEoBSSpBG
QDVq4WvMYGDORLs4hEVUgI2ImGejt1KB3hEhqZ86csYEfyG7qW/UyYE67k8BVlV0NMQxeF2aTsvv
Wb7AmLfdxX69q0By/n6eWPcCyY5YaZLEgGU42t2zeCRMJgb8ipMCpRVHTwKxnmSd5/HfgkfC+JI+
A6RaJWR+2XTICg7bUv+277egQoLJrM9P88agbi/88lLtp2mXNwp+efuv+RnpqYhVUbrydjSq/bdS
bKpuyPP4rehUjVbTA/WMYLhJ3HRzwmWRWGiPFzm9T3ofOJnsxXf6NqpMU8gnVgmOjuYlIqYBmJZL
xsepYX8X4lPRE9MJPgI0nfRVwRyVBVf7/dYGXCVtvVqv/3bOhZKir+NWRLmQ2jIloXhmzmQgDhA0
hR2u3BrxmQcreblUoDnfQXJSm7XJF2p5+mO5XFQacuuAxtBJPl2O5muUVWfQXPN+iBbm44b3gS9n
ZWZpV2/v94JRsayEK+bCvY+E9/FwIPA9ezzR7KLTpcXdTPY1qfHQ9QllmMX/16Zks84pTKJM1b2v
HBptpGfkrywZbhnPkYtY23jeqRSexQoutUxbhpkXEK81E06lrh4FemiRbdFybCzoyh7lme0oTard
S6XI3oCfrfAzqpGQd9egCchyWE55aWPQpkQJNTy/W+NzzXzXUcHH893LJM+BBw70RE7fRUykOoxd
YfXKEylhoGjINwDpAxm5YJ9RVac9cESgIZg84YR1cXlGOxJqbi2MPcI41EZr2fa+KVLNLnfOHJ2D
SM6jjCSXHL7D+fU7iQnnuupD5ZC8qKy5laJVwra3WZW7hos9PKi0wznJYXOLfBkOM8TfvMtxEkfV
hpO1yKqwXeJTQqWjJ0fMCMpHyRYtH6vH7z0G0tQ5bJZupkjcnSrEx588ZWg0MVXanOLLACbk6IOj
GMdGAk8dDJRWK/9+1jZDsQ4G0uoUyzMvQ3bWN0gGddQh5/6mOrTNaEsfWyCTbl6gOGVsFa9hRk8N
w7JPXG9gcxX8FCu7bADanEs3BeZKh2VCHp3f5Xlu4C/F5Q6mwmkLxiOhVoBcgxvs/8PAstOfYYm6
QJsrLLybSw3PV8fVJHn8+eHhM2A19S4fHglBLxx1TtzO/w/+i1Mz/uWaDTodwApUed1kM1wWkq5+
EXQwRVKbk6MYcFyD0b6Y6bGnenqdvQtN/hUrZsBHCdZzqMNLiuBCu3wcqDZv/89rO2Fdf8Sd0LoM
cL6HuNflvh6871MiALr5Nt7KN+AuPm7sFvOX53rYN+4/hHC0trPjQm4b0i1xMLA0G82l/1loHXlm
nqaKziR9mVYTlj7dpu+0OQlbBGTgkrp9yWh7uiQdJuY1/pJmGg6JFDsat9an/2yn3+ZB0LHvzNs+
Nv/g4GciJYmXaz06f7j7D55StGLDOAARqDaBgdDWjX92SlH76mMbUMRu8do/ymP8tvVkyzSFSq+R
Kero/t7awemcIF2XJc4JGDDkGwKA0PyvTE69gnypZHz1tOfMmLu9JkvMrcaXdl5GYV9Q0iOIV0/D
9ifsryiey1x2X7I+yY/Zqbc8ggKRWDZMzzS02dY3ecAy2C/yD6v3TTuwW0fmAQ6mhZKJRZOfS0Ku
T1GV1ruvqgzjSYf9M1Rakmw1sd4r+zpp+sb6nhwqSvITWTrO6UYm7tcnLdAS4QlrvWlbcBu0Is0T
I+5RDtyW3Ab1xe/qsrBNV0ee3aH0tELPVANERbXmWmCaPCxrC8bRtWaufJLCq1lJ0hb6EFpG3a64
YVNnFFj6QV/zIyAXsa6dTjR/0RpZDJuErk+lFULSvCACuv+sT/VsdpNkVfENY8SK6SitfgPFEZFd
Ob9ALz8w/ajd5lKm9e/LxOHHVlkaVtbSZjwz66AZgdYsuSvLjYDR1p6KJavq130GChTRBAg+oHLi
Y7nRl5iggT1gw0XDwk7lH4U6XYyxuLdOL6sqTCl4V+nPs7WHpOGJkU33gtdd4eOtMx5u1LfkViRS
udvCYiJUjHhFTpxW7NUVjXSPqBA0TBxpljwrjNjW7/Bce9Q7bo4CJdEX4xG/aw/ATURAGjXeFgWg
8ERNnEHZj2PeOtLXEjRfYpTGL/2VbhDB2xb6LKm1xW9QgwCWm56l+AbZgi2OPdtzLw+wBtjWNIWk
xz0I1z3sk8/DurSTkteV5Moi3kOU1pmDOPeAWNRA8TTQzdfT1QHLQ0vAON22OZ5rVzZ3wdBMkyqw
sh0giCQsRBZuJcIuByp3/Jp424oA5XPcaUfCX8biS7y2R3bhm6s2sQlPezb5v3rpTz2P5OefjOlZ
5tLMpsvP8/7cce4xfv9q0zyzcSc/OLloz96lrKjCVYmrX5W7ZY3XuWnA43L6IIXWm0/KqUIPbasI
8nipj/bn/dYBukaHQ09OMwntU1ZnFjWvVPc2oFCnKUlx8qws5CjY2ywA1z1VVrSblErmUL3pw8qy
eUJXK7iE456PpGcDVG31+QUkmyrnOydmzF1aofWWUvqew3F7VPos+3IX+8RU/ZApvpOTPDaufIn+
ePNH44aJw+asfCQxufWxab7Kn8jEuuuQKY1L7UM1mGtW8Y4fYdT/FP/t424jmQVLl+TZR650onng
vtqTDIaA6+Bv5jKXYv/Dph1mh8CieF2LhYnIAkIt6em4w3DET0nc1aVdfqgNNPGTUM8/hYWcsrpr
SJ1V9Bf0ovt+vJVs7pzH2dH4svFfMHmcYU5omUJTACLZA/8Ku1+XMldY5YTt7mpQYsEyvR74bHCx
BK90ouoxrGuE3ozvr/k+8h+yzdm2y8agt4Ou8WzILUHah9w8Kq6RGCxy05qoXBgU9+eSugU37TR9
9JxYr1CDIDPiZVJOaH0cEDB3RAHUAPsiasK8Lk72rO0RSMmzrWDz1uRNT/xQYvPEH1NFKTzjifrY
gMqXLwuOwYKH5VTVE3ESbck0sAvqv52sbYNa7aAVBvl+eOJV9XQ0EJM3O4WAqArhA0OFrcfYIbJv
JmSOW6gV4x+u8bCiSsYUyqmssQt9h+YXtfoAtpOoLkITmMZnupZS6eFlZ+x3qAd0kcz5kI6Lq9qH
auRSOBuR5Nsao4S82bbQfASy0CcNqV+lJyIKACIQY/hx55nR1sE1UGODa/LukvY+dojE1m8Pz+cL
/IgfGXtXCIqegO+5iIUxmEh3l+vgeh3P/L81klIq22cIyC7YZHWb11rhSpQZVM94vxufZW+fWalx
vrU6242G2UxC4lDksRITaPTkpPIA49g2T7yLY1h0GzuRFiBwaAitp7W0TUhyT3oV4aTnXWKxrizx
0oE/MvEOsJwLlegtXyLjaBQerOy5EaxQmUMj6MZiUscxlGgOCJsbSeIdRGJzchx8Q6suuLc0OqW5
+ixj1FkCJVQEVnYSYVmMUKMkpqYG8stEdSKF4L1oIUb7bafFYrzGhqfQy9JPLJE4TnCvEF3bsMr4
QKoWLqh7f65wIJaNxGmc+peztJuX3SpmJa4p3YTYPRC4GfTp2Udg/2mrFiLc3S2BxY0oYS8nZJ4+
73ksr1N6cM2b3WY/BR5X6wzzCPjH/ucNRCVWJoou3IUfQKgnh/5rTg54QNGD5+1sWqJFhkotRPDp
aFbeZAwwZaeOSCo8byxbjS7bES3JuWwcErIPO6JK8I9GX51BsDBzNh0zkBscwpm2weVhv9kfOEzM
ptMbDtke6VuLw6VRX0BUDdZ591zsj9wYfxEvnB+4I/vfUq+KLCQ8b7wu+wzMiHB3qHYtaluPnton
85bQRgAXAbIk0H+SaGLcRSzoP6QZ7Mie1NgUO1lDr4p/9fha69IeNxY7CHOkI6sPeBHkX+QWw68r
9LUNQ86eWtlCPsfUbM26STls/1zFRViFJtXAMGeNuU8rAKTrXYVCN1uXjPw0s9qXsm7Adz210yhR
HeCO1AcsBRiuZlnEoHA6iOyZwlCl5DXnrOMcNnEXzGhzdSjWzSYMGbls1GIMMfDVIcWgqaSxJcS4
Pq/f1JFOEDO6V8+OWmB8V/T4s55XKTXyZSRMCpcsVmbWA7TbxUt/WVgk+fzkoisnCLxEL4OZGi/J
asue94DMWEH78ID+HEqVbSjPVh6ZL/AeqsRvjvMFXIG4/m9/3wl2fypqCXFoZqAO/3N+Uozq0oMd
4C6s/QBu5ecjJQDBLsCYdNnNiNNnqQgU0iD8bWjVwU6OSz5hjk1VrMxHetrIpAv1qtLc5mzqqtdD
piY1KDeqtiPbC9iuplyFxJbN+MscTT9HMgrLvcvIHL91EBZbNqfPrWDcNzNiRz9jejKbuyXdsnte
NhC30jPFfxIqFUKnrOOFukpXV7Jmga8cgbcLYAiNSA47vX/5zvuh+QU+MLACBefqRM7/gnVwa1WS
omVYrOf2Q1IarmJDJpEJ1hAvUfM/Ay5GLZz2RXwqXp6aMt9hrrZPhd/8v+NlSlZY/LRS2ALJGaS4
Jh86UD6g3HU/nkBnPQP4cRRFNG61Kk/KJQtiuvL81Y5RwvjSjKtdCakwOfCFp9oDDi8HGu85NqrY
1j1Yvfas+m6ZXkCoYH21Qqutbu1TmAgVChiOTk5XvAUIIc/aQmm44YUi1VHTn8+sk+v6Acg44twG
T9WlIla+FgrHlu9jRGMLXqIm2aLA3iFDSt0jHWX6cibN8Wd0qQVk8Sz6BWSOBsyOo+lY22uIslIq
ug/eF2UuQQmaLyBjtVdPoGRD+m1pXQ//XcIF7eNAHvbW2bdew9/Q4MZ1YXe4wWYmfk0NrGvpEyLJ
t833lzpMlURRKiReBFjpqh9AhwfHy7NOCPG+TRF6EnAahOTY5LZb+qrnU8FEksXyX2JYbUd44AQ+
bl5eFsrZPU/oltCjDXd0pUe3YhykhpVrE9FUyE+fW5gbPl5sx5kBYqxf3jeekybkhZmQTMHKdQSc
qcifr5OxWJ0hCDo462IYBedvcL0VDJod5ODgaVUhXa1HBbhchIFEV66/396YPaARg6M4qzYGmHLP
YPIQhqehXS7DXi+1Ws4JmhA6Ne5qnCmVuT4+WU0hjOE0IZr2m01wlpiFySZ/e/WMon5yHjMvTiD2
ZzH0jHSLJCMLLgCPqE3pJ3aKTEe0LduvKbNZ2uqnF1OEv7fhFTP4ZzfhCpz30D7QOoQHowKf5Q6X
ljYqxkVC8K3zY6WCBgfcELU1wFHn8PHM8I+/GjlQLlyep83mjEC2tunyK3GG1tb3Zo7uAKDr6PhH
hJbRS60BY4ujhdRLaGWOFOKCfUlsk2Q9KppCph/eOYljs7L6zS8x9mNXAP7rcalihsq4UUxGIxaL
q2oM00FNIc7s7zWK/Y56fwN+e7doQDIakWorlC5fgOLk7Gh+daKEyLaByB5SrLKcV4D2PuLH8THS
7JOx4XAkiG6vh4iyUnfd1xsmeqBl+l5NWB5l1IOaPD4qij5uxr43ZqJexmM8pSRUA7bCtQCuRDGp
rcWZY/Ne8+ody27d7hisS84REvCajC9+JLW3sj1InTv0b5PyH9kocX9cWqTNSHis/qmuy+OvuPgL
UggbFVEvy68gJNu1keBU1SwcnW4f7lE9r1GpxsHUBbFwbePpTzblEH3CfwL53kGcVpksB8MBCuOC
s9BNzVN73OpFl71KkJWSekwttpt3BluK+uyhKPwHxSTna0RA7ytve9j0LjIFNHJvHA1flNSCBskc
DZGjBdh1sL+aI9+TISlAq4rncxj6ZfdqDi3t9UX+tYEusiiHRTYdIrAPTaWWZdc1sh3VrpCjo/Xb
gUMyA+/3HzeDtm+BhrE8md7YvlN410JwEsh4l6hu5yqwtyQOf19QVOC/PZCA6UNXH88ygGLGM42m
XpfdaoyWnfvEd/6plKlKynaI718a2yvuEBq1viEgvQXZYTYtFEL6Oht5rPzIUhsPbWDdNGIJ/cAz
9VgZcajoAAhor9d/sjqrYvn0SNdDDTlyOg7eQOI/aAJ+ahgps6kIW9sX9nxbNUAeE5obemqN9ulM
1E3avXl1mD77xZR5fOMThMbmyNeJ3VfzQWNrAjYEH0og3LAwODywjyARInStVSp8RY/zxQm6YWaD
WSiodwPjC5u+MkDv1VUENQch+rWXcgJlKo9dYVmigNQqSz/IzVH8mjz1N514A1VKBekrfieAQvUA
99/tO7aOwzuv51K5axGuOTYTeti+vMC//HMCldXlUJu9DsFQsFpOqzrBcB9qixlhsSJlcIyh1AVB
c+5gQ+NEh3sqKaEasRN0IDqjK7BXq0E6BrzYvOh9ZiA7urGOG+YNxGwehixyYhZyfgUAJ4UrEQDa
ekYKzyvZnqYtiYnUNPo/HcJJi3Nk+l6nQN/LL0yfN+jLo+nbg8oo/lxPPz1KtjtILCHJzJ2O8TCG
oh0Yvn9a43Rn3Fz6Uabd0loeWTnDl4N80iTHRp6yJIqfnMrmuFiWx1f4T19gnSf/h16e/WwMh1kr
SadpPRnV9nbEST5FqHhiPaWyrqBj2TzKDnW3Mx5Ziwkcjr2IPVfeDJtTwUx/h+3QcSY2Ob2sIzpk
0bb/Lc28b0G8Adf43fyyffas6XVs7x6n9h4RgyL4iFsj7CneCTErN29GXTqkj4kCV8My+nTQtNT8
tXS02wq8B9T4tuDJ3FEiKUQVPtxntQVNZlb/JtG47pvi20mApSoTxrKQukx+lmL/MqSoZymrE3hf
FJpTLOPKBbYJLrDhYftuA0LTO5dnbVvDq19/qn6xGxLL+h7Uchewoz3M9oKa9wbngRCpgvVyb+3o
gjwNKjXAHXKtm/VZk/pBEKQ6RS2CTPHoW26xnGq8DuhLae1Ma0tpmLy3fSl2WY9Zk4wFQBjvgOfx
rnI5jW2eIlr8BWoGtKaxrKadR15CETOfBknHekUBHe4i0zBhHddJkxFeBqLrRju0rgOxDmr7F0RQ
ItzWAByVIF9vJlyZBZ31eqHGqkwaCGiRLSfI83we5YF3c5q0mv1mtNQFRgc7aFCWBKLwefHEAkmu
hu4quRL0ZUwDnfHCD0o/LIlnH2nzClXqSXT8MTr/UwzcOmhy7sXDrGyG/nLgDinNyF59SUNlyAFp
nDxQLSTU9I+FYCY3XAJCUiRvW5Ug4k1CZH762NkNOy3ayyOEHA27aDi+2GkmINE+4EqV7IfHVklu
8jmati3Hs6ekfXrj+cGbiGGYSj+evyKQyw9OOBLJIvMf/DeEFQZbkPJ8hJPCNsPLLP7CFbvGrECc
cLYxGrZrW1S3cBQNeqxDzJrwklNZ8takhhVulqlYXGERwWjPvxdW90H80O0tAjMwS/J4JeayMj8n
Cx+Fw1u/5qezJiAsvUGgkH8dPmSU0L1ucK2WbXU5Vr2QVc+3YOfJOD786Pwm7drfpydNkikYk5r4
Xh/YSN8tgrlXMAK8QVwl0JhV5nTP8FG5WPkRT8gVErEBTFvW6mNn5MQhqoRW1xCNdSKsErktZkqs
IgPjAyi0UFs6OtilB3/30hsit/Ia3/3WRxBrMMHw9AWrLDaBhbDfTbk4cOJPOAW3ijIzu6bThIvE
hP8nsbFw2K1MAGlMjB5Z+x3HRb0jv85crQgVee0Gy4AEFq7UfO5CNgCTcCVtwVuQhsaejcIFxbML
KHAFVPqqe0gI4MvhsEddpEwLae4lnswCEM9IuIAAyCOmaTaK4/leotYYN0r068HaQKgwVkgiLkdu
dXPWbD7tlImwL/sf+sI61LJcma8aF3v8/TOF0ZhskD+FeCKu4Jqp0s/iM0FxwYKI7Dp1fwG+54Ch
hxmOLHb1dFrWIPqrIkG7kWvQUZPjNhU2GFqhK/Q/8zqpxMsV2IlJH0DicFU/a/ymahKnmuWRMOj0
MoBxajiJkOHAw16XFX6YuKABdMJmwuEBd9B+fmPr7NfuFwsYX4qmZPb38vFxemZKmXrS8B4mbjXf
TJGdSfv8f+kTrshDLVLj2i3cU+l4phJ182tLcAwqXdsOe4aVMjurbDaRF0YRJchqjHmnW4rLXEs2
U66B5nurekMPhej+HgQQHEgswHWvPdVn9+oAR9JiJXb1cmAk5XB42bPe8Dmvy2tA165OCCYuYkY1
7eU9fIJeOnaQIjjtQSNFCJTZE95gbf8ezVYjVu/+H4yVt9IAYJNs2jyNuEuGrRMQh5Fl9cTr+wbr
F7K22t/m9jYge3UnfBhJYQ8OLeO23/DU17mZTsQALJ7VOZPWbcVBd6PmignHcbwl9KJvWxQcPElR
sjeFHtql4gmBPGhTRCwkGPfzPx9KbVwy/43OHlriP6xuPKTXwa72QVSBbI0jcFac9Ew00cqWGKTf
tCcUzArtN/QOyuP4qKfgMkUvm2CrZdW8yJnldtTkz0cpfliW91YL7ne6LqhjtbRXBXqmaJyV3YYH
NS5mtSpGAq5a1ZXWAqguouqZo8oZ6DNtg+rLtYJVGKzIanFl9Thb16giTukIfbrIXxT4s4OFgqJ8
bVPtkQ+GIYqjDx3+kgTQPLYQwcqHbj8z6VMW8xMLBk4B6AhdRxRgUeMML2amdQ689+5olhPh2yuQ
jy3nJ1cn3CC5Tx3+07KwqLcZCs/jjOOKTHgs9hN3OPEVazHdEZTPSIttMwyfgUD+f5i//eMYJXyf
MojaeQz+l0nqeS44EMxJxIR9b/oS48vcqjcBzA/9gejBwNPM6kkS3L5FjRLMdPU+GpvAd+1qfGWq
LoE03W/hMaAtB1NuRn3cRBr+GeuYaeQJgDnuaEhKrOtTxcQwqRcuCW2Fm+K2gdnwM4RZc/JnANN1
aQk5To2HTdoTZoNnLIXcCpiZQDOS7P/Dr+zjRk9RyJ9FmyoYlxoQSNQk4+EI4a5OF/ihim8ClZ/P
QaxSSWmOEVsg4I0UOaF8k3GPGVUGN77jLKe5UD5JTBfniuygLKP78Nkz4exsRRVe/gsj/R50UnMM
orIRwspwYQzsDJJUu/nLW0iYhX3kQHfild1yD1cNULzSoo22CqxqmThe0sE5yEWoHNCpX5PG5HPd
VWG4ICIeQwocN3TpULHuocT5akq6dNHrpjrhqSiaZNUpcP/kubmumGiljn2v8IzESNCKLiY0s1dH
rhjpxDmyzB1T9pYbe8SiPzOugWaCus2NAXvIYTPKwISIAusobKgKQiCvKPNbz5E5gAo2KwgxXOAi
ITip3hxc0r/J9XCi1w4/RmWwLJtcihO729oG/4W8u6KT1l2XIszHhJa3TNPA98fm3qLwPeW5/mU7
8Gd5JdXExUiwbk+52qXPVB/Z/hFDi1usPDIBONT7TP5AzPl2zdbKTZQFw4yJxqWdQPBekoxbLydT
T+Xh7tVCp6MZYADI/DKqWb7BbK4AZ/+vVFxHMAzfUXw2vT7PVRNxGbEI/GaYfAkWzXdQyO3L10JY
cIzXg75XU19m0ES3m0JD7lKOvlPiWcxG+XolyGjXnWDhxJDZkPyywCksf4rCjgwBDIJ/g/w60Cj1
rswM7sJPBi3Bw10dy0QyPQYjjX2sUfTjNFiQI0EXDU4AAo2n9YjjRawjhunJA5II3BPhsKot7c9l
AgZ6qGqPgGgILgiGvYM+tRgotU9SScDBF1giwMltaeVI6Jzy8aSAeXhMabyQcSWP9NRp1jo+2i+K
hbOjKQlyY+0Kr8rDswdk3+32LCo85Nqjthk8GQTO6FIE5OC78ajkHI5DZPpyCSk7C/yb7O3YZ+ol
E3fEDNutvINCMSPtHS2itMlXVQomjTJ05bCDEjP+6R646Au1+FQ73nmy+jdXmMwos3nIFf3bSE1h
/AzOy2OQ0PwiAzUpFmMvSpLMV+wW7jDgiqWKk9N+iHJhVD8GShNsNEDrHwTT6tDfyUL3o2cBsCEp
mTVCn5Jrsjgx8JRY9hHS68+//3be65CsPUVGyit1rqM1J6q23mYTpZCsOc8kUgs642Fiat4/Of+E
ZC0Erc9CEu7JF5zxffKb+OpxMJ1AjaRROSXoA4kSWEoCd3HbQ4DNViAurmCeqIlzoQgLtQoz0W6M
9UwFDNWp+BOuCuuKXxYWIVnMAFpNxB2scKC2Nj+UFN1Z738wlkxcDX6Ii/pK0p4HPJQboIOk4DZA
zulTwoLla+R/OW83kyelyU4jQbyP0firNilNL5dvOFOCZtGaB0DRLui9T8e0zO+ecrwAHzzIO35n
+B7832tZhmt3xTJ5deRPEwC0E931Ju81YSx7ZRQTilhH3dRrk78/y4dCFPQ2178VA5yXuc7cuxDf
a2M6wRTcSjJ4ZCRK9rjxPhYALCOrWwOjP8K0THCVFA1Lb8u7gVDkuFm/mjeY2VFjjn7sqqeju4bq
dG6nRDfKPAjfMU6+wFLrgY36+KKOx2q3r5wSS2TwY7sWnqpZf0qvZiOMmCFPyr19X8gbMiaD7JOb
NtOPMTkJ2lFz1gMjLERMf9UUUpWz4X92YzlYRBEbHwplstPsJ3LjHfEcSFMORyTE2tGdDqBAS6f/
BSVsE+pn4tVz1J1PCP60BsYrnXhRv5tm4QRhqqKJtaxNDpioxJANVRg55FZF+e08ljpQTjiQI8ur
rueZieQNzXUhXO1UxoIxiezRocg10GW5n2tcnfEyDyZGPWYkki7eWNg4TbSGTMJx/fJiy9l5WDdo
GxH2eLswV3J5SiLpfkE6gGbTL7EA/1yfao3YQRv/7HB+Yy/ieSaSnaxU9UCufgIYBpc9zg4c0MbZ
yux3JXDqBTEDKLrGUkyyZ5HkujSxi6bNIxktSbwplRwCMY1QDkOXVaED+Bb4W1++Ddn/jNp8bAC7
66ynvg7J9GBF1eP1mw21rfDlq/rdg6xblYR2YVr5x8If+MjW6259LtXr+kgUnkLKCNG6KqMnfgcR
M7/MxFEbcEXSnwnMEsjZAjTqUsB1rbD1H6qy38rNM/nWfgFxxCWc/uCg2ddl+KfD9mL+/BbYf6kh
yVH+3YuZskjxPkYzfsbaOlf6ngOIM5BXT10dY6RXFyF9ukMkQwTK2EN9wZ4qGfs08dEUnk1B2OGP
5ruluMYFVNF4Tg4rZbmdk9a1DeWs11CCyOZ/kQJBXZ40C6QNAGSWQjha9uSaHK1chpOrmqNcuHTX
eJQl/eiCt1vWYV9CBty47WmtvFPREVb0LWUefrWYTBKViOxvakzU8TEB6NxApwhjIP0rKziv+DkZ
TB4FD6VnxdF9j/0J7TdS5YeBdRZ9pFKYarPc8yrudhU0UJsfEgblUDBxSte4JDDGa0TufZLQdVRP
dIrUzVTD9KTMGHwczbVmDqe2WxENscpbqTSG91/iPfHX4ce9O1MOjJt7S+XZ80EvfiJyinfI4+kx
wajkQ1qLukHxzIojiwdM/exevdzsOyWT1uP0bFXYRhjO7RxV69URymT70QXBqD9Pdp158VW5z5cM
jmvPggcLVovuS5sE9xMUPz8XyYmwstooISsC6MygE1Dwr/XoH77RedlYELHQjydtDKw54mEJ+OS8
pnuolxuD/iObSn+qF+A2ESk2AX1UdheZ5hW+5KRurM/OJjQ8UlLjX143RcU+k7LouejYeqVkkGP1
QEawVeQuKhNOVL054PIrN5hp9VPmkoZvz2vH7QmgQ3jz2uB3csQ2fPCnQ6bxzGNp8zQ9hS3GzuM5
r8l5A8OGxdyrYNieWzCbRNu/xImnZHrRvTfICkxSw9Nzk+0zIPSTrrfop1zZJ65/B7TdpKgBI6vO
eYb4uEIJ+9BSoQ0rJuSlDuSz9DStcz0WJ8nceBGGIHFo2zBajqTwAIgXJ6KBCEy8Kp/uRVqyj03u
IDRgPyBK0fYBilVmuE0AwwhiRAfVLr4ntbGKz4G8yYCWVSWCfgDKHascrTWlFhd9FAwiN8CtY/Q3
lKdgWKcj7RBT1VDTnP0hsHK06U+XPkm9V1kUYzMW9gs7eKEciI4aUkZCg3wFMqku9AIPkLQg3/yJ
QvcbEU2R5WRcv3oi92/cG+Bu9GycjWW3U/sGEebTXcwwE0UnEKOHEVyQHudXANSU6Z9kWwy6AmDW
ydSp+4eje85TegZjjfqIA9hwCzfjM9wotomzlrSX1diY5T7u9kpYHUsHRFGxPARfscDoE43HESud
rLSbxhJ6jqgX69ck0uHAW6MdfRbhKdlPO8Sx/imfUo8G5O6cFosiCs/DJ4pj05rn1K2vMiR2WjIS
5rFQWjxrYS8wpLjko90Z977dUwWtGJ7+UfN4Ta881/+TEl4cMxTkxdwsMxS9cWFmuRo4thVNLwYl
afjz/nqEcIZLa6XulFSDJbDu0Yt/slo3YzsZpsSSoLdW4t92VspLwiUJpqqGnw0TyljtPJjDnXhq
0vsj3VDRmPK0WXZzr8ap80hM92lzIene24DC49MmDpmMp0kHP3Awvxrg7KCUt6low01V/ERMOdxY
+R7hiVEfTMxmNrRuU0BugIYecgDD6pOX7Pc2kzTSgheKfX90q1X7Jm4Q52xbtsQ5NUh6Jax0/nEk
0gfysW1NhUHdEOENq+QrjedkbTfdkaUa5dIMXp4QufMYSj5H5TgWaibQLkbuThIQMTCkNS05ORmk
hnRlXf4BtglnTUhlnugTZQfw+SABe7+WF0jbgsJ/0CF4ODqzVnz2PP3vKSNSTmirwOCclNjOG++5
uAjavM2W86JDm1fWeqKwJ7C+1jNAl/OSNMcscBLbH9RC10YEVawHSOevx6XL+0apF8QHFFUux/Nf
ByUS6c8++lyPM2rN5YAZYQCODveEBhgtt1MjGUBdH4bSUObnWr8K6sjBqTIzC/bkkPMtTwSG/gET
5pwDlSx8wpPPvaTJWrCqEThoW60dhU1Bdkdxz5S4ibhZ8aSfa9ezDwOpglo6AVMiRc1A8NIu6x0J
s2xtjj2m6yYB4QEq61bjLAudDeOIIlB7J6hMW3l/NIF6a08qSz2V3RJ0BXsPIVVa3zVV/4K+pIlD
SvIXMn5xmnVQkR4/RFwdxCn1xT01D0kGYEuWW6bXE3qP7cR0317Q7tGzT6s05zMcJr5Gj8QH91hM
Az9DnGuKBPY7sQ6tXPHzYJkew1o2f0mpzjVVrIFTSsqXoPTyV1NI9rXolFGD9VrpLGILUDVRux0s
aL2Buv1OzElluS/kawItJyowml4JSDCSsQqsmehvhNjYQmaRnsKVopfjhWu7XdOHbKBjjNc6rea8
iN8myQ6zYCx/My/8etQlMfLxpjeBQm58Bc1o9RdgGlwbktvXkGrAZqoFkFBd6muf879dUcsI1YgV
uyCSlDfOGyV2ZJqVpVn1R9aYU9iylxV19YZWZh8butLz45bMEatsSrghAUO9jBzUg7QPM076igeI
2wNkWZKaV7UI0yG0wymwWdhbxo4DHRTj9IKzQQ97hfz4bNpevC/OsUw4SVr8kro9rTUnW9fdw2gF
YVLYEVgmB7f2IZfqBmJkkQ69HgrDlF+V0uK3UndxsCOP/8oNiwRlDuze4KKeweqDRLEOfLujYnf1
v3dNA/Z7niCl7LDzO7CG5DVbgog58qmsWCkIt03IAeC3jVZRBpaRh0IDN/TT4AtN5IDIPl4qHWqV
GscjihuX/EGYnz9pCK2VLBinULOBGPJkhBevqIt1CfqMwQOi/t+Yz+wM9NDoNCyjO7kDHKhq6fr5
0BzxNaSDnT9IvyjmABTjJtdM8jhPUPOZlIrMqwEMyLyyJ362kDs2kTNapV7Ebckn0yUSttz9GAg9
I9E0ilPVyyxwP6GVKlFRlSK3VEoZLkIdLVz0F1BABrcSewa9w/ZCHxmLFycIfaOwSmgWdxFhnd0l
rXg29NBcIuzB5YbXr4VG/rYgddBmQgIqlv2SyCJV3eObzyUWe7fQmqaUIpZI8wkX3/1BurLuyQEv
kBrb5nDdN9wkEqP261Ggiqkt58XIEz5aHyRRa7GoLZXK8G8srzGWEDpWve2jARctufL2DNdAuIG4
RpfJKo51MQqXVF4WasgQJM0tlyZMV10dDwf2x+9enfEI7kenpF9r18RdKIO5ezQmTX4NK0wELeVg
cHHGgWrjMvTl0x0I3WkZTHOg2FlWnsps48IlriD+X4P8g8utL1RH0i6f0dMp403rkwJYPmEGQF7k
jx2O/vrTpP2Qix/Uayya71XF0oRg+h9doHutgV/7MSj8LoDNcU1ZXqQ+6Q1w/rW1HaWu/NIowneS
MARHYU7J0YkqfVgox2cFstNANCeC1C5jkZz9SJ6+c6zOfs1nhdXKW7OVNb09m4CDho8b4A/7LWAG
bpeKSVwuPgiNDFyFd8oWOLdmRYpnMtvy0NJ+rIXgxI0yGKetsWIshrZA39n1veZfNO+yzrleMlCW
idS9X+kcStB59Eew/cSHJunQxXUWZlX3sF0ImgoBeIbI+sKGq//gL7yTm8makVuWUe9CVE4NHPpg
D3s6Fy3oveIA4dXeZdDEjhvtqRQgisBYoAPdknFYvcbp1WSxLfGTkbfTn6l9j+MqAjUbCi+o5nbo
h8cWRFnnUV6+0GuikckpUwDgTg/UkJPX+NRgrkXiCitWm1D/aOnKjv3KerEuSaEkKI3BIya46Nw6
llD8J4iwoCVWnneXwote3lVdGfxBBlKIrbxMRF+BXUKTnrLlCN8PeYmRyDhFEFZ/VT+wojR6W5HE
tcZmG5mHflx8wFmLk2D8X8JBvTAicf+Jk5F60hV2A+YQFAHb/UdwexkTbBujGzNytvmmsseT6ga+
ZtxuaLGlVnxrIFyi1CeBZXai8qkHXahK7UThz5HxLs4JuSaGe9tQ13rYrLsiIrss16Wa5HJ+FfHV
yGzB6kPqKgAVgp5eZKtOmjN6TgRTTf0mOEzflbTGwQ4m+J0ljWOZFgRB+iUKjlwWU1AgrEZ1UUKr
5WbP1jEIOkkchwuEJMEHGyHiuXS/jI9KLHFRQe1LkD7VYOUDNqQb+0Zgdpuit9cYlC9CQqQOWpaS
gJUPiKudUOtjjrjpzc8VpuF9IyVkBKOrKEebPnUL2KqZO7AJQ+o9P2ynpKrFt9SNyHVurcH6Si+f
1VUa3R1vdPQR21Ksj1ZyynH5dTh0Jdnfj+WnYz0qm0MoYI03PceGLETQbf3963Qqu10DVYqR6yr0
qT4q9Ryt1hfkXqeu0lO908HdKEX+zVE3K7hJmpRvbsSqfB/PeIv52Rndi6oV1S4IZra22X5HjWjr
+UAPG9+Rna8jVOhAwSebz3bK9ctA2JcUrvIDBw+ic/LAC6fFKsVND5VAP+Go/Yicss7GsWCJ8pcl
6HfWLvNFhK95HcO1a+quCFTwHq7YhoCo6uKCfR3PXpzGsyDqCfSq1TBrMqFpUq4RudszYWJRb3dH
deBCy4JvTeqPHTPgvjITTza8aca0yLX2F94v9sBhpfqiDb8X09WqYa/fQ7FGb/rhvb+tfmE9dkeP
SK6n10/W6xvypqKjri+++OGuGkjn+Q/SV7UCgnkHruVDxRGnnt8l8DKJCXKp5/h0ryxrwlB1KzrL
ATEj81zSgO6uSkYToza6Ikb+DfmFGzcREXt/Iwcjy8zzYbqeDCzUyFp/4Yo0NnsWNqTVCD7j/Y/N
q/TJqSjOqUmQAo9CvyuwKHwsxkaSUv2Qjz2pqmAZn9qsPNG/LQFmRM1wlzmtXRMHuKWG49DtVT4u
4c0W2v5EZ+tXpJWHrVyI9Q8J33WWIOER6ye3pw3HwXA/D3XOiQ3R2wA3eRXFmrNvdywsooi6SAne
no4snXHMXe/Vd9QUkJaUe5/DH/aDb8HICBCydEDyHimxENVRTiM82na9Uon0l6PwT+WLrSHrrVpn
eSEcufO9Ivo8rMq+91DiKTpaigPYkOvBTWZweadpsKqBbNDwSb3oLzBUJZF6BSBLW8Ckgahc1nAJ
MOBGcOIWK/3voaAAWg4UC+vGOdH2empXK8gnoeomZPur4ZAHl77WbLBD3HQVKMKQYvqoJYgkGECF
Vn0VXhRteoxfZVnnzIW/IGsfZT/aIzZ/6RJWgwEyozhi9uOLN65RpM5ynXY/6Zm4tYJj3armr8+C
rL0oS/D1ETkFVZhfIW5yM0LZtVcNgwh+NzKpRPIrnvTKtJJO7m9LGoLcwoXl1uj4d7k+Lp4IGdmg
wfZHc3B4ThfxB/lcpX3QolsF4nS1ang0Iyd6S9wK5Osinup2OuCvXCHSLiiHQ119qGuK8JPBfVIL
q8VObR3FMCaruOmc5T3PCno6jlZpe8JN/ebucF4O8oDlIxkdzP6A/PgBmLYVFbwf8zd2bc1ZPpU/
2V5suSgOhp5P/Pzy/KHtlsBl2TucPQvzSHc0aV3pOMC9ASBQk5I+2nqtvV/VeRQt4+wXxFnO7rKE
jLMo+nIXQykU/S2HMSh/2s9vYLQEraXVKOJMEFVwFvN7/g5Yh3WiHkWWg0sUGqravEFc80rpxIM4
OaHrriooINiGbr5isxjsKZ/wKOlBjAeJUtP/KNHfLyfdhnHEWIR/+IyGSRvM42tUtTh8ipyUnhiJ
EaM5SnkrVZ3E7ybrTSjTeT8wuEZaJnuKEYYcU/8b58GjKKy8WNn5qhiVon4EgRKbGh/n2WZmPK2V
CM0MWz08nac4FX8eK/rVPEJvBlfL8GfIldRajlp7TwF7iePlyoFGR72yNclqMOOIQTibk3sj58YT
Aa5aGl8eBZjpOyl/OK+sSjWT8mBzyQnGJR0xeQc3FSR7NikV53wUvOKiCuaWvfWxEicJrn+pJAqY
zTomcECQJYDkW00KO6naxsJb96jW542SMMyBDXpeSHo+nbUe2y3n2EaUN/v1aB+XMs5tWzf3B7ST
5qCvTj4/R7qNObr8RwwjPGogfSlKS1WeltC018hcHPuSR1Eh62F0cbN1lkpTSN9DNK/9g3drxpmo
oU8nJ3JY1CbHdH0Pw3kizX9JORibZ13YNrOGVtcv09zNuPH3kDmDZwPsbKSZLlxa3yUhoRmIDDdW
UgXsUBavCbhc2LG1p9yy+XGkZF6L6rEhdp60xOSA5DpqQ0hIL1D4R9SIbQsGQsOVURfunjdeUzzh
kOMgLcaQdRi+oN9cRSZOWiTJOGpycTpjqQ/y7RiLfqiIWXCpF0lwWcPs4U5aiU9GO7/BnDE1dL6k
1kM8qYtTjYG/ndsn9E29SMAldxLXD/IbgK2gjD3U42bIMzau1BWi/GwwjOaEgz88nsRPQHZv8pZ8
MB0UDjObNqJWSqAQEe+1R6HmjHvu+P44ZheIIaYqO81DJXGRahTodgFXy0YLPKQw/hc2Kkmk93Zl
1LJ4d80a6LG/x6PGODgRQP3PbaS3+uLo1rhL9apTJh2k4cmcRhV2Rw4YEqSwjNcztnfxgJ0kYs1R
8kPMvE6Mj9NYlZgC82A5Jh5J6prf80ODfX1fyxxVy+TERHd375jD8KSoptumnMHJi3P21GCSAgj1
ivjhn2h5BNuy4uDow1MG1KNw68DHdbBTWd2PIBVi5rLwPRgJsXJz3CDOeXSdh6r/Yz48W/y+XZxf
g5vAAkAvqjwbhbisKlqQQyEkMwylxJnd+bTNmewe6VQj6PwR8m7m4Zn+fNktZdHsvQOM1r0jcuj9
y699Sk5GTbPL8dsf6FAZOiYbDwGllcqWpbrbSMnnJOUbC3jy42XtrECIct4SyaykiOCy1FLG+x8S
JQnQ6QHu62FxsuZMGR+Ozt+TCjAKSF5KDblnj76gMzoUf78Wwp6yp4382fYeC+PL5HBRGcBzSQnv
PuTVSKTVFIQwMCZEdD6UZ4LUQVBipx1C5p59VJrRlyAsb5h7xnFoE4MajbC82T82p5zkI9gQ22rB
/laghF35mWnTTeA2OffWiAOEi6fK5zssciAWAxob+4lvDT/Ss5h6SKAXcoJeQseodXBZaQev+kW+
lmmBInK2irFNDUTwSOiWeHzwvhaZnO4r2pWjDCMqsWdeVlC9qvJt4OtGddcJLD0JUQeZzNvuhDnd
G/FEpdgQ6g2cs/Bk2dx3mCvY7zgB+n3WT+d+HxLjMl20g/xFaGpfmZiGBBnyv28RRL6mJXSsQmq6
CtzR1BSQPZiBMEwuCyQ0LQZBnJKg3zEiDWDd3z6Mttk47vHdb1QYiOvHzpCfIX+RVVlRKou+0+9A
58VsiR8cZ1s7YKucSgC/jqZsylDphYQUBLL9QaU4YQJzrSY3zazUPb8l9X26juhtYldvh4x282Xr
4PxWFvlgu6zPZlhEVEQ6CIk8AdvIYAvoto9IZFxsTUzZbFrViCOMTns2p0GnmJsprPGa8DS9k/w1
gEsMrRyU95IE86g/TAxdnWOILA3RfZhsRzL/vawTXOA0iZWvViVz2FaOaeTCqGbBWOTxCaxgiI7F
ooPO7065WlFLj0UJ2joOFuOpx7LZ1Tpz31RBgQOttq+ZeuEcNrN/ldWGnjyoL3lkIU9ZH+LOHY50
TsL4a5Kf4aNQKpMA1Nj22tPNW+uC7MQszkN/TAt1a/qrdSQGuDsJ0AAiOlbxm9/ju3n9OXkiQuJ6
PRshmEySy+bqlZ0TEt1aDPh+Wdfe1EHAUujI3OOVtZiyjWKxI4iDtGExx4mFdqb+f85ttldQqT34
z7mqxBbWI0Ou+U8IEtGBdBXJLZTpQlcc2el2kvdcCFHn3c9l6FbNkeSksh14Iw1Ku1UHwkcTOBhY
iEPCHMozm9PtM21o8u1XNC4X24xAVzHjnV4wgSZEvyQm9fRl6hUkPZqzrXFZBFF4glMOap6W2Fd4
NgD/yLSY0Li1vzPppFA2MZSSDdaQr2aI7BQOAso/uiDCX0ytqpn28arV3/yMkbRrbn6/iSiMids3
2+8tqMxZBif4d76BpfI9vdNyCJ4ouNh+0Qk20y2Ssvg6G3HrZ3c4+DmrpHVAWZljNJPkRQPvrB2/
jmlMLvnmTriuiy/05CaVUfnKc1FGTUDb/juHFJQh+Mnl2A9ffUmOYABrh8KTZTbg8ibddNATmnsz
3PfLK5hmNF4hus5F3tWoFivVdARuFvJtqtWzEtiTA854KSgWxfcxqNpDDlG0aidmfI2vXGt8rt7H
jElzmtbYDnL1eW0ojqPMHLdOrI5ODDYtAyWcOn2eyQwmo6CTHSyRPHTlnPS7khntRWzpbdIcjEJk
RlLCArQCLdPLz1Yz/1VwbbVC2BzSy6YB+5r7eHdF9uLAzA7z6x4mGItQBn+0IvqMA3VRT9en29Fz
RtWt0IbSVbkIUL+hER7PIwUgIid7jTHft3cw+zQ7lwjrF7i6grOZMTsBChoYZlg/ovLzyUEv9QxM
LdiO3t28Ws0Na0afbGxYQfHGDpTJueAtyN2vx9y2KjkG27O3DSslhr6cD02x5GTtDpIrdIo4sxM3
cENB6K7b3kNDdVblOTTNrhT3FQvdDUFAlM09Xp+H8T77b3ZAf6w3JL8k6A1bdHe1qhq7b0gvB8MJ
OwMlv9d6m9rI7pa49M8ZvF6H/LSfld2wN4mc5k9xtZTQniAaix6uEw5KidNVoRmSzGSYXY1Ls2uR
7f+RwO/AArPEmXuQJSoS4HlujyEtCXPimZU7yR6w6tQXKOQyfO4KsQHOcsTC7zdj043UNyJpoGKO
vsbQEPaK8W8ow/BF5PcEbz2VnL5BawBz5PvNAQFlLseMT0fZ0obybMGXRq5ta/YTPA0nmlU7WKsJ
xzQUb2asj9vBGhZeELmj2NhdJ6Ldf9odmnvJF9+WGJzxTqL8DKa9mwiKQ6KpqcUgg7+fwMZ90cOI
boLNningn6hAukMwUWsgUbPVNrubHuwYNqLPv6Bk0vQ9msbbWBSr27B08kmoCeINw97VUQRjyeHM
0ZXyg7nS5ZVSFNaBGqiRCwJ0lz+iJwExwhqoo9FGx5hqpzCTW+AIvGLsrBi/a5eejx7bROggjGFc
Rwz0OoKfK+lFrbVjktRktuxH87S3Dp+fenDMR7QRMvL+tRZ4/ne6M1vRYRZM3wBMphW6AsaUsiE2
H7LH0BOvTzg29zQhn2xd+ewcaGQ2mLDAqDzCUrmBn+VcuLukf72wDP7WafdenywkovrOT2HFKynB
1k4C0dLtkV/pUX+fWLFdxQT4iFpvtGqlodVJMJCQopptDuCzb+jXRVAtL1AQQpaHiU8cqBo7ztJp
tCEjbz9MgqMD8NbJsOsO0h5Xk/JYdPMKttlnWwpBzEgvTAFbXVWvjSQiy0w1lNwf5UtxZEpBUZKE
Oj50pl/yp8os9epSGea1SUX5MBXuG9dgSFMoXLk0yTlJGdApGpfhdoZL2o1hXUKTpgJMwI/gIvEH
vYCVpo0nwZIQyc7S13gZeQFnulTysaRdPUgZUjmZ5oKM+jgPJss2mY4EQbMuRpabRtqFesLnZR4n
yAzf2MiYzoL4SWFE1OTvb+2/EDb54SUJ9h47WABzlEJ64O56UDJhESMUit/TSIWS7v0OjuhRiTIl
rFx+hCWX9rToqRivNZGWlXDX4r9TEaGYInp2n4s/DBlh5DLTZcdalSg3z43EXckWNuHOTIkLFoRd
fbdGdERutd3aonjD+YaF30B7y5Fk8J6HrOHXW0fWqDnQQGPVPC81jZGhCwrdl3SRtI4ADlEKP+MT
L/ud2VuPS/hzaYZJcny1WpUz5ubh6gMByJgyJ78u1UiYluq4r639EI+j/UWNdjgS9IovjB9PRAsA
y72es8wPqLJoQaJEMKsHy9/bk2fmx7Y/uq0eeU0A/G8Jfscbst4Q9Xmfh+LOdqc8cL4nA/zG8++M
xwoB5h5ywcNSyKvw1emQmi625bmA6/zea9DfqYQ0jbNL5Fe4TPZwZ9QQJU9/J2JjV0nEPqz9vuLG
i5eUVEu3QBcb4J5Slz/i2aoN13pnRVdc57MsR4yBOyI4g0fI9LGLC5xzCdWxrSgVZh7UnLapD7IL
fhqyhGDmvaALtNQxbz9v6RZs59eQNdLzkUy1SpD05Bvw+9gshZOUSXROyjazhcCeXt0UpO6kYTWj
YMl4YrQkxO0T/bOtSh4KmfzspcE71EOGH241aHgRfJorYD+hwVb3MoO8Emjo+h/QGSS0xvLX6jS4
UxKl5iyOeR2WeyTm3U28wtKKXPCK6pMTUxt7i+xoAH9Pgxict+7dAe05QfZls0y+zKZXxl9cN789
FvlDGZUSChDv4hueTB5H/w4fQJXKT6wOCwIQ39FkiGQ3XGWga1X4VdlVN2uWvSWa97kt/DoUCfon
qhgrRY9ti3sVDYLzCUuOXMo0mJIofJCzahQHVpT1butGyNtcnzsfK4/U17zayHQVoqo7gHiAu9b+
59FmVWombWBmBD6ntqyL6TCdCxF4C/7/mhorqRxWqtTrJ0QFH/5b98UQFqX7f35nv9wLEWcfPoLh
muIuD0IavLkNECfV/JjzRqvPvEAjrZNoMSA8WGRbvykMUUavRLS3D0YmAx4xXkqT/0cZgUEMziav
b5BHcd8ba8Z7eRMKMQnUlBQAKFD4Uvm8uomZKTJZ03Wg/jrQeTDvYvAbYD8Z175m4j4KFahSmX5a
rE1uMWWR5m2V+6h5O3ehoVMZP8N9zPBIBxetqQUmdivuD14yJEmzhATu3PCxnWqSOLvprA3UuHLQ
z16Yt6uQEabTXhMKdFd8XLTvklRkBHlWgTJhCAr4FCYVeh1bjI9A6uKaPiMNfBL0P+2Or5Ckmamx
rgbpqzvWlM/Z75g/c96/xm/lYvKRwtu006B2YVuqraCogYFkMPBKewYBjXPGMoh4IBxmcrVvhFuJ
U/JCoc8zTOXpHDa3dlXHUUxvHxe7rqdN41WV4tgHs/eyqAW+cH+Erst5/pxqnIH/xdl40Ji2x5ZA
Ek72yGjmdsd2untNoQ4UJ5BMmwdPrDwWsDSpqDGUOzbaAtNRqBRh6MjU8IQBfpwu9Nowus0Vu1R0
850gjwp371l9CaZJXmo/W5cU+a7k9dzy09zXeyRhD3/tT8PubbNn2bubg0gUBJ/CDZw19tO9LK2v
/CMwy1yX0f2PmwpqKtTgWIIt+Ft/CN4fdpvbxACHgeOLTbwRhfn5UzHmTSNbG1QaZOZtYg5NSzoD
jcMMV5WjTSKbxE/hUJZy8hBly3l8wxVgp2T1LJXYUnjOrOVGRqidIzgIpJNZ7xJsVMa+KdUjj/Ju
GBsalVzBFtg2LHPh04YFNWdAHH8aCbbP30eH5/QXGvLT8AJ9zeSR7qhmA8EnPVwTXxctXLwo04EA
ybiQ3Zt/0ng5dunIUJL/z1e+W07ykKVYr2Xia9DAbIq8q6/6WJfOd0wtJ90H9eAH9nKerg2u/8ET
BaslEAfhwgC3Pi94rSnf2j1pXqF+9tH5ovBwHurxi77s7idyf2s8xyT9I7rwYAB0+zJGUSBYptcu
6uWVevQxR4Bi0KwtRWXGcaKsoYtSz38H+NhOlpEDrMG7tE2seiH3+vSVkcKwEeOw5IUdN5qzOBIO
AYuwWX/povbeMOG00wFaS2PER0QFriOH6w1GdyxrKo8TB6aB7As8i69Te3y/gT2c9J7UAy9PO+/Q
dWFDzoYzO59v8Lrq/itbPTsgUqAy3avIhBE6RloD/bjRfKQbaR/qX6l02vwdc0R1gc5eTGO6YNAM
L9NyFyH2VStP6B4AK54wC03Du+lCPoumscRSSU5QSu4MBSMiDo6okNiYDkeuVxMwf//JDYaAB+uY
RpmGEf2q9Qe2QBaHtyr/WtrFXm0fpLR23Sfl2pv+yVyHCjpI7TrWTWt65pTCx1TcuHtthAYlvjsL
EoXObCEBuNJy4GUk1hTaev1RT615H5Hz+TPxIOAa5oLirIHuHAmuMJHDORhson4TF8fzhqRT0UIp
BOsrmXA6FA2rgVy+E3TsZm/c2Xuuvz8urTx7RFeGJPsja1R3fygYqHHhDqtrp9gRn/UayVmpSYHy
eDwD7TKwIkbue0e7bbuW+qnTJ1kymlztH0WXPK5S+JQ2Wc6ntoUTIUNA8uvoxmM0n72K3fmT3y16
I9yiczRbZ7dYJlHKLYf9Pe+B7Cy8PPTEqX8L02bUoEScWvF6wa89212FVxOUnle0Wsg/h4zSVIm2
T3mnLIEPGYuEzqexqTE2QkbJXvxCdytwPiRdfGeN8sdJ8+vmkpGYUFQQhgguJI1hPyAA8+U9jT43
Zz/AWEkhzWnK5KkbpNRP52Ubj5vkB8SGTvv5eL2FsiGsfjjV1l2BA61shO7KCbmGtrq9I1cxLJ2/
FRAb3gXfI68SW4hhWDB5mpdORjc6P2/0PwhJ7ardK5gbzsu/GodRgcPHUHqHrLKrdJEe500csB3Y
PbcVGDu63bEFZ2ZGDMotIBmSfIpIU+RlBmfOQbLzHQdEz3s7PEz+aemOTGuEUNjyPg4MkJo80fjr
eNvMYD8pE8Le1WxkD6EjzalYQ53kr7OserrSkOvK92VEB/SXo/VHVx7EM/vjhvbn6BaTaQzHFOLG
LyaeysqXmmWBv+0ZFi/5JvbxHtw+SNeD8jFUEDRWYzUldZgjp3NzrNMzZ1ZhyL0eHwff7kxYFNV+
BL3yKU+buvdplCL+0TykByzhwWIYs0MaFPwSCGRTd0OvnFEKyFe2nhwznOKeWccR/vFe0JBwrVZj
OT6e49SfBN3ma2GWYAVPQJzyRBDZGmgF88VYGU4yHrs/eQSnicLpFY/Qju2++Y+UtsUnPpz1Q9RU
wAngQ3K6WIzHqkGpVT+aesH77Z4NEjViEXSpwQCy2m/AG6qC6NRgw8FmGyfzaGYlrJ1cWbM6LxNB
gNeLTMfIut4mNz3fhqXjc/vGb6Bd/zzz8Ra1VavBwJMRK0kZL8cDXht1qROO0zh8/+d0+FxD/0CP
JDH5My8tZYuSRkc0FvoBlKJPzOjBVCYnXLViprDcDScK/gRkzlyg6LvTfo+64mLoBS3+x9iKQfQa
crcmrwuBU/1CSstV7497WXcGl5nPOSWzFNETmK8f92ZuPDQzcFovnHl8PBJ1Fs3hKGcsqVDs6OUe
9rs31xsl00NNK4lN0DtrAG1VQnLTEU13BCTf8XcN/1Q3h+cm0+Tksg41WNfPVEwa8oZ7VQ53uEgD
iyKe7l+HeCEZNmNCRvvBtoAHNw2iO3yImN0qG2TAtEC0VdhnBqG4SH9FDzRZysZMwFU45N2v1sIq
NsS4bDu1RhTWm637c5YfUgKuM7yAsl9Wvfe0Rbb1DTI/iwI5D6/BpXsAffJsMHYbbZTAnQa8hFkM
iDlj20rKyD+PUXcUo6dtHzbNC7pI6d5vncDA3SysO37Rjh6LQks0oSzr+DVPoQG2adQZ3LM2Sqpk
6qzEddPducKKS4ZyYquLSDb2KuDSfudWzxFox1ZTfksEwLha1IS+fPZzIIDbeLBjLDk8wjsb4x+8
q4Yz4FQL23FvzmQzr2aGNhkiC+1MNurd6BCGtF1nB8Du4wAzy4vrW5C1ukX71Xtuv8DjWZVxxQhK
GiP6eBQK7xF5+japFMaV8IJC09LDG1+YH0qlSg2Ob+9yae47QOmt5ePNrE3lLKC+IimfsO1C4B7n
s/P+cAB8xqaVWXfQzSZ1l3p9L1GoXUYk4L/rkEnaydBiQZsxUVcvuZpmngU2NnXvN6MHP0eFf3NG
Z/gVVJSeSKXuu/kdGDCIQzvKrSpkg0Fr7BqOU48olZUJvrnC4Gl5LJOAI1OJ6puIluN1+/0/C0F4
Gz+djSvgvxwZ9ZjKm5ZUNv9tXWTkJqUX1gfurgBGkJf0a4GFrZCZ1Bzt0tUSrUmoHfCtN9EGW7mc
726aZCeWUSyLpxW6p3NrogSX0hGBqQzeU9LPJtoM7k0H449ORS8O/t42Bu5yUKEk1LnOSTGPNrPV
Dn+YFgz2LjtzlnUufxWQ7hu8zQ0ioU/xYsdLBLzR+h6y7QCPDCx+/Q30SqUcXXEx1DS9m2xauAi9
MBSpi5wLnPUJI4nLlsAkBSJS7hh2KmWSvzcvpT6PLDe+zlrucmvfZyAFjhLKeiLuBxPQiecHWbjO
91GAOE5VQY4QXyleIvQCn2+tE4XLGq4+VrDXuB2G+yhcxeNb7dcBRtkQGJitxtyKSidUr+tbXAEy
0Ae+5LT1emK/m//dlcgBUCaILZgRv1sZZvyUjj+it+I4kZCY18u99chUxhRLJDYgvDTR6w86J173
/MZCefmOvELEW5DM2qZ1FQ4oipJV7oi2+CtxZo58cDN9ftk1yguhyVbREvvaeuxLmjvPiZ++fDiW
a8oCc1T2wdu/0CsaHparhHvOKiseaItfiwWKCXJCVhs4uGlLkA1X33FkSiEvvj6SHG7SzNvvmUaR
PBoA3LX1HqS5WUv+xMJH9eMenEV3zHIoyZf9p7Ojdr6Irhi5YuM6rZR38ApRG71e9Xq5j0mXbSyz
GQzJAlN+vYKwW8e/tVMlBwEPSAx4sNf+VXewyiFOMa7q9ZjQIJT2QTApbcAf1hg5uuB7aYZ+Ieez
Y4UYUOrQYXLfTnWOIDJCFRwVZ6RqFsSXFYLqqv/wENz3cxEsfWuHBM7ebBHX07Vi0yBRE8ix5xVQ
58Sbz/4F5srUAhB4df3usjxXXh2BmlMruHaRtr9MtEQ1MFsqRuI8kUollAfwwioWEwu8BdoXwHqb
HlZfQ/XDHoNNEVzcdgEpH9jWbFHURQFrysv7+hL02SI4808yifyr5MkzDJ39NwORnAh+HGzB0QuD
4qW66EUVgG/pdiV+JWg0Z9a/brIFH0rG0nHnSk1YTPi2e0k2+os7QOytUmeX0/rvk4nslMghD6X6
RtcbStth1pzZdu4qNTk4tNU4iyyNm0/7WK1pGTPtjgrZf7+kdncIqmPwQKjyaE0oiFo7ndAGQI8D
wYlMY8tAqqpXrp1rzO2tEeichXGwylf5WsJv16wFU/lJ5h+o5iKh7Rhsy9vMOGp9aexsphXcxCK/
qRA2EIByK7G8iAFNiJoS9MXEflf+jN5wypW3V0e0iFGVwkHKpHmzIljk6DZvKf/IHVYbL0GMEp5v
nmwr1XJMwMrJi+HuODcL1gdVbbZpK+M9YewB7GOaEJPu5DjmSVsapazVXuecSe3RSS5LMnXoSgpN
fl+3T7qvNNGnK0cge5vCOo1eReCtQwY37gbgEtCb4rgIGZhpYawy/WGtBjLzmdf/wDlgfRJ/q0G1
X1F3U3HQ/e/ubeiljWxX6JMMu1QgAZ/bOVYKVz4uF+Ur8JaON77kY020v3oLArZQ5P2+BdlyB9Pc
rTJ2GYNdSwO3G7w0GY2svsBqRnvPOrv/1I8P1h4zBMgiX1jn6jr1jur8FKNCpPh5mBSlFQi38Yvb
nxPS92ZjHWJO3q0ETvWtoDzxEOSjhCT+qo36o9n1sU/rSdbslJJ6cJ0fBoZWn6xCUKrtNNPByeZN
kD665WDAb+6GhTtUGgB+ZyudEGFNXRDTvrc4osRf9IdWkqlx73YLS5C+20+cN6TEIjjww/fh63sh
KlYMcZqx3Dw8lgJp/NhdYyWvwSQIod6XQC4kQc4MK4/iJkWSBlhMSTDsUQ0d9cDbLxD3JZ5/JhHx
duL77lwSNLzjQxscKgGL65QtLyDj9nKUVN7f52v0Xn3qllfs8PnH+pIocUgs8BZ+HMoAeXo9DHD+
sSepLZsER9dWxQbF4IB7pvxI08vw9+uURv8k8VKCzPqVwj0u2RMWcw/6gxW8aim/FS7PVlrC7IgZ
/TGBlk5noCcub2mIDkLkRdRipLdFhpr/940q7v6qh67nhFTP26gcFyunR+3eq/UO02l19L9+3Apr
ivHsjcebZQF6XYb0FeFvh6hH/Ay8mSpVCg8oO3p/JJ8dx81VLbCxIAXlJNMaEcO2Ke3xwxuU5a0Z
eF+EYFtSsFQAL9+TbqADSLSeN2o7uR546/vD+PHgmPf8hRlBMZOm4OCCvVmSr4xIwrnHGZ/Mkpvc
MpJXJvCgYklp4InuLFCAlVVFflNYpACXu+Y4AYI68ck/mmtJHAHilCzeLZQy6DR/S61Z6UrmqI1g
XHkJMyOC6zJq+P+6f4iYMISwg/lE93Y/C5UGCID4SKV7+zdYjXQRlAfCm4ITA12+YVzDQXnSTXsU
0trUTPutuo6Civi0b0ynRjAOY9ttCdZcSmSvHOUEMfLWsI8s0MlE4cd5t3RMdH0vTGG1DwYzhor0
jjpJXQPJ7k5+dQQhLTOTF+fZv+ODZ/kdZVh8sXUJQRFUGld1aMcVz0jxWn3li8O/YbFLH+idbF9K
tadgvS68LepN1WXWP3QqPyBgA8+D/3HBIlXJDzF7H4MSXVJFcWFvb7oB4tBtSXHJEcni6gHiaClP
KryEXXKQEFag0/IMtkDoK3IdBkYTPsqQrC4rzAoUv9LG5ebYv3J9fIMDYGm1MMLP34sA6x/UxHdp
pYdm4Dtaqx3SPA3MMBtJAr6OGc9JkFeDW1vQNOd41xUVNdN2+JDI94lBwfcjv8I18sF9TKNSknQt
MA7XT3VltDHI18QGNUSLbDPAtSd1OiB1TK1P/xR8A/wdD17F+Cpy+Fn3eZm/+rDzzI/JCouaFptT
o1/aEosAPKiILtyYTHwxfTcfGFNogB6jOibc3nc1JdH/kuBzsEJHfoeJjMnNuD3RAcThfQGZOcZE
UAgChjeZu+NZBXS2fpkkmdg9j7lZeKmBXeH0OoSjemMQ647IN4rT3JlzbI2sMDR03OPXOz04SpcA
TeMyp2Adg4TUPFjZGyTS0w+d3o/NL8p8bOZM4dHZHq1nMxpMVJNMZAOH1B9L/GrrQYqUQm+hkVDW
1XvKeYie+L5yv4u/R0qo2sdc7jlNG4iDawwBJCji4wJCCF9vsEewq6PgThfAi177xCHqCk2zXc03
Z09ldD9pI/OhQwuLDduor6eDKWmVldCLqfJkqXciPItr2JmO/2QMHt8AsDyEsb1b1k1WbgmmK8IK
7uP9hDTrw6TeuNsPzwMuVfUTtLnJuBySMQMCYEe8ZJ0dSSH5i6C1PUPKe480K1cEyS43Aau6P7EH
pat+EcJqDFKFe9/PHBMDCbF2iaJtBWlzlwq1J7Hb0GW9TtfwSekYABmMVwEJJcPsS+KIJnR5tGQA
+IpYNm/mcMcg7SMnLo3ReQtJ7TMH1YmBarTke6MU3fIxTm0a1P/MpTO78PGB4A7YXQA/qUbAmI+K
lz58lecoXpxHTGCxAdh4SefFT4qR80+v3dD1OvuxjeCbsfkiSzf/k4oFd+bY1BCgvdfwHlkduFL/
ymDDiazsPdUe5yidw7VrRRh8j63N3hlpcfCKTSqa7LQOzjVMlfv039oNguq3l7y1NqUL1Eg9D+Vq
eY4c23aqAGVZZ/eGkwj0PkyrtVe83TuFycHxVrlCqY+sYtODr4GhzmPht6QW72dVaF8J90HYBGAH
ausxYeU1yFkAUZr8gol72LEONwsfau7QW8sTRDdKkw1cKeW3BcT341N4G6mp6srxcSBlxUfsi/mg
R4a0htQbLcxbm0YlJduvOD/P13rLcIlFjnMZl9iXgiV6/ARMG17n92HHBOXBLXrLO3g0Ic83poFA
Dj4V12PiQrjPd3WxmkRWyfCrBNEroMtwRHRCvZLw4uFXuo0fwkfgu1jwk2h8DlKcVhnqSa7pkuUz
+5LO1q/9mpt0Y09AzpSwMKmA1BmdKgFUml17AUZASXN7F4Jvv6aEqG//l32d8y2tYWVKozdGr59Y
7ePN9xrnUPKbuDN9hmsVyq//cixJElSuPCjnNkyuiklhW4HCelH9SvXp56vcgQQE95RvwzMcmVLN
lHe0uHyK5UgX1sp4q00GUrf7GgWSXrgA0MqDnoefcemJofF4CcLijmdUmFdata/GBDpH2znsrat9
2oF/bevB5iE996jKeSTLTuRUi9RofcQsJ3QdUA3qid10+0P70h6azflYPMIC/cRWAexsRZHpreHi
fR7/5gF098UR6FRmxYr5WJYZBUIxyNZDaZqBadmVRnxDxRrs9BjjqxmZqLiOrQ4BlCmrqisDTcxy
Hzn678leOH2DRAxqFCXMCVWhG5DquFnQ538pxJ+gumE1eEsKNzAfoE55HdWzN32E6asmCU2lhDzl
rVHGX1shiLlLNEX4lXuarA3LAtJnafx5oGTjKEVzaKawsAXZ/4toUPaBq5r7vgUgIf2gh8fIo768
ScDUTKgqFBlSAqj47uY84ohiA3sPl8EgtcWdD6i3ig8XFTOHwwvAl2t/7qN7AzCs5LESnfYVfea9
ZQeAVpMNw86dKUfimWaOPg/+OFdag/ge22+Q6P8XuJW9kGthBJqdKtpyElwRNerc9ZhGXi3HBN9n
gjI/NYWcDyyaYHdRV4YAIzuTcuKYNtbSZrkBOv81puSko5Ur4NpL27FuZElpk7unE9ZJ1o3yyNPt
1ImznDYfOIfyTvz17N8c8E/20PKH574G0RxiGLJazFLOHoK/4niELKJrA9lyB+eirZxh8KoGfWqo
f00WnOGEsLBzucqaY8tHgxYj0eqSw3mlRQUhU9hMozKUGgj00lMeg02FSHXygPbcoNao3uHo/miy
2n8okCXBuRol2mLqttk3B+GhMqeCSZYNdXgQEoK1Vj4fDRyej71nADliIvpXd9t+TPN71/xiyy/L
qXrLy9MOvz97Mjtj79xp3vRhMYiFXR2VsJA1hnUUnef4oQ9GMHBQfwZB9QqNPRf6vd0vS0uOYXOg
Tgy2dNl80/ipMPd6itqvMIno6G2EpZj3CId6RLNE0n6rAteULB4ZrkqEwwuWJ4cq2P/87L0SK1QA
QCTUxk/L3V1YQeCCRDqbbier99aEhiZzTHIaIZW/9M0anjf4YbuG5Du9xeGs3as64Ilv3loCtrnF
CbuTuEeAtYuJMA13k6Pti7b58pU9AKNedqkHbYGz8SE0meV3RDNv4TZqiCeGI1LKM6E8xJ3QW9Zg
rQgdWyPbxE078zCIotks0Y9q8Vzz8rXz63pPkP1rAEd3zgmFYZO8xvG9r6AK2oEqCjx6JVknTeIl
OkWUPU54Bzu6kikW2OsI5awcX7Zz8rPIbX+2EJTCMvV+J2qhAH4A0v/95Pzt5LN805MlpjNNuhAX
duaN+tqSAcFK442NE4B4LKokvYDYVK6IoqEvOi6qwblY8yfKEKwYMxzBUew+9vZbq0jbBKjQXk68
Mukk0cM7Kc/3TCae/PHm5mMuE91cUIvjk4JYAiJY4j8Qjreidm6ov7oujbRfgUnNwc2gcqYx2q4N
pg9iKvRKW9fKXAPLooC644N4bXXDh1+SfSX7UFz+1wkmKtDe5WtNwYFedN91wXh43eQw02zAQMnW
3yOvVW2HtzpQH65fSsWqhJQt/+CaxI9QJwIIp5jB1n0mi/z7jxOvBGLZKlFqykCgkT5r+EGX1zO1
QMzEammo9wPsTcMw8+zHFckpXFx1Y72yL/P+SOtXCnLS1y8P9fPntseWHGFWpeQY332nolM8huQR
pkGC0TkQCKhgy1jq3MLivoez5lspRa5J7RmXL/XLTh8pHEb7hmhJPGmwr3+3x2ginttokZXTbGSw
2TZnexpzE0kOZg7eP9T+gCp/cH6BNabb7nHA9P0N7gTPuX9ASZ8uPf56qvuCSCKanSLdAzJtHneL
uYxK96Z4i7jV3S8zBdiqW7C3VTHt1c7m4jf7RsIjT2ztFJ6FKFwfrTDV3DXPiW4inae9w8QAi405
mkZwY2MkT1g/Szq5cjdYUmAVV3Mo/JY44N56qPnGJW7NAwh6cciG/EJ4E0BDzkKTZKTr+C07X4oN
7VSktg635+caUK9CEjGTuUvJT8DpQcOM4r3Nk96cLPfn2lUUlTDv9cYF3WL6JYEKe3L5uKMB/G01
5uTRHSwu2T0rmuWGNdpW2Fc9QKlm9A81M9FSclm7+FybwuTsRYsVR1Nlp9LVbFItV/HMs9sHSLZx
xF7hVFH7O3gqvxnFra/v+5hDsDCU01HXkkyXpr/0vWqdkozmv6M9VLMuVSrSFmHnbalMdtkX/+Rl
y+lLVrxBZbcQ1ZApCwtG7WHyAevsXFcmE3tZ+lhD3R8GjKT4eKYOHXWamslZbJs5sXYIDblGYm1C
06wt0chwHQdB9BgLd4J5yu4LNM/xzEpcTJKdS58Pkic/LmT4dRSWLKHLnVwGj9OG1jbhEgK/HLJ/
8IPjlBbohzAUhXIEP3MZhZCx4U1tuZ32o6qenLs7xU5liNeCMZdT9rkuG9fE1iMHj4wC4tNVOE7U
psSP4R55SweBJHl1QCkDK4YDwhLG3HK+7w7T7vN8yRvrY8U296DteMejmZJ9ophMmjv8fT26LrsW
ufMpfNDBJntMrwYBmQIfcLK2w2RxfCBl7kAEyyhGhEYqe0DrvjazIz4EV6eDLH91ZUy5gQ7Mo3SQ
DwnSY4FjKeA8ide2Vczkl5YFLhCFDlteD7z/s3vPXuq45wWgIQ2WqEXVtBIiHIWV/WovK/XAGmWL
mnL4ZvRM+ARIqRuRt8UfolZHJ4fXUg1qH6ffP+SDDzsH8GRdr7h6LpWhGNOf1dLAaVdQe2nnOC3p
+ksYorqxMM7kfhduCaM/CHVUqpKprGcX59Rlg4ATyNmi/GUXzb+yDMKmoBR0G4dTDPGaEy7SdKjI
QoCt2jXpvSk+AizHfZQqi4ADiExiB1FsWzpursVWsPwm1pGSvJofjAgssFpgdcZDR+I2Wm+/Id7S
87tbT4xsmH7AJmdPx+xu9vvx/RDnjojQAjJRJ12e/YgIAyNFahnt85kSeGe2A9HQxcBdNq5CVmA8
sRSpCa3IYFsaOyfDSWlglmiTT6l8a7xQAAMy8pR1E7tJLG/yCom/T1ccscBi8tSULxx8DyooOM3a
Mta8YxVbGsCgJxgX8z8OQ3IiIr91I3xkDt/OxIqosJlpIJsEas/wjDMNee2UlpSkcmoxKovADvlF
jAyOxeCpJ56/+fnltRMRd35qOhH4sRwmVWqaxC+x+Y97VFokpS8MNJ6A01jskEPHWn9wvH2i/pGF
2P4ZxbS7bfOkTpTb/Vx7purWRDCoIkMa2lVP4G4ALLFuQrtVxkp6w4NK5m/LpugSq1yggpFKewEi
R6xJ79Z35ibR2XTzWDPbm+L8SsL6dCrbeCKtHW0VkCgcH/I6M3y5hV2D96oUKhvbFdX1866Xuzdy
6ZfXfUE9lzIg7yHobhFVpgYbPxeYJdprDFTu06IHDFIzmoXaqEbHk6W6r1Jckksq+OiVDMZuA68A
KGqQgizKcRbXcOEbbke4zkzuSxhKaZUokUS0vln07kE8oK/WETg2fk9t7ti2sGVyrbLvHjjmQpYN
9oSEUeNUxR8dMn84YfesfhXSPZJlMaeMPz9SofiecGso+hzY3J6H9opP75sLQK+0X1dn+mCSbzkE
4fDCS05r3sxJw402Yl267hzAqyfU9qgrJoRkNQurZzE8iDX5UOuOJg40yAbK3RHnf90nkoG2SVhP
ik/0lsLAqx9rNDbfut4LEhrtKfgOEQOdxEKkA28uFQudFn8Nl4rK0NfBH37GdHUA8hbcp75yU0v5
+KLlmNBawYWqDMu3NXG8V4U0TvlKGpzGTUV3+PrdlTX2Za92hJ/CZyHg0erYLWnqBO7jccsdOYDd
bAornkerL0Sbi2KP8s3RxSu4ouELb9v9fIPvdQwrm1cLbKynwSbfnxIaRLCVg/0vLhmbE0zr3Vou
HA7A2if8WClck+4BLCkCf+/rdANM9Kh/i5rhIUzKFIqUL0omMBRz1Pml/6u+DgrnoF4hMZ6PFEEP
tL+0RYXRnK+AllIrAr4+Hk1EvGoUh3zwtxn/kk7MEaxd2LGyCpAu+CbtGPMVtrt3934N93LWXK26
lsGige8H7aMLKCos6eIgBT5p9DnxtNM7Z5jxwlXzIhFaltlhLe4mgBmWbOFaN5ifEolH5ycgEKrN
/ITkC1Cvqj0cC1+9w1+2dibARPZu2JY/UmJSv3eZVplnBg7bL/XlvvfN8e7U7MaRNOwXVvEUrIJX
ckW3eJwg886QzsCBxRNgdTEXuaNcCVvaSFJGk86en99NC1ZQYcwV5yDzgfdoLgmIanwGFbzBH9V9
d9SMInyaTNjK42BYP7uOW6JHGJw8zMgocDE28PZsogVrJhU0NwnpfgFRO4E3LUAqmiLGxvsEqquv
ZgwVC2EhepDpTHuKQKGayKpybl7db6JCPmp0JzFeaEbZjwQW/afKYqSf4eJwaej3GmiRsuPgAfwl
LqDhhWIBjzwQPYLXLQxhn23F2MMo3pykhoe9HWJHeEopZcMCOK5mp4aHpc/g9WLiI09YHTwgD4ZJ
VMHd9PRu/RqV+GhzKllKVmVSuQg5pbQRv2MzIxpU5Ana2jHGxfm+t/Aggyi9a8BCCiQwJsL2rZe9
8Gvl0CkXVBh+yu75X2h/deGpiUHivZr6xxkXr6j01+I8Hg79RDtGKeF4406YXclRrjhgbPhP9W9m
GnW8xIT5+9C+2xMkBIOq7YE731ldj0OoC6VojaaNaaGOaMNbumAkfEU8OGCbygTUed9ATbOCqUaH
rH+zaGiRB/Rsron1x2bxU+rY29X1dFnXfdMAmjX9Avni84FY9IlETko5M0TLPnG/7kxiM7+Bbb5Q
/EJo0Y3zM8sVR2kqXZTZ6ZLm73BkgYVsDtXlItpWWcC6Gwi2bfuMc/F6nR8dT9Rjm9ugAVJxT3MU
bUlbi+Fo5Qp+OKT8NyJ+ItEClk8xxnc2IaafGT6fQeUgMkK0S0rNtA7wdtCCq5ZK3/4fJXOCbNuh
4OEBNCPCWitbphBMHyjrlAVl9Uc3IJS9w2SPbkTckk3o3T1RGFt5ZTyI8jOIMFUFPoRTq7C4Nvcd
cONL9SGTqWNDEiy5YNUxLWKa8aO+bL+t3c++j3yghRUVeT1o8zfwtCV/vFK8DANXkIYA1EB0pcGq
Xl7SgtMZEZWgy9GmnYmwlGAFgO7m5QqblVlGDK9EZgRUJVOPJy5prXsHE8KPguITiCPzkd/Q8LLE
fer/HokiJUL4SMnivw2ZsyWm/6w4JBXIl+6Jo59itsXb1TmT07RNUfyUWtLiWEi+NJf5OH4yn+HC
5I+86eQMmrN9yAIYQK51bg4j7ue3+BiwRaAuX+nanpo9vHlQm45WZ6F3WrotzuP4Egr3MmuVvKk4
7rx5TmmRPiGaTrqKDM072PqsKJBHrM0NV1YdM4DmWn0+ut6tgDYpXIeLzHDoKG+XJXe+BzelmgxT
wc9pLnmYSnrd2f5Tv4LaT/z4f+wwhmsDg0oAGy8qsrKNen9LW91LP4vyzu5E0bnZYTfltvK8pqgP
o/ovJWiGl4+F5XhRUbPEdNmvAbYv4OKrfbL2B4AgRcP8U0rSBk4Uez5myZiZCi7QOGqJewEPo8Y1
t65WJbFz4wedLXpngos0XAKe+cIqyEDMOkpZ5z0yb7PeV7QHfAA1BI8g9ECM5irF9ThMYqMUSdJ0
zMxwYWC8dB7AEyczSixWZUcivrOl0HoYJfGTrQr/jXxCbaoG6hwtHq95jrK4+D2ycvDQanAZ1dRI
FtKljX9LjWBdZC0giQq+CwxhQV2EnWeTv7H3vXwkpI0tg66mysHOj9lBQj042msLQ71KuZXrdhaA
Exz1l/By+2MK9l+uYrIQxsltKehfrjhXtncaps3T+FXROFi6Oi9vIH34is7ZEuIEUgA6YBEdCPKr
Ws3cllEGpBp5aKxFcUO+hby7qI+dC16eoHkzLs5GXmzu2pmhhXBS90Z+fxNogt9+cwwsYfv697KE
sij32Za/DRfh400HNahoyT4cU8ItzJxGm/u69PTv9LIrv3IuO+hpy7nQyWNwE+wFIxnUQQGvRGNV
7kHoouoK06P9kov9zFfoH4Ps3RVIxqUiZQA+JCoLbVyPrIFWm17SeSSx5+YiALuMmjMcLElCm/XL
2v7FQNmHVsSRIZh/b93O0Wyzb4zLQ71tpCVscF4uWN8rTcpZO3KUhfK5L4m3LlsydPH5ue7svYuh
hw2FPSzRj5iixxfY9Xx1vr9UZiMvSva4ubjJHZjaThgyRojKGbzEobsmVR25lJseCizO7pCEKuAN
xit+LDv4dh3CpLKj9OV9BJ2WZGDbM1K1KgkCKR29flAZNVBEZcKCiYrMBOp+HDlE36PI05B2aeTC
2yAIY6kqg+klLZifKGS35QV2iHti/EF1z2EFfNUPfUq908RDajdxDn1vFNh7CQl16TFdwUhD1ECj
NGOa1zUHWk5+xjf5nSaCwC3C9KDdDtc59RwU67b3RaQ6wPbRySGYVYK8t1YC7EfGhLmwy+3TShya
WKGlEcB7BNsnRk4ryxUS4QZhXHU2J9bUj8bokoV6j1lru+Q9cprK0kzU1tLhSdyLyhf4+EBT8ndk
RaElSeV7QZJpiTI5bxYFIiSg376OQW5QFzN/7Zmqr185A6JxdrVrJM1izv17mTG4PMsU6yX8Oblm
H/EX1IytytUQLQWlXnpXRIU3MvkcaQakTwoi58ZZNkpDJwpfecl3THUChzoxSlT4+Wsr8Cm/sgJW
P1Pxpsa2s31yiyytX/k2DbfyCO8wmB7mq8xAAYcBeeR1HZuwzSc8GHRpfqq4BUekgYer0lT+nOLq
PgIWzE7Etn1s+6aDSP/F0ktGmgMrULR7IZGLFaKZXQ1ohHu+5XdIV4OjTnISboC01JajaY8VS6bv
ZUdGKkOZfch/onHI3aNz9/VBopsKXSkY3lwIXmgtJ4QsSYg5HQTjaQU62y3aX5qUxdthCkBNZmcD
2Pcchgu33KwZfJ9VHRL8qljn26TIjBJ5TUy2mtjHLrpKNK50Ek2GVpFVx0J61O6EOpggbLhGoqqt
E95Goq9ISj76JR9IIKvC1RKpgUkEB5XwqVtrXhQcUqofDkucwyH1HxP2PUoJvyI5e57cFyLLpZ+I
rGoYoSzJOq50BiIr1pMgIcgdRTW8BZhggv5SRjkFM7dHV9ttreHg+mExTxBpr68ymB3Q6N7KCo3X
xHsPh6cStKFJEs0OXx7BqjxRKMHWUSgkeiQelRv1JKQeK+z4ofvc9sxvsuJiUFDSVlQgs6Uei7sm
WSxv/zMUI3X7sshuTCO7hqXLxPtDcKocDfJOCPf5ORqdCFLhN/e0Nhf3R77esDRXuddaKgHORloV
pM6BSWa8zu2GIpeVcSZORpTH7l+h+klmnW0AcsMKmyyzcAPqLGtYsNV2Q0Nj3K/edD91c4qRpNnl
xZ3CxA4i4sAzg3J4xQmL2G700gn2fozKGDKoD2Nozedd0rix6dV1IhVoe1alpcAUsZux5NtO12sX
Rjt7VhFrfNHxqDAInVrVMvio/jba+DEiOmq2vB6y/DDYwAbpvnW4mNPTennFHzFPS2J+5yFk2Wpj
3I4wQ+K7ahzflPmNkGmqkVSLiW66O7H6/7k9K/gyaoZgM364ASDczoh/5UpWJklOMZCkATDSogRf
jRKFShv4gjvV3VOzq6/7PsrT+rebeWVzcjxp8T7Kye1soWw77XAgLYPoopBnQniOkFfq6lPnz1rj
Oah4ZjMRcHb42D88ItDN9UxnZUIytxoaZ32mYyxRyfbMiQgqxfk4MxzigLYIwl8pxvnLWK1UkmZ9
jbLztFOnuun+ig3S4WrLUiu3iCxeeVsVpVHhrkZhCo1GO7tBMeJ3oAbcHOSLJotNyAX4SaCcXzK9
FNfbXfoZkZ8IFBbgnOnJu4YqvkF9UEGlERnG2jzss6aH1+7A/frN0ML6KV1HtUI2ErPup9WE8zfR
abjLR/DRj2JLS7gaRVgQccf5Wq+uP+cDNhd5vix1PI/deG7dYPWL07GfToRWEsL/q8Rcu09cyBLw
GsTT1uDs8SqjLYhTmyv6utIC+MlsQVMAFqpNo76JmkvovzuBydKBd6yaSAUgGAjsiOsdmvkk4t4Q
W6tmUnPnGY1/EgRwX1AYKJnbmk9SsdWoPUX1Q/pOCz2kkLaIv1AdztwJ/m+WN2iNlV2xDIqrlUp5
KUFPmE85bpLJtNFD47UmAopyLnat37nyBwepu/k0zliU4AiUeUyPIIe7DAfeVvYTL9sNTl/FcSZX
YmZ2S/4mTLyER1VRSv72hpXgrNv82VjE0k5PEtjuAKT7psTfBeV06tiJYHLYv6dw6INwcBu1LnJf
5mePymV2hDYhFxkUZUtAkAEcG4z28Sg5CvvkuCzBZ6Hzze41q5nuLsiPmwOJMTi7G7DX0oMEY1tp
cTgetM22Y/NvTLIcWrfg9e1UAQilC4olETSMAc5SUjz4bfLjEAxzmIjerJuTLoiMf12r07d7bSbA
QVqpPfEdckGJdoh/F0s6fTR+/2+2SkSr5kNjrqIlJUCD+ezeOOzm/AyqC7s5BMA3GXIY1QEnpaal
u3iz3quvNF5vVUm01+9YGem/byfDmZVUMGy/N8XFowLSa2bFrMW+XSR4AXqP170OiTwVpCdcN6Zy
JfnFNxWy5B1Bw7Xt1cetXZa7OsLPBtIHu351rodTB7eyWxunr/wMkUD4PeoWr4pROJH8SJsMykKJ
297xbulMUESG1HYQj4pnV/bdvN1R9eCOBHLGWL4jEGB1CR5BIkVuc2lAdHd/4y3y45ufZ9rdVZqb
v8L3iFj1yaVC4oR8L3txHXbKYpw6A+gIxUJNuGVGOrcc0N9Jj1UxD0FKOhUQyf+6gS01UhzKO4mr
WhOZH1r+BzktcZdWY8S/MzzX2mUuZTKLwhjQLMR6vmRYOh6PgDz79RpTD3Cdzz94y8ZJyyJJEiHk
i5DxyKVm7VM7qU+SeRy8wAa3z/3bcXlsrjOcovOsQdr534tIXX2rg/peRaYl4Ld1XTOGk+UfJsww
QqJi/Lj45U06tahfURhdc/5dzaZ/MS6XMPzibJ2zSnkOfg7guhIuT07KvMPbrmEsbTTMGxjNrJ/Q
WlJkpqiPuoFrv2cJCWbli6s9PWAxRmW1HAejyZso9lRzBua84PPPABAEWLsSPTK3D8UgdS23DJmd
5C/mlsoWtK3hVd06O4yfMGrhkk7bHoss2TQgN2EVM4D3+8IxzGX0rad6EtvGki9ni6bfbtVkMweT
A1Vt2wNzKpChm0wPydlpRhSxP4M38ANZwvvh/M2QMa9egaSz6rPnM9in7xk99SfUW/K+BBrIt4eS
BrFu6X1uP0uPnsrdlCiE94Q6ev3dPOYAU/cNoly8pR63mFZ8HiXFJo3GJE8swwaHM88zRy+isOpN
xWCbk3odJ5vSjGeU5S9iV9UIIxii5GP9Gzc4mFvzUExjRCpeXZcObKDAl6xlupQtU/cx5REdI7XV
E8kkw9QQD08diqPzCcb0vYK95zC9cXSAWmXPVZRTOw2tDxO97aGgsSDHu7+0JrpN5wIuYJShIFXo
Ey/xUn1mBNcBVrvIaHZEGQWdYmncesBD9ispc5II7eeRLj+g57/fr2/GeEW4K3Us8DBtoYCdmEnS
5Ig8cAdlUVnZpofYwuZC8vo3mtwykoN89zOHLKkihEs1phB7w5VtjUo4vWWpQv6izOw62gaVSUNs
p070ATx9IT17tJUGOLjI+UMxRY2jXVSGwccOKkQDTFj7u7Iuw3kqvQPXdhGM8Cl++1JwJlOfwFlu
v6CtUut9IqHqQ6ouUVfAwH8zd3O0QgT8ugy9EzLA4Bn/60DItehUy8G3OUQLuGwo0R5w0a0zfFX5
/Int/U31JLDwIITQ4dZXPblz7IPzrBSaauums0y1VIJK23ULPFcdg6e43m6WD7P+SNYoNs6Vsqsz
Ef6HW1Alca7L8C8SPQiWkBtC6wV52i6hOzT8C5N+uIh4irxJxzL0fCkqp/EiocInDivNYHZ9a3fF
kBdk3V0hSwHm6AXFRolib9OYslxG1b/DoUPuvLYU1U9KhQ73jm94g57KHG3qH5zUcXGorR5JZ3jk
Ueyl5LCCgZB4jQiXzlPFnA1CJjGp9X3TdSIxyTrnwiG0BBLi3ocGbivD176+qJC7RxsSU8Dfhjji
d0hkE/zGsy5RMZdnWpcSRlYDPv6EJdf006bsCIm51/W1/l5w0jbtXiOsnjv0Q7pJMeDsnLgHF9ww
TmzMXMTZ1zk+ymJSKJdiY91/Ow61CKpcec/SG+LgV8o8j5a0YK8olO/tA0vum5lW6IdVKM8CEQ5J
8lyzcUki+6hjMFqNHhl7IyHKhVx8RlYl2JnVXRtxYsviRMp+yrPfWoZiduP8pLzwdNjgk8/wMFNY
7Y7gzspPI5a1ez2/zB8A5BbSIjiFuObRaRD1bn4L3JaCpUwzn2mo95U+uvWH/gaAP472xM2eTEGp
wc0Nli+IxDRW1jdH6TTtvQ96dAkJMMVsrvM46sdwUAZdjNiJ8qQVnuK9VwUT3PAG6pBIHrkGjAdm
F2fMa2/eoDhd2fuxNr1moewgww5evS+Ge2+BpNYw8XruPf8L/9NiG63zqqFeH4luZn6HLdULEPWi
Hl5mPBoXuwQ0lYLlRAaqWTxhO6YLxqUIy4RJz++dfSutZW4SsryeK5WXpmLykmPrkEtqe06AgCM9
DXRGPNUJkqzj7luLmBOSloAkGIPzu+l3inWP6Ows/77EShtJf3HsNk4tQ/yPRIix93GEPNBLQGlI
OU7jD915sZs+CvXr47P/ibJ7XSGhKd9vuY1yxFWw/VWYfjZNMipPpWTnZY9hPKrctzEt8YyjGlyM
yzjrQ7KJSRN9FxvXfJf8fJwn+6yleXpS4PaLVEja1fM7lT39FhcRMo1jquRRkDHvzi5cawZThIb8
m+gb72y0BkGuw9As8ZG4xHwdNvZGQ5C7VHt8nbb1dfNqmwY47/PeQXZdn+kgUSZQAEBdzNi5P85M
+G6OYSap5J4WPtw8F/TYbIbEJHBB/5z2T1SvMXZX6toNQOIKwHdHAzCzGSMejHXu5X7hMBX9BhjM
bCVvj64kkbArL8qLvgpAKB+sOLdHOIl6Ogf4YaPBW4xp7soOgxWUL32N8OepK0lXXvYS5ZT+eBI8
onW5dLBsf1n+xjmiM09rPFIwNJzPPJ8BfiagKGu5gMiQZpgjF3iH1/IPMs7VlH3Kg9efu0OqSawc
Otg2IFT6X9+NyibVtrM26P0Y5+KfHo+N5Vsf34MA7e7iTfc2aEAT6eXb6Tre+ujhpk9qNftqnjsb
TyXbyCNvKnRAOlwuagvzSWQaX6lIR+uIi2Gi8gGfHYsb0DwkX9SQgCqYkMY30etUVLgBKx34IdAV
5T0pQYHaAGaiRdtxWkZ3zfPVUtZUqjd+QPlrNbAeYLNFymvKpSaZMRV7jrn/dsAKGao0zuT5+U4i
Js67+hhj72D90LXBNaKhTpiLiPfa4WMcWlYoZtsc2yrNK4HUVKspNkl5AD45AW35yGndgyqhjU+i
qMmUmbfAmVN6aIzdWyFl8qbw/CLduUwS4Tv4vEIXcMTRiuOMgKFRdeRuK1rfWLBlu60Qo40n/ypv
siSIg1PWIezCVcC6xg2h02keT27IdBUUazX0qvApakM/52mhJN6iuz6xcPvS7TZ5d25Q3fzTFWqj
MmuqMIpp8m7y2dvTMZ7hpBUUGfnC6EKTy725TJPhQqIwEgGcQlYaBccMm9GmmdR4iuoWsadSu0QD
dp0oH0Bn1G7cdTcLmqQgS35A7K7+KWAsjdZTdj2fShYBzkq9/fyIE3Mds3Ax4XRFoTPWp+AFGK3n
yphkBB17inepPF9cRnNNddV+YEkSDHxG2UNHkCLQJQhjFQcrwi+3CBZyOqW53eJXvBzg3jmzgLqT
VDyMfb2Lo2/rXQ/QBZZr6Vv1HiEgTh3izmXrjBCLROs8PmrFSK5lbS0TRl8L+dnWH46TLCIIekl+
8ESl2hIao2j2J59TrZ7s09xNDl9n08rf/abrkNW80nWD/SmUATEGpzhcDJgZSt7tk1pEYu/UUWeL
2P85vt0wQCB/p49v5wzrpmoOj/Z5mOcmuG2AFOP9015pAmeY/ycgMJhM+qb5CIXsRBQ9e8aRh8Vh
+jVFaN2jfzjGNi3IyfQljdW8UB7OzMiDI4dDdkzTN4RAzWmIbpcqRlM6AwHVya3tM1GMEF39d83Z
/EV7HzP9ez7z3/mCOFO5UT9dJhWzFAhxSrlQcG7CcfeeKGcqN0r8PVFGAC2MdngOYYD086qvtUya
SbdkijIAe6UrTNweaZEjLs3n59+8umn0c6cM8zGX91DzS15mFpzCbcwF72sif3OqCgBNT4RATY7T
wXxTr3/3fkOLHgVnyxFx0mFL9Qxm1zmD+Ju9/KdKN4ZAvlv9ad59mZfOHO7FmHvTv5vk7IhtanGB
WIMIOO7sRsvLoIpzx5bbaI863aYhzGUwenjSMXcbgW4oG+x45DpLjb0npc4UB2i57hxxEXzlqYhZ
pbQpYz78TKWpuBfQSBy72nrsQHYmAySYs2WScrTqUEuLREmke0AdaXuXM+Fox9dWibzTmryd3E1V
Lv48bJ2fTxcKdPEHujMvp3eNdyzRHWRLOvIxFGvv3/YohCFwUMc/PpBwa6sRar1fgPQxtldBzT9t
liyvSTuYfjYwdxjWQs1uxLieJtsjm/QMQ/BtMH+Pmn4y9H6j8wCDSHc843CC/HJN78SC9b2Wr7bD
MHTtdmNxRfmhhElNOWP8pZd8qcEX7JfqBWSvC2HAuCZeDv20f21qc3m6jszihz4Ytb+BAqgKwlNO
ZgHs5/cm3/F7rpCh8Dr2KXNaAQUZBMpP2cFm0PRbzgGHRgQH+YWqhgGwA8xF10jiPnVxoddpOVCD
s0B+FP0FBLAgxhOFYjPy0yinKbEPjhZ0vX969TWVkTCMfLXIOeHJZdHqBae6D88yQFM4aOioTzYX
V45S50QRnkG+5Cm2Bjq3nyRh8jc2evwGg2+4LeDOz09qgZ0Xk+bBvu34YbF8Z+lwe1N8uJ1PZUuK
UC5HiVU8n8PDlpN9aogd5Fc7tAZWDw2Ov867ZdTY9t0+sLNUJkbhtSCBWFMk4hpAlocNBsSBTQkD
EDDpJDv1fxxTRk5RAbmgIBTOqqpzvmGVUBGf7zRIDZTSMyxgcflsdtMl+o/KXVVltX8fNWfoxnT+
PfvikaE2MjPsI7W/t3+d3O5v9CnoYPLm+q+3M3xjXO1D6R9s+hJEMYs1zN8uyGFKHbpd1pbuGz19
mNDJ4R6Szc+kKIv5jpiXE8ZyNpyYBJb2Uh6XhgoXWg4nCn15/81tGyKVCMO0Ir7pfQFQpNFMOso3
2PSmmOwdqCmb4/AlQUWnm7HeP1aY4/wDrRCB4S9XBXZKdwoD+V/iU2PRWy99qXzb2TtE/b164M7H
j8IMJQ2sykSGX5RsAKIrTdF6JfP3kky/3C0Klrd4LU8ybW3QgBNBz26Slf86j23DhSOQPaP8TZcD
c+8UaO22upTRjrjBondcMraZp8YSrj0ketn6hdBd8i1h3tYQDviUKoGF3jGMRVwKxKsv/nnQ4JmG
evGwSwO4nA2esVbS8EW12lJ89x7cfDJlw9jc4GBNpsn9p2rrNpyAJKARxoCdE+N1Z3TzmDQBITpP
US68V+7TGh4wbrMbvHrq1sAumQr1ZokPtmc0QEndbnl8xC71d1RyIpqv0Nt8PXN47rLnH6jfEhxK
PNaBJIZiCSY6hsIKGjy0Av9CCq3G5ib425hfRsNx/ourJ3yaufc3wvrowsKrjeeDPsm3FrPveSq6
Fphxc12r30DKfvfKldOULw48ENehOkcdrcmwgTCKZpO8oUZNSl3awZ7u0g6DHFYtKC1RVcI/oNfW
XjCqLnK1QD7zCFmrumJuAd0gU3E8v/w28fned/N3yfv84Ac7ALtAwosr4k9jjtY5/dK1PoP8tp0Y
mvSojfrVd3/kJX9JzmzSBAfBDKjPYCcNKiEqjX+mfEASxEq5whaOwBtXS+0RmE5I8dTU88FLsmAm
NUHMS89n/I0ZCFnXGPCIZWobDqqJKeVqIdqVB8Oy56R2oYHAx7oVe2BtqvncvNk8nWJceApdOXMX
qD2sBl5agh/UvN/q5ahG2z9wBoE+nJ4WG22CoJw3HHGFWs2L6vG9VWYTXs71cyoBKhe5LQCfGDYZ
f8jrTeeUyo757d9cj4gEaBqbgawbFM8HnfHmCHTDqeUvF5HDGLFO6YcBI+ncDoQv0CQwwZVlwQla
JHP3vNpcpr+V6LQhDJ6ZY5fbJV/lApDgOJeAkYjyTjt0gAkJ8uAvh14vNqxp7h5lJ9eI/z0sPJRw
LH+2bsKVju7ZVIOcPK3eVa4CJ9M0b9lrDQEfEDUffvYq9INaSZj3cf7bhYVtbG6ztTKF2gBC7KWP
9qq8ro+IVVfijigUorkENoP1krXj5oRgn6YWs+NnCyw+3v2IrD1zCEd1RYpvYwWpUm59M0ZmkBo4
vN/LGR5Uj5C+OTir6Q5IzuGpc87MRfwe0zI92Ja5Mu7paqQIJ76TXEnhs2DEGiKipIn/TN8OBJPG
4x/D40GIdOqNT/IKgkgScZDp0H1FG3FHDwuYDG9vP8h9n4vHu4cLjMkTwOskFQSqfZqBrdfi+gpS
SlAxzvC9X+8TEIf8i/jyHdL7KouPvheV2y3zUGQ9LvpJoMsgNV2iqgy0K5Xj4t7IAX/7o+cNbtty
Qyal3sEzCxcs394zBgZjRVHjMX78diPjKL8MpZvfHo8TiPKlEiseuX4aESWc+JA7WXWPhZtECX++
ofHyu0cod54V7pbPU9Vih6ea3UQETfnsbl3ym671nnMKMPq8KfA4ZXd1ooL3ZqggJ+D2fBLtRNBd
Sw9+h2To4cXthgXkq4r8gaQvgJbDf67MMDgZyI88s3wVt9aUdJOC5SFHrs8VIpA/FTsvXyt/lNFK
RDBznSaqMP9NtgTff5EmJsOrHN5EeutQjJWpi8kOvAcNvEQxgyDO/1GjIAQY/db5aI4oh3rRpwsR
0f+u6uNs2Ceiwe+X9LrmHGGWZIbyYqhApk+yDemQ4ZWw0Au/50IG6jNjHOni2Namr9rrXQX/0De9
8FGWOqC8T7dC0Yov1QwsUjot05ISeUKCSgtqqyU5aPHZ0kJxUvRPJXRRq9S7AnBS6d9sx2Y9AjBr
WopdGvxIJQOxgjMswB2suecIrzwR1ZQqQjmO9YZuhMb1fzVySRL33gHN5Ci09QvmYrpr/Uzel1MQ
xbiyPBLQIPvlZOe3G7FV1vB+12ea8vzKVJ1gveHjoiU33wyQgrWEmZlaH5BKRI5c6bIJMa0j+0wE
jAfscIUCQYxDLQxT+2rG6AzcQLc4n3bVePojfEa8AZAbHxdfuT/ulPTQ/9qVPnNtdNx0BaRRvm6u
pgVdliEbtoJNzscWcZOSnmJN4SCdaO4xWbBUXUPmeTb+rwX2QrYZhCNiq5I8/GRsyNmzNZfnVU03
uAknDb7SwXzxaYJMgkvE16KGqQVCMlquKYGFZwokLX7eAEH46cf9LbY+lx880OXMrUhXLug2kXK7
+Qd0gDGYsNfK6o81Xyhz+h/uJ1o68Rxjf95HcgGxm3GZ7b+aTUQ5bOZ3ihkBpcQ7lk6vchaYQvnb
DfEJUo25SGp16ogU1s6JNrkHWxiMHLtQwB00TI0C+I31D5GqiGEtISdpHxQoZuYk/lmHNi6zQI/g
wPwqddF/xRmVLLC9UuH3sNJSbW2NP0FEeH+AFUrozDI5NatbwMxO8F1HDaCiyqlrsiRLfoJcdYJ0
sDu7if1GUpeDMO/er+5xumRny866cGLBA4RDvClD5gGMe+/PegW+g0pRfMXEVb4XYTw9OjgGT3GA
SXaFO1iti+eEwrWs8IYNoBZyho+jjKxCiMmlSKIj8YFNvReMfYAYZJqCJuv0i4HLCZHQme5UzPO6
9KUD8OTJCuFHJQsSmehoZuLRGrCyrnAaYTMYsOleN+C+HkdqtWZYKuEEuvrwezMd4pZA2qKe+pYa
+tr80rbgkdoaUCmjiqWmcehazVfKhiFex4JBQ+rF2UqBtu2TqRNN2r5PQjpt9+GfXcYn3Ssm7DeV
ElI0yL+KhNTz+kSDxwiVOA4oQ732eXuhhwg22YIqNxkVlxf34o0gawyb0rr3/pe1i/ZZTZ4OoLb1
RYFMk0LEZPIXuYOuJPZh8lOw5gsOa5TatpLruM2d4Y2EEpjYPErpoAQAN5GNp9NiwW9MjK/tq2nK
2f61z3eGVH+nCUYApZnv4cNjjuggiZsZV+KPQkSdPS1KCVy4DsYeZheozfNjHBPPac9XYCe/1lf5
+MSp9Q2WE6cjZu5PASCMnO2zQtv24n5FleqcfpTdCRJjSkbx70q7FK3X0AGkvG4bdDxhThNA/SDZ
ie1r32Sd68aydRWyP5F1PhVqsfuDnqN5TeWl3Bx5v7iMcqUKRys9W+aOiMQWPWRych4fZp13yb53
DH1eAKp2KZAojDCg1OhPv5GdW/+yU31B6i8ndwozASa2WeS/7JigHSbQsLK2UEUwm0upoCHPlbDd
4rKYapbyUci8oHzWXJqz5z6fVut7ZL5PdWO/zOyJxMMaGhiGrw4A9SG1z2OjtHeMI/whLctLsNf7
04b8H/SmCtWBr8B7CI7xO0l+yNqbAjIO4rdZYKsguzd5ONaymYILkZ9OoypV/CPNN/lkVnba/K1E
ThlrO5LARYOQTeceyDvKTLPOG4Z4T21hUQ4G3wOn9dXEXC6H7wZEHTVCxU/BB2h1pS+VIsCqxvwd
OpY9A6St2RmR3wT1ONjEM7G2E8FSrTwOMZ+VMOUHdLLBw5v+BcCxv3P0MFIzrqmDTU0NYIyU3efS
HtbMM9J4UaDAJ11EhPplVgeQIM57AOA5l0/sxiXBgQQNLCYZ3I3krMP/1hzjNFX89N4wDSEd9rvb
bt/9Y7Ydj6ktNyfOqo1Pln8sdW7wJjoQBhAWWpFizQIqfWmLkvrFtB9WLNzU5hCTKA06QGKM872j
UHy9PV8kTuBSP9SXgsu/lIXSHL1xEIjJiQ7jm1GcucMjEq29Xw2JbYvxsFcl3SDUq8bP//9ZPl+4
5HwVcE/XExkHut2aVNPELC/UeJePAyqV7xA7ZQ+XMLFZdJz2qfLxMdryZoljL/eL3Y2nNak6v541
O1mv43UMNMkljlGBFblhbXhowvlNf5rd++oHJqXW3yRRqfjNSJJk7+HwTv6RuXg/UdeMWO0stgi6
eWFKtbPNLILJZoWBBsFurLjFDzX3H07I9tKPTdTt7eaJN5aREydl1qdIRKrMoY1V5hE6QlkCz5Gx
RS6bs4lTMgwIz7qJSn50POCr22dWnK1jzLT5sNwgCX0+DbHRl5zcsO8HD0haOikdsbFDSwO6uZdb
T3lbTC1VJElYTZB2b/BayYN8C5yFr3YgIsIZZBz8su8ogis7HXOfpTdJ2pdk6u8punECR4DQg4qF
Lr9lDPqsQ3/RGwsJx3agbF1eG4PT4UADW1sTwIrM9rBnARWfWqT8qfc58Lg6TvhYcokHT0nTG3lL
qMsqiY9fWlfN1Pel/K4EMWvTbmCoNlK814vSV6vHASkpIqxPpFD/55zmD/1fSXN42PxyfS5W4iul
MeIB6BvfVTcZwlN2KaiD7Agq3YmH1nueeoMYaB5OpO6TMLGFcYBx6iQXOhJOV5I0ep9+YH8hsi0U
sABLKhyfI1kJMBge83iBVgIFIfX9c/2MDbfobGEnApq3DIhhLxbuybS8rcCTnXudQVtW0sxJz9oN
dS0jCAt+OGKv0OqhbrXvXdjMX6llL8dJfcrusxkagR2cBv3W9p0tVaajNkqPXCBtJMyUZ1dZVQrZ
tW/R6mA0q5fFbzD/NTCdjmLZ3M4fsL0PCl8YzAcvqoQvfxCbF8JxG+3NPC2qRcdknQe2S8CA8Lo3
0PNV7kjnrcCFPIsnJ1vRFtVbHEhU3t6LOgBoI3rNQZ+ETm/x29WNT1qeQl4a1di8AKSWjiContsu
psxvQvzdvHvTZ/4UOcDt70lHrZzoibTK0mlzjiYx/N0uIL/9TH0gc7kDvZhxBge9ve+1sMzVKvFd
p3ZtqH8KMDYZaoXrIdomEeajo3wBza1rmAbpG2AfLxTFhaFTvN4pHnbEtYh2vWE6j/Tzj5y8hfVK
yWyWWG8FHGD/LxndCOS9eyMmJfXTJC/uJhHawsSCL0D7e6WTyG0czmUOUxaBGD2g/JpItBThTMxG
XoWQj20NvVg2mXYC6zbsebs9TjdrSzq+MfT8rytKbGpyFlxCWItLgamU2DtSxF1a0xDrEmLbmaCP
jmG/MjUBpAjsbR5byJPz2RL2Aog0k6yCGSP93HgMwzrfCIhn8ygPclgdSwABdaaon5ZqvzsxnZ+8
28BgWuKKx1zB6Bgvm+BNS4wgFf91tjbErqJC4NQJgYURh1utS/fGXwsra6PCBaBELXuO5D+PP1/y
Q2HRTFLXwNfN59sxZsUEaM0ZP50Sw7ua1A3OCF3MKPr12VyAzO0M/m1HNLf2K8aTMKlRxfrKZeYl
EgxKTDWwabnMJYhjxoNNTwEfmDCqbyxhNt+wid6IacB//BruKyOYrOiBhN+toMo0deehmS5I9JMe
Vw8mIZpzeroa6Oc8fGlzdVykud2Wk2Z9j9bFFUGFr3h0j/fMcFri1qXyaIt21thEy1Eyo2lZLdNA
so1ep/9sa0eJLI67hSpdarxKqUOElc8RvZsK81iklavQEzIc3hauOIV/VCTLuHtwq2wdEIAwH2cc
IJTn8MWZQZMD/LngLujwgOJ3aWaBYgtKeaLDbx+nQegc2sILRO8opc8fbvyHMyO7xkGKqF8KmECg
uWPy+x3jGipHRWnJ4mH25wXgaitbyTsevpktDnfAPUJAT3YACK60w2TM41NZE8WZnugx5f/oB8KO
b9mjyeLGuOEoxNidnUCJubofRcPRIaG0M+Hl+WJQIOWagtdA1DdjkVdKvYVhl50Ff4aSA19jJ/ZI
NyGox7r0C7mKj6TALaaB6sycyQgyBvL02Nikv1J04tbDfizPE1K1M5AAP0SsqhpnmTtB8Z0k5H5h
x0ITGtZGaYqyTmWPcYaII3bwXzjfYBw9y64jU5VRu5Q99L+bHeHzU4PkG7Xw0IOqQLsRaTflBCdN
62HIdbuR3zyYJ6e7MR4iN/3Eqi4AygZcVSxnYZP4hbaQ2NofxwOMhavJobHwP3oXqVqrksvdfwj0
V+mWfWx+vvEKUQtergzGXHeaEpptDSUZFj9xRljfr9q2ajq2Jg86CwUAl8cj0UGJ6j4RA1ZiMR7n
9Ny2qQTVOdQXNRrSLOswckDEwLBRicOyB2R/o2fQXiA6QWsVa4uB/wDGDzZZl53TIg3/CFJC8tba
NbAootiu4lXKzsFHHD7KdohlePRnknqN9EUFPsLvKxCxijPY8bWAyalDRyfbZH3HaGoKMoyClgYh
xyGktZquGAKSrc1g8AOlGpZPDZrRU+I2gRiB5KWju7RWhFoNIxQkBlUnpC38237qvh1vmIIfPzuW
lqlNpLP5zWA9l0oyRGZL1mN/+FL/mw7txor7tfwxm4gp4WlY5qIfcIveV5WL5BlqnxjIu2sRjDsM
NBZg7XPmfIU4XXyUbiqpLk1l/MvqAKFewsQiwuKAfDpCiswKRzrNH9sZlQ2TxPr8b8SF2WsortIs
ly0HbIzvPZ6/lr38e+YCkZUG8MojxtR42ZCuop5s6J9+xN5e4AzeMyiRYh1omh7w9ifhwP5x0o0z
CH07F8XU7apMMsjqLiUblORM953JPzZGDy2nrKFUVjsa+tOnA1HgQOWQWny1CeQRUSeaDR8eP8sT
o71bVfBTWv5he7yDy2Cj9SGgWD1a4QIiluw2to42ROooiqetUZxB4GAAoZK1S+52JSi1olSxT+z1
ALgHRzvvcKYGvy8xkhlx28UUZ1/nTxtfEv+2Dj4VHTLLd5DqXVctffNuHTY7kAZ/vMMR9U+fFgsC
qzXgSm98DMZblTgS/cxcqpGmIK4ndLSKKnWFGGMG3e45j3QW+9cAGciFBsP43GBb/Sn0qPZWv3Ba
L1cq3yDtN4lTQ3zjLFNCpewahjQckf2y6tLppcCjW87HW794xxOEOHmL9pxlHun5QLgwS22/gJ2J
dRrFGQr3pNvzqh/AnlUWqIesTh1em5dehkPTyd2Dad6ChOPlkU+wTldNO7iWFn+HFUQEeLXjgIyS
2XUbFqagUPDdeiPgJR6BB4E3CucH1pjH8pRI0Fhxh1T7n4FVPR2jD5nrgUqOGNbcJaiFFkl+uCAm
bC1YS0S7XgRdN+aPSQ3xsLgHREEYe30x3tlr7wM+n8I7TwHuyVCHn4nysT+KokcQWoUavQVmJZdu
QC5wsxnb2/AlK4VmVdZqY/gkyfNMwUa0G0+yuBDTbRq7DS3/iMd/rQpGE1udhOg8R9R8qXgrR14I
1SB+CNgJ/5nsXuUgQW2b0e0pfTqPCRohBRbRAtgB6TIB3Qmao3ifaTQMagBzpF0LVuI0/AUSf9Wq
/44cBt32ObUAuI+DuKInfxJf4CODV/+cophISmpeK1Ktwyjs0mnysM8FEiXxV0MNHvxclh8UO2kc
dnS01bHNzZGGDdS8nhbnUqdBEuR0Bc96erWOB2Nc7sVl+DkWa9KckKTDs1E8IRQjjcUuPXLY0lNj
QxrxDSx7q8gjQwzf26ub/hKTE0a24H3Ja8ldXl8GTU5jJ4GEyz8i5JxuwDQExNDwhYWZmameuwJW
JVT1MzrMet5p/AzW9PiXlj5nIZgEOnfinHTNMF5DxK5QM2EqmE97vRrT/W4I8xCvWdjVl3U9xkUQ
PWDNAEm7Q7/sThWvsUaAZXVXQLxq6H8+W69ZGXrpxJvVShOB5dUNG/uoNNuzveb7ZMJfGzwWv3N/
nOE/rc45EbdfHHNawWbKSL0E/YMOwWLDRdIz2jqWeOJyXHcYfqzVT6eNGnmz16rKQF0xmLDRiDQm
N6Th9kBvRUDD7W+5cJECycYfdGi3Rwy0UdBjhEvtwsB/MozTF0aiVUt7ocGjRlrpn2QbcT0/Zme7
UqXM8tLWp1b9rzg0vCn70Y/Xnn1HnKLk5Y7ViDnuRvTEsMzfxt87X33fPeLbpKnquAeaGR1uftXg
Fpl1BJTUtJYSsRLxjdVCe4n/5jSiLw+nIhsSXa1+6LNHvHBVRTfbuvH+7rs0+Fr4M188qDvnsUci
A/Oe7xtpWMjTaP8zHwueKVemcEQ/dZNP2JWbQWgqoxyRw6GBtT2QZyhxXbnswscoYVvf2Vl0fDs+
nhBVh1QZLrZp4wXRFLPi5UFoe2ctjKcI2wRiR+c2czx6ZhuLUgqflzPfRtlJglk8w+9GkM6s6Meo
Y+ua1YxAfz1BXN03XlFuRSEYLY083LqmgmxqRkInQ4/me9AXdTUsfEHX/IYQkUg5mDDfhDM7N6TD
y7wwq6IiceZ6FvI/bh+VjnpyjkvheLFbYIqnZOUpk+mdQ/ao4qnmqrGpwJgdzWUbiPoSbCuaCOS+
TtPDCe8xApZavY2sXgFVU3H/w/+whVbrlcFYC9lcJpiP/uoAbHyC/ln3jsY/ZcvQu4CjJ1xoDtob
VhC1G/R+/npDUXelM2FWcw5iDDienn/35NTNC9eEext4bhpMYJklu+nIQVpUlawBZW1MCIsFCsQS
gbaRPHQNF0ROGWvVG90xo7RykbWy4pNyMRpYPXqOULPZKIGAxUhMtwWhq42kXydpVg7X3QZJz3eb
ss+FisX+XNwrPiXgxU+k53ZyV2vVsbVoG31r9qHNKZer0JyUkLCsItTgjzZAccs/h18575AxMjvJ
J+4a4eH0vmNJW7g6pdCC3WalX4ortph1muBJTvYEBmo6cMFnG9oUeWcMvgi9V/yDG4EUoH79Vh4z
BGlDwnFJwjKbyLdJAqbNc+RdsH9yNjjEfkYx8VU65YnLds4g9olid0JuZMkiNuSCet1EuucMYaBk
jDwSyj7IpVQFXWjNF0/ywmMKC4O/a8jAC1GHEdm/YWwT36k55D8O0rVa7+A2y9LWL1+GgV2MrAZ2
IDEUmO9dPSjOcE9Tuqcnoow2s/buqNliwZiNSAuygdJns3A61pV+vsiBgV4xzbNfX4EZcLwW9Sv3
qDbBe4IFXUNyngXUgrMCr/ZZFUz2J7ijsICmSlO6OawKQnU2YK2u9jvifCKMMZjRtepCwRry/8jn
cBEiI2t0N0CmhQL+4XyeJW14YkAbZEUUAI+6zRz+wscqhlYkbDQzwK1S6KIDVYYDSS16LuJyZgda
L1FSU1eDK5aYTqbaSqxC0exnKXXd4bSQYmgFdfT0f0XvjQQYBPBdRgQHiyaCHZQ4wW31i9/YMNgO
lVUKfd3L+klroiu3NBrF90Yr6fXXetPRO+DTiRiFC5YFyGDYqAgq50mbL4MDSkLOcEFUHII88dB4
C9nFVu0hlmVCDAV9XtZmO5bRoGndRo7Nh6iq5Dq3h4zZrSaiOFk0bp6qDv4UiPyIOvDIJl1F01Kz
E8sZCPhu/rtUEKRw6ZA39j4VII575ktKsM0h3DMi2EZmLV4bKCO1ey1Mpa9KuBsiy5cLprKwsZ37
NUPSvopnZjhLzXQrc0YlSSjCCuV58qws5hPWHAweWmvEkTbsfIjbDuF/WhGKxBbi5vV75XA6lzsP
MIUNkql1I+vXTLuKZ6wubniS8QwK+yLugnyc2cmuSPbX2cnJkcchOyLsblIXj2CDIKAt4q6RS7TM
MxRbObXDmlo1DdLjktLuf7fiYBE9GrYX9nsJDxwM6wyXVEKn3H/RRRIvYRCbG8yevfguqf4Icoph
L8pMoL2Fdm5+pDuBuHMsebqJHSxA5jv59tooqNSRB7igPIvkZsgMQf5HGBCRJUcGpfi3fUXRxWJf
OeCvx1Xwm231acIF5usI8YEsE+4KaI16ATCg4js3rdRuwywkczgK1unNDf9e88kmT4UqHQjnoqXI
z/SumTB18LwygN9xSoYFraXURbCv10D77h/vPSuf4gI7+cck6gMA9DL14e9U4De9kZTnSxkB+DCp
UW4oa7N5ag9tGcrNHHk74y/FoNqhLYe7s5OvLcYY0QZt5hAsPSWLUPn8Ww2GDB5sxA2njTuxlaTT
rMQPgj/6ob3l1ztNkEeFU6HqCjqubHz5/Tu36X9IjTJ/Tl5q0CTiOwRnBlEWzEzVfN6OdCZZ6zVv
AnHz/KX+wibgykwDsS84QwH4LHbk0kPN/8q6MNgCSh9M8BA4bc2BbPeT472Nwb37A68Wm5AnQ1fx
n3V5LAZgozzZ3hoO46sGmi+mqcFx5KoeLEPy/gQ7hDmArXTHpuBKLYpx2gecXo67DlFL3/jWxa0e
Hfm4KOicO2ci4sFYJtjs+t6Mf1BbIUgt9n8w4hPoftHtZkVlp2FYa13GNaHcsvgNAV460IKiqW+j
PfqS1TWAppoJNEq9mDrZaWdDBR79K+HXCT9tT+nAUcIEhNoh+3BuPtXnKVzA7fIt297dW1kv+ys0
utFGEVp1tew/BQUTvqGNzaA6RzwctKLh6ZJ2i6ZnFJZmsLTyIsvUNCzQj5ttg95l93y28JhC/jQ0
LL9FWYVwNPf6mqBUbAFGCf0UCd+aw/EpVhA3fHQfLwyLDvGnpiZbb4YZ0/uOvL1J8lcYso6NYhNp
i5baXN+RC59hQxO4KZ8A/jtlaoGIFkrXmcL7wGV/BRhHmokUz9k4W21HY7T74od5Y1bzd6K4Z/93
6gCRuXLlUmj+O+uBr5ISI5yNzYgQ7SnDJuw/GNCTCFSIMak0jyixY1mMxpJgDUuTTJCcujWK39iF
TU0Yt0LIMsOw8AK71Mc83Sk4XHqoU2+Dc8OqsWofAp1+pZGaSqpWlJEypVQWsMvA3zTQUo3cbdaA
5IzAA94gA/izO5Ghr83DGZVdMLTQtf3TljTKzqixkDvFf2LfBsenJq98+AAjurmPg8teg6/iVWMP
tvxhas7njwMcPwutngd/qaVRcBsGcOn7/B7tIuMhAzz5zUfloOug064FSuEd1fZTTAeDNsn3Vkew
PjWEacdOMQ0K3UFTfuhvdhe0Gic4RVa/vMdhiMa/3tC1Xbc/2vJGhog+V2wJdGZlmx2lNiITrmiq
Hk2m3srwetL9rp5vH1bIrXPGrP2A7okSB19kpqsQkAZRsZfrZfa0AQwGjTDdr2w6Y8mthVAdpKAQ
IHVJgEwTwzQWBRJJRRZbKGj/tIp9PaVVoFlH8keYxxMZxHg0OJIafSb62IgOgoFIBP9w313otisO
vv3YrB5Ffo9bPC2+VaYPgTW315P9fxwxpwDUlUIrLQdjKi7nfUwz2O+ekc+zmHVmMEZfRIpzexgz
2Lh4kN4nkF1S75Dn2bs/iw5E3nUIiCKdtHtue4/bmDt77NT/fsjgibDfZg7QqGU0GZ/zz6a+TbUv
d803vxISbduB8T/dS+Z0H7wi3sN8Yow/tG7VjgaSBo9AM1GL4iTN/WJird9FQOkPTBp5lAdQoN2Y
/f0NKqpNJG/NSZRKuPXCWqOF4wbkiALtXlCEwyc1Vl8YxeanmT2NXBiHuuP12GwvYmOwmvSkvRM+
TbVjlcYKfcdntAzPfj0LBIc9vfXDK9vsg+zBJSLKpWybgqjoUPR2vvIMoVr2SINRX4u6VmIgMxXI
63Kp/1EdTmeRePjheTmr+tl5+CxCBR13e+vjf61p+X9XwtvEwk8dSl3y5v44j6RdITzPBdhy+Flu
D1nj7qlOnDWf+9P6bo7g8tk4UH8dmSNsGADrKT0j9IYh/Fs8GaIa1Mkrjmr31ArbVI5VN/5e7dnq
c7onIC6L6u7BL+BXwXVgaaxZV9q3fRH6F17QRaWRtBcKL6ldI9w1REtBUXlCVt+8d/m1P1k4Eo9i
OOv+phZtoTdWvzFC7QH4j1bG0C8cqH2nINHFS62fPHn1HojurSBJk+Q7NsCc/juUzLaQ2eReorCk
utdEINpwNGADEnm+lqM/+xwDf4qHzXRLpJqqYfhH2adX+5Sy2ieQ0gNOXB38DxyF2+24paxR4zii
mtbQ1FHPn9gbQsqwYVtjjPyqwSXqEYxJ6MS3t+t4eDtz/sdUo4FWRiePKaXBPmgFTWm4RpFowNz9
H/2ao++rh3vMBKc5i15I+3izl6AZmGQJuzoTZoevcWu8FiGCCJ+T+8oyJruO8jGfYcTxKf3LgXaS
QlGFtzHBucx9hR1DULqHz3KL5w8zmHY/Nx+zO9oJacqLDxysGAL2E0D87syIYtVQCw+FYlK3zFcD
zCeeb4DTMvVDjhuAxvAHvdCBY9d+FiixaOP/NCJg4JoTY21QAvIQvFbjNcX7g4kt/clhvs9GsI7a
aZ24ZO7R/QYO06Xv12SaZKA1uV+tRR48gp1u1cTDvrCkohtwdhvMdtWbGV4Vq7i33DICr4DZJsxd
Z2/MLAA+20E2urT0Lru2+NkDGh+tBbVFS+J/L+6hsJgrdnvFZkH48D6xQX9pWUWtL58h4d5TeX0d
/ugOqa4N3XFtxVK06FLMHU8Si3gsGgEitIgDq3VkyCB33D7Z+yRsErZOCj+JmbPGbWaCcSvXTCQa
ziZxJGmEzvCekCwt85mDOi+0RqiTNAMpsCey3ZiVulsFkAdo8o66baG6MwNj3PTSNsTfMJEAJ7vj
/rOYa6hPmWgOB2xg8zm622irT1Nz8LW5Y1DfqRaVR4OHoJDn6Z0w/OauANBPGMuhWDRWanEBStUv
vX6R5U/fLOctdWEY1JQhs9q1VtN/qU4HbCzqRT1bIpsb2e+pBAAwxqK4Y+Th1CV+BCyRLsqg5eFl
o1fB14mWI1LSnCNwizo2zf1DDLOyZUBPzlizXmkOx6AJlYlHfHnJ4PaG90Ojxe2+/6YUGCbajJon
rmxgTSwakAl41OM8BBEFtG8TvVh2rsSVjwL3vkEme2vgtmx2OQsqxietK01Q35HioP4g40A7JM0u
kg6E/QCba0gU4ZFTXXVFihqwxvpNaHNWVqHbmaQ+kJZHRsXCmRZH8OKp/XBXJv8C4Q0mtYTpUZvb
0SZJ8vwl4xcG6cE0RxGpV+u9UWoQleqPb+jFycJyvWMURVNn6Vie4Tbm9UNHSJdJz8stxGY3U522
nSe/3/Vb5Udn+qW+28T09cb+Eh23pAYVQpF+SFPYgw6kAwRCttowk8OyRHZWKcHgwhOvcoYwvMNk
WNKtPCWi0Lpi4iBPLZnWYF3oiimiwUfWVvgbXy/dM7DsBDnJgIORQf17rlY/8AvPxeRAwrkNDMqu
DMCmn+mpeoVmDjXkTxEYOGp/1skXrFFKqdBjtucBYCyfmp4j+okQ2TEa6h65ioVHJqto7WO1LsS3
+EZFZiCsYjVMwgmhRUM0Oo1JyvMRCRL4ARqlouEEiN+ZdpfUjYIWFuOex8zimcY49g5LO2JjvPh9
r5chzHUbT9KKorWftvY3tTob70bFsljdGY4kb3gx39CN8JyKSFwk9NDdI/6A6SFWKqX1GgREv0f/
NxZst2bfhiTynOya3W92log5JjO7FkPKJ3fwsTp/3Wewf00rrCD3HcaJeD3tO6KfhoComKELU4oQ
I3KSq85Fg7whUvFGLMiEJUT0tXH9dSV8sAQt/0j7oNFw86uRX3pfPb30VbcIJBdZCLGp3qs9OmH3
UeGD4DdjI9yPpOH8U4a32Jqaqj9S66yTrqmczHopnVfUXcsJMZL3rAfrgDPV3IdE2G81Vs+3tGHN
IY+R+XF6awOFl1dtF+SsDV0lq63HHIU1syG5cAk3ygw/sbO4laEtYeCk++SSqec6xr+z0Mf3Y28g
Ur4OYaRz84GDL7DVqodk+kVo0AW43ZNRiDM5Q9zqfMNS5UcY8p+6/a21yUkOLzgB/wHF5IG+s3l/
YSZJtgilidtc5xPmyd2vc1tF3F3aVm2dLugXTP6CFBBV2+WMjWsDckPYiQ86BQbo6pd4Mcgz/yoU
PdOAjfM0wXXI+ByCbkZpVkI5ygBOQW+wuvnCZ5sqXSKG/tTxf3u28NBz4eTopf+BT8ZZx9aoQMgW
KAc/RdrnuT+8YeNmSf/PPVLA+bIimd39tOuu1BpqsL7nWW9680Vm30O7LwBIdFELpdTDnEpOpcxt
DYqymIkqrX/+za+vYsNgq4v18H/KinO1kAVdmCCeIp0Sred+dIylqRxrBTYNEWMaIoR6gTZp5u2Z
IR8exgrVXNT6t74QAoz5JZnSJecMm4Avvj+4e2Lunm7vZUWg79tnfGnNJwblWwvGcz4QCE4ySz5a
51cNDUos2POv1QZPVtYfMKIHWgsePPV1W10gIWVO99fZhVZtu8bz5BZnjI2HbrMtz3xOofobP912
T/wt2hFH8LSYxHjNX7uT8PN1qT9OX3MCHtHQpdsbQ3f+sIo8P28q5hgsDx+YTtWcOtFia7PvIrBG
LfAVcYIvEaMrGtTbL8o3gG6T+neAQ1WuL2JJ3t0jJntR9tiXNLHD91A6dZYG1XijPAyTBRlCXWAo
6cfFT9cXiQFSt7owwj+K4j3RoNz/i/z6tB7nOCEPMxfMciOxpevTRegriF0xMVsVW3pTckj4yOjB
/pGnQLAtxrd/AumuBWfwax+qwryAN7M8KEle3jJCmI7h9aBDgf6T/sxpCiuGvC3HQfkgNRSG52r6
ywV7CM5wRDaheX+yAG0Napfj55aSRYtgYHyJZp0xpGeIU5wDcpuzCeND5xpjGhW0lfUYoa1sWryf
bN+jijmhaqPpP7NgUNvJ1n5wvNgznOQR7CkSL5xDFGm16qecZVPk0M2GVPKWyP7z7kYCaiVehvSo
TbAuNYB0JRmTeSAAqrIeYDH75hlbUcdF5L5NysVuSAOs0v3p+o5kPGKaArgh3sGL0vw4uOpFEsO6
l/FnBdpI8FQVUiWXYoH33VoEolvzmnOwAALwoHFY9WWpIcSzdOfygyZ03GyrCMUxyXR48sW5GBxg
ksb+D/MUcczguRpntSn7KMC+LETSY5KZODu+edOWH9WHG3/XNPOalQH9DYjjxMya7tm+GEUHtZtL
Ejnx/mz2y0glCrJguZu/0fB1aeIh3sK440hwpgRVLS51eAkzLfnRctkS/Pl0TszfdSYCapTTbtHp
UFPnHpAosBrUj+2f+KvboVljDCw+TDGj3oqq7AVqklTjcfcP/mu6rIW5K/rEuUH38J+DAM0AzaOB
NTGxXZzkj+Bxt7uzL0E5oi+0DvUVSnKkvkEMA/Qk3dnWv2pMTdBNAGhDqqskZXheSuKwlqK/ucyM
h7OKosG49ELGw3/T3v0DXnGuo9gxIKWQ+DGMCQKL0P2aUa778/R2ray8LKRgaohpzlVEMjahFDF5
uLmxXlMheXTc8pcl7Y3EZMBXMMNwf10lqKOByKiTPcl1bfe5pJX/d98GOEJvY0QArWEXNsaEX9lQ
+5vXO7IP2RcYHooBakMNqthE7jv3CjcRkXZp3/Yc1M3XqLj5Bqhdppx3t5wqNIJyk0C+vxZHae0Z
k657Zk0b6qP1A7bX2MnDtd6eLbZxL9beNwIGfRf+VQ5IGTjaM4KPf6UzqRkCvXHIzziLnFH636Mj
RdlLWgGh1eoD/+RIeljtzHeCiwbo/x4bFjyCYZOifD0a/J4ZoE/TspUEHvn0G4ZqVGHoppNXJCHv
7CD19iwK5GtfihcQFrkjGJArHvzdYiifbnTksktjMfDlPfnnoLl2ic2pzYLLTyBb+s9bpeM/I31D
uMjwgmIbZS0s7pSvC/i0T5HeHO23Pxw3mWz9LKBd10f5upzUCkPNh81yb6sJdmevNHp7X8LNx7RQ
2JlAI8LT+jYJTTkZemWckYAC020LlNqZK4xA8/FBf4+WQYC+VpIa/pVRerjdoOdYkDzxBwAZNdJf
z+EOJ0c+jiZeyaNBxMF6uY4TaYJGFv9K2ZTyAP/fxYHui8s7awi8Ub60MCellMmNLH6h6RTCYAWc
50MQolQ+cr84mJH/brtie34Nrtt8OHAOuNazl21wmSBr0H6zHurZeqocfUKSZz5jMeCbmAtlAO0s
bBvlScWgquhFJWLMowZV07l5MdwHVIVbIk3l20vr3hm0sRFyxklEzRWWHjJDH0hs20RGgk2nFqiN
sK6fbAVZtdIshed6Hht7KhZpSJ5yZoPTnzXIpMdfukYXqXA6aLfpn8bV2A20UrrNdc3C/UvpqO/F
mLkQw80JiPUP+67PnSMTolLJc4LAlTz5QmKHwr8jdTxWUAFyKNqPGN5EJpRaHJCjSDfwDccSoVui
+nEawCdaIlW0XnqD3f4Y05FVJSErE6xbKFHFoLyjo9ONwCNPOHLi3EmEs/RoeWf9qR0cge0tqENS
kYeuVxc/8lGNaZPVWvuzx3/1N0szCc/HH/AeU7DeBjUsg3eSUVWIbHmWIkYHTrV7ZGH7+SC8J27j
BO+JSG8yPTfUbGHIfmjqHjP7gN2cz0ocS9alY9f6j90TJgSdYByxgWQuAHXBzziMxOBv0pV5p2ra
A2rrJ+0ZuEag4t99oVNnVrX/eHzrBgJwYhxHZt/4wUN9XCR1Jfq5MtZwB+pVnzlVzsTfiDSRyUZi
AvIgxxqMjI5M6ycKstap66+zbxucODlUqzN5y7BVQSXyO/RInZLg3obQC5IZbemQ19BYO8a/qet8
t5xphcuw+6BYoNvPaOV9EtDHYKDi5338L96BFtSeVcU+Jn5TSfcz5RDqbvZ+ZiE/4wec9u6waO+S
OrePyxto7C0Bg8UFM4fjuuRi3edxHUVP0hTHOhbCyYICBt6uK+lDKewTtF+BK4SRW9drOkskipaj
nB7bKzRyzSpDx8nke4t0IkXdHinixAi2BPZpOhT7fiD+w1wZtNkQqLQ0UQJwjBOgPoJn8qf6xLMM
8xO8Dfu8wdC4LaoPW+DwPyuoFqEQdFkKoUIIP1HYBYGfArQ+0Da7o8WT6rRpRfWlB6jBt8cqvd+n
64dPisugdBhJ7nf7V30vew+bPxfP7jsBpoExuTSgg0KECVCWWnfM5zMz9m3HzEWDqkqrBMWvxwHW
H5l6SvaUUG32mobYdhtgUaZRfmv7IAg0ZvjsX2bDwCSsN/A7Z8UTryCUO+loLRKILzkyB7NvAvVi
mWTHnRbY/U4XH4NmkKgqsR/xyNgLIoLkBbrELzX4jKrGTQzw3MSXX2REZLx/BgBTLpdwvlSnxQcZ
yQHivWzojf2LpOdXsZGBTsGHYKith8D1aWcuF1ezvH5UuCeF6menU/chy4jRwCnyb63KbnAjef9/
08c58AJaOsQZmuRHDyxSJqfpWEqWYRO53lcjoOXkXasj1pWWhdf9zrqYMZZW4riCMghvKBJvrdlu
isUzIABtSg1kGc6I2oHXxDVSubUFZOH1W0nGGQQl3U3zKv5D+Do1uqzN9KatQK7D1OqJbad4efFF
rfoTXYytSX19X6V4C16x6wCCTvcJb2SFWcR2EUJQyHo8IIbMnFW8ZtyMD9Ixm7/mCIviO+RIBUqd
tGcJByZxguTjYhILfLvsdIcwbRfqRsSTW+YdIRZO8Wrhx5T1lhxNJ9ZqgUcVtImYSQxgnBDNtseP
hOIU7uksh030aRiHBcIDWMrq3zvnxCsGF5njHgq4mXrIQy0CJeEEHkCp/wEiyRjexYoNHwACFOmc
aJK4b/JxaSgGHq48HRZQMiwC7ZtxTHHdJoyE/3wrf03NlL6hQyZGyr6cbiXtKHmkrlnXg09lYDF8
ZSZyB7EHwBX785cm6NL+RkSFfpr+9XTdCs3CQ7oe7WY7JAdw6pm11MJHq8u6ZnszNdVRNzUY9gJ6
hdYNwk2uLGk2jdAGaZBDWd2dafu21KFOWyIHxytahXfu2X2O8UJI82oIw4GaUxBMUT6qIMhUAkjB
iz5yej7YFB+Zwqnt/+ECH0Jygu0EwqeHNR0MBXM1WGQ50NFs6wLBpUszjoxFQe0278Fg1kJgufA1
+2RY7oyv+mq13cfA71ioFuOy5IWs589fxnot7v41AW5hi4UF3cob+Nwhtj1yFa2xaxtP8S0HN1r4
eLS3Ps1nuQeMyXQ9FDoCWwtf2iyaq4BJzz7d8nWHdI8xtsUT4F5cvQ75eeZIvbWmdDg5vytRXiUR
VIK53UzmLpHRmOmATZpLMpqqPIWFt7hv6rfOlbfniC/DSOLioxZwzbJ1qfakZy32TUN5htNp4njA
xmSt7vNHS200uTbuFYw4MB7HffvkpdtO34FFXjoykHPEUEAmRF6sY7HJ90RqPjqqaWINRu8aCuMI
rdHDBYl2AWSIGYIP6lOMGcYNAp7z1sCLWMtMynmN3PsiLNPe/9xvNba214siMZBM9Vx5TgnlqkEq
rPElWm9xgKNcVSBeS4Ns9LO8l27olBLOnPFMhiTzzXTHZ/aHP5gDR3V1laoMz+fVe+Ld4ra9eOyx
MvidawuP1zuTwiDYjmcyTjofgplXbNbh9Ia7HLCUFxaCMjMMhXp00hl0wjNDJmklr440qDFcZQNR
dPrtRU9wxVBBH3VHOsdELZ7Q+JmPEoSe0qd7tq+wiMN6cqYB/wYst+bTy0PyhIAvxi8OwP/gireY
aM81HAudWVooEr2tzvIZ+enUhxV4tyCYtOz0Ya1Yo6xbgOg/SiqPOYG0cYQdahFINRFVuCthzn8p
sZEI54EzgCBGvrzmCDyyCDAbt49XQ4843WitYl9wYpLkW1VGP4KrS1sOETbyt9Q1Hnf6xeWpcwSF
vQ+vQFokjooOTZkwhOVr/ws/kLDWEp72VUNSpe63YGKB1JpopmNXf/KDYWbOUusHFFkd7kMYwz/G
/2/OHrEPN+OT/UmbxVxpCQLg5dsDAAuUCA6PqN6EV18ONLn2p58ESzFqqtAbjwu3A43tsdCdN65n
wDx6xI0KGB3pfmZ0e1stDH51/ApsPLAaeqX7ZPaqzS78esq6EVczClvGb1KtWTWgCK3JGR4JSPEg
wroyMhSPyE/AKy5nuPwJRyhI9yQo8gdR+VUUbpCYsMMMT8+P/AZyxvoIVG/nKTmI1LhlwPAyABPp
wDAK80HXoYXzlCfuIESlgm+yu/qIbaOYUDVYhbSsCFSoMYauZT8Ig2uZHia0nWRJofpXWz37w+si
pqo9wY3F2TfnohuWv71Q8ChpsH+WHRI7Ka1LOCXWY709F2TevTN/c3VUiHXaD7a/Fver1DHxjFvs
3Xb3ZJcdKJ9Nbfh3CK8DEuOJkzZVdVVS9hi5nO842n7ygBlASoa6d4yzOHBvYbq24kzbpZa6ayxZ
GZeq3aK5Uk9Z9T7WL4qQ+vqEvpxcsxKOlVoUR/oJErb7EpnIsqjqqhJ2h65su16s1pJhzr4dUR0d
m5Qg9neJVqXhQAYB/o/ksGlptYRuXU3i4eLjvEXbpDxIZUfMJyQPnwv71ubg3A6rwD/71AAVfjDi
sqihTvtpn9g1GWIDRAUQh/+BGiHodizXOB4fDssdmdS3kZtsM6kzZ4xZ7WwknClqDkjsAQQQ/4Ut
Zq+6rC21NihUQxPFhctzAl+Jmis2IEJ8RpD3e7tt5gdo4j+3h3HtWQ3It7KGsY3LuZQGTzSTE7rN
uGsR8JGQl3fEaG9SkfwUQ5jPX2osI7YB4LjjTZzrP3uKwld/ys9aNFots17lTaAxuqdIs622hQ+h
/lik/IljkpNR5UWkCr3FIwSY6raU4RLnbPIMkgHKvpWZa+T0FnVocb6K6HwQ1DOGLEyuHGXSh059
3ZBdWAK/4BN4FJPOGij/4udajcxCAj9X8jXEN/4PAR0o0loE/M2DHQMAoAZGNF6Y6QJBthqCUVz0
Nax+qo/xCf2r1BTs0egNj1IHSG/V8FyukkD/JDor6FkVlgG63S4wjc04GB26qyocq7n0S8tmjuu3
twblLzwSyw+jgZc/y8vo40XXCNkAmAJVFSBXvYOKlii9m9AKFe2ivTqHA+m7nfjnN4j8/91Ux+0S
TCRX2DH1NaYsndOPe3g/DU5Eer2TeTxO7UMAf2DAvZ2LAPYaiIpErWDnelC711sbCGcJvRwHAlD+
00LNz8TBh7aPOsvfGEIiWLS7+R4NXY6+pON193aF2dMspoqRRq5uMnC/KqR+zOlK4WhU2oLuD1TF
l9EjAngxytvx969ySXgjk27YI0QvISs9Kdoabh784pIPyWvYWmuj8r7UEwi7pMpRm9pHCTM5SaeK
HPPjWIG9WROlQZH8MfcEL5oy6Ud6D/jTCIgxFp3AE3dG0JX8yIzIMW+myMqVHyIHcJO0k4lBtqw/
xglF6GsHO/RxsJ1OxZGVQnDrbBtR0DZi00dzJXpJwVzRKx9uRoX5e1U5RaYEiZSahaRfW1OgEROD
aEpY60goAQgd6iTtMEIjsKihG1ts+4q0YcMt2LRqriwcI22aPhXUbJu/mo3j1z03K54lO10xf2OU
EQQ/TZvahnT7kNBp77eXL2NiDcufCeOOgGDjpSplEpD3/p6TwoMlu2X/Cnx1ldz+4pSzEBjFptRU
IBxSgjOcQX2P0mGgA9mted/H/EhMPsNAH1C0zG97tJSnbWhXuY/W4uuSHA1FlU2OvCPETojp5jq0
mlul/ClxlheFukNzX0EFPwRmzybJ4PFKKQZfDXTAUBq9JC/QCeYr7TUi2mZ2lIj8808ZnhlyDZQx
XeziIEshEKHt2DysYAdRsNfcmmuv8Pv6DONJLp/YyrKNrB0GVc5DR1hUStPJzk4IHG16uSSZ9MMo
gY9IylOL4znlSqc8XwzH71UllhGlclWbk3c3JgCITjil9Xw6t0vYIHwsYwfoUyZzGsMNs/E5KnZL
uN70WDO2wVNTKtrduYtsVs0xh8b/g+5Zh1KFu6PX2NwJejX/sIE22oJgDc2GVGn978FZg0iKtuhO
QEpDHielbW7FftEtvRCXB4qpP8hqVMFpY5S6NW81Dqtpn6Zuq2ldjp/hWLqIsQDwNppgZnU8N+YC
DtdvcL6BFDJE22IVesZDEFbdGfvUCDaB7+0EdKc9fu81yPnuskYvojL2530bALVmx9HNdH1QO/1H
mRn2JP9vcgtmjJTVFOP73yW2WE9n3k2s0ShnfeXBi0xKZGY0Oe4XfdobCCgeFGdovTs8pRKFJVas
3VCtm81GYRoStzGVN6A5UnxDFU2CkkPqFxyPKTCnQ6lsZ15zejnXnvwyi61zFyinXun81+snhtWz
8+pbKf7+LF92CoL2SaBTrvDb9sJ9ehgen9d1+Hh9xOc6KenYvi0KUMuFrrTc8IIoAjABE8ixyllD
6oFpWjo29aMP3VMNZpbN3p4RwrUoNDN9wwrfI238uulUywmM1/xAtNhJ86HsDW+nTG18v5l7qdrS
nvbyUVvdLvTbkdmpyfPCKdWIiBENDY5uU73Oi1iqglhjiVgDUmphMZ9IMDoubP7apTpGUdu0VcWp
DY1rwjJ0nGNOhgSIFpBiVY2X+OBgAFAFhsZxizcOnFXk8ZDNnwa4zc7KR51qVuEJJIRR8MZiQVc9
/NtePlxk3o9zwkE2NGCht+c346QJEJHAVM01GejTEe8FcjkhznFRZTC+gYGBVWTB0JRoVsSeQLbl
AUWn/735cgqsRP4FkMUN2LbNUJOUtenw1j3YJOOm0MkWnkLvMkFT8aNO14wkXRUlnighpNYubD9R
1fA6VwC5jMkiJmTrG93VozrGi24ajKzTLb7ayXZGSuX5v7Oc/6Qq1HSCI/gRGwyjL13ihq46TIuC
c7RpxugA9x2GRJ3CQa9XJ/g7Gl4nkWlUMsPN6uJhpSNeEQt09HFEiDTjoQfq71TDb/W7PERzv1jA
L9uipnA2IqJgNGDtYn4HddBPO3GmveAcT8qsQZUh8qsAQW/8i8K83O+yuC4clWPOiphyL8+/H+aJ
7Ld3yhcL6YAOJ4+aGX/tCkEChhjrOOoBH1yUoQDShNLdCseFkeqXcKzzEM2/Z3HgrA0ri4J+hQkO
L6YyBXY5uEtMfLtrVKykq5iGqR8h0t9qEY9PULSox6uiLzU3GORWz/S2e6P2KjGVNJ4nKqtq2tF6
QksBeCy2+Q9APplBPU8cpFz+I0wLWZxZITTNb1ZMIZYV0JrpGOo4WKSC35ittvkD8mSng1eRBqf2
VUOaSo/Ug5XTaonRlrF+G6r3ch0sClobyxNp2ssNiCLxE+WgRQ5vPfxiqJGCSaCldyYhoXsm7YW0
PZhBWNYGbuCTeOYYzaSxtXLnW9FcBNTKr7MIzz716Ksig0yy70UwbzA6csPSUyAO+FrWQBN4QMCC
jSfCfL2b5kGB82xIj7OoU7voC7auVZns76RuGVQXbOfLzyCfJwoFk7HZIy/GcgtLjoNyrYtXW+qO
161N7t0DHP6NtPEU4Xg5UHbVObGbrPIVl+sGchz7Okb6e5h5T28yX8Xd2U0+g1R+xJv9gk0So0xP
qgnLbZeNf9qS4s1Z7j+BvzIF9AhoZLMblpLQkkBZTadC9EOMTJMJnGuScYMjrJxR61vchhfhJZWw
56iDzazVCTg/Lv5KJXO7Jmd5Xq7xH1TWQVLpyigotXhquQqWInQn/w8SqhOuAg5ICMwYPPvttCQ8
GVzfPA8Dj1JpVHg19bxmkJh2W1lc3A31TscJCbr8Sd3cNvYb+reNd984yZU9fboTb7Y9A7ojy6gW
QTUsaqQbwcoYBKZk47gNySrWvRD3EAlhKV/NHTzTMF1kYxpRuHFlQrWhD+obLnDJpxrNxduFpAq9
nqeTiB2KCfhZe8KgLdydpovNeb6yjVz87wUqLSnqQiF4HAQzFNneBCTwSL3gl5e9pBLSbL2K/79P
fgjkoYw7874hCuChhQc1mvUDSubhJUjarLh7J6x1v+f8tKNEZl3jTm6YUIpa5M0l05khhwWDdvxZ
D/KMj+qlBKiUIReC8IAmNvh8yC3S31EpGNzwb92aIczmhb6UtPeW728dbCC0pZjx2Q7jetvaTnW+
+YDXhn5btgUJ6yqIoe2umSWLGFXd0n4KVB5PlAov91Lk8lls0c/CgcV5lL8Sqe6Nv7QHNNf2Vo2k
HWkU2BKfZ3u3TTntszO9lN3navQW7Kx+oRvfr+J/It0zDVPE6TNn3Xf3Isk45xVrG27vhf9AKMZq
fCH61oFnfifsUWGwYySPGR4TQi0xb7BKhpXYX7z3jby7e/h57WRWh7Y/ztB+V1DAILxjS7cyEw+W
HxVqU2qCtFlQg+9U9ZrWwksetIRvEJIoCQywDjbETz26H9NW1pnDHkCKoWFq79DMb3ahKginEMQu
uVsW6l1mkSendAqva1OLyf/d1f72+9uiRRvgZpXH+CtNoBGxqDZ2KxFy395T5t13iweVdwDOQv/p
dTDvEsbcXn3en81Lvylmp0Ip0ieUJj+q52Q6QOuSxu4U6D+IHoJ2W8b/kqkJJ2xrBciw+uL2J0co
OmFWCj4uKHwvwvrkBBFGITQo8tfoBv1rBDwgEu6kAb0JkPl/VHIuhk6x2oLRKvqpI9iaNTgoLcf8
eJFP2hD8UOgscHwUOgN4mYRY1nt4VDRxZ//up/ny2CYFNnbPvpUVQ8vSPuEQuWnpHSghwUDmOELB
Jpgpq1vGasUq+mp6ReWwq6LlXYgyNAe8cJmlPaYQtqYQaMVl9vCjGMJxPu/HxYHt+pbzozVLvBr9
g08Dp+FDzvN06w60Fclf0t4IF/uXnbXd3k/OaOOSj9uJr69e0P5ShlomceFURI+ckNhFzOLKXR2G
8qwx/Dwq8fo6RfKn3LSv9gEpdNWgb9iX+Pw59WaeGQfDyUEVrtE1E4jQwJ2zLugDxa5vL+IXBlih
sbKzJq+w2ZLtUmmgCDorO6dBaV/65vGVSkJE7koGJYJ+WGJ5RF/RFEclZKoa6HJhA/xOS1NJ+6K+
SkVSej2Uv35+xCoQnlh+W0Z/bvJc1iVl4QXn4MY4BJl8wx8aaP+1VKFa0Ov7G7zYmJ+eSuVW/9im
hwir0kIgivc2jQVlM5AD/oH1Ggr+GzIhUgC+t6yuWdLPUD2zYwiHg5GXlEz3uPyQVB6ZrLe7VSxf
1+uAyqzY2ZlLllP5muEvyyjXZIZ7DrKnb/XwfM2HBxsxaEnshXYRxigKOZBCR3RjuJwEa+IVDwLu
yreO5SxSCi9XFnbBz0r4XphdUuzpejR8vH0HgEFytjKXIRdCCKY0KOe+UXUb8noJMwb9PzmttZvq
aHOmhAeiaBnQXjTIIjSJYI8Q5y+mX/q/HkMcOWVtkDkYjunp5N8OdIdmHxrm11WpbaPceNYYvH2c
tb2rsetmNXUE2nukQW3ExGMhnS/41zaXFa7LIXs7u22zX2hjW5zhbli3WkgemUn+72Pfu+LwEtNi
T4b1M6Pm530x3rtSHkekYC1ctu9yMuijJHkBu/JKSNJAIkq8NGmAoLbykFKvrFUNtFaXoOGRk3ak
PFg9n+2ygXonMZoNjug5cmzPPTFedDan7AOyeVSJ31g4IYe7xiRJWB2NbI2NGBU4uu+03EsOw/Kh
lMbivUa+rSkytifUJqUNvIBWmW9jL0g1FPMvwuRgBwsRX3HEgFFB50boOIRiewEm0e9uijyPrZfQ
Z7+8Vo5jzUo6C9cOQDOxgyze89emYjOOfvg5Hs/5YrnvAxEAmL4NhhzzQxpYKvFkOm7xIZQBERvP
a6eoPiefUl01jq9EyBx8hBOgy8ivh7ReGVw0hAeJHyDhxZacvrKxBc+7EZ2UOo8sh+f2buPGPCRl
DhIGeZqk6W/hJ/wBBKZ/ooV8FYXLvFS7RsDIfoY1l3HTE8zeYXSk1yLghg6NIbwCzk1TT3leUX/4
mdRsQMtsSBP/OYGhYinMT7sA5Y9sVxPtFIdmGkEjqZWvwuQ2rsMVTrn0OVI/eEhSB1bL99Tx87gG
MrYMyEjXKsmjC3wzLuHzNPg2HZCcRd4gPWLkcVrlVmcTMMiTjfwXvVjdumQ35hSRrbyntaYUs5pD
IbZl3UgJqbllaSVXzrKP11QJ6RccJGHak8n9LR0z+MHBbD1dMQpLG0mhZPLIiX6rB6u8ZQLq4ylO
PF+UZ/TLDbqtubYuei6ighEzhB+x6/LmM33KGxBCsLsZMo9otsO097PxTzGBRc/tZzyvdSb234uM
tXu+FcevyaAqg2pmRFV4AR0iIrbf0OLhrQjtmrLGeVH2lKD602/+p9jl+F3qD3ZkOAduaJLs0/fA
y0BuYpwgSJXwfGjYOcZfhyeusVe06gpzkg1yhD0YanatVN/gi0Oyf2uBXSV8dRRZAiwyAqr5yxkm
e9F1t7cKAnWLwJ/+SDXABwOhcN5hAA/FpQhiRazIIoH3eVDRUXK5coW+KGLmrbxlVkxxtcLxbhP/
RlF4opCwImougJYC2ststE5YM11YN3m6cbwSmQS5HE84xa1YNPD7mxp0AVc/tEQJau+ydT/acdj2
33dOOJxCeG3gAeswbmBNes5fqxHN7f4DXsn3oS06O/hLHD1iluTNMfFu5NmimlCGyFTU93kud2U4
c7x3ZvasfWvaKHSpOUQWziN0C5CMHDdpW4El2FoRTK80LKCSqJsaO2n9/kLFH33i/qscKgQv8F9a
qpDMQW0WxGYyzW4nhn+5qxvATd8s1mcNWJYkI0h5lGcMEg9lIxZT/9hvJyImnVccgQWIrhnUzMTE
wfyDlJZeg6Vv4QP/BOCODvMEBqM0yegwRoRgsxGKC33ZeKhs95jxxTYvPf5gf+JO6vXpcPpzIRJA
UCRtX9xMTNoSfmAn4Gy94k9Vba1c179sInlWcNIWUR4goJ6I1O/T1LbPLVYdmJnUgxwe7huAveQu
XGKOgsw8mnSkq0kwdUuzC75HhSL7ipCRf7XXx7OpErZWHe2SkakHzyPQ3ytqR7VZ1WogGCaeR5jJ
VEiBILpttkG/6c5YkmDO/hRhR/Fan658wlxgv/pOyOoUdGWhp7jcQYPJdbB7JW/pE+rVCwy8vHp+
laJjyjrHb74rGtSEXrDxnglFI/aIBQtZcd9VNa4HtUj9o2WfaPNC2lMNpRGUXivQvBMHEJhoi1k3
nppJH9fhdwOwrzne0EoCF6eMHQWi99Q8PgAZyo7evfR3L7qUPpQz+Ky840IfvdBwfNelDSShTJMN
yC1WxbvfhYEU7U3qbfNU96OkfVJYozL6aikmyeGY6yd8tUp58N1VsUFDmEejJqGjPWs3qOyl0HDf
RXh7IdeK8Wxjw+j2cOHsYt+VvE/lCSnQcB0jdNGu8C63Sa3OQw4+qohRqz5qofIeIkm62QPK3xKS
pWLpN998qrTXrsU2DHQ+mDRqpEUQgUJ8NgEdLI3q1RPyWk+Da5rCHUAMQBybJTCqMfVzileM2t/s
Cd40PdvoeJJAEkCoIUBJ65qeRouYJx7ZoVsJYc4Q9njmpMt1JuNJzGzL+aKIVIo6ZxiId6MY4+cx
volgHnVgiM7V31H+g+xODarabDSj7j+8mz5pQerIWNHgTT5Xtep4xh/faEJSn9EMqQLO9XKjHdDH
C8P6A53BKJJSvX9XxJOSEUqz5/kldIo/ckYenNDckuynjiOQ8nd9gRNL2l++RCUEx1jM4TWCL1m3
gT2DIUXeGwmYRikV7L3iCXK5VhtCArJAF3S/60b8zrUDwIBqmC0pnlbB2fcrYg88o/We7C5Mbv54
v9hu4hPx3hblZ7fRS0G9FlRPP4w1J32JV3bOyA/5GmgCfXDFq1s50d+ltGczVM0vh4kWsizr64D9
6ZtypPEUVW6WmsnkzjohdeLtpdghL3srHaGXS1DaoiHTnGCHmYJSGPqROWsP0rwHWMxR250mOOHT
Zkq+XpUk14c+pkLZzyj3p3+ENFDCgpANB4oZTs2lMR1eo7PHMGp9M5WHR4sm8SWoR7DXhmjpHTj1
cwGyKrgEzb0019xzrxIUFDJ/kxlovzvRkNi/cWXF9joDQAvW3h57xdWCtrkt3God7f0TwxEquq7h
30IHkz7n0SlcyetbfvBCl1gp8xKxFi6B2AV2x26ud8pg8pZyhMZaQK9tltxcATHBh3Y8VlMPNN8b
5CbA9cWF0g/4Q5T/oGqpAOcP7+CZkJ4liO/kQYMfvy9w8XiWytmhbowu31x69QiQPFHiZnpBfhOZ
7T0fGo16EXFowZJgAWX/86vIAd30onv46sk1Gu2UgBbuwrj7xByK8JML1+KNpSJHwqNGRu8/EfP8
7d21sO25DafJw0fYcqDAdUSVNKwzF0jXrRCwzTCrhTo3U5/3M8Iktn2pZBNdQZoUjivgKz1P1HD7
Cn8njX572MN+FLl/HoP8bMrk5KreJwYp55V5xGNdwKR9FfTql1NH8TbSqOWQVxYkjqKYq4XlmC4y
Fw13AVkcdfXEG6ZznBDSZOFjCPDIP8WU8cCj7oga6h3tUcNnxKkAlk/0kkLWnezFfiOJoOtp4If1
q9UK4nahXJzqlOdAeUOGMfa6+42DRRv60xZ3CB+//jhgbpv2ImtaNLKxoTznJutXaoQD5MAlpwCU
VlU7x3zK0h7IW2dhnlOOO2WeqbjJ5gmEO1XeOuxodIjUYLnWywcU/zoAHYnAWQXKbyXPBr9o/VlI
36NKfKJ5xfDG51OXZiGg1iaiBAo8hJ97Zol1ecPhY69iTuDIPjBnsmKkBbBgshFPRFJpNyxYGYoK
YG1+yJL17QqPJtW+gc1yZnBCvDhQE0rH7puJAXtMFXgUf9TLZjHhtVnlY0Ze+KUOjO+iDGYoPd3m
0XGnk6ai4Zxa5D5xQkxfEzy3xve+ilouj+qIPtlONUrrv7rDVP9dSdz2BMg0d0BB7L0al8Nk70mP
bS5BrepBIOVOMaQ6U/bMKvvi57dyUFskvemWMVcJ+wZLm2Mv+C3dCKB3DQ41BqKYECVusM8JDuK7
vdhKPU1u/SSq0BHr/dmctUynjH5kXIPq57kty74HYXQF0nc3ipkueHQUpX76qOJFIRirGaeYxdxd
Ky05yhp+BBELZhnVl55ujRCumTLG411NbGjYTx00oriXQ+IWHP2n3NqvZwrLiKWUkbl+rQUcRyKA
e273dlZblRW/rMJlNs9j0kAi7aSSf0oGzyIXBs7isXagsRrnnM+7xDWbFRjYGlEcVGkt2A8+Wlh9
nuQ4qMklgydajePRFIPMQ1QYFTmJWsGJXe3hmGcUINFmvbVsl6YLRBhyD4XSkOw4jekP58K7FiBI
OlGWavzcif/S7HzKQ4CVSsAYaahX/6hNSX4OG7fRIq+YRYTq18Hfdn8slRgteahLwzEE+RCrYAF+
DziDx0h+Ak8omG7BiwSxnf0WIOJB/jAWxx8NR+qa6nXIz1iZ4OYIhoktS1Lg+oQrGjnlfLkLLb4L
JLh3OEyCFvVO4PoDNkWUzNAPXyLUmwidhyUIBcEKy/jGdm3ACxhjhKPke0VPIVlaP+T9xpY3SiMx
Am1FkqYLhnq1fdpNnHdWlpIQfBu5mNNUfVFybCPMyOh9XY+HC+IEnCxVlOZ06lvHMa84TzlBF6Q8
Xw++VDoon20jeRTtcW/qUYGSaGkiyekCHeo8wq19lm+Dr659KuLeGyxNq+38iYwsXWzs9MeSrUZL
mJrbhz83vowAs8uCpbmXwaxUsbMXuurw7Nqy2JE/0bY0srMsXE85z19W6Fcl3DQQf3arRKDb/oYX
1fXvW59Ta+Nd6k7bOoG6tRIxMteYV+4fPOJk0+rBznuMY4xs218N4V0kRxfyWh7+OfvnHbHPlRrW
Ds972GBrY+noR3sZZ3FRjmNNVvVHhUvyOdVNZLtmwYoCViFlGxddcXjKz6BIshfhj9FuMmwTpYu7
mTczIezTsscCLDnirLafgCJm6GG39mjhHAEq5At5sqcopgQNjLU38xMczb4catKMoo1LqOikRUzK
W7msGE1H4MZjqz75yRE1A9cEKOxoBlkhoY55IUdmiVQyQsbrCu60jwXufWL2UNzYOCnYNt6ln8o3
+bBVY0fLQMy4VgVqsvcwesxMXcVYaW48Laj+lIkJq0rYzFIkZxx4ygrad8CcIrAXLBtLlB4uieMu
jKy7MbqPYJyznnZd8SZqw7W/uOxhoJ1AdkthlGa7X2qVoAXZompXR72FmQ1uFxewdmCrSdikHrx2
dNbVxx/WKwq8QnEY8RGv6u+E1mjQQcuiNnNeerrNwj5C2Yue3B6jEjb5wPGlinl0KqajmDokbOCn
OvvxWkS+1dsQqqWF+cHUy4jPhL2HLsizFNDvD8tgP9mVm0fs5Hnj+kZWrnksiGMD7kZRAjmpluFA
ODR9OJ03EsYt5r7mou8cmBq93x1d985Rk3UjhtlsY25l2MxHwkto3118NycJ6VhfKnD4HMsDNjuX
r0Ces7pchThZpT6CW9IFj7BKUjdFJUIi+PqRIUncAu/a8yfk7siavYOGqbadQBSQWl8L9LuO7c9e
sUo/ugLZZeenGXNkk+h8Shp9yB21CpoW5wo5+uOX231dCHwdgNTpyG2jH/arCEuw9ckTYAIWDAmE
ZZNPdS/b5FFSRXGm54PvGRBknNFcvzBTIcZiJ9UO6ZuSo01ZhZUFBIdOYJ2paFM765mbXZ4D3whe
m8A60M7oagvM5iy36uFgNjKblrnS4/He5YAqGIV6YK6CE+V86NaH3x31j8a57lXZy+MV0uXNlrH/
S3JMJ3H1+s48URYz8lhx2aa13CBWAB8OynLYPiHG3wVBdGgtFlfDeG7OI8+ZBizJbqs6/MxEJ4xp
Gsfy/1I8ewekwqZD1YZ2BT4kIWq0QU3QjG3Jq3Z8MmWNXhssPI19QDDaLIkYV8je+5XIlGbXwkSd
2a5ZfBzrIPr95VZBVBtS9nDbcTJepP+0nyQIiwLaPzLM7PcHJTIpyRV28npiWcWuMr9z/s5SZ9za
BYGPvvy6r2Qila+XOgkk7ZeeLFXq/urBh/Vl0NrooZt0MfIUh60ffAOSbGS+VmKmCvoY+b/VFwIg
PuWPfoXJ48OIwdGAMWkXvKEsBCvAf0+4R5j0hmSYr+keVwtjlRzJAoqLDip8p7LLNRzo4QUqf25X
BlN3OCFsiKlNHssJbA6XViNA22cujTAGvmy5crBFPyNzGFZ2ArkbIkwu0pt0C/gCYwVQN6rhOz61
9wuaIgxP9obnpS847oePi17dKac3mummqhjC02NPW2bvlCBlfAtO2TpZ97PaNHvklHmihm9mJjdi
xurZQyF/Y3GHGB6l7dh49S9CqDfPFqv1vx5gphfCGfFmRCJAQzcoY+FhvlP+qrPtKDBcoDm38574
kb7TQKdf5xbCLxHwAXznYJAjEllpQY3UOTmYoRuTxIQK0aG4cLoJZETZbCvhwnwjJTvX7QH5msnu
z9MrKzs0F8MFjUpZbEhGmDDwnq8apZXdzd7PdGKCg/yJ/wEbNRT+4I3wFMyL5DtxRic3dczqYdxj
1PUYTTiw+QXWd457OxjLqTbuvLSEttBScoA9Jh0tpY6P5uIBHwMdJtNbfrcFmB0KRBdDlqgfWg+2
nsNgBJgfLOSsnna+zNXvytAwJ0jS2M6Ph1S83ZDES91kVOyZl/l32DXB0OmhFZigbnPyZZkGIOXs
0h+D34in/4GTqWPzmhl16Vne/uDFPnv4A/TCcv+Gq4nAOIqLUMQBgVZnO3LZZG45LS5o2As6w1sq
Zys89T8zyHgeYhKaGBrYdHe/QjTpTV/hCL4n+K/jpCFC18JDR3nbGwdPgdkxyQzNb0l/1m8ut83Z
k0MgXTGhx24/P5sj9RFZNPK4mPfFnAjaEDI/oWTY82Z8Jd9Sz/FXSOD62ft/DtF6aWISUOhJ4OOk
4BJoVa1oZkcTYtpKPPeb0DVdN4CUjfD3pt6Idhh87KIcfRFdFQCALv57TfDINWgx1ru+XIzeRPX5
biOZC5H8iAiqTxX5aENXLndmT8lYtL4gDrdn4J/ealG0mhae1Y/2bbvcOk5lxMEDreLI8RYMOh9P
c8BslUQFy1+Dv6/+AoVx8b4S3LPwc+lX9JG3xYRG6Ie968F+tqiC+ezVOh+U+7mQLXkkpTLseMpo
tvseM/XGiIiMWf8L7p47komFNTaChsnZvIZPz9vb4CQykIrvCduWXf5DKVHjNyTkSrveOhtaaNg9
3BSrpgTDwxcSW1MISqz13Z2rr24mw1Gsdj4XgVrGXy5RkSS/q6TkAd7Io73PYD3WvOFUGPKt3q8Y
A9TwOOIA3ccTtBtfWx7WPBZlSURT23dbPTUSiNHNqVNZJOBj4Q38OqHisnwIIPhkEJ5CzBR1ztRA
BFityB71YAp5TlLdfyC8FG1ViTY6IBYx/g/n285HHHlUHPleGhMn48UB9aDblcZ1dzNphMmt+Goy
48Ffx7/AVsjovAyICuQtsE2EjkVzLsN4SrslHZrXGRf8WFJkqwqNWiJWNtTB5CBYxN+HWKDfU6q7
LKsfeOSylEMTJumaoTDnBYGPt9LGRBlxkLR80wcZbCxJJJCIk1TSp3zYAssuVnoFhDVNtR16Za1J
yT/+BKD0vkxAAr39oEfYGwb7LRk+CIUi30CI3e96WMge89HejiseK/Vp/KaKv2jbV4Yh1J0M+uK6
ZwKTO7PGPYBpvpPnp3qa5AdWxvjGLgGRXWtPWFZc9XAyTSBVZIuSdwkvjM7iYPwvXw1W0cZcVNe/
hWwjMglB5zYJETiRpds5J3UtnJkSoIspAf5Jg+JRpL2TwnksIhG0e90uLS8zsKN1ImiD6vmlOFwf
mrTJgbhtRfQTXZfA4ArtmRJnXN5E1eDH60YvaeKdVNE1r9JQ9Ul5A9zMQ4rqaARulPwwuyx1mQBE
DWhP5BhN2PkPbKZFNz4lTseZEPd5OYCaFWdn26Mcq5KssTKm1484iiqhqyk15QpylpOkX7nBSHEh
i7n91UUQ+NJrrCaldlEuWLGt0qz/5dnMmbEc3JgKiE4Xud6nSSdWDpP2b3ft3o7cyZDImwtDSFmO
fMx/GvzNn4ad0JKMNAT7HrCCh656ovvoaGZmP6btU0jzm66X1pdxNfVvmAmMUk8TFRtm6qZMVXva
TaTM4SEuPLFYKNa7hic8Q3d0/E8OtD4byHZPzeDCWdz8W6ana4z0fOOKA6F26YL4hsKAbtTRxBfU
eRIPc++sgBWyPfYBp9Ymh6cSiy/fgW4xdHMVJISCrDkA7pocd1301PL2Ku00rO/wiFZI5SHfkD0X
5fRaZNIA6klwXImujUdWWN7WtMyWKHSTElsQy/IcrbFLTQFyEoBczbQCP+UdGintp90ShEMPx1bW
WzGbT7bp0dwwFbhdGh/bfgWoJhiAhZuHzKNWb9t3y/CGcOZoyae0R3qRDecysLtuI5oRpqUOPcKm
F3jvUmtVEL7lAs6e/Cgruioq/Hw3cKRmhEbo4zQ2KQwb/pBQGdPn46/LTLDcCcFMZ34l7NhM0Ozf
2b815aNROCMWTUl5AcipAlpCMJ114VQ9ZSt5TQd81oVE6sqhkC76q5IySHyVZ+pIfv3nRuzhZaaS
RJol8oiG3GFJQwxmm6ckaRoZE4Rj/b77fAA1r+3HlkX+1tTjro9TBGRre84SXkyZbY5kHlGBEnXP
xDxlnX8cFSKoOdyVsnw/LoiXtCPrzdD4hxaVgglVHZr9z2bvvdtpNdEQXAMHZqjRjNPAzAAFSAVe
ci9TxmqdE3pQA4jtKRo5W3B3LdHBSRaWRkKlMD234iimyeQ2Idw7Y497w4X1BEuCqTWYRfMX/UEA
Pm9dxBKsiQnXeVmn3StdqYQsdNGeyfzNGsWJTYS9oERqUzoNrwe9+pix7bo+7ySmP0iS4SmSKfPK
UQmp9DSNES6K/4uK23rX4cR5XvD+uH9pnLypJMOx0kDEvj/isLHscW0aAS4VSIGuCJHjJeGTgefd
lcfztTtZfHvbZUYNMUDh/eUK8RCIgyzxAFvkFkvknKr00dwdvqoB3ak2ytuaP378mssz+7mLsxw5
jfYti7GJZ7CYY+iof3BddoXXWkl1MQRO9nKl/GgcGNTtjt1iqtKuSRx41uwWWyIWb8KGgVQXm/tz
yDhIZjeyXCP5Hon2rTb99gnqimIiaSdvKk85VV/fOhoGuoJpY8mjoZ9A0fWL2V5q5DeCTvsQQ47X
Fwr66xI9+2lqJyFa0mabCSV8sqyQb6/BpOxYOGsuBPRF8IdXYtzVu/ICt5CdNTspxuhjS6KOtQYs
FsO0BK2a40J/iamNZcJIZRf6tS6Mg/LYj1HgZgSdtJiZgsDWTga+maARLDrd9xhyRnB/AFs6Gjt8
iIW985oDeJEGhZ3h5cfKVbFhgSjxuAusdv4kkM3/g6oMzIk2YHo6NrCNWu8275Qt8jmG371ICurG
MShVjc3cn181pUWWKMMhRm5r0rf6tocAWuCxMFJBjx6/I1z/Eb4rn9T6EN9CHRcMxr8QSJ1BHUCQ
guAOgEtlH2WMc7XLJEBy3uCkk4tFYIImwX1VDARZ4sNKf6KIGj9E8KwgxTkJmCxAccp3VHErRYog
r/yKDLurltyiMT+gQhf9P/BQSzalhNoE0n3ncTbVrMXD3ks4cydIgHhE88pwtE7ZH6swCrbW6kx8
AcO69n73dnC6vOJsYvj0Z7vUCB+GdJCMvg66q8eU/z9/pbKsPTb6LXCDFqqY08OrGvTIXDg1xeFn
XMAmkg8fOERk2zqICXtRN6rWJt6xnbnKuhjFNQtknxcuFkZwIQvPQAAZCbchSl4Kb/Vf7eczhWkO
43O78nX7PsmkH7hpdi47QyTUyUCzJAjIF8GT05GGRtAvoYrCu5WSvgKZwsNgh4UDDSO2CcFvTxis
2yeQy6uc6Ea9BuB6k/vhLfV7pLbuUVDk90ZIDMvqvUEfOPhSWtKAI6/DsQS3up8CM4MsTehm5tzq
YmiTYbI7Jw75CZZ18dJfnfwq4Gwk/0VWmaBFXM7LPotfG2+Ae8yuq49ih8/ikdqaJMbCbhfX2bKh
E4m+xo97UD1KREJxLv8S/jLL5cK3PRLUdvLEZEL1Lv83/Sa6tMjMJtc8yu81PQrhnq3RNJkNS3+C
Kh2GNncq4kvVShHTRzGtaGOLBq35ihqhnfeGppMRuE0tzTPjlyJtDdAUnFLvQWrNU8a/R4VqDaMu
buQGwFuX3GsSLBBcDP+eXbtkCuOFmTDKoeamBii50qHagIJzJ3Tm9snWvNXHecWjK9KzvPlY3xu1
/QjUfIWVuTvUEb2BA55Ez7IQSiBM/GrFWnl7iyFx5TFDIywcxEqSJdT+Ti+VQrMJNrGw8p8OIF1l
o0CYoXKKRuxRtFqckcp0iW0OHofzDB9niYUAOQlRvEKjWNA1nKpCoKL0WbdQQim2CggGZ77dRrEq
Ts+xUkW+u3ktgqAWCFGxJS6o8bdbzAbuTiJRQfgvObYmRW6pyMWpoBu84sCotHZbSIG8CTYDEVhV
DQ5KloZx4JgVKNo1rSuUcjsPLcw+CHVOSvRaAEOIzP9EanARPmqggJkGg4ydwhr5C8XuXfvl5wDM
2Qtk34EUP+/QapYpLFkH7JFPKqwEUmWiS2nnVslsfE7hSvrRanDPkSCMMD1tngM7q4AGFmMUdS31
LGmIYLq9gS9MHgRQcxVFVDbX+jQ5okcsOCIjxETQ0YfgNn5eaRbQlL3Gl8sgZ1yptF9cy/AYLObG
et5s542RfFL1QjX/OfP2d5JASXn70T02o42J5eVihLm2rqiywWQo5sOve4Yl6LJ7hEc3l4N/3CbA
qdTD/G9EPM1Gmwm7GhG2hJmOtwIqSZMmEmzN+8nz7osb8z4xeHHgppjQdZskgyNKEz8eAVZgSb/i
IvXN/fEXQ6cyGOA0wsIEimcj0qPqTpiHp9pzdcl4tyRKAhkMRETVLEKBFSAuI2WhaxgRI9uvxK0X
1+PAWjOPIhHlmHncnMDMTkeIi06DNhgdbFsroWeFJS08QuhNE7GmmCrEkjqkCRbGS1/IlBOskRvh
BoB0uPSOe2Z1W/DeDAkZ31axUcwTLqqUMMqezRvuJE4UgEFLVyz2JsBLu221RGKDRqDw1SLTor1t
UsfC6KDxpR1/RSyRBvDzzCg4XhSQ03QVnvLimR3dG2V7wtl9MD5vdXPv9ghgFtf5HAobGGAApk8N
6dJOhBi0ckYQA2C81bFTS97uqaLdJN/Rb+sBRjdf0AhCNWHu3FXQ4CJmh4JCAKgvILP1mvKPAFYE
/eaJYjiLzTve4T6Q4ntj91Y+S+JvcHC+hOa49DbErss+PRzasy18sW2rsTY95QoJfiKrDK7A/jak
tAP1tZc4gMH5+yKRH9P48AaZFIZDo+IgXrJl5NwD7CjA1e4fDLT7DKKhvrnaWFIsTo+tjZE+c2M5
dn2/J1JrZUV+tXE7WgQqW0+1WqHFgzktjGanMAAs7SIoMXLnYbTvPc1Gf1hEPYYCgUp3osKZDDXm
kZzQOOQ/l1QNS7wuyBJTlxP3kzEJrtLeNkL4l2mFMkBLDBmtRf9WeDG12jh+BKWGnw4Nu04ahDLt
LAMriPatrosvyLgKeIbnGr6IWDQuBjNUw20DPN6Gk16urNY9j6Y5ktQrxNglWThj9mx+KxRr8oK0
m9QLMJq7/M7W03/hQTO+P/7Jn4EBRWRCTkp00IaV8p/3s3Ewd5hB5Vg2aqdLq/tC5acXHCYriazS
3MNmB7ZvoTYx3TmTZiWNiGeYJqfyIXcK86RyVfB2ptB2Fl4Z8t1vPkp6N1QkNbfl579f5gGThH2l
VYz3nXgXGeoGXRYVUc+0/sJ+ooWLVqjsW0OjhnB01y8zr2IBgPr9fGcQOxXfVOmbOYHwuLPn655a
TrAyy5t02LQt7aYPfgTV83e2DitiTOJRXmCRbIPejGasRCdvYWC4ettcw44AKIkEXCq8pH/M3MXQ
PxjIFpkhQmP4Nu4bZKcDfTVg8m+uV+hDC72wjHKHf9rziwzEFdkXTKLBXK5ABeCUQBrHIS9rgSUl
kEYbHLsaO+Lj3fWuse1ZJ+8p+UvwsSJIHVM/X4IAI/gJL3gjG8nQbh5MIHCf79VUaKimgEyFgPWm
TdBwys1Ohzfqv4tEmwA3xRnMEdtiwnHTbTeVTbwh722zvAYXPsSclWp9TA1NX+94F8fi0guVwxF6
euK9UCk9bZglvFBUVaqbQ+Gm6o9JuEIUJxBGsauOcrPeK9rQcXaRa4tPcFmMeSPAfpfoBi/n177S
TNX1MSpr93XkyUdRu0XUd2C01eEqXM2Ljl9Cy0fQIp8OWKem/MtNNW7H7mRZPhAf2823V8r44q3z
TV7O8kp/X1nUAksdxeoIyFkC76wlulLAQIjuZspLrGohbAi6TA100gG3v44AoMYSGZpXGpB2j+rc
RfDqLIc7QwIUdxBNhTvT9BLSeK9mCKmMtezHpsx2Fh6v4OUfdbAmBvs6sCQ3tUakbyoPBgNhWkP8
EqeG4TGZxxamEjBF/pbldFCyymIGZZ4VPQ6S0NKXcelQ6/1ucsHc8d7yvqalaOUwoRcyezIGGtkx
L5iR/7q3aqnIffW6GEfEJ52PnPnepfKLZLzDbOs/ZGvR9qm6TCVbxPbxj0tg/ycywpQhDcZnUdEI
loLd3f4mI6fsyWKcQP3YqbpPUakVexCO/uG85F+A7XW44zp4u8riQZP0uijLXaXyRzNVujA2nvli
hjzy0lzChZ13J4rzrKobMCAA48E60QEZG4Am9QNLl2uvejVaD8kY8OXdVujmkTepSTgV7MTM35JT
mzbIUyM9OTZ2jG9//oLLVvI4bHTqnFx8T4vaEvRuCZ6DQ5NKKBGyf7hr2blrJaklDFkdAJmD3l3r
4ujweB6vLUXGYG9shtLTSYbzqqxVfskuQkMqCrEQ+aDKlq1bXW7PZ/Sit2iAGZROBVisTzm17nlZ
pFNriwcAxtQGkkfO2j59TKADNK2sW4Rp1dfRoEa3U657VIRfOHN5/Bju/o3GxL6koylVNMU42BNg
zdeKTFhkXCC3ZwaBj7XKpjFga6rOsVF97qb5Q1mqLFiKdLYUE+QlHyZtomVG0r/hukI23POugkwB
y5a+NbAkP7AkY4HN3XY6ct2EjsWlcbdAg+0ucN2sG9eII+eJBsBTMGzvkPBzwUHoVkelyf+2PbZI
1FPNQbLdpAJKZAmC3Q7JtqkDTYsWen/Em5lVAigzGdweWwbr9iHZiKaV8hFFbvG0/3dcwzs1TPWf
VVYTkwLMgy/gQo9jBvjf6w/oHl90s8KyzUX1s0prh8Q+rNsV9Z8V7TMq8aMakAVY3fa4jB+uYOyV
rH913uxl7L0hOL63WpGIv/HyEVUaSzbhRdGbhckS4dwEuhzZHcGoNaXl/2Rr/UHGJB5b7vUcLI4W
twJ7MSBenhP7xyfunPQIIPoHMbnRyNhoUDGNlEDxhLppF1g+4FaT8zlkWJ4STp9MPcv8D1AayJ7F
SezIV67fXJHFhQXiAPLrgOEgzODLfHewSsZvdskkx9CeipK+53Cxek6TeQiiyjHx+EcXiDyJN49G
gn59UOYJOL1H4gA2ZOcXAs3vfsnQgQFdxqnvGLnIdiw5rlbLXgKTGiqIo+ZlvqdRf6Ff0jkNm8ix
07eh0Pgx8uD1TmAf5YNLxtati9R8eSJOjUhPwM4C58hl31DEL46LQtc1BUmXVA4GrY05bNNIMB7j
MP1/GMQ3YNe4rX4m0pcQhH+4na5VlD2RaXdHpja2hyyddOunOQCvcvwyooBwmwNEpACpCmo/sCmC
eUONfML1GyMfBtNfWadf/kP8RTnH48AqAVWj3Qhe1yLEjDfK7wqI0b1ozi3DwaJKGjT+vyXgBvTl
c6SWhYF2IcvkrgLdyBXclmJaSR6qF94x5HrTtB/1JQOzfGaMYTy0iUFMA7Fm62Cxdbc3GkR+lnYK
KfXsEVdoa7dqyCuzW2VCWH7us+ISLXWWjVgU/jVxtz27Hz8jg1qYkbm4jebuVCcUYrTuGTjbdB7q
ySLFO4SGSpQFxhDEv19gIxbSjsxzBFkoA3fZJafzR2BmUkZhlDaitV7O/umVOHaD26Qz5bPfjlCJ
6IbTPNrBo2oyY0ZxQN+IVnEnIZ53wxU/lddy5IBNl0SD4P3hFd1sktgvbs/QC8U+Eksx0jwzIKTb
G1gImwK5KQrYdfcoWQbr6kNm6jdhA65Ey5pDA/82N1KsJIvEpjX9+7/nix+IwRkOdfapJPRvJf2+
MZUpG19XO3o6sjGHRVccRwHhQRfIZyJyf8DdiRQ5hpMLH0LUSm/TxqUS0ygzuwTTcyE4HhbxSUhq
pzfbvLy1ew7yD/SzwZongckdM3kiKuozChAqUkAkn6Jd5UbboLwNtbosHu6WF1KGesztGrLNJXq/
Lx9sPRqijoAmgCesiscEwQN4A+GGRBShuwM53sXmJEum6iiRJmCYPShtpfNHo7OW3xDmSVrE2ivc
ofPD7GCmLVy5RyB/fRlJZJ3kZrzNokelCAYlCsNNU2SXmP+XPnwKVDnpdPCGMemhq+GzENAGtVfX
uAFi0CLWfU+k337YAllT3ui7u58NFXVeYxTrcEMxxG7Bczj7mPHVRxNoCAx1hvH73PZssHjuhhJM
GBhzZrvLV42CCXJ4KVozYO9CpP67yjfA7HWsriKkxcJgQPzSswC5Bb9YQuqyRH5msIHagiGQ9yY/
gpmRC5ypn3o6gRHlAHmsqU0Oz7k1pStA8BKVsZ5YLw/LZ/OX6AguFkR9f7lHRcoOmqFrBTIURxyq
3C9+QniPNoQz0eF2CKbsU4v/yiB5Fl+ibKhqOc72qQfOJXpPYnh57V0LuJOMQNSzBNZc46Bu1BZk
15E3w+rXFFgIX8kCSJU2pqGG0Mm9X22MZoRYRmnzc+HmgepJ0/nnVVyCYlW7HCOD5uxwPTnCBtH8
CcM/f0X7W6qCxjHZijfWyUQut6bseBHyY1jNDWQsivWFneDRTJt/fg9ivkWKQfX/OtPO1+1SildF
DunWz1Ua0qa3v/kmFvpYICsCh4/AjJnitUdTNjqwwH8IfpOjKka+x08RDuh7nJJJsjRRJi/tY0IO
+nT5O36VECLSIrUZqtMU2x+LA93K/g3sKI+kBQ/DDKsqr+xPviZ1gP+TgzI47NPrq9248YW0s1qX
oF2zGtyp2mNXAB3MLw8F37bK++h1+5mQWIs1rvHtSqkqRvuLflw8kIrESaFzhqmwVJo0uO5nM3E5
nILoKycplv8O0UbaqPysAHcwjiKP+5+OOHtC6CIrToaxQrZOlhd6xtAuNH5A2pQDE9j9zalJ9P+w
sQNlspig3jWJZhdLdcyiF1Ho16RDVB4uQLmBw96ciyGAj8pt8C0b5i35YUxUitSpcPt7sUtt6m0J
dugMyVJmtaNb7GFvFYHSdiZzXwTFmcmYpqA4IHjzw+yO04oMgIJNTfH8TQ2r5LSo+kDnd19jHfDq
KQ9orGDMIAK8HCd6SM5im5XBW37ymlU53Agz/lnDfZwlbZireSVrPYe1Q0wIQ8mcMQVdl9IXzcFL
1eZOcbcAvEjv/HULo/M4BTxHmV/UIWuMWUlYTNQXOZEJkOPAkrJzW0z3bEf4WYIaW3aYx8ZH+KWh
cTvChuzW49cA8qEaipqgNZjpKEaTiGupOswrmIh3qtalSwDgS6i1fYcpmRHrqjcPJNtGZdOpEdEv
tJfa30ErNl0AwbohVLg1A1E8iOGcncWhGdwSzbIQ0Tb0tfMIKwc7igQYfU3ZCl6VqtDbw1q4K0UQ
FbT6YoCv71ZNxzfpHKCPyVoj0jr9v2TST3bi3T46ePogudO+/4QjSE3VHiOiXUBusfTEekzX8VmV
6DC1coG9yYlUvO9DliCrfdFUzeM2+tXITUzNtZbrCsZTtlYaBsFLVvDDUDfXBv3UYhUofuZoqmc5
eUwKwn/7bUU/4t7VOaNlCBIxyxnSngkx3OFKAPNGewB5d01mLlNzKXASGUnpsQsLE3drL3ZLyIgU
tiBcpdUnKIEsw8UmodQk+kXzo6lVTiMoT3eSrRR7XImGN0TVnhaAPW6PGI28mFQhanSdtykuBaKa
3zuRnKtXECGYfOa3NSIw0tVgsRkAfJRHvbXs/UA/sDqHQKBqdihoHIx2COaNXR/lX5suYcRrwXCY
2FwUOfMBZUCmnP5edf+uIyUjVbpngDNdtHs0t94yZwhOPMh1D5x/X0Cd3EkxhM7u0KPOmhPXoYPA
F09pBVYZ1N561rS2lEZF2yUZOePADYs4XqRfz6f70b0pP9bQ8vgqe23CpQF7OAUHndegefDBhV+h
bCtotQc1Bt7202etHhYkT79x3rugV0luizBOf4ivM3D82aB8bAQa/2LMJSzGY8xhTcgR1sjYB+WI
JtUUS+mEbbcl+5azWhzoTb3hZ21QSfSLrxposjOgA7ykCij3EPSGCmicv/wX8WM4ndEci0UX101n
pf5MLvDlCHA65iClpUcyztUL1NFZTlF8p5PXz5LrM5GbS7ER1S+XXO0whDFb1K7gnvuXATtU1GuW
3EM1904tX1ojuk99rqYfizybJaj7Zag+fLqMt2DrKxq/paN4A1CJ+CCJsxaO7S6PNhNv3fRjW1jU
69morPVj7qNrlJxwUQZCD9AnGUxJZpnkZfvMsJ5TNiRtqrttCQf6+4bSvJ5Y3zA9ASFK2D1isfr4
HnA63Nfqdtf1bn355hu/PT2dYmFYoosYX5Ap+3NdXAeplUq12r1BL1eyJ1IyF5sonH3/WW4Db1c7
qRV3dgEuqV5N83y/TGp4ZwhVRHF41SQFO7q2E8GSt+G49Zd/0CMniiRFrdLTmT/2WmEdtIppi2cq
E0QuYMic2RKgoqMJPz87NCLj6qpQYe06INta/K4Zm2BT+hLMFnn78WZFxNaOs72STyWkv/NYRfXZ
sME1pKCzU3z5OtNUjGbci5JVLiGyVOy5KvgQdbN0bwYoz1Z1QjMs9HEEg+gsqV43+BViKcgrcwHd
R59KpRZfH+uppRsNO8b5IuEW/A8lItpFAbfYoGJ1zVLuZpI/RrvJbYVEtvMjjZPUjV5s5hv5i3n9
52doeJSGCos7KPmutoGoccxIJCpAT1SCW6CEuvgrM5+YM+FQpVOGaS3yCdWDSEHKjjLE2peBm01O
MEnR59yamPV4Lo8bvDBWmT8OmUb7kzM/wkx7BcSwaGt2R/3kN6K+ChM2ERR4CSMc9E1SpnEt4iR+
/6yYFkV2capit6HeG8Vf0CBlL+i7gZ8+cse7gzHx5AXUPNjeENyjUPuZvONFSzInUKb86hMwa4xP
ANLbWTfy9TqCggtgxmIjfixqVlyjEU0Mia5cXVbqV1TF0S8X4uHlVZhNc3Q23opkpSoV8Q6yqoDb
AaqXDBtPMBJE5H7gJMAL8/vBIfg4fviiEoFVd6Nf7Mu4AJrv1UrT1MQ87z6a+rFT7Gy5H8PmxYoZ
KAH/U/x43FF7+QEGpPJex2tbCDs8Fuz6ElWcpQpNNRWQxyd+KF6hjUwaw4I1W63gUzlG3yxaEAYV
dunxf7U0YlAIkU/BHbiBcoWi4H0A5mp9x8QnwBB4LToP8l8ZsxZnSde3GZWJuH0MZoD4MSGCCsIc
ClaomCLrMyIR9iOvJEVEaqYLE3Z1RedhE6Zx8VhoxlrFIOS8Bjp1qVqCXo8jRM/I7wW3/zyd4Z1u
Ky8RS20dY71za/emtqyB7F7w7pSozY/q5np/A15L/6l8mdLYQ0Wek+z4Nc0c0wYZTEHF9pbchIr/
oJ7k4U6q1HaR6Vs9OTjje8PRSgwzA+m8CwXUhSGYVrJzP/zhWP42ZAaMDxG7NJxZ6xKYAYvhbLFC
KwHXxqfstuUWHHnlGm1Hm5p3NYggp1TX2i5agtl+qRLIdWDFy5Vr+fEiB6sJBTTXEfDNPggYtlXn
p1Y6XuuXXYnqPBeOdtF7z2Dap5DmtshtFLBm6p//Rt8oteMOETD8CBaadcfv9zoVegpb6rVXk4oS
w/51rODLPbs+6Hhmk9kZOYhRmPhITZpZW0HzCPDcdQO7DYoBxjA0KSZVEUloI8ZMjXZ7/Mihg1pG
ZCD2sZTda1I5WqeDUSJRxgqYcwNmsVUHU2fKN9Q1EPe5rhNQLNqGW7rJDl9sn4ccnVo2QBMunYiP
m3GM3La1NV+NU2nlYbswHXn6ojWH5myThhQuN/gIoDLqXy7TDytqgg15bw3Tyxt21LbxSzaO/GWV
7qkjrDxaFyrBL6CvqwvY1AuKgzDODveAP3ACDFEC2KmBq8BiYzpyRKDWkIU6H3zhMQIJDS/warPW
mIBFbGgi44sqdAN+ot1Ks7PU/BuMr3yXk3T6Hc2T1xOWkRI3OIIDqi2xkSbnfMnrfItRsRhF7264
ly9WFDq3nstIx+t/UFGinLp+4Hmw0P/A+8N2pjobHftORoAbwVzobHLKe7jcklc56KqIPY/Cn2KQ
tRrDIE2RlTeYTdt+/4J779LOJk5Rtj52MUZ6FM/6xWu/Qxy67Y6pOmKXxbfQ3zskdcuDV51fQnG8
EUYvFnosbjfrdSCQYGmp0dHXNPZaEKlmiK839YoEuklxbRqY82FMlBBjRJm/s/hauTT67Unxln4A
YnHznWlwgZ1+SqY7neFeatRcYFF/jmrVpLcLKcyrvh8KbcV9oopfcPHasow1xykX3nU2UhRXLFRn
Am+zuPHFaNT+Kl4/+YbpQQCjB2oECWNI8KR9tJpEdZ5uOS96y7/gzdWhR7Vr5YmnHhYZrvLcqvy2
Hz0i8qXRDzJjK6JLYrfAXMS0TE9vhAC52O7SgHGsldh0m8055cLWQB/j0fP/2upIroB7jW2IIftr
pk1HDSrLUQZ8Hp9EUTeAiXhpkQKowrsDxeTnRe3o9RwTGLmQVhlQYR4AakgqXKe0WZkndt62cxJT
WIV2V3zRpQou0myXc+UM2/nSTzLrfQxNQt0qWMduBZ5JKiIpN8Tt0bQhdNi8VUAovKqIHHnKV68N
PfRy4JbgV5Eee77dQGXoYiTfOX/MR9FGwBSJgTEKIEC+TBmNaQnFhiYilIgYdI3Kkj/w0yPVEkOe
f1HU35hqFFwOa144asY7U4XAo9Q8q4FrtTjdYkbsjpfmKJUL3LZMt1RTMqnI+MRTDiR1icZZHxP7
XpAOv3T/8BznmJWj/2oYGbcS1hyZqFd6OL/jOqMqdFIgoYfpscFe1kZ+ECKYp2lps492xf8YOc/e
NFP6ABcbHZkUzq8NvQwFmJFf0UgwyaI6NFC3JvzvOJ199IdP0KHeE2jKhEK9umHFLnKXP6J6Mh1j
2Etr2ndfo6CEwIdVhTmMLgeljcc6gKzEJm2viSpZdhT+AoCWtAw3Nn5LnGoPOA46aud/k/Zu1owY
EjCRYGCcLUTeogHe+wKNZH0XjGNGL981b4rfGIc+U/yO/BnsDfHwvtoNHXpQe6B3KFFllBcAtWFR
Vro/Hz6iyes1e6Q1OSH5SM2jKtAnc1JQoht7dHzURKNUlisUUylXebYXlvW2WLC4HMNlGI4D4u8q
XeMWcV4FxLgtqlzmCNkryFpkPmvsjnh8mmmb8GeQ5sLTbMOayGlA2mHYiUp0XPQj9JLq6eO67G8m
M6bjByen/ePLZ0ik65315tcyD1ecsqH3Ek71/0KbFRkMmNhGfMqUTmvuZE+B3E6wGUHCLlN79hoT
SgiaH1isxJZShWKPkVWZQEfq4vaC7eHeZ9gqvMyrlZ07woam5gk9hn0JloTN1wuKFkjOzJK5B/n1
LTBhZZDeekCv8hWsvwQ7u+11kVrJ05bylOUep9MgkegT6xjod7JqtfG5hEFsYLmBciXJqbN4Q2qu
lpNhxmxFVzyJhQJ8+tXbjUSl2ZdagzodiB4o7cbDMpkk6YYHlXETGjhx74BQVBM9mLwUlJllX44h
wAEnRfAE5VlD5Rt4PKr69rMTZXl1WHc8oHXtd33D0RT96RzjIeE5QcmRGFD4KQIZq+bripKhB8tl
lZUPraoNYBjjllt+TGgtXKk+/Ng0Y4HKnP2jyY3ScLas7qt5xl6sqR3jRg/Sl5KZ51y9hqOv7nN2
gdfwevXkFHS5iRgNEpRsHdQvUEZlQ8Nh/UUd3HGIt4dxIM7oM2P9PcwubMCsiqLjEVAha7N7Jv4e
w2bD/AWbSlDjmE8Ien1OoxiU4k1Qs3AZnybrCXDfCKdqR9/m64ojD7lQoH16K4ymeCt3HG915M4F
WpRyJbXOqqb281y7CH6/B2NoXuxpwxusZkZ5YXqsnMzuuYEPNbZyHR9NqOjqzwOdpbmN15vqMxjy
1bYgS6eoQRdfgBHdkNeYjluTLxxxy2dvNMc1PYljrkflje+XGIBxK9jyxmR/cTZWccZIBvcyrmqD
WICRmXpUo+rSSSn0tCoZYVF7XE6xX+cEFFGc4ixKP0QYP36gYho056UiTpxhcB+EpconRJpGDOCR
MCxLTQ4fc6ZL1LJG17cLBLrCrXvk3WBRLTgWVath4togcW5TnR1LKBqojoP/4R8Dk5MwWLYsKZMK
CKXF3oz6djYju7fc/jsZOmNIDNAmoQHxTIvb6dWkWX12oBQ1auwdovJf8PZiTkRiw28ZYByA12ou
SHWL5uu2ONTrl/NcNj8AmdzeMFffl7SBcuz9VkIYl9uXd0QW3rBWw1pCc1ad8YwEEE1uaCCRnJYR
r423dz+0yie0PkfawwhUm5+NzBCfRbWTNFKW0gf5Zk0c3r+LtRsATtGyqH/H9N6PzBe/nzT6meei
j7OXbPLFKvWNp5OyIoPCeFR5M9Fu6LxAXPEkj5AmmHIVNjolSGFgUNU5DodimvrNXoJWvkSUPO/h
snn7U1DIcIn9GQdMg7XzNCb5PZmBEU/MxFggNk/pdW7kxDgf9xSriqXRorpoDovidBCfQZkQ1cU5
hgIvaEG++AmJD0yBXI5/eCqsqsE7A7QTE6bzQHYJLjLzH3EDXhyndMmJLDdHF4wMtlUhk3X5yDYO
XRlXKcA1p6e+d4C0VFSm0HCjR7RGCxqwRWbA7VkHDkFW8IVYl74TNdE3pV/pjFTmOl4V5USqCMEC
cekbkdE//fUVMnongZyWrDE+tB8wEnyIv2thRZDHQPsAIgK5tMi00jq/FdFS/zWvnpf6siodl/vn
anXl56S68sqYda1VqoI+ZFQjT7qHH4S7/Qi/O506rHFSkwZ+ebvXytb41Xt+HgCIeuS8DpQBI/OH
hTCARHzB3Gx+0Tu6rtlnuvpwBRrzk0RYCXkeeNOu+exu5ltS3UrHuJIn/qzmMkvNBX54s1cflrvs
OCeCGaFea5y0ja7lV6aZv//PeEaz8nAfbMTPrb8KH90+EA/oIGCeQ/pY30yn6VrwR7gTV6K/+plI
nD7ZSpHTad8iPWYTi1l9Okb2Fj6TfQGoZKYbnzxl+vXlzALCaxVtxbF5m39c0BsAGuRFWiNQIOFS
zGasOTCIDDb1v2z8ikSXPeIneVS6jtoDeeK/1hwtYDU/51EFNZWe5ZttC0S89PuIazRhfqC3p+lp
MHJEeaLJX2xF4DUvn4VXrr+WuoBbqZImdQpEOwywQ+dGAybhhKU5c32e6gwjTg2lUYcSXIRDPrxs
wqiZ78j+vLxYnwCLXpAuqMB6T+L79zv7jb6wve8jJoaZF64DDbYYYRD/aNqBE7MuDppFKEX6JjgB
2bMtbHDr1O9gRn1hSPwsozkyikLULPrjqsKi85bIVTCzi36AaZz3nouZN9AHxKXZ+L4yMRgFH+2O
WX+FQVaUttx5IofpXKohhArhpU0sPrr8LUT/kJGhjOymRlZpZh1ZrAxcktCzJUDEsZMXBtGBIkxC
hTDs0EtiKElyW2S+y8qWL/O+Tk/5QNiA+fDYB/yLJZIx/hdXACcMu1ieTnBfE2StMpdcWC8rOAvB
+X9vH+BWYTjvCyxxT76I5M+7IG3G8qKQdp1DVYJCUzbVLQGhnwpjYIxa9pTLwzrKC7LVQ3e6tX2q
gaXTZ+U4/lqALp6YMnUHG6MGAf7R9rwnrchWPF32cQ9mX/s9fL1aQmc5bnQT4dFV6utm7sPgdbXw
kGh7WfcmTr01REYpTzoeQ5WzVWyCzHgQK4aWCq4RXxSt7mX1EiuL65EIcp6kq42AXNaGigCbqW19
X3DAURxRjHvO0D7OFWAXsrVUNIBkuwOHJXaQFvSWEwKWlZiYeK2cD/xovVx23z3KF4ve53Y6MDeX
ihhmjpm5SkT2kcpKA7ncayNUgaI1fQc4OYngnaruBIXqKI3zwt5hOvgSFtt2mF7bLtLOpFKrTy1I
YS6kh+jfX9G/Op2rp49/fRKv0i8Zs3brJaqjB7ns79aNGBrQ+ZKl+EYnl9KoUY1sQmC4axn2zHQW
e2klHmIlOUh37F10pdiO/NUP4P0lLIRZeYSCKo6B0qwUHOIHKOEphVtN7Qa9xOZwUCifd5GANDry
EZbWibh8r+w9m29YNIwBmVsOwbO1IBvlLQfsGLqnNRg7rKTePqUqInLwlGQ4HcFpH+LANlYHws9x
aDWx0LklMoIs57cF1xd3bS/s8IyH9OFfS8mb7dndH/a7AGlrcyLFvwmrHIWbgUtuRDUHju0A4a2q
zoYHqxgquMA6kQJZPhBbnkOCp3i2eFkwR1rnXl0WaVdaAY0d0k2rhoFPe7LDYKmc2nmKK9wvHASb
rujz47wTX8fFz3fnxJmEwrlBaG3wk0MIhtMcWr14oqkhBlUwV1B5NYmQvfyhviM7RjmXMjQAoeAb
ABwwbwAx2gAUDr6o3ICR1KIXINUbT8cpktIm8jvomvPZ+COsJRrzx45dPLIlskdNRHciSBmGEfzB
Ryj1IwViqoAoilSPghMX8iitbnzYQeu+DKqtaKQTVwNIu1LpsPiBBkSt/17Vq2Nrup3VPmPME0YL
VVSrNxjNGpSYPe/mhdyKBlIkvvSUuWfZlFYCpk669KJgXejIWMRRCX6zVL7Ts09HM26Gw00NNfBi
+ABZ4sSw+pRBncK6fVa+YGM+JUTkDQitC5eJ3wxeM17EJFAK+XG+dkkDAUM0D0Sz+hPS2lL+ltqp
tB244d2ex6Av/jVbLNaUoK2YnkWkwdRVAM8dq4FJjElZZrKgnjssSIMORoo1m2uHxXFMeTpSPRvw
XxPCNz4n4jQIdb4AVc9SUiwcLbYbKn0GY7HWVHOmWV9oh+rY1zLzV3eBx9QyegEmtquH2kUdJa4i
fFU1w1gro9VpI3sFwK7p0fLkK8tMgCgnhnMQego5+3h6M8oec21WuPUWA2r737+oiX7VOpQId8hB
M44cHZkp4qC180lTXomhMPZkSetnjuDDUXFnmZX/Oysa9iQKS+ZEKlNG1M+f5WVyghfNm5ZuLLYg
tvu7CvqKPuRRpEUudijutlvz5theXQPBkAxX0rsHG+FjONkOOuO1B+OHy9tjEqQvMLI3aiF9kcDf
BFpeU3kIF4RZMHhMZ4hlW8GGsiOje5ro90CdL9qitbSZD33d9NFxYmVCBHhmicSO4lh8fa469bmo
9265iYkXi3u34t4YZRvkLq/Id9UQa4PisRdX2Rqnp8LZJp4sRgaNGwgjAKGQlnXOGVWM14qpfIph
ZiLywcFautjllzS30WFwul25RSu4Iq3C+fWKFv5Rze85ZTr4zWC/d1LfMRxsB+WoiYPSu8l3PRlT
Rk76ImqwyTrfL/so1zpS74l3xnNED7ek+ifVVNp15AtGp0OF3oHBDGvxXOlWiaLEKjkXsei/fgTm
Mk6QDJFadX9vt6uFyjIrSQ8aOzRxO0zhujgy7GYwgy5JEazmFxMUvD/384yCgIDQGJyuNAfGh3kk
IVOKbFtSJTPOwswHStCfm1anRGtFQK5vGSwwFdk/iwkpRGMuM4MGPidpqijDZpCsNfgmC1xZW/rS
5xoIH3ah8er3C8xDVmgUi5CPsMZX120WIZEJ0aBVAy0rcgKQTy7VVVqCOp9dD3hzYNGTTDFMHWk/
GVwzTVH90whRY3UNyIkNDeWOUcz4I8KCQRH1y+xpvh+mvEqCJHnJAhb37YKOLb1dt/VOFO7KU7FF
MAL9baL5MIYfp1lZ0LvtVR3K34TMIdOv16vo/DkRSxUDne+aNJ/hZCkq90EcPvXhkEEgARDP25Lx
L9hcj+fjOzTr0xeQcUPSUc5xEX//JJa7ED2P0i8CoqQmF2V4ypBdjCwzKCt43+MojRrWyGXZDoBU
vUNaElq7Gael6dAtthJ4tWJr8QNH7ytXBtdRlBjgfpeSUu1g8RQqPBRLJHhxrrqpVmKoUlXhDeRI
QWz0IDX25psgkjB2Mlhs8cJIcuy7lxn2Q9lflwKULtdehfHKVfuR717TV1ETKKBp1iGyGVm4uZq7
qaf/u/NJavLlHdsOMLmw/9BXZTMbHT3a+YgYDKvTYB5uVotJT2OYynPIGGYWtBfE+T5QnuJgw8qj
jyNrahDig1yeRRJJ78OPvNgSZoItspKLpMT7cnmiUmfygOVYcjKZbbCFvQQVGMNTgKWnephXx9xP
NhzpVKBnBDbJ/cD3grH4QQ+QuSSxo+xz0d4D1Durn/llJO/jyRkAtXNmCOF4P/xf1vKjYKbxjqLK
z9xE5nsXqp4NGC466+NN0VoRfUUoJKIwv/lnqXuxT8r39xauyZWGFSWhU2wqpOCVCGiB63V9AyLX
ksfKW/Qr0A2bkKwOXArX2XcXgoXSWrYRko9MWBS9MueLtYdPP8XJ49+EC3AWmP7LG/oPgueMcfq7
PjVjKNxi4pT31a5oImgZEFNovF04U6ONJFPPeBDQTTZJsjnlHX6NnqBnE3N3nYJlnAcdBbx0obLe
J01q9gXQWfLPDa7wdftaTDmUar7DCNT5w7IVDlNDTRS2REywPrl72ZRTQJLeCjEwqEJlCfHJ2EjZ
8V9iuN//me9i35eXQhePmztD305g2nD3hGcrRALUdpH7hDYjqcpx56eXQtCRA7XTUkw+mL23vVLL
DkK50kML7Jn2VQ4lau816KyGG0amC94rJIOI1F2ATq6R3yJkUaLSKZjl+zL2fVUsZ0RxYz4d5xDy
UyPDs0eivPELDrVnxlxzp3QjMy0UkfDTToIZYIpN4f1wju9mjsZ2jp2tCfgJB/VO6Uf1dVqepFMz
V934IQKKNhAGVj511ts8OWP6aa2rgjl9Xtlim9oxWjPAbkJqi1SszIidLgBpN7JnYEu7z9N2pZg0
w3+6I9eoUGyjGBNOZ/5QqC3nCLF2tWDbX6Mip0Bc86jzARqJU5ngnBJD0RqBDzs2nz9AnvlNBCRO
GchpnofPwiP3gwRKq70cY73z0AJMIXkN6hsMWsvMgi+ATTyIgKUvWSlYBcQ8b87Z+Z9A/qxJES0H
+4ilKUkqqXnN42HfyLrVlDwQPhjyDVYL53NdMAIr7ApTUuoycfSS5a1QzSipr9klcuUEl6OlST8W
edsM4kMIcNdTTKhHOstGd2YDD+nQnrloEHNH0qQCUkrtRE7Jtsh2GpwM1bvhCq4B9R++i4fxfg5F
aoQctNnLp4etYmJw20wVB5ZXItv4f03agHdS3sNgpyweT6AI21+aPUlK6thqPtOBZn+HAHfvHmks
1lhq5Mt/nRl/VyR1HPe6+B97XnqLBDWVeZn1nNSHwmSMAg+uypJrrgGMYLobIwAX42I03I6gP28+
WKAlVC6AvQcfSzO1BSDdfjbRjV0zuG+hJMTtcNwi9cvAVrnJ1hbONdFeLgj3uj0Aj6b7YdIxXhsW
JIAiJYjch/i6zjXzkEqaeCj757ZcH/OiatmIQFUVcXcjfmLET0eFH30UsU8jWTASl0kESy0wYsme
PucLWqrdC1Pfx9b8+vc27Txc/+I6BeVvCIFRpS9CRY32lsggbAS5Ie+qjwCkK0PPjDX2qCRVwWqt
sX65A7mCYnUyWVrKwc7HPgAAb9A2sn33qtpzJNFgjuxvq1W/VKZGHmBQ848UgsPe9jEn7iFBf/pL
ORdbuAuSQ6mDjGNDkf5nZkL7clieTJd5UQINRlWBWpgm+v2kyJCP3rkPQMGTWL8VS6hs1M8Hs082
RTkZtV0s2moDBRsBPUZwSbT3cvkVWx1Mld0L6A3yHCTMLaTPHCBK6bE27JlG69LZwHGcbVlmVpSH
Q0p0ToR8XphOcSZWnmWc0hj93n3DrTL9nUc8KJXTdv4RuESVuBZwdviKEKk9nYiv2x9UytOMYqa1
nCeXWvTymsjm/yfFoio55elfTiPk0JvLbMJORO6kxe9Yt38zmoO3Zwd4JGJKsA+Kd7pBusKwluAn
dQ6aLkPf1CM+AoRA9m9BZAJBDU3hSwkudaOnCRlBHN/XHrinqvWoWbuHt5J7LvQbUttGggI5I3gD
KSW8bTexk4Y+PF1gXryeU7erXula/8vd9zmH8sEJQ01Ce7du6GvktGBVRCqkBkb1qF79W9MZ1wXh
sGtWMMfY4UwjU9zspWdAoU0znEv1fNxYCtO3Bu1uLKbRtQuGyEVc3863++jp4uOMan7arxa8Ge0v
KrKLTQgHLETRwV+jiihR9szDF+07yz+tyaKQ3TAjWB7TU98zY8gPP5A0FhfJIF41CPv2bBjLUdNu
knmK6tQPJcNhO/J+C/AQX4sDg7+6jxdalkLdAW5QItUflXziXxajWd2iKlluljmZcPY387z6Nlwg
ybu5wirrfTxJsVl+W+PCLCGLpc9DXU+v1cIIkeilF9PIIc5gFJsPRzx0Bhur+r/spu/SzGFz5JrD
bHu1vwZGvgS8rH2wJFzd4p4jDZiG3lVQokyRr1IiQ9+iH/VbiEKGoRlADzlZDEtuMuY2MCP/imIF
bITRFY3uClYIANo6x5iwDcedTNVqyV6B4UeIRnA9eW8YmKa5GQqnrZYo2CQHNybLa2H+ktEm0T/g
gDodg6Hp4yjRqQLA0hsocSUjwPYyL9N3cTOzELqM3pF89OA//pf5PuxCF7sSlFJmfCn0dftAra+H
mpKIEk7f/fWZkgCqrCfrhv3isSF/wRwXx04mJDCo63hZ7C5iRZDr2KzH8r6eFFb0i2Ncj15gW6W0
FaVFuo9XunxsyJsF9vjhY9Wl/+KkeCErEk2tgcBnGaO/5Py0jgrR6lnymfE7gZCkubHSR+dvvihc
X6nmFKq3k9j20gLU0+c1wbii7GJTfMFHfy5CBcfcMhiy3uoHAgfacC3Z4yLMB849udjF7w3bzfp7
2FKrRdynRINdt8gkqLIjwqyo8XBRGVaP7AnWewIu40ctS48cXIs+mq9Bg5kNtdZc7cyMPbV6gxwb
7kEFSr7erhvgGnEGMck2kd4o03uFRmCYOLHhH0S1QlVuqJWShD1bE0wrRBRR6mjokm9FtMlGUfSH
JQFSVj8d0y41YaZo/LsSRLGRJ3dS0IGpgJWXhgLbLamTNMRIT5VdIZtT/UgZUSU1SmBZU26CSOgb
XvN5HoXbAGVZq3k9wwDdGIEDJji5pW8PZylyRptCZcXkhq7v11Ms/uq5goa5g5UIQt8DDFs5v4xk
fG2nLz4ItV3K6VgRotILrl6YBXORX70VQ8EsaEq0+KUduboMNybPKfpzpBppcECKiLsRPCGgARsu
oyLwOmS5O876CqHd3BR5QJWKr9PhN4yKrwvDIhxyzwEXgj7mSwwMaE9kDpyWva64/nbMLCXg26Mw
odKGQYD4067X1uARBASY3GMXzTXFdLmO/c25jFQWIi3kwFME2d9Bk3RCNerj71yJjNAd1OqLuLvt
YHjYhlf1apLAiJ3iPtNICm4kCE5/iMeWNYgxvXeeIgnePUQvPUXdTwaV19YTqRmg/9GNY3Ov6tQE
br8kYGRbLfpqK/nK9FBDZeVDpCbwPfqnn1jqTGOCu3zoH9GHrgbnWorXHQ1e72YcXvQ+qf0w+3L5
094XoktEX4pYCJ0Jg/50Ukij8v6Ny2rmtJWmlEkFdyqUljEn7CrV0Xfru8Lm+0dSUIlr/Kx5kTfH
h7DrJ+BY2ui/SOkRVvrG/X0ZnzjgPCjBpPn9pALW69bzwtPLGk+rNOiLZawcc/H3geLONpF82cbH
uLa6hu0p790dn/7DrajHKG4l48AgsuhjYP9zN1DpsbGVJLXBaFYctzw1oISPm4ieMKsBozn3G9HY
QQFXsVlgQJ/ObSXGWbLp2mAmmSqym5iUhK8jj/HafiuRL5lf7SEn4j9pBH7P4BA45Tio+DFj00fM
DS9uWEPuKkFcpUv6Q7Lg3yinea9KwkZrHgzmMjIj63j9cVF98ZwTwzdW9AYQ6knhWdlWiolXXJwW
9Lbmlv5Vtj97EWLAwbdiWEyMNpCkX2ETzuqHqh5X4RMCRsTCJA57xILmgD1EfjIeU+DVtx2xIbwq
1HZtUxct+EjG43ScahA4eYMNiJMeUT333DKSqs10Ll4dbqueNgHGC+ZPdqIfLi5720qRJ7RQDl5W
RczlGpMlC92ZIChIX3RrH5AdDEkNsIXWPXsljhQGirp2BsmDefFBG7iMGV8No7iJBMtce8U7/bgh
kStGz4GnmLcByqNfrclArRLKpwROo44Erse0+HDUCIyU2R+CuEqfe4qsxoiziXyjgE4rHiL4fYWq
XZz9AyO2ppcUg6yWEJkgaY0TLYDQnAoG/hFKx/2GXz9eshAPBIHEr6Zn2azqzyrKd1k5eZpTBIQg
gp/33GCJ8p87SZTe+dcXiTkTfpRjkgQf+DHS1tTM85pV9sDyg7VWlwdgTKt0TTl4Z+1ajgvLQtNI
wm8OKUPgv6dum9GpJ6yqh/cGM7ayeQyivZdnnMpWCZ+vODGFXEoLXCTqVDItNaBQba2sX54yKj3Y
Jd3FgSQezTa+0hb+8kOzoNqkVMEx9wbVN4DPhduihUXBV2dLnGQkAJFqMzpXO0hWwKI9d0KEExJp
YZ3y3NKc4v2CSZ3trORYS5cYaoDxky83k6QeGzfQwq/626MDW/6Acs6x0mUqzYrXkIixSJyBOE+s
KDgZ7oc2C29QvV8i3aCbm9Ttamp0sRaeHLwCwQtX+fFWyKGJ3u0BNthyDtNGNBfTDvxXA/wLbEV5
W+fSfl2aObYhkSgsYyQfoEIu1KCL9wiLJbvoJtTJf8vqAmhorA9xHCtnykNxUf9xkG0jcCqk2eXP
fW+wojDOPFR/f1N33LvzQCg/KxHTXddh2tFyURUcE7Xea7KDp23yjv8fL3xp9k6O5Q9JcFjsDe6e
JHvT2Q8aSi5wf4wg8PI0wsWCQZlur1jU7izYu03GozUTXc6jSdrSyE0bvf0Y0MpwR7tUbBh5Izkg
xNsflDX6Fgyx7qDKzlBQBFH+cMKbMKJ0ndIrowxRLC+qQBwgmOITb6UUDs8sVHvD+YyrGm5o7euW
kl6grB23EeS77xu/O6dkkEQkVuMQpU7hQsfKfh0SO2JmDJxlgFjV7ZP6M4cwVyBEuEyILBROdLB6
DA7877gTWcAKnxPywp96i93H5dQF3LNoa/VfoIdJWdCGQAumh19BzNygvgCjtJwqsKTeWVaqCJNx
l/iSENZOoJbUaO4XvZhrsjTh/8ocogA2ksrkOS9+6WRpUAPenIaC2fvDpmA0X3RCaHBwAm7PhGc+
waDFAEXgwspZuS2DpkIokyjxms+4cyXETf1FStfeDpuablQtXjbqyBONx2k4tCLoOrE23vR8pWVH
APimVcb3yY+I2L6Y/aCbhas/Kp9OMyfB6fkPu2ASRodEB53KLcfJ6+Iv2fTZG1BBaZ2+kE1nzHtn
5wZ/rCn2Q2BSNDrfbw67fR/XbokJmEnqikiu8qpy5wUtztf/buVRWza5RbHTS5DHFKgs5Ulj1+y3
Pedkne8rYI1seM2rp+l8ayt/GqGCx4xeNstn4mWsL3VJiTzEuvWw6Y59M4BjkHeW3pTLX5UNP3Uq
cuUcmka46tDWc5/27WYpy6FHROY1XyA73ujP4m6TkSJ+LshAbJK7tcy+WSWbNh5fsJtYgo5VzmS3
4cOrPby5XphU0MAKn/FRt9SS/Xnoi1LrH2F06ACN0z1MIRTyLETNGclXziNHRC//wVhwV3F2AmeK
hjGbdK9u+6mJ8g3SQLSuoqukhTRC0llbhm9Z2eIQmJMlr7L8R4zSp3lU4IwgEUhngEPZQXNACBx1
1KBvjeE5I5WvRmP8QmVVw/ogoBcQ7PrceQitHc4VU0UQHvudj3ZUSgzi7JB2VlrWwLTNmouWf0HI
n4WL9DnOxfsmX86kSHVrtyISeCidvSkTC03oYs4GQbG/zm7s3uAW9ZEn3Q/tsmIw9e4HA6k4AHaL
HmNjy9YWM8W1ObPJV+/Ww5KiZZaZBFhr1Qc9QWJ4v36QQddWlNMewqQkHTWAbO1ENmDbKUyoTqRI
buN+V/ru5fcWxAEmUTsidGbCp8GU8sxkn08aqyCc8MAEG5rlI9dwVPw8cT9DkwWoMhtjDyjQbZCw
O4X0deO0Wy0vlmPlkU3orFj8ElzBg+kC5LqO7yVaPueWlRpriBsjFE8KVqQW3yDOjU78/AA9zZ4L
4Hrll6PKSji2C/6+KRPStE5tTHLUCkzUBbtr4G9oR5cWjsoIRlk0IVLBiRH4CHhrgBo7qiwPyE8L
//N6SWro7anqop+bUX8dfJo+8J0PUGedt4LhT/3FTWBoKYFucUXERFikZAe6PpFlo8ckHIOPBF2+
+zyVo/Jdy8hGTAdgrfLCwnwfeyhokREnxTWKr8GfAEXvi6DKk8cDuiStte+PJb1jkh3Vdz3JWXzz
dPnFVnUjtF4Zphw2uMLYP/asclXpciQ/mYpPUA9GGjledIM5J2Ka/PIKGZVdpI7NF8SJ4+YLkbW1
xI8h2IPzYI2oQxynwUFXxH6Z0t74ApXPrQsIgyGwiNhzvUTcxyLH8GOvecHKJfu90vlN7sG1JZad
oILoqNtuWzHk1M7ATDoKrnZDfl5peNTrTxIMdrjtmU6toxvVBhnxt89FQvtgaJuPA8lxnIXqdVSi
xnku315Fvoh9je9DN5ETX6G+zXcrOshIQNmxsfsz6ySZ+Bzmyry5SEo8IipKPdV4IOIyPANMc4PV
CCVx2lfj5/8OvqHM9YHJ3MbUNOK3BAOTN8v8WnlstCPTcwM1CSoCF/cbUlk8E6vaMKj6sB0aJ1e0
UM01lMBh3AQFsWyfo3rWT9dBOrWsPxBshFaqHxdRIdNzLkb/dmMo+A1nSswBcSQ9eM6iWObKZlx6
1qkGeAxKHR0phklGqLJeqtjFJV1d6tXOeRoPEkc41/0J+7iSf80jrP0Cal29jVcxrFKtjAuyrREf
hy3ZVtIpv8zGooJOaY4V2ajUW2VbWcEv+14W+nW2LqTMHvihxPaJAOb+ezJJklKU1s+dYxIYA9yG
QDTEt485CEoGKlspXUCnZ7twao1zGbIyeENoYlCSNvTHqGfTBUOP8RZ/zzZ2/SQ8V5y+LfEVUAYb
zWDTJuZjGxFhpCmWGU8aNGgdcszXqf5xIWRw4nBNqAKfzPo4jQd9eky97asriGRPsqvil+zgPDxq
++7gtYFl/PZhSQ3MqdBymgBBdSWxAVXogtlX91aENskxbcCm5ayOitAx1jVOYqryWQ2KHit5C4Cb
6xUALoOYIsQh/lWCavmKQ3Watp057N6mKbC1eKwwGeEoeK2SD80Cg1UcZ196sN5kw+wrDe3LTGXB
CrNjrgpdfTByaN0xFguxRJUw+13HT6Efb8ZFJdDh+QVHU8nYo70VZjvjyAdEhBfzg4X/Yhoez3Sy
btWAo4GGXQd1Y3K/gAW2EVNwjg7s5cmd5YBXxqNDoQQ/fiYr6G2KuxtyToRKXBV6z3ASYBby7e9b
Lvqri7H+7uLk62+ghNTByFNjwt3RRL03xrODo6Mn8HDGyScZc+dZ6R79KJA+jqfOMAAWs6MJtTLJ
Z9GdOJEfugiwThveshV/X3vHV5JH0RfT4IK2LM+/VTLeV7HpBhVgTmyDBEAbPTXlPWBObSRAv6+V
GEmhn/qm5SVK9go3PYhuHHdbhjME0dxUWiyNSN2kdiNEO/M8d416GzGFQlRKSkhpPNrc6LvWD7hA
GPMFnBQE9d0Bw5VPepL7rLz5njA01Uyi2rvnGCSb4VQJt1y09dPMPYoL+A3YfXXoVAYqZd/h+5iW
OUUnpltC6dRMuYt6xF70W1FN7GroSmwFTWGGp9ba169an+fvrDMkDMsjzzkftIZPOatO8hCoBzPQ
TYIU93DLyTcisQG+j4WbZ0b9kTlBIvq8XmGNY05vd7H6MHIecVFLyMpDm6HP+kbjU6pq+RBRH5AA
0eeWDtU3NyljckXbhUSK6UprQhy/u0E/pKXYWINYo4R/mao1r77zRMdarrmlFc2MspeQit4gDZ8S
mf/GDw7ID5S3VxQu3kut9lGH+jbaTSdej5l0JkhGotVc7p/kdJIA7TXBtO5rsTeZM2ltey+JTZ1m
pbXvHUMGH0MMte6IHo+xuN164GD8ZwKU4A6iOK9Q9RMz2FSo8VzeOf8qcCio3EUwph6Kc0P9AF3N
1ah05GwPX2AnvxgvgVvy9GjgGIgvVJ3h9m0q6PVSGG9f8Qz9MMYaB/9gBNWXEdUJtI1EuunmyjxK
RxL0V0g6ukDxArPGb4OF3P7MP5ba0TI8uGIzQc47W3doq582HCY6huEz67L7Pnf0BXVHKj6FOzkl
r269v4xidEF8HTSJcZIicdque2DOTeF5Cc7JuvNhSQgrEwkZ2OVKRxcbQaSADrux4z1LiYNyACaE
ZnFwcYn1MTA4Y/M8EDlnrYQiNGIopk4Jif3hyzjYCeQsoR94/0Psdn56HequiExAUItRk+hzSBvV
zoZCxrxWSSriwMQr0Hr7jRfcFrIW0bhdoDN+Tq+AJNNsnxZSa35/jA6gRjptTgZZVVgih6MpDBOb
MiVsORb7jtyfSeN45P80N+HmW6n3W7Qp7Nl8Us5tZRtDOSDd++AnpdBK77XcOdP3/IvwAcnJ9bcO
aMz9XaIA5VO/EP+MyDsVkLa9fIWLpv8TYHeZ6l1Mr/v+s93Kopx8EiCp8Ts76SepTSjMSlafCLQg
B1amxALjSVrr+XT8+X4rVFAPPhBJ1gPGAHTKDhM1OEJE3f1f9MyRwOElUxMZj/5kK8IGPp/ZyMXl
UuuVr5ck7Rqa8wkoYjhwNX49ponXvamE5QvU20gIQ8LJd5vyI0LWhNkxd259scMGr3zSi7myxTNU
1A4lmW0K/NDEPUtX+CLvYXMMO6Lk6WoK+1mnYMit79lBDDk8UOXJ1ETBUhZH4Z9XQfl42xi+Mi0A
zdKidvHqkWSKvDTQ64QV2djhDrN5qS2u0jLtVdRLmVkLfu6+n9T2dIuL/tQIT3eoicb9D4LK9QvN
4dgwnGwHPmRqViwmQYgeGic/xmzdkY9bhbNmBooZVqwyOaumk5IBvfQ/JezrRYw119cFtDMLNtv3
5h4F/YvnecRJhTsiEpO2if3+veCR/8vh1rR5tjQS1LIz2iHLR+ty44pSxkSk+IMgHFKAH6XV18HQ
/DLbhwKBfZXBuJz2JcTl8znlK5cLOuu7NWAIBzbXE4gFUruMGnk8sGRJne4F73sybP6jVqe4OcYC
TdzrZ4UbmzjOIj8Mz09UdQnd77sQ0APTNJbRoT3/gOnloKFjIucYhKdVUItLhgtFfae0RtZ12Sx4
LQUr8iZPrfqzRssECjUZNHuBFniDqQh6WFhnVyjdwUDrhph59eVHIb8k5c4RRNTJE5R5kqE9SHXj
GKr3jh1kKs2AOc6khPTuG2A299O1EYiByMBg30qBiD6JgD+IYIXpgp8lwE68t6fO5gtuZHr953Zj
Lwd3buF7r5Qg0Ra6L0Jx+gEASbUgqlF0n140cghwdUCql4Ev+oG0LMkWoLztImIgGLM8YhhFP6ZE
p5bDqMmqD15yKf27sVgNlzelFu3FYJLfxjt+6T0fdrZI4KvvEMdLP9rtVSjnyFbfAZwRpSzjevkt
Ste+Kh9nEIRLD/fdeXk0rzo3rgake2G4A0eTszzP0ApTM7u4iTD+SLxjUYF5SrXvUbED1762JEXt
tlQ7FJ5ByB2ASbLarRPQgpJxkEhqN8sSUIT2e2nnY6MKN4RsGgBoaHkCB6bPqLEnwSj7N5ai4Qi1
3JVImua+vG2cgkS4CrlZ+wysQzJ21alabHBbe4gOxfYoWWX6X7T3lJDhj/yz2PQMDMWbbRrKtz0o
Bwhv1kcczi+Fd4z67IpwZxA8nb1XVQXaHQ0MTLZSXyyaU6kfUqbcZZ7X3erbkoAUgvc6rGRjBVeK
6YbMmFGHdq4zICuXdmVMOhnS7o+m60He9AF/u5BekqRp4/cFQ8cdSpK8vcmIEWWcge84EVwPQ6ag
L1F5WFh1dd/gFsc/oPL9J8Un1u/cv+sT5c11amB7AQjVu3M1oL2azcacbwbGqRy+JbTGyYVhQdiK
pmpofJ21T6DMisNc2t5SE/2kF6AxFWTu8AoyVY1w1ql8hVMOQnJHn4QjccBAPFNKBz6PPgWnXWMB
vdVIvLxCg2o+VXCjIG535SKbQ1A9s3bC8XLYIIlMt6vl6LThQ/70GDNKzdw9wTMowotMWnkxUmdP
KDOx2kpEJFMKJzo7gVwcq7ACHqqKzv+cz6hB3xL2I+yWy/L2VXKDzo9KzFDWt1woVHxcqUgwswpq
928NBxBfzWBDEiGCKpIKNWbSr8MTJuSgKZDkZeEwDQZgz/Sd6UyzO7isbbF8gDi5ITr/BtUrmhwP
9mhDXwpsdBVIlZV6MmiR9Eb5O3NSLcvApYL7/QUt5DgDnHC7SbFPLRhOw/mFDjYppAraZIjB5qlq
RVrX/TRMsJfRERLDKffy/KlMGb4vU3EBLiCyRocDRK4mdZ4iVQvmfNKNdRNnfd3/sA3ik7wtkYPy
iDGbaBbXuezjjgK5FasLNAO0AcYdjeZrWRysCzvEpZ5tmlaY4D3xutoHXnNeIWKhUwE+v4B3IoZZ
Ch2evLWc1yBi9KCWJbA8MY6UIX9+1Kh760pF+ykX0iJLU/GcEs5U2nuJ0V0TBLRo7dcaskF/afZY
x4/6ykZWhbBybGQZfZbKtFgS/qigmrgFjTTewAK5PViHzcnZfn1JMBKoQ1LGRjJ/4zTJ3QtiEgLH
HH9+KNno4M2lNb0kJ5EUPZaiM9qLLLmUOLFPusjpQd2+MCMCxqzZ6w6V69SBEcMaNUyoEHjY4BcL
h/PEq6whqryIpJV8YSFa42ZByskHbsYQcCvzf2ypf7nxO1wvlBoI/qmkpq1FoSVuKGh/xHkSlRqs
iC51Woz7LXuoHbcaMrgYEMSpJJ4m3MKefgrrrWuAuRw9FbEmvb0KB0SeNJUjUZonQAzvsaLWJ+72
15yIHfuJMP6+x+75n/nBlPM6Dg38iWYhE6xK/6QZk9dUlwl0tM1oTjsRkYoQluVLS9GLvopQSqOo
MOhNiqZSNXQgot2MVUlIQtRC701mVUw8u0NKJvdAC8PYcab06xnNNumWAj+fXZKsGm5ecwbCPeCY
iuNFcsPCQpnGWwEH8zJ+XsVTWNavutUTn45Cwlgo45yKgBySrxJaYiybO/snk9+q68yHt8udO0Bd
jctyfz+9+TMXmczhgCYHh6hNPXNPnOJUOWmn4hivuuA3BVEMyRaXMEmdLSw7EhPYsMIKaeka2GRN
bSPr46ukYD+6cA0SAhc80nasO1o6g5x+ht0+KccEmAuMhJvzEfT9yRJoP1mZIgPlcu7WCAWLPzc8
0FVb6NKzu8PIOwTFUC2lKJeTpXWlXwGQdYePynAEIr0RNP75cNw9YRT8FgvzP+QDJ+0HZuScDznh
nVD0CJ5Hi0LQ98aWf/2whVnAYwtMnaouqeiMLR1zuL4uWOJnN5QE3dmh+LXwWnW8mLwPkktK3jmx
K3FkHXodNjZ3kHjBr/ZbEd3/sZMuIq7Tn5AqF/ZQCXs9GQsr6mIZpSAkZNdwDscwq7bW+m+GrQ9O
ObCaOUDKGJFnf3utHuzOeiyjQQNc3yzJMLW/KXcNTd8D6gPILHJQH4XvkzycgW4hiUme0DkqfBFP
iiBwjOrHSnLCvrJ0a0ayQKkuqiGLGWTqdkt5UZxaPdSdmO9lmWaZ0qCY0RHyJJ9+TaASV8lt6EiM
/5H8zvYtsXv75Vmu2wW3Bi7v9VckcBOnwHWnL4OXlGJg7pDi4eI0h6x13h5gU2u6jyHIDYQzqY75
hLvM28x3MEmbqlEs140/owLkCu7uPsZBr5432YL2kor4gj1o7qdXdj27lek71ci1jPSkYALtTxvb
gLqyE2qqkIUBBQXCUYPwKd97QiyDEgcoRrB3761Dwhom2x7eoGYsedfol0nGlByUw2+F3fCfAY+L
o+Ek7J3EL3SyJJEhzZxO0LsTuDOzdXB7FZzKev1BgKINOKlcLQuJ1AhtESQkC4vf8vysMibyXnIG
qm3bHwXjWU4HBIb8hr7IHBQikAjhIf2TlORQebK/PVxHVCsSPozYnVrmhnXH8Bam92VZ9knfneQ7
gOWwzPB9yPCFzJeilEKgsv3KcN09ITyL4MLUzw8NmFLI2dpYHnNgQ3CwwMQIMeOxo0WenXr03HSy
zBXBL8NyvaJ+UCU6NsfCLql8p5EWvipkzahdJ1ov2xREMgrNpfePZ7f/a0OF7QpFHEcI8uwSpxL0
SaPbWOmFyzDNMvdEuj3/FFa1Kudx5GQylimOau7MSOubotherSVdXBxVrpAReAVOsQ7/vA691OWQ
rhuU9WiVIUUpS49FpyLZVb8Wv1jyr8k+udb0b1zdsaILatH3lI5f36mKQtn8k7lZIU5qLwmw5aBs
nwsiPtvEQzHu2Wz8zgvI8R6T2TTyI0SmPQgTMBk0tseJchLCaCOmDOPulZm7auWH3XmUIntShwop
YAKgSnGse/KlQjHYgBIrkKkEulsjL43pdTeabqSbZR0KIzySProDUnjkJmzGCA9iDM6Ff4HpbayO
wOeeyO+kCFb2el+oiatcmhi76QEBxgj4ih0fYumLuMFqO9YUyJJcUKlFCnrhI5de8g444oWM7uE4
GOrMI0t6d9IyQdGHock9mCIlZtRhijwfR5vFRQIiIo5VmXCELycU/+OM0IXuQ3j8eoKxzxiMzaX2
GkuSoSfppjYq7t5iQE+BjdRgSWUzTa4yvmhtA4Fjmed/clvdxhPjjJ+h0Oq/DmiAr2MujbFp6QyD
G6YH7keRpsgJWat/vD57nZo1y8R7N4StYVAQsaSrodIgwlBnQObzxnK9SnLCjmXX4bzOjR14mNdY
qxKc8j1PBqyhiuSz/7DuDre2wY+wm/2x0qnxnRd1RQTXbsJcHM7hg9gaHnM5knfL05QWn7V172wm
mO2Mab2VE2PJGuNOQ9UMBRToeUlGD6K/oEy6X80CbKu6q4XtU7Dn981q1GFIuMFem432abTx1K4c
al6MK7JY4j7qW2I+yNX36F6YWpWCddKJOpNmXvshrXxAtYMpDfYQRm8h33rLu2RBIHCbRatnGUeO
iCuWbvOzvDR6hbG/LuIjbb+AIfowhrBykpNPXdAXWVcIFNv2sI9i5jJNnFma53cHexQKd9v0sTMI
tn2xyCvjWfFFrCougwSHvpkoJRy0UOvFZdbflnp5ERiLqJNjF5zGMX5+U46LYiSJvNM3QlyLKMbF
0bfww2p9F2Pl4RS949k29HGMQXZ3yK8U0qGwbC2Voclf5m1dkdp6YwBGXg9GbKYCIh99ZbpZ01Ux
A3V6DtOVCRRGEnN4qeRS9iKTPqA0aJ8iF1pdFUlspOKHcJPZcVrLKLqPc3cjdQKCC9PZzsP0f5rD
Kf148EQJOynWnGaxFku4XoT/OrM2M+H7xoDunXyRN6hzfZHdV7oY6QQxis1DfZ7DWMCMpD3sL46R
Y/zS7+I524WJawoyEMhJVWuBtHPXoBVEdzlkx0ls5n07RbnDB8anb0skxJsI23xeKdhHl2yMmMa7
86bpb2H7MM/gsv6aeS+Dk6d/KVYQLvJLRRa6o1WqKI4pCKDrzm9MmZsod3gSJrKICGu0waQXx66k
P6DV4RsYM5Jekbin/QGGQQXuWs1UOsxzCbhUVSH3AJpmr79UTfukKdJXxECFHrOZGwC57KrVrwlH
1RjHUF5W4biQeWNHaryvPMUPEDr2e2hdyng5EF3KgValQXMAX6CzegT+vGzpsvXJTG8ZSXXh1PVB
UMsMRZD3ZqLSYzyUApF9CT78PGRk/dnFmb23evPNSAOmIZD2QRq0fqBAfuhzlFSDB0gD1lh9zGm8
s/H3DVOO1IfYC8m21jcKOcgYe4RuJ/JK5kISjzQVlFVJuEDPy3QKN1+3kykgFEs2DhN3nS5hJu7X
GyXKrQM8FlSGtKOP9DE6I3L0krQGCxeKT2aWlCvV/euBAJxd/w4/1buLNjIw0UJywTZW1wUNJbOJ
BWLPgk+cfarQ7PcuTEFKeNoYj+R4E8sn/7vys6aR4bE1opCMurNBFuDvjFbnhV8XvUQM+6hB6yKa
q5HuAHlaYbrkRzWErje/FvfbVqO4E6Pj+wnFLfDUOg4HrLmi895cq1WMWpYHJj2NWMBr/aCnRHG8
Bnckl1g/BnCvx50/9pjgyec7JOwpoXCCpeGYp/Lup1UMGBq/7qcw/J5zocpCGWrwlUxk9cxIhCPS
LZSOQK1rpIWGN5FXWSI0cm7EDCL9heTDwFXx0DgFpGGJkFRwesqckwDBUuME3kTmEWFqNch+l2Bb
u2QoeYJS8aiapPMA54xh99wdms9RX1hgEa0Hk3sz4NEBXxMz2iC5Zfbaon/LNG8ALY4xHs+PDw8r
heJqmZJpm/j6vZiQRuE69QJ7Twahg0RrVkg8b1DmFFE/zziTTCQFAlmA1vhyNk3mQbnAovd9TG5b
Qurgs4xkodVo//KCU25PWSlVe5FmvD0WQrIOKV5AHH/sol4hJST8I5Lhyps1ohyhFc96MNj+p72E
0Vg4Q1nArnbmU9l0vf8rwj+8Eud9CaTBDgnk6VR3yo72aexCYg1VS1MsKrlN08wUe6sfXjXZrUdj
vwr0Jb5t9RmSU6FSfY6uz62mSEKrKS76c8eW940gTB9jH5fHdZpeZhnLjIcMM+iGRUMPAMktuY7E
Tx3qUvD+RTWSv3oELikeGZhOiiSlV4WmYXT4z5Fzr+LqwRQHS44mBcUWaNUm+QZmWmtaupmplnD0
uAZx/bzgo+CwBvm3tcr/3TRjqVEwi8ciZLbNaQqURjC0S+wiTfUTAfEBmdHVIPxlXVekq5UUEaAZ
423MVWLiu0C19kopdeeCq82PsZ8r6wzuNyQDLO+8uNOtupwKIaAwnX/fTNaS/gesPGsNoPyNqVLq
LDEElK2o4k2dZewdEngKmB8wEUW0HXOMktIfWiTjSy6M8Txp+/g5I9KmGLNh7usYaC7FxV9dOAKP
VIM5PttcWKoCa6oj/LxFPR+xZZmqwuk8TqekBdblsevTsE0KdOGC8I9nAc5RAx4nvfd4m5bovNKL
Wj2E31ldFhQVZOEdi87my2rr7lYflQ1SakNw4zE6H/NuegstEIPXcLeYXcfalUWLND+lotJi5A64
8sH/N3PlzLQoPPqpBzzz8MbW59K8x6Hilp2XTYVGx+RVHorv3L3T2rwwPJkw0dB4WnP7p7FfrvGL
B0nBuiM5S07VcyhGojmSbBd4U0fY8stbnUTx+txVzZlT4OZn5jzgSeOCKFAbVfGpm0YEFtqCJrGB
lDN9O4MCjyrOApnn/yCONYb56sICPtBKunfpDSMyU3z5KbEmUzVaZokQLqFopUfk8MbDBj2jt6lF
2Sh0CXYiB4RsVuILjJWORJwi326pFDCfn79KhbRXS5uHw9KaVyrjMQJ5c9szlE9F8LoGBwd0OhMQ
4F3Ydu/IkaoWasQr/rLrigbgkmhsi4w3lA8yjRF7UKmtqnpajNW5V0hZ+Wk6E+GrsHmjFQHbyZeE
m4v8hhvYGQBMM3q0kt8DBxbrUNl85ZCsk/esNaHwHQ7IROJipYrNIEDEFqfcLRXhoPr1uvi5jJul
7dTUNEM4rIeWkXZBa0PKhHXcTzpedRX3iaBTZir80j45fBuWPwSrVgHtZiMRD1zhJ+TyodfvR39v
wdr9eaZCfRoRU+KtDBqR+J9qsoFlYTTA3NfxrTLXtZX7lfIHTqyEGiWjjWIsetaXIAtFlVTxmZZV
M4je1GyuRAIgQhUaLRauW1Fq3ZotNcX4vRDP6sz+JHlGXuJxhCvq4eG0+0isUugZ9wlJE+KzsvyT
Set5jggQzzBKPC67hLCF0MTU6sA+HWFXKGgtcV97/ztM3witSWCxyDeA9b8nqIZ5BTwuVRcIG3A+
d6FjTDlch9xjZyOkWACLgO0H7LoTie2b16Zsie+L5QjSULtJ1hfTQneMQX0Kj5zHsGhHu6P69VXP
YX0gdehEUJOCrG15rjk3eKlm9nbL6sYT9CqVm6m52FXN9mtM+DcxT9pZGF8QaptOYk79MFniOZDh
iLqk0r1iWR4PVi5hI/svN2yLdHR/7AJ8rT17S4+xwAcInfq0FI3bNXz5MASDjhJ2g1b+JDPpT8hj
TTmnDa5aSAM3sqqXZx2A9Ayu+8TWuaqjpjl4DpUnsLTXPXeV0W1gf52Tfmk16W/emNSCMrmfdms4
MjhbzB25OocJCe+H+mxtk9XIFNJI08cdoMgPozUi32gU+SqWu94EJJPmLcTtnjcot11ZDTdLRVvR
GMyq+MnjJiuSVFqkoexrS0SCSfm6oK3G2JkO49+OsiEzl6oFQi3uEI5Dku0DVtdi4pZVQSUU+pHv
O5rG27HreWBnBiRLmF3kl499iwVHjVjlmhqZbCpeDHdZ7vP774qmzFKjP/w5cvg0kbDmuM5aEejk
lAF6in4b1PGR+UZym5pNVQSzY4PmZlVpDLpND2ghWHVJ8+ErOKwVl6iEuUKQPyReX2xgjeaI/ki/
G8mKi2B7oqMesGzuJ+sPFrhP5zOjqHANdfYW+Pzzs1afRd2oVkOiSl3wDc4OeOcMNL7+HLx8wfC3
9K0biVvOtf/WOuf1xF9z1hvmZLA/g+wZAjbI2L25CIHZ0ZL+E6hfkkBJOJ7GCW/ES8+Zv1Ihq+t2
BT6hGYLEnsQ9IqNJbj4qlEQH1RoG9QQ0p61a1oGl7p3o2hbSTsIjaMk7KAF5hSJd7CrYzlOUTJ0a
K/55fux3h4mXQstx3LWFNRvvGjOLQmAjoHHb7C5zzaE8sNeKwHUrHbYdd7+D9YewEBwMIH8CfrK7
7V1xMzXy8/xHEiYw0hmhW3htdp+Vn+PqX3BiBxd/Ic+TimIu6tOA5BPD4xUHnvkGm0zZoeobcIZx
zUssA569cgYnFVUUMIE5azu2gHffGzurrF2ywSBr+fh5hH+w095XM1djZGtQPJAKWGyMmqlLaPML
9rVyzgqsCrxCAsSAckKEJ04JFMBsCsYBknlMbhUhUKdaTLfMsXEJ8dYNVdTCyByp1LKiFeRAVIme
S+tt2eI4gxi7Aicop1AEkYkHhBw4g4A48+GoRRpI8KtRfE0XmLL3byIpAcQd3xzg9EtlB43kKlfL
i9OIYw4eJqHpgUP/ylJuuiMMt1L+sKso6V54FrIYhmd4XW+HK5Im410YU4fDwAsab55+d2tZfChZ
IWl0RIfsQm779sdZfe61w3YOgoEtOhHYorh+OshBffrg87R41ftegfelnOFKy2c3epXPPYjkk7Ql
r9w+n9xqsuKEVcoG+Q4urBjOgI92NNr5wdwwszgfOUTCIgS+H/zyOSLh90tEvUctJCAjN6suvRVV
lMsuxtu4IjVSO8q6tv6Mvpmwx1crDOLrCvnGtWXjOCdO4WBzZoTjWnpVBC+O7fYGlGU0dfAfG2na
Vsk6IvAIfzAQ5uywpOWfbJxXiRpxJeW1FjmBfMykLYrcvXhLD23bfrMcNqTDjAF3dp3/WHAYTOz6
IrVKwCOoGptqdeFDOkDTG7nge9mjuGcycqbREhERqf/wgzeSExlt7gCDXj4x4QSQ/6ngvIYyStBs
FKj9lRuKcZbT49jhkQ8/XI5d2n0l3WbSS+d638SJt6i6n/MSkAXrpmUaqmaTMK/nnt3Ct0AevRee
3WYPt9fhB31LA6h+UD+i9gl58faz9rhXQs/kcOJpF1wrygCdfEodgCAUXkf8fcUagacEFxAseQfC
CNgw/vqVKRbBw6krivg5Ok+5nGUdTRbvDFDez4s6HB+REq9lcSKezE4SwsuOjUppoT7hw1XgmX8l
BCDapSJo/R+Lyu5PcEN3CI6wNks3+zFiAnBpZd4//f72Tley9rjI37t2dDcmuKLRxWNRpVGbmsM7
3+5pMIUtVcMG/8TZ0RvcDyJRE35gijGhK+clWUO5BM1wNFyueTsYHv3I8Nc7foRw1nuzXajX6ezs
wI3JdT8qAVcFnD4Kw1v/lEj0hmzYvyGoTqTv9ctlUAEIwRU4pl1oxTogTfDJXig/diYN/Nb8ibxl
fZ2M7SC/DmmKYRMFwgXsfE0ktYNKJ9km0TAYzjjq9RyDeFPD15LEBY3PJEdjcMQ8g5eOh3K8xXMA
EcrHHFKZugbaZ3xnCf0u8KS2PBF15bx2CwxovdMkpQtP9BGOwZKH4exUhL3Z6odhHCmh+ynZ5HY8
/8AKnCwHlbu3JyZCzI5L+CTOM0dYihI64SzEsiW4bLmDdRGqUdFC3ZGh5MdQO+xKzytAajHYl8wK
X8/ipsUDRnsyOn12YQi2AorwNScrca6B/m0pWmwmjPGVR6VaSVqdOxd0L8JNsZxPKRAFaEk38pcl
C/2Vr8FD+FgRW9m2F1LAqoQRRSWmjbBg0nyZXyDY3z9y2wWS3hUQp7dKfFtkPiNyEgesOVZAc9hY
RQI+2+BCFRvs8NMKcCYFldEQR1o2JNi3UclMMRlhUZdRgAuZ3SAd481lfJENExEoqrEopMFspz5f
xzzVw+WAdysfj4ujgMaYf19PL6QccafxhUbYHURvaMhTJltsa/0Pg9eHOwCt6lPBSo5zGH9G6wrH
XDhgAHXEoUpauL87yI8y3HdqRI8U2HitUlK0LAkRHqYrJdmqWi7UrFz4XOX+HweLncWLEzhoAr6C
gbhxgwL16w8IbXXczzaufxDU4ApoX2OHDbyz8jLn9OPZjtbDA3Ad5CLHnVN5bSQ2yS2CBr6oX/WP
drOecfEMXhfjWB31fg2xcZLg8Oe2yPp3M0AxWPLR4BOmsl1KAeB89vUW9bxzR9vnI2rNAmsxuKEu
xqImXyfhljbxA1Uut8KuPvcPbzH31RNHOrT0AzvRu5SzBphH4eMvfWxNz6g16Ofv6v6GRgbVe6kc
d1DEdzYGjAhVyzBwqwEx+t1yo4YcsNoK97/H3kZIaESd66EuxqRaiGQcBPxujDa1nGaiSgn2quML
uFyBwgf8cKn8ZTK8jbzs0cGFuhw9Ol57qFyP/l4Ru9tRZCMzSqYvUZEjJB82vT/SnYldgL//fiCH
f7+E0dlAVaArCbPbpDJpi7E+Dw6DNsN6pWzLa1qi0mQWFSly/lK8+H2uU2aecgrEE3vqU4KrdURg
nJngsgqBfMcFKdgyojiBSJ6BvZoXBfauOAwXQxnZ6UK9F56ktSirq7432UJhhzZchcq6d2jUH/sG
fn+3sLqsNShQ2de5J2lYCsdUCQpWjMwXjNri/WWgxZp6J/13xA0Qw0sYC633dlDYE4FeD4QtHQ3n
dMt0IIjeJghSXCaj/ntvFe/LjB6Ugk1Diyl+G/OsKFkgn/3eCjNuj9wdDhme4oVabIowmYUy8lzg
WWATHY544HigHdiHRRL8Ynx5xW1FvIMj8dsmqFXt8ib9mEvObHpa1zIyATUnZh+4TY8dM0TsRLp7
NeAvXFMH1xPdcyl5j/8BF++gTMB0cjc2ichR2EG6NvOi0tA5fToJx1gHpmcTXzzmyVoinOxOw1Jf
OS+8/XGebyDt55kpJdEPDw3ppzViU4vdBMiA//UqcgXJacVQZm1rkFmYDCHW2uETclaRJLlrzgJv
bAj1Se0j0JMNc1YmIy5JUwq2rcY/SyDRKHjRVoONTKD5ZdUhZmmzheROP/LKCgMgFXAz/6S1acId
v1vN3AGh/DMqaImMsy70yQsxcw0OdDrC7mOT26SP7utL1b46e8uVEhlaR9pJNos2AVHuEI7AFpR6
p8pZ19DgbydhlyBvNBSqLyaxhopa8UjJl7YpzkF0AaPjd9W2Yu6mvRmsmT9nG3WBUjmuNPjU4aA6
PZeG/4GWsvsemEVMVweMIOPmNPi9cIMyhV2RJZQeH0a6bAg+LMU9aDL+OmEB3JbVAPpyO4M5ZH83
zbMSMKPBqXnhLf2dOq0Mvzmpj3OMlpR6uaqV3zlhWY3yenAvpNny/M7Q1nG7tn4JHVab5e+UWCib
M9I9MUjXudNzTekeLWWTAryJ7YVwlmiFcIMqQLziB36Sl60aH8Dc/g8cnvpf4pKpf/ElldjBEFCW
yjO1R3cb5gLS/SSXXwXXBdDbW/AV0XZ1kbNZKNEibVxrjTymY1LItjUKJFDIFVh3gu4Gm2oTwqy7
IZAnZt5TjTW96uFMv0MJxmmtTAPt2SEXiAQN97PjnvRKGSVgqIWe1PNQLWQ5yhGrJdLdh2xlcT1P
sDtMiLqRXofRYAKDW8FsdK3lJgSO22BttmpGI46Ft4vEGHWFQuridFumfc4hfA+AqY7e7Ux6ss92
lbgAFN78gQtKaBkmFABfGrXwFFHLigTVCKNqrVFaeIewQHtI5166RULtI89SVgxMwopFX1g8HM0s
CmxCkabaTsc+WzA1zLLCmPkE9gfgvmXCKFFnOJ6EINr+QPvR6or54RpPKzQ89yZZ+3y5CkCZXQSe
SrKxQJxeyPgxdRnSI4Pixx7ebX4mVrSRBHpANJ7G+KaavtvWrTg4oqiJkLNTsySwa75bdwb8No38
5GCxZABNTEdrE7zl4lGy/356uTIDUUtBe8QUnFfxmFeo3W8OHI2PMlmUI2e4t/ByRiGaispDvszu
lW7L4j66gAWX/Cn8W9TZW+A4Rh6CHfTFBSuLBQe4zsgnIAnRUoDdMgDZm28uvTzJHqVe+R1v/j2n
AcWvLZV80hYxRorh0f99XJDlbgD8pOj7OwesG+wlp+ZwiThN2ojo5lo4ZFGK0vrODuw+kaTLECJF
JiTOQzob4OGHNdnW0FQb3oOAYa3TpMaeinDKNJayzmCxDSaUQjXn9HHnttBpX699h4x5JM4NRfIN
K9q6B3s5iSMPhopnf3o/KpDTnwlFXpJRmZMBd/JPSSqowLSYR8/te7NIEXbIuzWB0DuP1ifpc6wj
kHuI0T5dYC+0b17Wv3UL1dxnzAs3JhQqw3Mm7WnueniqhqxTKP07+JUdWlMLdCbI3efI/vhiWoRh
6tbbrknIQK0G0SPiu6Q5KuverCIwBHEHS4hIvEDpUWk5kuqCkppf8RpRHgVge9BcdLmsVipQFm9Q
m4DQgYZtTe9h5+LS7xwrkqnY8ItzxHQHS8aHFaPsMdMvpUcwXftWqUvVOGgVeIAm93YSo2zRjKwT
gvYgyHIUH5KIDxpVaOLcWQ897cf9mpighAO/Jp3TnvsO9O5NFQH0hSqD5+jGfE9P0n63CyMIRuRs
WW4hIvv6LYex7TT/yaBEplTa4ZbN/4HHvfH+uR3nCh2a8DAiN9w8u8fqL+suPZ/p5Ob/4MuD9DIV
I2F67Dk6M/qH/inXrm1xp/+6rqtlEm4vI1uLdz7I+AqhyjfSm/szSpx6fQwgZE86L9EuQh/FxutA
ywonAvYTAejWIcYl6YYE4qpyJeAdvorlmaU5dPCyo1mRQeGRFCGj1vzscfrM7bdIwPL8/JU6v8mN
fy/YxfWrSkLdV/tDR5nO2DdvoLmr2dvH5TLIUcotT8UuzTHYH+xXqMAXc5Yf79L2EhnD8mCEw0Gk
jVmUY46mNN4Ti0KcoVt1HuipAYIbeE+KnHUB6ijQMUQkI0hyRPFvzdR23UwM8CASOdbC4e7G7Hz7
c4sL9JpIMAVWU9mcnDyTC1Y2eESK70PUjM8DVQDrunmbQtmxbVdmIxVR9ciTpCT0+XGq9qWuWTzY
ygoismfFCo5F+oJUdGC7bfU4VMV9HUgH0rqWiRO7eYSbCiMCd5ykW0m1DT3Uc+f4u8OLZ3jVC64P
5/ccTquCIsLVqGyOVe1O112ROEDqqWceKTL2EDSSJqQQMjjoZ/VprbL0GIF/GmwYUXOlNAXAknMU
PmFhaf0uDUNL/KCyMbwg/h2ni/qqFfjLwa8pVfae6qnIb5JGzRrpEfWyo8WN4uI1zUwDJXktp2Cp
7pxfu9jYbCCKA/JrsqHUjiyD72rLWbbvppJsvtIP1RXWqpwajNNxTZjLsEYgJjd3TkK8By3RDwF+
eiA6/e2VJg80wGx1F1truPZDN1pq3kEzQwogkHf5vxyMkxFqK6cjAiqwAKZ0jIx7rjAGQITBIjPZ
z/dZTX4WyedSbd5xQOPHNkuYx4dX5q99O/VDNujYe28YP6O5bkQqAkNxmNmLcfkXzlIYrIDsbADV
gZFuuuKOZQhPQw4pfNdUldZndGZz66gUO769YBW0tSI4nAG50TAaikdkAzxvOdCaTElD6naMXMZ4
FJR8zueeHYcqEHVb2zqV6G068YZjF89g+C46MT3ZGkem8PSNQixNCaKZkjGU5Cs6ikqtXDsr7jaa
Ret5h0uHwNJgOZ6hEiXspd2XpPmdxoU2o/+0N1SkyPzFNgvs47GdpbTmRwQ/o7bs0hDwwqdzW2CV
Q/P7YibQoMH7O15EWdmQxtnr50E0VOXh0pZE/hz0s/E/kVxfXrCH4pSEkY7deUMuBPA3CGFcMjvC
m2vux1qMeipZ2OOC+zbyGQn+eYfce2gLkY+8TkALWJtLN6W4TYI6Bc95rJG7apaHieb40M8PyGJE
GOnPjIucInX9lRH+Cm371dKD3fMcx+jmoLtAQmQhmO/ybXF6AXQs+GZxun8yxb3Z0aUKayxpXu3n
d/n7Ory2JHolSYSMq2oh1f1Rrlr4R+vc1SPIJIRNRPDqKb9PFqlWwQyZEHiacofF0z1j9HpnE2g4
5yZY0cOs801d3sR5qmcbPRkkpgMHeRPXmaFo78/cqgElwugx/HqZtYhzq4X2Z1DXczdXefI+JPLh
6sYMkkZPQLcKjtYPxMi9yW5VpWyY6a5XvGtEsDVS00DJ3YrjXrMIUWDxd2aM6ilfeu4FV8Qxb89g
7PEN/D8CorVWM2vgbDGSj4qG5WsV1pRfMWoJU65f+SdE0W3Gb6NNO82ZOExI5d7/GX0Rj/oqoAil
PH1Vphswobx2vQhxbrVuvO2rNTdapB+QpJ0buzaJ+7HOxELIQTjuBbK8tECmn/9ZosrRBRw8Rogj
cbD6KVgiYJh4TViONCBGlEQOUYzQ+8T9ytK4WKUtqTh4ItHltpCfpeMH00ojY7o9Wnf67TTyn+n0
rjv8YwqYxzqz6XHqZzj96aufDySjx4/5hGTOxZCAkIaROVIkSByxXLhY0yjJzaG5vhV5tPWJriid
TW6D19qO/+c/MhO120QH4r7r3n1gIkuX3yqzRnQ9M4ZyWdM5e+omUBZ7Y1VDbKrv4Yqiy48LWRgn
VN/IKyDz+cWZ9GDSg4E06ahkk+6acVTb1tBQUS3HRuS8hY1v/l3Q9WwzrDlrolkf4kpcws0UM084
T7Fw4nXhAhygLkHWavwcYrQy2sDpIvUrinHueQeGA70SLg6axwJnR9KmdJ2jZw9qEdGdbbv1y557
VtsxwkAczemKNHZR931Tac7gMIzE9/FTuFks6jOLXVwY1S+N4t4vZvx22hJ4vTgHSe+K6gexNcKI
tHMY11D8YB8xodRR3bIS3f6XW6PeLqBDCXo6Uz4vzBLeDkRp5klclEo0NhI7WFfqWyLvC90F070A
Ektxyslf2jxWWQUF+hZguNEDw3Yae7OZGq9LyCiV6s5FtpmXepw30l386Dwjk02Cpqfa2g+/PkcW
hhjL4fctvJjkZ0Twhw2cdpjxtnxbPR5X6mGYPdz3YASo69oSsewHSTjjdj6hXuqRCvShiFMDpqI3
5gxjV+soymxBQtiUmbqJ4GUpsazm9UdVtYk/IHFkwF06gkHD2huIcYy+53QaPJa1J6SxAFEoUCeq
ZLWRUBoPMLD6bwriPweORbutbvSstEg0eMBJzH45Qg1i2g5iiXqUad3RY7cR5t9R6RsaaSJJpPVX
v5c/8NKeJ2ucE4IqKyilRWSq6hY/79uZFPJB4dGFph++iCeyWkLE8qbeD6f4p+sjDXYtRl8IOR/X
N6gW8hYGfyof4zokxTgOibSxe+lI9v033Oua7JB7WMW3hc6awttoHYXVPahY6CWNPJt80K8+SbHm
sE2N8+NhQ0N+M7bk7kxAMKemLzW5V3G5cIAhajKp1Z20PotcUOeqp45Y7e00XwuelA58p6TkQmGO
JfmEFh6JgSNjBQM+I8lN98amDTjdHTYitOjVlEHAICl4AZ6lauFK0Kjyh3erhf8yuhNAqxUO2714
2AtrXdqUxC/iPSr0IxffTu2J3unsMjnbcnf0Q+JOjk1HtwYEpWIzUxB2KLuaFIm0wPhVQmh6tVrJ
mENKe/iXzPtDNsFDqFll2ylWFzGSrQEv6Rkn5ddgCIb+0UhKLHBUG4jFe51K554xMT02oDTYjcCJ
+5obLRCgiDS+gOxHLXpvoFLQala2QF17UCUpy349IOdNBfxYuvevqIkxLF/fRLqW2pFisjcIAEjx
N9FiMetgrEUJ/nuU20NlARnYhtuYliYUbQKz7NdfRLDqHjESbH5QzNviGFZyp+o40JDEC/RRL73U
SauDSrVkkdddVQp/ZPmPHv4RxDlC4S3hqFsgCoWlRenYRrY67ESVgP8T2IZRe9hnx8/SMtLttRN8
YyP6bEhLW3uZx1VBLuixn3+jnP7zb6o/C5+dnZcfQJ+4R7CVtVzsr60rvvKZK5lcmRzz6csmObLm
W/Wn68yHMo4HyX4/OwWuXBK9TJN1GNhDdBbHjaOytWPY7Nm4T9Pkg3oOO3XtOL55lAiGyioo3Wx3
gL4hUFq+o6Cb9cK8Sj615XLFQKzyUSslMaVH4L5dHgB6/PgkWptADN7ROFSBq4huD4nvsnHjMUnf
qMiHXcBNg9Mqn3KfwXQ453a8ChvSeIRDcKOCXQbHMrVOe9+b5FlzNhzGBEv4HTfxwvI48ZIrkF3/
2QtEJlXlZRj4F6n4BcxqDkYCzhxFYI1Uc8rUlj4QZUyl2QFas8T2gBW5Qjz/fg6cJBr9ng0FBwsa
bvHCqlaNBDMttSLa6c3qUibeSxaKXd3ICn41F4KS4RvupwJzVNk/y7IbDIM+7d97w1svaME1ew4l
nHu3tPBUCIiEcfp6FDMqWPmEvcXAqiUCBwLxhc9v3iZJDZoIHnT/pX1j8v1Y8Gs7YE3dPRFeVt9W
TGAJ0CST2iJHsb8aJ3i9S6CQnvld6Y0Wz6v9Z2psiY1HPIJmb5oLxWKL6U1M97ezeeP88RQBe00d
LIeFq+7pZSzkxp5gF6lhf9KXnyMJCHfxe6h3ygTnEZ5w6c+/wDPS5EzH2sXo06tP+SF9qEEW4LSa
HNkB/6H/iDh7KJ1qfV4/J9wP4NSL1sxvp3f9vqvcWn5lUPvP4uCNP1LtGGRCtxc5D6lb8AU89ytA
VVnclyJESsgIilrkBuZm6Z3roZj03828RkuHoa/yON4pPBQU7oVBZbKgGPqdgKRtbns205fZE0sH
rM2nlch9quGnF/EgsgDxdlFe0LfLNH/w/ih/6qgFv4cD5FX/zY5nJkrMKm8k0aARMN1Rud9Q73nX
RMwr2jsog9Oxe7OV2yIeW7q/JPZzdzqaFJ+E2Ijd37CDcNnZGnsLPv/oS35k45AcU+tH2ACpIlxK
1JwIRJa5Czi8Jd4vyuYrnaldWJFFsF831NRXH6geTfKkVYVEp60vrOZXyq2TMkJId62TZwFfYS6C
se68Px0Q3gjm8f98gIuUaWBuke66cY+saKUX7dZSAof+3oCglMZZp9RY+iQW40u4HZy/Q48kZsh2
o3B5wnW2cxv4YaI48OkCEdTHubAFX8cfkWJC8C6zTgn39xqreJb/49S1b4hRUYDk1m9pnn/98Sxk
vYTAvDpjWFeYWrJ2rA/iaG71Sg22A5dFhkCkSx0pwnL/QtLKSeCjA8tv+6eQkB8qAixbp07jz4nY
Ch0l3n2ydXqMbC3oDWgBmq7EctYNdX9dWtgh8oeBFangQazzRbH2U6QC1Vdt5ypzHftb0z95WWiA
tARloj9wwbWqvFypot6qelFBA6a2pUG58a0coEyOfvcoxKPEh6Mx9OSDpH4p2d23rM6dNOklcWxB
/+4AwUJ2RyT7LXKz1nWatr0mYEg68Q8S+4r4nXlfVqn4DhxoGPjoYVFPltS3LWD9vBaNsyP/UlPy
26U8ZKxhBHpO7p+5lXOFDo+K8ortpJA+Rfxke4tuoydj7eNUhhnMymr7m/QNel7xtSeRtMeqaevy
DjQAmO4ejRo41BFiE07QE7NIwx+bdciI97NRTwGxXsdlEyckDQXVSeW5/5PM7sXAbl2/lejW+mHV
9JT2Ica8FoCW5eEmBHSaNTBT2bJYZAScPqXBUhLQppEdIEXEeBPY2LEZi6Nfq4+xut4fYAFqK8yw
VYBkX8A7qFSgwcnLlkQs61pRKpm2IPm7jXvl2U4ttRxFM3C/mr8v1z0EaZkkcQ+i53k1DDkN7W1B
NUeqD6J5e8RZkFLw8qN/lcocsd019SXJZTxA8T1UZreCQcofGp6JGX9hTeYif3wi77h81tjnBNKg
oCtpSGn7aPeVMBPy3osMOXpQNAbFWiQu2wW50W6CY/yYZVsz2PuURmSF25BhZVu3w4oUcujrRZVz
9r50LiBCq3KnuhZfmWXlvbVJbzFrm/JJHjetv3/kbCZ0ZIc+Oko+J3e2zghtxgl8dx+7VbKOtp1Q
thibuEHMERsgVdqyxIJrkgPR5CVPY02FrT1qHTZiqT/84I4rI0nZ34BDv0oThr6YZYkXwiTcM7ty
QEdA/UzYsH87Rtr/BrXIG+7aLN/EkP1J2R1hYl1CcWuy7OYC5Jw7KXlt5GHH+7xs2Qy70yH1645v
ipCyknCpLIWwSVq04+nkPxY4kDKn+ozDMmr3QyOZ2IViUz8gTRXv+C9e1s0wq+RqMtYw8/1wMe+O
gCmgSHSfYLTgU1pBCerrdQqCL8p+sYtJGYpJ2ynZwQegUNH7beLZSo3mhFZAgPOaW9TK41Y5aQvj
iS9XJKoxtr7J6VjAcaaQ5iisAGRQavfX6uDOvku7KplYAub4z1tYEw5fYuGlZIxGp+HSN3gISEpV
Gae8qh7PoqVXJUWNNncFi7S4kAFYy2ixf6MRsEGHNMjkYM19RqdtCTJDt+mpgjw2yYtuFEfGHlay
L15AJmHkhV7fru0S9RkzFFUTyP2xJuE21YagNbr+GmM8SiKF7l5VdsoxNl+H/2agCTe1YYokRtCz
wMxJkTyUQX16wbl2myehQ4Mkjcx9WPsh/pojWWeluz77P8YpgnACvIyguRbsgDUeYBihzpR6AmyP
dzZSW2B8nNBC7prYdqKC8zOBmC6op2Ts15mmNZB2GWxqxyG3+e6WBrPoyEVz3YxlrPtrsq3yxBpE
0Dt0O2OROyLGUpzByh9sn8zOgl6DY1JhrNAaTYT0eykq3h0ncUwnG2/P6NkPDPVwuoF2tnxPWyiZ
qOBfq43F7sRkULbNSKoP8Zcyz+qPABAnHFGKLbqvP2x26dWo2I/70iuGZF4OG8mpoPJtrAsr8gDe
8iiQyXNvSUu/R9IiBwQk8JHWF+PcKcdaXtwDvrWisUHpQdOsSXrPdZQzvvDtnZW8MMW22kjWa45e
U532vq2U5PcTYuFyuFy9U5XGh5Cn3yTBIjkNAUn6uBRaA44JIvrGpbid0hkItiUav9MnZz8w5SO9
kmvmsBeNAxQ//cxaTaxRXCx2VKh79SS3oljlBwJNMV7IYTqnX+LVKXDCpv4R2t1LKqr+Nqhp3Znl
1QkE6DWPPckSo0C4AkoZLwjUNjEKn0Gv1LILU3He814L24SGkBibykCSfyAsitLiomb9JyGKjsh8
FdNFiN6b4D6sbBNeHIT9fo+xBrDcrSXmS5RUVp1fIFWS7F4pwa5RRUuS9Sp8k/QUzU3Xwjlf6U55
48iwJJ8wKqynVN17CeVpiC5zRYh6jKtMTZDa1Bb1ke6W9cgRMkQw06ODHZ+eCJs5GwUpaqu/DKHp
fWEiHg5EjpFOUF1m0or+tuFCApWzP7SnzEBaOOLDkDumFRR3F/IGl6Ap4FGBlXC5/ZYB9Ss4EdpB
py15GbDukMi3AJ7LJUCaGG+2e3uic+iEulIZZFTO8IA9pOSjYfGKjZuW/wSqn1HB+agy1XT+21rO
wQstuYLTY/AUsoNxgDPop5vLiX6HVP1A6nS7Y+Q7T6H4XxY4H5DvrXg8Dqi01yJi9YgtH7R4z++O
AtIlCw7NqYoUzOw4a7N/PWuLdfB1QoGb2XAP/3Gy7HloOJ7myNyaOhVESMITPSiQu0hMy9C5tzD6
V9dSDvoYUE/DogsWjigPS4G5WE3nJ1CQy7E5qdZRKBHuUun8hkfp6iZJaNnxeRjbtfc7R1OrL6PN
RfZFQBrDfFep8aIK94Y1Ii7/IrbcQSZd53ZBgFr8hvcDGBlRxjEypkeyVw4VGQ+yN1alf5tAo3AL
Id/B/asV/NwJzVF8nLVfGLElnFVNQ6JIFKdmhswvfH7O74hqpL54S3B1xf8qQzRAJsN3zdRmTil/
+WZt8CLKqZwLeEtX19Xa/7AmLLr6ahabNts+agn/F1+40wwx6737cDFNjUKhOnuK7fW8lqZszdiU
Zyo1LNa5Kx4aqJdeXO/WXLELHHb7PIutu4iE8edeMg+63dFkXxXrFk2jLqht6WTtWSIKQheaINIl
LOCBV0BLtRL5hkTHjUX5mTH/IPFVQ9a3/bj3EyHMbrhrAtky3EHI9G/8f4L+xLb4Xf7u2aCFpgnu
fLoMzFRw7TYze7pmn2aoTMqtX4IpRqN5lpXu3Ne9WvnUz9T1/WnJ2IOZRtpPzcfxSqdtg8u+8/B/
AMaEjFXE3HL2BN9SEKYSmDvhUpf5IQ9A6RmC/zAXi7WOXAXAx4ihBR8G7eZcmRQ86/zO2Xer+Tzg
WqDwuqagjzTgqrzZfev/Gm56CjoUTE/RyArvav1zcgxXURTuYcyg/+Bux5icwDnJguuDdooddXpP
pOrhgH/mHE8f5QAphYfC0v+UOPMkMDH+aGOu85Ry7u00KrY5nULPoh1F4ubyNh7LewsquAsFnhn4
YRF8/0WuQuBNqcW5w+858t2OE1kUvVex0852qmtbRCFubfws5H0a52MdUJhlrUFG5vxQsddZN2cZ
JTw6RGFXWucs6MqveEL3TIXLsYF1TNja6awYk+T14kZS2o2gT2fBxHsOhHP5RzigZVL9YBEyfflH
/MaWwxupIe8/y61nrOErOQHxK1+UPP1C9B6jVarndnJEMTdEqhQg/TkKQNCHNb9I7BC0bwdMEbfn
S5GoVFkHF9Zsr4wyKhCUAACzHuwbgXeecuTYEKAzTYdpF+4JUc/DDkgLb+RLxKbdQu3MBXTELBjw
uqSNzibBq24e9x5Mj+mK4si4SBhFkZtZUgJOaalCuyePDCHTx9tB8l3Wy5l1nzdMEoL92G/pSuZV
R290/skNHt/xYnnGnZbg1FAzB2xaJnzZTSTUhw8aMylECqecL4fCtAiDz3U8v1YmcxLFJuDtoM5k
thTWFIr7swxQN2riAkDd+puUv82kCx6XSIEYSEACHf9m8GgZvrQWbrXeNKFP6wcjMjA1rvZMA/ga
rgPMwLczJsYzbgLJMHTHKKAMvy1KsnKNH1FT9zxK7gewSMiHPoNn47Yzjh1NnCXVvdrYrR/L79lp
eYv5tTfiKYlaStEJBK5t17wLG8ToBRWItql7byGKgBBCB3kXaGJkZ+NZb6Cdmdl97oea5t7v82s+
rUmKmtREOZ1rUa1YqfU7533l4xeSNHAb+YzJ1QOdpTeT/Qi/Kfg6oy0jZxNHNuY4ypWS1FIMxBSR
MFvhDieJKSfk2RBFx+VwYeCW+bQvrSaTrrsFm6TjzdwnUGdeAfsH0Mt/OhMMcIi67evbUKuEdEaY
WcgsuKovV1MDH3W5gxO+NbT+bPdgHxG+ZyF6sFiyFia3HDxszOLpLYJiUnGF4wPNEe/crX0bKmES
V77qa3Dd0DKX/bs7P5C4FC4y52/+Uz4mVp9Cuwtewq+r21V2VeVg0cAO8YMTwkI8AZtW8TtYrQ9S
Ug5pvXrYNXke45vswb0GNwu/i23/jVvTGqgBSrZBuoPw1PRzoEuzXBY4XrmIxAOQEsQia73qI/Rt
wIpw0MirpkHZ9bAbaUNf1pzbhywpAOT71FLLSWv/prmcoUuYlfHfA5xYEMZsZH4zW8yEQhuClpx8
+/6AXu8KT0InOWiB7aaUPAjI8X9Pk2kVHTry0gc3EiNQ00na7fEmb6SfKfgpYn5Dn4bwrc0OUGUd
PbsBayiNDszE5Fg+p0ROe2sroa0hF58R0qiX/iaD8uqhL3fLaGPhHFj9P3FDGIUQUcV+p4S8/GC5
ejHlittd+rxftvCVhLP08STME52uF3vmOiTJTfd3oLij3s04sa10s8SVg8yVdk3sJJCcfWSbE5UD
SoQjTIRPkGklBS66LKrnasa3PLOiUKjMLjJrrr1kaozVC3JEf2fwqlNx9jMD0/IXzFrQ6CUZfPZm
8WjwRbc3xps4mEOyBj+WcLp030e9FWuJ3xbRbFlXXoadY/iNipjs7WVygH2GGAM5Jyjeol/Q1Eoo
6qpb4nAX84fwZnyXHMczJbu5+691OhFapCJoAf8Qb3ck0DaSRLqiSeRYeYb1CkPxXEon7O4uwvSL
GI++PKhbcLkaUpTZp7hAmMmPKQaGpMJK7Tdv7Ue4tXb7Pc+Lf4EAuXnKB4AiaKufjYRmQotNjoWg
OUufVHGHJFBJsYhgE1Wy1MxYP1ry/wx9zWA1omAr6qlcVH8hyVnZqX6HXUmkGlF/D++QrXsuqy0M
NVoGzrRbYSNDzzA7UDzMA1hSkqJL4YmH7OreGfTd7BrH8JIuIkDgN4xwuPdLKw35DK7ZX0necHMm
fP6Hnu+znKVUKONM8PLcmtOQHhiCjqXzn0xGQeRyM47sBQh+95ehBJKVuld5Zjoe3QJVYWX+oFuM
syt7odatbufue7DJvF1x2CYRVRE4hPXbk1Fbu/Un6srbVRuQv2Lu3YoASKB52Ba+8qlqVKi2VW3s
KDp+BaEJJd6Jq/ZaIb346+fapEilPjAzRDKVaTtXpBhCtbv/WNfn5o78TYVgIIZsCRTHxCLGQYU7
JM7KezJmuh0c9pB9FbkIqfJkI+TvFetaDpY6HHp6ltIDM6VFGfDkedUU43uc70Yn+C2W/ym5w2ca
AVaKJs0baJBvt2zvRUtpRqLfPmcXmqUspxjl2OiHqdUY5t6jVsFeQtGhhRV6TUm31OOOOtENm142
iIjohHK1eeW6qQ84PxWoar2CuDHmzplnW4il4nrJ/T1o6Uf+2f7WsUT2rL06podl+pKDdUKNUQlf
UX4KA14gSCmP6ZRFoeYmuqSIso2v7Ap+OHP1I+opF17If2hSMnQDZEUdTXQFb5yJQI45iSgSlpWW
f/2zfSAH8UvfcsVLEElnhYLY/4jstJJl0yLIezBtHrIdp0TFFJIvsDLrH/Xjg+VPcXrCywchbPrR
CPkEW5duyTh3cUHAXESunWE9rPVHUEc8NxVdmUa5PA/hLwOxcRNQMqILN9vVJAtBRV0zk8SCUgWO
jH2wsViRHTSikYhrlf4KVemLVFUEsHOmHpO/UoptzhhyKSdM8D9FN6dVGDzcIeUVd2mgsiFut14R
h2yX6kxXQbqeImPWj05bVj8QU6kXfKuFascI7G5XM/pZGlgqfxFe1GfrUrUWTLI8pJAjSQ2dezNW
pJr1bRlTgjGGA+u8vDdXyCP/2G6Xgo3GPLdIbmAWKS+xkab2zg+hRlkzcFYw1WmuneBuCSXcY26N
kTktRtWTN0Oq92tdFbJ9ZhHBXPSpnNqD5urW0f3GLMcpc1GTCFEHTNUYdeY7mBCZ24k4us40o2z4
3bshsPFFttRcdMceJKjpVLbRlyge22wth8muJ3nBV4e/VH/0bOs7lmcT3VychseQevazIzziwIcD
/4BZcBuaV9D10EENDolO/tt78/y4vGwU8mC/hWm7NLIIbmEyjG5/30JXPA7MqQL80mEOTLNiHazK
vK1alUMx3crfWW0Jer68Y1E7AgNGploCo1QqRsUdYeBQWuuoW3Gu+HPNIvd4Of1PUARSMnDfYlSJ
O8atOlY7ZljxRj4sOS78Is8vLmbPgyWcWN4oBr01+KJ31/nkP/ZBuDKg5iQjRPFb+W4Ih6cfAnCd
B/33b7l8mfDguaF3x42jt3urxtMclysNWSH/qcf9196u/tYcufL8QVxonHDCVxNywo15J+2MJUtE
/o9KX2u3Ck+v2YyX5yeKOIYB+1oj7NWkNBqCfSHFScuK7bDr+T+Vp3EQuwIZmtSJ4AOGWRUUXdTj
CSFwHC+AIDadXwwy/p+9Atabg9je3nj/qKxpfOMhu3x8GWZmZBCtVJ4fdBd1+MdfSR80DNG4528S
+SswXUi9oai0qpG6yY++RdvS9xGdKMQpguNsVO7eLb1A/s4KlBR0wcM9KNNzukE8dNPZNMWpaqhJ
g0QYADsE722e1QS5FUKVoMzYF7J6Kb4Hv2zp/HgWde5vHhOmGLqOWoZ+RzjnrBKosvfOc9AfDeHE
u2SYxTGW3O/g29fXGgtu3OSSEKlYA/FU+xjRAlQNN+BYN9GdM1SdGx+FfFnt4gPEQXlxfl1D01L4
80g6YHdKsOCW+91qwZKbQQpQ5npAnrMONVf07w1Hk9rJkrTpKZcUdVb5PD/FCzsWPNmQx+Fw7DQX
34s1qUCQnwQJ46epkmCSSpKVjW12mLMcKomyYZZdIVnr9kFFdLPW0jbuwD8age5btiolpq/ib5yC
B/Lu5/L1m7p4llxAxD9qKZJ3luUqQbOVFIh7w3V0gyu1v/gVQEda6MnsUTZt/7XBkbrcvHKx2Zd0
SpsDvwCYyY/afVHpsVubxJuV1IEZ4qRueGPHaWYYdW4xe6RIKo5s0EByq8SmU/1u9Y7bVcx65DRM
wVGpvYpwuCf9aiHchp1isBdyozMF5YjKs9WALpPbQpSJuRDL6xDjSFdYnGEW+y5CY3Nj1GxVcuq2
wJitouEvZpYqL/EWi5/s3QXGR71JMCpoWkVoWcO54UYqoj1hl9ioqZ6IDUY4NsNPtK3tPzcqQ4Qk
13KsNLlvibp64SEXqOej5dubqzWos5NPeKDglXE/MP/sCXSF0XO3atf6tBmtTlzP67iv7vIYgt/7
Om4nwUCXX5Li8uqT4nWE2cGoucFgDHFBXiEGAy4aThXdUFLLxooDsjshcNimTR3G9zMtaKl61GAd
FJXP77XXWNhQqUTicNFf59cd8IJ6HaHeBJKgv9J5xSmqL8tqknNW98nZrWaGHA5x73aH2XdtanA0
6c9vSG0zUl88dSkMhuYsO2wtEpd/XOISf8rPDhGIPxkVz103A7u0GlWXdrFSBmRSkZkWXQh/RbaZ
PnwfCx+FFgTDwF0ljHrHUBe1YEUvl/BUY059xFy6GsuBWXLJMXYV4P/I5xGpK5KNY/WLg/lBmxuN
GrLQ/Iv9nuSMduG4pzhyQyj8mPJuSstrrTkVyfYOCcr4JgBmNiu4dJGG7Q/bZ6+YxHNO7VguT4It
O+NEJZYXrRiBbXZYzSS3s5A5CRphJ1NDrQ1Se8tQRrqQgJvrHsX/yeu/yr4DG7sQx+fEI3Jo/Ms8
bo9paKd9OybtBpGEuuGdAbHoVfVwCkztbEtiyR4F/OlbQpuSr7wHBdU7Q9UXeUi+MdP4zShzw8FM
d4Yx75DOtyw0EHh+AeMbx7nN6wTbN77Svkk+kXGiKv85hloALny+wlQBWJ+O2jrA7nd0rHDF00Hk
J58RGrFNsBbOcVX++2P5wbmRJtiyCbUqJ+NsjfM7mfhGMHa/E2hMcK5eAeOT/efYp+qIGUGG07B4
2KKlru/4qiAJIYlDjqeCH4mmrnDkX3BrbQ3y5HEiiI0cFThbNdYfy1LxI4t4nzmCNVb3Anca3u1q
GzaIhf/vUkYrBNjnUYadJHc522KOteXANC8pY6np870mm8k8WkDmsor1LSBJhGlpn1BhpGrEvWXT
FQS/AMc0rdkPIBR5kYfso1YniiVGJFKtic9bjQcoNWqOnBfrT1A3DSnbFzpnJ+ibaFOmjWzGYWTz
kNAmJ7v3clMdbsrNUTLb4T9vlUX/cQF2MeOvAFji10iGWT0hEp7klFtmy9UI1Ez0aTneC0kDanx/
Ze11lN241EZ2oyGSdaBKqu57IrBhAfn+2C56FiPHgi4KPnHhgn1RQvFVEWS/l4PYyYc28tFyvlRa
icYlAzSWTtYRRQyLuugtJ2GDWPYTLLeeAn+tJ8GVex/blGwCGvh4ylVSO5qvLbML/TT5qE1rbT9m
xthZBWrP33ZkupVv+RcgT70vxJQnDCFdlqEMt5aCaJBkmHXwK1+/PabxMKamFAnxhU0PmU8Qqx2g
jiVPe5DsNLFV0dy4iHLJO3h7OL/d91tdC3nP0WOtUpaapd4BWfwSJH+JKfwdImhMwrKy0eDUZPGl
Dd2CuOL1ItGqcLv2xyaRv8Qk3KPMz4iUmG0mplaqES8Z0RjdlDtRfY/G5IlhgPssXvqYmjiHn9T6
Z+kimq5udMrDX9IhPMqK6mSxeeJ7cStJyP6thnSaLPdtSA/gyDuu/pcUBlDQfFuqZ8ppMJLwvGY0
RsxcLmJfRlV+ZShtXMxmAJmluNz6M9yDVJ/5qvoHepAIOw+BUyjat27g5B6+/6rwpeDcq9S4K+D7
GSxKwMrQVYtG6wh5MNBGc2+U9Xeu2Lgjydl1M0R7nUd7PzjlBrmAooYzcTKURXYWUPgav5zGHJN2
1eSqssqOD0Aa8y+Wrmw1JHoV/BzNMGIC5nExKtdZHQFksypLN8W20SUqPCEg1hY8RrLF3JjXNhyb
IsRV+IPGzEgiqFjzonYeZo2zs+zYN6eoquNDFsucDgPXiwS09XAAOEH2QZbLnWZLz3KlGYbEeUD4
Q5MI2ne+YlexnVL4eauJpKtwurGPbhO8OmEGlInpZu7f4GXDqwTaAo5MfYBZOMMFV+xSxUBh855B
95J18g/O6xAKaJtISv4U1EY2atPjnAT+mlZhQAdHPHykcCJEn6P6GGfMbX96z4ijuzwlHq4B7DWC
H17+NYVRy7ABXI+MeGdIQFYxw8dagUJSvjjm1H9ZfRGJEmxHL1PqzlkT3cOouprzZd/HW34lay99
AbYsMhigKVrwHN24NL1wxgyAEk4S8RI8KhQODmjWjF6ASM/lSJTmsFnouf4I5mNcZz+/U9HOR+fJ
6ruCPGVXiPLnBMUu2uojJfw4wOWwb0oDs0zEiY/JHAu78KRyVeRNUJ6eNbUF1I22tZtACJxaa65z
HkW4otLCyMl36Ua+qZyqbdxLx3p3C4KYY0XWuYg6NRB01tX0ak6SO4ODjjeep+7etGwWFWY4LSVB
AIzbWekETLR3lRmYtjCBJ9ijmCiQTsAODQLPYpHcUM4EOzmu69GQ1Q3lBOhppKd0/ymB4Dn8GgDi
eqFKlgsrxtedpwB0AeK3H21Wctu4N6Gin9IBQinp2bw4cg0dzsGIGgfafJ1h8+DHiKvE9TCCMdNY
IZzJVsBUF0Cfc7nYMNtczTQkXBA//Zyp2tFe01aY128tFSPBzb1FFY+xwD7QKoGAarhFBiGO0hvU
XJ1IaX5xU7r8KTsxWKpRe6HQkKfQfY7jiNvyUgj/DrBOn8bpLuI14hL0ZdKDOJJxbUgsheGeKdCD
W8oiDKPUl/3FbsL2ce9GkoNHTWZ6OGK5ECj6V9+dQz7G+eCuL6pU5MRrQ3toaOvdjzUaGp9V0h5G
5w3Ha1Jwr7bPMUDuuNHOPaVKmfTpRZclpzWvFnld5ZDhAg65vAEe+Nja4sbO3AyH0KbO5i/K/Yao
caymIMWvXtt1JDuvVrtFOe0ZpPT3Y/n6r3QBPhqac5jxGlKqvV3NbWmznLtFcSAXHKn2bwcEDcDT
QpZncYCCuieWabGzaLJT7r+CBWlpzeWjmNhQbzwmLa/MNtzmz05FJbOyWiARLJzRp9YxatOw5E+u
dzpeDnz0eLuTP75VPcuaCxWW9YBS0zAm4mhp12NjBVniU6OSu9W5Nal55ZeiwsePDg2NSMx7MVC7
yNVG34JrzE1GC2l7cqF2YdLI5Swf1fnzet98En2AzV1aZz4X00Zpz+f1EhmSZNoChnnlbz5wSWAb
sqjQ5Nou8Y2YVOb1z3mEfFPBh4PezJu5sdsN2NcNUlRGktg1HodhfAorc5miGX2CNyV5NwuSJxxa
afWoT0vgWJBHJ6xv30W/85oTjFwD5q+D2aNIFsjmeWkWk4JvsFz6p+16m8tYxTL+4D274/H22ojq
1CXlBBCsh3aqeqp0b9M2ShrQDfzifnbnW+y9Xx40FqFc6jWPvJJQTyO8AGA9kZlOM7tqrg1rdpBL
/T0OHoqkZqdJe8+pU5prZD/dHwQszFPRTSiLcvFomDkqWrS5FPEqHHg96PdGaiSvz1s6UP96YRTe
WWiZc4zBUNiUCcc+uK6oFl4hmBZxUSBoEAqQULJWaHtdUZTCQbHZCeGS7myDifK7iMPoNnneziGW
xJueIsr0HzrpqrIA3tiQ6XxT6xQ1aHuGl/5EzKs7Rcbs5FqaOmuNzbFNQsp4lLrfEVIGYWX0m62d
7Kusni8QN0Eln5enOA9t2f3/2k7vv0z0CjDHGfhvl5WBULiNJGf5+2koGbT7/MhJFH50waRzGFW1
Ty6tmmPnTPmCGYpIKN/Qf8kOVapGR8krzm8FuBkUvosjUQTdaNpus+Voc+8jgaGxFP39OaFKe9/f
NZa1A8fKm6uVRG10nY7TWT/OucLlvtTxLPSQGJKgIHawOgz7gb+v3wFmtZff1chBTvzbo/4niJZt
3F+98gfIoY3gDoIz3kEFPl9hGwVDVCc7B7m/OJdLHdhmdKpGf/0m6NxK0naaxUhYrqR+9EKAtEKL
Th0UMNC8j2eJBxAB6XUU+6D0aiDCgHfM79rMbDD/lAa8RGD8uGK0NCG7sGImd0Qk3PvRt61fdbGn
L49HHG2RCIzzZWm9p90XaPbG61agQYxHPGAj8i33SKsV/na8OSfeEPiBijWX6OfbHQFFd24hilZA
x89z+kPJ3CUnoMJu+nP6GVIXl4LY12UycYLnGjBO7eo+W+IeILGXaIADWZCUQIdSX7tGXLVTVaKq
v2EsSECxI+NmEJY4MhTY0xieCy+ZaUHo32MLQ896E3AIYjDAG/w3DCbE1XkAHQtzGgw0cqotjYwm
Wpsx/LfrSKrrBb5U6BXvKGJRAK26QV7Ydd9V5UlaFyDcIEfkQTIuvZ0BiyHbzvvz8vhli9dZrzGA
A+oRnUEtuNuCcEZOojiFpXaTfZ742WZmFUClp73hkHgYwEmeXwoEnsIsAlU3jEuzlRaQNnqOBONk
QPlOdMbMncVE5bBoMGZs0gXlM/XZ+r8i1Z2By2RgVLn2mINL5L8d62DAJuEbtMFx36mOUYKGGBi/
K3CKtBRWuh+yIORsXgNHAN19CNmzKiIQQyknmoHX8CZgISlHuBqwDpUSP0iDIkEafTQ/zaTVa/Qa
Xevvc0QSTcVYsg7jlQ3kwrv5g+/QtYBwJKZP8vgb0bFU8vrFJ+N2gGO8FpIhdLfDGMheQ7NBH/fT
hKhyAGBEDJS9aHTP7CRwLsugaX0lixU15QNpN4C4AyDRdUQKC/eV4r3noaUmr4nINzQdGOEX8BBS
+nRZirbPFixUznIwJALZW33e60SIlfwIbweV/p+VsaJEjrhk4ZrmmqMZ/jhnIvM1HPDsiCDpbyLI
z+gXIjvtgE1/YSHGUDWQGt4LaWyIN5CcIkRxCXYESGFks/kkUPUeTs5eOfEzaka33SV1upplvkvD
VvEM24gSKX/p9HYIzYzwWkR54jKawoUU+54Z3cc+/wpw+/WNn2vWfBfkVPe12xkGGtm0PAWXUKR9
Ub0dwi5bU8P7v1ZfNuUBikJbxDT0FF2FfhE0Pd8jiEYzmRUAO6UOlnE9ULRRtO+TP29mZFFte7Cr
HmHvHhvh8ZQ0MaNFpH4RT3qLuk8Dehd+SonAhdvVwDIVJPz+yq8E+eADgDcCLHf/i+RL1xxcNhnu
Y8+/20cHdJvJR65XdvpRQIha/9NPJHb0cHczeE0fV4iuIxCNBz5HG8Hk0DC7vfpV+siPG++BhVgQ
vCfsbknOs/sV3hBiu0brAmdQSZD7wkva1JHdxMi39/w9j1523Zur8LhSqfp5VtZkaTDkEdOGvbe7
dvHm0GAMgGQ0GZFhZwSI2U5szuQ2z7kXeaeOOX9UVbBpYdGJepbcHpFwpxpwskURs/k7uws3QzpR
xsH90yVNdRxNjK5OpRRTOSakqiLcRHkUHMxQjQQaMlJyKnPAvdACpsTJfWoWkeapJbM2SO3f11Q7
SRwAFT5drNPrFblJxoGp490xFm3jhvi1yydUu+4nhFPtLMehzkqzbSBMS/WwhaqgCUI2Q4udfTwa
kieXdLdNJfMYTZl4UMjfDvqcUJht65ufGZyzlhtAaIspXSt9q3JOyH/WNnJGHsmSQ5Z1a5uRKZVl
DNz0gCOJzzOOiFZqEjP+RVzjuACJYAIIZkCC8rWwXTVkm3EirJJ1JUK9GV1QmkluVVYEtxKwUEXt
kKJxz4CNZdlA6hL67l/MG2ElD1/MdvQCD4m6tKcJL9ieYV5EkR+4OzEwO/n47M3+BSae6E9bQCWP
7S7qqwAfCzYJBIgC3SPnsr6gyLgV4GVYIWrqQ2f83FBDVQ0w5E2vpnO3Y3EbW1PWNwCvIlyU4iYw
+omdJ8Z+ZvuErr0DI7wHHFGcTgH6+/GbP/RlyvqczmtCzLrMyDCe/hAuNC30VlAwuW4D5t+OzbBr
IZX3lPbxBUZaJHqckfjW4CXlkWkH/BdrkknRBHkLgsRWfqOvcMwUcMOOrPgxrsO6xdQZPOwgCI0Q
YBL7VKSpUfDF6SuxFvkv4UfEvVqjXytef3hkCI8McjywChjBexFF/T7HsHFHu53jdsLFB8FmK2Xu
joX/qx492C6vEKl8VWGoiyGQHyGiqofzekXA6O0C3i/lqd4TwYJ6xAk3VEzVhk10diAVNaswaR0p
uVhWed7XLS3QXBTsBv6AKP3dIlPHniAUsBGleg7F2mZw0ERu0u7ho7wsCV/Ermc/9YUCifERFbEi
sM1z58FDWFP066wmNQ6RFrNLJ4BNSbHqILr7Ob1rmIr0g9vg4/Gb/kuhHkquD8CcpC1skayaRbcl
LsfG8pkYZEgN7ypOc8ITwkj6RPnbZq0fH1ZhGtHTJO669ULnEUHzJmvEzqbpLBJhz2JVQhg+z8RI
RjutIqScNzC9z3POf+M6ROXCnSBvvkAnh40VnyM0K5YTLYlFldyNPFsC7m/8PATNdEb6gSFSueWX
U7Amh0O3dFhE8HvQH3ih/yPgt3+kRIb2/0iPbM4ixW6IjxBLui2UvaSs67dd1PBEgIEnQCb2H508
dEp0Ah1WcIUjbPva3FrYUHZmwC69BJOCfkesctcg7AuHPR/A586qxqf5AoKGR6+WTVhF/FD30VTL
YsPB9Uv/K4Gz47JoDrpGAbNdfIjY8FuLsc3IsB/d6hi2mQu5ienEj078bwSR4i3nLl0sDr8s/Jj1
PzuxdYTOhUDAlzfb9i4kdcb4Q187fykg+lj2bx+byh4evlLxX9RAWcPD+YaJ/RqmA+jm8TE2bOXq
xHdS64ieXDsE4W81KB7q1Gl+plpJMOTHfgQq4iteaJnXqZ3DCdLn8PqQTaMwy0RkO8okHp7GEMzi
a8JYkFAngQw8Mch1n3SdWOcpDBDbZSjs0jUGBA947/qAvQyANK9O+/7ej9sexUQZMu3q8oB78OSV
5U7vekBBPEXxApV1kEGeD0I0SPjtof5iVCq6h/LUrnaXkDVsiihc0zwez8aN0EbXjN9u9a+aOxUS
PFTKSKLgqDZNSrVdDF7qJFZLW7xTvdr2wSl+t+E5bhA5u3xZ9ch63/FalFFuldA29/gw1B8sLTu9
JB72zYyXcLFmOapZ70q7FCyxQ7A792cxyxGcwTCfiji+YKngZGlSD04xlVnaLez8rUbOjl4RbcTh
cjzlGd/fNxPsLIAelQmyQpIuquHFEbQnbZhY4+J1g6ZCTin42ka+VGMWenbSWUeE0H6KMrJkblUp
7LlCC1oDnReWQJIDholEBMX7Keqc2p9U3PpviSkWQw1/3T6P+mffCIZ3q78u/ZVF4qCupcSfdaBP
o+1A+8H2nSY+qQyGki0SakBYj0RWWfs2cIy8mlnAzZer3ACRtW1G3X4/5C5R3n+E5w84q3A1CAGR
EymvSFF0TnlpOZCWHK43pV5+Val/ixIoEughJADy/tJYktWOTXR/xIUPyhD2onWA3tC77WVkQ7uA
kD9+fvXQ09YXfdoQuY7R8DSMhRAc5ldVangOwE08RHd8pBqNyJr5EVaOrLiaXXuvaE/Hls7oEAwj
0wMggz//5hFWIX5poXOFMbm/uYiBfl4wOnDtbVC3ZGFVXojpvIgndO9/wNA3Ejbv2I/5KuTNXyRB
dLpzcyXz1QlO9WwNEjK9Cpa1XuyZsJMOVJ0tT/hgNgibASVKhkCXL08xUXwh/x5n3tSNE7JKGtBy
R5fC8nMtKEwm6sGKDJ7GHcWmP5HtYwGeoEgqmoyLh0IrFrEYz5Y4bDby9GOvjGvF0J+chsfKQSGv
O4LHtPga1zsKmOYoRW4a4UzVQzsdrU2vc9hlpRwP7UtaYpCaNx+VKeCK6s7lm1RdcbM6v9hM69y7
G8NTOtrZiOJdD7AsU4cMcwo4yqjuud9tR2EcYsNR8mMPeePNtBI030luZMu2tNmST29vU3DkUug0
X26awtaFapTS00UKOexl3eonCQdZJ8XByKM1CNZcMtvKn6idqajLJPUFob6TCrmwNz7idOwKrP6a
ysvQ5rS8j7URVsVzpJrOB5QaJktGuoBXBdihibr6/LD7NbKOaayJb1FyJJrv4jLybUyEA1IZl3v+
pCcmXiiTWYzjPJ6Snam2s4g7f/NA4/lVyhk9JeC6Q3OgPAMCF7M5K4NN33LTLK6c7GtX7mXB4tfs
Fyhr41GMscE0L5agDGznXCBB9fq0tuPaAX9aYMuOvj9ne0IQIvHdBelHj9XOpvchJC19MiFvr+HO
2xsJ+bdnyAAVTuZBJ8A6K+GMJ/lwv3fdzQn+tRSp/EquH4RSCAYDlkC066Oq/dw9l4+dveRGsoSf
T/xZu83P1OAd0qKm1849gnaLDP8Eh1eZXZvXaBXENfFFnyw8haRx6tpBQgMMewSAmiDuZ8RJgz6Z
lQfvX37Td7tqsI3vT9psHAtUw5NYXdKAV5jHpKt6FdBaycjPthA4NiuOTiJu3tV7w3iVgtpStDaK
E9DD7aI1qZbSxvLNF1+U4vd0HleTCqG5OFuTMVZF6FD1nHAapl9SHFjNzEVG3ff3GJqbPprSlcpn
nu+mLheycGIDWAx5GM5MpFNMc5zsu0rmlHGA5Ls4koATJazlQGEyEk4R3pLPzSNHbz8l/UxhUpor
66Or87+KCoakH3y8ClC+zYrrmT7tPy8RD7mOwbs6EjzFHR/jlxgGXU5fdW//k0GO0VG1QWONtI9G
nIzKHRYYA02Y+K2M/0JVI1U4brbNnF/cbW3O3c0fJYR8ybbJ4YLbU7qqfiAdrxA2SRPt4UKM8OW0
X0HU8szpXKBz+g1P6yF0hLPqJGDrHigYM82u4iVWwnOCbiZf5R9ls9nYOhvuwsxvjaR48KoRRXdM
f2q1BcBAgjMtqiu/DAyagQQEdYQnsy0PvpEUG5jrDPyTNFZyATw08XMwJUJjTF71jYDtTlh1CIOG
c0SWCZkel3IFeQmf0ihv3Dr6A9qNbCE8dSutd8Ml50hJCTv5ntqJTyYNdfK7Th6Sf6tAeCTCPgMK
Uq7i5B5EOdObrvGbtMd0gKK3RXr9GJn/y92dC/CDrwnKGNPRrLuX4bnxyi3twHl4STFO88b1zAcK
J5i639XbUzVdb9H33QfWMQaS27nhn0VmRtHXrEv22JiyeqjXYyuyO/39MpHTAh3giSOIR8Mo183c
pyrAUb4rksG9ZbTHT1CS1QOz3JGQg4tQo/FpeT3lzl5KFHHF53oxBl3tZo5USzW9lU8xQhgYLPxS
YjeymuKdZfwq6nKjp2/h7527hZbTZLgykQlIXj8WNQGaWklCKA8xNAXnYK7Houhg54gL/gIfPgAD
czHCVXwJqmZB1XU8K3jsGxGoXc7g1DUudN7d2qNVNbMxuRU+hurgabwHgjUIc93FxnpEWxI2yquM
EIuBpQex8AbUsdJ3gdVKy+KMLoVq00j5X8ECLa+GnOF/Paj07aMT5dTDNFUKfun4d2dTFiEb/Qpk
n6aGZVpEyBRfJF5N6pGjJWwx3AS5SvKP8SrD9rEHHVX9iA083wjo+/bBEXJFtkntB0o/WR4ltjk3
lJZUcZpAanVKgW4kaVF1sZxiM7QeD6FBcmdZzhvgK9g2llF00he+1bxzJA/PLOjVycjfOkWVdMP4
mVXkVPZ0RD+6oYDwhDB/JyfADiZrqaRCF6eSIcDfvfHmkVd+fu5Lt4xd3oaTbaY4BfrqCm4ZnvNl
5EOpm1CfNfseT3v16KT5k54/sO61d/jpZ5tHdhheBory3hFjW/nIQpZ8CCLtTVcudX2K5N/+OC6g
U3Cy1RlHH7EGXPfodI/NfijnUju10+ONLbsn5YVnLOASKdu3usZ9hcN2j9hQ1Ba8DEekS6lVzdk1
8VL2tD5fZg0/DEt/HhbCfBfqXwcQajSVHUJjLrLmigS0roWHCajltn7NC1fn0fdHTz/5mTaju1JO
YJonJYWxh6b4IqBq+1d72FgaH/TqNV0Ho8Q/brhGu+fGb6p1znLny7x3JRuAasSDmlfrP+jKtDsz
+I25Vgz3gRmZ30L+h9wmVl578OExRyrR/hRzQlY29zwrMfPMBLCqIR+AFqbbBm1QmBMa1ZzGuIYt
UBmFbocVRFAntx402hZePNUU+F8/uCOjIK3LY4ktweP3IfM0kLNvfWo1rHHn4DXlNIsZmggU54b/
hr5bdLiLMdQT8Fy3vIUGOknifIxfnNWNqPzJHoY5AI491YGz1+rYQOuSG2Wc5qE0rceEG5ZlUi0t
sI2oB7DZIAxE4VC1ytokie2uViSisZ4twxefKMFdVot0ZObrrO1/PcqLvCef3VEwlxA4Gu0bZjn8
oopb4J3At7BUVmTx4zBiIW4BbamKKC/Xi+7tALn5petCRNyBMCUpBdlD0bOLic6AxiRNyvxTZ3NW
FKWyihtHXs4QC43THEGcbl1WYy8wUVn5uhig8MyNNks52nhcauxzDNk1yfvbMnWozLtuA+y6njY1
NSBBsZFCc9hp89mbG+w29oAawJrTvb6K3nqNSczQRl9xCg6h9x5/2GTB7n0sDRS/TIyzRNvsp+ms
PfUuekwBwJ01t1FOUpH1gd4BFjXUG0HECEOO7d5e0w5T8DOIDAvypbGYfa6Oh/qo0WER1O60AGbM
scsUs845g0hvUoZWejnLTtZOqSDFR1elWqOK8oj8u5BhGlon5b9boyywD3JUZ+ThVYpwimAO8sEL
D4N6pwdTEZVQT+/tXXw/7v7U2ijoqh8O6F1weDgnKTHzfi5wr/PCv56wmR/6nPmOgA0MZahUwplL
lEqfbvp99rb44auNiL0jL9xoOkxwtq/VIKGGs8B0qt3TbJtTCucPrrjOhp/oGrytN+rWxKJIfZl6
vkcplof14BH/nJwlb0wpCqzyfRufPN18trVEnv9UW2vCGrksn8PHxMT/eRlwmkbVAoY0t1PGULVI
1FJOB9gt3PtBinAD18QBQS4eqh8lWJX4ximNVkbYY/6RsxJDYcRxAWS4B0Gsc8dUnOhFGzidWOdS
OStKFeJtn6iE1h/IOWROCETrCcPcXq2Z2Vsc8J+OiYpfTsfb+i5n9zQJn4iO35yxJfboJyIs9ccS
1p/JxyWZxuZCIXtqz0lmRwJCfUuITh/ip2XNAyBUmWGTgAyfRQJWijuM9JGMVbqKxNUH1OKCwCoG
w0x7+7bGiSmupQ7cBgVXsbOE56+krCS+HZZFYyGwzbJ4hs2o1xdIkFhsxaeTTE4pQqEol92CL+RB
ZBceFlcds350rFeRi7yzxhsouO718l8ttBONkg0JLfZcZq0EZ1Qhn4XtliS/frVHCIEaXWXJU/8n
GNLrzbvPtX0xQ194Oc6wEoY3IrnVz8v9fu+s8ikfLeJhpwNzZsdtBUm3VRj9hMPluHhMCyUhZRj6
oi7XS9Uv7sAYGP7bhUWgpK0y9vgK5CD0HGnyRiVpK9fPy+G7CrGQZS1CY5HR1mmRYTUSt6lRqs9F
m7lxlqa2ulNGINg6XeDEenKiKhfsse+oKUNMW0faIgQ6XmAn2jsw2eiGDZKxct8LTDGMFQl/6/LD
UgSmI9Y8cB/3UZcS9vdLhgV+bQTI7lrwyYvmWHQE9a6jNSh/2VI9aHBkVdF6D+N04u/AK6tAKgWC
wmO3+l1UEpeDaHxtqC6+EUF6q+9okPR2upjtd4dfMhjmkSrcr1jqboEmFREconz6WJHnkOHpHMIb
+f43sahx+FzAYvqgHB+kKNYQN/GAbIGD6Bm2mJqATtV055cVagERQqhQ5hCvpd4C1ncLaWackhx9
AHq+nVkyfAnLcY/8mw9OTo6YzN5s2VGWi2kVOKEj9fjc8ca+Yilv9buS4dTy+rueEFvOOiC2okEq
T3Ka/A5ETxIbKtyMSRvySIcuYJwEcPciGjcxJQ/STcLkgdxzKP4jCTRUFm19+dA5LHqwgz22lMm/
XUrKb/3nmn+W7pM2tT04vhF0ODEtdHIJqueZCP19GSiLfPbQF338T0ksqxkCHAgaiCPSzVKAte/l
oZL75Vn5zub+fQb1pXl9LVp5FJV+Yx9BJZvHNUksJD1N099wXw44/giP+owUivCnybJ5eCXz/1bV
LX8RW4EtBdgRcM9VuvKMV9/GrlX3HqeJsWueoU7u2tRDKp6wtfG/CJ5nTEpQiVb4vKXxhxz4t3Ep
apU8zZSsDoPsOiLWeP3CtfykPf7fvVoEr6li5M+tnzMzfnN9zbGoKf5vQKJ2Hl4zKW1di017pEB2
gFNhC9woqA8RPRqfdTkIbCG5OEVnc2/BRwdbBQAUfrB2o0KyAO1+MxCI0ZkWDjtaeoq8aihYbW0P
UaHjHux7VCYLQV/Boh4MG/74BvGa8KgqB8TY57wvk8h/ypFXNTVblLuODc3hyln72vUcc/92qaIj
q6+t8Z2a5FiynjKU3Lbfye/RMs7eaz4GW3KdZLTat1e1xJfNGFeu+lJ7L/Hrg7HNlmCLJ77rAKek
BUxBym9TteZvJ9NzukFr5atRfGqKYh8SVWaqWl0dmHje7Zz2eoNrdptwQhz6w9dlyadt53yrwgSS
MYQOJ3zNGmhm/dZEzsG0MwLXnVSXss0Zkzy9ZC5k7epnjrwXVW+NSA70AJNaIybJRzHGRWRfZvQ4
3GZeNY6QdXCfEEnWpsCcPNP0GPSxcEUQ9aoXEUk2dlCIBN3MZ3x+5IMhVtRFPaB3ySN937Lla/Dk
BvOCz57CMur8+sSeOOeMH3BCtznG5TgsQ5iyPjxj/72SnVoUou0jXJPAxByMxjNY1bjDNnju6m/t
2SJxeQtiwiNbeJYtH3+lGRX7qBu+BRQWewbFhOIX77hDwweT+iSZrZVtVMOJvt1RILZLbCoON2X7
LWSeHKYBcGJ1hNlTp1vkqjr+D8PRgxcEaTCTyh+lkPkCtnQGJ4rEBlUdDK/22Yx7XDKEZw2G2Bwr
cLm/BMAn9wU8FZLUp+HOx/EH4DbAW2GHbG9efjoWx2czUTbiHPlL3nfKRTxjmT3HiuaVs9CXOYmp
J12yAgQWqwBSdKPN3OO9uX6GTNRS5AdDhw+mOEwKVpW8G4CrNlumy8CrxHaVolJh+OZieBdmIIbs
4/ixDBgA3Z1LCtKmFbQA3eSxwR3wmCebDep4D86VZdaxsJ/ow2YXtgds78NIBofPe2f5Bd4Osj2C
fn+hUjlvhxb1Md34yiVKrT64tRMN0Qwwz/HR0bL6ghxENTY1yVwtJiOeND1xmI3NS0UNuap/Z+e+
mEPQrpBcezz7OsBh1J7qEZKEiF7lxJ4OgRcKB8Zf9NegTVRvpbWI6E0BArkf26knxBe3F4zFE20B
frYhCJmRizqfgwiNXA4kPAoogumN5SwWi7aADJ2kjBzJybGiBYyAXspbowJxqedCQXbwAIHODOyR
im7C5oJM9XMaeRy6BtxRgDM/l3RRTcY3Eoq/lDm/FPj4LSKokNyURW66VbFZ2mXgVMwnFZZHhGe1
fEdc+imf+9kSe8LymBeZopWt2904ZgU2jcq2A+Abp9gOH7mdsDL+I8am6N3uiczeP1S9QoT8+juJ
eEp3liUbtFEBQE1B/HtukbQAni6Xxy+3xULcEoXlwqur4bb6LeK5H4llotFVcdOcemaZFojzjJ9q
fZaKuIdjF6ZI1ksBDJNx9O7CLbU1cl8rBp7tr6FiGyLBzeQQ8AofLDdbWddU32gfdQ7SDAkthbLe
umCr1bzk47tETALozYUlq3kRCT7m2aAmTDrutKhGFW1IpOqAw+yvOOrBM6WZ+KKlu+ptupNoxJVu
fDndaBsSqqfPnKIE11/xTvC5hjdhzAx8o+j+LgZg/ctrVNYSFWFQpCz7cldy3AagKVmQTVhbeXop
YHFfSkNCSEskdjehrHZYkvRnS9WMCylhnhhLYxIBTcg7dosfx0Yyh2v3+aQHIlfRRIuX89DtCaU7
/rFHotzv9nWxn6mSjfOSf99nzYA4lDtVF5ET/cNyGcVHIxbYLV92HILfpaApmx3WdZTu/RAQ8YSs
4N1oqlZ4u4m5WFwZYpRwwcUJIkzvE4V01dkhuBF0o1pRgd/qDuPTiXI8j6kkcUIPYifGZwbB+lMa
CO1XlRMiplOfJsI7y2HIyKBYvE7l6ecfEiAeEEq+KFXWOQ4GF2o4XFVx0Qa6zZ6bOoZCp4bdzjPo
t69b54oOLEZffEUIA07eNsZ5NFPa1U8p0xWFhEPQqqsO+7PG+5Ie4dmHtb8ZbvNVedTAc9nSUAPG
EHzRf48xOhGo1i1JPAo+XKruu7beBAFdrNB9A9t1kH16NtbYJU5IXTo6kTorVe32a7ZpWykZGYXA
Yf4hBy3f3a+DhWjDg2le1bP4wkxOWUFtzNeoJo+OYGrwlPHpGkRmPZ+8nW7k8atZ5AOGEeRNjd58
rLsDFpw8UvxJ0T8zixQtWi2znboV26vWbic3HtAX9Wnwdpxh9CnTzygDox8MwIORyU0z9EFnIpyw
K0kGcthJXX/7uDYIxY9aLxAZ/Jnvza8N4Q2DxAZQMDr8LMGWAoGigMXqxVg6umNDQGuwcC1w8tII
D+hFDVfFlI9n09l2u5Pw+YrGD/SHvagD2uYUNCvd0Z1iAlUaIFPoCrqedfzU4KUFQA+sV5Swznfc
31fqXG0SgO8RUFXQlfSbG0CQHvUc+neK33ikAOBJ130yB5qH6ryaWGERfH6a3+Z0uYPMLQP/Tof3
UUbx/KCXMWJvy9Ic6Mo80sea/WS9JH26q7XwxvdAU9QImlLZoyZDt1fdXYTn1Atm41xTuXhd9jNU
qrkdHSfhacfKwRXKT2qS7rxDd2V6VSp7kb0r3FdOGb8846bgBbfmkRN602Au3PSylTdfm0ngcY3G
cxobMZIBwmegA+CID80WE1YiXMXwA5OOS7KgQeLaHxiVPMkZkK+tMglyBGBgJ3ufxkcU+GyOg1pV
r9jhBl2RgL72xgFRQN7x8ftmGYtV5YFyo/UhtlwML+YkdTqUebJEfjiE03fCMrR08bawxbdcBjA5
90iv2ZT3Wsuw/qXEsP6xiY12p7AlOUowIM0D/gaEUh4xZKiy/zK2ntckN4dCld/u9enVOywHd9Rg
cFevXhJc/oAurNCR3tEkGgBZ6JcO++En4uJI/E8Qe5Bm9535EvkDerdZGl7aYZ+NThU+aG7aVA/a
Pr22TE4c857RQ+6dxlwfRT7ReKFqS6W5m5wZQCaEBG9npOcm+A32IWSCt8toRLhCxBrfkXwZqwh/
MvjiypVINUFO8Hsc6Cr1fJm5gdSXeVyujUmVIMOvKXCvohqtgXkfll9RtPSBfGNb1+Gm7AvhxwYF
i6PnI26CLaSshP58L9ORLM82d7kRH7Aa+MUY65KKkmukABLBsvJRxlEIEityQdXDMWi7MrAAm/+4
er4vYhWzGmtpEoVNqOlirRQzIvHwK3uWNsRv4a5+mTpf2NA4JKkA+0W76P+g9y/MVrMzWwhkiwnx
ZyeAJXutx+LvyplLH4MIjL8Mk0mqXvQkR48P5zgcPgxd4AsjzZViJ2SakhYUYQUN6YTFDjd9JhJN
YGRDJ0PDq8Wp80Jz9K/qj0sXDDs18msGtRu2LKEfD10y4u0UYojPb3VzLleQbTy9rRQuhYfoZ/y+
iTPa7dZUxbh73XyN3Jay+oig6xgcJbXNWFEenK1buGjjIHngxWkceCaOGezCvhRedEfrm2U14lKg
jeK6fDhd6gyoUTzl5RH1AuUGTicYe5tWExdg0NBeEDFfGW3Ksqcnr3l2tQz52SxNR0oMe8441ctl
TG2QiYYqH0CjwumHIXMMsgFfA7cczpS6HHfk3Bi3J80CPH6acHXHf2461nKKGh3bK0nkB9bV+w/k
o05/2CBfmO7X5rYsg+kLQ8uCod25OGxAO9Ay+3YJMCsf7pvtJtpK9rNCMoGDnt7EtKFNdjKkN2Wr
krzgBm8PapUgxv7Gkc5/aulYOXJtRoM5DVMXFF9N+RCrmgxbWkwvfme7ojXvDaY75VYn6xiPC25o
7TYuaykCB4nGn23l+tOXo+lDEZ00Fk4mRo6Z8ziKtp30QYpuUjmAfvbeWjJaeb5RW9RipbQ/H6WZ
gsI0bwm91L6GTwtoo3kfxP3gwTZuu6T5zbsWmz739Zt6Xxg8qVy+83ZhgRu1+XDf2sLbtF4vhtxV
sknjUshZr8b3Gl0BOIzf8QrBXXzoPSwxZCuOqYLbxASvM+oxNatSBwXFSbmsF8FSjxQJ3BMDReCY
qbXtbac1+rQzyONPkq1uH+K4E5JWAzSE807WGYB1mFwmULUqrKTLLYLyh0nRZRwq8H0S9ArDe/7S
f71ofFkpxlfXu0XdJMykCf+DYtmgpL7hHh0Cfs4xWwCiD9NAvbh4NqcocBGSHDEPs1+Azl7L+7f8
/qMEW4IwiwKjM1kWK7c8NKoQ2PXL1RyPnY8j8uva/fAfCThss5qwCyjC/d3aQgeymA6YNPTb0Gg7
SHvH8UgcTQoYZC1uFgGRpFVugORH2jilBcV8Hc4Di7VpwGWeH6NAqgT0sj3iE7Z8HbcZvsvJrEk5
bSnASBYF+he4Jn2tIrxwxThA/Lvg+JSTQHy2KMcwC8tZr1ihErq51QaOJpK2nKJAujNrDrhCmurG
F22WSRGp3/gvie8LHiqkvpGa+gji7KamEB/wnMKNzcuJMpSfLB/5ktOM+HCoZcR8GoxtBcatWteF
h3rR6bs5uOqDrkepg36lvOX8J9sEJJXYlk2iqY4XfC1eUSJHRXvP511WScRrnvdBJrNrAwwtcY9j
uYUQ6jML9osC7nNKB5oIKhrbZT4nyYLaQGVenTJAEeW3cXMSBWyoWUsctyzAZ2gdH5O7VcNHHWvZ
9/JVb/rPuIKIWRVylBGSgTF0opR4tAEbTIXoUTWmu4lFWUjaKnPQ+yG43mwzs4Zq8CeuDpDD2BLn
FJy2gXbr+3hrLRJZkB7qKk7U9THdmNSi4rSlryvml5kqPBkibI5o1W/3P/+Fd/Cwx0dB01Ms16bI
Ad6lhDXMS1txkcOww+ATvubz/atXHzFW45bMQSszPzlCPwVSN3b+dZZPAE8+8OsN3kAPPBbW3u0I
s/w0Bu7duzarOrdAEAykpMQ1PBy98C5mReUJFSa9176uThDy0sN0FTsPhMiyc3XTtEyw/fMJaRIl
hMnJAFi+jfnUAfCL/1RFZIYizf1+zq7U5e6Gf7gGGlrbWXR+kfdIy2UeIOPebacHPuZ9K+YTKLP8
VSqSWi5+SmIZqfDHclreLqNcZkUplJ5L7nJPzgG/nA0FPa4gQQh1L7vqVNLv+DacfCjTiVhLF7s0
bVDciAcxuIl64kr5i910TZJuhpGUZG37on1tFr7DcVcvyDfnfvSDvMHDd3Kp3Xs9uVe3yN/BTW+G
I37CKQJwRPB3ZegSjlwJeCgLE2WA0kssrJgQpEp+EzhhxutRgMgyeGOENRAqY1ms3kCHyaWgD/MC
4l9TIef5pSIBhTAKfDp5GoHVFaPE+ah6M9vb2jAmtKzcP6WJUE+iUri2/6rbICjz4VyZwua4T37t
+rJ5Clu/5TOE2wJ6vhL/0cHu9vQVyoFHTBtH6zFZtMhwPr21yf3knQ+qCF+FX4GqELzf0+QDsje2
05Eml+ZwXNZD1fLayPYwL8cLMTNbESPUNcBZaW6We95yI+JWrS46b8G0oUiXiJHe9DGkkx+urHLm
QWRnuwlRNz7b+2NYVdWYKWCC9FneV2RS5W1a3o+KeXqvjgMPnhfWUZaXODSWCoIn4w+Ub8vifTI5
PraJzbP6GhiCSWI1lhPf3QMdll67CXP58dacpVVoxRr1/OQ2afCnt7EerkSTSQJMvSvQ7Zt1sqXt
ZhYdH9mqDf+eKNpJvTtX/4JEHlaqUfNGIg9ogfuodXzY24zkqza6lbrDGp27K3eWJdTJck+a/15M
CYFMEOHdtsxn95Vj0rEMfVEQo3jXL6iF4Lf6qEHTk0kTrD62kukAgm4gx5Mq3+RtMM9pjca1czSr
VaPqQ1bSivgtB1Ay2BwwqRXCCQNy8j4H9vWXgH17uN6jQP83kRLYbKA+PbtwvMqS/0eb0Kc+nPWD
251W/3LXeCZYtwZV6FH5LQ4pdfDKDgiqr1ZByXGNZkZuyKwmP8oAOuZyiSJQPJ82R3fC67msSnI3
N/QE8Lezkb7sTPp8RVUsG+wzAbMSUxIbXK7r4azHQl4Hgx/1tLY9ph4I253ejI7Fw9NmxskFsevD
hntcyNW2GCwMAC+WxjZxmZKn9A/WNkM1NWSxnfFXHIWlvt8foKDPtvXEC/N0vUxiqrShIvxU8+eW
8wsTAntt5lswB++cVbhmKGeS7w3/pI6x9kwC2Uog9yewgdPqXf3AR7WXthyz6wsgMYFLOyi/0QxC
741LdJydnZKDy89r6dxyBvl/rAjg2VbCXMZwWLYuiCNyFNL9i0sNbGHr9s8dzZeXIWJg0ebZeoJt
mdjC43lvI3cXV8MAVQIhBYiP5s7KRF46ILZaJ0pyV4aNOKzpFzvRruQHkCjnOgTlm7+lf7EFCQBl
5w6jhZ+6ddy43Cc0ro6uqONrfo3gjitJlPa+1o0z188Rhs9InGjnH63NKA9tctmnw3iC+k06rQEc
5TpPNGSpmIpY1bi3ZiL9w1646BjN/9b68ctV2hh587MLG5S2ZaaspDA6CugNh4OOHmiqmZg6Vl2c
2nhzfypMt24piQr+gQxVQfhp93KT/OY0VZg7fsLcqtBqBj/aP6VI5YTH9XPhRQ/OPzuqoTkobmgt
amZgg0mSt6UGKL1YBbNc9ei94/fWoUMV6FgH1wOU4342yP4vhCFJ9BHJ2ubG56RMmDnHC39Lg6Ko
NNzKhd11u+F2ckFRMUaWe1aCARgtSKahg4R2rk9UjRYpusXHx0wc0s0AgTszucISh1BdU7eBCqp+
8uCXSjNZALzzK+cZZzpPp7M6CKMyKy35PfyNjJPGpvObLPGk60Ut8iomdo42qKh35yGCjIJUfVcM
LpHMvZ8ZiCmYrEaJrirFK+Qm5Ae/eQjHzK+fBvGsl9o/xtTNWX8Uaf6xKIvzYFuvb2xoGQk4YSBd
xw4x/OlmpemYchylKNPs6hJoqjVUnobh6xQ7ZjKS0TNpd9Yo+0xw6JIfQNR/BEeGEXSWmHSJtouV
0OK1jstSbXTPIlZATnq8z0/UWw67SneRcvZomk0Epj4GsePvTTqjHH27wfmvIoKOHSg40Q5QMIPM
8y98V8SRngVX8L4Y4V6gr2lfNFGXGW7gi0gR02qqzsVuSTsZkCXLnPIuPVXmjh5jje7YsDQ46gfy
dfgIiRF0LIlP8yyQ6e/wkqyPodhiImQYdJDqdoSUvMXEHwyq9ujynGaz+DAFVQ+AYPSUNQEIDS2s
Y8QbjGfRvKRL/oiwvjRG6Caqvydwn4Ffg9IBhYp0mjWv/TPSPUTXWhSi7PZazyA7V2xoD82hvuSm
Cp1dRLMmf7ZXW7fOQfShOhwk8Tr4D/YHOI4sFiCxukZ4XfZStAs7OcWBZZBGvv2C05KhE8tcJ5Gc
gy1Q6T8C7nzcFMdHmMgVDVVGs1PHasHUV09SyjpqO9VGNB4BHX402cXBDFR6dFAzLcM8X7uU3ZFF
qyqQLfSimo3cQf/cN1f99XJ9SWzAk7EfFbaJljwDRE3TNCk/CdekyNFZLhURdIVwGHlr1SNS4eNl
UyqMPU6S3jUrscMVi2bvwk2pR2HiMSaOk0c2t4M6/zCsHwgqAzI6F06lOvP606WUV3D6NVF7Lj8H
a63HN3n+jIjeQkkaCk+wumLrT3c4b7aOmj48OPAgNeyE8UFBzMfhdlDLwUdgi4QktJDkkSP+lHk7
oDNy0ch3MjvmtfovrVqEtDSudAP2IhjPDinrR3mCzAv5gi5YyceQlMjQURGCGYhMV2Lq/keiYH9L
q/Eb+clDf3n+V8zkktFGmYZsqIPUOIKSW+pUlIDzS791LOCwvQpmYttEmCUyvWwJVaS6AY2HZHhl
KrADmCkzvuugpIFp+/FhrHkm4d/5uHBOuTJk5AtDT0INmapjPzPrEP8JxMNr9uu9PuPOq5PfGsvS
oGVfflhVy6ZJAPz/ozLLoTQ+aPGRoX3p7fpfzncC/fzb0ouYZVVKUUXHAyNlPtagOV6Qt8ZtxkfB
rE5+I+on2a0knKgAZpTJTlLMy/UImFXSIgVaaLI+eY6n/HB0Qfjzs6EVimYUKi1TUmBGZnUCPudc
+N6DmThKxdthi/8t4OrNW47cMwbOWA6faPS5SAE5P04019GYpx/o8Xi+TnaQWiBJAdYYWL0g/qn3
dACW5Bj4CSaEiwEUEjkqhKGjcBtLEtrPPjBJwSVILjaaxwg3M+AjIAKyhUWrdr3Cfj0due4tpzrp
DfHDvo7V5XTylPm4SKj5i0G6Lo2kGHMkujupQhRHJRu2D4ws/fVtm8JbijLdSgeeh60iOsi/pWQh
JUejv7303GZlhVvYcAhUDHraz/Sb37C8wuSv0t8fR9YjyYeAgnvNbGM9aFb9vsQrFWD4zExWw7bJ
4WWL13c4hFREdDDZcaU6udS+6AulbCSAsaSoG/zuYHihdFsHYlPuqi5PHZdNaFVgG6FQMrxF/TWK
Agqm9t8zFFYe5nKF9YkwpvXIB666HWcUfMwEh2/VUt5sRizn2QvvHSFHeMSdNMuUjbK7YMWbT1xN
llSy0nPnTTcH4W5HloYSPzHCSnQ27oNXvjW2bkUYxrGw/1Fo3L091mddoi1H0MmYVvPXCvLy6gCW
W5WCRyfsjmbmCz1JaJklfmEQc0imgpZVwnts87cbviOm0nR+Z5mFYxFbGcUVT1tVjGsSv4Rs/cqz
1EsKy0CIvE/6BzKLKGzQPLuHjHPVAokFCsp4keI84EpTKAx0t9lbzxK2v/xoAD1vpMMmyOd7Iwtv
3auGfOrb6e6H68Pn2Ee92W86J7F5ONGhnm1ArF8Ui9bxKg1Xt2lf95YbBQ8uAm2OCVMXxyEWaXpY
Uv5KluNudmUxs5ZpzSXoXQoZ8ws9YJLhkokAUOfiasCyBhIFDym6O0cAO5tWVVsDEyGGAGriQ+gz
VV24JdsQWmaWGYyI2XkdA+ZzGjoJIC9tFx52+ZhVpW4bXXzBonrKl6RruZMnjjrGiw1paeCuvR2h
NXZ4ybP9aU9X95G5RyjKebbs+KZT6eO7FP3vHxxjFDzI3U3feFADQyORhzVSFMBgJH3PQQRG8Tk6
s1J3fdI4bv/Fqa8tH6EltL9wO9Yg0RVgd2LYbaBQEbm3zEJbDMI2vLYG7oLyh5Q/qn35Q3BjDB5R
4F67Uc/ZRZLP2vBApRBALjTIereCOzG6PPjtC8QMq7bT7CDqd3Omqq/9nkVGf2uC9+a7ntB8k9st
EYfxKra3fvheiIWBv6HL5KiLqNRa9WPabucevc2xXEIKTRePDMb25zI0YBS4qADxjwm+C2X68qSR
x8E5oirWkW/7IALfUfKCdpwDgbINL9rriZkeWIYhl/i+OctOKB8L1opSZlNe0OWyeTSYhFclsdew
+m1PqubR7Ab+Y+U3OzZy06q4qXfZP6opl7A2yz2/Fjra1fqVmztMAenpNruJRan3HmQC7qmCVzxD
B/iu0LP9/Mdk3czlAsAHTLy0abRjSTs3V1yfIEqyfGpeuMdimB5/CdrOeeXSLwHZ0gRGuYqsXvpE
hqGUG3RLimXHMM+J7D0bFOmAHTSTHh8wt62OaH1S0ao5iwKygqsxFkiPFLUWFi2KwwNz1uHs4Q9d
irLfzz55ycDuCbOSfy68wd0ffZfM9ZeEJvUZESUenbEjhEB2Z2W3xkVLLbf0naMBr2B4q6+vtjvm
CbuJ19fOqIjWEN725wGNd2LJfRhCwPFSYNV+bXWkOQEzUrDCSSBmj2aN6oG0F1qA3zEHMkAbWFcQ
+eJL+W9KlnwrSYHlENIBGIcHxyXtejCU7yqa+4fmu6hJlhwS8Y0HljCI1B9/EjK/ycSwq7RRkbw2
Pfu1CJf0DdB8Cla4+3L3b7tVFr8ak1FeD32H2ZMOynOHK1X7VG2ElMBytc9twCmb59N6IJ5O6T4M
BMFL/pyBf5+gt9opyUAjbI6rCrWdYSPWaKVhd9vtaJItQ3iMIvkDbWdRyda8uoQIvpQzuozksj/u
/6RiqVUbegzW6o2PRmbYpFuUGPYrLRiEbTD+mE/pjAj04qKuqLiYrkE0FDANnzVFWBCiQn+8jeVE
PPfAlWxLsamOPPE6uLhQ1bW7x6DwleQCAN91kiufblegm8UCocaZFiirbwKmfcphUGVkk3W3GLgO
FpcAR4qwANOmUepZz7nmV4YXIxSOCg+yF8uiSEzwKQtRNS0P9ktK5/a2jdwTVRjNmh5dO++3kM2X
JGszxFLKgWn6ZIvwDsLaSqhyECAI3lCakTkraW0iPCAIsJi3Z6DSv//xyjQtE9MRwsucI7C4q88B
GVuZrY7DHrv8RattJ+N+7BWSuZcoaQtsia6puMMFIBo/8YI2JvI9MADqwcYc0M/RmIe7ernp3ASS
lrH/NhuzKuzD8urlnIwTqguvQ0pkc4C0ixVIq43g5V15K/sL86DAbRaToyIJVvML83MQhf3PM5F5
3EoPkBI9xPfL/6gwknIn2vdgWwI/IjsT1ZcVhP49QDhDtsJ51gF8vDdMR93NoCX/BHSazDuZBRWP
MF471PZP8qgr7vLCpcu++xT//HBhrqVbtLk8vRI/HPd0dPRD4AQTgDaYUzHbLKdqGgxFtWGERm5E
QNdz5vJgfkKBShscY8H2DIcKKSsdpH/zTZaBtCScczcZKnQ25uhPdpFY01BfmtRMt9njC9rTRxXm
m1N5ZqFgKNak8lXjAD5LCwXHQAXmPmM+4cehsub0UOW2/Gn2ByIMGPx1KMoAgz5pTHn8ST56X894
3AnbPPFPg0BzTiVW4OEoTydOpsz8ObImxx1kt855Max7Mk+4oRH0cPIjdvHdlPaU+QAXCeHv/jjW
3rK2UBTaaW17hiBuTfrKS+Vy+llB9gYyBGzA0PhceYesOEIo48X6Wj248XSPFXgEDbV6DgcKbpND
DtCy5BXdTQ3egF68fe0xs+pLwbrZdiA+mKjW5mM+uLALHpkZfW7sHxkhJJkq7pTnjmCyPuK/y7GJ
1KBH+NFKamySlhy849ZnNoQ20zjCyrbbriw2D51/b1dMqx3J6i9880A+GhC9PzoL0JWUg9NSiFj8
mW3AmlELxjQBFoFJXLmdKNDa6sJCPbicsTuwlx9lSC3gEdVLTUMN7uy7iIJs0xZ6SSDLRad0JO6G
qSRGQasKJmPL6buo5eY9n8MqvYHQw8ewf9z5T/ATmYxL/HVDeSfTJw/0etStfMWVjH8t++vRQ1QR
RmKUeTseTyfTEYqTVcobLHRmMaw4Y4yjWQrAY7LpCCVJhuSPiLd5sFyMt0MinxfkpkiprvxETdJW
gsGjvSV1MndosIMo9rxQ2hHXgm99azlWZ/Zn3Ri73bux80islpJgLfAOxjQtcN0iXtyXvyTh4Jaj
ESfDbvqDydOjJgNrFhoSP6DNncfvjGAG3zpH3Kb410pyLUyL/MZPoaX3+h6TuWijQnfF+VEi8b5a
UCNeoDCCqMTu7+VirFAKhdDFbybOAYLKVim6iDmV6auL//RgJOPJT8BI1vbO6DmTbRypewE5BFuG
YzEfX/uB8im3MFK8ON0lvu7JRgdSSdx4T1+tOki89iD+5N9AxKxzT4Rm8/2+jdXtY8cwepTNThAM
AVxFTSb/5vZCE+ucv0ycxMCx5DIA4SWTRnUPPuPp0muGxdrJ9/mnx/4ANq3GqnpHeSMU8kClGCFe
8pcQ/r66NSQpI/r9Q2d+mSv/C51jaG0MB8l3VyGupVZ6F117KpLGjUj4+H27P/4umAg6xfRrh3Ay
BmqwBpHXogNopCkGPJKI9LbwlXPmSa9PeORXeUwvfX2/HPkNq4NOaUd0qbOP2UDc2HHbLDTwW+pP
r31nIWg0+oXKEHsX8T+eenuwTPhov83EXtDDiD001L/p03+3dprfrECZumaq7ERZCFOsA2qoE5HS
VOI9HHayO8mkAB8inSftP/Vz4v/D0Za9wTCiQa+DF1Ep1UTIiG3EC1o+ly+6p1u0IFH9PJto9Klj
XBjqgyaJ/i8AEvMxW2so1f5CvSH6JfWwXj7nk8+zagVuYFys7TP6yR9505hT9ZdaoEPoXrQkTBr3
cxW2oS3v6yyQEZX2mIlHtTfIi1JjavqYBPB6yKbcbLY38qZI0p4u3bzFzi+3kQF3D42bKsaGm9Iq
us2CZLR4yF+8yebjuTZt14/naIOWNumPYeDZG6bf7bkNPHlOSUaw/CfxoRvTrRT9WEnGYhkG/NIa
zQ/AgbWTpfB9I84dqNAqhTkbi5N1FoNo2ic81tT7z5gJ06H8NXl7esF0WQTuTbw9jBnPSMmrtsOH
P+vHn1hd1nyAUiysrsRrl9uhgaAAGkhaYZUypeznZDDhMyQoDBYaVD/U2I3KMQcab4/c6VfvWz+5
mdyzhejR+38pHVxG7ne6v3ry9Kp1TKvMW1hYZVIKs45gCh4S1rsVQUZQDYBydYRl1Db5XhVKhJHe
WA+xpeuWtds6uO0d4NN1y5wrHAV+F+R4tjzKzye0fX786N94aDo+M9OdSwohFuqN0Td3ITUAAA19
UQPoXpyvmuhalb13ZHS96bSuJVwId+59as1AQQtwX+KXhLZQ4lOGxq0ltBGX2nkIr0PKL5BRU1+/
ebSPWApZcxcUCDe7A4NPWKRKQ+kU8uzOdZhkc2Jo/e/N7bm3PbeQ3fYBkG1rGQ6E00mRPyuD4ZMl
9Rw6L6w8ppXr1bY/mOPfG1eHQTB+ES2CasQLhLbT0j2sfU069FeWgMpwxk6iUV6UKKAAEJpCHl18
lReK44vdvgMzcoojrst9UfzoQDNH1D4W03tlaUBs4ODWtzkmam2+GkH4mVxtNUUVOQOFs7Zs1NPh
NX+6cQMzHqYS7nUIVSnG0eq46OX/mSamkmb6XEXN8vJKjzaBx4DmOqrPUYKl5/hBhnz3IT1jWdNo
yTXhC7zxB7ayzMCTfjRdFFa0H9eFvd4tUcSXV71/vrqXGN/ElTpy3dB06P0hH9KnviKoKbJhbZ2x
UNWCczfP4vbZuEOIkx1jLiy7zUeQMY6v9xc3dQY0QmPpLyb3uO3qC7b2Gw4JW26ErjuSkRhE1Xuf
SPje6bKGJc9F5ck0qpg+H10kbVKre/tO+Iq7srjeeljGvwxJzqnYAKFfrSVw4KMtvlhsP9zy+qbr
xFNwKvhThtzp73HnYWwguwv09BrJFsm9a74sJ/8dPF6dJcJRB0pNGbW2yW4X/u6nxxbnA5oJtB+Q
CGC+rVd+Fe5cKrbC3hJOAwAQMwH7V/oRSADlKVefsa2VO50/Pw8kkmNctoua+fTe8L7S6A1jkqVL
5JPCZO/ZCrX/KezFVdfbJNDY4V9aA842WZ4Dy76PcWi72t9R4/5ZnfeSENmP5LyQCHpz0RJvidWU
gFlWW45Gg4VuJ+eQgZcHBLDwx8fkRruZWw8IbTgJ/Tqx+XNwQ0w/RJXcL19BWwlMTZL5lZQa2HQp
J1XX+WHOjeV8H2YB//Sw0LIGzUbqWGaeoZXsbhGtgxPOhbWu6pY5Bvg5D8Jsd4HRb0O9AQF0X5RJ
Kk594oWd4/umdLeAUI/l/lexeJmk7+wOVTs1NLSl/D+WwdE2jjtKRs7+eFX0E0mxNqMerZdJ0KpU
9cPTTUb2XiZqmKusrU6pAgG7VM9L6gLDQewswLOCXRTeNKWDAHSd26YPu5nwZpcLoUzUdSsOG4Fo
uUt0ziEW1CSJ1VR83gDq6uSqtY+0PyUvwbFy9m3vwRJLf0VX0yEJFYSDIuBbr2syGwaSwlCoNhxs
V/0dWWsRgnah0ImutZb+PySKnVXT8WLLVKpdDmszz6F6TGhadsiN5fu6DXGe9QXboX3tPgiTTwH0
3bJIZSdt35EqqQ/egjaFbdNTlmMRCbpY587/hP14odVHnSdhu2tvAvgrUfT995qotbtB03ikD48F
cbSvUhVeruKHtihise5lVng3vyZMRnDfKOv0XI0NFrTwbVP7j5mYDrUfmNz/IJcr++BCySAdnV3D
CaELWYKMIhYcQ7YAki60xrqc0SJ6CLElrIGHw9Nr20AHLw9qgQr/6cZa1JCwu4Yut/4Z+HHNOLfb
n8EjLQ89ERe6NDPd99BttcnBtROa28o6UARd6aAVQzDx5yuxMBVM7p0K1aSvvlLfdGOapogIzfQj
fDNEkEnzhDujd2wKB1oOeQTENfi2rLfv2uL4aOmQprnlyZt6wEtmZ6jVCCq3CB9VjeMqDhSSiOMv
yuUq28PxvgQ0Y/88UVC6UIHXFxr7LMmyx/kh8c2X3K/cGL17JgWJLpX0hpk2HNwQACJnJzi3HXgd
zMzujWa66ap7kkIHcaXn5xO3rmHEDBKijMnjXOeHFHtRTMNyyla+Qf7XgYQNl7oVA3iKBrxpHlde
yFN7P8kwV1lR54IuMYlhG1JPFkdRciNDZuOEQS4OMWQNHBKd1sDeHMplCLQeab0Jgv2Jdx2EADS6
/4ddEiWm6t+EJf2YuhtVcNUE09ttr/HiQowV8EbD0GyhH1RHT4Tv591CkNxcjEeN5ToimIAmGwMw
YJhMwYoylMbRKiSL73/Y60QjvwS8jtYov+lmlC4+d56CYCeKJWmBhSqq6tKounKSFQDO7VJJE4lk
RfSlPdjRHfpH9/nfYrCQPyq6YMG4bZssXKDLyRf0t9fJtXC6s54halqHV3EIJ2b3OkIpSgY2P8CZ
XgjmcM4DLHsRyumFkmQ2td/9/bYaN07nnhimfGDEqW9jqqB1sJJjgtm540kjkiK3qOMtZl962pF2
A+lPpko8EdG7Dc/38XdrpjN841zB/vMEpAEY8XbV5vrLFx1KOZSxGaMmLzKs3zaDnB10ltuRZRLz
U7UBtuBk4UZ1nLAe3/jxCXIU8zzr2cmxfAFxkM5P4HCsCPPTS2GrbmY/zCcSRD2qGhhsogiSOOQ5
m/r1uYTigj3oX+igjfRtRPTWNuLnoyDqolbE/pY+IGfgkcGhVJd4AtX4EEQAJFbX/oim52CZ7uKf
92tRGrIPn5OGkjf77lNiXtWsdO+7qn4Dky6KhuIc6Ba6vcPimKeu6Rv7m4dLCY3v5ZmzA5gF9YeG
WCnHCnfGYPGGTXlkBhUnSYNVSEU+M3MChzTwfpXd55tHVaSiRIdRaV4sUboJSRUODqxwDt9mIi0w
dMbOETlu80Lnytvvkyi82lBQMDbmCkPpUMX2JcBIBpT7GpEtpDTr+ncMG97h/sXQ0JQFhVmvsJsx
tSBZ67Ib2GAqeSVdpXal+tIA9jDLbElFNIfYJ76sAE6yNMfuITDFw5ZPFjnOMoEhE7Aq5Mqc8YGz
jtixTaNLWovCJbjtDRC/pATg8Ue9kZPkN5hIwigNfv0jB026CV5OkgYvj8zQqAzb9xl6chPEGllH
1GnjU0GLSGeeWxaLHfmEs+eGw0/RDCp+INjmq037r10DLbPWyoMdklp3qqZ0HzmiK+X6A2JF87gn
wAuchWdLxVTePyKOYFedyymD1cMvgSUd3bv5f8GJDlTaYPCqTvDq6c0Evm/OgIkqVhc5niJ+Kmgl
Q6kfd1nipEUXw4AS35KcvNCTLd29NkgKK0E3Eb/ozlZEU22FQWw1CSYfsr4eG4llJVQ+1exC4ZDu
FtGSNFsOs4j5HeWCdGMUdcmQamVNRM+BDy7hNH35VblOHAERLi8gxnI9a4r+OxJ8hCxQrM/C8JNk
XS7I3ABFt/r/lM+qyZGKtY2hLQr7InDYgjhqDwXMKZsoCFi9WAwFhQl6z+OE9eE5RhfHziho7jZR
GQ/R6q6ZPcRoAvhR52gW+LnG7MtHKbCsasQ5RnZ0MbwsJ8zGaGdBDNVSBV90PXOwXWI5w46+mCJa
2U7WQMQJ8MoXp2BF04VXAqn4bqcbkcUZ/uWOpJ0GD/p/pvMCrb+T3jCKJBR/L7RsPuentR1dqjWX
C+gSDkw2VGIMsGAGsf5B8zEBl8YOfY9IAP4Wejn9BTK4oayiShJ2ZM0EfsXxBTtEEqAAnNRmjQJi
u7JN0UAxffVZoJz6JiX3q1i7dejWIALZkUiY9n5pvbQ9G41DLoaz+hLvzS94OsrEawYguB9xRAwQ
erlgcUeVDGzQVvjtZi9KcCVa6CUXnRhBG4zPI0id1uhFVP1bGOSosXrayOpSsHrPX5Ohrf7ux5FD
nquAPaHqXXENitudayWUt2qhWOkDGFsYWT3YouBuWilsvK2NbnGkRtU9D2RVCn0igCBkUicD61et
Nz4YrHSMr6fQoCvVf2pI/dutluGV7pztiExFGx9+XIdYQu9G6uDFLsH0GABmmYfXs4mmsrAaOzQ/
YFCwNySGYgt61A1vm3VcwMzNNq/cgnAJ45qhgdRYE1lxjrlp0t/39zya+2B9AtjH8tOXH+vY73hS
l3S6sBJ6KhtVp/2Yz4SzS4ADynboGEP2IJpJwYJafY/YiEP4XiG90X58STt2nfWAq0+OTpoDHF8N
tDgye5QWHIAzQlfpG4La05F3gPdWOxKw5uq/TKb/XDg+kM5wg3PbkMKn3bF4T3QiJSC1QfgOG9zB
WjGhBoK/r42G5mKnFyZ7+P0v+w3+OdDg+LJzQz4Z+qOrJVnTcvStjEwvDjgeD5qRWnmw8ehh3UCt
Gm0FK1Ks7sC9rOmoxUC2IYKQ1rdBcyHqwwbPK2WI/RIaXF3iaD45wuRGerRWKzJUWV8R+58b6+qf
/emoOCZkiID9OtQHjfiPbB8je60aGyuUCR5wGNMcP/bum7v9xEvH5TZMC3VH5mHwWuYFkloVcTBt
7WSm43/nKB5k3Wf/e/XgAluLvGkOzUtco9NJ1/GH9KOfRZ63+Xv1f6I+nelwYZ5v12X/Qzec5CjO
IC0f/AUbGI4gceWSmUP3tfITFjWQVjKxoMnxI1dbCae2s91o21hWqWxrd34jx1ApCR3fxZbuTuFD
qtvHUZCkFySkh1JIDggBrqNrBDUmQ9zR90Wh6gCok62COGzOWBaG6a7JdczuzCZ0rXn5dzPpd4nV
S9qemF4qKzbblwjTRxVW5j3QJCYSLXfncz7YTIpo3HilKz0/NL1z/vZkDTIigCnXsVbF19mdT9Qi
n0LtemUlG26Z+CdcEgI0p2yxk6BBn1fi6hnSStRctr+dpOnY/O8kOv+8dmRMHVzTecdzkITVSldg
Ehf0FlMG5opy0yB7mQp/fUBJ0Nm71u1iMKA0rLrpcDI2bq5KKrqNNA8c/mSPCkqPS+1Da2dfz9G+
4q4H0JLVz5Fxwkisj6k0X87/ctklfXewFAGcamanqzerL0A0KwogNb+7FRgjZS4Fn2O6sj7GilmG
hMUR2vwkFLparEpOiAgQo/aiITTPSp3cZJ4KZ6n5cLxusRtWRicn1y9omcFVkQuRruHb+4oPyxCl
kIwRBkhG/q07AJtNYo4UU9Gdm1uC3CjbvnxGct21wy8lwLEbeO9Ch/PopTqyyH1cS1onheqB9o3Z
SSkfWf+nVmS0dOZU3eTEk5ImLKhm7LGW2Bx0qQ/4Ng0dmdxfdLMtClBR3BRHS0W5im7Nwgi9rK19
u0hulilFMaRNoKh9xhL/CVWWDeWIfTamtzSqByfQ9Wwb0qG1bbYRf9/T8sW4FHIcye/ryW6/qfa4
f+ovvyuUl7sS4SkipztcU4CynwtPb+K1Tsnhuf4A8WY9hrHYgbUlO/fBMHQzN3RnQuZNIQmcunmp
dAKmHRGq1BLetBVzDT44DrbzzSEuhQndY9u4qbo9e5/Qr+epa9WivCPMhZMXWfTca2nX774vyUSk
FL+hBKCulJQRRgosEZ1W7568HTLt/wA3t4Wluh+kjE3HvYKw81F5TTOnDOqjONx3F3x6HM4DXVsz
aso/cGmP389+Cq9fQxKr+ei1z1oQfCTvkx6oYclwrOv7uXCixHW0ehTLKHFO9Xl2Ow9GKUj5bPIJ
I/4iC5Z55SX9/m7HA2B/Py5qvrTDjduNN1cm7rrv6k6cGAOm4BYigHMGOpO6p5d/5H5Gek6InNB8
MUeYy4r/qaVfQTw3D4YNIGfSNOdkpMzzW8Rl8nq6inma3bdeg5R8k6TUcFtik+MKmMLxtafPEe0V
Ps8yCv+ndi41rhMTkKyNRICLMKsHF7C/OTkNKB/fRIu9DEM56yv3vLWihI+XmiQdhAd1vP/17pzo
mLECHO/iUItIK5V3/Am+g8RYWMCHvjkfYyCUk6kZwWTbfF/E4qa9d32CqoCefoCD3H9hLmqfVTBZ
z4EQbbwZmHo5gTN17QZCnSQFagTEXSC9S1bZLKu0itp9j7YEqfP/qz8iwB3LvG/hQDNaL88l+nTV
zANuz2UTLfd5eLSbmGbxgTyDOlFoPdf8iMrJpddcNrbHGcfUdYv01Hn1WJt4JfFFYDX6K/1k/8HP
MP0XX26zVlRtBVD5ZteXV+GUmnTiUkoi/8udrxl8vsyaPdn+cM8u7GDDM5xCPIvubCaY9nvq5aX+
1XSlRIjUXk6d1Jr50L2S2dHOgdGti5e1eLyFXXXr3gFXBe5qLtrafMg6IsHImjDoo8yJPfCYNP8O
bhONyiQo9igh1I2TPnpFjxHrKxRvU2ek/3zkJB+vuWmX1b33GJ7G+QSJswFAkWeQPUCo1U0ae1xq
yWND2KMDrkdYtS0s/24hbpQm1EOzIjZTmkY1ciedjogGxRpBI4NpKtvPZXL1kSPem8ay2Dt1yc6S
A8/HIzM626KDUmCPoJO8SpikoFVGuQl8vqfLAKXu3RWeBe85NiEC2bD6q6M2zqqqJMHMLpi9GQQe
sskFstfDS7J8FHUM7lSo+PKsddRC2rJyrTAhiC9RFkTVNY7VjE+NoJ36xCvh0lYsPO95tpCTVuCb
r6RMWOWJt2pOIZswIW7ZWe55uJp3nE55kPaL3QeUDhwE7oZPkxpAVvEyEd8PhoJQuzEFBBmY8D8v
v5t6rDzrkYoO+Q0e/a5APP4jIrqKoAHCV7elnYjzFPnM01CulZ83udI1i5fr8FE6I7VaKTrm8QoH
XojMuShaQHAVmuKFeDQsERc17MmxUD7vlrd7zqDWaiUcBe/REAIgXuM0SzWEuny4XqG22UIdYEwx
L/z4BY1vSxr8G7gbATRAfNg4nNrL0S5OKOJYyedxRzL0jYhO6zCMsf7/lYjzEjTBMmIoar8+4j8O
ZGrcnSxsai12qjprtVHqoyHFI2w9O0OTlZY3BiVp42MO9ybUMzB0J4MLyUtc76C7qMYaFJBmIr+x
l9YyL349+HgM2Wabg+emWOB4VlRhVUU3ldG1FlfsGGR6WNJ7DcWrCVV0GLGfS5FUSeQKQoF3+boG
y47KmMk1utOIeAc9J0SN9o1yQEX102NW1fC7jFPVWqjQpC7O3Rj1mixfoHPQFekqjEKXaj4Qswzp
Q4RhtLZZudIv4rW8Olm6SDY2MBIOdrxBpGlKQdHwr2+lLdtBt8ABdtg4cv2hCcNN0l6d6yCLvVgb
JOI1qMyBQBRQ7e370XirxcSkh0ROAkoZ47bqskDqUwUfTuvqcl6wIMGMg35C0X0Os56DMDuC1NE0
7wOSfznVHSyRE3tRJktEdVCPwmaTIvuqCSgZu/C85XwSasU0ptuDzuQZkjK94+2L+XxFf0IoXcOR
RQMNFJjvQhvb4WIbsBvira2BH2zoAkvOfaSMgCGAgi5/uHOmnslQL1Efm02clQaNY+ejQQ0ls4Yd
/ZStId/4qgayhpmCxnSl2pqTwBNnaryIltYBdAgiUJqyDsH/UumnwlGuOAGWjtrNdiRUnZ5kxOXd
cXt1it4lI4cL1vWkiYwusF3jYGlzb+RIi8NzNL1FZyCdnv6pZbYhpv/2jfxCLZ3F09wBlmAWpWib
2kNwKcoe751/y7Xq87xSoFHBaRJBM4W2ymt1myx04PUCSUsPxz8Cbse6olgyImlqbLp/QuAaQRQA
DyTcTe6E6soYnfAjG2fD0z7JQH8Jcn3QGb/x0zNGJ7iy/giw8898LHu0rkQ4UWpCit7seBWIc0l0
4/TQcMmVVvZ7w0GDRn38cG/ZUHNv2zPGMASePS0uaJNGKZO0+5c4L/ciXSKuouIKwBU0xc4bCHtV
9ha2jxHQ4JgZnCVOOlAG0Cp/fFaZO3/T2HfZRfq/z/D5Cy2hOkY3j4CiqyyjSvOSYAIJqoDS/yHL
QziTW9mTXqZQiHFPQWG0Guy9RPXaGxlGBIKSOihxMXEcjDZ3X5ZtQ3aOWhEBo4X7iD3/jjEYiGWc
4Qa48mdrEQHJovkmwn1INdtWtPC25fQPMIJ5yNfIoYtpi1qHkU8lzc1hVUh7zsK124hod5/N0TMV
782r4ItBQz2OisY1PnWnnPCsUeyek6wbI4yhsppYpWv9Cg0c2bjdfN26yi1ImTAYnt7GjhA89GUU
f9NxcRthIgprfcyVsEafqH5XRKWmWx1sL5G1YppYOilKfu+FZD0PQUHUsDBZ2bSTuSxz1aPFb4pt
N+8LlARULsMsDuq6yoQQtj7ctG/BIDSEw8M6KhZ/5UXh4oYg9O++jwo4dUOv3sjiDJH+21Q0/BD6
uskr8PRyQhj1D4A8CSdjNMusDd79yA9jyH9GebRfpolv9BFQRMggJNEDNHPPPPpAq2WBgB/xH9N1
Mku1skB6jExHNrLK1RlBQRGAXAZafdxy/r9ILWxiC/lz+hQjgQ90qFwbKccDqsOUabGTayCflee0
1b6y2obFJmBsM0so9YSt2OcGDJAf4XHidR0zhZimBOrKeb6nfobjtStydRAydTln9egghv3XqePN
9cXWgrpyHYI0B6CJHFLkQZjuB0s1uyDY5YPtGSpxFuat1uE0fMfFtGKEj+UrSacTDZf6Jsh6s7y2
2QYioRrla2v/URfVZKVLaiqX5jjqTOAGbx7Job4eijefH5PQVhV23XyMVBUJSn7cSp9PxUoByoBP
lgvaAqAGGeqZw1lilCF6fO+NagDvBeW1hMhq/jGF7qz5g0BdRqbMArBs28Tovuv/9c+jCxFWl0B0
y15KwCi5VN1b9Ni2Qbz6xXnxAYNbV+ZRmtkdPRyeglDrKdjJ5b2iG438QOo5KMHbCqSFtCpPmJ9I
8dbtPOuE6rRtdWFnFfrIE2wLWeG1GXnbh7vJH/tKiZxq7EvKQ6HLK6+yB3iMpPvpmVzOKDISmhxX
jgKVoxs/17HID4Ud9Cp1xGg5pt+tExC7XXFlgQfKyezAnRVO57ImTc+lav9uZzzXjiJW9CVcuNM2
rhgTiSp4iXmfdSfrLywzI9XlLFY8mTz/uZvXcmz4kv+l4fe1gwWiK+YUP53analR/yuvCRCj2wOW
x8IqtZM2QL3CdoZrBn3LJIEQ37fDk9SSUWF7fIXgYPcOJ7a08GSKAIHIvadeBkSSDKYkSTCxITg7
9GhZULL36MWnIAk6lnSWqU3A5BHILHIiDihkhZKZl9KMrJi9qE34+H8q34S+IoJjJoCZCy3VNInv
amDXA2YMhuN02k9B3ESWLGvV15ng2ZM3Hh9KJnSPj2Dj835WhUW9A+CIqq08k07TLpMs0JU6+LSa
waoRWmxjqHl9AgOm4zqjqkxAW85Pcww2gH641c+DtjKEv2DKML9zpXLQtuPI6wtSa7vgdCczgYWR
k1CqFdytXVadyt5uiu4G+4jOFi57lXENP9WK1Gj5+7EOvJ4vDvIbE09AAlCOSytZwFN5a2wb2gTJ
OB68irNIefvUCa7jbqCuKerZIZzNKfKJpOMhgmqljyEIh3CEhRhBKX6JObilrvvAWcoz8TwEoZMA
DRAKnXCHqCRvwLFQoIFjx34kTQvlFRhVJlbwVGnUvLvnqHz5RpnIw+6Tno6bDEF2XYxWvBzkLhdK
P6vAMFvjxPrq5mM1LjD8EUNzzNjCtyRk+roGia3u4QZjEJSEHeI2ilVZTuBptDe/X7etR/m0LFsa
FqAb+390rT5I8bZ8GgiU2wmzL+hk76vi73ozZSFnXQ7HdFhV7BHWxPW0No9pRue2EcDfdC2EIXzu
4Trk40ck59MZxW/cUVhE5wqFjTrNC9k+Mjbx4R227RaSmhiBYHUl9mLqpdZVO5JCnwP57dTzkRu2
spFYJLboA1wBlWor0j5emA6jOXn19CnHy1ehl4XDXbRvMfGAyqqGd7s+4QUXd1++ppHLmaZxrkaK
ygxh6BSu0r767PbQ6Fl/aiBhf73mYLw5+nW/LA4aEoy6fREsZDXbrbOn01bZMv6JJz7TtwlnbjLF
opBm9hMmlHo2okPMn8UWdbX5H/wZLw9eCGNhvzETbISRyR2LXFspKl3pZpDyUpSW9yZF4ybYUSTu
ko6JRv2qqu+TDoGlTdJwQqzGTqlYzBKTtyLIVDxN1svRzSEnAYvEqXiJGyjMzM4Rscz2kPnBg/iO
wSusL6vLFnU1/ziwoj+as1S7IeQV0JGRC77b1rQD4PT2Gfo2zxwH1We2QbPTg0ibkNjqXV/B6AWp
RIbaSuN1vzyy0umbz+2V0K0XM+aY3zCNhJH1pKp5AGjH0Hk7BUgpPUJ6EXVG30FB11LVycBkH3uA
3gaJerB3qPWxJU3YfNcfGWaWdcrFC6bDyOYRpjJd9t3Vdffj9eOgQsxEezAbR4+39a+Z64vMeoof
PX7Glq2086gjMMne3K/vt2reyng8Exz3hs7MZfrqjYUXrPjmhHOgdFx40ywSHcXzYrQNGwiLNycz
a8VaqjrkiPeijjY8PDfbsqH6FojxGkwnqkSb02qg3+1W9VXrT6H/LatpMlqOm6y20m1eX3LLE4hM
PPaHUsXyNCehSionxv+p2bdBicI4KVE1e2dZgE/8XuaXlDwr0IZvRWF1L4hJzTx11vJxkeL8NtQu
rbbmpXq1dvpNHZpoL4vOeS3DbD0OXK/sQSzRPCSJiA9TcAc/w5N0mVooFXI/0OiU8ousVjiitvBV
xjvjsjZFjr+8vtmt9fArUlvkAqxnVQyCaJ2QOW4k8xZkbMaKKigsZ6YGGQB9Z4HX8o0BZNzNpzWc
SuAF5Tnxro8GIVWyi4LeON9n83o65j2brSi9M5Z7JWSDTuxoRoslwovDNiDxppuGjTi3AcLVJYTb
RrblyFamKvnOhT+V5UKpxwr6KqMoDqiAR1PV04oZOGW/njFvxpXjuCYXKDmnL2qYrvXji6qfiEbR
txBiZzytt3MRVWNouD4MPUo6dhxrjARKOfmBVXQWa+3zkM/9S/71zFgfCsozYjm/+cXbyYn9cOQJ
LfNHfo4Z53fKxaFAthHv3j7T2RjwnifIo9J3QfKhmc4k8VXcKmJZ350MsGtq3Y3hWznOFzrRaHc6
+i6fkTe9pYz6mqo9HlREeRUMgb4+Lfts+K12NEU7kNlsrfOf97NbFQYxf5HiKlcfJ+fnM5ym5TFS
10IPBRHNhj8pKxLfWPNPSXa2G51rmDd0GdxE7/PeIGioshwhcWmkh3TMIZoEaRLlI/5LWUvm3VLV
IacPomNR0jGFw2qpAF1ZCZX7ge2A4JzCWggIj8EapxQsYHoJtNdoDQPka8xGzZxMjI4lj/VL9Ljt
2fRAnWbRJFFf7deQUnPfdIMgUisH2FXYHwpd/+8XIOxriUusT08aFvQw0H2JxpMG6VQ8Kqn69pX7
niIyXPtluaLrgocuhvAjYcQLKhjYpt0q0u8jwKJ61C0s4FYyOKdDhvgw7m1Ahp+I13ye3IFnSP/w
8osT2r5XWa+jzEgg9GXJuLAJC/butEfYGGI2jalqeNLh/oC3S4vJ6FIrz8WyrQqhtbVYkGOMh05a
+Rbtvmr+B2/+VwLHMcFQmSpwtrgVQa7OAF3wdNTkhKG9paQ167Uo9NKaFJKfgz+n4+3JEd9PtP0i
c54FJCpahGWI149IdUo9clSi7RATVCF4ILJr4x8m4S0/3H1tFTj1hVST6sfe5zAyYR6Qg+dfZWWq
MyYcurLJBDQm+7XPJ9g/7J867bHJP63ORm2OeWpXKRG+IhywMD1Bm/6xx/qsC7l0lO3fmqHg0mKt
9+tIp1+6M8loIPNJfgtr6hpr/bnPSUw5hzlwPBxaKiLzd4O+eM0NowFKO+Q9PFxFk8UA/myghPrY
+Fr6ZU3YMP599q/kqHiBexrv8C/TVh8YYro8g7EseUeKatgFIYUTU5NytMHLsW1pK0IlJeIPZ+za
/upUuA1VuzM2bjFe3ey/n3d3ah2DUtRz0UFJqhirQr/IuaC79sO6mdZhkH5lfwI36bRA17YMX8Q2
oGRRL04B3LAgZfyrwXHrA4S51VyJ2MZ6e0bDvuB+g12Vp7S+FGyuW4BSzY7VHK1ks/eET3DY+DfU
skzCIsd9z+J8dmtyzbpXM4LQTTXrRCG441BKmy0SRvXjS2r2n8RuJHwybsMBiRCmRO2NaoZkmMFt
nruxL/B0wq+VcRpMPGHEOHcHcFVr1XFspFRlAcua2OfB4c6kt2sePO5koKZvGv5o5kxv1wazKydf
/79518hiqNf56nKoCOChk+gkdo0iQVaywYMU4ZXenuNlYbxN31MPegcUAJIdTNX1eMCNfmTOgYVJ
/lXKs3s4QuJ/hMe0YhdIt+ovRTklwD71LOYdFT9fO+9oKuzt+y+je2u41fDeGN7SIm1CQDbhh76N
Ss9VJcNM7q2LNxXzJPZ66mo2kFUXaUHU9WLlW19dUPSQGm4+cUApzB4rpQQgl/SjS+83A48iuDkD
Ijz+pEoa9Ymo7hrlKhUJ+vO51KJ+S4MxrQ9gdlmRxNg2xjxSfw1y5IazE2zPLSgJVDal2YQneZ+6
KT/2qkY8/rOSSs4b61c+rGbWYQkqLoZK7tG7Fhwt4JQYOFAsMKipzhuE+E3xQ8JPTNZRcx0rF7Ou
wsLCSeJjELdweN9Cu3p1qd/d8Gf8de3sIn5ZHiTVVP0rp0qH2mbRmOScJziBppSV2tM5ylJNsfd5
nDJ9SetEX5OMyRZr9vKBkssgcXEd/cZP0fnHB5D7TKQy7BKzabsRR0DwH4iEY7jhz7bvkEW+JKWA
kYquapSst5maW2Q7ofOXhOnXdklWxXOrgNjLnJYSqMFxjGPz+LXT1KZpOL9qiY1s+DWPRPgZz3Gj
4SwZ6x/4yriyutEVgUjIeixGOtG8VPttSL1bVZ4ho3+fRkK5C92P+PcpKKbzJPqJtaBb76hZvO2o
xbvSDyWIj3BxJ2x+4LWFHkvH/2QdHtHrVKSC2wL8NAEdxkAyB/ZJ07QiBpXr3PnxYna25qnYhSbb
uJCHqmOAEiirNBcUV5VwuoZjI1SZi/xXVtfVgIHSUFygD5VbUIclX0tbpFrojQ/7lTYUs4A8dusH
8DeKW2uhZdoNqh/tR/EKvRLGZiqtcdn7qLMBJkUioJRs3DHSNzbHIQaTRmM5kTyBnBy4LJNvCvBc
ZzjOgVrlDw6Pq/vtq+56xQKreQIg8V9RTtFrT+ZoP1QYdhJAkQKjXbQgrNpyYaRcwzzbd/yh3Kzl
qILEHUy8ClmR2WCU4ChowAZBGpGKqeui0ztQ3nsew3PxfXmEqIJVKClmyDkVFWb7XmiGSnL/JSLi
gN8QY2j7KgxbjZ5vmRyFTQwXwqBD7H654rItjYFf4AbfQ5PjfZJsnOEGzWd4MIaltB4Yer8aAiax
B7E+liRRPyBWTBzDDPICf+IHc/B+4EB1GsHQH53k/x4dimrwX3hvoTTpCXfPKzyT4La1bQjIaPrk
HDFY9wVffDot6bsCxDkyGCMCNQbM28ULssfTcVLkmcZvBUnlgmaPO/d3n2EHrTHOGthy4DvrDBvE
dhYJ5jGKb5pffS01lVDsi6mxI3jh/w/bEUkbi2uT78z6517wrsKQAxDYN8QYJN0oz8Gzw/2c1F4e
8F062dT5HcBe/OZcWhC+CIp5bu6okowoNe0ZnNC/sOpBXwAyB6yWddbNJ0ku7rofdZgZqe0Ge1CE
8VeA2xBCljNixrt7tfrFs168ERWZgw/StWJC6Zp6B27/cZzm9sA7IMEJNmSv7TKN33o4GYZGxgb0
Ep++tCjBgM+hFYWZdA+RgLvxX/vUT3/zM/8R5xdq3SYAbVom5nxitSc3goiqNx5vBM/4OgaIy4O3
NE1oNqsdD4hGonsNnJdcyAyNInAratmmZ2VFc/WTqxWHNjwE8YNxgRQp7wKgvgIEyFfIHvZv1+HN
dd2i3YKlJHLqZ12mImGrnRPsCuwoSDUjsSfJ9sRHmZVV9HyIzZlVPi9znMJQXain1XydIUnHQpu4
YVZMiYY1OhIVQ1ddJdEsSF79R/gS5wz2t8+PEout9I7N+/dDpnRxiXhuXxpnE9gE3mUNwwK3scfa
BoAw1+KmAGGgXElmb+YxJZ2PvcUBPWDioDdc8wuDueQ+M2KtYMryOj+2z6WqQvknlhvc7u7Sw5J9
WeoKMezu2PoEYfSIX3dRPNlUr8edlml0My3LLZ/mAfBmLnpo0kgft2RHG8sOjRA8YGrGEK8u4adR
97lxWbaGquD4XXZxaVdczzN/u7suZwexkyhwep0/aZFIJ2I3ICzKXloMJFdQrklIOZRYtxlyzODg
1X9UEjP/j66yiRmyM7ilRBFia2mNJFrGqtl2JYcAc1uYaSqpUKu95E4F81/kyNjT+cPIUYX+WNW4
2JR27DaurbCSF75n/lBzzFtOb0D/sifOi/IqOeDTnd/8OTdmZaO+Uio2tzKT7A7nOR1mW7ndc40F
Pg18gpQ+LiFTYjGjWTp90T6+NaGkT9SJPBfjK5TA2Z38GcH5t0Zmi0t+/7YN91evoy04OZOph9r0
hVKLe98yVDKyu56p3/j2hBJpcXVOQyfKhVrPireisjO7gJzj1QqkdYgMqCyH4nHTqQApNXuCgw4c
Utcis7XfplXMpr0bXcVC7HR0yVBEl0dJBFGUXKr+GYkDNi5FS2xb5pf2aH1XL00ZYvUD5qjgDfeJ
rM9R8MYseCvhw0BTjUmNFwPRdgC3+Qrs5P9So98DMhr4sg5/ZxNJmj8wKuMae6gEI5nUK9ojnzX9
CXTlh8BgH2SbmN0KZnD8YLoJi520RyZPOhIe5426CjvtOQWG05Sm0nzuDQHEZOrgbP/YYkFxmZJo
mYzSNqHnjQVsT02CH0cmgjfOGGsz7hqZTLY3a/JY05sQlbaIlpw3zj/FIIkhjz54mB2k+i1lkGuy
lVpz2dLZN9eL5B8aVAMmoKk8mHegPQVr+3qeQInaf/ifCzCI6WNK1QoFH5gsmChl+9sBTaqLJgE8
LGL7ps/7Nc70AqygtomMUtrM/gnffG0PnHDT/0op+RFQvFKp8agfJ5RcEfweEAmTKFgEJojkzi7Q
XoPb+fMXKb6o9jvyCgSo4gotJToNDXoqhZAjzuUefePXk9eaFNjPYaPFyCKmBSYKJ92Fj1G5MxSB
c5YSTgeAEQbpBPGZuqcV6CbOFzK2PMlVY4hEeyIWy9U0t+keFmkcL1L9OoQWardH9eCxZU6ampR4
eoVZuyn6YcbW6EuqlwsAXe23dOOjEzx6k553CTCRLmiSHgjUuIjiXx21/xZ9LPKdlLop3OWTTVh5
7UTelGdOg8Uy07jD+yGF7zfY9PSmKNnlCoAADESdKIkISHbjE/9XHi4R2WaLXoqJPtQSh02xtd+y
UYVyrD5kndv1h2Rhyb5fZu6pVckqVFYCAfNSSXqPq+Z0aJs9b7rw+cNNU2DkB8ecfRec7zYOxHhn
ikwIgQcLX40X8YXyX8YoZikyhx+hoaWh7TB+0iyw+d+1LJ5PhCkFPki9jzJnPR2YOx+miOekq6KQ
zbM1ejrE8k7WGuExziqMnqmOxyfjIRb/UopdskSeAPSXtAiwm/0szi0AxDn0lFeSKnhL5pWiJpk3
MC7h6O+taOO1CsAWFdCtMiL8PRnG2LsmNXv02IihPWGbeoCiPRzKWyE8IWWqxguNL44KizJ4U7Jm
GVQHUkqith+INew2PzmqYSJQXrwoH3Oru2AV53klZ0ILEZihbJXnsj2Bi7wQtH0r4n1nP7pIweCy
K6zgrMW+Ewu2b2T9BAmT3FZjZmrOAdEfKVIsNuGti66l2YEzHYDwy1tVx+WWGBQI8GW/0W2ttxi9
k8P2EWwmrJEbFXoKzAefXt/WHpU7QHTBPO+pk2rm5f8b3VRe/GYZJHI8+KvdP2aenIZpvoK2pABG
1K2vXBObqIb5BgOYi1abJD8tLRvN7lVT66ARo8eZJNCAvpyaZ5CiZb1ok/GN2GLpqz+HeeRgFxYs
qg9Tqt2i1Uh60Q4x0HnNyrFW6SWP6ezFYu9PSm3RmN+Zn8lncR2Erdql9UawZfNBJcKt/fwbYBzZ
tl23/KF8+CYcjbrGpE5FmR6xE6Qo9tCtFp9flh4G4p+LKsI0wVEmy3O4FY+8RK46Zjf5xi82sRzA
k89KFlZbGMCOovDRvO0rE0LLNNzA9eCxHEGJ5Zfs/7vWRUmleK1aDfKjPSIM/v/PMAVeEf9yOegV
chtdH9zjqw7/APe9Ot50ClDTSxjwiAIl3IUVt+r4zbZDsSBe+opwO2PSCmBexNXMVKLuBkHzJSKV
k6bBg85543OuclSZS3PBryFCM+iFiGqU/ND/es9noHjXYtetYvZ05c+yiChfnGMXzi3REl6jSlmf
SsK4Hao0hsyf2YKwlMhHn295adP2TbNLh0EwV7+fpNYhfC0kWFn0HwCT9E1EQ8Es3SeS/CRaLEun
xDp3lNi5FULOwWcI1iwLScmtUmsWTkUw2AO93XiQ8/tzHE4xRcKar5MZyuUZuFn4VuGk6wOs/zsr
gG3Tko4xjF555oqPDmKXkrXMP6LRZbOiM3pTsWHy233gLbIdwpk3tjBns6x7GIxuz3If2NAHiSMi
/iQjPoBRrl5IWfo1+vAhAAA1H3bS6yYFfHZKdgPgqsFu+ahOgzZJftRHBM35WuhJyVAo966UU5Uu
PrxdgvufktdE0T7nItOGk0jEuSusMBj7GavOmyy2YwoPdW2FU5d4Mz8uw7qe+MbEztluM5HSA94K
9x4hId04HVykEPxEcJuKDN1TWo+0Rx+X8xukBOErUfKNAyKhFwJzyI22mq1gDuUgWV7xQxPmXQzq
TFLmswD3/l80WDJVRdx3qNE1sSdd1HeAqk8IK17q5BDAis3P5Nb6474o03oWlbpH35YRe7a5Hkn4
SzPgRkTauoMnB6385WMDO+WFyYWMg36Gr5lxOYuUYWcpjK35V4m9f1olsA7sIodStUgWqj6PfGwJ
BW8R9fo74ZuFIVLsJh9wdMs0B9fT0ERKd30KdjzyD2NM2pULoCfAMZoT1Wb6klRoHi3qnKpjOQi6
fnovYDcimqfuO16MUSdmMNshK64uy3/VwAN7Hsxs3HD/dlBQ/ToRZACoG/N2SOIwOlVV46IMgsfS
GCx4YZaq6X2ODLJzLhWxmONBO4WU4S9SyK+4ydNrOHIbMroFn7u9vz7CsH4TZMWPlT9RevBHCrAC
K1Dalkm4BriE2bejc8VNFu+bjbgO0XgA8aKsfZ7bAEPGGzb/g6f9t8IAT104lxvbFkS8wKSvg2j+
jjZgZgnabcPPT3GbQ1Oi2NIwHzggsPS2nXbXTTsF2+zVRYXXsIbvajPGMMdbhMbKILYLBLTpmI+S
6p6BJgalPPe6eq7xcpk7lg3AcjoEJklW0troVvkQoS7KNuTuMMhbFC9mA60NUoSEqC5UhdscDLYY
pr/3ZAhToCYWa060fuA6PpFV0yBSrxhFIHuV4KqvloK3weoCUH3D2cAoASmFrTaK2jVwD+5tI8si
MYwlHfOYDJh2vMb0R/T9Qx0DOzF89KGluYlzrUeMzCoCPzYaXcOnmeGZBSBDm/y0HSFHQoTT0wrH
68ipJo3ERI5xEdD6Vr9xJWZ/50SDTttHYTUzvhFw1sMt41+MjHepJ6YSTt3PdE5QxsPfStrieNRZ
VG5phdpkivt0UZOEWuBXO95GIzeLp/g+nmNTUgAUTzVHyPCxx8jbPZojD408mHuka6xPE779vA2j
vFAheEJh53eSkqZJziGG4dluq2ikmdq94am2cKya4/FoXF+Lrv+nAIp3h9oyngRmPCzkpPx7JzZT
quCOrFJnpTSk6t4tZCuYAR10P+lQkOuEsph2XvDqpbA/jixWzJbS/Fpb0Ce7hDOX+aTm5EX5/myp
Vu8HIAHgqQtWWuoq1lZfFqfXpaC80aNzLLTnh1VPVGof9z04iaBAgkkAvOYc/PdQ+3XmyfRltlWc
kQ9XIIt+ROX3cEBOkTKoJoCuP5Q4m1HFfm/ezpVZYPhYiSVnzjiAysLLQgTR3S8r9FMiV4vqLZJ2
I0CEFFFNPOZJvaaXZE56qmOeJ+UNIRyaNKKgLgaCvBFfwsp0b3L05P+T8WuJvcVJ4yj0HN+HTfDy
BCs3rVJt/6iRDf6BldoaFnlWNlx7owtp3XRQNw93xrslaf/wWsT93lSs4aAWiUhcbqwZZZhgJgAf
QdTBfwocNfyFUTLS8dWNncgGR99D0aVmhDeD97URVtiYJwHBQpnAmthJiTX2a2SKtY3/r1Usj1LC
X4E0ZuNqSW8LNK3Crjsm/trMKxX9aeHOfUajzlEzPEIKNcH/NLqBjhMy3VeiNHSAd/M3muIIc1LM
NeFKMnUr7Fpbkfo3AbC3lyx0+07OZMhVrsFmai0mx8/C5f4NEQdv2SHaNhvDriBcY6y9MJBuGIXM
7jwUqeTsziTue5OcF8IhserwiX6A6T9nQljW+AlPhQcMTxALATrBL2VQbgJbd0m+vTjtb2ni2vMC
u8ddIkex5CxRyyvdm4dxdcu9+6tEH8ZBvE+NeIXQEtePXZGur5rx8pZe8yaMxIFynvxrxqA7MxhQ
lWPXO+MO3ISxlbdyRHLrQ71nSmfGn5fMT9jlM3IZY9KVgX3MOOxgtsQBwGbsLB+pW30hRi9mfxKi
5E8PeVYR3Tp91wnEOqPwur8XMIplQfmjJt96SKWUDsvhlaWg5hXmNivGcdQPW7/bKKFTSUbNNU62
qPyLT9z11iCoRqEHIcOqo7sNKOZDFRf801wtE+HtbV7QsgdlvE+Vk3J+dJsPG4rARAgMtOF7Gby7
SEDHLsaOiAc5HrbUCTeAyAWV+Dlhnr+IzX5RCDjWC7MXWRv40PkJWAMv/rvugOcdEV0uEEEVoOu9
ae8lhx10NDxxJI1Qo1j6sCU+iSWtYhFPpd6xZIQe5pgO9Lt4SFWGk/9xnyI91FcljA38MfJenTRN
2APUrCknmsLV2aO94K59EFzB9QpgCy1fP2cN8OUPqqdHqc9kMTlYS7ByzRfYJk0ANoSAiu3Labwd
oYpjGy6sLj6wOmJ5Wy0nEp6tOIqmaei/WRz7i/McPfW0xiJRjE9fz5apGI023iOab3uotCPVkG8r
8T+rjkPcF0CdoQg4ErZAzOp+dOc2dk+5amfUrrzeSrAtV4e3thOpRBPDT/mNfu8bss3zDb8V3wLF
MgZXi0yj7rzkq7gUTjzOdwhRK2q2EHtg+GPY3OWEUaQObJX1dF7aSU2xDVjbUit8Zs6m1s2Du0ms
ofDdRhU8x2+QImcqCTgAokLwtmSp9X6t+qMEkkK1uMKpENKtRUW+aiMjfqmGerSpVokDe0r5Ph5s
jp4Ak2bZlnY8zvl2UffYve8/rzRBw3OaeTtaJMKfHNAqfDWWWGxPSjdAdQ7LspdgRw+UnKFfGx2A
1+j3uGDoFSMx005LZrx/nf956htfe5q5KUwgGtIwHBU2oAgXSbD8CtWpgSzKZQTbK7dctN9eeeth
+d44o5PEu8FRZK0hq8n/BAXv1aFS6YbPbaOBh0MqRpqpPTWDSa1vsdpJKo0STliMqpWedj4K7yAv
32h2VsfsdSuxtVFFdyw1En6kmvcPAIsjRE3kFPvX/dy8wIDeTCt4tpTOnLgdRb/ws8FSN0/nv5MN
2nuBeufKGP+LVhBUOvYKubIvT6usc9Cr1zMeJPHfYYsWxf0/90zZjZslkFVKttlidTEgZ7ReKxUC
WSinSiBO7Cdhglt7F67KL/P4Wxeg2vqiMFGORAF60bEDLiYrHdWy5R55pm06K0g08869Fhf1Ga1h
KopFUeTKQF/1X5m1PAsOevbOwsynWFnaQXNxM8k8nZn4YCeffsPt6WRPardmBDOZ0mBwpi7z+qCo
+k1Qa01mXc/JpvVIv77WSkJQFlan5wgNpy4nDVsIRI9AF2zfc4EEgrLmMxfAuwD4hJyc4NJWrbpa
AAJZVTz/q258jKcK4U/PTi1nIJeDPlhBKVUo2hgXCOH37dyyQWs0KQdG3ABZMX9ywqlOW87HD43r
w1e0cdju1rwRuu2rNdod1NkRwWSm4VaGqlBVpgRhMxBdiJVTspgfl0QCZC91nt3t7LSkrYcqxI3o
mrsqxc2b9pqh+b+Y+NsNYKYbNv58HUqaGfQ8HYic07U/eG95KVxd5rHLBtMBzTcoBxRPQSU6b//a
l6xZgBLlgl+2MrhTtSlJ7U60W0DHe3vFYBSNud4JGi9XqoBUNk/sR3IRuZjalpAKNC6Trv5nHdsG
DEi/GSxtsNAekik8NFzYUra4iMhwZXnvim2iWpYiO8tInDfxvBS76LGJGxwyGx8aVBEoHgWr97HU
NRjIrQLSNRWxSrGbuRwWTlgchTaMXDmaVPAmbetQfx1/JEZ7l3OawpYj3Zb4Ie7/0fMs1BQFQZ2a
yiSpdUh7VCKi+xA2XWmFr5ThYSQ9zs0ECOi/yCurDVR0/KhIBXNOwlCsIdRAf+LX/+beUaaDhlkx
GLmblQ4Op3q+3p4J8iVz+hgUqiNgpd4KCZG8/NiYkgo7FOHBnzYkF+/x1Lli4RhzXuy7EO8pm/x3
DY8sxUa+qr7pANyDS+T9dsn12tQVgh/yLQQe4eSOiZ027BL/KRaE2zvCJWrNSWsRX949v6tIK0Mq
W9y6EHulSns5/WODadnBq1arxQTf2GSZJqgop7tUOWGQyyHyhJLGj0UvU9MjbpcbymguGoW/8t7s
AxHnL2o+CiDM1KoanXWHy/R75FKG6loFYRSpnEvJvJUnDDr7NCIoDCB9aUhF/UUFRA3nZ4eQvTnl
NsACE82zLiT7oRRskvAI2mNF4EtPwcRGIR5qhh22mgC2/yj482P04/Fm2o3+nDsVQnd/AkVt73sB
qlD0u/o//h0A4Cgj6p2DONKVKMczFrOPRoBL9mZdLfkSrpbmvkTcFAj7qvGWk+VSNcXeQ+OGLDd8
4snAUJDo3qleN8xOPtPkhYsT4YmLnL4NSAYWbmfs7w3J+hSoSCdAkp+heVr4zA9yuFJuArLr2gIT
Zyj/mZj0sLTcKHvdje1RsMNmXfs9vpQGAyGZl2rI0XYcdaCwpTGr0az/GQnYPHIYRLnpRdgeDyQj
GVeSR8XFAEmF4t8GlL/O+5pxD1E5v2ShupmIF3sudCMiB2hncBi+81w3G9dRLZjMidxWKetwYMrb
36A9oejH+7+wqjy4G3Qog+biPlxObSm6ozvXFHTPnVDabDZAUTayHzP6mtjwmc4qTMT3GB8h19PW
SSZhoAQz3oo22/RVMvGorIIYwW53zS8shqZj40x+lgXVXDx9GrxPRMdIpTX5nHc6UJsN/cPFdjgB
A/Kxw/ulRGJmghtSCuN72AGnrR0z0ZWnCPEdv234NyFX5div1qa9yn4pAcN8AEUGZ7Fiktcb1jBk
XxfhRjAxWn2I6EqScnSH7ClkD5VLrmSirqkopRgYu9ZVv+OWcrQfziP1UjwN6QViAtnGDdrKfK9+
M3BIYarLL6TzSkg8CFDdDgApOvzotLDJC6WlNJrIfa7RB/bL6ZYbScds5KFgRTPiGAycAERUqe9y
6ex6h8h4BR0aXWPy8gBIhbDF32XoMwTTgHn243+IRMgw+T+GjpiALizPfPtU8oTx5m/606A5rLFi
CXtTDVFrffY/AKCVugGQYiQo2t/oqbPyjeHGC0lfJ5boJ2qWTb9EUci3svDwb4AN5UIyNHBSgBx8
AuepbDzzZZbl2UJlb396g9SVdWE+ZawXbmaneqE/YH7nqhN2vHfDTaz+eMIjqMPqSy8KETRUP3M9
q4MJghPwVCuoPcvgZJFC6b4u8BjaPaV6inMj+jM5cC2AFWcRjE5Cd/N04zxLObAdcOuooT3DYKAU
WBrTqjJjT4ca5G7Hc3XF6An2v0IVk027X+3XSRnTLMs8HEafVEkaCnAmmjweSRzdeYqZEQP/cr8p
uEAjurJvWmyL/mWh1GNYCrowuzahiY8RUx+NJn7hSgfexutSNCm4vOHtm6mdJ2bLUY8DXwzi2vhN
1MNkxMnmrlO9SbCRSVR0sBOxayAsYHoZFc/bqgOfG51UNfVb0Dpj29Fz9vzVvO5cmTzUFLJ5Cw14
ECsQlqLYCK8qrqUpOwwCDPAdGXRjmZtaqSgMa3THez87816WX4r+nU/9W8ZIKKRQVrcJyrjE6lr9
q4kP2mhKzhxZVWVV6OV1xuzhpvHvGBrROxDKQVNI+q3Fcw1LxmVuLEpOJpm7Bg2G5LlTQpz+VLp3
KQGmx8jwU1Gr4hGp3qQ5arOKz5aQXZ/wpQIMukL+dOf87AzMHkwLe5XN7EWgP5IQE8Sv64lE+Vbj
oL89bOuBr4l0RQcWsWvbz1UQ3QDoWTfVKbp8Q8s+fS5DS+1GASM1R5+KBF/PIsgzIPXx+uVEyOSZ
pr/AG9Df985+txdxogoVpmQFyq9XU41kY29GMqVneiJkeSK5miy5AGjBuZf0E5hrlqeUtKYFoZGJ
y5kJTb/5lpZFUwFf+sFrF6soIg0pVraaRLVxsVgjQPQdRfRzJ8HHh5untsyBq5rTUWIxX/TZ75bH
bCcf+vYQSYbb0OIUKhM3TDaDUSjcbNTBjwJQ8pk5eMwtQut1vab23cWU9m7uAtNdK5aP80g6+Kv1
buRq4Bu1j9AxsnyjE7akzWm7AF4tCaqa+EBcNA1qgN9c2yypsRwo6mquzHb/KQXGAVy0jfZTAlvd
6AnlkPcoJFBPmGMCFvbO5arz9tjDA+gLZs/02oCrc3CjgwxxD3J50kDIKp0KnVOeVNuJGRZefYAe
ohZ+LtvgBhVhqmk3Jnv+J6KWqYWZPt0bYIM2ru+m1f2crP0mwmTj4m+dJGTv3/5LclEMvq/4C39v
mu1d1CaqP/uNsCWRNDcT1qV8AR0C1S1g2elv3GckyW9vfBMjPDjkDs7KMHGX8cNS1ci9RKvoJ28X
0290I+BxI8i4d+Z16wgQbHD//YCXuw1VlEdGlE80bXGsEXrYwpnYhgEJOmyqXkcJ0Xi3G7TNY437
Q2dGpeIqMBNs0+nUihQ61l5tXTwK81W/sSOa/2/MJAsLacw3UVPlCOs2yas81c31ksGNMUEJ510e
JbDprYFYOt7xIYPAwEkMqXogupT9tf+gHbdMxUSELEJ83sGvj8MqSlcUGOT3eDRF+Wcdwibe4wIs
WbQxl3+EEfi6ON7MDcyMsh0gsUooaJSrPaPeIWQmJem4SfWeG16QXnW2NvgjTrEhuP9x6crPRuW8
3BXdyVaY9npw23fDGE2YH7pjr96HWddFQP7D5rxA6XcB7RmRPyNa5Yo3+y9YEHlpq+PzDlUHnxQ0
3GXH4jqqIKrJ0QtTxn7Cw+a2pF7KYtTUVTkkU7uvZK7KuQowRQ5pG7UP+XcTLSsuOQ2G7Npw9+Jw
kVI0fwq2CY73GWSanRKxw2QZD8NUcPJ0V0kY7JBZjnH1tmn2idzVOqvnVGduWLYwxesDycf0JuXN
sxHLPwj3/Km0Has0zvvwa3/DgxqqYpel9LRDxA6/f+99fpJE52AKfns+Adyz3MCwVzRddC3LcVmW
oaDjqOdvo7Mc9+dkhXQCf9KMz8k7GHJuQ2Ql/waSAxXgGxM/8ZjOpuNR5kSj26TBLSOlQp69VdAw
S1TSdT7oZkcHcS0eeZDHQ4Rvquw3zcHAm1pbMD672i+wFyIu5YY/ZRacZ3WwHnjoYiH3Tmvo31wx
/487KqcFcbAI1ljB7lN8BUygoemvs1DhYC+4JVllwJiR+wgD2RaWQj+nlzhF5PswgMrED5LvVMi9
GPgwbNIZrOfX7laC3bpreSkBo8RB0ZrGDjsCt46paxFRocX+eiz28nETpWdp377QtQ3MCjnIJTP5
tOXYuFqETjdPikD+rq60nhbjte0jOOwS3RaS8pHz+y3Ba368xdQoC2wlCY+bVg4YCw5gENuAd86e
apAW2F9IWi4D39ag+wqmdJ+9ZV7zMc3FzkT/Xn//vmXwmTYOFuZKq55AZq0xhVwIN4KYeZk7I/GX
m0wbCkxg7L/R3LuRResvp04N4We37KjP/vhHaOLnonfh/aUFuWLvYWAT8HG9BJJq/ItBKA83XFlg
bPRbRTRujncjJgCbBylCRu6G8Mwo0N28ZkKQstsRcRuSWbP02X+zRh/uRh+3vRUjnvEU8qGLDoAV
l5q+663YI5sLiCWjdNVNJ/Hly+NjrDs251wVhlIhdqGZK9jNXJ06h0zfUQuKPpZiEFSfC4nH6xoJ
zqIYYQeqwx7gvNxg3Kwr6B+kxC+XStgbzdszVsWcvb6N33L/Navhi1zuquQXzgwuuJzccDFTypMC
7UN3z1pieR+W2jQkNJl9IMbfvC32nKald+fFugunZ89bYnZDxixwfLmLiC02Wm2qFuuzIrn6Hnuk
/9e/6cvOfe3UnEf8eE86iWmd08IHlsHBsu5leB3Z+MZuyTJOY9UpF8vnu0euhiIiYf3Dk64tbgVE
daB5MvKeoiN146DqUPxkkEGZbm7j32jLaAA2qixoitpGRD9UQBY4c/z2+KmrFAai4MyH3M4xm72e
AQDx0VIfibMiyrsV43R+QtBQqT1jbT26W+9Vlhs2tV4feolClrJAYf3ccliFVm4KEPEaHsrfZKe2
q2EXpeKaop1ddesSoYGTdsWkZgpCaKV9DVGPWhDoJpXzQIkBXOnHMYiBrdpjs86j8fLanRy6A8oX
D+NfQye5kgecPgZU8qEm1BH32njj06Y5h+BMHFgr1TyeKSNta/yFCGF5/9O83lUJAEaLGXxJA7jd
HsI8Nk+HWVJzJyrdaVLdbthEPEFbscJ7Bf7fkbq1/ZRS4o9oRZMm3I4IfLhjLSnGT9Naxa6bYF20
Qt7O9tF9NAByIID9eff8IxwaCdcPGukqX7dm/5d8uHMCb2cCbCSPOzZJ//WmtPxB8HWVzOXZF9JP
pH4WV1JUh07bjJ4s25f2h+ZCml9Lat/oNwcsRobJaRqh2lvexH2sN9cSeO5zciIi1Pps1S1bb0X+
lXlYRNv0l90rtAI5cJVCLZqJJxGAbeZRt6Enm4vXfCuVjaYR6ZEv7DWbvqxuDi/flEiMHNH827pQ
Nm6eQFF/9/LvDoixSM+STFvav5b8A0R1mf9Qpx8AW2rLR5+cw41zb5bw8LJ2gw6rKHWOYysvBDqd
vRUbyHlwpXEcaXIUjZVA9I9luUHtosY3WTNOdhhXpfpTxu5X+/+E7VUQsRribnERPAZy4KCT889/
fbpYPcepnAgQrjs/MHvlUOt/LT5RAwSoEWGaBgr1I5FiIXByX/tdZdkrLgmO74d8AwKXDy0O+GFW
2TtfBXcQy7frIjkLIR4TUUYZQ+Pfmimjtv3LZWl96GL2GGMpqrIDWbZMK9DDnzJ5anT6mG/gA8Dg
5lVpgIr9evrQq9J1Qq4sdM44EGkDOPFt6W9rRrS8sn3/qD1J5Dd2fAGFWz6VAnTWcFAMpS0ioCjW
UUP3oLRRFHOdMTPv/g+6/uOPjoxQeEyRa/cxc5DWblFVjTdknGu+YPAELqOe/Av621KDUtpt3xx7
2xSWCjO3s5Yan/6lgFyE7y0PVUG9AGr7GZHyvVZTWgVuweg9EU2Va7AToKicGsbFoh1SEYpAVzrr
VbRTiLpNGF5vwzTYttDbmbFZkbjkJJNG0QwNhs/hRW53hRCN+u1jviQiOJ+0SyP41muTmWVBzoLc
ZDXyMJTSvsgIVAyJyys3Uka+HLwYy5LEZ/oM8JK+2l9u/jHQh3Mk6Db791S2mJvkb6hloWryVK4L
yAfzQ8Q+mWo6hNIa+ETQUqR5U2GmBbIhZBxtjoPu0TFampAwBmXs8+Q6vXDDiOd5kMMd37ZkZSpi
LZWi5fX4OP2ezc9pmmPcjh2i4JdjkWQjpw7OfGY/GIcDtPvbdvgPmHVGYNTxmt6+nbvOz8jCYaAL
U+IHlzHAMDCnyJ/SX0m4DrvsSrm3DCKokMDgGHBx8EHSTxk20LZUtYgnREjzne03W7vXollV3TDY
BvcfYZPbBrLoo/PrPSYoPTYU2RzrqL17Uor9itjys0Ciu1zVMQvHRwzpo9fB8XC7oxlpqjZ9df6q
DoHMKQGCL4avFrQYtjgtv8/4vwNZnl3LiVa4+3XCWX0aOytoaayXkUXfkNx5CXJN0lBL6DiDasOb
mQMRO0hkNs7Ose1wFd/X3v/PTsjI7pJ/gfkujWRRnPz/VtFXymcZjtgGYYVJp/jbMREk2NxA2vh5
9zOhhEJ4VBx0I+TaIlFqt+n48jUTX1w+YJJbJMorgAJwl7b1alm4TcVMrRp/xZmSi7RqH3Wh1rY7
R9W+b7HqEiUN/K/QkN5Km+7JEKFrtYcrTvOMDnrAjuGgfAvGApn5MNpb8p8bb4UYRF+RXMA7qH+j
qWwAfSzR62nhO7VffTWIsf9I+1uEG2y6pN8OfL+C3chovkf9/qHokbchEhQZ+QVd1Di1DGmLX0/u
5wWomi6Tju7ARr+KSw4oSqlUixOYyGb2PsI/2/b0SgQev+12vUhSuQugeqzA+EnkXAnvH2IjO7W1
RUweirZZdHL37ZnorzNti4/abqPMj8F+bM0xaXLm11MKF13a7PdZgMjJsN3yyQoAnCOv7fdRAhta
wg70X9PBplfXxgBntMT6WmEJxQd1hAMDI1YUxorGeVPlPYNV+BiNkBZmVqWdfWAkFTQOXS3nwdqK
/4NHCW03AneQxhna2RmbGi60KXcr4bcwRvZFbiCxfS+kexcwBgMOPqnXGfTGtLSfCsgT8CnLMTum
u6aMc4Rz7T6Vxrvv6/NRSZO/yF693QI/QCjaSomJZTmbkmsJ7G3c6c020ElVspoIt1KiIoi6KDnE
Y5xEwM1n5A3fM9ua4dOU1Ags55aZvtJpb+nOTGjgPakyETendoDhmpVXf6O0grMPb0de3XBpOtjZ
6eW2lI0pkj4IGFLd8QHJ59f7g/K/q10HftkeCnxTubA2PudA8FWDlvZy74bSJh+DI2F3/+ShxLcA
H2jeFT3SCPVVhGA8kYXnRCXZYjh4Q3XgRETbFd8vBKRmTCmktYB5+tz/wbCP90UpXkc77irUVIoP
S3dlVF4EA1FLt7v42GnTWpDcst0pKNsGJz21kEUww11bu1KsZT9xgWSARFOjyuOxxwA1aHskwYJM
GV6ZrGX31mh9tAa2xobvVNVTslZmj7wOQ+Yhsi6U1M22w+59xZ+bvBknwOg0zE5w5cOO4GvPuqDG
Vt6kTsQXiaxDmdu+PFVQbQgStz8RioAcPNVokoZG8bXlAT9D9f8awn/Q+j3eu+vyHkEsSYWKm2RC
O1BUzbtcC44GCFVg2HEPB2SslGMXlZ/cRgqcuaZMWAOfEPKgXwJNGIGWJWmSaroIa71/p59YPpZs
r7o9tCvpt0CmlUaVdQ2BcxR1crG+Reu8JTHRBDrh5gRjsTc6zNpAK0pHambLkXpTTgIGV3SaK8tC
3yIqii8YlW8F/U7dySdCXi6mcAh6D8Sa+9IRgHTHB6UeaUCuQFJp3W2vkdWCyGN3kTIwuHza9vy/
uwCEShnADFzu+s907b4IX1EwTfciTzRV4ecCelFHQ12OTDMft9MegUJaXwGcUtUeH3yu0TzJk+QQ
h84G1qKBTFxCOxlyNN/OlF8+I+uztKVjvZVJZPZSj9jDXwv4HQSZbWUESsgqHGcKSsYQX1+MwWTh
wr9OaVUObH87z9vhSosbO1VlL0Fq27aAv7RBz+rk57KU3DPEAa2X2SjD2mO8jHhKx63xdVLh8qgR
h2msTTUjugou5kBQQBql+3ev3atGv5nYvr/8TSFcacgMPpjkI3BCvhn/P8yxotv3bEA7EyPb+QqO
j8y+l4/JfyioXRP0m8Kp/wn29+FNk7ahWDB946mqojKFHJGojKS+Prp9NbheX1es0YEG8VEoIVM/
DdIzvRPWzq1AEDrixS7+0RqLRAuf0xB1c7GhkY8V/nGXABSwGKjjBT2umTr9XZCnPxcKjbPq9Jfj
WBRPsDCLiqU05497fz/X4Hpt6T+9pdpVLC/hzKELxym7XdZnplKT1bOi1AITu4adh5xSItu2SRTS
6VQZWAP+NjPmt2wfaRXLG+/VL0XTSbA7Iu42skoQgeUcqs15ITS3Njdtx0AZXiPMxncbCwJXr5QX
YMugQKncSSrU9d5q6UX8a6kibqjhoVNB1cj59FOqUtNcboyaoSaUmKU1YZw5c6O0dKKOudD3iXAN
V7FVBSOXDMnzWRTGu6jHicdD7jyzTnHynw3lRMN8NMzARUr/KTqfz++jrEOqDGdQI3tvis4noRMN
m6b6bgpXrjbU9RS8zrWRNl2qQUW33eaCz02WkSDI+gnbGaKM9c8v2jFtmxbFpkR/HWF+s34gRdpD
pPEKJvrsA16J6EJ3+ZsWkmLFtFRIO6Yc2kVSC9AHSk8OOib91w0XIZbvMXINI0a/JJTRkXL93I6H
g/EuAGtIJgG3R5JBALrPddM6hN0Cg4PVpxP2u+TOfy91FIl9GYtOU3rdMbuajCGY6SrNnXRBwelO
t3YsxoNZ/YwXlgMSta/jGHnytclNfnb6NoI2FCkx2Xob11N10WmTcwaE6EH6QHJGH+RtlSRXcFm6
AbGK16MdRd6kdD3ZO54JmvgyJ+R6ZOohVvfv/HjfhrVPsiJncN7eImsSxYzh7BjK3d1cvonLy3I0
ieJ0f3u1hTRsAJ+7d4XU5nryZTHHJsAqmvyfXF/PiEmTkf7ZbkLQ4APZKJ9qlIXAGp1Pf+3fYKc5
R3CEiUBwadkbFya6CaCXAFKu6DJVHKHT52jqZFZKwlGey9qqYIocHKySBys5k3SRgVVznyBWRfL7
TQvpar+hAAWdnXg5R64kXjCIU40toZoDtuI8qlwj1IBoA2VJlmAmDGZ87iJ518QoWs1xdVl+ONWj
nM6DXswcDjN+91GhoJ2h8KF++HcLpHy56/CXz7ZFiXE5Zgl0jKa64zlVpmhroNGwzIxXptpCJY7D
rUOg0Xs2+PpqLv6TnczLu9Q8cIub5bFkQXJNGPDd+ZsYq4mPYBjg+iGKyD/u9BnBCseVJC9q9squ
Pn3v5yPG6Qu5c9ANcZepKdVP1QhgNlwBviRxn0uwwEIgwlUh/0Nlrlwbe7+YD0RvkEnk+RQtcUWt
nWTciaEKysLcPh0SUPpM5N01Az97dbNI9XDWc4IURMrlTulHcQ1WkooPM1Ehg2kqQ6UuzEOJLzsN
B/00XFKxr6dft0FI+9SqBg5kepLpDUiUM5bqH9nP2enV+MlQ0ieS4GBNtplDNgWV+66zv1GYMejn
3+9I6nfqwYHMN72CmaIV9aOqn7ZBshXa3P6gMJlj0jkxNAch679nRFZXAez2j7JgycEfrLZ5ZqMT
dFA8p1TbVbqwI8OK9rXkMJ+dM5/m9xOno0mQc9YXTovhNXClJ8MYLZhJUgLoF/y+E6AWtHMaLnRa
meDLO5xlMptoGmPOL2mny+G0J+yL8lf7DU2gKDEWEfW3E3yEGWnXOWrmdzjUerXfTGhn8Kb59c8c
oexAkg2zwcAmUy1AJq4aRHCx8ITkda0LqHqrFOzvtu00LFt2qFdHCBePU/snyofJ6QR+pVqaCM14
c0pgdTPl2DqAYOhPiG2pVA5f7ttY5g2Zp2eo1wgVfV28gRhK4jGDy8Vu5A0id4EL2NXBzBOApfHi
Q7Pp0s4eWI/0M5wHzj20AsUpTY7JvfEkiv05+anHe1gWbJ+n/Qcj829of+tHBRTokei2IdAk2ust
yM0pnqzLUwM6V6lYwpb+7uhVNUMAdE+lMVy+SkIy546HVLimLlOG0S8EcukYtQF8qKbPujDJos/d
7iGed1mK1uL6SCvBZaj7s2HLU6y8z8N6AwHECPTsGAowYGT8Mi2AtvjzbAfSdIwwHSqQTxeQBFIa
rnzyLAYHGJ9K0Qxy/n/0zxWrtSgodRrZwunZO28h5w6McQfU9jzyNbmChvVrVF0QPybW9fScEYa1
ywdIN3HjzApSxMyx+2ZZ6IPkISEXNEH2Y/BjxVPANgk0pd5f8QUw0ZwUr557y4jgZz7rMswRDlDO
mcC2ZRXbmTsuP1uhBo/V9uL6CZwvI2OvAnBLL9vQPRMdxqYm0Yq3C/IMxoRrM18YONOyWbMVV772
R8ZnYFSWdeRL0rrh570jbVG3zDaMdwl8MQkEMlhFNk3jR3nD6DnAO4weIvgOrcoVMmPaFuYP+br3
NtNwrTGExFL3DL+/zdfEPxvDEV/Ozg4B5r81NVHyt2uVdAnuyEh1RlvMfH4+PX/etLe8Sy0HbymT
y5C2fYCB6nP6S7HLCejyRNiybsGF5c8cLcMd9KAwjy2PkyG1Vi4yQlMgq2frzI9pRYMdxYVp+Fhw
BJMqR72AvqnvSXTxL5MdR1A6npDjx3ufUqhx8UCtWE27H+BIpi50AijiGoNkeZpz/E31yEm6PypQ
FKzJzco3Qdl+fNRwjR+c6Rp2eDYETtxByQeumzvb/LajUlITtTgm1IKv+R1eKJFUe0GIeJQedF+p
191yI+h3GuKn7o/JqbzhdwDr4PCU7An7l+HZtURgaRhowFjr9ogQsp6dlfSlH0HKLyUDuQ9pHuuL
aji+w8s4mSdjbIJw1gj5OppYeOcIwH72IFpIAkeFGCNia86IsVs6NS6WyzprL+mM3GsjbwbTBVTE
jE/Ua9epnk5ags0KquElkhpuZ5fyimZY/E4Yjdd40jDdb+/k1x+OPoKxe+SIjm9+jTvKbvb4+4TS
DOrTNhd0x0WmFkTNQMSue1U+c4MS2cGBWzoebddAarrqcch7UGNDV6M2ivLx5gJzf4biHthKE6Dk
vb9l2OFZsVbpqsDSDoEKnwMK6Oe7mVLqSmkRugRGp9tUSH++2cTkfDMzgQO1ndQg9xCUHn6FNvqf
wE7NX9SMd4O8rnk8K7/b2Hdk/SqvWruyAJFZMofMPgXXsUmWLimz8o2Y99lIQmh9eZac3ZHBXJzn
bcfvlSX7TC2FGIaeiLGhENm2Vynr0usWHy2TnsQpOiCbb76Qk7/yvZTahZrQ8DFOFlX7IE3crbT2
lQBnWuc7cjpoIJrXrdf6zAb7FWY9hwRA41Py7tVwNuKeSm/uNqnoqKwmAcI7Km76rk5KZXSGNoUZ
svADgTv6aGOVgVvSYO6hM5bMJf1nUUF/YYpYBgkb3lzMJ64QDDISWS4IgEzi4Moyy7sAeywTwxll
0CzWZyF6qiGPdBLal3dAWMR/PLVHya8aeEQlau4TtVleCs+DIlS2VSX6VFtwYjmYa9Bsv0S2Vo/z
j/aTQnyvCO1iqj8VvrjP5/6cXpuQkZwA+i1+6hU5YGLaunTvuH6dlFr3U1BPfHmWhHx+tlHJ+xqI
v6sVbcFz1iNB8mIDe+qKr+ow765xraEW5PHDATXg0vNpGoRdG1D24XIqXVkauqsgyt9I65YCCUr0
rwxbP1GOuJgTTDJA0huRihbh0MnGIpaOAqCF2rLYUjjbcSw8egdHzF+a5eqcZ66r61NQLNwOsLzk
KjiVRz0JEndPwC+WAZYa2CrjJPj7XNHGQkg9bXMccRGOjpIWE46QDVOnXfsBGW/iJibavyiHmGf5
0imDsWAjMOz18Dj9N5vTEYyVTyk1wb3kBwY9II812V5k0/qgiuW/5ZX48MhO6YCoapJynuIz92a9
qxz1FitRbMYwtz55h/oUZdpr65uliCFacSkRB6rLj0JmxBABewBaM5wRT5u84k0DU8jgSKlaYiZz
wsqQp70jqZKbIlPK4H2QQLU5sBbDjEaX2OxTy/GA/I6zZUgEASsD3k5x4KloqaGHtYQSExRYNlRw
uLqgyotsq/OVHPhIkLl1rFOkFkJipx2vjlxmjj8DmBn1Oz1ou+Y8PEMKuncM32HsFIode7Jxujim
hRDu5ujrX9YTfgrE6xk4lHf1FRZcgKpZC0ViVJa4pcbph7vqprRflM3ole5EcPeZpVLuhP+4191q
IAsw9ZVm6AC/DWtyxxd/ADeDtoPDpUOprHnFosrWwq0LJfSM0evrk50CtkzqNzIP98/7XAc5KAws
KQIX1+7cL7gSYBJL+HxN0NEEPEHhPGlseh2XcmHgwqJWwaeryjQxpuIhYeKTx/LsgH7EJsriFcxa
n1K9g1dSNBbV3hR4uVTZHM+D9haABszs1Cf+WlwoB2SjL8vfIx5+YUwFux0oUv6ao+ZhdsbiY96R
yctOBlBrhNOqUqcPXzr8D1RVF7ELngy7Nsol/9dhqMuraZQT0kDOnl0XDkey1/OnTLYhdApFiMMr
t3ZhzR2h/zqDiGjflXzuw2ObyNfeE7Fjmr5NC4wo5GG2m9LPXpA1eclJnJo9HucBD9K02VJ+AT73
rLWm97GRhiTe5dLkvzKl2KybsKpcUZ8gBGHe3kSuK6O+6f1Q1W/42Ip5jADmRfZ9NFnuP/OH/P+A
8R00/Gf+duek4oLBlJxdzuXyHM+FVF+OKbEyWDj91zlR5QvlELjx12iooQJ42xiQESShTjhw/OOQ
xJ+rsjQz8+rtBBSmsDUmiJQgHCN1d/1QOpuJZTOKgUzviZ0OGoaoo86K66fLhGSd4a/iVzebRCXK
ntA0BGvR2ygW7g1664UUFJLUUrQXlRBm8loqlgtOu7vhPLiY0xy5IpxyBPsgCv0WFIjnA/W8x6e6
+g5BzM1pkX0cQQa0FM4FrWm0DX73Xfuznphrsh3GWop1hO9KyrWKfFAWjuCzmorUtR4uRfgY2jXc
wjh09PbH63fZiEnYQ0sVfa6kjB1OtLEvQE6DpAsDlMCU+mpozLQAJvDb//azmx/gSWgX3rjBE8+9
6nSIkjwWXE3hC/2S+fBqYAj4Z8JdppriTVzmkKGRey2XaLslDpgKRsyhVqoa8HhFVlJbK5Xg+K1K
k6Z6I/H9u/bf/CCwzMEPxt+LAeI+OWBFXUIjryHZ436Epbtef1MmzF2AO9YhNLUQMeVWjJdyKvEM
cLvh2TKfZiUeKEMRjn6WzDKgLDdKZxt79ATuN7E7kM/COTGeHro4L+MIb6aP1bIl+4dgX4ss1w0d
+djeMUqCC2tgiwf37Dy5gv9XSopEm+jrPMVb3oSqu1/BKQ3bRgLvmavkXt9+i5dto272pszrRGUO
iFr+GY/h3ebP445yShjB7c9ff9Z2TN2Vgif5UzEgn/XkLv2hydWe716rQsy/GuPhEtFgxe9MRtal
rr4N94G3UFLgzNy7fgFxNVCIttDrR06bbE3byWLQnO7LRo7rwxfjRUosPpN95XcrStXZm8XFnnPc
kuwPPSzbg/xkOrXKpeRj8/rH79yAbuo7zorIL/ftf0E97LyzLUQebH0U5hTmx6yao03bCde88i4y
Y7H9kvTzgRR71DN6QeQHiMAuMFJ+blUE/Mzzo2PWiPrcWemIs+Q+qSplL4/aUN1ZZkq5pu/hULjQ
hfXu0RJ2MWsg0wlVpHsUm/9aOL5hUHyW8AuOfF9dUIQ1elrLIhm1m6Y0Jgd0Hm3J1fL0qhtt06zQ
GJ8oMKB9vSPAWjoqXzNxQNCF/kJ35RcKyttA51A8n51rT1G3aUiV+MDqjxCf0MfLb0AK/nhkPdj9
kPnJinkLjSAvkXvKPDjod5uQQcLjPcA9IiJt7l4hIvfUJdk5p1RyoXdsALZRkX0lLdlwcofG4hYn
fdOpLB2MEIwUqpDA3vzIw/8Q7sWrWBQGXkhtF3I5Oh04UAtShSq9tL6lbI0YzbQNwhLLGRCbisNf
cunKkNFiwKjLewIfUc7nfVCB7m97nid6OJ4ou13SKLECGkxf3DletcQM2DQVHByYfsawXAkEJ0d3
SQz2G4ethhBKFsTKkJWhP0Y3PjzmBgxkk82J3jYm25vPaFxUUsS/uOzpG8w5CF/qhG/q/MZHCmB4
9VASNBrLy8MZbi4pD6hT6sBNTzAJng7p1YsQf7P0NseS/s/yb15yORN87fv9zAiURObiOcQ/rQGu
tH7oaZCDTcxI7ahjeOSh2i6/a9DHS+WBFNcOndo7ruxRB7VILTrecwGvAm66fm9rhORcB32RZe+S
aWW7JmyB2Qbs47BWlJY26bZvPPVjSFWMBWydkOS/t06ubyXMN/dghg6UXdoUqtcsK1Ai4VzTc+sn
R0eXOa8Dg6QMklGeYgfYanzIwyX9I//HCCYo1cJ/cArPDfuRZJZC7E0myCMz6xeqFo+ZJ5ul5ycR
LJL4fsWZvhzV0t/X2O3vNv0+6YzwT6n2XVLov5kA1gvTqOV0Ts14ZvHKvtckWh3oAAexraWPkZKQ
WAEwoQemIyjy3Z9aSD/pqx9XSweWxw03YnQiFKUhQlJ7dGfP2BJf2+Z8cc59UBcJ4BcxfU6gWjJA
Mk0BYcskGTegEVprRC19vbeYNiQcwuq0/UIbSB5HHH7LbatMUh7j8usijBoPaC2LCafbW+RH/rwA
RMC0sEly8SpGyWmi6elxEWILdm+muQTj0GXTCB7Z889kXFkKHWZ6CJaGkP7KCmAF611UY1VXkn06
rOGDzddUwrbmX9Hj9+GSjHyYYb1sosEPDVbUJyIV79MGgQ/WDoGeFxCw4aDakr91AlburP1yVqyP
gQjvHQ/GB+8qBqMAEjkAm7JcY48Mx/L6FUjj/4yxeKNCV3h/2YEuF1N2EOW5yIi9XaynOe+/ZZg0
sOOdMOXEm6ie0Lf2yIbhMxb6jXuqHs2cjvv9O/guCoXwoJPJjv7YXDQvNcRrUCRqEPbPRZGRpOIE
OQnS4KYqklchV+6NilFxaRdRp4q16k1jGyxBlVZl4QQp6/hiBlqSq/v97FcjnwiKmoDxB1CS+C3N
d/DHacGKDH3bgtwWvdZxqdmDnj4E3nWInzqClywAa5oNBmdOSlkzjQWu8vE/bacFR4ZQeV4NBZcZ
UxZS28fSKnvf1Foxw9n26Sg/JqpLm8bBU53NBGTAs3PcDohnpLUoqv9+FU1Oz9swwtyUt3/uzUH+
ttHZFRx9U//b5caZ2jxpSzDTF4RxJH0QeE2YIplWp92KIoxFqirVt6H8Jwd7vXT8A7N7i4sF+pen
h1sKpSCL2qJhRotip6tWLNZMYcO68yy6zzvIw8Wf+23ecBKKAE2rg1iGPc/b2A2sMobAA1CekFE2
+tWL1Mpgi1YnAUYK3/AVfrODdW3Zueis8PVnLPsJt1eIexR9PpFEAFOA1n9tZ4tjzhBYIf0m5gf6
/mwLFXmmVwl04bl+r0ILDAorj/kr3rCno7Fzl5UrxcVmIfTbd/5d3Shvj35LTaN3/oLkeY3H5e7v
+9rN+yzRhX1yB7ol9JDx57FtNb/DyZIF2gKCksYa12xOy+MUhBOt6k9WRSI/bDBp+Mb3TBuF/D4n
N7CiMa73jfQ3ZYgq8xb6vqjp9tFUIRvl7OIjJQfhzJ2C3qWt092Y+spgD30CplKYnHArEF1S+g7i
pjoj++yFNskek1xhPLpVJi1KCr5fjD9RFU9xW3iPJoooFJqThWTPSWmBc2ecG6LPvGDipvgtEkbk
9Y09lKtxYuzpFgxQymerNL24xY32Dh2+X68jDa64REQG+EMgbYUIQH3DpX/efjfsEeJLbP1z5XDL
HZPi47nHKjtYEDGYN2bhEo6qs9rihUlkX69jiOLB0S4V8aJoAr8LYL2WKPe07Fs9M/Z0/wnazBL7
xqjpaKue6iYmtqJcSQDvRo9K2GoFve9UUljN1t9LdNbfKdy7SM9c41/0Obr7XAQgSN7MpCUXITpN
oyKHyH1CuxvlR+vz4Q0oZ4lqKwwz8gYi1XW8V2cXu2pgFGpdl+wkNFIW6x16f3qk3/I20xnAJMgk
LYuNdPSwolmNWsNq+5KuzeSSedXUN852CMLXVgP16c0nEv7rpivaoP+zFsJPbrclyPNqL9NMQUv+
37+KCl+RIC7CKe1frfUsOfnJf256Vn/2NRvYKiQVA1oFgkEMOUU7J1qwvyzxffUi2vuSE/ia8aYj
PaYYRBZcXE3GEghH4J7SKnaLjwXcYFz8yWh8OiOKpbB2q6TYK8yq31VSuJURuvkUY/LliHXOrXRG
iT5daWh2Sk6gR/yHglAoXi4v0IbB+DRqN5bjq8NcbRE1kXSc/+KxRlGRkq7jw6x9HJ+796qrgdHJ
u2bxZqrNF3IJDPkGgs6q1IGcitdW5rm1n3JDL1kIqulKdeuB92RvmhOLhuCUyv1buOTUb+Yqbf4E
rngnX4WjXHobj+1gmGPr8EPXRLZGQGwq3uJSDDPXLI5riJ62kvb+ZETN5lPdRRtOXNh0SweWVFgw
4YPqd7ncGRJqLRKiI8sZO6zOL3zFqsiFCBG+j/vgPIWLQWjF1FMPr5v1eVZDQnOyCx9Vqniv0P66
i1iYTy2a+Uurr3U0fLtTAmPP6lGKu2LYXsbbPjiAnrsnp/H5cqqXrbnpS9pjYkTA+VnNGrz3TSrq
aVGNGhbsJkqMKzNMF4gmh8DuuQp0rBqUUXs7vQL1OJk49porpDrrB1jRcX86zaIvjNiGNsTrEgvn
lJFKpN7XW7WKiVb7sa+Sq46ajm++W3WSaabxTVhoCgC7P1c7GEXX7aYkCEaMS0qkWtDE//7K0Jd1
MwrWE6AsSK+RKV6aIISMW6mysaaYfI2VBmi5AA3Jd/hpY/Ic4wVaRyqVu78SUawq7ODNlHtOUkFc
bGcxPK9+QbHJ/qbbVjyksB1H5FprI2fAmlz3DWDqIme5RT4WLfKfEoZTYwKmxeIKfMeY9mxJ86/L
qKVNYIMbRBFgmbwYgIAvzDQwepWXJq1DY5Je4hBElnV2hzv7UY18HxmctE2yHh88wvLznjqvBRc7
2/KjkVuvfokyxwe2DLIlNJhhhi1IzIU3Ph8Mrut/1BozFoJ3t+Dn6I6+5TU4HzVSdODXNF2/my1t
IR89trYf6zw9qgKUWI/6fIC9foTOL9CX+o5QMBYe1p5tKwCoW0cfvPjjGilsd4hwUPUQECb4Y+i5
B4goZA52pdy0PV3fHH67QrhRUxQcdATGzlu/bda6UqndwzfYnQBg2uSvJA1IhALLUGzH1O6llzCG
Z9yKTuVEAfsBUmhB42R6rwjG6gk0X1BCfdwUurKdlk9WG2KZftBZrWGGioi+3MvgjCtxtRJkoVfa
2D0v+bAmqp7cJ7Nv2IeeQKFR6PgUHT7m2cohMAdeXw4zfxX/ezWE5HViYxh8nM2rONRaVcjRxuXq
CCnUsp71r5EsTpZx+BtLTNg/8gJsuF/QpVxqbK+PoX58gPXph1icBMVRmW9y9RosAzR4vOkkFE5M
G5rl8OKVRtEL96OIv9WF/zpamKZZYy0n4TLCaVKzaZGIHNhu8K3bphEZycO+rtpNThOsDxiNgm+B
vq2aoHn6fwm7RfRik1+C7FZZNQskhFgHLOkDFsCBDMlAnnGYTYJKyhasQkqpCrizoYI+GlhXG12L
zR1N52ThkambF/DQ0z2lMda/hEIhJiu1m+SSoHjvG+9ydsiCGaoOz3PgDMezxdrRtHmxsO7IkgCr
hZqzh9BW+mJDa46uZcw2KgcsSojr336Dd8bw9HbbyaWhFZCn7mid8uWAQReLCoqeAmsUhkkfSd0S
0S9EEHH+WhCkKUAR1SQcT4FuVJSots1LxFFm69NUxmVd5w1hM1h3rjFllied3+epY11m5BpTc76n
ryb/O6+f5xwo/EEu33NaVECA503AkyvgaI9+BQakcy3DKI7BNFgJh30pnbKVBqpWoaNu0TsqsRCC
JT25DTJs0dZ8GM9VNXF3YBSN7OItezPLxVKUo7vL/KOWsV/ly2qcmYv2WKJU5ipAC7qqqiFY5KKx
5Hkof9Ye+y+2i7zQTzNFTveJbT+K5MvA4KKB51zNYq88ZaRG8XSZIqBL/7xA/86yVBVfYb2FU0NH
847Oubx5TIztK0VuWEjuQHp07MofkmBBrOQfXwOs2Vhuo9Y4AxRwK7zkVp6giYIZGddHynQXNM8x
8K0uNOmGs3QtLHqt50nk+gnPrgRfmO6ADEu1dXQeiGqNP6CmUEGKWt0gl6BA1buidtD92J5z+dNX
3k/sDEFw2wqvc3UufIsLcxsz2cxWbblm69RGbbvX8kUDQAn8HtiqIUSdkcrNcO0kcXvFUwlHJSUs
q7iXR4SrDtMHXRSDDtEuGILvM62Zs4hR1iquDyJeddihTzYGt8cSFt1SNZklVjqhBP6wYT2g7lVU
HcjkyRVaYYp3MY3D+dxTArG9WnEVzFsXPQuvQEiODKf/XAsZF9fgnn7Ff8mt6TJpmEroGgZ9DwWh
bppXnNzBnDLN/LONdmAydqwnNergRYEDLiIQko+U3/AQM7Z/nCq8r6Q3j2b6h17C2x+8h+hmsgfZ
paPvDXZdGZOwrDIFEp9aVMp+agXbc9P9xONl5wp9TMmyVUpbj96Z6/s9MEWnN8GsI8S3UDMExGBl
5Go9U1lsHSqOlNUj/xgWXuMs+rS8g3TCI7/VMPGSMMO+/EV1RYK3ZKTta56e+Y/0Guas7nwjY+Rv
lu/AAsJDc3Y73HfUiR2QYE+dJeHgID7ANE9Is4KjYLNmXO0LemZqItSFigQ8pKXzQ8u5Nf7O6x+l
FdKOwzTD9Z4veoZnw92ulB3H31rso14wPwSja6aS7eu18ejvDc70QxfRxYaoUczslOzo6mVMYbIZ
KFu4PFCEeX+cxSKjRFwEytI06wQL8isYsGo4E9Lq7/s//jTvX76ANffpfT+8wHdMDs1wD+k1BAEI
lXPS8o4vKfbXJ1N2ApiuXY+j+C65ZAN1Hah0+BKcjRya9FPJAcWmjXdsrjeAmmFeMuvHBU04zZGC
5brKLg/fpwWHipgEAZZFHmRKLPBUuK6yeZXz6YtTchfSPNYpxJxaF3RVm2kgJ8yF3ZTdXmcohPu0
QstyaVxPiYkA2LKWhd9NKUYP0n6zDdAB4l6DohN7UsexNdm1+9PoV2KNWWoFlUshqI5a4mA+zg4P
tFA43g82rMzOEXgTXbdwtgcpI2sipBbssRqcSJy4JAhyGXcjbCmH0AkyLuzW0fVL9CTvlzWHsohP
mX7IuqY6OFsqX0ZP0C4cwyrYu578fD48lNSuEzHJkS4XrruKjd9GDKCzrFmg0p/YEZU9Hyr12BHt
rVnp26M5Ph1Cx+ayXCWK6iJCHkcvYmMBNaYH9GwF++kus3yvkzzxxCDmxt2wp28kJ/Lq1t536Nfc
vBLC3OR5PIHFgXhE54CxXVgBHv48CHQ11ssQoAbEsmpyOeVcT2wfoiylgZvtpEWyMEQF/zGzHl+H
cJ74A0ruukB9TucM7paXFq79P7jm1mjw+yQoq1KBQzaxOdAggvovSDMxsZ3JwsvBK7EACC/0O7Ak
OPFSUDcTe1RccWkrVDZPCKU+vYG7vQFjBvGXFRgGSNZ06t0oLfBcvljmTb3O1yfRZs/YPCbZncbN
8pGNuM+pCG2f7icSPgSLJV/thiPkAdxhOokqTv4S8BecZs40DuExXJ4HhK054t3LXRzD5fhjDcK3
bMvNlrCFvdeFdVuCrkDVsJN9R6hkZ1UDoIzL+NkHZkkUbdKEwegxXXIlpG3oAqP+P7+XAiLMEFgf
v83JvewNuFBc5gYZ8xCtOyE28a/YYv9I0zbA73KMLeaX+WK+9tUpPx1w6NEjbjt4zV68v9t0hxOn
Xl76x+zm2L0G1iw9sJllAcN9uk7g4FVSXxEoCJsw7WZGN9PDLMjChcpJFAM1rdlabtvW5G99wmXV
GniQBdo9/PA0wWxwdWMKlk2GqFdUVel8uIg1fYXm/4rG+X7A2Pl7TgCmehiFgX8qv8wWl5KEnX1M
Qa9vbq+qkqTWd/J9JfEVkKNTV3rnS+3SaKGEMVXsvDGbmXeJJUweidRZVyfdgO2aHQM9Ik0VnWI6
XE5udv30xJAi1qqusIy+fiforrlfuLTbgjYVWvD1lipNX5SyyIEce6oeQjUE7HcHJ9hwB2U54x0M
6DhyElRkl3gQjHC6mWePS5CPYhIKzgRVGlix39gIvfaF/46+Hk+4KLLREPT4ck6H0VYIPjpT/9Np
nJ7fPmhvY8sSFvg/kp9Fjz5FJkd8IKuYceqVqY1H+N1+pPDFlGtkLk8lfNSjOM2RyUZoiiSu/5jr
uNgrstsrAi97Qp/5QAOS11wLLByt8UlRTz1wdQm0wPjBkopuAQ1cirlbzRRZL7RNNvb4LlNdrgQJ
G5RoX3cL9BAtrRGAQjJ8I2xP/b454cPCrxBH8J57YIqg1VsmCa7pGnL6uG7hK7iFD2nM7iqP1Ttn
dOmXBdt4p3Y/tblsAxCvHwGMzNOgVioGQWAEEU2KQoGlWp8YYibGAW1GZyBvfptmqf6QkpXvrl9W
q7ZMx0m2HHbI6D34Twzy4R6DoNqFBNFAEYc+DEF0FAclvWSrGUIPWVapJW0IrUoAC/60KmtKemIm
O3u8GiV6A0Gewn6rMMyOZqXNrmuQhlkFnXoh70HEnK5ngHn8gkMuc8Rece40D7CJN08jbNfYuMfw
R1ow4qlf5MCWU2dHo4GizE4h3Mv0eL6hxlxcveOi0HcynVf7aj1JXj4GnU5XA9/d8+SsEwv18hJo
RevWnqt5LuxZoQnlcFQtUVd0jhVS2p+U2o15Awpkjucn9+mv1ChX7zMVzHagoDI75IDz4U+V4zgB
CACc38YTVJReOY+ZfhwQ4OkYkY/PBbfWHAGLPf9VcFjgMQ8vt5mWZQseciRSKsfkehZPtpWT6QS3
rhTt9KxrHNCpflcomGGz/ZkRDG0+RwO9Na1bbLsITrUcOtBVteIEJGGeYZ2JwOrYxReiQpJ0Zjku
h2iU9GSyuZwmO7REiLpbkS1PNCsAxjg1K32bQcWTwgGtB3EL6HkXRfKMcJgZSg80HEkz0JbmDsae
NaMjAw9jO/ogdx4CsYEJoy7AgUePqYihsNSzzyFD8LcypsifAzrJ9KfdAtsvKiiaaslb4pr4mFh+
uhyYTiPon4LBKS//aE/VHHlqJTdCbB90V2vbcl0q6o2PZKF8UoRaUp1jEQdmaj9b5d79/Vy2oeHH
wqIp6cjqbzHT60fRMjkjglrJxfPlLLVRNuvU3xb5hY54P0wn1XmxoTvVMOvGIsIrT+oyL8EpSHi+
zVdBTdK1wWqrwTbVgtwZfzz1ccGtA9yq5cJvmAD7tM55MyOSaOXx+RnCGCuEIsbmotgNNsKCwz+K
nM6ZJWxz9hwB6rquzB8J/4lgZmsmfBe+MoFJcSEtjRUefkuS5KwUkXHpLSNsyEby0SsoTnkYi/c8
vZYZr65tcMekm53kVor0srXlAAbUiHi053ipcWUmydlb9PqyB6RgMb27NBAs5lWr+kWgoalSI3Ir
BNmUkt5eXxthMn7IVwakQd8H/edhBbfIplpIklqSvHhOIt2jia4r14u25nsGAbrnet2VWB2oATEJ
Q60w+TD9dz7unW6OTsNHC9uIKBy1U3g2GKDWIOy8Qyl2ZyFmxg3iH8zUi0WmNr7CKKKB/pqOU/1A
r+gysXldFiM08Zh0TM128f0e9v71T9p0aeShdHY6EEF07TINWMYR9VxxbU1VQgv68YSuKy8zeyWW
RPVxyTA0zwB2pNJ5h78Ge+eBd2d/fdvurcLo25CCMkPc+mMoirgCaDH7cUN3g2+ozT4GHxqC3oLB
dugNAUb6AqOsysc7fSnxVE8+xGyXVLprGEc9s2/rNt7uhCn1FZt9HmZA0l/42FH77jJLgNdzBBsN
9B2bol9bM0ojhX7srhad0ajRYzZj/6bL7+AQLtAAccwVWXwOpLfYYxqyFosg9+kYKb8GG3MYTnmx
zWu0J0JND2wL+1emOJ+qcCDiSoTvp10HCqua7Eds0Sc8qgtAKeWa4OAu0mqteOz5POsal4Hj/BEg
45eu0bR8RO9rBCf/hER6Gcsel3lZGIOpxn3S0TOcliR8DYycZobckoAhF7EZWzLIU4q5Xd8U32Bh
90tBO2C6IE4IrEeU4BYuE2CeMMVtKHkkeotYMmICrYrjRmBLQ/0D331sQuPtJNYbswBAiG0uTwS6
8z0Pwgr/LH+b7RgKK9AztgvHIj8y03eXZ/HZfGiFvne7aLfR6E7aeYbFF/nKSvek6voFVxyaScCP
79AY54Znc82ihFi2j35azOyFZUbyYSNK3bRqmSSqmfZOUFwnX7YUmCB/tLN9s6+wgBkbMESN+EI+
OyHj+HjW55WdSCkk0WOTWibAsBYgK1kEmJPzfs9Ss8q6LJYJNIbwEnXrXvjrEaIbxO9InMOYh4hN
ZTLgws7ay6zNZpFWs8hRwRWR8HNaYjTW1jswXR615Dh1KFN+C8IZ2KptUy+5V+6Nbp7DugNL+EGu
phlFSsKHpFT0GcU2Kbbx/bpmv+NqhFmhO1MIaGCiqmy83aklw1+3xgSJ12LjtHF6JZoOhkZTtfZE
FQDMEBny2113+3i2PcmF7wA58WFgKho0y9fY0WbGck2N/8u7OuuFZhe/4D16BoTBpnbIbz7G7ekf
gujoBXCeuC3ao0IZmKwrXJ/gNY1b64vC8nkD1RyLzOgTfGMBDg5g0X0IxwEPk2HHx6kH8rj8xjgM
2ntmtqQ1Y/LeKpyBu9WJmmH0zJ+43gp/sImQIYJRpeaVxVIiZD58CqVEpcfIPA5cQLtEioF6pa/t
feh6ERMIya/1ALZSczw/5Frf/xMTvInbPMlgHgKK7ecvpr72wJBzXCp4+nludPxAD9BwoarE8cXr
kbvTfM8y+sDd+f9/f8coz7zzCPHvNqPW5ir7Ki3PEgKhO6qmw7IiIPZe02DtxFS2pM2mcLPAS4sY
q+kuBXInAka/wP/gLGZ58mAj3yzDoDFrCDv6urvjtWNZZygWOJSjXrRs7evaGpFXoMbLvrHOq3c+
kpuq9xsAomSfALvXieoLw99HSGGCKr76MuhCTwXxMvbSGOuSQ2QXf7V3ykny/oZ7MzKaqwYBiDhP
VNITnDSXL7NsPky6u78Fja4C7KiPFKKQZJ5TFMFgXTUMNmpdf6+nFtTS0/GgzR60Fsb7GhD1SI1h
i8v+46WFiehPnI0S0zVVUGqhYtfl0/eo1JHi7WwR8EylHz4xqvhPnqgkdEFG45UMzBMnr0zjRDuG
WKnBhspNNGa/uuDWEhnR9b0DsqRAEhHkT5L3bIxIwFpQQFAWkwxwRiH3FIUMfULZf4dDI/9TNpZE
g6BJmwMQefDrxnOraG24vw/JNRx3/nc213IsftoAWS1teRQKNu2vwPOAYf9b5B1/Gwh7NuQZSa3Y
W8YMR3rqyRjLMh/ia67DIE5ON6gT4u+P/UUHfIrtLbfCu2ZciPVRiqvONPHjseuIk/sn2Jv+Zbhq
mdPiyriaw4opUI5aG+lMrHKaD8/n2HvE+sPOZRZoY5Pa28nd6SoGSdqgADW5139Yfjr4LMB0Pn4s
oqPrHAalXuwxoX7y/axXzlr7KFTF66H1Ws/Hzb6cdjEI8VyfPOQoBk87AD7DGCeK3Y5xrvBTtPbd
XJ7hC/iNMGtbXF53W9Gh3dDnsFeUZvck3Qnj7wY3EANeAJMa+4C2mlIQU/iKuqhncBUCLzXquBy4
W7v9iYM63t9Er5FYEj2w+6LIvjtGaLard24ognwTyLDaKaOiqS/B9deYnKZeAObJA6wY55xOh/b8
XvuvcixOQRsaHjK9Hu+kqIGEYo7LBVx1dVK3kUCxqUn1dcwfkKl+6s3JdfmxJzrZtQAZP9iBHE5d
mM2UVk9PssIPRyWayW7Ar7JWlY2JelDWELIyPJnzUKx7ctbTCtxO/yS5XkgxAx7e70jYaiwbr4RF
9GkRaxvCbop05Nj1rTyVAWKfPdeij2nW8OSmyZG8Mllm1U8o1GEoPisUbLfd/rtGrrxH1XRaRgYB
Rc96AQKnaenRtOneWIN3EsHhxqH3gZPy1k6FeIwMpVMktg0F86sDkNkcaSxRQemDRtBypuJol1Qn
DOpPc5c0NNU0ovddam4ya1Q7I6AVRoDlWPjkp9e5lxcsex0biMbwfE0UxLgoeiRgH242u1sCykUR
zigmlu+CIZZ4cHAX5iTux8QJYB6tDsCi7enj35ks6pnlyK0/4Tf/W479kmloi1BHXlpAvlrf9eQf
2PN0r3s1TfeOalmV/Znu5hrl1Ch6ltHLaJQCKyOpAA3jePxzyTwa5Rg/kkrVF5V5miAgFjS/8MhH
CZKruDAhcBdyvKQPg9IwK9YHL9to94iTTME0oqsgITEitdZTjkmrlZvVZ6d86B0I3txdXFi7Rm0R
jssQYja7XUaGkIveIEO31LEZ6OAqD+emSP5VsDZcazXn61WVUDsP0J+ktuQS46IvVHW7u7RkwlwL
Lvz0ByG1O209IIcggYz5+sxJfQmtB5CMDSt/uh3cI6j7c0KEqniFxxnQ85pAq7s4/JGLh7p30pwj
LTJqDspCpklYCX1z9rZOy/KyDh3ixDWzkrzzIbGSUG18xG27xg82aD67ItOTjhILniT8yqDJblCT
Q6ivLdhtuQzPg6RiOS5xM8y/FVXN3D3EmR60wdbYaYKOxaPYEK3fZFoZWaK7H3pckcwfZKgpTNcF
/z6JxjP1qSBQOQQppTKQbB9ycjcilVy8LTkFfxs81KuiwhkKiVKCH3z9s6e91Y9Kn2FIZUE3UUYc
KHPqLUCyDukq0TlOiecH8jzgLI+l8q0ipOpVIHZfhkOaiV/ZYXrH7++Oyjv01oFcrORUk8vpWf6T
D9/1kcFfeibMaMftOOk4oPUUS+C3i2yjex/Vtb87hfYCeU3yiSsUMV8eyhgbFLcvAeMr/9ZLNZLq
UJSfZ/Ut2kotvenfgOlYjQTIfPwKN/80W/tYgNw0IxdD+c9O9Sl2yDwJKgNcLAKc1erWsy1qiDEK
0NDvoUF/KvMA2lZHwRzPXgwMWGQhxJBvQ40WsyZKJE4kBPmpQx33Pm1k/9zCHUo+izML0zoqM/mY
HYTMPLJHzCqO6GJNFPvXZ2UpqU5RgeyNWcjKttfF6bIlwwkxER60P3fTEXxdHfNan/r3GQjegbn/
xAuDrybVlHRMeaJ2X/M1pNDpZrS2fN+iIP43KHySuJvUfWd088gzRN828WX0E+WQrhFPKApDdRf5
eK9VXAe/cy8kpA01bA2Tf6Rt1ea+aVCPJJLKmoGuSbcReB4UeWQPHh2WpaEKmtEbgT1hWINMsH0m
QxyhJsSt7MY3xwnRuO3xgLTRHjUzCG4wVbLG4ATfLg4kBOoiTZnToFpWO9unmOAaObrALGcEULaz
oeztp0KITriZtqquSUgbo2/iN6tuI6T3xwO+e5p28NzOotyDt/zxqkbToVV6MosMByC5SLGj/8mc
ZTQyvMbUSJmnn3liSn8/517DN4f36Vxtljmtj9eu7G8K4CfimuH27f/B3hLml1BNp2mwvH6SuJEI
st8A2DdxlBkVuuy5oNWy5AMz6DYujUlCKQh9W9YzlRP9J/vlUkZy+ZYkR/OcK0+HzQTcb7Cm3fPz
5mjvv3lBo+YDgnwHya3pEEZVrjt+DGorhiDQw7JVc9kTXOhdeCMssBSEIV/3RpzviB8WQAmq8S7O
7qFJ/5PlutY1oi+ywPuJQfTRzxQU8y6r6FJ5physb3RE78YTF157c4IClYX7+JO0SXWEQlB4Dr9K
8KzUvAB1tEnNsCkM+RGMy6fyA/Q2tt7vq8qkErwG+pqOu/3TtNscE7t72hoJhjd/AqpMmZO5PtfY
eJhVeDriVZSoLOTYZ7nX16r59pBwSxTLK+JAA8+Exal+Kc1ZxmuZ8TzHQQzyBCPp4BXsrr6yh2J8
98ecVJuKgY+1dysgygpgkECACqjbBhJLjFU0+5Xlbd9yeQkJm8QDacPeoCvZWu/KmMRASxk4H2bH
YoF0SqeLf9d2fN/yYwSj9x0f4VReieK5OfGXLs6zETRIgstihNyOoMPefv5oOMeFgKsq/1oFvtmv
VtKUTJhYxPYbvEqy/qFQ/UAHwII4m3zAqCx6+0AFrb62VttghMwpeslRi312zv+iMlOxJxxqsZHb
gkN+4QNIC9WFkgIUAyEQruDniTezjPrtL96JUBuNXm2e1mbF6LDSH6Xx2Obpe2zStRS7RGWOZFlp
h3sJJvzbNoXJMkpQGI1ZGCx/TfVRibs5Zp360+9dQ2OEjCorDTaV3A9pc2G4sbtllA75XRsw6oSM
4eCMjYbz5QhF1+2CVAj1c110nPT+n3+0Te43rsRel8cl8zLsfy4yn5ve43rb2V8v4yrW6TkCwvUF
kyMRD0WRjB/1znAfd9vc0WYUUvBhYTbUoATTwpomLEP/jEl+Cp8i4du/chtQqIrQTakwYfAIn3DM
XdcGcYYeR2Ndn8ROH7auyKpNpJCrq9jvlUcX4WBJ8zYWyUNJllHnHl91nifAC+thu9yAOncSfvHm
cTH4Nl0DrKT7OHg/AIMRT+mn2TYazorGBNBcWo5e6tMSid6CTrpX5DU2ZAArKHvUZuXLgYQKFhtJ
oSL3UUylLj02u8IkgUVqPLl8KeCjVCqe0DNmU/RcLygCfmXBuKDfIt4FNQtYlZQVqAZl2mNDaEEU
b4L4ecmyd6vwLVuKq5hjBnqiwi39clxJBZowddLHdYuiYHeO4rcQ7SmboALBQgjza8lXCNIl7kI3
JeilV4mqMBAWGjkEzDsMfx9JZZ6IXz3ywzC8vlYCyA7CUKPgKAfM3KMxHQT4zxi0NCrjwdfOUrt4
9DaepD800lwslDg2/ysbSlUVd7wCoESYEwOOePL/33fYRZCfNhiA7vhbdXf2YWmI1L4+2hDhqssH
pKMdDtkKgZnusgrMbxu93RcJkYbRH3wxBlFUExguuObmAd2yJh/OtGZRiUAlpTlR/LYhHrMb2bdb
W31utiR9QlLMFR+vJNIBp5d0JY9d++w+zAFSLTSIIbQ+dunMLDkOuWdWDpOBM/8A4TJ6U4vVZMzy
ynTry/W5K9mshWfxIklXoB58/71fgqi/O9mLAPPBJkOrfO+vkvAhAdqTGa579Tq5n7MM20GTYrf3
H4Y5n9rIeTHCNG7ozXUb4+olApp62YNEHXFEALJs6HgtCI9MhpEBS0PrnQHn4PoVlOwWZWMVBV/j
rZPHKl1jWC3ykNXD+5XIwRGYUWVCOvDiY9JddHT0rfMIdvNSyo84bFMA6as4N6/gjEDo+bWcMc8x
J6jdY/vu+vGvgkIk8S8uy+hBq0FJUYM0ASNziywhDQr//S1LOmNpzSzIVoidQXko9NN8VNRzIP8W
33+vpUiPKpzr5hjDhDfL9d+6719yH4ae79EAeivDRj08NQn+v5iEeUbQ8OvHS49jEwOcTOmUUJzZ
hInqQcFnvH97V2lec3aE+OnzfWfyhnyxvxRCrcpl4uj5Vs8B9XkSI0nQOgwkGlVS6uivLi9KYSiU
Xe1HuDEVCbhsZlbf4bYWDTWjYAdFNiZ4XTXE74Ak8XgDrs7e8DznZiavrqSG8YhRWOY718/b/OIO
grryAwVr31eRVQirJAFliinPOJUCTnfL+KBUryIsX7wjFR3BejD+jEAxsF7tDg+tZ6ziB+GA8vKn
ZnEW1f+j6mr7sm3ffguKy34KUIZMZq/cik54PSUP+FYqKOevtD/n/watuTcTUyDRN5+YF/Y4hSAF
6/ELDZQqzKVbd1crKGCRp7EmJiGSExnx0ZIgxbPZyPmSc6WQWsRAlUe7Pp1L7SYbSOVWJxt0lzeY
+VzOW0jJFcU12nJe6hVJBk324cQJywhrElqpgDGXJoYQe82KcHEb2ADCM3mMsOI83hVsZmeYxIpU
Hq/JAb3vbVEvuQmmZ4NHq8exEUaiDqDx0eEhYCBu17gkzpzQv3BPktnOPMMhtSy72y59rZT6DZS1
f0p0pC8ks8JJ+kS3RPyOp8/yeCIPzb6CL1q3mcmzUnchLnRauN8JVwRv/i3DChml8aCErFK6MO3t
TO5Q+QvSPOZ0oTIGvg19urL25+catQLmX8CD/nJWeZq8knSgw8qtjwamCdIOg0CZb1+ea7rq/OpW
6aaX7urs/NnBE86bCA3TQ23dL23Sf/K6iD3RJxDVwTl+rWuzO3kHY1xS1cinumicjpW9/luwewEj
jZgAJrAt0I+Ud2HY2d+5PYJfZ1bJghxXOLO3h7um4uCQgiAcBydfbvDpVjRF5HeDlZyIRs8GXhk5
JGzzmCek0ga2J/EvqiKB6MsGw+yEW49JonDntN7Ti2B7Be8s3X6lpl71KUsAk2vqVAjNTckWxLKz
KHuIjii7vy/MjtewujWVM77wBDyk1i/ka/ZTH0kVlSBDbp6GvVfNnE2OXNPaCUgh21PriTOpvkQm
O7ZfEMmR8hALMxnOmVKrPAhuCQV909O9Ao17LlK5A5sFq+7H9T28K5nbwI1MNddsLfyLEZdZ8mRj
Tf9jJDXSGEUBOwDzdalOxjUFDjDj0O0VR5V4urYdVW8jKkX1TLLRlZVtQ8+oLH9LLsebpz3q2iZr
BpW6o5E9vPC4QFdSPSUzwgFKJLK/f9SASYNSxx5CiUEMlhfLWmBo+si1K8e/MGLYc/+4Gqu91OZw
jX26hu0+kQoANKIJ2wFQVN5o6bqWhUEOFRjiDqKy4YvSwSjR4woycou/RSwmVAM+Q3Dw2Va1zHUp
qrQA4vikC3Fm3li5fVoLf8PLlPkf2KDzDgMq5bzpRx/K5Q0YZtzwcnFVZOLvaLtZRwYVZHnyjGtR
nZ8Exa95fYVeG10NABBdDA3E7nfywHSuMvO5i62e5v+UQ04tAuG6Pp/AoKe0raqN5ls3YNhZvW9D
GAhXsIuYorgrK4yf2ozN5cIR/AHDWklMEUgkw5CBHCeTkLRWoxPK0LlNoakQGkUTq1h9n5wbZRMi
OO1xjpI7GkLBlrLlWYQAKxlK3lZgtSb47nSyhRTlCLK5RHJjn1CJDDwPIOtE7CpazHRHF1ZF6HGV
cv2OB/Nn2eDHq89r7t7omqgoG3RO5eAeMGUfUaqZwa1vefvTwwWbe+CTEP7GyvcBJ0z2Z0o7pC0H
nHDYkXTofwTUDgJf9PhgpSxGHuCqVuzKODfIiw419ldzQ3L63WTWdQBzflrnjbENIAfbQIPhJDmH
f4I7oTKL7CkzdhGq10iRvKhmc1HDi4dXTQ0rfUl8X1ZEQUi4Acgd+llol3GKDosEJZ3Z45yjPSfE
/mK5qHWxrZmQJlFYs3LBiB3TeJ48HJIEE7SPDsjwAoWPcil5OLzIfE7cRYRVECZgg583wAmmvsXm
S3AvkY1C5IjKq7I32h+I4ZAIs5tDYCKo1ppNIn+D/WcV9my73UCxxH55/vBYuzIGU4wKwfN+QAR5
uruYqsvwqSplp1TYh9YdxAL6w4jdE0K8lnLwrPBfpAV/ksm5K1fMRQCEXlZt2UrjjTP+JWfQgBvy
40+hti/G4oUBw2obFt4r2JVQbi8syPgH1ZgSHHZbQgu1n9Xbdgy+8SA0jBqItAI3JxiTL7ja9Yg+
Kg0q9hDzkUfoYcZhBKTsmhAAzgHTjVuClaiydd/QcYdsL7Xe4HcNJAmlRRdOg7EURTgk4pRDNXZf
dMVBrEYqOPQl6XFNOzNebDx1AcNkkM2MlMTmfbWoahnvSP5FlG6R5AGiB5/zsLUZJDK7PHRJOiDb
gL/0jfbS8LdFNh1BZV2XQvZBALLm7wz3nvWb6sBf6cY7C4FN78DsXNKqr17e2omWtRQO6lOqrhHF
LZqphVi2srSZu3nvCJtbGp2hc0jjB/wojZtbcpkPtpMBYW1P4jyN05XKqohqCv32dfwjo9lylpcY
tJuug9gqrzbQb0i6neOOWNEFg2NBPsqQEvP22Nn+a6rShHQhm9CwsGX5C81cNHLoEALpDq7uKshj
jnWyABKdyrgQI0LsfJAJT5QJmOk0olsGBvmT++nSQAEfFbIEzUWOQKCeGniEe81JyzjtQDtjNGwb
6bPzTsaZUOBGgU9i5MlfkhingbQeMaMg+fLtN+VeUzoHryh5V0BjEDWKIuooB6/dqP+OZKnispXR
K+BhqgqMmYBT9aRJi2xBR6zKSL5D4hDLQfKP3Cga/ZSqh5VD8asc8mvv6FM9Vg40MRKVdye5xlil
23dqNxHtPyEbAXfFcteMPFjIz2s2TWa3szt6QlPjz0cJnR74BK2s7Sv1IYPqyMp5AgT6RuYaAQZx
zRy54lwfX4QZtp3e52nCCHurBH5G5tMyHEZMYmxoxwVCJEXTns45ZnPaDQLZrmkCZXlVy/RuTZDk
Iyz7HZCAYTbL36Ab6UkqZnL7gZ/oZX4889/cyqXF5NJPRo+gP8XGCuyAQ8jSf4a9AhvqQ5cZmSX/
tqczwxtPq5bWkf/GxkJpiZvsd0NQaF/ESmnN3vCkV3LCeKT7zqgIGyLzFhLAfNOsoYm3B9o/lgEB
l6JNroXeYkk9UK2vbXEqZgtlMyTz0iSDfZej/z37biuO7Qys++jKu2H7iHRxHVrJ0XIB+mq18dgR
bwyYoKTpWKgzaKu4232H0i2afwzizqCTM9BtlAov0lBw+zSLk8ySW3ufYwWeuS73ujgQ0MlDwG0n
nc7QZMZotriZ6TonK2js+gVC1tO+9z3qqW0DbJ9Nl1d64Nfbu4/nSy37NvxD5OrCSu90n3Hk7I8f
ghc/FIj2SYljihGFD3GJDfF4a/7Mfc5ug3Nbr09aARSPQlMuwoH6pyCBhXW9FRUKjrYv4JW+KnSo
ZL70rC0O+RKyhpF85aC1ZOCS3Ratel9Iy9VJqFt/fq5Ep2dOwsqBvyhQ/Yxn7pkH9TzWOlKsx1qg
G6E7qGtnwRRU2au381WJ8E/di9uxgsVRFuhfqlNRmTbhtNrIijRZSXZlNU2d3dsp+/bZrS0WAttA
xfQ80Nfqb5Y77UebiHctcK8oolifEQzn9e/d1XmZnDIAG3SebuF86EyfmePwBeIEVuMMLUkjaaQz
RZB4917yKDny+KKXc4RzEIX44oIW3BDl70U9pFsiFiWp5a2lr9EaugTbp58VBNHyvWYDFLG/EG/C
F3Cmqat6ieifg9HPYCdNZ2rVLDT5R3BMikm1N8BauP5DW1ClegIq3ZmUnYLA0LK3SbSJdDP0FOFo
qMSl1HUuvXLENK/+ejemo8TiQnpHZPK+jv2WycEjMap+RwSdBdv4NF1D14Q0Jv9iGgNlJ6JqVTXd
R9hjNuyTNYvy91aCbadMSQpdevYwcM8rzZMqvooPQENuCqF6uI/v83+rD8TB1j2oxfDOU3m5ZhN3
ZX0CiHz2L4sYqY9esIZPVGX6kq7l5LBy9kK92M8s7DeTkRrcioJ/4xRdDLwYosyU6JHQueGX1ruG
WklUWN2E9rXKa4p4zG7aNuWfoIUHR3Mg8qTNwXxUBZEdY4DKeL32z/rjep5la1QSlL2moHxO7A3j
aEFpdAL1cvXK19bcdWhNw1AHRJDPa85ZA3f9NOGgi8uQ9cIdoPUcIfzkR+45HiNEXTrL7gO+WCiB
LjJIlNeNcmsDY/9k6ULprNXiUsk1UOAnXc9y/FyXDKzj6tcvdyHbG/YJWXXrdpusNHfU6sQ1iHfF
lHktsS6+gflhp/o3032fqj1ci+biKg3iG2nq7z0eUcYFzaATr0jCpog+y1M4ke+XUTAfzdUYgDD3
2hBtNbbk272XbdXWrl2ctGCOtQDG4RWBhrSXcgIux5+eGyj0UXubv7N2x3vLsmW1K3ayXI4tx9yE
AEjUcSWPmd8WBeEIGGz4nhCFWaI2gtu4z3psXgvuijZejMSjO2BBOnIFrLEfHatibtQcNo14rtIP
46ai3wlNInUlq58uNhPTIBORzLHtIKh/ukYV35HBDe2viaQLiP9FV7B0/5ApjEersQ6eXzSK+YSC
dcpk1xZkj20e7Yt9ypeNuDY/H5LzModETy1lqfPCY8NebeDZd6L4WnMz4ft/xc0/M2mD1rB/TfLu
DgtI0vwea3RV3LPIDE5EHQIS6OByqGIa0jCu48qumRCJ+sOI64L0Q5ixDzLgFl+eJ8YpIUdzqPq+
rEPA8klkBo6kCCGo0KnEgOog0uMIgw036r5bElxAwYprdB0JVUKl1eaLJ+kWpeSxvLjBHLLSvtTJ
9qevqAOIZy6vs/ShJeOyrajsBrtxnvPoDGoep3SaGhgsyv04lbzeXolPbv0fsMv2OL/fhCSVWEbg
jb+IrWCTnVuTUa11glsTpFc9/IkFAD47kE1esdpNdmEwSampvYFhx9UXVCiNM8CWf76ME/ln7wyo
8ExNzW865fPvXtWDQx6i5lDDXpsaD9DZkXqB3CKGRPy93rSpt4lppBhdGplb4Q43W/6z0AhC0zw7
G6y+Rbid8u4pVy5f+m8/S5ScmbPqDO6RwI04ZdWaQQnm95oVQy/rxok1yUNYUpmDxVjItUZjBkFr
ZO8l0yupsgkfAvExvkw2IPib01Wtqcmi1pe4QZKr8MVxfokwo0UuhcPiRYQvMfB15rSgxnK0WvIH
kql1UU7MYYGjvqGtFHl5GTvYvP3AK5kBuqyAmbc+HHBkn5+vugtzg73fJr8ZElCsJDetSvFQHk7F
7nB9YECHXg4EUhcDp+mVd0i6XQP1SZqGMWSUYz9mpI4TeUbA+oOfVs0rmTFmSIvjH+NfexCWDO3X
46pO+y/yM0Nae2nJyWVD+0Gidk8eCWxL5Mb/9WhMsAx6Dt4Bk0bdDUH+vHu67sZw7tkDIEq5ByGx
/xSWTnf9j+DKL4Gr6ykpvtnb5Cra6uN96PC7EnfRM7HNJ2MUEbSieV12dRYaknYljrBykuos0ldF
AUA3JbgF+64awuuNvnkv0q+wpoCLV0Xv2xKUviZz6h2MSxKELOzPYN+TO6+ebC/vqCKUzJaMOG5e
zUA8oFf/mvJBzsDpcui57XJzptK6p3P66L6eJV1uwfgk4yh3MNT5rRd0HG2U6Zh5ONlJ3rYeK5vg
P7v0T6hrR/ooZSX/BZML4+i9bE9ZPpDKAn1UC5p0EmWd6U5WzmSLkE4nCsjxTD1IgkzmYGuy+DCL
AaRjC93wRw47sZes6ypX5QTw3zbVY9E1EUew5S+WK29jcxkqr4bRS2nJAb4gFJbJu1kPR3Ats7ET
9Jv2qoeDbnJx33VlcVXE+pAieIm5zmSizLW/R0jj9J3OnVVZkJMUXr2x82eVIH8sMVWGptL7z9th
l78fF/WghH+HvApw+t6F29XcjpYXOmbVley0XSNXp/i7TXrtGzZnAq5fTQ6wsCCouK36s86VrujG
nGBo7P554AiMM6JFLq2OhAK6oT/0lTAenLmTKfnULvtD08mYxiPvW7IiFpSBGnUQq/MqKQisM+xa
2PxrnZXj2U/uFgGzjy6dlQXcJqpYARw7RzJjVPQUx2ygah7KMPCCerLjNchYdp+0vHW7nVDe3QPj
c4DKkMOSwhf3ABvWW5/PDJ6tT+lkFPpQOSk3Zf5jTJlnOh22oJb/u2vH+IcxZjm4/INOqbCr9UI3
GlD79UK9A//XLzUrns0MXpsToulGjFB6Q3FF8QyPt4QdRlsAPoUE9b+q0TVNEgIujRP0LwuA64EC
Y6waRRF2bM/YH28Wikyg4pYVcyna8BJyN5yxNr2FCi7lR6jsesDyN2LbtB3OpiCimiYB74G41wZa
Qn1y+BF7dnhj/t39+9kiz/FCeNBhs/OoolLpOK4oGZsTmiHAtwjmSrguy6h7qUF/Qp/Nhs613Ald
5ejVsfCnQwfM/4PSeVuq700aUdbicK04ie46/0Tfx3/waFnnhO3+dre8aQNWujrNCX8o0Nc91D4u
xjJZBc86EmwV/Kp9ml7cDxsfQNEgJeQFvfwYsNWuFaTGIRIwtWD3IkDpWbYS/SHLso4f8Cduh69S
jpXoNTXzH0TX11RpA6Z7KEtnRajq1uuwmfFGm8yAHgwQZ5VRJpWpdCfVb6LhYA9LSl3uvSaYCs9Z
ij4Wg71hTQExmCLsb/6E8XiGhVak58Lo5vx/xWwutQlH40YDswek4CmqN6KMNQWt5b5/7NMt4vqY
cerllgol8icEPP3QjCdYigB8utpwQWCTGFhqPwy5RYESHthjr7AzgrpQsd5GmhcbS8meXuISiu9x
x8kAsKcv/xSCYgbVld/gVBkP8PH95AgBViAgvYmmH5pG39wOwfXg3Litprrq4WUgMKYzlJ4g8ipE
YjOv98zrZnAS7CcZbGnpSVXLOYhRz2rWNJxIycNsCiZec/yIx7w7LvC4RMINFdKxnvrFTMBF7KgI
Ksv0RcPkP0HD8i7ECygFp6SngFTqn5yik976raC/fSUCNNu9bizM7zi1bjIbZwqdWQZSI6WIKuoU
UhaX3dkisSrdvRuWmLnScKLBbQvg9h0CHJEp0yMlOxF4489aTpBtH/3TQIXykd5ARrrsLhaUtb90
21zD6ehq5KxgRxtDxIOSBrGDgUHRONr9ueAT5pRXZK2M6sMGNoS/y9GgQ2P9XIrNq+EcNkmnn9Lg
u1M2I8hLkkM0FfdWav6WkUJfS5nhVW0JCovbb7WXZeaR/wOaFYa0Bl2T5iEk43n1SmiXMDQ2KXzF
57HLsIjCWokM4nAfdKlrJiyU0kjOVPBs9QLxwTwNWCiZEtzbPG+yz8qjBMxXRmYqjkUznX1KRPgb
va2G933wYn7TCxK7l1urbFZ+GuZimT/LjdyZdI1gm4uotsEqgCefBY3XzCiHualGw0vxFLxaKY6N
k0V4x19rrBSf9TE5nT2hwl+QssXilfJcoNBQK9qvwh0xtBiJ1jlS9uRNf0vmAqmjmmdK4tibioKc
EVJNYdjk3sID22ezVQTvEsc/Yd5EgaRwpwxBA/6TaOxGBlNWOWahE/u/CHMBfZX4spejgsmlmzn8
fZ+UyEktyfMBkcVV/lgkv2fOySmH1d/LymP1hX658ojPofsbZ9CVhPt8H5oev36rtCTAsKy4/Q05
5cjWuTybz2EZB/Cv+FEeA6kSxGwJfsbS6btt7o2N9g6L+nm/oUs/4I1pcSdlnkGpkDfmJJY7O3m1
xSsIQWYthApp9EmDuPAwKx2x+Is2CaNH/0lBUDjZsVc+u+iC7iCXvp50TdbQmPwHtflUSOxWuJia
0wL3jkGpLOE0maEf78EdJzhvR33dfi/KzWdr19RlIAGK0ZSRQJiHcyhpkno1HVycPogTEyM3rKOc
1cCW9ygiHrdkUqzavE1eOgT+iJq9F9V7tc5GndWRMxeZbbpNaFxN3ONW6qsjcbSEHul5xzvt9sTZ
ayzyd6foQmi1ogpopANywyoRpzgSCoKdNYiaVbmFHGpxVKNIL1dNuH7gwCUlN6+NoVjuElhtC5th
kJo4ZCCQ2CjdMa7AgHERZgMZyV6LpfPir79y1wNjhsmUoPB/yRZZXiqEgOx3VDhAC2ZsYTctpycx
pl4/m5daTxHDMBNmRD3h3KGuO4p5ueE8TeMBHm0EEHercPZbEejEh/D0Q1CxgnND6t/aD2EP8VZb
ehgcYAnVREJZTADAvGFW3jreCR73KobWggTuCwV92sNojj4raHBQzM4jbUpMswhP4Xe/DaWeMCkT
vuVUAv5flpCNFJBNdirQ6+uvNnTf6SOf3HNRKj5/Q6HeDfBptY8rWygVxCmVtdisB/Dy8nafSgZY
WlCrcb2LDX8g0SCsvLEON9Lx88U0SpsgFwpGPpWzA4h6MHrakmd1CRv+md9lfrh+2BI45eESNDCx
F+gjz+NrSQqkIEIsz7Qop/vnx/chbnka2Lw4F6nr+4HRxglfBHhAHOHN02lEKRhLNdf5l/ogTKar
922IQkDPzCWDbVi+2QC3YEc2QQ7eqYtUNMc7KByuVAQJWgSDQuzntIP0iLdECJjzxIARBE6SkTUc
KuPhK0+pZUNDZsFnJrqgZai2PBKaIA4jgSEpJ0I/reuMBIhzZd3RAQMeeLgbLmKl7tkPaXGwxFqG
j7dcxIy3rIeXIAqv+fIYZE47BiVocbMlpnBIk09zXNn60SAVJeZuqoB9Ve4ibcN0EB1BiaklENFT
u/R8Vauun3gR9BJgpO+18dqF0t2Q6BLLK7/LuXcijDHLeitCa++2i8V+SCXa8Fy8rOxLCROSaD04
ojujvCw87KlUVoCtV6Kcv1nxUVSJnXAEr1jzo9lzXokqA1F3epGllx3EUFYEn9U8iL+EYlZePBwl
XeV5aS+nEWqRN/Fi4Y/+xcBXpoJJxW7gpREx1M3+oRjUhpaBqV28OStbGt0OPpyjEprrYlww8Ll9
TJngNbOdQY7NnOOq/DACCPyG6+qQZhnXHpyLPwUcYsttxUbqZ+6J0yosw84lWa1ItmLvfjVtRLVI
YezEdO8jq0bD7q9b5XtQqtvQyDUr3FdQzIoAbfxNnvHxBmZ1u8AoLC7ExQdU5+7wq0dRAbJLOtbi
MzSrGfYK44ImKTlztJu8Zn8FA+9RRuOldoLoBySfUMv0qgg+fKrw2veESfPZMUEJT3dkjfSZ9HWj
2DPhPrCTeTpMOM0l1O9dngYtQrAGg8I41vNfKnEj+1GAPz7J34Sv6IW3HbPLVrgWvZw8uQfejI+H
J7KeBIJ1HR7/OYaXLOaNkA8kF2xcezynkICTeFfxgP9/bN21QDSIDHnzxQt05AsZh68DaXBN0Zn6
0WqkmXSbFsjVIlwK2Yd8+VfZMM9CBhXtMpNH6iYO/JHaM5lrtm3QwKfmB68G/WckY7otFEoHUR8a
jHumUyRE2Sk5XeLdaMyjN/faQ9QBHKC6mmd6k1m+AVLtchgvy15Fb3Q1JdXsq4u+KNW9VUu/Fl+w
Cdp3Edu+8t0nMsc679CpxveXh7pKlDyxIN/bH3Wooeh2LvWBap2S/ezDFeyHa/hp+SQ42Ow6rajx
8XZs2bRTpWVw/+6HsWNXF87Up8azD5Q1Z4W7qMHdUyUfot68CNIg0AjdV3W1iCC+ELXR+8a7Ba19
nqMQpc7fvgdTamMhJmDjdJWUooZx4mFH66FIrhUZK/xguiYNbycQbjpi+Qivx7838Xp0VKD59qqG
xVho9K92oNHioIJV7utBV2Kw2tPbPSMhA53io+/vy8G2cwMENk6sR4WXUR0xiuD9uLHJeipsuf4k
w1z00YjBQv0KQYjU0T/ZLtFD8G46JZgKqqAoYKkxo6d6q6u44ebsNDLp9lqRqtnk9UZFYwC0DJTK
B0oM5pmfWDdPpLjH94Nu3WooKaPwPLGaNYbAY7Z5yrgBcz9gOrmDs/MNBFn5Zmlp6o9PgTOxiVub
P5TxLYkmz0Mq7FfehqbO0KYyBZKpRzPX2vlEg09AsPP2nKdkFSo2AZlkgJKp6sHNODCjP/1iKKTZ
+52JDkoeEDOuXGOHcEG9xTD6ErwHypK62ch978hWoKkwW5F07dDH1Y6Yvdoh7MNCeS9FyaoyZnXV
mSR42Yt3AKGNAhzPdYRHankehWa4VcuGNZ7EPUCLlDGXG7lGMgW92wSi5qFHK2y+q+mOQyXJ0O0+
B+/O6iJgFTHza88HFntf3MVLn8yMCdgNzsNrAMyWz68LvKRbsy2jvBJJsVKwfWAplxJMU/fj90SM
jJKkx3ZrTuqM3EllN1BOOOwds67ehy55M/QTPHjsofNI0XfnmByIqs70IhWqmrzUha4kE92SRjSa
ecKmft2nkx0+vtDIrjs8yM8M+7b0dW2KO7VgbKDpGvBELYjRKn82rqZ4lEgo2hm0oLr0y/pa/JPc
IXtA2lhLXacaGXz3pFebWWyLMTRg6MCs+wPS7bou5i0AhRKwfTH8fFeqMDVRHH+3ZH14VoNVfXNq
GrklA/jkJYRjPNbdgZMpS7il9vgp0p57tTEa/Uhw73QLPcDGfugu4cYXnK+7SvIOgOxGvO+L+tHI
09UWQzs5nyNY30dv1e4fBQDqWEkrRPFcZ3UdH1zku2HZBJpmYcPH0z2DAIVQEgCKBwgUwaFWAAcp
ZseFAd3cs+iCwlrATNm26nQeuTfs8HKzlBQQ1avu4h8ALOftv3RPgw6Wnm/CUwBbrqmbsQjJH3HO
jkmU/oW8r/DuDJ7TbOi9yyJ3V7ry7CcQrwCJQzSU3nMFEi2mA9LjOJpRiYPFbIY28Byz1llW3qsJ
aU2yDTRygYNzKqFAN9xEr5lu3SZ6pwHlHo2M3Nr0KkSj0IUq/RKNCfB2BLEsCXvRN9SyRYX55XNM
A6aSqofK1SboafHJyBvwSndYL4gcIVh8m+H8uhOODmNKvDsUzur/KTMXLisUvxQyhhiIlingVZ3S
O/1NMPCmnn47Ngw9l8HwZ/nFEk4z2VWhprWviqQ+WdK8H3BRHEhhATD8ApJDIAGynPUk+mZjYQRq
ybNOnoPUmt07z2vLFH4QtxO+UsbuWrkc6gj4QaIP7jFgwSJp9hLSjtTInuQyRKOfCufwPr+TTfcB
iuOMQZ8NBdZITQGG+vh1OaOqP6KeJxkEnk35AvbCRUl9pKj/Zkzq+KKIm8nhSCXu2RcGN41BngW2
2cN1Riuf4H9mbf/lyX+L1qtwcXbCO+Z8HbOaetD+Go5ZjyggBzLZmNFSbwh9SvnaFBEOwsRY2wa0
0NQvK+/M/Bc4pPyNDUSWazjK6ZZUMC2EswAqfqkAV4L+lo0ohjZyuceSb/GQvBRIP2tx449kh2KK
awqe5hbe8TlcflCRq9xiUc8ninH3CppAB8223XLFnu2LnRZisbUK29Z0XGO8yFiiJqGjrGQz3OEz
nngAwK3qah4vLrObuG6qRgBS3FR2BRU9rim5aTBBry3S2kqpzMwxYRpYfHRQfyIfWFus0sShByBb
lK+3DQ2CgQ3EGkQ2lcrY5sFNpR/B5dclwp7Xn/tHmmD1m9hqHY7n9yDsMNfkUwKoZx0EV+0cMRyY
arUAJeLRuj/elpWnfxJTS3i3uIjtgaZNBm/bgRULofxZpiU5W5rXOJV3+XMVBA1FsuJaGeCP+4LU
mC2SVCA9Vzp+v3i1HOcJPgbNVBUze9it9PRQZ5tKo3zbsqGdntPFIbpToU827fXNdnAk/b6eYFP5
AGYVTbcU+vgU16LtFmyrVDZaudCbaOTAJ3Ao2aRqTAcA2MaxdiQ8j9l9v190rjOVMPg8qPiwIPGC
qQRbesGX7c1qUQD1Cj6tHSmno50OOcXeXyfFmszQdvJlVOhbJ9D1imug5awAWQPeiKgMf8K4RQDc
paIvAiG4b8bedCVr99yG81OXaJSEXWpgjLO3tY/Ymcq4s4qJTabPCsqkQyxSy9tMiJjUmdW8lElE
Mt8fD413J2ozd3Ds+t/ckViVSG+st69BpMh0l34HXOPDzfmtqY6rUoo5E4jYesxstU2zX7jvcHlc
GXnQIeqhnsZ9NJs4Ut45U44xivSmvexVtGZM5f6zv0eIJR+ylHhVJuGtvcNCgctM1syPJ20rzLC5
pthNlZGe/FAFY5nQ8Ec1pyHcPCegbreYkB7hqzkzXENmdPdz4LiwbDApF6QCcfOsVxDrG5xPacoC
o+bxZBdMgetKco+9bPIuZLqCHAPvaOfDuYl1BfAyWl0Hi8JpEdzQfubmXxxca+lOASA42FDDF8C+
N+RMJ5ay2whbNAxL2hLsY5sADuC4LoCZZ6pw98lmR3nkI98VvAzN7jhyz4sAB6nZh3Lb2ZfSDZCD
Z2psEvXYFQ/MeEfOGDn47aESXLpbmC3ZM2NTeWGKEXxt7+2sWj/1vYtf9XDSlGrmFhh/lfi4HGiu
I9ePJyAXEwgYILL13aKyZkPsYAU8RCtOJjp+S88maVca2g6tdZD80O2W53gN1GbMsjSXcJOVtChV
e9miEZg6qeGWEhy4RadrG6ACHlU1NAF3SE/8NnRQDr4ywDvEkrDx/FSNfC80xt52ZFykw4DPGuwX
z2g8k48XNIQZVy0gOB4GvSi7SETog9IfFxyw0cRWQWsd1eYpevl/jf+bThuyUevLd4B7rK90qUR2
BhWSU1VGcUHUjPP6tEEMsMS5tDoL/wEDO38rZn0CYqJoOwPVAQCBQzJogylHzPbvnFRu1lP8kdDO
ygSZaZwFFiePVmG8zXu6odBToO++eUUEyRDiLUdDgJxeME30ywgNSt8C7pkKkDBdUhAntoPwDbpi
4n+cSz6EI+SbtrXCu7KkRpoX6LcoUxtYawUgatGnRBU5Mg+7Ejw7nlzDNiyNEbIJcc1v3C/nfpV5
eK85iZQp69Gn2dREBIW0Su489fdvh8rHsDEAkuH8wwo0fR95aoA5XAWN2A0AtHD1ufzmSA4EWzaV
/zCyEzV0xpaNmLp5LCL8Eha+nVqrZNwmPBsw0/B4yEQYHbg3x+4dOY6mzwz+SCH0Cx+DRFLASLOX
I9XA9L6TCNm8ED49Q4x2EWZY71DAAU2R7beb2TcOoiL9Dkw4O4WWuCcYrpvQNQbQga/rd4vh7Tt3
dXTeoBTDc2CHLmlzxXGnn42M2AEHO7EQwZ0tBlkL/QdS2l1Ft0ibPBEdyL3PSkptMdh1ggsbrpiX
SVF43Yz3lIxvu9Obu9ToZYuzkPz7W2hKKUYzZ9Mp0d8BwefuIwXk0aKBN+SuK9xASkXIs5t9zaAh
D4CIetQCypJSsNcQb9x3cHEFWGjuiyZtWibRQL91zZcrROASOtsXBYsvVbs/WxXvfk+SLOxNWj55
TbT0LU6yOmBShE2whff5mbuEzGa3CspgIWi1mWkqRVnZJUc0pS/k59frZ1zA6RUdOo996wjUZvml
3qI10QLAxv+u9eYFV06Uyf5yeT3i2/sm3QKpoixOiPKcpdoGrKaWZRjPMzhWGH6941+PE7focYv6
QRfo9Mqi6Q0OFr8oQ1rHtXwXC9wMeKnmyr5u9DIVS5dxn5yG9iXlkhFrwESd68q72ILQmb/a7Ntq
aPlqw39q4CdNMDu8p+0k1pifAo1lJZo4dwEzjkHf2OnasbI8MOqFgmnnF8GjCtN3sdq7zU1YhDZx
dA/p5LKBxgJHMUwqnPN7rIHDVklzZgm+am3O2Ga5cft5wB8Cjp9XXLsKi2ksgs54bpRLnrJTMA18
IUBal9UgrVPChWZ5x05hZGm+MKauKuumE+BDmnmeWhmmx1Sa7M7lRYFKKvHDg3KxonqhxdnTxo9P
ysPj2hRaCyo5nJyV1SNs/oygXxPWI6EMiG/f1pX3t4kp8jns6Mz2ACtFE2T3z1a8sCPKZ2P1NPGE
evugAVDzkM+cIDj4THwuX8SZ3wX5aupuiiOAdBhQN//s2CCIsudL2OyiiebDk/qrNZvqY5Matbz3
muSTYjOi98WGE5VXDwJBG6SNpi7wfvMYgcYeKmzTHyG2DBU37/U+lqStDkOUHlw8ydLvgpB6Tw3m
PTDQZyz1VjC70COQ/MGLIoX0aIokloIq6MHLXYkTVsQnFPNP788aikpoinwahx/JG8l2nwil3J1L
Pgr3qS453n4NTcYWgMunKDyduvt7NFhRR95BfJ7BKTGtYrA5Ea6WQol/mzCAWhF0olTOwsg1KX1m
PrvPggy2OjX+g4n3gqx9qSLVKYIKIc0XZu+adTn0pGl4ZevWE5rweDtM3C02b+QneMjwU/NMrEJ5
jFEawquPjTvsWY+JbsROKDuOGbPjZxzjsNwXgNpbQgOveDiypk4JehyzWR2wX0xsVpgXUzBQ41qz
E9U6/Yy/+YyB89oY4X9iMBMfPJ3xis9pAd3rmwnsX6g4d5JGwa2rQ3rbfNXolEgb9q+LAn/CTP8F
Aw3Ynuj8atJayHHu5RpzW996afrO5WisyjVeYm1KLd8QmIeNmJNE96etqbCiZy+NKCsAQxu1fdcb
E7vu5qKVIGzgg1h1zKmecpVslKZXvkBqxacpi7hGDUVOMqiYqgyqWYuGEYmrf2OKg/bE3mBjqeMg
Kjl7xSLYrn5TIhCb655bEnsJtqTNkRKPDgIEmwSPWch6eMyFxMxceH9x+SmQD/n5WDLlZAx04qKB
oK9BIt6m5Huoc/mwpV5XDE9mTEKWVnvIGYQTYEiqQsPPcpov/ntl9kWtZn/hVmGBELmMfHEo6alo
Et85xS8H8o6fAkx/aYuqeFh813COAySGnVPHWy9C6y8qxnK8YNLs/KeddnuAkE0BHBoreabHknIR
woshmvGx1IH7PTBHrSbbLhWFx8I4SK1k2705A2ffAbcAP8jl0aMlMVp/iXDQrdQpWftpJbK9Aqtd
P7DADZhM13Us6FNEPkC+eB3ifGs43y7OckOWuoFBKj5NjW7K1Xl21bzVqCGBRqbv2pkkdxZRUTvZ
tN3EiOJ/OyCefTKqQmQxSely7hwjOusrtL3lVLIE+ig2mvwsjOu6ocavyGfEDLOkA4n1QCW1kFyG
cFRrKM3lN3szsHY/uS0W4InguwlovEQ7VCwOtjV9ztb5VMjUCGnVZwSvHsW2CW1pKHWuGx4h3ZnJ
Eb4Zk99yBDTAMtSwPXahnTbUZ1Fi8I/vlihQOal5eXkGrxxe+RH8/uH6y8lAPRCJK2rTBzfacnUG
a99g7ubWfKgVTmWFa7PnqlH6Htf/HHwN3jdGhlTXOE9z11A2c7VzOhU/j09hH3Eyzf+A0Wheo7pF
qVwpQWQ90d9BvAcyMSKHm1tr261IeyUftiEdCPZXoiph/PC10Igolc9+XminWCT26vRrvvYfO2uu
c1dQM6wFrtN4vA1ZZd5YUMwnybD8V9rF3vZjVrLXglJiVWBYEXf5/u+sTQeUxcBx7vJ7NEqbb4ds
eXS8UD9VU9ATSWckH7Y2+sed0cPTohYjyH5XjDlNjzPpe0JU1yu23PaEkyS1PR2+I2K3trijHNr2
quZuCf8VjndDlZkxf2LXmn+5LAQZk7AqtFNKuXkaRoejlZ7EH4nl8+9AJpaNIJe2LeK3FZGtsmwD
OsCDiwoe/hi4+EPvM/l/OaFRUF43uhu+jSTAzuHqhxHLq43ixn+B//iSbFTzcNyUJpSdNpqJXY0z
B2fKfQ/zayE9JqAaLQldnanEOZ3KqfeQXJt+Sl1UNqU3jPFZlEXCgJDUmiw7b9byHtg/LX8vYoIL
T4PKM+CIF3G9UlpNdElUEKa9yO1w8/y0DAuU6ekyhOa5DKgbvuvUFZ/X0NBjgM8T/L6H2Qn8Fpzd
1N1z7uOizSpfJ8Uz3LzLMhXysZ19Rg86FgcQGKQMD/cr0Gd06lhEPDIpfVKOsAbc8OL7rPy1DPv7
ihwqFvqrYolT7Prdm9zO1Nrehr2Sk3sqzfZyhNIGt76N/Skle8RcJFhUSPHUAS912d/las6oKrAw
j/Kqg5jhwkEtn39s76FkAQL4Am2MCFKZsr6WgMjBV7YOlFKbJMgikrw1pvAqrLLEIsEaQzcCSdaL
QTuhivTk1J4o5tKmk0ISHyeNbqpDMzup0Eu8+GXmHhOeIG1QFoZ7PmtZplODk/dZziMg8CM5muR2
P066+Fo95zHWaJSFL6XdNY+DZcgrEzl/V5Zh68zUdvwiGCvlLvSawK0DbQV0ibXokQ+e1f+TnqX/
KGPPkKDWr3as4HiiQecV8vfcro/4/fFyhXpNCqoqpDshCUqqnDkXyNrmp/q4J2wtSiMCwBP1HHVf
09cIuef6tTebLTCwB119fAsW4g6DRogGhwFE1WdVbkm7IbADv7d0PII7UWHsyIYeso5ThEoxC9kv
4Ng4EWhDwUGCkeK26veOWf9W4LDzAv5Ff+i1bhSx44yBOVZikmkHQFtXmDF3Ghyor5jj//+cUio2
JpTr9Y1CUl8gj8SwLcP9m2vuJxxCN1CsOcIlQiOngIumS8haKKZ0amSK9zLF0hSzy4XaV37fo5vb
rAVK5FKoWlXwly4G1wdt4jlTGhxRl8fE1UaWrpGNxxi7HOuf5xBN+kHN6EpiGlLXoLn9B5Jn1YRf
SHAPpebc2zKWz+h47ExSmmk7HadGc7yhd+gzeUT6v52iu87hX1Udz2QV4iObSGGKwLfMGOfOVMV/
pBWB2x/vaoZeRG6sQQyQCMviSzkWCeac/QV5f0Em7nFYba32GxFWlmujnXfroCcIBuumX1WOPP1a
5aveh9bdXgC5E1Tj/Rvelg31PlVCtTmwNuKPaPF4JqGWpdTvg9gObN5mEudQZlJwedF8GtSUcp1f
B8HFiA9ZEcj+9W6ZRx6pQ6+bzmHygm8qBwxHc4ZBzTrbC5uaBc7+L0/vKEUNG1Y4wyjInJMs0pTO
UL2lCN7bOiiJ6fmeA/VW2UpHmPdHdfw1OXg1E6OCst7uIpghEb8WJDkT836EjOQnGjUfGNVUhv8q
Yrl4vrRpyjZ255rrqkFlP9dqzVPJCwcxorbboq93+yAHVi2I36nQNd2p1KXVfDe8vg5HwIjAwSeL
UP/rjWk5WMRSoYf+PdDtrwvKtbXajbH7hMYjr655dsJR0soRSvQs4YhPPyImIxRBoY68sN4fe/y2
Xua7IW8glwl5PQilN3RoCwZCAwOmWOvSEjLkVVaEvwXOK4BzCaVCa4Cg5Wx8uiVGVBpOoUh3yjav
vrgv0kpJkSj3mhEkneHx1Wt1dBeqEb4ZTtps0Iw7vDmhtVvhS9mG32xBZt9CoUS4fsay7/9HE9Ze
Si+dgULdi0rkNtmyVhLpJvycu9Ec/Yep0F4j4+MKjEIcIWoLaSw93eTkJqd59JK2CbvPaFbw03jj
t49rIObgP24YyZqsUE6K9fPOjTPdPfFIsM+iDioTdYH2K1FrYaqQ6toARhOv7tNxf3sePFUvkttj
i4H6VE/glEg2Nw9MborFNYrR3W3KnIrTNeW++BSS8Wa1Mb2y3ky1wzyfx3sMewWZuPmkPW1lmV4V
G/7A5O1ci2RCzDkQ1+EQ8AjrO+hmp4fk9tM1eHRh1RuCQ1ruftQsTRRx+UXu+ShyO4zSs4euzxmT
X2xVGmB8e8LWjCkJ1tRXngYfteaH9kzsIRkAQ7xzdT0IJaoo4X3XD3AjkuKUemxod8vNCwJo07+w
7TMjK0s9zHT7PeG4XE6P5Dhay8WV3SM1tH5fGS7FiRp22rHQfR4Y1/EdfymbNDRM3JCarIOi1GZK
nnuXjPAzLX2115zJD9xWNpFpJ+ugaI8lJbD1dGZLEwACPbWjjwt4isrwvKEbOfva7Y6tnMbg1uZ8
p4qQkVuwOu4PGWWyGIAs6eUrAufTu731CdXRifUCTca1vZ4aBSq8ppcncqUhMHipHcStFGnvO5tm
X866wh69k+K8E+rQOFkZeci3EKTZtFMqD3neKfZCqHpTaFnYMDyJg/FrcpPwSPgKA9fWJXaLmfIU
LCQl9weKOuRRuEToZfg7GsdzsL3V0Stf9ZNYovEOHelSfydXLPu2igNFmdpXcw7IdEbKlUe4L0+M
uKWdTgaHVAfNMmX3olNsGe8vGgr2PzitpH2dbPx4spxwqiIiXLUhdt0fhwMM90DL2VWPC+72KXht
GxdGSaB7oMQ1UtArbIAKk7LWagqI8W+UXDM1PE831F59fXvKk3KlEJWsZMPA7U/eAsjcqlChueFw
bfWYQa6oFdPvN2Whep/rdxDM8MovByT0q3kA7fgKmf2r+n0pY8kq0wTtT3W/lHmxn+/TqpqD6Mqj
AIYRfFyHAwoURDEtdO+5SaqckpZ/wAOXuS/aqbGadQxVhkwc7g52AUAgnv38WKjTbMlPtVZycAN+
lvdUJR3P8hAORJ8rBE+IPF+QXd5YyM5QFS4SPZ6uBfWbVfNTK/84Qv4zHRIp8jrMrvuEmNUzp5qI
xFwlkeZYsAoNr1rSBYIR7Gm0PaeuJEbU1MyisOs2+kEXelEcentV1L6WCnc/EZfAScmxtRsJm7nx
kVfN3NO1BIhKIYJH6R+JYismwAtZpCI8zorHQoDBAew6od0WFf3JfDqUKzYfZdz3A8g9c7WkK3qO
VFBE76894HLBnH9pgmQHcPcCC3U3g+UoEJC4ic870t/wTabQa5IFrkpF/Jy8iIaZaDE3vT8mIQP1
NbF99jjJ4HKadxyfA8lZhEUehG/EUMbrXSfjC4K/G1AklASM1BbW8WjYRAhudLYQNf0UwaG5lBkd
1t8LPxGowK6MxIypOp34dhLkyuazlPMxS0nHbvsG6C+UosZT9L0MsVdkGoBvkCRy0TajRJf6yfKM
8vM2DPuH6sso9QYKFahiD/KOvaJ1qAyBwMfVrYxj0aQzu9Gj98plPjnPnRiqwrxf5zCGNzuHdJ9v
Tu6kLGTOC/jcdemcMprafwjFF5aocyghhoBLSUhj1TaoNtn/oK+pCz0rLqMARGzluq7rXaZIrioH
n3f01BA9Vatz4EH/a6dbQlMl/j/MSyfOVEsGcwOiz/UWD1pQHWolfoH8VdsjV1eG5fsIBrXY6/ph
+mPH+iJ2rKP6Qg1g6ad5nDBjSqsoBkFqnkTchX4acTfs8XWvUlD2JGH3IRmi3kQonRq4UJCR0aZK
DxzMoVAIX4qcTZP5AtwtI8vXKszYWYlXVayK3LfkliQ7ANj2oshwJNHzFTQSMw4VF0k68uynbkwp
rqSzxP9ym1VVnYaWZNzr9zYdXuHEI4jMeA8ZBuKxTvgLrRz3Yovkq4C0Ah98wRN3oBHz6BVxrW6t
iY9k/lz99BfDhxUUQqcQbr5r8M4LwY5yNd7KlNhRPcgnAHLfT3OrOqgmtM/suO0L94efL8Sq0x1H
IHCOZKNgfdOIemfrqe88nXnXl+0TKsO1trj18JDbQULLTBx2dFd+/vkCyjTDb9Jt6qLRhNXEvYEz
iyulAOVCAGgcPkYhMkIX+owDSPyWaSCZqihRyKEHWPAS01sA0RjiP7FEwm1XWtD7vqtQ/ub6P/IU
EgM+zqGVInSyggov1aG0WZ53Ez8g5wom9i7+WU0cD00q8Lae2cRVr18O/kY490rWtWwMqbxKg/nx
ZClncxmPW20yMt17Y7RxhSdgjlca2e54P1RphHxbpHw5s4kqbkAJY3SuKiDAVC9U+h0JBzwe0q2I
vE9zX//gmxJBMgbrOjOcV0gc6W0h65A5/mx5wBaM1zyRiqMrgPVqupV9v66q5gFxsOjkNBVwZwPM
lIOOLlFeyPAhRpFYHTChvBtzxLXuxYsVcCAArSqVm7MAXsy9GWXXGffSEZCEEQZUz/wOPCCbGH+M
jLG97jzu7/cMUEQYbz+USpKu1o/oi+c19m+IKPOoXwEQzMFPoZZVFxt6on2GIwe7W8zFx39mlGdL
xNBeVepE4T2CZML9CYyL4sjg87xTnEo6bDXXNLXLGjjjzKGk4FUEHV6UVFn/6LdSYnxeLnZc57iC
nqMrP+obZbIHOXmbwnod76KUy25gXawt0oYB09kQ0WmXb3rPz77nZvtLUB0jPuLeoOEMWi/6bbV7
44AcN/r8RF59auLnIpS9TD7jc7amciTQBljx/TiffF8Cq641+jjq2gYUpY9R75yvCqHlrPmzXo2u
+upKbDIYNR8rsj9QeRZGo1MhhUe3VBlO/QfhWMgDaJxLoUp6SOnJ87K7EwTMekWQ4b6TczcCqZ2x
OCjz9WGGUmfjHf7nu3pFuv3k8JX7orIrC90Rw9JBbWBzGaudsmdfByAoHHXZ47/HN/oFxO09uNBz
ybyNf9nh9aileGJw6sPhLxmnVWm/OZu06sU6RMSd6VSwYX/YQANi+kNOZFUtNdXuLW/zd2Pgf0qO
XT5JJcs9VpcQKPU5Gi1QxCB3qV6smxy/apOrALYP0hE5jg9tKTK3txRj6ejO6N/LF84lzSaUEsQ7
2T9bDaAOfxO2IFEFowGRowTr9Ho4ZMIla+CL72eIES74omq3+khWQikJHscgc8ds/9F00PwXOAqg
KV4FbFj7PJrqiKJLW1S/18Rzy2TSllEjKzFJKbOjIm+kfJ8KH7JEapWIpBPqQjNL4EojoBe2wyMv
8vM1R+eyiDcWjki+TsWxd8wnNbM9ASJVz91vpFjFJOm1LJQmsw2qWNz6owgqWzipx2z484JtFzlz
IcWLiEEVhryooQuUuhgfyi5GjYnPhIfYgVzbFOtjWVGeqfKwKnLwvRuXj0TLyYdGMOCXXXmhtXjl
IFDASoBd48bCEW6A3Oup/OTckbZ8G9R4wif+uRizIkrVB580T7gFyisYXP1qhqnI/UYmV3rYvpoO
v/MiklMcRaeJpa9cDnRl3vjnSjgeGs+Dy3sv+Zi7j24WnGSQFkDHd1lmPO55dovPPwb+UR2tZP5/
h3hJInfoBVG64vqTsLwhMBgA0m8qzqStOiCSEQ0UsJWVdCCnWlm8Joizaydf2nSDVmr6eGzcsdfC
KuuV/7DdziRyUAWTAkj05vD8iJsSQYQkMml2FhgN3TT9EiLfLY5MrA/fZfLji2KsHgl0rm7n3N6u
uVPh15/SO3wAk9i0Ocb+Q1JlzhKWnDc9auWCL/pFHnz+2iY+32aASB9fr5I3yXVXePd4GhV3gwtr
8FYziP604VMJwYDlI5fLPTXZoLj8OuIUl3rkTaR5Gqf1C1nHcU8iDWILjQ53Q4vyoXbeqQgnJ6eB
B6dkhN2pn+WfOcpywyGlLf2eqRRg4g4edHtgStzf7kpYYbLgw9C2V+x7dsc7XMTXe731MTsoeSX2
PmufQ4ltuJmF6kVmyWQ2F8nO2a1K7jwWBLVf+7lCUDcnAW3EabAPw10QpbJXg4PW9NuuZrlkyb4P
cxcBWWw3nKvne/kKiHRtHCt8kCiR1GyaCZvHFBNbSuM4gC80xMMd05qaZKbE+oSaos9+eyiQnfKz
IbdQlJ3o8dTO9ELJhjLUigcXOuu9VPT3XF/s2dmyTj8qn7/eah17/uH6ftfU2Joo3GfTbvegZG6b
8Q11McXZIKoWehEXi4aXca43dwR0OJAVqhMiaAK6T1/6nVEiGe2ihoJMNgqblHVSW9Vav/3TSrdd
WR5IIhSJD92PecvKtu8JTf4MH0vcDbUQBKX0b0wg3LQVC5SLz8Qhd7hwPtjPkjlR6dXTLoH/h04T
5n56LRFaDg6meloLi4v/0BF4mHyXZvnizepMDYI+PtRlEbcb+NmiZgiZgNuc9KuUwUMBFHUxP7i2
5iPIldFX0ko4VP8XXaQZIaKeY2Nhf/urY6ZV9XHf/LE6dnYWz/i0ksNhUlNfSYxrDmMF8VL2CRYc
lwqiEkMojGHlksAaIVjWmF6vKEg5+1TuaydA6Da+8Ic0cXnxIhZVHh2nG5Zo2F/j0tN7NH+ku0n6
qTS/3s7/SMZPJz7cqSGDgkoqSvgBYx0+pLVRTDM018Mbnu9fCwwNIyR/0xtXcWPKcfTrRGyjDcLG
Vk4cgk2W4m3yC+4fW2W9u3ro76K/PvprmoBOx2FsFfKpl5dm/fEyNXF8jFM0k8Hg1UKIgDAxrBcy
yNwmkOk4PVoJKVol3s5ZOoqse28VpvaWnLc0tOs6yd+Msw/liSVWlixNwk48peO/pX0rtX84FR4n
AFBswbJoKEf1Fghuile4iwLKLWoHnk6149JBf+9n37FWb+wikV+SfKg2v4Zwavssp+fqYR2+qYOD
7eaBfKcH8bhgcaDWUbWx42H6xuvI36l06x/6HK3nA1MX/TYJJLb4NjcEfKAWhqW0xrFcwRUihj0I
c6jJlWhsPe8+ub3MU5nwzMopYTNm7gmnv1V7sL1UqceUpPFa6u+Lm9/q597c3kR8VpFNs5U2Lip1
Na5EfPMwieTPr+JwZaNRzgqMYRBPYQGLeu0McWd3UMjNOZ99UHmdNK5xfCZDKIPwYsi8WD8solp5
ejvgh17yg6XzRy6jlBMQbzKGc04PQdayrJS9wR/5JJMnLe6WC/P2zUZTfpWcCMkINsH55OpCCumW
Ivjwf5ExRy5IOSBJHVSO4k1JA+JlCgFcJ/qbyZKLs2cGV44z+SwNk3XeUnDTkp0Kc2RixKmUwIeO
Q++ei9p4kPCNfikBle85JEp9kO68+6xCgpIcnT3JRnAPOk8hc/NI3M0s2XVVSQUG8H5si2rjolcV
l3W3ktrQ/sMmqcmUA4SOAHGvkf/r+G/nUelSEOLLxQYvArTcMTTsMf5gK7m9js6gWQEQD1Sl88RM
1d94++vjvLATGGV+aMwOeBf/4rc+u1kRNVMx/d1e0nHilarFj9ChKqNYCjR1fmhZFy6o9VLdzLlI
jebx/axfwDFsQdSRtVqTbojhilBAHjzicfSyUuhfj6n7Gt3Lx/Xbrx8AsV3eIO44mFKa8fuaew6m
UQ7ysEF88h2PBsJHGDeYtdIVSPUQwDhcWamDoDq3IvuRgVHesO3a9/8TrdNNG5m3yJjx2KRZhv/C
vREs5GtL2zQ/a6BKTfrWMgM4wk2SkILn9m06PiPJoYS5EMSu7yal2i/+NKMAmo413taEYqVVLBGH
GlkQEVdWQJ7kObA6razIupO3pJLOuvSCcuNkNsdKh/ltVnsti5Vrkv31fCZAOeuogDLiAfVIHmHF
ZNvxxCRlly6nZWsh1/CFfpFgtmuKKIkOSqe1wdXAIVwOABi4G6HsYwnNqJpA80w62rSfmFSUtM3e
2ul64OoKzd8kGu2FV8IgQezPG0LZ6gNhKnxtey6JHfXsGhjUWrMxL28dxvaCqgIBhnK749QaviwN
t21GiljX22J/XfL2xVIiiaXn2b96HjYWRYrjInuHNAupTWrWuHBkKTitRsH4YKO5Z8X9VqVZ8deg
tKiQtmzLLTWNpePsi2XoHPbLQ607XkikvhhP/weL17WIJ3K9PcOnxNj2HtDPGet1pyCv5DwdwWdg
BWzv5vYLYc2PJP21Pwr1Kyd+GJ1SXO9lg4Y+cH906R7nhpdf3DIH192/vckjGwQmYlpDPPm9uPFW
WfbGHOwEg0Iy7A1WmuPuMIloueG3/6Dz6nLGNQNKk8TsfpDb08zQffQir1cfgiridbWGAVdYgGP7
FE68+5MkZZ9bO2ngrej8O4CwnJSuYP+DrdvuGMsUmZdC4B8Dz+7s7N5ZB+gQiMg/paz4FfwavF3V
k8ULhZJawWtyPujnv50StVW/097H3cq15zhGKqEo7ApzpFi8RVR/kJKnDb/MXEghBpI/QLQ024cd
UJAsyuBO71hThrKSia5TH07wSTZkcSuGrswC1wv8rOlicCuKHPWKQY8slTyBZeQQBwy+EFxJh5nw
0HXhNH65A0zBy8OQiaxHP1I9ZTN12mC5CTHodg+q9loBA9znj/nQme3aXtBJ2qFst2mz4tpCPGbu
SC3/c5zmhhdj6NWTtF7WqGkHFwfWzrS0W+EZgvLpDlKInEOkVfZ1Q4avUksl49TlfTpAWl5XGLDc
bTAEO0uCWq34urnRudVbC9N0ztf04jg+FKUhgyZSleinZRLx0/Vlj8iFwYp5iZM3dAIELTSbDM4Z
9iJRYIAOZeMaPMMk8utwj3a2dpHM+P8leU+H4i66R6lUCuMFbqVWj+h0nCdhYJvelL6fr5jqQLly
qnf+NRA9othS4QoINSjter+Dhqg7PIHKa2OTOOPfgAyloR21ASIXAsT1zV3o6cFDpgEj1GP323/p
NKdCJil0AkA300pGiZub1jJD+MxTeKHnGUu4hfsZCC/ON/bxNIHTv7D+9O4ny3PPyst89ZFu0iSb
HFZmWPqmmiEICYxLC/TK31HDxXgUHLr2Wcq09O5yv80aHn6L0bwuuEsaiVyiknGFG7JTmE32F+iG
helf5pfgVO58FL9wOG4M+/J1ZjVuiF+Fp5TW2thggcbvVLUPnPN2DBZU4DIPoAvMheBSjX5Xy5PK
85mg/LAjyYRYw5DACL+gr9JTW9aCY9L0cQTLvqVUw/INMnWX54vwX6JrT7ZcRWk+UMysmaYS4y63
2oLkSllAQKCmImUXNgxoMuKXGODv1s0WkEwwKvILqEqUQZr7ZfMbKGu+IwIyfpN5e/0bd4d7B5TG
n56A+tjOS4SY8glRnYsIvKonKKNKczjHnEvYuyKTcvmnIXaBYYLPvg6GKFqdQVX1Fcp9HbUbGvHX
+74vyRGe01BKvv8nlIcwut/9jVGyTCHH3zgABvG1O1Fwx6TX4b6dzuAyDe5WVz6g8g5H1AJnXU6v
JKertx32wKp073vC1WQ2dQvewRwDEePKzw9TqVgdF/xk1iAVGDWnnOuS/puNp05W46lQXQpl/PE0
FMoS2AyYU2rkr03c4dHrfU0XR2hdFK1K0dzAEiO8ZN7rnetVdIRKGBI3TgInbz1Z+lGmeDR0iYJ/
hWVdDAX6QBb4Di7WMj5XgT7KehFyEGcEarPEeQhrjdSBo2bnrOLZyXbTXQwVAQ/aVufIWdCJLPKR
k6eUZVzzMS7oNKcwql2uRcIh7K8QxnCpd4PJxckv61btx6N9Kh+h64U8zLCc8ArAx7sFRv9YG+3Z
aDFetL+kjV+ZtO8lr0Ejg86hNEATZgxaM7ru8PQzo2F/JaYJQzCUkTRn4Crt7+1suagyuwTdz3PO
IXOtY2ztRmyckwwvuKK3X+Z27qyvJ0Y9JETFtLrJeiqhVMIl4xIDl2pZE+x80dncwGY/gh5sJRFs
MuwJ2N1X2dOG9KnRKMzFj05gboIOEWeXRB5bMgY2PVdGuzmdI0SnwqFAGqIlrP3++po7fxnB2JYA
mdodKZcKb23EIkpBxfbQncSAG4WADMKuhfv8XcY6uMgG/ti4TtcwnM9k9jCrBC5BcWE0VoUbk9Qd
ZGrIX2As0KSJF1+CpWxjTxv8wvnBgIqpSTXIljlf1kkUFqVRgNAYJI7ouKCLbyDrLUJNBO5F+w5o
a0a2WlBj4dHDT33FsyYKX+Esvceq6BxwsocSxDggHBRJOMv4IEOxlM6UL6J7zq8TFBInfmD+LyUi
xKWWceIqPxMv/xEeWIK06Osg61550EnohZBSGRoGiCp4PIotr+vX0Mt21K5UleRyhg4HhcUyoeNA
EV6EXgDT10WYIUZrWJ/afac83HDihpJigZteZLcBMZgIe8G35dPzzRTJsuGFVg9VuDVQEDTLVgTM
ePCLoW9HKt3JM8WYWxp86CLe+GSc/F6LkCETliBqkUakp+WxKCPykf0EUf8ylixEggZaK5VaMT3k
M3lBv96YSphl2693lSdXx+4bE2QNEIRmrTWA5EJR/lPSOPccbWqyBrEiVGfCnquDqdVvW2vovp0p
Jotx3vkJFuvxZjC34995cDRPbnNAXsXQ2GsJl/G8xBvqBbknjXbfdyRLh9kHcOFRNaFFcodXh6Gr
X4Ie5OxcHhkANLliPTvNdaf9QwAhkQDqGf5BDkQdcd/jLbvxeorRoTc+rm8fx3E7fkgwwsTEfp/O
3NovSZ5J13tPaavWXAkCvcnhhsqmfg1jiBdHua/H4y3rH6n2L0s7kgOKyeUER/ywtKuZWj1mBSwa
kjbvkaNqMW3fESWcRZdEYKOF8j+VZyRdL5EhF6M3hBND3fhP0gcN3sUUQvVvbFJw4pec8N53XIk5
0wCjt3J6PGtrQ4LvjBSyIJczayakzf8V1JwT/N/KGHwqsamAKDoeGqEbnOteT76DZlqg4GpfaR+B
WyWtygq08GzKXiFNAaYBGdrMNqXRbRk0ct5AsqD/RcG5iAmpd3+DQCUa9vDKzWXtIF0UvWQR+5td
6ButEkM4GiHsVFt3P1D7F3wkoGqv6Y3VEYEu4sJxSueqmMPLCoZK0khpuU8AhKyi+c0AjR8S6E+N
u5IhsHxy3YyjueT2wioKUcLk6ld8fPYQzQo/xl2vlsPmj6l+Vy+n2s6uOFn/4XnC74kJHCdRJUd9
021lzhvYEiTUslDUqBTS7GQfKrmt1tLmM3l2kw2umKPykULCtRByudFIoKlf/WtmM8POS1ROyjFs
xZR9BmX7P1CCCpleA+scGNLPNfF9hL3+sVEKJT7qDvqGs7W0rhpcFh/yDjfI36BGTDe7/TgMNnkq
et9Q6nMZUlmkS3S4/os27PumTHUVASUHSJBFG0AhL09OYNw5rgLC29lR2GqsuuKozmPzbYtDa5fu
0Dg4P+MeyKBseqrYU8VaOVMDKXWMf8gMo2WL26rRqXrVWkfyQuotLp/p0Cy3zExb4B3M41Klj1Wu
MDrkwFpxsHqfq0cs1dhZOchJR5YFO51sd3pGp9JcSuKLvwsubY4dasg4uwglsdGqEdk/CeSrh+cs
QreI7DebZTsgeByI6zna+qb0+sxSq5c2kwO1u7cqINr2QtOy1lFl/tP07Gq4cjUug1XUHrJDw7f+
C2BxrqF7O35/DgoqS7tN/KPEGBImhqa8XBa3aRP99dr7O8t6ybbJDAI+CKTHMCqiwYdGPlExfRQb
Q7KpxwWOh2qAQkfdF048x+aNd0V6M3IjfC4Mevb3nQ43o45eArxcS/RJIEjcZmB1eZYMUxX1N/CE
93ISZGF5+y9KxHF6WBvqWRJkGVtPskjFvxb7IffBUF+tUR8EiCd+zJXKWccHxixum9PEXFwEntOW
dw154r1DLWJreJgT7V5Ia+6nwfcRgFtFsZ30TKaQDG/E+jMNHIADhUWTC4oSIywL3fLx0o/GyOVm
/m6ExlRexZ+vxculIlM/39iHnXeP7fDEPSjPbKVZyAHbJsTzjGL4SFzuhnFQZhSLLsMtnVx+dJM6
ihBtW7pbpsXXpCIGpTwNiWuE7rk/Zmq0XJ1i1Uu1adVVLPpdxHxgtLGY/ahZkrSsl1DDWSydW/B8
R/xtyjhHDFoHkjFt5KbsrGf+cj93Td6li60NJeKRQ1pmhNocQTk1uIx/fIRtXkIusZuierMDKJKZ
sgOzkHkMoQPnwH2eEkVZvySU9TU7IY057nryO8FrEUASvoinRXT7+I1dZt0v5u1MN4YfmUUE4O9d
WYVnxty/G0Trr1qAH6F1qIyTBY4IbyEuf5geQ+ogv67Dl3O4BACJhXHM3cutJCCqAn5IT3QHUZid
m9B45oyFCIoapn18gMgazCVwlJWIxTP3aerb2WPPx89iCD0xFLlEY+4/WVsq/L3Yi7YIzTvBcBl1
+hsdYuNsuD4vTLwmwO9MLYgYoba529PGc1PDAC3ccRFLYykr7PUaYAB5kyo4ba3cEraIf6kPFoRG
tyguZisvECYH4yENivYyh/CZmimGdzxBzlD2fbSSx6fQV82uTyps3abGkZRPJJyBQuIhQrkkeM0W
yWgBYANBIh7qrcwEZrRN4n/o8YYl3uGSD4TCQAg+10cyoS+o6IInlqLqnpS8/jKr2NjOPJPO/6J7
8lqe1QKX2PFRUK8Vfpi0b/5gz4hEWDsPhsuRI7EWmG+Oqz/1CzeSikmwpd5qLchtCRsjCL2uugjT
ojvDC0pcqe3FzH8mGqo21+8odKlfMSFFGzVST1POVjZE6R7QG0EdO0fYQ6F+8rsuT7bCZA+umr2R
PBrDfdaFOZzPumtojIiOOjFHJETSwWqSYENaITjNUMxk9T8AikNeKfFjWb5jhCRXpyBMPSeWXYXY
bNifYVjte3FWC9PXTw58l7PAwmUqtp8NDeb6zaPYWgRrnlnwq9Xv84AZsLxhGJ7pn8BUrY59d7Ar
n7CJnarSH+8L13w/2D4BXq9LduRQ24F1fqzuY/go2WFFaT+sf5yVcxQORWUkyOBD4nPYdTPLm0mb
hV1T8oJeXUe5kK6gwoC+aOCf7/k7I+pRxFvaHtNJvuEcowdtGkbBAGaRDPf/2UIkBW8tg5sqmr1t
k0472lDYO4bWsZGSgoMN9h7J3BOhksHgGOqI+98EibCCohuPKjNgxLzCO0aCe0y9YqeUjF4ddQhg
DL31vgatPq2OEsJcGFZstA8RtBli3fFrAbRAi8NgPtVp1auh2TeThgWzHIBLB0FFC9eqVYYjU3A8
iCmUMl6Q1BBN8Kt6wgGufZNML+ysRIFRpJ78F7rBGUuWs+zbAy+DLbS7W+SE2ShIJj32vVZ0oITb
sCLFlfd+Cf6AYyQKE14WNHOZymY1GHi/JTDyaQeTQNwO2ReHwSdzMZXFoeoZEBBpv/f+99l4zJo8
RXp/ysNSN8q1LlOD752mRlWht08O2ZP0nu5qZLN9uHqXRiwRCCGmca6udP0gzv5Xc1jtV+4bfiPs
XJgKaH47QjwLBuNXuDyk6a4Li/mqPYRtSdalcDX1ZfiEKo7kQBrNTfXtmlqB22f681VT6KwWLUi+
ZDU9zeBLOhbwMogvOY7oaCsED7aI6fQRDx674ZkiIsZxx8NVer3lHzi1YH9FEKdiG8r4gXS3p8Jc
Mg7hDR/yWPook1+yyyFShVVMArC7hudcD/y3GibwdrxYrRNiBCoDDNckT634V4wBmEWF5Pd5pI3y
bVnX4APFzaVmB/sKXlEOfPFUiWto0ysVb7SJTB6rDyjJDpekTtQ+04MuQJ4dO1EnYbLv8BzDIVxW
le/QJQ5YQ1t/H7GkYwbeaGcU2jKNB4uVT6tf7zznwUPW/mK+rVM91pt9UnJoqcUvVZSg1+5owqrQ
xqZN8fq3YAKke2qyek+tr2HS9gkYQwwq8zYhmc/NjkbvLPmMTCAfWEbJHq9OwptVucqZHINgMuwo
6JH7B5JvbhOf+fxTTh3XYbQ/casACv+au/ZwWzNruHsodq80YPDg+uYAqY6lUH3ckqfMrMQA+/mt
zblmI7ab72Lt996/NBVmwhWBg5lrM/h1iNCn1Fo3S2CsFhOPUJw3AZ7oj9bWvYi+XlOJzj/EgyY7
IUtyYkxpTBylGglqv2/EVEZ19DSWQI1SINV5OXRbNf94s4gOb+F//tdO38LiiQ4Mi/HV2Pix86kg
WRP3vQkWqWEoUmHzRraCRs81Pwu3V740fQCqR5Yp8z++BG4pBA26y0b17PA36nnW3+D0FrosRmfU
KmAY4D7Y6uk53muOGY5aCFKNUE24bCcozy2K/Jjk+ry1jLVD65Yo2GHfBSbbpeNzqTcJaOHeIe0q
7G+/ez33W9uFrP7Ztk0O2J8I2Ru1Fp5OdwzJD4Njy4yvB+Zi47kbfCXHSxIWrvPNNUW/ExHk26yN
hGo6w9Ub3nTa41Denj2VuHSIaK+RcbNwETx8HEcN/pFsIU9Jj5QqMv1VreE7fzAWIrbPeeCBobXg
dCfHGSEHAqdCh9VztD3oeP8GvoQ2WTKtL2IuK3Rw2zaoVomfpV9e6xgq+hmAhjxSUAqZnJVtg92B
/shM6Aeck+AAYPBY0rDAxW29FpR38bcsLExfHOwR/q1TMc7KLH0qNdaaC65qHogQjHbMAxRwJP/E
guVjZj/KwKJiwj6IJd4fWbAtFDnxX0fJLcpZiBSwKr8Zc2fLl7Pg1+VBeEs10+xFc4MdEeqUw8Xy
3gHIK1UvN77Pxi+ffv3sRn6GrQjAumE+36lmnzUCEZWV4ux4Jd5QogHl9OIxYRsBECLGedk/nSjx
pi8Q6qVQbDy1JoZAuAFowcvQeoFc2fmoxiez9YsB9tTvXf0WZhwlXGcWwD+CrMqtnb113BmgJ1TP
pzL1OqRk5tnwcnFIxMCBJXt8lq4o7gM2kt7OGif2X8nZ1KpNCxQxe+NuYBfIS4BuJcmTAyYIqn0V
F9aLUkTtp4Ix9CWPde03x0vpT21gKGhE+5WDOQ5SVpvzBjR3HvY8+auTZZwPqYcgiRhmLS/shVns
10oITD5sT+C6+T5o14r2YM/bHVnY1mXl0ZjRCEI7QzH0kD80Qj+XoZ6OHluXOwb9Uar81dcSp5eb
ak8CoeHd0TBmmiAwioZL2Qd+LLdwRd+2T/NlIM5OUV6QqwhR8bXAQcJWtCyi9FqxGFJsSzjZkyLO
R6Iu0hrnvI86uIkAxqWbWE9qByMrLD6eNzPEtQAcSPCBsh1rqh57HMoEftiQGflOoXkSsIYEoUze
a9zy4IulFKHHcTCAI2yLY9n27u9yLMX70bb43F+yYqfXc6pePA0tl6yz6+kjMojdEkAcfa9lsFZn
aXnUphWMzsQPfThPJ/1hG9j3gmDuatGn+vXLXPQOQIMiuZthCrzAwFOsOiBRXjkskcK+/OpsbBg/
dXyT1k3X/yxxIdFKfkY87MWHDYsiSp+Nxx6fQxWR+yLxW4UUVnpQERjAISyNeHdrBFpCGx8VGE1E
NVzRU5PfwooG93XGsDPQIIlxlZ56Vk7BscjW4OrS06FZCbIQ2oz0MG4wiHZMWLR93HmVzYkjVd3S
uLdWpU58T5f587XmPH/PusbVrVnXUGCX/8q9LOTOPu84sqKbEkyfYloGy4LFuTSGsyMFat7ANkxw
RibVHqAvwJuMRPRpt/n7e7ftFas5TrWKVNLO8xwnY1EsPEiGE/uDr5A0CsKgrQDUh1iuxAXESZwg
EJDYGWE+zGS9p9DOiJHttAO9PnYQs/f3b9FTlct4XlOqgWehyn7quOc0I9DEQFiN1bErGBa7RO2t
Ax/NYLUVJ4gWDzHlr1CteK5Io5hWvKgQ9AXpacJvUbcqDHis1eJocfqNec5WJ3N6iehNY4h39nTt
/vWIMuFZAQEfH9E3ofMPgk8prF0DySa6FKu+rKeCxN3drVuhOIYX/cTAKI+tSS4++HXeuJCBKURR
xkZYua9vDStFDsUuRCyOQMPq1ABVxgo1FzDmDVMlC5aHVeYxnDfjeilB5HI6rEChTZb51ozi4juw
cpM+p+m79LkA0KiUScx8Ki9b0J40TroWRu35tsD2YJMshkFGhm5tUhozfJHoMorTzGsqeW3KE+Hm
VFbnUV7yJSi1Rsv6CL4RjHXOucNUkDvkzt9+NslbjuEqODw9FlYrGbq5Qz9Wq1qquXXsUfWX+wJB
y2yC4ROu6wpOKpy5agAC8xgGJaUk8JqTfKFcwM6k95pswSFug5gjAa95wvzHs9eTRXhjtls1oRMK
Y7xNhSw5D13V2DqGd4Q5bRlU9P3DNBn/fYmR9gqcePVTEMu5EfzoWnxPdczMFowOU8CR5p3up+8g
XbAljG+CC6ghDnZOktgXU8DQz2Vkqi31xzxoY5BAwmGe+qzlUUP2xsRpTr5E2LEuuxjjWZCatqnq
lQKcrJhMdvGdwxFg6R/zRUI+osVuwSmvlkV74J1E5/RgXhVIgJB8LUWOzedojHBAb/AeJy6dWMEu
v8EO+7C4OA0ZMw91tyHpiDasKtKBDiO35J3wp4RQSP2C8ZONDfokzPh9MSmlcfAhwfwgN7gQ3iVg
NEmpxx6ccKzR30lR+mo/pHn5LQrrV1m6lgQ8kMOrVH8+Sl23p1ZByWMAlXFkZ0KYtR2Q9G5qHSB5
0e0Kq/y0wqiTIMjaGn/j9pO1yU/XAYUX9AI6+0ZoKUyGgmC74PErg0iNnx18bbWlOBYaqybzIAdE
3BPiIGUNLCQxmNlMZZ1xSUQzb6l/HMgET+hSGVgeBfGmgmHuxW69LaegKEkAKzqXjbiR3dv6Dbko
e9jI3b3DUXqNOxDgJ33G2Sn1gxy5yTOgmrx2lyVZiXaulf1xITsnt0Cbx6wIwjCdvdoYxi18OHGF
ELCvART5JpCbD8L6oJj6eliTeSTcbMiwDC9p6dpaRYjJtBw0OUhZxtgnhtk6dmWJ8CqG20eAJX25
G48uGFiTLT+9TIqTIBSrW1UPG2EpbT1mOLwyli2DbxkAbAEgtl5yG/rRLLWvryWG+XMJ0Ln0j38f
bvxD32qE8WgMlKT0N3+ZAIzJmBXp1RmIxozr3vhKtffk3tIftR4GWoff+V+soLRWIdrSSHVYuNTy
DuBmOwn0B/+flZSzOjxRwntA3Ify9tsKN70RfOFMC+6aNA73IQo4zBbS+VHkZ2yMnfgiRqD8rtU7
0x3ozdvCqW0W9Lcf8TuiJij9Dm6Ock126o5fwdd/2+JQvpEGGorOOkyMskGp/U06leSmAgaJspXx
3uiqLtCL0QdJ5QzzMk2CTCB4dUQ8XW2srdxVOPA24AGbf5ktr7Luq8s+Su7ZyZTuw/HDIMhHSArO
xG8KekxQAm2utM047rqT1U5mLwY5nZXvygg1WquvjvvcmwxhrYlYZCDrkKaitT6F/8X8wxQSit8Z
cN0eU/XgXXDavM0iKn8QZcQdKVkggFqj4ApJQYqpfPYQ8m4fegzfmqYcJL2vbnDUXUNv75R1ONCt
TPikCsVl7a94mECQ8P4wdsevFSF72Eg3qRbHHs2NFnOs64e389FPI/v7zq3Rl39cry/gqDgonF3l
NWuE/2TmJBOG38An73ilFugToVAxeTYNRB2danDX2/zNDUPxr3PaxKxOmq2obv5YVSmq8N92AXkI
t3XvikRKH3pVaE5iTvj0yQQXSJsRmwkyclqBFLVYYNxkyuu9xAhhpIL63e2wOguaPm0yQtEZ8+jI
qF1VCqvUPDOziGrSNBPnUO4eMYQE7/wKKXRmGPpPxrWnwKbPpuUaq0Fz4f+xO86FjLo/jhxJ98VM
W4bKer2rngvu+YBGbjoZ/D4VuR+ziMxej2jet2aIkn4fDxIvLtT45KwHjmOO5JPff5WYT+WUMG9W
0LhUgEnowXJ4dKfIJITFB/ldaDB3XpfVb6UjT/djluetIGeS7OIEOphFuydyBpBxRVV9XbGoY5ea
Pvt0nfkcr93kZvYlPHD9/fWuxrPocAhOr/m+ONF74Sl/Rs2yZyKkPzozBAELXaDq+NqWj8qhmIn9
Z5XtnY54t6djtV6gc0fZKQg88J5QwRj1wMBtnhOvQzyyPAbTRYc9wan9YtufKlY15IO3hfGfR2m/
wuhXV34gC2DuTOeVZfkP3ihRYGYgN70Ff+GnCpdtHIkffa8w4HPXjdbYLCRgvAzvrxUXAT9Vbimx
htakmRw3PMihiahxS/sc7uUSljMg9wtOZ2+fQCi3JhGoj7knHN8ueQ33j2Q8Z2F5d/sIlXomMC5H
g1S9xaX7RfMSAMc0vDEcp7lwNCnHkJ2PaEXz85Jo3y7CZRgfxSeNtN0pyusC9rBM8Jl0A1lBjtI7
TuWML/b5Qkziell90oUhSsMcI59gTolSvkXHMkFzHW6xTCrm7/xE9oRtmloL6Cf/QCHarAbl1eUQ
hRir7bLRe/ANkt0sPZuMEVl7MwqIcM0rtVUtq+pNZEnUaJPnuGJ6KD5xqC9ZI1BFO64zOO1c0gAi
fG8ZxmPlnrw/hRRDLi6Kd60RNPEU8x081CWwAvKl7CTQE7FfLpRk3YbMpvs1VpmbWksolDc2QVZW
aPgha2hG+PDjae6XyJgkgwaR/7LB5daDVzVJMJjo+6yIRJKZust+ABo/EQAbP/FcJyBuSeJ8KdMY
k+MiAiKDZsCo7aSMcYxokKGtB4Kf+WeJjDp5IRSas68/Qj27FlbZVC/Yxdr6h3GdI+fGQvXoO7fu
paa46s2o0bnzy0DzfNnMDAQ4+zwkKJ8J3Cpidydm7ge66Wxku+4NLX+EID6dim0HTprtnZSRxS0F
sD235WOMAmvGWdfEo3mX8J0oXixiti51REsH/xVU25bVKhftYGw8D68vPaB/X/pQP0hNijmkZv9E
oE8VbxcD61KzZ1OOhNfVrYG4guIOXNzvT6ab1M2sKx1Xj4k+JFEyzFMe1F5mowOOliIivfFz+/ew
oRfbHOfa44Cd2O8OwwqqyUcQfET+eSrzFD5RyzNeHQqVVyTptPrakLuM9x7ln9rTfjlW+b9WfZx1
1trxwdZZA790yFo+4t+hpXuX2RF2U+pmWNHAqBXHjh2gbumUpHfAMfhH2RGj/I8FHG+Z+fBwy7Hz
4NAIsqPNpaTcWXxtg27ilSWhX0ovTZWM1qR8CQXl2ZFhyHntPdsJdkOp2MfnTpT2r/jIA95k2lXG
j21Olbc5xlPm2auP36pi/5+H2Yd+n1khwjMfrt0zqCjw/LlVyqXCJ31l8zHeo/HPVQtfjs0+MkfQ
jPHxiWH7CtksiaB5pFf+ZnZmW/jHXVdVl6LRhiQEV19jIKArAFK1YFI6tJuRvSUnxOszFXUhIVrI
ox/WDAfPDIw1PM/t2YOA2Dtx/EnitULGnCOW9NVUTOlDHO2vSZLPuPEtKQXJiht/9GNqlh+09ZP0
F8bgA3uVSiD2dRqmAAzGD+gE81CwCMbSrn5TjNM+6gf+H9fmzGwOqJysFikrPXlOSpkdHSXip76p
orkPc3+4KmXftJpIs4X/wGZrcRdV+jTEdDzX3m8Tm2LNYw3AhpUKy3Jnw8KITIVSWFnyhXoAGZVA
7Vdl6SX7eG6lTdWQKg5DFpuAdM8a37LbYG4WjY27hG642HndEf0N7gtcH93cMNEcwhMPg6pLRo/+
V5/4CI6hUio0v+/wi2XZ9pmIydyfvOPypMdv3iBdvTJ9byszFN7/4Bq4jv8dPBFM+qgK8wuAhH6f
o+fzIg6bBeCXBpXqoryQ5Jbpwo8GjA7KyQ8Em3q71nt+33KmxeuBj9r+TEdxR9UjEE9a3hSs83yx
6ryaT+LKOzEEo3PdSf9tc30g6hYpDdX1m7fyVuktWRIsEtyGQb7u/O9qPavO/LJASZZu15Kxi5iv
Dqx3kXVDYJUnalbBBDFRQvZNw0toxVza+eyRjH5N98go/S/keuNSogqAXkjSeP2OOyQtLypRl0y4
Y/PBoznlzEEblUBjSFdmI9KUENGFcPxjzE+zExpNKKR3GNtbwAhpgnQ7P+xvdA8hP3CYTTy3WKds
Vb7c8PqtVZHnNis+eQlcHHBY6u4TGTAogzt3ZWAleT71d+JPTfOhqn5AQHD18AcDWGXgAnhQUhNL
FVVTFMj8LWA3STYlCN5Lyz/SYXoXDLfTN4k7Atr6qaFp5meFVc02etIIN6pANfLXHlKzq7eX3cyS
pgyL9dlyzO9U7EMgoxSn5XLH83ZStE+mRvx/x+8BM4ER/lQpyhUeqLhKMLWq8xU9GT/JRmi6Z5FJ
L4WsxBrRi8PV3/J58CcO8p7qsCXeCWe7Ho73txiHKtjsHzKl1X3rJNJXYeeQ/KRJqDXLeoT6LxLn
3iivbURLtXiVXev0CHPafaQ9b22iuPkNOecAL3tAxbQElN7PBeyJVoL++o+FY7AZQjy8xZeLoit6
TshphnVFNeUg4yoz2oNE77qTuxxd8RDd3oD7TQN+F0qMyIdcCBGuak86WpIqFWhP6qYX/VpPk0YJ
SMm2u7ls7Ez4Pb8eUb8AV+IBhpaoqjm9PzmRo3VI/G6XA89jbNNVa54pMVLdELEhM/YUQdr7RCUV
vR6gbN85VNYz5TIZZoBFhtq8ZkcY5PNsJR8ewZiVDql5aczTlh/wMluoMuU8P5LWN1J0YSs8KwSk
7Z3fsyWp9fWaIAdM0zmq69doLQSI5UBPqEDAb19eEIf6jYw1LzSkhQg+vuIlY130J7jUplDF7hKX
aMLpzHEL8SNdYzfgOTOn/Ew6BmLV2GIecszZG6PX42ZLLm3547dcK0kBmZs1neFBcmjix/QWGxsN
VCdPEqXg6uvw4eHbSeVrRC/DSNLbnVLoIhYhPShkRsxmgZq9RkK8iSBdjaqezS+in5OBaqrsTCOZ
pi84ZbUBljce1HPSg3XfzXIvDNtTc7qgMvl5ayvIQyPv6SK2OCl53unF7DY8gQgoxJhO4s6+jn7i
3z+PVbKm6SreQdEEwq9OTaXqCqNTqh7B/MVqojd+wGjaFldvW+23JhN7eaaSYC2pOI/jgbDnUl2O
o/BYM5O3Ip0bxwdWou4CHTff4HA1VN/sR2WzkVHyDMQ1+KJd0DeOB5BWu9EO4/JNhT/FFgfTNUK+
RHuKOKF1fH9RyUpuyO+RgRckwytiaRIg43v4GFRXIuXDQd/lAWyk9gnm/PLmPcAtkploFByndJwk
yIlO8OFvzmreloAldFQ+JDsOeoCThwTdp829/qYAxGu9Dquz3/ValThTp+R95e6PZPGT7Xw7yxZB
qy1vl64BeRagMFXAaxDYvc/HC3fhc1WK0MhwihwNcA5KGIzFV3GVrBv4cjn3CAWgXajr0ttni2/s
2YCPXx7bhMLB6JxvMouwnZmmX73s9SsyiOWKhIg6cC+YsCCVEPq6sU0RCd6zIyxRJtupfpyEeYVH
eZkRCtnhoMdq6Tbq5Z7pva7AOooPSUBGNSsL2EfmMnks8LcPU4kyqO6d71iJbT+4v80otuosWVlF
S07rrYRG1mbat2OeS2+Q79ihS5uXYbvnE8xJfVyZnlNm8/dCT+24py1KqA/GgSHvR9f5TYODYiMo
V4q0mqZAbD1cpcJJfgJZhWBIb4yLpaMTsLk924jhAY2C1GPP8krAFYkLzxBcuyBVxfRVr65ZFvVE
ea+4es6WLJyDe3zx/Ej2nbazr5hX6K2JEFf5URu+SaphNHlyCohT4ceQwaDTBR2X0+OZhGbGDYMF
cqSNdCjunOx406ibFdJrr9atJX7ICmG/TmTMSXWXk/jbqPZ9bTXbRgCeYjV6VwBl/8V5e6m9uEyp
5Mhz/DpFfBfUk4b4ADRuC18InES47xHqwLaO2iVKxhKuYn9bQFOD39eZ9R2Z/Nckfp1/ooY5coFB
J1CIcXYU32y3Xfxn0mcO0D5fiZ+IPvF4m7hRX30EdYnbbePQilTJU2njmX/YFCdFBqT8yriAwOc1
frcqYzOQJyWtHHTSj2JRvt+CHCpVBtkmnkB7wNwbyrDMEIs/3V/b2iM5YycODAo4ttoaV3J3k2gc
qyqUXNT8QZ+oRQauttZZ6lAXJVRrY3FBnltUmE9v2K48koqFjhp5Lwd0Y8hctqM8ycsWX5xGrnhL
YoBtkyhuzDcNIaUbwbe0VRCKb1TFhE4B/DzvCIKN2wZxWjLf6zsAb24r/8fIgEkU3/LRc3OazOX1
ll8Z6FEsJFvm8f/1ly0vN+O9vTUJLmyzV8CGLrQqESJ2R34jPW2YOBgWhiEFvCNNXQtBCb4Uk+KY
dx+2b24AgQ0I+sy3UF6G929EGCAPWZothkNIXJRPYdwLDQuf4UPMWEPVkC4zodP3ty5/Kai/fyVe
qdO2HpKcavf946Ga3aMHzqLVLYqVlq6VC5qCdUusVv5+yzWVOC1Zy5P8phMJZMMWq1VGDgjFkHbo
9P0UCrcKNrhPI78FGzz+0gBpJ54AGr5lCuPStD8OeXztttfKE3As+SLyFgkOOyRCkUghKS5d2dEk
hgSkA6cZElZjAbydMShl1s+qJcUyfELunmmzErwv+VYXVa/k+nqnhBz8VkVcvjjl+jgQMbb1nn/6
AzL0Vjydgw7Ln11zFZQf52BItrv5eDq4iDTtE9l7nTHS5H/gjWrgtZ7njOliSd+DfDfd8CosNJH3
bF+A47eQHnFRRekETyoNAMfaCSja2VM2oDQsMkHz9wDRtpkJe5TXK72EvPAc9bDCBvyeTNjt/MqA
MzoiwVJAGSpG7qTawF34lJxhKejqDguJ0qUEzSKb+R9V6kWqUF+6MwRGekVnE0YXtuuxlBHQ3yYf
+3zuM9RrGCmgvW0fXT/HkG2RUmHGabl7CjFJEqGPBfXAFdtxuXj7KqPxj2O3B1FnvdUWL581E2cH
CrQO5G0Exo4XHyl0uZUCCWgtEzgA3MYaF8v9QPV4ZfRGhwBI+coS2uXWe9H5wufIR363wlEmeQQd
leqGX5FPasjyDWA5A+bYYIkrkQZvVBgBWj/sbMgPLAV+wGRPWcnSiRQPlUTubtiFwNgUFLGvp3H7
vZdEXJngjt+kPkSgRzruII2uznqdBl31598buYCleH4a0Ag5GciTl3tTQGclP/QWuILJkreHZ3UW
8Gmo+v5qTyakkkwnsOTCMsLf3uU0SlOO1AdqLfyXBU1upIYSNbi3coYWL3dWyAbY/wunNH+7TCqz
yJZ+dO6SxngvdsDG9Eq8BCJmNVcayeEVEEuT4W6BjjSktsrY9diR3C1Bug7frMNcfpUPvV35Sh8Q
81Js07sLbJDbTMFTeJqR+hDwGI9dBHS5CavpD4i5cbqrMRLghXbaVwW7wzY5qHDhYbn8K582dQBq
HFQo1YokhpEGK/KcFEV1smHa1Xumf2jmCN789i4Qkn/RnRTPjeZlh9jtYWbWfoE+4/iiS3SCApZf
q1cD+3BqIp4jmDDf0c5kp5mDzm8ysfRbwybehrHw1C99IONS8djw4RFQbopZ/Np3hJ8dbjFXqtTb
2nj8ve8tDbf9a3SNAHrj3LlMNUT0I1GOvFB70l5eKTb48Zcsk7U8hkj031Wa+K+pG2jN2Pgm06vW
hIHOdvTTTXndxMiscgelpMHb8ccp9rX5elj/1AtqMa30lGxSF7FFoA2Objm5j2ZXSWhukOSedqnG
7j7OfL2+F5tfKkLRnhR0zxmWrLzmTak+G/5ZkEVu1lgOrdfb8r6jUQOStFpOFFCWxiHlfylWLTaC
GoJMs7+Z0Uw30swJ/qtzcJl0wDMiWzqjPN8Bh35jVQHYhZNSSmiBJFPAKr4lfAJbZGLMZfqcPnfh
FZgKNNba6Zq11TvNHtbogvuFlKc/VIkVP7B6lsERhLJgAbmZA1EJsJ+eCC5xdFKmUrx3Aqmv8bpc
t+bEPjp08NSlL3mbITGx1dKrgPEHB2sh8k0I0AyYvpBk6dD45cyU+zPBw23hxQLeYGQyIQL2CjpZ
m7d+ufOJPK1ll4eEyXxpwYK4RZfZ+6m+V9x+FX8cKnSMtR9Z/Z4F31lQhZNxrvjgk5n9+QV+EXkK
N2FCux/s92TLZklJBEJ/DKmWkmN040Ej/K6nIuSgrcg5Wsbi7/BwPyA/6BXSieEQvHOxVqV6GIqh
xnpbz4Ktg8QXEILolXEGWxxRyJX2qIUQsfKUiJUt/nPkOhgfdzifyaRxhwBMHCuRfbBJwRRg8GDJ
m1og8tseVcZujQj+k9Tlm18QnL/2v0Bnau1jij+43LdNbJe32ZWZqePFzAgr8mmJprUhJBwabn9y
MK+I+AEjiEWoxSrS6N7S/Ku9wn/TFCe4SddQxo/LWcEfXfYf/Rw5IN+4CzGpxXvoE7n/oR+Nwel2
VVcTf/8KGvDBao32G8rgXxUU5Sis0S7F/i3UjHMXNp2gSQyDsmggNKABKDwtuZK+fDmJQSFsbwsB
UsCDfHqZOk/bn1YUdCAMhyRET0SUoUWchNyQ2XZ/ZwRiHArS1t3xKshC6lx9lz2nk623x+fs2QjS
ndopk02IK48SfQmTtbWBJTvc8WYRX9yG34VfeAiYdqsbmLknoSp9+uDHFEvBe7Hdy1HFDOTPqeCA
eQXE2i2lA+/7uFr2M0SFQfTwHyZR/fG05uc0GaXQ21QAzkZu5wOEgxAdJ26QMuVJ4B1f2JbzzgXX
hb6Dp+7VVCOYN7JZtDHiqVqmPYJA3kzkAm1V/x2ts4vjWRfrUUkO7D8InZy+eHg0Zvizd5Sf+4SP
zFvmcXrNO4x1XvWg1liGNWet9dQwHjXw8/Eu/KSWjXOvgmxv1a3dalX9Ogwuv8rs9w27EWLQKWYy
Pp5oBDS5WS0RFvhx2p2BeKzHN3jWiPU3if50Gm439GNSGb+jMsbXH//uMuG+iZR8lO//XkxUa5ce
EMXQrk8aiCRn0EEst7cBJwCG8GULPc2YaaQYyoOe3Bv7cCXhDPdIKuQcVAWh0v0/jWWeQSglF0aS
4dZp7t4cbehrLKysdEy1bZOcxiBCtnTkFWTpJ5wL2CYQJn1Mbi/WENbhXFv+vnK3CgMdpoZ6cqJY
zgbIIn2oDERrTVk9Vtw6d4qfShdo79wNtt+d2RXKiz4syoUhgJskl6bIo6mBBCjVnSQzLPN8tnnF
9krPxGW3Mw5zXRxK8htDCpxXHxYVxy7fIjFVZsBrAXtLTbogAqfQwM66inVJt+mnrIBt5pJSJOpP
mW4t/Fs0aC2nNafBfNCfOitMwZZz3S1nCN6J2OGmScXAUIxdyZrzkULk5wJpD9/VjCnWFRNS9mqH
4y7fgvxIg2+kJs5KCeM80LaGLoTQSiupiiKo55WwjYX7FY+vNlLB9ZIngQVzQKtWIKXO4rIdYgmW
QnCRhjjAym327qfAoqelCX4fi5YPCFATYUYtyS49YWJMmtRDE1I+aNsdEF/dAamEnE0oG8jirUeX
ImF20OLImfbPxqLGT9v9PXPVPiQ7GE7xx4p86AN8bh+vY3pwYlJyBRRwr7QJMi/xujSYHn+l9N0k
3CmV65/bB5r74USeQD6sjeElLJelTl5VGfgX+JZhpffM2GGGX2/4Zz8Egq2CRjco3qdht8Fl5wvl
zSdzlIrQwQexc/7Pxag42LQ1gC8BX7eQcuz8rHERxNc7sfa/0eKQnJUV0+/9hI6gZJnNnBFlWLlk
qqjnwWPP7cCtzmF8G1hAxGXeWy98FZWcQ6hSlJPnZnbxyHa6erP9c/guDJ9s0Of5zd3tJ2HOk6BF
Y3+MJrTbCh136PUlTkN2qHgLRSInOkwLxNNaeGdtk8iQCJIbWwkF40pR6U4rlZBHJaWqx0uC89D/
UcFMkl9ZZbhiV8WP5/5G0QFGk3MkltGtlPeVnGSCIpGLbxk5JbstAZGoZPbJeXa2EoCzUjvUmcma
tbDXd3Rji7pnCzB+S7dCmJ7DUlkkvqX3Vr5eiNL98kgeWEJsWHgafbYaSzu3MhQAV4k7yF+AGhu1
1ggYfMVQtASYQ1B8ZPjXV3ygOmaNs41cv2vjZADM2jJ1VlCxRzhgd/AhvB8QIV++Q2oYuOLUEMRj
XUOfxYtoU8CYpLJ6CV5g3rRgw5wVdhUa02jsbfvT1Cte6Z2fXRfrdBS+KFKX40UykLgqBjxlrW3g
gqvI+1w7Pxz6Oo0XlRCw2Fx7wBVJKdze5RSQdCx2dugF6xCseHL2KicdjN+gKvkO/SuyNRaPn0Ru
UgzJE9ToFQ9FXfatHUBwutqurKt8uyPfyy9fzmLtG6FhU69cpNF7Y11Vw/6veBptm3AJbp13BYc9
i3GMqUme+pZPzSMT1W+q/KlibWxn//5ZbiA/B+OFAyJZaeMLzKDdCJQroRFUG5gZfcj9AZ5sJ46D
c4fxt2ZQbOO3Ft+fvUj2r5JC1lDhjb33qxHRRcmPgEDtvhJL344Zmy3pI0BCbPFwhedIj8/ANeFs
qR5433COu4JVMwxNMXPaVgAM/279Of3utMHkIdEkbzFmACfHZu2Y3TP2crJSrcibTEwrKItc7YSO
dsBu84DbD/yLUHOlMpl9xQ8R+rySKvAfoYTLRk1KQvwbxjHZj9lUL2w8qgheMXG/5NOHFyKbNfXS
njPHfMbGL7LhcCIlvXaQJj7i7ubLxpkkh4DzWInRmD5xVSMa2VaM0XC7exM9IBiRRRiPi2StiCLK
fGptlBSW9W/OqnXrJyozHvvwsM4tYlsOj7mU4heP8Zaj0ljMBsONu0tFxPJn6p39EZLYzW13uT5T
6eQi79sEfNJm8yz6vAkmReffk3LJje5hNpeYt044jLpkLkkr5mLsRUS5wHpCRAhdFwcbWPTOJCAC
qB+EbMlVFtB1xMa4rzCny3U7UCp/7weEkfLo1s7kVq/AT5cUCRBblTg3OiN+mDStHwhJS4jdO01+
IUoL6Lgm5mTjwcLvLdiFRPgF4IfJv6nf20WVsSsxHYbbaHuUVZblCM2xi8mM+PLRA+2nR/0hxA71
BKFzZUE/0yN6nllnmHGYmTiaB0oGozTs5ydfT562hAMmLVKYYxnTgX+Z+Cuzv0/P6fJbTkB2ZFx3
IkhCEtlWWj2d48qwCa7iwuMnhi625EQMhDXW3xWZ1WDbbU19sIgxxpARmIYTubdxyZbJ8Rzoa+EG
6FCmjaLbJ2kmGlIgD2RAtul/0mSdCzRokYFr9ge8abu9UyHBX5kTJmDwUhLZHIY9oe73v5oamVS9
1noOOv1Jq+etLrQBnT60UwBVk9XxbpUQUDdRBWZXIwxEISArtPokYNAVEbjCSSe/1hD09ifhkUGX
mtuJl1dxq6ObtyvxloROioe0f90OYzAU48Nd1YrxlxHZp3nQ7MZIWoufafhScrHru954KJ8UKDFw
tNAxhKiARSNaRKsHnuqmrg+ZWW6gsnxEHlMpA+mUNdWuCPDa/s4DHGY2BUEyy1Zf4o81Jgy1L61x
XsqVo7xoYyP2EN6Vz+qOZfIk+5oMQ1SeR43zkahzzO1aTqwktsfZkLRAobA2/CClqzm3wm4D0q+O
c3/YA9aIE+86JkakmgsYYpTj/Kknk+O4zfmn3ivW4zpxAriasWurysEtjJvHg9w/J543NeGflyM8
ji6iDzMT1FD5zbIe1gSzYFW/crL3oXQNMda+pPsGXbsZBa/cOyav959aaRMPUEirHijQqtP1qpTU
U4I9kVtHuNPze6fFrCcfrvGGR0I/AM7/Fep98k8NxQUrVjgnkDAIFqWHLPTp9TAyel2SbhnYapKs
/1H/kU2ozi3VHiHyKgToTz8gTb7vzNvoAMP0QeTIS41Rmzm3U5+YZDfNz1aK4V5QKph5wgSdxRKc
p33kIqz+MeHrgXzNr1KgZyx0wNVDnsrj3Jlc6KvbNvP/W9Nlgr+lwttwZPned7H7ve4vHdUrvaq2
nja+stu7t/nt+/Ol8+h4VHlyWcMai2iSXK97G4naK7tMw3x9mFxw3opvbdz9WKrd2B/5kzgRj6QG
diIztQ9g9b8qnfBOEh4IiV5LepzXpqqivHzjju4moDuWU4tPbFbXSVIa/YRk0VMVZ4FbphjlL6Aa
YM7ftyFaXiYtfBh9HU5Kwm6IyPbR04xeK6SCNUCz+kHIgO2dbpOf6A51q9f6vLRRukPjFy//vd7F
g03zxebtd8u17cvIsle/k1CIsZUCBD9dxKKGg8/WJ1wawN+6ZDr2Wax+0dxcn1z+JSFNTUmuBphc
GrhhFnJEGFm2YpwXp2yUI2xM1GWmc0zVRi6C4faKTPpuLEVzOeoHxQ1Ioy3g6D6NJvsBEgdKJmL7
i/by4npypdsJLDHWdgyk0WNEeHe2Ms1YlDgtanI7D2H07hVg4yCVr8bmLczG1vQ063/dfoPebn/6
XpMTV3GMaJY3IWrEczOYNpCYHgx5RVZ28n5w80+NsaAKCQLzXiyKQ8oDm/6K1bYWQzgGNzO4Cw5y
HiGXAkMe1eafoNkFkLczqcTSQZIQBA/W+IqWKmSdufIRbH0MfUF2tdA6OebeOmJGPjE6T3isTTWK
D5G8PFzuWuYNJedl80Mk2YKraityir7McehUL0fW6p6wy8Ha6T73d7xzSCduVpTswxyVzvXdt+so
uLpO/lyAxHF90SfSnatJdbg0lgYJ55PJJao13bExoautaXIqXBZQhDbFCoCWCLKsz31zxacdJi8+
ua1RC8I8DA19hx/nmBGnfeEtd/WBIajcWRI+AGj9i44qe/6V6vcZTHoMrAMenxzbwG0sQlKFgrf0
sVI1jYApo+9GSogWuS0F1rpvwWMSDf3UWvzXV6Wt9j4hFuwdkdOEK7WfUmramEnJ0krPPTwlhmdH
LZZst70tGAME+D54l0FBlqVqeXYXsXbi85s3iiqNsuZTPCpu+tATNOfuOIk64ZBIrVqz6RMP33E8
I7mg+HLXQPihvJVnVgRUqANKNQ17KpP/SZRF1TnstEERSovd23WPZZ54iQCG3jQqgfEgbjbLTD9I
Oc5ohHJYct+C7crYVFlsnJGeL42tnzyd2qEZ3SXs9nRezau0N2n4Jh4vlwAgVnCyCmHg2iNRE9wM
8mYQqE8/xg8+9IPdLGPIsHf6FfY+LYlYpJ6TXWb34JqpZv1rXv+zL4bl1xdvMBXkPsVxb/Y1H9/7
gqz9/q4Yoro4dKrtiratC7Jh7CpMxcXrAe0y+C4+Zb69IvuTqkQC/fhA35g69girFaf8sBLA67qx
9TNj6IWMD+xqZ7zv7/Pn4bbk1HUNpmVOhutyc0qffZy6YbrshPRk/3tn9ftguBAcprAQYmYR1+Uv
+TjpD3UpwLX+1xIXAySz5O5rqF2pgS2Ngqo7nVS/cRvVCmWr5CxL3AWRvkRfmH15P11Elo77pJkX
QpaeKO8Re66esIRqcAUopOmv3niaeC/R2oovC16WLWR/TXA6oDjxHMORaTDQi/Q8PJjf7q9af54J
qikilA6qEZCAaj1Mqo4OAf9ItpMVhpC1nr5yqHOxZvy/hHMDunErGvlikYVzNaJ7iwhCQjRiURHt
LjMJsL925se65drxA0eUObk2quNdYq7ZMEzQoCiH1rOOz4M15cjEF0+YOMDjODgc6FCpP+j5g1bc
N29FmPUO0zuO80dIHgCPdX5aFHdMyw72uwgK9nROpLyUHjJo78ulLzq3lyhSApGD2F3gKzaLQOaH
9WnhaYGda0xl5idNKtlDhzb3RI3568Epush5NyPLUJgGxsxnv8UgXWqRnuLbNmqsFSkDbtTBYS57
QFzWmMqdoMFWztoLTJJzQ3GCjuc/DB/FGj+UTP4FZwX9EwDJUviB8VpFblwplRYCwAWI7AuvFhQv
9f+YhZjmMd5ANiR/i655aVVnPFAyeQUKKf7+roDJJXI001De0Rn5xtPE7O9w2TE5ZoDHNuSwUkhJ
uCj2hVTjReX22e5VF8Nmix/+EB4VPEWQejx4iWVlIDkd785s1YaB8xRmisXT2mk+a6bZUEFlAYXQ
YCX+ghU1npnPJtMGmQnNvNlDu3tpE96S7dzDBas4yWSR6WGXHSA=
`pragma protect end_protected

// 
