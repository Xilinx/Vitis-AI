/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wP83ygnX/eTUaSHKbCQu493HQGAwls7G2cE1jwWWFu/TGPNci6l5pnaXvzAMAfiDc7+b/Qp/Y3CR
P4W/K4m62mlK47g++9Y8TBiMxeAuPO9YDNKl9J9ytIV0xrMOcY7VuG5zyNb/QS2pTTkPKhrnahE3
TIO31pCkXR85AHy7uH6bsIbGkbWQQcAygLr17NLJO0NA5dgEPWVhCPQSzpC1HwDDwqnvG2DOryi4
CeQQrBM5XRrHU4kpSCEA0vyu4ocsFeIYrF2eV7o9lH1xZg8eQMY1TeUQCvRXh4i/rG16KsFiyrl3
JQbA+LxKwZMn6+rBUbAzhTzoTuJgQqwvtFELUQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="AQYmal0IxtZlARGaEAWRIO32qUIViEwMJF5/818h+X8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1103152)
`pragma protect data_block
EPnJf6MtG0IlgoN7FHoPSwbtQsZ7/pdJZ35l5+J0IExAQNiu2m2wyZCwUOo2iszQyjlfZFInl63E
WZ6TVh67Ue1k1cDhVdCXQRadC44LGBFVS9DrooKeHqgxeVbaA/ZHO9X2Ua+COICoJECS5COzz8US
7vb/QWskpqyMAIBM3FndWWAV44ZbnARSfAuRjgIgRb0QIuAoUEkZp3mqt8mc7hMtlR3zcAlj0Esr
8p9WNvFf5oS9x+KlyOZ0y8rV7eccrsoSrmG8wivZaXOIgoYdgW/tWYG7lNHCGRWpusUsAJrnWx3v
WWO5L/lafEkx/0t7ahGFds5PL1YEmL+ryQ71wL8687tv8QkU5IzteAX4Sth/yIDTMKazJiv/bM6o
EonNAfazzd/3ydQzKZx8lfDy/gyBI50L1wOeD4ePk9JtS0q3RQOGtdgHwM1yFxqQ4CWLZHn3mNxN
jmTa+ZwCAbpSVDp6m7lVWQTbKnmKFX8DpM69qrLpUczEdrUy8lqeYP/yISPNb8CQf1H3JVXMFupz
1mwWKH2Zk8LCXUbL9FNtmWKG++lEjxQ/dRveqgzerZdhIlBkwkG83Qp0rt71qJr1ngH/BRQ2rulp
KuISgTQrKSCovNzkZFrWjUxb4k5orvPNzwlNzu/XQ1vNsQQ/W597L6YuXMHIeRseHrpv3i3kaOSH
NlZUuFFCN9YeEyg2tkwkcesrLwu/9nPzSkkjFNqEWe/eHW5ZSZ772+eBjeI29IWU9fAqWm1gOjjw
U1OA/4YSG5hHlnxEV2Mhf5w4rDGFEahlMkHCdaJURuJ1Btgz+z1ASRo/lz/GF5lM5NAnVrmHVwvZ
lYn3TfIGBzUPM8I11bdM84bgGO2ANpmMHUeoHxObYxksmQwvGgmVnho3dCDseZPrfK1AWYxM/N6G
FRNzanRlF3px3n/xRhVOt3nPcCtlDhiyZO2vFpf3nAzSjZqDJOLxD9Vz1ZX/pTuqORI0o7LjM20s
EqmB+46PROx/V7MGAyFMO4fBfh8Xt0FoOKEe5MODE5mn14Im7dQ/KmdYlFHoq04aP2poZ5uSf6XT
wjKnL1aLrHLMEIp5fG/8mtkY4YKf9aFSPyefABT8A7Unx4X7poOJWTm9Drn1jEd+/Neq20sYHpPg
AUv99TO1dBRuu5MGLqvULgsMSQYR6sPubC3NcrzhLLNLm5QNXPCOW4WLqcATdvsDvseOUUt3biVJ
7z8komjy1/sPGpTSKmXQZCGYo6XSeBpplNBkWGdWc0j+42Wr/QWckCorIRG4JI4MqaCthiX3LD5b
aa7BFbEAyjB7TT/jNJUsikclDbk0xmbWMDuV36TonRreupHUP1fqpE9gzwmCamWWT/tF6+bkvVRx
TGafVuz+EVzybBIcdiNd+/RQroaYYZfSrEV3FvP0FKH4oyW8vRXOxy30Dcb0b7q9fL0nnF6kc45b
N74LBcw9Tj+d4E5Mprb1N0iCDPX6VRUW+eFIDgcDcgdpaCzK3lsllLMJNATKraqBPxIOUjgXpNtH
XJgIpRVfKG+/z021EXJGgbIBtw0oR5Fio93D21U0FFEtOBmb85qFeAbs16ncBLcaB5GtyExbsyMI
z0CMz3LcWMjH1vTrSdpD2g7hchai7lvEW/TTiqKkl8gM4m8NEZ27AEs1Vh+Xl4OceLNKQRn4vm/3
hC0T5PxzZOygVzIZZkr86YzuwvS82snNghaIKchRFn6Nlny1XR3URK6axR0JMa6QUsRLKI0wBcDK
lqyyh/ktcIaE8T2z5tX3+9vyDVK2+nq+2LIaR/+1wxy/6DiaO8o9hjQeTspsEZnCuFquMvEC8UQ5
XoDtUj9BjgfB7aTDUIyHaFYGd4IxBzB7cnS2G0VVefUYaFuNbUt5kSiqANHVYDSxK2FKgk85xciq
/j8oqbZNAJAM/kOFfW+7ueAZfpBC3NZr02ktWhlqBYyOHYLdpmCUPkyUihO+t28QB6p7E/eL7rOP
lj3zAIj+y49QwqKfhgM1ovI8HV/TrjBaIV7wJBD5ByIOzIoXJEcfF4oxvJKFOYqbXeVWnWRmwQnq
Kfzlw/wAbtO7s0hQO/FQHOqKh+D1s2lrNB5ihf3lTYv+bGImBM+z0sKRno3iVsOx74eE+2Z+HtFk
mzkmQ71p1MdUaBmF8OivUc1ovFEyfquecRw5s2XXf/TZcSvPuZW7+hPsJJmUl+Nuz7baoEbW6Oa3
5us6Nn0DY2cH9fs4xapc85MbWNVaQ+zmLONVDpSjvLluHC9xpIc/iJRkcFXZIb0MDFJfhn2WSX30
6uZv/nI8w0uHWSlPsOVYikmzQtPlqqSeMUvaWqvlYU/k2ftdKaryJI8QyNnBKIxcQcIKwoUc2V8I
hKqTPHkjMEQKxrkl+TMir6i7XhlS27B4ghxqVio8O6KB0aWwZTBZEZH442cbeFYdT1gDM/zeqRj1
b26SWwjXhAF7B0KyD913RxMtYCHjhzuDA2wkckMrBZL1SZj/dcXbsSHjCSn9g31G5BgjYgGwoG2U
T1N+z2h602IlIxq5uck/Kea1hsTV9qhZp0E/feQx7+BMZaB98/ZhDr5kOlvpfpQUVZc/4PHG6CL0
hZ5KjXbOzqR3CQAlezg8WOqPjQ8C0BXgCYB+r8JV/quLrdDGA/66zxonMWq9vKJGJvTGIG6Y0VIH
w1cBeBdpKGxl1Jnyq7YPeD7ytIts5KIWX/V7aHl+3zly/Q7wPggB5x0i8xDJzjUqhdzA95bEbV+d
I/hIcULHtoi671/okHD/GiA1SCWxFe0ffeRADLCsWvgKjaoyM5elreh3m5Hbbr1DT5q8t4pIn3YO
SlQBROM4KSwe9NCe+JyYOHId4wIY3LlvvR0RQBhGfzfRuYxrpL6kDjzmQb23K8wmmuylSd5FOkRw
SdQDl427ihLOepK/qj/ZVltMwcsTBcdMBCW7F+Y01oAHvfj1gUlDE19us84Xwh1K9Q6OcAD+lAKw
M9JA/sXmlTlQeDFTNwck4egkouGB612S4NjkWzBRCNA1whNpivnRbhkHn2Ui7ZpF6tSmSnP24GZo
yFIdzcNlyiiF4hkYg8/jEpvg3xeN4g76SAMRiXdfN7bUKTOhmsD0QZq3WUXDkPm+WP/NjP1eIZ9h
uVBCIvFtOtqHMZ8Gqb0Bd5OGLHEmEIbu8Ep8rloSv/JTCKjKDNrNzuAV7aBWdbKVNUqWm81T15hu
rD/mmF3A6chgADNBojV9PKZNgy36PcI/lRfDkzFIprP4MvWOEc6mB2A5smsRtZ2FjtP4B7P9emyi
kMue0TN+wQupoiA9iRHiJSsmVK3UCIcy1y83iIumNuqXk6FEwRwfRu0uRO1Yq552A6+6EuTRwZ2f
3WM653VuBarpJgtl2uxEjbKHs0O3eGvRffjaK5uXT7tmmlxa7HkGN6HKgcnzCnEX80TfEHvjrRSI
AY75tupjpva2cBJ15A+vHrF6mtMdI5NPFiu9N3Nv/3s+13OIyKLUCQpIPf/3cHEmPMlordj3esak
HqYJBDN5/YqyFyh3qcTFe7A2uPQmRoQh+JCueEdyatKX8w0ZUYo/CAuWzavU+pSPOi4XsMCkQMsm
8lj8XXkNwiaYY/d9QPEKllmwikCSqkJL98fQc36AfBZuDjGGa0ZBlVhUI/AUHg35nYATo0Y8Sfqa
e8dPYIsLjGdAOLPDCvdeau8RkpUCNq8CHxcBzdNIEEPNkB5kACwimGUeNOt1gSxDwRMv50b95iby
WJifjtnEWAQAauKZN36ttNdchAmVNf2RuQL87ysEV6aRI5W8SS8gvNFLuj/fpli6aby8Kfz/TjqP
Y+dqTuE/QdB2TnTh/eV5e3lcHWTwOlX6cor34zFKDOvLylpBaQROz7OITsZ7K+flZN8VM7Za6bvi
gtaR8uAZSVdvY+0BkSwC0A13Jxd9P2rk+b+8dIwgJePJZNuXYx8bFfh1b6YsiJbpAdpiwqgZNqOX
iYIXG2WGoa3x1VukUrCDcJYVC6kMwlrUB3pljlRRiv5gfYMdvLDsX2OgTi9TrndFzn5kJHCGPsYg
NwyI5W18pnWXDSPNV4g3O9qV7rpFLtR54bUkT+gVQCnFEraNoNACBG+OWisaoBLYsGUE3x+x9fru
Zy8ZV3aaZK5HUi6HtGIw+W7eP3p+cBcVm25CBjUGx+GiWoZdwiSy87nJ5hg3iUayBbY0rU5CRCzW
JgfVoFeOuHgdJmplj67tg1BYsGHb3lCWd+s+mGNBQVp8phYKtlHdLnR7O7bjSh95jM/SW7l0Zzk1
pNBrREEZU+7EV9C/5oO5w5iI9YcVSmVdF7bUmGgQhzJloZwToVq3X2z6p7amd8jqVGrMTUhizU3A
qOlXRhDOHnsFr+E7/pzfdVQYalX1HDeHJXSI1yFcR8ipwbz5dWDeVHVpZvmWHAkywCt6g/H4etSe
jE8pSDi3jQTV8Lc/xyc+IVB/TC9CFnQO69CsxdmvSQ3CvIfnw+WIiPufztuVFNJptXqvk8uIRofy
1DGLPcOA5fEjiWovSVV9sHG2RvMnxruZAm1mNi2kKP9WjbwkoucsRUI87PlhzdZOsn0tm/3pDRfx
kqymz+Rmbm1iQAs742Ne1vcP9ElebzvnFMPKTrsCAXfc7tnMdZVJW5u37+mVjeGeL02wMil7MmIp
9e2vWYGAvfPYw3auSt2rRJdQ9kHwbVgZd5UcqUiyNqmJsjQH3n1/Ik+NtQA/EtSLIOxa+uNE6dH0
Kqphg1xtJgR5g+ijAPPJx4/ktI2cF5AO7wFmelolbL5bFjlP2IviDxr3TI2apIRU96nVafLhZRbk
W7rWl8LDEq03saguSAnHQnn+koxi0ZWQ8Ie8parOdrAWc702Uy0ASQXOmDxwa3lcZeZHIxp6VAoM
tj8JxFdc7sihKH433KUIqSzmklmsblumVxVIMoL+YlOnwJOk6LsiWtOICC4I6IC0W9eqQW+mYCWG
RDxcCoU/VTK4iJMm7Nb7pyAelHaJvYYdaW8mF4hhA/fqMQ/uLodZ4oD9edc0YrDfyr+rJkJqdqXA
dttyrUFo6mDhyCk097MZWtZF1SeZcSh3y7qWe+UC0LdTX/18pf+UY5CYG8I0qzFlmWTDnbA8Sqp3
g9zoj806gR4RALBdqr6bl1HO7iOj9yaIYL1nwQd4ykkaojkoa+3NgLFybmctn8ruPHlPUdlEHtd0
4jFyZ3il2kbEfjv1t2VFL6TPh5xawjQnt0vHMoQw32VNaGeYjkEnccYUOKOF6CVNc7j5HYJejx1J
yTbzP4pjueuhozw9tW9dgSf3jUbvxDzDyRvRv95UkdUAuEq3+4P9gnPSh/8C2W0WDrW5Nu6kT5oK
o8AQz4WVa53fqWEn/poQgo/k0nPrMidQgywSo3JCPJZXmgvyqChm2EUCgWyT1JRIVxTrbGWbOGV6
pn/6X7iv4eIBmrmVM0KsTLu0pKbZjvtCnEPAMQFNNFxqKOQbf/HaCYXv4wT00J9S8YisS+1YJwfc
iWMNeuPoVZtjJTSj5KH2/0saGJPnTbe4QUnDND07pOosadPDV9bp/u5pVMjaEA3LL09C7m45RQ25
k/PffknWyI90qvUsIvriCr9bymmesuGtdUMMGGX0VLL37C2C57yA6psTPNEu1mhZQvHG5vgXH3d+
STqouEp0rHkaXJfbEh0K26e3wC/VecFl+rsYwTOurrkPut+4bmqQuphokRzjN2wfYIy6oThqDAOn
ZEUjSidFmSF0q8/J3sbOd9wtVCeaEIpgNoOlT7XSzS4AteHjS+g0PimX3FOwhI15Z+cIeuJiIu4o
VaW4QeshCLucVRVpJu2rtDkSsK0/VseQB8ym15iEaaVR/nOYqOikGL8Gh0hWI56rUuitYghfbfB3
Jdgy5HPiKUqxa4cm6Wf4G9ewsi3QQ/oOAds2I9B6RgMGlyvTAlECvEJPzFPe3QAbJr/2top9ZixF
vpwhVN8v2fj+xMQLNJK8X+joJoVVqTtmoklYa/P8zjcv+vm8vWksDlrimJHsRxB98Kcur0UHQc3Q
U867QKVybse00H7ehgRtaeH8pNilDETG/Fx7mf5HNbmZlS3CIJH9q57J4Y26sbQGJ1sONEXTEtSy
yrukg5Fa67kXfA9FibQ2Ucvccm/yzylQmR+Bf61J1Itn+Es1FYZOw0dlR9cej7yuQCNJkjbi/fcy
mkDiLWkkNS1ftOmsdq2wtbeFJ8VEH9TzRAcK/+3IwC/0exsdDutcpuTNOm+V9+ks7BYAz8NdkmEJ
0fAK9UwhSmukLvputoyLNncYfAoKPQrHdv8JScfzT6f2nXzdpglabqGJU5vbH6XWYucAYq39NOpS
nY1TeQa0V6cQXI8adyqKFsjUQNVv2H7zs3R2YjxJ72Vt+WR2lQ1NRnXzYmVsImKkfSxKLQR4ygKT
SWrGzkt/5lYad8e1LI/mNjpofl943JaEUX2VOO9qAiahu0w+X2eeF+FW+A1TI6JE/CglOMKk3xZ/
eyMur5TiXPiiEpXPjtugLTkEZTrmgujmqrDDYjoCfqVQO4OEqk4UnILj7fpCVZCPuOsdzgZAbrHD
yfIo3eWS3WNUOk/uJ5VQMyMzcZeSykJzXCZSeTVOqjZ8u0Zuywt+NfYNWzT4pjaJNMZ72afpTM3W
/Vc595obSJ7EbgQKS+rfYp9pFBLLlqsnCcG9VP6uK3G1xkj7Mycn3bYR9BnwgUInmNwTMrOh39IL
6doP5a0Rv2P7/Th8qtA2pvr90P/efOXtvGoEVu/XKV1lpZAtCszEQxgOtvR9O50QvERNRIB+huHw
INQmVwZnK8gsUnP+C4fJmuQVXOo0OEkVlOThfl7KdzvZln3jPbMVkNe8R4s/AgFbeImsKqJFJCaP
vlxAVAu4BVARUI4iUMA+oNAuCrQLf8VXH2qG5NhFitZU4KWp86ImvABD458Fm7ReWNDerfvNCAVf
PDnw1q4U4I+Pj3RU0y3w8lvGAx42QrGGYSm21Xbmd30tTORC/dxDtjTxGcN+UVEdBJJ1iuO+5Q1k
sorot6VaYao76ioF7Pand+htyg87Cz5gbGXGvmcYtZIvFkXRTZcuZyIYQGUvxeDQy3D+Hag0cXOg
Q/ryJDT1MQICxIBZiKjB1D6uE8Q/dpTQ8Hdl9v6L9dPznjKi8WuR0/A+BNwwGUgE4wo8nm17KUeL
+IJQzSWc/UcLOBAFLWWec5b7Q9uCxh+LPOB2o+ySe3ESHkR0aoHIiYMnYX0G+5REiKlo2FHCuXMc
jkbI5FwIhhTZYrbc0F2muYA8qJA9Dn09VR23us9UwTfSDZuDskqTtC7zju+0EizfL24Pvhyef6jg
I5kd/IARJgr8cGr5wMyRptTyoqHMr45oKNGxXmBkvfCZ1KjVj8o/anyUnNKmuvoTjH6HfD039hfJ
zYZNdvqKb7MI8GF8PFXtPzGPrTT3O4WMrLVw8TsQWC8NjrtuIGQ2aYI92iYrRs2J82nXIsAwEZbO
lPr8X7yEFUfmgSTk3vTzWZ+Zy+M+WgX1V0iKSQApPjjAYoctt4GPuWmobJwaLot9zrzT20dZeXjj
CiiXwoNV+yg+zWY7xklzsatwFVYAMErSmG7ohejwQbDlobW8QkyFv0MatUKSYiGjQqwVFwrk9EUz
g32Kp1VH+UltPPet3VLXn+8c88JgZt80eykoxlULBa5tV5Gfu9gGcVM0Rj90eZH2lzlxEQBWQKZI
GqbJ96cMMfxwTOSdH5YR7gAXdZMmtps4e2WGmJT6mDBTz1rXwgiweB/O2LsF4YF7YQEE9fLWJcz1
EQyDeVBCu5JXu2LXaxcnjGi0RhXXeooiO16bScJWsRgGV1bZkyAncxtBADMYPY6Q//XjsWSzFpdP
hRmAiYVgdaL0AnRZeo1XUDp2GwI8vbI8htpsjEJzCN2tlD5H/Y1bqn/J66jcUf4uF+LkyPRC3ybd
n6sTqHL8X270g+/QYuk+YCGogAfoTjIyI68aF5hHNUUQSrWnIKuP/zdd/kRKr8bzSPQFBVCPWjAX
K06yQOvGwLbb1hLsTCC6RHaD0LxhSMDeCieNLV0iZ1wI0Wlo7EFTYmjEJAMQtBQEKdebwYdmULa4
vVzyLSaNL2YtAV+hSZ490ZHMIbONSqCCrXKkCo/LOW/zdWfzux3s6RcjYecVw4xzNwrKTVvnWByP
cmFUxW7sZFwJbs04vaT2WpbG/s5/ExRiJ/KU6WlOoV0imIZHHErSTDAba3lTbilWWBFIMG/RUJWv
Gg1XlV6NYKzR+XYzjZUxGZGVJm7RtHW9XVr3ccrQaV3bXsukFy3gj5qeK8XqBG66mbP0cXXcwlSH
mzvWeOxVMkkLAflNni/ctJwEAJwEQ6f1MLuTwlt2z8zIgzMu1vnu3HOuPpYKgaF4JdabkwvoXOme
ShVADV2XTOR66jHivptvicI+w+xrQVUtnHN2XC+efYdvBM6tNP7ZpRw4x2pMj2nu3nUpRtkR7u7K
LX+DNT7nr2gMo2AVtrv4V+WGVMq0pPahCPUSz2yGgzceIK+Pz0fjsRDXrfY3/eueRe9yqPRmaBrV
3zbknc5lgkCwTp7XsxS0jKwb6Mnxfo1+F7HmUqEiRyrl44Hb1tzC9N7bW4EZFaDuXnCS2ZnQ3f10
dB1kL7Mo5XC9b6QfmopAqPMRA2aPV+e9c3sOtESQEr5S8TeTZ28wmmxtxuv+BoPotdKIVQ+WchPs
S7OteAbWKMgm7eb8instFp9GptgP+2w1wp88GKno3bKEQuoCWJmf8txSVyKoFZPRdKPZ/9nYfQEf
hcG7bN81mD2yZ9kpZ7tdog98+VdAetaLzgKwVH3rVr3cs98oHd4HYzXUHKf4t129qLcmZvOkikXX
1qkFhhZzAG+/oNBxyMbdI7i6yOgw94DIfLu0X20/qT2fdr1w+/pO+XoWex10TuJodpTqC4nRIM60
t9DgJBge7Qz3BPYVVSjeh8weLO9bKbIDjXT5wq5Y64hsKQjRL6jhk1T3QpzF97HcqpZi8NNVH5BJ
J9wUyxyThupgIhU9bggDBdwsHQLX0LkYASJ0JxZq6MdoNtikmP8ioc3EeuoRolc52xIGaVXuSMNi
Q+twbUlue82kaaQwVBF3lqTU5sNJxWDPbZNIIuKv85wMV7afx1n7uBHQlHyr6DJich+Q63xC2gdb
H8rveOQqiHfm8GsJIjDFSbf27tVuex+HouzjUsV6i5iDhBADm8lb7mUVepoWgpfjEOX9OfnOD72O
csz7p2JIICta8SUKx9f7HfgxH+O0CxYWk9llD6y+pTZkv0IBSbc4dNGCP94H697vCsqXEilg5FRh
kKaoDQ6MLGqf/O7gN8GGOXq/qVWAnzSVGD4NkNHBd+fxCxdEB2/KNrCFZBiQvkIq1q/9gtYTXcyv
x1bKifeD86sltSgmxVwLiHIiH1Y0bnh/vFvUqERO2FefWLfHZFaOLk9KhsR5C63xaI9te7pqBWa8
EmrTQmg7yWXjbQ6jd6KwrMhIm6zg7gbTYlR/GQxeacPqcPtXmhN3R4VUQhbseflf6yhIfvecZxju
vRXfJNPr0Ha7bqaVd5rPCivenVaAhJEvCn0NAUsswK1OOnsrvR4udK8+KNPsy/FaIuGwPE+yTsyT
PWLmXlXBtDao4swIgdhs5aI7qDg/MvKV8rc8VyC/qVUqyg/OggaUzobSptWHN5PXOr3KCPAJPJkm
ACp5ZOurD8rBDcECZMbTAR2uCao+jA/QaVFJg/Okck2AsV4j15wZQJ0B0SI5qlO8AblwJXTKqbtS
wgzAAjKBM2tMK/dfg1MZYlgGHZ+lhoaZZJqxKKzFSApnuo6oo2atxUjaVQwKhUorbPFISWvrkoDd
nozGlfn0Pz6Dr8WeO+6KFiUxBZII3gzYESDoTDQerjChK7Bs6AguRFClbu1sCUV8TCmm5ETc+rJT
M1y/0JY7/eQr7mlzZfZLV2cKmsa6/DFXaFR83ET5iONSWDFVA31j36LGR9Yz328Athf2LMjvC69n
6iOv2N4p7nPktMqlF8gZY+FHW/GlcCLIE0o8FnEnkKUn9SL1qXsi8cNEjBPVHMxOF9Gh/Yzo4ZsJ
N5OmWEp2q13btcxAy+J9oKiTONLoehklOLpvfN/2oD4lhxCemk297HafYnoBhL1m/6QeeyNbYA2m
7I9+zQY0CcpzYFflJihM/GTETNTSSxvz5I2K+Tf0UX+SyS9zSd6eW4nwvw5As/ht529joV35VDEb
Z6hiQ/rcRX2m6ZyKGI4rAWQdn+enI7bVIatnY/ZN5j7luat7AASaKJgnOoZHOPIkbKixaYu0o+2W
Ui0mjVB6ycyq87FYquGdLJpfD5mS4oVUOcL0NUZK2bb5sqHaJXqNHv/ZYtnXI49aKodcl/FpP0vO
HQkdlMRa0K4+FUaB6/+qMJwGvVEK4eOJOGFIxekbAqPM8rBMCFGZHdwyW5McaxHw/65ZA3+sWuWD
f7Az7kNhB7+IDLVdLoLNAgA5/EVNnH0YrUxmxxN/jifqbgWCJkrYEZALKeI10s5lM2KDWtzemBlI
21qTpfWd4ApcuKOrLTlI7NpWnIIv48Qr1RCHLMZCyKCPhsKGTJ4QkOWlPS26OSrcDwAW4Xz9cfmm
8+cgTD/W/fV3Q5d+MHbFtUyV74eZVr1eteei0QFRNGfmx6hexsANL0owkXRpdSLPOjsfpwEcOkp7
xuvdjcyX6ueLzPIAI0E+kiuw/2ASLX2oZiigPDb/IGwiwC8i5PAoDUo41N/N5oh4izMRvPk0ZJDE
ku3lCsRCUSLh/pSrfS7wxhu/qxOcmdNpJKepANT2fb4fJxJlWvQHRkGzVZKW7BVy892ZzXLQHST+
XyPhiMKypB4IBLPl0f/5SxE/FalLrdbyVXurd/ZmTJfSOZmoYOyA5fhe/OUrpvUZa7bl3UF/uHrL
7VMGe5+RsXhHdtgKK+uibdrf5+eMh/s29mWuejV4IbS69ugdfcGLCh0T7IYh9nTEBmX0pl8+Dwy4
lrtwrbs0eegGlCKHGEOGR9D7LTVAJrbh+D52xV4TdIfiQdQ6A9ynoenIrGHQj9K+tKiAPYMobS9w
lVG9oauw7vJYAUZTYM5DJK5n/rkjZ6vlCWP8GO4GbL51W0JDueBSM1je1J1Bf62+2sTCOdk/Y4Hk
A6d7g4WPOGklAN6aDRGFVtXHSzPs0on5n5iuz7S5IhPKMp4HxFigL5FcdqhX9cSl3M/Xs6RxaUZy
V1T7Aeot8buaz7WVZrg9xCvKEbF8/uuq9JxaZ/Zk3gqBlsXl6U56i7hVkRaVYeriNDWxzokOqvnv
AWmVx3jQ0u39kEGWkYka28a4kRK4xP5fONO++BLvu9JhZ1G1xWQBLoeiqL3txDe9ixDypxf0yQdZ
Asedf88X7KSrilvXRuhXp4O+1hzSgnW+HUzjYaCWTjnlZRh+54xYUCAcLjDAwetBDmItV5LLRzs2
6vh2EDwJ6i6M1YHq/00HkRngTgGpzH5YveLodxMC5RGQ6QXcxdegOfzTVDM8R1zf+tp8GzjRFCGU
wk4ZCcx1ymHm5bT/eGK2/YbbTf22ov3YqGQZEqreQSvk5z/kfnyhxSFyRxbetail7JOBxs2sdcge
V9vHSFADSJkiwz7L/FlrMrBtS/srt91w8v3IyB73pO2U6KAHKyIM6TPkZzsijaPStH0WxxWgnG+2
01gsfLdYuX33wweTcY7K+6G70wlcnWUOXlBpH6qN7ge8cpFBG4NlPDobn4p2BA4KdeIxjBMfS1W7
D21+TbxRnPq3TSBGog+e7GOOYvea1D18d7u2PjKyDLUWo3GqlqRV/oRjbxyBwOauxvQYK6wRs/Md
g/JEK3ggWJ+sxLr9wkwxXy4ZdVUT+JKu49a02bP0xulYtZSSkeU7dEBqirnKEjiSeLHwvoFttF3M
6gaH4jOrCW1xc+ur2FsQmSX5p4g7jM+zh2dfHeXSl93fCqpgUe+n8EqEjL1rDScY5u0TR6v+JOB/
opj/oo6I0Xza5wO4GYg4SdoUDOz63tHWws9BPX63IEjghnjITCIz51DX5z3Dd5J/0Xg5VPJCUsYP
/EjXE6gLw3NRr3zZ3Gyz+ZfHRHA6EFbFqWMDMaolVv0r/FCQdkpN4UQp+5B/iSyAOxlLTeT41gA3
I1Kfysv6zU9iZv/LaLCHpLyPOyMe8JSDUqlTf42UJSOEHw8dBX2RyVrPE6g/WZ70DbpmrQfvWTnZ
WqnLKJ4v/QFyUiMSqxTv04OqYHrhU1h1IaAKKK3Y/r5OCpnWUEPSurMXZYfzRyOuyGJEgqSEqW4r
S0odAL4udlGtiQhZ3L0i/L5UIlxTgcmfZz87YEFoN9nrhQkaMDqy8h0fMKqzivGnPMYJ0IL+dFYh
3B0Nf2E2bYDISuTrWhpBBD5eUJJEm/Wiska4eYk9ZzvY2xn1Ipi/qyArLYIwL4QpZa4ELgzFNcB9
cUEk3pzN3GvtsT17MTpRzwAXDGmPZVBcjRihiyJz58Mr1CebDLfHAw4ttvyXFIpjI+c7eD27KUby
/cV11IHBB0fc8yFSvkfKVmf626wbVO+m4aeAsSMAN13SCqTRKmkL59JagGLUUanFWECM8KJcw62O
8K4H5hJmhWhH2NDBU49LH4VHkJHipHH5A3GOdJRL1fQ6gEKvOf651X2XdffdiIeSlQI0DXuymVq4
uZSsSofOfyYe8dcb7yoQnjZpU5VnCAn01HQ5yX2OJh1SQ+8QSo6tYo5Z2L7eHtBSl2sugKboXpML
Zyde9YE87fBvxFBamGIWVWHwGdDN19WpFXb1LThdckYEC5dhhaFy3efefVvRMaMRveKQjqOkustC
L4Beqkba+mb26Pbg2P5Ugn0h9W+BP4v50TaDMxcbvb3lNRZJZM7urmDUYwT8sEMadSst4aS5C1yi
/REE5A3XtE7yS4agBFaC/tT1XatOrlwjDnkvo8/8FBFMcCCSBBm352JtPPzSeMCIJbZrxPYXg8oQ
IcNxg64xIBg3G8WtTAKJ6dCaiD4m5uoVbf8AOWGv8K/PCeFYPkGSJbeXZ0wnYgPH8VTqoZvb6nzw
SAQHbtVrRGf0jbPtfaXlgdWvIFzGrpOwUsR++F57eb1bWa5eqTnGuNMwLfinCFxSkwIWiSpiaP2U
x8y5t6eOuQnobkDNIOyNGzh+bxvZA6GV8llBo7SQ2iJwMoVf4Wixak99W3C8X4VT9CEUY5I+YlRS
tBx7D7gnzJJ3NPkhknDfmZlnEuaVozkFi7IlaYrImEsl8samW4HWVqbb1opT3dPdRoZwWaT13NCL
+nRLzlSRTrQO98mmJYHkm/jRvt2Go0FYIIGaSald/rpK8VoK3kxTVnLKNuIjnx3quB53JloPqxra
zxZhhtSPcfVyLebHQHcVhsFHNW17rsTLhjhot5+TuKv3go5+6rGB7ZF96gb91J48b2tiDVDb0kQt
jvLXmC8EdLw16Md28q/+IdMeyMwflh0X3dy0JsivNJFBvTpu1Vvp0+Zl1/c7Cq4qi/X7zDHgPZ5j
biSct21fvaHUeq/n4YZ8ECu8ZuNX5OFxcazZi33ksh8MYgI7Ab2NwhH7xdHdgUGgWVU/EMzvJPz7
pds5YAavoD+hNtTyfv8hE4Z/BgHGrZDoyV/b7zuREgyzVoyvSUwpyVqqvqmXrnHMh2dlVSuZ4tqu
OIovH1fZ5L5PKIgFytI34XgmJBspShZMk4fVpO8KUl19488m5jn9DbyICyBDRoPlq856zZeJI0iE
wu2QPoLXAZFDrkirUQWzNZbgHdQ2C5BkCwSe7lVDpTxPS9CqFhzGw8NoOewDFcPanhaPQnHkV5Ov
Iwa62g9mQYLelfGktuvUO16oi850o0+PgwtnV9HlZ5fHylr21CFeyh2QKGfbyO5Utt6TXvAJ1y9h
2hqYZpD9L4mMyrJEZzyGVm+MJ2aiSt0lKi1LIxMaaKlx6vng8tYc8gMqGNTuliqyvItjIQjNWRux
Rua7RxLJsTRYZ/JGd54euTfrPjrQ+BzSfMQlzuEX4kZSsmnZAiVvHmJiq+2DUYnhZM6mB4OJiWh1
6CeCflw0j/Jsugo5vLPsM+bJ8ePr20asX9mYAB0QYoXiQtSi26I5S0XIBwmoTe9duvOU8NlEozGv
tR43/vWDVPzV7uj4B5xTk9pWhSuvD5x7JYGb1IkJZVlYa6GQL1WGoXrMqHBQ6ziEPvCClsb1F0du
KKy45z064hb60wXXBFewNeRsDj/AUDqskAtidazznbCbfHH1g/yTwumQSsVc1IDKuCD6lMiUF0qa
Scg32qPzSaSAeIzlqcKFauMQPCBEfPeK7Y8/R9+8k72qRhqzVfUHVgdJpju8GyXkAh5+5Zk1r2+C
WpFrHbGdLd9KIN26VM/iXWm38HmvFWZu0GUXrHwyewpBlMoF9035capXRYuWxQYSki4wCWGtjFdK
Q5AaT81xfnIlTafWLCrbEqE3agSmXAbBJScV7OPGe4QICy+YPiMRqBaxaBq70m2uGwCQKY5MuD/i
bnTizk5SVN23Dip+jYMPT+Dp4w/jnEbsoONRGnksU+sVaeUaiZnwRDclqsokI3nk3jU0YqSai6GC
Z8+gFspCfKSRQ5q6BxudA9KQl47NjDk3Sh4wBNe2Cih1fbBZZ5x5+03w5+N/6LTEXVDJ6dm0DtNe
UMeIBQhSYahmgm7W1eyZtasDSEMwx9a45gKZfeVbyzqizddS4ndaQ++lChyFPXYMjNrKeG2z3Q5X
7ufrKqE6OLBBaSlSQ1hL8qADatw25xEOS7yK9BcbPOGwroqweNnOlyWXVuZ7ktl0WNj8fMK257DC
4EJdonsycIB2ptJEsMYX/LOZ8rUdRLHhAGRxTqgj2esYfqgEv/0jFhK2dB0iYTUevsMHMhKRTHCB
8M1JU2QUHmy0wdZv7JB7T4O7FLJVJMTmmBlkPSJDoaYgKPiMTP/oGm2eucKju4QP/6vY+MqnWFHv
FhsDqr2T2zbsh6oE+NfdV1z0A9uB3r1sfBOQd+Vus0ap32Yl0oEkzqqLjeL7gGtfE0Kcz2CxuvC8
1FKU5iXQ3dIXcnGwSYpHVZsobHtMe9mMPAE79FPgGVEiafnJvRfxhW/6SdFvfKdK6wHBjr8TR4/S
/4JSKva6AWZeCr9+x69U7ND0RUp/IIN1qqqmUlAVVCW2sUscMiOXmNfegBx5i45fkqzzJIwsodeA
bZB9aze+HX99Qq1CcOWD0BiX+V1OMHNyu9bzXOCW6Hg5e9xT1zmIk8hztKc0I8r8cCisswZdSLHL
g2dHHe9jo8UjeF/craKg/Ee+6GIh79j8O/XX52unDAVQ8YY1wPdVRt23PC67bC93oOvcDJrbQK/p
AlMM1C0nLUq9w/omH35sCBpyDpcdNTQI/gQmAdwfz3d8zimbf7x8eNopN5ArMbCX6EXo6LnpGMX5
MxChyoUy++ZavqloAqGwWUPhFwbYuHzgnYlgvrv+xQtRxg/lkrJ97bjVMgblnFrhCkbG3li6oI+m
Y/UPv+eq9PmTKYTyiXnnU5zO1P3DBKOxf/Hq3LgFdrPWPshzYeRfgk/WjFLAiWvZqK3nrGi/E3xM
JGjanqNbM8t74jjoOeJ8eG2H67nuEieJ2QECpnFqvs7f6pD45xullybjVrtEDsyXjezFYxhBG0TY
CSTMdcdaQCFJmLCIm2xV+8Lsrh0W4OL9u7ZUDFSxEkVmo+z6gS5WL4ylw2uWwbtcZWconEI3xB1e
mO+iN239EPYC1hZg33UWZ+hPy3GfdFSTVAWVONH4I4waJGjdq0HimyR9gehG7geEGX0F+4Oredbr
3GAe0ytYmF3+pDOS1jF9pOyNp90kBHbdcWTnlLjrQ4sKU/5G2Y5rDetwaDDwOCkSU48IOCksttu8
6ef0oxwUmJKzWz9BxkZA+rRG6G6P7xie5vqLXe4heEy1eQLvtQVaYIGe1vcyYJVDsa9hT8vHyV8u
n3YCUo0NnHRq+xr6keR5sNDWUAAGGaQ/6JGAUu3N78nWZXoXgLJYu3qDMeGfk2UvRV6FJVAvw1ZQ
uEa3fAx6arT7wBCCyIUcvaEB5PuhYTTBXT0DI84+FwgdbTeHKLyWmXqBMALoMcX13+37uquWJT7h
oM6gb3SgQtMGXCXIo4Vf4VAih4JBKzbEPAsOf5AiouG+ANYmhgxZllnteE6xVZB8xtvl8xgPDT2M
Jt+8HSKtc7wP+hk1lqC8yvK/OZsGH1gVIGfMuqHm1hYBXfPySQWTMwLaDyATqVSLI/lOvyagapJl
NJOi5mnqj43u4UsUdPFSGNQxQHbIjPdCf9EKqWHcQmq0wSv/KScD4lmrn/FVDiK93a1/C0mWtXSH
c2wjaNeoMMN7YYajLbPA0iTOl9SsAvaLInKbJeqYoQGPDSqfXbmYVZtYgDKSnFBepj1We+go35ti
ARKSa1UUD+SYktDeI9izsO1/fMIzxZMTAFtdsJSaxv8/LDZZk41TnGZ936xDumR/SlrDsqdhaCG6
L9877EdNVv/DFY0v1wCnaJCJALvBZlFRWJKJ3sEvsOajFsgmMc+YytW3e014Dk/278IrDCRwReAV
gO+HX7LrxToyHH2FHSWQHz4LPrmoDl4zRzKJmndXejmfhU3+mjRRnr0ATIjUd1uO7y9F3190TFJj
ahVsqVS6pU33zowxt+GVFU7BWEUd4WaOTm6KjtVbov4TKmvGxy88mN4010CnorLJ1gvUAje3yvac
98EUCOFbUPH2bdzsNdYeD+S6ohG2S/q1eSY3c87So6WjyR3GqangMVbj+uDRC3y+YrnG3M/b2Uai
gMMxQ0N3qA3/IdTt+wvV5X6W46KaEWGkBLlG98kksN3PPqmbUJx3Q6VWxk6n9tGzedvS1HIxAqxT
Puiv7qrd7sTg8gHe15YmY03cJFzEBBdBGGe9VmGOfxqNDqRR9KP/WnvQdfB7GJpNAvH0Ii9F0rOJ
XHBcQ3ucQEOWPLp+mX5EocaZJ448KuEwsJABt4TfwMtNcrVod/yRSI9KCHUeUOcmKOR8LSVGMw47
N5tJjGolrvamCuUF5RSXN2mIIIaETWkoLos9mMqseyDgYKqs4pTSTfH2L/BwXAZBRZu8vvTPxWCF
QC0ONwfTu8Gg6EYen1bJ+hixIZUG3Gmw1RsH1YuVwTC0yyZ6rILQP7l/ngZS5t0SauPS3MAUxCBL
tL5tFhDOaotydY9gVMroh69anbDm0bY35KmavNZxI4YGm7P3DSrS+TOmORmrU8UZ+QikLKJ9iWAn
/qVe6E6J/dCrVdaHGpkcfJh2T23c/VWV3+Mw7BBQZV44ezO20iXebsY+9XMDOrx3rxukj4lSGPv9
D1P0kMpfRM0XGAY59brlyg5SlGFsYSGzvl14OcaiIWSG8y1VV2ciecvZ2zMahFHdURXf7glw9fK4
kVGmAnJHNrd3BP0EVK6qpPtRtKalRoL3bC+jP9+tWj/s/qBowcN+Phj5cyD3KJGfuTlGNyljqAQo
xkzrXjxlQ/Zv+BD9y0TbDqWJOrpoBfQKWVf/TOZfwT/PxNHzKniHsoJuL/GU6wBBEriqhkaGQJsY
tVk8pYoXb9Nn4GMILZHvWFQlRryxnngMyiA5rMTL7KDbdcBrcybI9oZleQ34DqcMFvQYYDknTk2r
leFUnhOkKfigxghOwf3305oPZOp5U7gs3iE6FN0Nq7ulGLG5VVH5IfgLJrgnkKHNzbtPRSv5lHEt
Xk5BIovaKKsHZe1wgOAIzUYj5mn5kygYABUDbgeNLbq2rFTUNA8oPT2Klaxi7CN/b8GKVoK5CLi9
OLRKB5s0x6aKydO1P2wXA/PZmeD6BtgwfZ6jgGdGK5ABw9QilRX+dl3NGTcyfsCnl19opcOpcbpg
RfKXzA0M/3bNk+YPuSFmoRKfOKnycx6TAZw6Lz/0L4rMPDN6fyPZ5FqEhO2czo6Ilqctw4Q+xaEf
ObD/Gl0lssBZ7NXn5lbCfkOnVhSaZT5ijxAmUQNmbGn8aOxTcUjqioynIabuHBZJ0bYjzR7v8itk
huLUqY/n+9oT7TS3TSDiAmiiBdE0SHYakzfS4vX+c8Kbf4hx+ZDcLcINnRzU6chbJh+AxvDOoDD7
NlGohsixYoaug4PyTFJuwqmWcCkto67iFUR0Sfs3p5Kk9ngUzWxEEki+FwGLUxPkBudsDFVaxzUc
3lTCEX3MQ74swZ/wbxxRf05ZT3RLa8CmufFgqcrNaWH9mKbcbtO5bkNmwA16TZoLWM8MCyy0hM4x
IVYIKVTWucWcx3vPbsQih9sWTSJeBKiHXoKKG70oy74e/+H6mhI/JIxHOBJ5FAXYNrqeJqIk3mXb
iv3G3Lxt29OsPhHBZGnyEZzr3ozYJ26wUhcUEAIhQRE0tIAXWnwM9HlDmZJc3RFbK8SJahbSKWR5
U7ZG12QYXgII5X1JCKSEC73gEbal8p+bfWiZMfNCNKy8yTUXL7iSocU/Zggw7ZZYRvzvNhuVNtLE
bgS/LolODB/P+EehgbvCXD/PRZemjULu/B/orcD/aim+TAoxu3hJPIoAGkjSVLdnz2wwBiagHoyv
lYnKzQdhHLUyvLKRTEpYeWoeuXIu2/zYwPln7Dk10JGgA4kOF0OhBAa1jNUOX6qQXuz03AJ75dxK
JMaRAW5emlKpHacLGYe9rXeTvTW7K72NqO8oBkG/JXkXXZ7FgzCu6mRDt81Y9/O15WVIs9NBnACm
NxXBfSrQYI7VvJzb30mEZ5x1bGNmLahjGZEpwYEfqoCYb3dpvvRDvixWrBhLPR9U9f/RmlYgWE7I
vVdN5q445wC4Z62cwysi5/wgWj7rwWY+G0JEqlc+4mIgkJrVRGwl7l/9MVgCFmQJ6+74/Fwujr94
SiUk8Yxk3hzauifect9BsiklKZ2mYr7rngShvSsp0Nf4cOXEij5tvaA5WCawUS4NWRcLaw1mF7dx
UOcG1nwKV1eadxoOeKhX0qP0Og4+HeA9KrTlpojhLz4ncWvCEAX7khH7ivH3FzHNyiaHEoNQ0ITX
Uo1bEQXTqnjgoYfLAzjTdbnpKkx0HG95DWXMp/CBXMGetE8bEO41yzagTp/mBgNy+0EKqvEQ6a1z
lxiMKhKNVyrsG5tTPjbMOTSaVb8mIgyS7d7TsvwJ2NGy0RUG6I33S/8kowcEkT/SCp37diVVVKJK
QFWcsLdgzyogTrPg8Gr5mtXLpdkAd+Lf10Z3LVl/2zwdgjoeEXhKm7RzrKXzusYrssCAjaB8ISmO
vrw3yHsJ4DQhDdtaDblvl26638j7d9qq5uZXphsRyYOTJPyxEYcaHuK1z3Mq5OLjgpN5R/M4BhEa
Z0NgKkS/5fEjM8QeqXdFGif1XfVUKIPrYfpvY+FXqvyH00DVtho+DN/u6FL/MD+hnszOInBXwjdC
tx0ZOLySEkQb4xiJgxFXPH96fw1/xNrYPrz5WR+Z7QCMmVfB8dcodZQj6+j0TnIpDbVAntexNpKC
PCv3gDXcScu4hjw+7NNrvGv2ZOuUsnqiIkXgQkumaZDqGMznqRJA/L7Bhi+Ng/Mi7f+FReazP44e
8r0La4bdSbPmos/x0FB5PzaYpMK3Z9ERmbhRJR/Op+HZsElAe3BhNLQOnOmLNa5uqqtFveSyP20e
PmSPUgNmUJGn7t9sqkAYdCfjlkdliNqVkEnCwJXBX2dOtqVDWurNj8RviRDMrSUBl1MVzyM0XvNu
iabzYgA7svUvC5M2fQwj1tP2M4t0shAbz7pz3Q9gm34gYz2Oey7uCqixbwUt8pk0W0XAbgxr9lbt
a9oM6ag4u/k9tVM9ypFqt9B/vYJwi96ewAkmc0TTbFeCRp9dh/9Ypm0lpxmuVimsL5EMR5ajfb3g
j4/TZoGottIhHwU3a2rlZ5DNDBn97NS15fvqL0/Y7vXonmtUCbODqzd80xRsG1L47C6BaiWomWSg
syTtJjyVl/aVFSrIANlYDTNkYur/kivSOXDRoIRx8qin5spCF9OrdvwFvdwN+MCsWuDCNZkO8Bg3
yzaM+CZUThClHkwr4PhYgEqbi9+5zZwf1GIrIew8ElGKEi6pKtx+tE809eqrHGsBcIamTejX1gMi
FIpZUz6Ise9J+p+R0DRrUO+dWIM6zjYwRArpJnLhmHBQFEiYdqIqZ0CLqZS3w2Uz+9/qE8vgSAb6
+9EqyWXvTvDDwW0M78hzrhlEPAWAlaBZqxOZUcPXrgXtO7gDTWRovZ6JT+ZaCLzy+mXF2FcbRPjK
QiwuOyKrBOQvPCNqFad2R8DYsnjVcVoa+MwuZ/XgJzP5D8pp5w+ItUS4Zmg9ZmPHHVHfTGoHeQy+
bZnJvsSXL75XnOGCQLWIZbeFooKWPR42AT7MR3T3x6gfxTXIu1AYAAkssyK77z/8VSxfZSNDOPuq
A306vzxgFmwj1fAwD/p5R2WB7d0V93+nWvs+RvWWvOu6VZJTNWgEE4YJJ7+l+AYTNderNi9dAzI1
GIwIWkiWWhLRGoBTi7s5x+nUhuXqzMXdEJdZ0Tm+63Bk+kDqJOjLdtklCNSIsYC/EOiE+QJYwTJy
tYGjPDYigXdQ0en37hbHvuvrpEe9ednWKHW1XdKGevjx0fFXpUgI3CDbf/MKFpcsqvNK84OTl/4n
Aw/QziH5m9Ck4pShzC3BLlhZHpzTMLhgAYGzDJ8wNKopHocv7MCJHeb4wgN7gPFiCY51X5+hTOSw
F2i/BfwaDhpIgOpCI+n11nDlifPu/4ooefrSiT1sRSdtA90q0I1JB+CUXogSEnklqgcpzjIeb0P5
vFFEURp1HNEX/W5NDhTRrLyVLyVs0kTJcmThPE9E4r5lgHiC1qBiHMOvTfhsmTanl+UV9u4fR4pZ
elfs0XSIAl0qdYNfMfQZSMajoCq5Yl0z6WT0yNDZPYcS4yyOs7lBL/vqXG5gyjIRJwL0RpqnX2cc
c91cZ8GxlQHd+IS/ooAFOmfkDUUxpBpJ0jamdTRNF8EBAVB9vEd2HO/WYkt/ecfWbFmpUHDbB3hh
OpMLzNAYXJPVbe0wHnG/Pg461sofH4dMqCGle06HCc5dGwmM9RPrUJZVYTRGmjubvn3GNMJd4Wvc
qzGyfX+olzbArB10baKktS5UCmMKvWOWg4HO5Zq3UMJ44v+2QITHRf2pLgRJQsaDMuSO+f0gd6u5
oeHTmp0u7kwlpuInsQlompUQ5JG9HB/ucLf1h4hr5/Xg6Dv/qu+lVwLW9BbvpeRKECFwkoZS+YsF
OF4ncFnFC00gR8RfUqWFCN8r9fF7BoBsCX3V1WsuFdgwLY5eCYszGbDGB3EHhOc2NoCuPSdZ4VrD
eCHEcw3Ggrw4VAhpCaxAMTaGiURCTw6wWagOxLHKRRLAlLy49OiDGed9vCoN/Md/h5AX+FaOO4zK
dGqzb/NxEszhnDVFmYIfZXFxhWCzUSMqw1j6aSR/sSYxkgIc0z12W5s+mq+BWHaE8KuyUw/UCu3E
YNC3IkpFKWKP+mIp6KGtMSqBRl2kXyEnIosNxs0DNz00dHMDhCNbT8ZCAO3quNDHa3eMNc2W+jGP
KlGC0TGbKq8ojJkZR/eku9iqzObWK86ZqQ90hI9dbnvGh6EfWp3s777LYm+QVFjaubMcWNcuvV0B
gd3fStLUNHiqa6QUhStRN8nUY99oCWCeMdHjrIYN0dmmC4uBIagiYl3qA0LyqLEMnKlYp06PYAnq
o+rGs6Fkx8QD6LWxauomu2J8QDBwSJyUSe0OVTUAxGPXzK4u12WlA3SogrhTAfBiBybap2R10Xsg
ombBCj0qhcIqrrc8WK4XonsBacDp1YE0cMxaKLqDyADRXRb2gCmy/cU44xv+JyUoyga0iCS3cOIh
1D9CDoJcRl2D17aoh4NUlg3wQIRU099eIBDapThht7xXrKPhxtfyZV29VOb09Vvm/52+TQ9hy6mn
mITHGtfgSUh2n4qdHaByAD5FN/fhoIklhAm0FrAbjIAXZ/50YJTZ2VGIItMnHeyNf8tvOrDTYH36
EUcZi2NrxmxJ0to0NS56dAfQosHo4P3u3Y/DTCI/XKkwZxcNJfdL3/VnFibvaJHecmrkcIR8o7v2
CAgKYhBX53/h7Zbqlw49I6THqEvaBpQPOqxUFI8YNZWvQqY5ipEdlw4q/zZSbXQOBj8+6iP/mdUX
GawYVYkDdax4i7zYvcN5n6MSnMIdsJpkFHeW0ZOgSUtz5H1BrPhAWNTrN+bGKFxuG9KYCM9kkzJ2
DkDl6U8FEOWB8xuZw1+Eikr8rF5PlzdXn+4nW4wgcotC2lDksTiLH+tqgUwIooYo/5nc8Exd3bY0
2wCEDEqDaRi9aiLlGkDwZlC6VSHaUKfLFtk8PkOm+917eOjqnsjOaWzsFdGd8uQnR5pki0Wmk2YX
O03KsrWXs+ZyYKpUn7gquJbVQXbOGovrXmJM9uil9Q/DyHr39X6X1HOSMs9Nw+ka+5Wi/JD3vwrc
dBFcysYnhC+twDzP1U4M+C7xyitEyDMhbYB4BumE7rZ7Ylf7R5pBaqomM9t/An7qs+nP4rkT55mK
7tEXjquxTZsbgR6DsMXt3CfE4qEbkoUC6hMAbR2y/q2Q1USjkuhFe+PXfWRu3z9iC+5N4tmn/6dd
XCvZHfdEqgFj4W+AbwGPCsSfXXh5cInnVqOR6nEVSAjONc7Hyq4cXZVmra+iuEIDRJ/8rcuq7HeB
Wy0DoigP5ob9frZPntDpRiiHUX6o/SI+qHEaFQqV/Iv1jSWVpsrSlAZVxus+fkjPa2vOLNgmEt2K
2QcFhPAYtck+iVSHE+bqRa9roSPmD5mV64vygwwyRVGdD+GMy3/g5TZsO2eloEkvdjSEMVWMLvlL
w3AakNVhg7kez+3rhDCFZfcymXDB7YU7+VFfXTVKLp0+znTfUv0vyWskWsocbs7F8SrTvEgeu/5t
pjitU3EQ8UWxZtLp36Y7QW3UXQi2/W1T+BUSgQTH+fPAy+O6WgAJcsaOA9pmwYMPn2My3G4ZRofk
I2ZUDS3XS7jYIN3XnmsNaas8iR2+LeymPWk8RBLtqxfJi5k/u5Z0VbnQ/O5xk69jPW+xLZE9mPdj
65+dVUA0HREXQMO0+lzcMeGvzp4eyV+JGz6XlUoMVQ/uwjA4odbwkKkjyTY+tvDiSHbMhS5Zb5TY
LPJ879HHZAQDbn9cKP8ZPPv0xDtPMOv/L91XPAI6Vl79W6SWyt1ov9MvcOyU6SYMPPsgNzILq0v5
CJJql4r5L+7ADl4AHLKtEOZEnrof0IO0doxxj1m1zauWljXyBmZ3b286T90rwYBfKpuB9XTWuHix
z+RCr0YeLmhKZz6cU0YLAhbEdZo/BVDzD8ZJb5UbT2DB6Grpn8aHKkyxXRHNLyiSip1KnTeu6DxY
BE+5PcFZ7CCIixNLFOFwLrRa9E8soSxO33jB4t8+uv71wox1j0v2ugMwW4LXhH4E3JKj8MJ3mD5T
XJglgsa//sZJzLTvOLMkmgCUxdBcIin0kfxje721IrsdxnR3a0XFgxm7g9Hn/gy2tTD6lWUOYLqS
QSirarlE0H7UCnWROgj94EmYXV1yb/5Oe0Ku6PC/9kXNWBxDOXnFtloV7cVNumD8rQr7TQpfddpa
WfS0tV/KCaRURuwT7r4jfB18436VeCpOSwL6YTgXMWlAee6tIioBeLYLuBte4a5oAn1AjWHFi+KZ
lzE7Wjq12IItb5YL//679ThRaG7moS4K5NaOPtLS1kbnpqw1TZrsHCtT/B3wJuyqQ17OTq+LsO7h
CFBButusiMtA4uSFcY0Wmh5Hc2vv9AlplzrnZ3Az/dy+AFbNXJRTg7cj+7pBGptxGlJaeWQ41Bdm
c1ZuY+7G2g6ZWgWccZNXQ0Em5qxLiRrWqVZZFDXnR5mfa6Vzi8NKIMW7P7p0/9RJmfbcKqqi6DAm
ecJVsl1KJ5pF7Lm/by+Z3UHqXy+wk/ESA0FYX5lLaBKKleHzl6UuDLUxg0KOBs8YaDStsI5cx/XO
vkQkiHnCA2hbm9EAQkXAPUYQtGw8RwBAIWRnEpEQuu4+FVLE6D5frD+xiAyNcY2V3WmHLEwjrFK2
W5Gm2SMhyoXDEDG1wP4iJYeWP3ji5XQc08Vu13J55i96ZT2vH22tPsHDiBEGziXS42sdhJ+WYPVA
8RRvGm0MrpZJcBBycWbFdeK54YAqAiePU1x3r/Gy1xds5h71hdIaKSMIamvUS3CtdkA5SIsEPzOF
scY4qlOt7NmKjPVB3sCT2nQSx1maElgWwXRXkiseHgsEt9sePqC04tPKyjA6FiFq9TW9YLUNmcQL
9g+kfsvLtH8O5tjREMeE6KLCNM+MLS29X9Z4yCcgO7JeSOHMjLyf3E4lc02qmiQpV2Y5wj5goE8n
vA3JAo+in48C5JEJxfp3daLF4MWhlHLRUaHPZtMyrD8+l07zwE9y9j/b9jgx0XLT81x5NeE2r8kP
PBbW20u/A8B2Y3etP0aV05ataB708r3gVee6f5AeDyPGFWBbbRb99kyEQMhsOHH6bvLLabHo6gS2
c/+L4rLQQIHo5B0nhv2+q/PxmT+HbXcMutSE/dBdTkFfmvNVCxfWpVwWtu6APsaBCIEYX93BGSyo
cHGyvdWIqYRTGGYNiiL0LtTuv6rQ89KDhy2eUB+CCi24HbyMppQmhhn9TtnWn3J/hWqoFdZ8E3Mt
AiPMTGal4lMcgXozrrR9m9wONOSnVvWXwLdtsEprbKFX5fflTNl72LSlQsAgcL0o78uBrzex6FjW
nzx9TUSe6/ORFxC0FtS0ofxQH8lCPD1CZudOr5HmsEFVQB798pWbe6ew2sz9+R+r+Y4yUL6x/zNj
JKBoAeTz1Jk2dQrEtUlVOjIqrc6WU71YK3HnsqgZ6WqRK7CPxOJ3+H6813rCLt3hd784TW1Q7SYJ
jBIiGzDMfMVo51QROVz+Jg59O/6u0s6xJ2QFDC9YHvFPAqEvCTTm957Yq/wabwLlI0N851g7xNjB
1nFx8SRHMze3Ev1ZV2srZ0k4+r5blzaGL3b/va9+xZTKL9/bPlRnpBRx9D7iW3xa2kH6yZ6FmZuO
0H37ey1BQZXa3vy3oplMYKtW65d9P9XaP6TyIOD1qfLHGdFAkZGc9UL6422NuagB4OPXs3fCDuKQ
gvGby4UiOOJLY7ExhbP7D4OZ23REXFiBSti6sLUciMG7wq2EOLdrynGA3O276OaLTPNOW2IT1BpB
vO1C5d0u5iMU1LdezY+4mn0bvq160vB0e0jsxMb9nT/R3yPC/LTcB+sa/NHnwQmpcmD+rc3+U0H0
tQvglmzkHylwejDTHZL+b1Q611JMY5rKUPJssttNMpXQ0VgUj4f9akXd4DkXuJ9qEp2WrIzPTigM
bl5E3GGc4aVcVXjRln2xKg+SKsdccd1YsQ0zRe6TYoAQYj7nPib9mAsneXTSHWWs6yIUP+s/hQCT
behOaOsGDgGc+pPT21OfducpaQWs5TWPM52cHQkqPRGQZ251hTTfAf+l0n2Z+hJUD6FnOSOwUbMO
ChhGKbcDkDhXX1tqs8ysPEz9j+fa8mnPbpgb2V7X+DKSaHsAcqEJWM8rhKdCnP/otqS6QQvIEXD9
YyOXArniSZlMi4O5iZ+L//fHKWR88PBQfNVK/4RYZ2xB+OTxdmOEMiaQlu+KQys0EOh5WIGWAzc6
gUJ61Jc2bGG06IiGf9k9M2M/wU/tPoAStP4e4SkpJSyLm5LtHS+m5WOmO4HZkLuBws7UV9axCxCP
0kYl+h5/w1YCvvklN+Yu0d3OwJ1+cIU9Zh5w8HdkynCGkGYgd0osgKcPiqb7Cdjz5/rE8J9s9xih
jeIf9N5lkv6JoYg/gRD/utU2/+SccJqH2lHb4CXPWQpJaZWfCkX6zP3cLKObLgvr2KN9C1fH+s3K
ulGx3fc9AdtO/miMGF3/B9/G7ZOkbgJfJkCzVZzw4SOSqiphkuAkyMmfN2GiIMaUK9wiThqXNDEQ
ttOWT30M80UXQWPzmYZMBRAxxwQrYdgzCmxOvEAy677rJdFdq6DNYwjp47F4S0vos0zB1RcbmbPN
FbGiifVBMdIIt0LswjiKKqy0BbnK8dHP6dA9OsvgA32svHAblg3CC8ikkHSDCx04n1qyUq1COoAZ
flAQar/hudNGhDY+GJVk3YGAnugfmUrZi8GhyFE/34G8ZUmbVWMjSjjnGXBeCC3dnbiB0vfxYDID
7TOCt7dWl2hggWQs25pn7P54rv/qtXassx7vhB7N215q1zOr50p5rXIpqAOmJjrouJo+WnEZvTqM
a4P7z00llv9JlyGfzagVzehfueB1b1EsskWmXCkvMRYOzsaqOnG7mfpz5gRRVWcx559nTsGQBrnW
JOZwiuyGLKsu1P4ANMbrga5kMZixrQ8uEHhcOcyZ8QHhOBEbbGxBSIk7G3+7F0vOCD9VNZcjDxfV
4V+5Vx/MwYrIBmhmu+DAwyPz/V0fHID7FAFfnUvOAHYFbrNh0OU3d0uugpm7E7RRdsU8sDqr7Vbv
O96ncZLq7sLQYioGdmYtxWeJgPKRl9rkXaCqcK/qVfdePxM4DbenrWefuJYTiTsxVFka0xuYQZap
SmzhSk2nzFs0WZktqLmDRtU9R2IB7K8tlbRBbu+maVBYRQ0NIMAeP56+eWfeXnsaAiI1y89/Bkz/
Q0Ot+8EvKH2B6ZgJsPHHMGzKu0OTNk9EjIY0RxnXA/ZH7AOEPe7Rkw+HgQpAA9zcoOCLvK4Tjjvm
7oDG24rJjndNKOyOA8KUWmtf8YYHIbmW+Vi4eJjr1u82na/Mc4EbKteSOxDqMKFgrNvtKGHlwmlN
dK+6nmIhAqJuxKvtvRAv2xnqG349Dmh5kus+0ie1aDYWYk1OwcZeufhDDR/AvRgJjovt1YIfGXBk
g7AbKl3b7vRACuDAWJZ+EpeLGRqxpxcEyfqaJrB7K93MR0VAZhNbLLgZk9puyfFLPk5/3hx7y2ZD
6cFgztuXz3eJ11NX3flZP46g4gCHOQ2v2zQtg9Q5sv7icM9li9SbZdnjUlnnsizt9vU58dIBEkN/
+FUD9FeHC1RV1Qs6+rVjf6gp1i2PkxYJrrYmVCvkV4VRVrHcIBVDbe8H3USGpcsRO0e8yZDdnWNs
rczqRQWISsdpCbQUjiUWFpudZckIjin5Yi57fxwFUCpYhEc3NXPHbcH2MIxz6sV4ZYMcJD+JZ53B
GfmOMSNsaK9e6YV3a0yzMg40fVUdJzEz7EIHfTzWMMqutNcVo1bJA2DplFyu0OV3eDNa1iFzzOxQ
of0yqgnc6j6VHVT8wWcUhR1VxtrO1QuiEJLQyjJ1+ANwTdIMwcaTFQkWSX4bm66zVIDv+Qjb+Yo4
FVp+GUyQq8rXmznzOh5zKMBrwodIARHvjGdXLbuOlKWU64fAXSvVNGFQmmAAPlEY+qM34qsh+hKt
w92EXLlwXmRpjKtgBY135G0J9eBVihMo5VdTQMZ/Rqo/zK+MpeVpRyNVEBJyN+wY2nfs4w4AT4Pa
lI+XSszXltuAbI+2CLGPkPw7vv4zNpr6SO3yKL/9sGTeF8VyGqEofYHmax+UY/o33QJN6asKv/3x
J6rK15PCCKsflCOM1/+qWjkdi1r39c6NduNj/LrGqq4A+7VVTAUIQ31j/oP0IfAXZ5qZPV8R1rZE
vEkZ6wU+GeAyDdL9pmUEEwpjYxNv2wtjMmlcyhiVnNnHKL/vLFjqAlbw4505n7qvuLVnOqlw9MCc
7x6rS2F3zLEahQHXUnoSTQZfr0/Iwk5GB/wYku/8HA1gZ4xL/AjbhielpZeqhvzWFvF1/YFL634Q
9WSIS7OC9wwhh5MjxDXNB0krDSqpUW7pnSYzG52AkaJJSKFn3txIe+S2hqCrrV6yyRmKo/QMY8hK
foI9QedwgaA8c9p0bcKlugyt/oAueyWrNNQwyEbh2cAGfHwG+nE24SGNcBeCm1Jps7Y72IUv1xn1
+YWP7Sbg5hzvD+P8S6IoTOzb37f0QaeqmCr+dgUlvFEWVh1yEqLr09EQFAK5WhZm0gN7drSPktHS
oxELdxof4LpaMnQ9raidTxRqq6UcSRCgOBb3RXYDyXkjwPKBeanxFSxDx+LMNplCrqApJ8jYaOHN
Tin1+tAWKoS1G5lK6VzNHZYbOspLAgjwBoDD/7JWAPkNEHwqYKIorGwVDPvp+Zl5hOMe8bi+8dQo
8ooH9MyW+lPuhocZ/P1wUdEW9AES+6gup/7Ml18MnllL54g4KWPf+VzmRWC0w6LXvTmxpUSJ7Ylx
jkB+6EyozO6pH4nr1rclyF5bWUKUPL+LnFhy28JHR7AuEAm85aEfooSRdkFhJq8SJqPHN1scP2Uj
6O71Ap7SAST8WXyysdfBbq6X417g+i8ZclCIPFw1dR/Q6oLPhiL+btLRl6TRdnGRUl5ncANDTAEk
fHhAzLwpR3Sv36asMqaJXdV2uUF8bzIMoeSe/91+Eg3b+GOo3ktBoMmECKhxfCf44F8xUOs/KxFd
F6441iiM/I3O7UX6k6L05K0b8pvYBmdgasp6kDMkEZmF0EO8Z+aiLVTN3W1hmVAdDJYZuQ0r3MZo
FpBTLQqHPf+wdGOpAwRGwQqU3fD17DwXoeGHny5SUV/ypYN6sPZ4TBDHn6Q7CCW+Cq5YL3qrU6oI
axFY2THT3fJaG2ipbFzFVK1bGsWfvqFLrh3HHrZRO2jx9S6xT8I6ngFbn9YSdSch68bmyaxJ1Oj/
89egnX1etf/hcJULQ29kVfWHf3z8hDqET8HTUkHm+xCBnY9QqnmZOkQUyqYvfWWTEnXYqLSK5zMV
oZAWrQZ8DolQSgUYCuq/AqWCORmMSYQ84foxlq9c6mHv145i15MWEGYJuI500HRz/5WGgVgSXYzk
A95MgiYdny1OPLTbFcqLL1Dh10m/lv7AESZxApeLWxNa1J9wRuyk4yYC/m89hgvA7sbVZRJ45/pQ
ySuMajIFlHstFx3voVN3O2h8GPhPT82G8uPox16/bAcr777c85bQeDje/t+AaRIGQNkLc19g20zi
7J4YXCSgytKZa0G54ppQwLuLXr3nXHtsNjGTUEtVdOtV1hzZTMztpLquVXZ9kz7Mqz8mCMAxSqey
NyKkXpCfGnXDJrr+IRf2qxDzcqzo3aVW53Tnx09zLXfGLGyViJqxst18ERBLCF0yxC5a+x3vsYuv
aW34ZgLojlgZ+fZv0EF8uASxuGRXr3cLRWFN5T6xtuK9d30U0CJjqkTRX90MmBgrvoxwTjOO02ew
bra8qvLZz6/hocZjFyFlWngCxKkzhNi7eJNxnkDwK72GXw8hwsurzotNgyUu7YJGfGFuh0O5ckLg
aKnSLVVNfRTM+T3Se0veULkWi1WowT/viRQjwl4k8uhg4GbYzJvE26DRHe4dtnpidNro1qaJHBg+
+yTHSttyskOmnWBnJtNJjwyQiyeAwFrVGlB+jUgEWrgrj7pkFmDTwnlVyRYB5kApuBzp6a+GxLys
weioYGntwqJ+y7molN/0qogjR0T4gucVHcZBa4A4j7HZPk+b1gfcCQvDc7nkKYiw8O7/wiReNd1n
4W0lN9hWsGcCpr9KmhKySA34WC+vNwXjdo4WQLlQReorNZHhr83lDHteA+TgObvga8fZbSg9eREh
y57iz9WQsADvba6aMkSVDJ8TgqN3ugWD6MTJi3XMbjnt2lPhmjpB/2qWhEZ4dmH4/8prG+wqNO2c
TL1tkgT4Sdx5cegV1X+KJWoOog+SOA982eRRyC5lftByLckK2osBY7GozYay2QsHUIymdom+ahhK
ic7ql61Qycp1ZO7baGjDhcVkxN2QHR859H0yHk1d8pCPy8hgSKg6alyoIjmQ78x+WLF9wrAcEKgk
VzrtQIcqTMnO3H+zY7Ndaynj00YPzVtM5RpEj2nB0nxf2/orFnVQCCfPvURv3LkUuNWGvvqtKyWY
q4kUPozhL9Nuo9jh/5ZFS1J4ZlORTWtvo0nZEqiMxGQm8rhpZkFQrVUL98IhnBdZRs7bQd8oH0mN
t5qZ93/WYDJiMM0mLMYb/GDWEVfhqJ8H0swdyoniJz9Nv6mAPZPzmvwrVXJzu92eFgdWBMPRxAkY
aJg2jmj1jqF5rTKmwoIxBrIrccDsJzN7eJq+9h4LPDFEVJhYjeZCpSd4mkBRA1rrJsF5VmkBa8mj
pPa2HuDEvHPH82HaWrslXwdji3oQAgo6OscK6MBTulCYn56EqCvD5Db+ijkZ7nFbQVRtp43KUlAA
YMkiGVUlxdKF9F/ffSV7X0854pXDqkkZDW4NmBR5XFmLz+fgdsX4igenpxvfFL4ZlAX583qCW1Nj
hp4VQ0upsw4+WUgFbdSqG1SGZVvZfNDoyLsybY0BaFVmJnfP5X2fpGt06LZKGkMmpgJUG/Jwkr3H
i5+o8N7S4bNEfYPKW+6MGGTzTIuQERcZDxzGtA3Se5mWoZiegojAPJHfUPxrSo35aXuYs47ZOrvE
MROvK7QvqFIgzabYv12Tp83vSubuCURQlgJuXF31uDKn/khvUzYWuvmorHdo7JLwXAyL7+wBX0QM
FElAn0Hn6dbD8m9/66F/odGmEG5GooLLjra/QGxB/kB9gFuXwS4LdrOk8cXNONXbnUKxUS5dMn0J
e77f/xcudJo4/osLn+12DXHs6ndZFFscXa0si1wQCPB1spoDXozc9qcrL+PuJJ56mVhusEj7Hcx2
uEtu1fKrYaU9b0BbFCODlN08AEENHVAFbOmkJevudz0tlU1daF/wU77qteaL/RZSJTNRDKguHnYW
880kKnjdikC230VLbHIYcpUHRGx+EDFn3sQPIGJ0P8HVvrnhmpmi5PJerRFfsG964cj25MmJik+C
uACsaizRul+Hgiq9R00mqZzcynU/Omugr7ORDNUVbmIL/DtWJYzRojdDQnewZmcTfMSrRAcFnYHk
o1C93tgR6t6QYi2mn164pAqFQ5eAbW2GREJGI17oLh/oBv7t5BcvrglN0bdvDLSEnEdhAPAgvHj9
Y2ykAlK7KFBf6CUnyJnCUKBQFQiC2W4HpNetNjeduHiB4dE/f58P25NxaQxAFGTNOtRaOqngpqd4
34ox2cUudiiwmfd/bjgyFu4lCifhB4CTMPapNLmhqOba4K6JE4RY9jBN3NScfUS7WEi8PWiBwEdW
8rx/F6FFUroa+S4hPgw3W36U4RAcU5j7sSUvQ/IHt14k6yDq3B4YuJmRDu5AFiboAqPRNUELO7cB
UvYQ516QDj+natsZ0Uh5n2mU8TF7Lxh6jOStumsc+xxNe206SEKqC3Nv6Cp9SPIgI5UkkdiuI8Si
9vyJdZRjXNSyJnUefKrDFw2DGmUGuIr4k3lQ6ooPrDKaBUexXswXTfQqIvghq4EuZONHbDwv432M
te1p0iPQ1pxMCS8i03+CvjFphdSlUqIlkRdcmSMNpGewGhAhETbK4c2Q5qI2YOLnfk3Sq17pf3wX
JCsbiE1CXii+JbobHG3ijfU8aviBC16tD5fszdohFL1LN+/NMtnQXXUyS/pnMRCLZARBGa/+Bzzv
TvsTuhOx5XZGpq7XbkWlBcwNWjr/PKYNHd4Gw067LB1AcE6uYCHd2oDPwEdOFE5LSGxmGdn/dr9E
QjDrIyhTvFP+Ye/AsTvMlGHZa0Qy/ygnwTqs7u/UzqOvZJgsUbVWZpqs4IW+39B2Q6luzwbssLta
e+dK5C+ZIC8gr8BM1NZwJx8QirG7vKns8Xkb+Rr4NpmV1T2SxO4EHCLxl6UuGks7SwXH96s502aW
zaY5z2orKXXOVW9QdDj97M3Zr2cvDADEXvM7bT7BTHy5jNd+umfW5BzLTDbRFKcZYQEIx9nPzjkw
KCqgaP+uCFxDed8BwZnv06i+8L8VyJw9hcCIIu89OSHPMXoOJjTxvfXyDYb1oOEWjmmDR+i151uh
Bhvelr9ryY0d1YjQdIEPJLdl6UzWibCroobsLEavIANiOcSOYvGjkVZhsRiKEhc1p+LfTjmtpMdl
lOB9dLYPscH2tnGSSyi4FY6/7KwxqiEGKWPJuY7F9OCc+1CSP5z3c4y4wnABt3dFy0NuvxNs2bIu
jOipNIHVWVlWTl7YIFaiIdppRb1KoJ7uTG9pG9+RlRHAwRfM1ZWdOMjiD23fjoXHKgWAeNtPE9NG
evWKRJGMV2sTrJmjA7/X8pBV9XLeXUBcMooV0FkMoG2wJlovWVvYOSxpp6ww6Eo+zrBWeRGtTna0
0qxS3EARk/O+hiN9+3+k1Y9NMcgBiyy5xm5w9ROooucfpkoQcBDum/QbYgV0alu/n3CaPx4B1ZFy
1KLrLZ58hi/fIkpMezl2PM7eITcCDXD7uPUt3uPeljLTn1c3HDcZm6rgoCMAuGK/sm43k6A+ppjA
uBTZhyDORCcsL1XY//+RSWDej+Ipdlev24Awzjoi/DC2xLV7F3lJPkwhG/FSAxOj/A3b9bv1fT9S
glAD12C0gLVOWC9hMA1uwUXiueZTap4zUjzs+drcNg6Vnxzbm8P3Z1/pgvcrduL7Q41moDNLdtrC
VNDetWrD9yzonZJy0T4aRNU/gP4eFbF/SbLbJ2tpD8Wz+e8mER3WUHisG/LchdnLf8WqT60BNU9b
UM8rbCxlMoexoXmVXSjWGtmJ9zVbUKgFbfa0Xajhtvj0ytZ+F0GuBR/+HKyB2Tusc5HiF4qqEpR2
b5GeX6QXUCQ+dhR0R66d0xoAg/CuS6Rcnugy09d4WSiR9fTg1GTvB6irm2xZcoJ3AoGVgGR4LftC
EJOZlF5J+KqKXXjTi5ut1RceQHHcbZ+bIxH8szoH5GUNWWj4w8KuRUd8Qvkxe8EFamxQwj4pp9/o
/hUFM3ki9CFprFB8KpXZ51HDn3F98KS1MmlnkF4aAQjV9//ExgZYwFEUMD+4qwTRtTDzfgivZZBH
Q5YI/hMo5Es+Jaq1IcPdl9HQBh+uctZV/MhbVkbFR+58KUkbP0JjRJVfCHGp1MMk+QDPBUlXZPDB
TrrGKtG5btHerIDMBdNuQ2U0O9BgZIlQYtarydL0DVahKxmznxYn/TY9uL982ZKgxSt1AfIQFPa2
jtLSYbFOiaDNKrBk8ePY1pVjv52LE6nzZQrBDSHdAdPW+ErsERgtSV/2fIe7oFp1VmHJF+ufEfg+
nZ43Zzqyb7O3We0kL+DQuG2m9pY2SoK1NuRAWFgGUOX70BYAHDwI/mjgxYQ57qqIhcsMe4ZXvz0f
UUereo4TSqiIcDWp3punHGNEk9VmrNz81pHbUjOML6KjbEDpswbJS5s3N7gXSdwFUoKWS/ZHBf3Q
MFDMUOuduGSQHm1NhvFMOXonMGXz8OSp8bdlLABg6d4bP3FIkEG73ytwvW86uHqTkreb4GPVnVEk
ztMIdL3Hoz9VoPiPgNeIr7HNo3HzGgZ2EQsS6pkkj1H/QI7WdayVDnJxMdXJDzKeCGdmLT6plKma
p/5XQ6Bl/l6rKZ1XXujb1ZFo8fIIun2FE8qHgC6m5RSZbgbn/aa0Mq0e1bJphHwLYEhXyVwdk3SX
4iMu+57YIRGYBWiVodnohAs1YauIwbKzkn5CvO6+yC153w13s34M564v5a2Tibxnw/Gc7+DKMf7B
JybzphHkIVjIqJBwBVYLRGD75H5w/ntG3CyA9LRSF259+2ryJQRDz8rSvLpbeeb19zA6YUNg59ng
vaykRbhmsmvwsqkEbk5kLC28RHOmxkD/kPgGHCWuFWgyJnZdSk5l79T/Leu1FzKLx24bsRloAkXa
VzcFKGRSysMOLPXO8JDzcSasIIzp0gpiocTL/L2qKoMPSIIHs0WisJcCUjXqsMmKe/85BgkhLI0c
nidW0AV6cT1EiYz8NhKczTuc6KvRB9j/JLDeGYknnvLM7WYSg2OLy/J0snKEcncJ0ETuRklNbgqc
uOyX3hJRfqsFHWhxQyo/0wB5HqcxtMK4trFfEFTa94qN25bCtKiKfxUEMZ0JGOpQ0RRHeDBGK0Wb
dBncCqYFJrJvYiJwYQZRin6YPuA0VqBWmVYm9gQ0wrIbtDBaSd4kwJ5/gbwWIy/V411ijiUjz11e
41edK+qGD/eqxNLcP6J1RIUP8H56NC3mrQvXrDY20j0Epla3GdBgsj+TKMm1R8R3fh5Ha4g0JOkP
DQkWBv31SzQ4YGkjHICVaov6Fd4JQrGg2UWk7u/mxl5vEmCHwfdpHicP2qCJ3wt2CV/SelULc4sB
DqrMV4NTnw6ZsEyYlcLADgjFMylmbuxFjuqQfRuu3t7P6HkcZOxawAfgaTjvqvlMh+96SD1iIpwA
kQi0pVhw7F5d0omEWSFGQUhzhJlY3pdAhxL/8UB9JEudOKpSo2pnlD9hP8w1b5b00gF6HrQ7menz
He0vTUe5QnJVa0jayKf31HO8PC+JtQ5ZPPokJzZjDW/Y9OYFEezN5iUpPJUGYLWrsxx9mZavx1Kj
U9sQ/l8Sfw0Qct/4iMSXHdUlnGP+2G3Yeukt3R2F7JFg5DX1aS1pVedT+RJOAfas6fEFHz7BYypG
lxaXcyIOqUjTALcRe1asb/rtmq8TlW48UfDuQB6U+Qe98WvIwZtlpFcROOclKkWa55UF41DQYYfD
EYfulH+k/1TUpd+eg9ZKQL35cx+6LHRsIS2j8ZUcUrIRhDRcntmbp4Ct8vIFUy9L/clFT9VMyOzb
EM1Zum+hcVdl6c1xgnROa8g/dnqz/54xdQiDzmR1nFZwSp5eWKbnH5BZg/zimvHh/6FaYtGAwQ5W
hBXxJaugodDQWu2mEbpv7pOHdhe/iK4KwjbrwiJXIvuV0rC407twga3AIcRchT1E0m4DWHB4oLlr
GublTfi2kROblrSVqqD0f7pQX+wjXzlrcoMGNGXBDjOf0uRmKkZCDkVZ2BPCdxB1dr+9QO61OgE7
5NsRi54WLkktXEraVGaoqvZ8TM1PuF0uuTzP3JgNxaMN+fTTcnly3S3dz+U6/YyFu3deFeO6kB6y
4x6gYe9AZlT02AzYZIxiufK1x48Irbph/MCaKf8m8eT5HAy+mKrnNhjsXYVdhEGK97rlCRfRTBu4
54MNjx8SffzFxq+lhRPciM6rLXTBF7sZZj3LG/0C0jvAjcENpQi/EnFXjRDx7K1MPsadsHVCKxOn
g1b6QcDgFcjNbPnYS2qLY/wXY/ePPC7L090KFVQxjsfHQmHp7sOJMJrweu9gDQU35S/OOkZczmnn
EPS8AOR5OamA0hl9uHQ52MjhRZGdzeJkExR9rwLZ+uhsXSBwyke5go8DufB45jujRTQZKTExgy0j
3gjryOJt4SpZB4S2g9JUxxLgsfmYHldKx8eQ5gYC5nnxgyNM9x/ITjAdMVM5tspH1YZ5yJMQCgI6
ktB8PbEVrXG9wR2PSJN/+sC4sMoVBuOc6nByzr33bnUmldOzBGLv2VnpdIMhIoRp9s3VsSdV9bNI
MZYR0GPypwoTx8MeC66dt9lML81wUO+bqvfx0O2R9bdn3ey0ocK5yaHiv+j2HcJrnQeCKAq9EXcu
Il9NeWJRUAB97EgPy3hbFH4AnQNdRUZl9EMjuYluIVQ6t1RIu5XtohCsK0N88+F2MIiNkqsFzaPk
lldAvhYO5HyswQVixrwbngc0rhjPKLASml4XXqRfhuQW9riZUq1CkldbSva52Y+VG6u+0g+hraiG
xxRK7FTJcQQg0nt3GmTOs3NVCFrVC5sruNfEEDqzn+OfdGxGSCYoGKBRsbzVapOxdWblWUeGRXXn
7hEuW23RGet+eSl/1RBzdtmuuf+3jBqS71Bq3rVMV8D1ld6FdIuGcmf5rv+KuWk2beLTtYytFTW7
P+32U3qazZi0ooVFEzHwvmFlyF8RHAM8DefAL9eG1C4HjscLLnYRdNTI8dq+hh9cNYraiumRrpuk
T/9a39uRNmEAUZ5hvOpUNnfyjGkwsuQH1zaSQVAAdK+ovx90m6dO0/n8ioNzIvtVlw8eOMoLzLQu
c7KKNyU+Q+uNdk0pXXCPCVZBxYHoOZaFMLH4l9BG+2QhbhkpgPqeUX2cA1Gf3szARA+Ap8iQRgJn
jRVyKv4bDHeUTqhyZW1ZvS3UJizbJNdRefDfXnaI1HiBWR8smQLnZz+WXXUDMGuK6n3nvtoaWyKw
AWxEl3amLy2uIrEWMIOZfFohpS7hpOfDxttFB+7/QRz/YxeD00JkFuks+w9+3kP3ybPfGKKC0xwH
spuV+SgaEMnyVZ8p3wI3n8wsFNuy058hl2gi1az34Hz30x63QMeG0L3kiCofFv0Nn5603Uj322ZO
5Xl0VkfD/KZGTVwymtvVzFoMxEZCWZ1hC8CesbpXnOqfmFPyViO1RjOdto07JZ/74MlrLJOFTgyf
pIkQZ2SIgQdracEXH0P5W1rnjvUWEKUcaCQ1x7t59vw5F2mPaJLVDD6vpugLbZPdClGFl2szuTTI
xVauRPDI8rg3Ee+WR3z89HFebz2ImyXLiGO5YsZPAv82tJsLOaUUywLCBoNDl+90UJxxMDxcSrTk
olHk750zUgyJHvtOtnnsqlksaqb8l8SXvU72yBICKT8YKOdhvutEs2fxTJd1Yesckc6XLaR+v5FR
b+11/rzIhx1Wmu6cdtM4vGzOXLvOxeO6ST4XsT9W4iGcwlUb6myZ5torXBZ+iYzoGyBi2COOU47v
QU11uHh0eCsKydFsOfxCB1J+ceueXgPx7NzSLlzUpWJks3oyvIkDHNtFoSMJWvrJwKP7fHubsfYQ
/2wNIny8JVxZhCv+ciV43bzUiDLxQ6gwbUFrl+QBgcIa7rGy6JiKDWcsU3QXFGzghrW1V3X5+/xe
o5pFFdPNDBHFfXcToUxnYgFATydJV9sM4yJjmSagB5wSj1xN2/H3N8e227s6flVNA19pA3ebnbhD
R0xrinl0W6seKYdaSiL/gdPpn2Q73jt+2HmUhCZeN3i8MKkev0A8GKnrl3+RWHmQWfQvHM4S9Q4T
pR84KW0nEucyH1FV67xtE9q9fFXOXK9N4DMavvs5ztbskEHG9OQD0ESo30gs8dbtiZ8XgV0D8fPN
PZ+DIInMqOq0MdZ44mHH+za+lp4drbvUt9+SXz+9jbLxgeiqis5dg7Xxkf52RIA2VlFjIUyitagS
MGOvUAURRcaQAW3jmJaNvL7f+4fduNGBh1WPeU1Dae+a+fNkPZuAfge/FAdDL2fZCVBDX/bj6Lnr
XhSF1u2VD0zqb5Q9uCkKrOKOLWVooPShF04z4GSVkCPOiwQt9TENsjNUM6tKWnjyWauvczpg9bvY
QyRaz3x9jXPZupbC/BPrv6OHFNQv63AEuiEKlEqoz341E9MAVlg/hQH4KpYCLAXABEbgR2PZmnKQ
rcPuLn+RkW9EVs+dmhuF5XMVkhYZpYgYjvoLuAruekLG65gqrFsyVIsIT7E20qeGGKWIAhfHilyj
A6ccgWGFrZIIBaBCehENJfpRsOKhLMub5GRNjW4PRuy0JqAU6IqeGulasHszTXojb9qe+O7ciSe/
NgYTmGEM6SQY7Ae4SceJWuH/LfKSX92k2S1V3UD++dq1Y7pQPquCDBAo6SMahyI7iG5qwfKUTN0D
1RI5M82J1+HiyG3S88xy6R6pgOvTRnsjVxT54jVaZWvNaENz/+cQT6FzpeCVbmiRpzoIcI+0gQ8j
bS0qtmq+74PdGKPicrrv93TUY2i3+jMIf9YB/85SyzjKp7h5vr4iJmywnlmiSrKhCkK//MlPLhUp
mSD9OhbuHmrLGa53DEijBGHywU38F/wndLJA+U18cN3zfJK3DmIqRuHjPcbCg5EYE7WTbpaQcsG5
GM8B8RzrfqYFOv1bSBxFe6jEVSi4VL+quuh0kOWzinYMA4GlQ8smIOdSYqMSJpYH2pnR6WZiC8BV
8qTOpB7uFoDy+4lBLyvyQCYnnFLOk5+k1s4exr4VoiVxWiZUh6AFzZuaFGT/bCN4eaftGzk1uNHF
7fFeNI/tC1e0hnALjBDzGGFy24mHOL3YZRcB0V3ULnaok2V3MtI18lly3gL0SXniFJfvqzjpgtsF
ELKpvpJ7E4Jh4BFtxtXZYZdleFx2rUVV1csiFgQpcXvsskvVJMehQm6HlJJvFoONPvcCRXX19sd4
/oQWFc9TrYn1BA9TImxf/7CmnEtNqjzN5gQplByX9BRkfGZltwzVEFaVnFxH9ZOvWs9AtahQohgo
OsAf3vGJ4pB26vpnjSRDnzQgUDUE3d4IYUcwqubRrXnQlBTyMZDcdKT8RflJ6q7FVRn3rK6EC77L
Clzl9xSi7dklS/kvRZIw0ZJl9s9LxX555GhZyk5MPm5Fnkh32rCI23SUjZ1n5ZGPItMPsn90RYD9
ondCFxOzdW5reSbMTA8UCtSwzoXmSvbP0vSkb8Ka9+2pcdRitlNCXMg5wFGW+btWviqYaeZiuTOF
X3hBxNWvmJdgxTRpKz464+HxGInhWMtDd3wDFL7YwvcDw0ekdYuRjns2gPSSGa7+M7OUKslhqf+s
cYdwnhxaaYyvQVVGXmEjxraxAitTdB39QEVkFrR9MKVR9G3cqlCyREGUESxI3DIUZTWf0JR46Exl
EWjOdzXsGLXhUGqsVqPQuCjV+wm0ZeCM+7nwz5wbYxKGW3/65QDGnNp1WK5frQLxOU3RuqRTpekf
s8E+NKxWSASh2MWWP+RIardRUO2cLkMKCgJMM2GzSV7kYdp0idQbysTL1TUunmzSMQ1b/sFiG9gK
Hpn31Hwj4yLtsIkVnYrPvI1+3DbFBfh6eaGha0eDQ9wcxvpiALfvmsjzuqZvx3Wth9Qoe9F3Ri5D
cdmFjmhZQVCd+lnoh188sUNRieuoU7OZZaKfYEGcbsFCE5kpL7u34IpxKlbpenZrhIg8KPfZvlCP
AWZXnNK22mAbKjkhtFKq+wMTiYL9keQlpneFNfUszBAtSqpI4pxf4jmP8ivAWyrKL6fZcEo7zji1
x4ZS2Ou6naxFZ/CcX0N4YbsuMW/Y3Z3fNZNyB9zfB68tBL74D+A7fc2vdjt5IcWTQ83BGu3VG1GH
WzS4aKVN6Sqyzx0dpowqCo20N5o5donWBJflWaNJ9FeD9MERGkj09kJkbdenzd0KnTA3o84V1WhE
6lqE3N9J1jAW3kZ8bo3wYTIa4D5aZMO/HvNRkl/gx6A/oLFkXwUHqUE9mOgm6GdogqLIEU1EKvz4
Qx2VbzXOG4rkr7o4RvFVv3BBiOgQY7nZw/DlVh6yk6Xc2mVF/tc4mwjlHWD5Oo3NMsEm3wyB/nGa
daGhZhfDnlMdEbmfApHicFpSpVKxpVu0QNtRkm/p9ENQF3sCfzpQSUDEgbl88Yyzj5nxD5rFmSgm
Et8UhXnrVLqfyrBy300aZDgOH77iCwLqwIFahOShVYy/RQi10p9No1KpHlGhOgGfWsZfNhBHayGM
n3LoNNuQfBagBiH2KdZbfWrvKG//V5sibDnBEkcyJZ/7X0QyOQBkTzZeV9hfVk8C3bNbc4GB37O9
CLWKX1KiYKyaJ/oTh/GlaeGaPCevou3UcWGEbnyPldyrNLG19wuAYGkgBUYexSr+fJV9XBqN3dy2
48a768uAR15z7AbS61dM+Vho8kO8h5Jmwempb1RH3hbxkRT+UvTQiDMPWbNToSlj7qtIFqtHSPSX
Fm4q0l1Z7MfSE0+rXeJO2iVh18l0mEsP6P4UucGbQ2wq5ufNeHHaQSsbtBRZThEpob8sUBv+5XS0
HxVhyRign36kYAwSdtcG4HMo+FQGRPcrbnhhFeDF63Po0mRfFTh1Bi7CJWQyAH9tfslaO2yS7FKI
BB5DEFYQaIiYHX6h6tj2TcgzvPAM136N5YHKMK6LFNIQjHwS0+iCFu1iQurpNtBhaNL0p9wERSMi
6Uf9eL7EchnzWDBwspp1+ZmxDQsVqiZGOQyKxjae3Rhr5Nel7yl0Y7r9SrpeNjAp+LX/X2ZTvuM/
i/N7PyZFP0+96OgZLdK6msYF27trk1Jw0Kv7pdk8Vx4LWsXe8cA7rtuObL6KNoSZNiJEQksTCgM7
nu5wEziTY0ubtRKEbmogKZ+nNYri12cND8Gxym97tZti4SIpBE97um8Ogl6qYGQ0ObpGFuR3RIBB
Vgz5f71TQte44Nb7GmPqAxyaW5/ooqXg4L9eKo3u7lQASOVH8p7vegrJjoxHTVVhGLO3bePSf6Cd
vNZ0/Txjon2ogp0miT5Td3WTsCmIMT7ADdSOfrL6tfyXFbkhYtfu5Uj784I4KNV/Goi0OXgpFOwT
7slLQKSbdQ5gEI/DbbBSIIoC7IHO3iC+JOKEtuvnxceYgDxlWJLWbux7bX+Tvl0eMiOL7QGSwV2I
Kxv1NOPXVEU/PUlJdFp976SVK4dOxhscT3Qf1BHotXsfm6gZ6W36qsZPPkPXVFxoFkwzxKoMRFMv
2+M25Ps7JtWdmFSL6TUzHwLiBzA9DFVPk53pPUhatVjmP7ONA3yY0/FSikdXK3ff267bAED2q96S
vUGYnCI02pmxg6PDXbAcTOLSpFGAR9Ak0I/+Cp/b+Epn+C7MBKCeZ5HjqYCXCBdcMueKg/BlrXyi
8k09B5XCt0m2XlptuhWbcu2cWEHb13YKRbB1ElfvwYtTNHfSfFrZ/m4ww/X8jmlbPinzWCg2zAs8
HL4fRv+ZA4iFK08suR3eqML2yRxHGPwCIYbcjohuq08UjH6eGsIE5Qdhmh48yM7sJ1hP8q+0ph+t
y6z1/Rw91DIacrJOlXtbKIY0cP5+62kfghfLc2L9j8bA5pEZ6y+9sjC2SAs5mWX9Q7HW5Q9JdSWk
d1QQO2K3XCcDrGXCQruDmKgThVOwmQYSePehRElAVetz1aAdGqGaK+COuheekhRzEA6LLNmlQk/w
jyJJQnJ3IzL324+9zCEWOJLMyCMwsPDBeoEKtRrlEUin+JXzj9ivrFJA85h+5zppiGhXNwTmWWAC
KJMpg6y9xB9d7aFBS5EEzgB2EvCulKM6SxRwh+xMFByWGsb+NwcV4T6wTHY3n2tfl5BRtcD2vR1g
dAkwiSJBEanZApg0OtTIegCU+xeSJCvPLgsxc4Hw7cFeAQQZ72VnZTKjOkhzNSvrAtcb4Y3jzf1f
tkChAheyFXh3dydB8Ic0KLKcIrlr+heDaN1zpelgeH8IuwVbhos6Vx9jJMaM//ChV2uBqaPY7OL7
8MgsTEiiHPp4Qr6sQ0APFdVh8as2ABSvlSXEI7FEDDA7ADIfE7Mtei9vTu0UAuFyEutq6m6v4ltX
aGVUAir3Ef98lrBniSR2QyK9OfkQ85iwMjfIeVQV6dpXKxvXKiSwu0stuY3bHnre76KEIXeCEh4V
Anz09vbTAuzrY4S6KFTdokMI8RtCVGzgCg76AWg+hZrLFwN9BWxoWvaX54S9kDbMrUqjLu4b6O00
l1eHjEbq+rvD16Bh5jGFL8rrzftcYVCecr7oTwV3T0aJUMUfwQa4zQoe0OtlsUG3fu19lV7eJPxV
HmEhjvNPOYVCmY7VEAyPg5JIV3rDwsyXo5nfej/JspLF9B9JQtnuNTJDJcQFRiG0UvzVb//fMpUl
fa/wMuTUrV/tt6GvBu4lSLBNgLQiIAVvDjtxVDgXJ+ZeZEUFitrpTzdA0SzO31TjpKDXlqm12ics
RfAoDkJr2mPdKCIqx0jRwJ7khSLTuikFjjFJ3KJ+JMySbN+5z7HxpCgs2+eWrfKNtb4vdkRRxteV
wKQzpU838CDpzKypB87WMWxGvkBXlW4Ll7uwtLYxnwFAi3yAJsNNBomsjnpRMA3VnDVwX0AfkKJH
YU53Is7ChYv7I/2j4NJlZR92vcGRHdrKSJUo9PpHcoZxYuxW/COPK2MV4CPUWARbAJZSNNF4R2LR
XE/wP1uQxuFiPVtINENDJH/U6ikiig9xtiEOjG2KrPOPyImwfPBm3coMraXB7bfJSxsbdDqEzWO0
lg110wRQzeOi53iOBuNUI7l7Nm8UHw6SM/oOA0snKRjv1PQookTG/68uiLgEvDSUofM1u/gS6mB3
htIX99oj3ukdfcMd8MsXyEspBMNuJ5hgWDolbEsMqr5KBJymPs9Ew2ys+iIWIkp22JjHakkP/B1Q
TGNPybOXpOzQeUhdE0nKOo+f1lBDyq35pKapCB2eiefxir0ACc656W7XMfNy0GaxolvvuHjv4RCs
ZWxEJw27lW3zteflnlhwpx/iYbzmSFtwfO6+/6xJ82R6lzEbE1+rQ2/CulapemINwQwsaLdTbApp
POgSeJ9+JICisBBGQ6kfFGMRWEJuVa/IHx4qgFioH9BJk7XQFnImxiAbYNrmads1ZMzYw5LBTjVd
x5cAX1J6Mnhneu97L05+9p+OPwU6l9GCmIEiI+RQEOmp1fQcIjNcjMpvH7VNIGvHVkk6CdCzz6cx
p7hyMbQgyS7z3J5KxCw8pEJCj4uNKjA8WdBUcczzHNwr0xcqguRIC2appZGF6UQqoNbw1WkmekMv
udhCZC2+UqGZj/67rS+q4vs2Qw2PhGiNyutsruVUF3rMSG3Bqi6fwNQlzWRTCNZyd+0afOOug23P
Xz+DCD0mZdWCLrYFioWj+78Xnucu/nI2VWdEPSBae6X47+runPU/fRsdcYcl6MOlgSKrULXoiUeG
tindGsPMqW4r18QivZxjjiOyuF4BbTHOO9c8qm9Die4CieSFYoY7tiKUVeSmr7F9WszaM4gdZhaV
+35j04NugImDZjzqyafilEz0sQR6LkdvHltJQ112z6gwLfdK4qSa5hIpGP7yQNez6pCZYz/U9uaZ
FkWdHjVqKEK50abYlFAiFf+kQNKOjFK8/6Lw90LZrHtK72ZuOZ+k5/3mGh6EBvmPH9gl/nns1Apq
M1P4QPA8oJnzuCS0ONHaf3xvDPjUW5GaM4lZ4AEuyLNg1I02e6CnQM/dvGpI6cZUFJJ2jXGsTmrH
NCyByCHgop49MZpPf7M7h/zBpJM1Hqsn8qZFKlkao6QWqh242bApByEVBdK4z0X6dZq+j7qb0A1s
GDg1mlxWaJPk53HP/uR60vbOPTPxuMEFF7+3NCmWBAiHw3ix2V4H3tpGJeO1T8/ISDXK2RMFyKy7
QzWmWsK4dEdQo7QWYuLdR0DHt3NEmC68itGf0nFfdXxdlF0Zh2uOPPRTDCZTJHmZAN8mqDyWIXBZ
AUsoYG5pqdE0SM8ZLfQwtbgA74VE8je5isU2tAOcxu4FZQ0jkwkr2QKLlXh/KRHZ7wrf8ljES0MB
Aql5jILEp3VCKNpR6xMHwFfgd3hMnXVSNFKFt23ReyiPvtpivNHhtnNs+ICMkPH6P2TKSao2gRvB
wK6e+zbVrpMqhI00G5gCaNdSZ9ZImusLdxw3HbO+8RrLUuh3lIeH5FeTi33bYRqyEWTr0so3c1nA
B9YRTRUdHPfCWXFHPLg3qNhJsJwvsH0uVhH7T2aB98mkgjLi+gWwEwA/UxUcsVl41Ne3XL3CT5la
neq6jHQsC+e90jrLePlr7/PWJH280Un84nHwSRhZ1TjOlGoBw80O8W1Jpixssl7i1HG6K5PNsiGM
jD1yC/9B1djrQ9H91+HqtYWTabWQ6/GUd75xxsgydNG1rIkIoddKbht8yoQOEZR3fiELcMrAi+Mt
kvVLAS1yFFuVPkVEVVClWZyj0ZldijRS7TYHEByo6IK62F4SZNoMejx0xqEXtOxt1vt/nni2iTll
CG8WqMhZW4v1wnGro5X2iXQrRrbKqqppwyEyjz8LIThdG9iRrSLjDNj3ExxrCsk98+6JehE0MWRL
25ZlL/VzwDdj0GU6Lw4o+owRXHfSvS7k13LebzBpMBo5orjLGxl98jZp3W5DYRd3fumKvR6XueJo
hAC399iH/TL6KgKUBBXrj0BnBjUywxkr0ISVhN1uAD+w/H6GV9r0jLSMbABODzzdcyYp4yy1Kk1J
07gHuTVIjXsTalgiaWR3FoaHbn3Dnw3mfRZ0vx99SvxZ8aRg7jF69knASMRsYPII756AyWNxWsJD
465EIGbAPIcu8+MZUcvlRnORKjCBQUUS2h2VPWs51ufnoFmCJS2/T3yIb71ZRO3TyLJ0E+tX38kv
U/g9q81PkBMIFx7zhLZbKBEJbLlmehgI2MaChLcxX0rvPwin/fCwvftU31YmDvrHWy3O6NWR9jju
VIe7mtQ3+Y8Hs33+sEWr62FIbB2vsP5IJvAxtoPwPtxh4LuP4LSh7zPlJWcEQNaaT2pP1Oh2F/QZ
d+PF/tkvB3mFN/sN+vOUNrelwntKKbQtPtkSzWMMk/3UAtMrODzREo8f0JUqCguwc+MCE/wjqmSv
uXeTKsbblQ65wRh0wDdSH3xWkPwgDxTfAVR2o0jbf7UlbN5Dr+AFmFz+rqRRs4tIzEabhgIVeRSP
hr11W2R+WOfjmEWhdE2GDNU++4QE/7saeubpZ6hyMOe1oad/j0/H2CGFNtsSg9J20l4qdTLK9fju
ZBxiQLbqSFgYPIwOv8fuLmiyKpgFcmFxpWrUbc1GfmyISdAuzra6wm9A9sd6A+031Ce80tBA4DBA
5gL/FHh+NHPYWSs5L1QC6jZXwI5Sth7gRm2vrk9dpon8BPwZQiKvr963a3tCJf6rMFK7TpC5xv28
aWa0nqSmjORifNj8jCCkiwaBeuW8csfPL19QWCQgXFgh/6tDdYE7Uf9QZjTkhHs0SujdVXcWI5Jf
lPxjw+0Y/ZRjh5RxkSsqBVJJAxJWDHi9JKXnV6YCTAMVfNco27D1GbgZlehnVzUaOCc+eeHWUYAa
DB3x3YQu4zDpss/8k8VAJPrcs8tjTn+LVTQpucV97RzawgnFdJRVgG8CDKt1jSqjt6hwNRVnzRQp
YxCEUAUZ5kkMsBcm9RtxjI37KlT6u7vj0RXdMXeHfwGS8xPPo8mhsN4K3QpC9KfpTUSkU3KhDRcL
uFn53hvWu2oFw8eoTIBhDkgdRHr4ZMDb+/RYbvwkgtWAuone31dPXW1zNkxgO5c+32nsYTjdQUsC
sRP0JNpsx72wDKqZHilIahMik1CpmwH4e+2ljFgcAcu6+IfaJL29hQMnRCv7nA7NnClsEoX+WBGX
dGfz4LIAuAQoE6Q7SSbCWfspw0rpeHJwWs3JlmdUYW+Nr6BY6n3ZYHXi5R20dhp3u/BaEufOnL0c
2TZlL9vQ2tKp2nzgnPg5FgeriEf1Xm/hO1RSrKnOTR8+s2HWSPmj4JKU/zTNL4C64+olRZAXgyCt
Mxf8DPqxd9oK6OESjJSlpZ6tcJr9AYlhvrUMwBBYTsCXRy47X99bR6B1yvb+KgPRr+y25+j1vDkf
7rZd9qCLvAvZ+kYe7dch6a0GqcYs+f+WAJ7uicnuIt/K4OGSHoNxWu0S1douSiYEzxVC4u4quYIF
y1Sm0F8iczJMV15blUchinSZZ7fIX4+B7qOTU8vNwZpc12g00HvOwFgNJL40U8pu5uFkzA3vDtze
BAV8i3Jnrrq5k/P+T8IJZcPtHEne9EpXHnCoh9hMBBWpalnWLcj8suEsC+e1qjMgPIfVKa4+QZ13
vyxKHOiCGXo0Ea/9xv7sKnSW0tOav+P9AEgd4OtoI7h+NdRQeWON5WfdIEjyHFR8HZfzAb5pn4/a
RFrQoFbcFpdIZc+yg0gS0/kBwI35vo3cB9EyaoHnJFTLBpn8CwQSGVR5K93N7LnNVYXEm64Q0rIj
fg7iBP4YeRnn/jBbR2DZ1/ZpjOf6px21hYMapzOC7A3Ts3X8Uj85ULLDt/B788KbPt1+SYUda+fq
4VLMmUQyC1d40M/HFT5GXY0r9ItYqoDzAu68Fi9ixtjkAJP369oBPI3/11VsVhSNPMGK70dX1LDp
iXiK3wVF5f/vMPZPbPH9NQRP/oQHFbjUmLedOUGpbNTk+vyZB71khi+0kZAdb/b6kIMoTxu53Ftd
Og0maSRixnZDcqk5vG0Fxtfpd5C4Y44Rw/hwswEAmwG4+nkx28rvoJArY4a6yLkOVT+eQz0ru5qL
vs37z4RUiWgSG7OOGtqacArEpZf9O/0oPWdWs5zBKb3cHbESzZSnjZk/T/ukUlPKGGMt+0FBL8Im
4IRBF4BbNiSP9ojw6UccIrRnMxTPwtYpAzZzthFKNi+zWNbTSRZ2JXusQO7fUu1Fu8xQsSzp6l6Q
i6v9WIu+QEWgUUL4xbc4RI80IzAML/kjm6Y5H5b/RH6gWzs3C3fhYXZ8lSBmEKqCq4S6A6XV5/aB
VflktSPdhtyCoe64ZDCX9T7QeJKrTbW6NJAZ/lRBtORULTENUsSuqw0KGxXDs8S6kktqBK11WjEa
pePGHIy9+EWoAwb+ay4IMBXKi+kq5Eho3fSc/k6F5rCkzs6kIc3mhC7blz/tsghawiSaKx+1tP/P
zudLyR2Y2w7dNXQjovUdC/TckWCKIllY8ESsD31A/zv41sPu6mrU2RUX7JFEZqra4AO41SEyAOcl
Kyh3H3YEA6sMsnnG4ZNpBt5kEubshLi/7cUHRpR0GiUNzlTRytV7QQ5Yr8aG4RfcKNfp0iPoUrc7
UuuI0pBXtj2kZTcCY+HSU5G54yDEtMPBLU7Evq2HiGCv/PYFNCYfnyFFE5+iY0UmcMVbeh+JH16v
cLj9GQJ3Ud/VnwGy7uUH+TCRCCq0/2bCfgYxSChzQtp/AOSpgIFHIiAuO0Wwp97QQRnFQfNKjIRk
rIOjoLkNewNNoSUNWAgt7TJh4z8b8YMztYDBj+wzZRiFXWNYt/MHI+PrUDULpn4HofuUIb/dpTy2
zz0X80Tn1C6haCJo17B7v1+hgVHsz/fpcgaWGmcN+498dzu8ffknLjqeJae4geCGb+Z4GQHu88Yg
SyqfezRX+OThpyqtPOqf0LjpGwyEWnazjsDN1ZBQ7stKQEJ7Q4glMHO7AL7odFG7p9CMVHNnA9JI
TMiroJPjV7HJVU9jndJH24i0D8+xn/7+mizT4Y2DMTnN0GWenrsrHIjyjdWB1ptAE+G9n7pwJeFE
Xa4IPtnKAGM978P79i7DhgLjhyYFD3Fp55x46p/3kbo6ZHmyR0Arl/muXBd2azlrdxYiCsL03BSc
P1MEF9oUwaInG6Poanf8hKUsZDAq9TV3n7gGWYEyqDCYO/91vEAV5JbYjNQ1sZkuInLGUeHRVKk2
UeQG7FbcEvMe+ciNA1kUkr+ATPY+iFZi9awF8qmjnPh/Nmd5Qw2Q77O/tjUac9W4jNzkVD5oJTXB
6FbMSfcM9bzuetHGdlIydwIPH7CySTi63kxKweesU3Tazk18rL8oGkoNOslSNe0JVma2eF8KQzsx
gc7QsS43rRfWiLqVFYAVSaUAqYojsLO8MFS2vPXLLJoEPclt6ES0Zb+ils0WRyAd9GopaK1Ix2bQ
/2+9Q4VtzDyiNJoOiKUaFUGu5vzC3BH+ief2Cl7jX9f6Y0x5ouqYeP3H8sPV+7XRW4PMFBPVMdqn
FgosEYdnXSDEOKOOHTD1ApZPe5zHc61qAlZVhzr5K5CBG01QTuqhco3ekKkMCBoRknVtdFCuJuq3
TbZUrDbKA2X0EYKwyZ/XKi9vpBG6EwgQzZIuHpY0Cm6NJEoYm0WLBvd8uTQiXla7OO1TPBy3F24l
Ck/OMsxk+WqVK8egU1qov3TU6jwZN/Qq1ZUWtw49BsK2AiQP6hJoyQPiiUsyhal7z2iXckwDP0ny
kxsQHxUsZtOZdPBUkaHC12ZefoDD4NzthrEYdMj+bP5AygX3fWwDD/5qKDk3RJq5WiTdgaxHdP9H
tHabYyvUi+6X/kT9G4qX2IiolvrRXxV+0WHSJaAKPF3v0RtUrpA3TRfAOZHTLlLYG5O6jc36jGiP
OrK77GS0eRiva6l14PqrETvrHMGKW/wUJwb7UJa5J5SbEa2rePIj0qV7FgnP/3gYtvpDVuUw/riM
ybtOQEvfzwVU0Si2dPz6SUEzy1UxaHIjcReEgVLKYJVHSKDWO9BZIA5PBzfVkN6Hb6i+Y/huIXrf
eLZ4lxThP8ALlVaaqfmedKHFvyRMz6aYD2nrvPQqh+/cEmzPbWcduH/zfIe73WJAunTGqEtvuXpx
krEJij6FS0i9/zv/tcJsXzEzN8O2GYLDSM/VKw2vqOl1KzFrbfnu6k62o5LamLb6F4QhBidkx9cF
psx8pdTgqk+Ram7dat4BbRmRa1ybLvQtdcdjURovzvjsohvWh2RlHkTeK+jGEwz90k9S8qdni/Ze
Oj1STT315FX2gvu6ROlfsl7Osc62xGDwPlvk0wMZ9XwnqFqdDBUUkDQZh4p/DWHZOPWrWw9xECa8
ysdt8fhEDRxwt69VeJ7TyqrNRsztQp9w7WHPMX2At26SALi61839jA3Y7gcG742Ibk895908/fSj
XQMTShE0pif0XirhVg/2J6Y1q/zCJZzy0a8zonbSSNtcn/0QeYDwFDSR3PWHBd1V98gRPPWtZlc0
X8YiqOHoz1//2gzTCEFFUuTGA24YxAb4i1vM4d+8t9WUvbJSbqI5bXxdFCjyZWjVVXJw4Yx8iI93
IBftkvAx6T4++5COK3WPke0bxPiidSSTUA02FOE383Z2wR885Wz5NFzMW1hQKC8InrMg50avasp4
QTLCq08teO01dVswoqOhzJevT9VriZwbdfDK9CDz8IgiB9AISsMyeCtS9uvq9ju2HlxKRshSqiJ3
fW6zSmZI9RqmHhgUjOZsp3/HKKH0lYyHnskBcBRPwEwUMQixmwwd5nPczjxnYFXdwCYkwHl1KNCz
AZgmSDLJAV1bQuLYIt8p8pLCoHxgQuHMhmBhouqYpByjxpfmbS/LzfhDBxZemaDWiKMuXjTLmVhj
Yx/f1deG/hbXKR5j8QK/R4D/Gy77rnRg+aZvmj43vphDCsl0uYKhqyezTH5Xe/kfahFcysxC+3x8
5KxHCheeZkrI8GKk2EOxUUHktv9DqQ2A3TuVHdGzkjI8Rm0OSBCZJrdTJXkAggOG3t4EzeW9Nf36
xnFvuithU9ZwRnrbMlScscqruHrhgged6iQC0VlyrGRf4y7EnDjH3VTWbPp2dkyxkFKAMvf9wt0Y
6ZVgXHSM3LF2TVa5c9q61QmmHAlKO/8P/W8G9NuPulx66JY/2+66Dnajk19hN75hPY5lL18GPgkL
Car79DRX8ikHMOOZvikEQLrYtBVXoaviCi+0xZVlXx7JiKdiHxB2AkSV7Kzgym+SApLYWDo3LuOF
6ZIM7/MSmEfnoqp/gC5a8DshOSXSJ+e64z2nP6sHCNCx/Hz5+DCj4u/kpASeVPyArS1vYgUiT6aM
KlydszOmas90EMTXOgf8NX794mWZiQlr7NpqOxi7+PWSBjQS9GyCWbXzhW8vK1t2D6Z/cqAtrfA/
j78C5etK2OQwdpXiDXCnpwOR/5OVetzMaz8+MGM6RqKJItHUORnwj7EgrcWaHK4ghwUnfoyulRdi
2L93DKDmYnvLdlpOWW/BAiJqQTJvjkY7nLSAYdWGk6U1BVlhiaR3jRO2PIKwnOcl6qHW0jeU2y8F
NCxvuH2jdojYisiZZMJYCEULjVpLdyOYJhQI0Bl+WuLx0AOTmQy90l0euCIzu9OzsKrXZl0L+pHc
hYFyloqr4oD20GZS14KwQOLKi7DhUKwvwCPe8WoF7yBzdzRKG7SaH1MsMvUUMYgbPKxs3XAmrsPx
7o7U8Uh5hCxRZWp4TFQh3UyIwcnWLIexBPzNqfK8XOiNGOUmaLnZObot3OgX0RARdMiFlA1vjdZ9
s7KTQhkpbbbF40vGZLUBSuh53xh16S/5VI4wySpFv/00dYaQK1qHus0ePImDSSmGCMjtvEz/COlB
SyyudbI9H7xznoSMerPrczOqh0577DkBCOzFgnW0grGeV8ulQc1pDHp3RwTtGciNbKMEaGqI2AV2
qULGL+kSvXndL2q4CVqH3qAPV7Nt28epc98NCUZZ1EehK5Sw9weO13slKivqYkcWkhVV1yOfxlcC
imJfNz/A51JAhDRckkHXdY09Yhi53bcZfw7r7yj/O3RyvVx/0YyZznyzZsnAPzHeAM45F1TqClHD
2xnuTjZpX5l1X/H3ii0tvRwOupXiE89MkAp0u7SU3Rh74onbK9NGE+VHUqNHhLZZIJ0+m0ef7r8A
XYO9UswQkF/6ZB1GRtZpaFvql3wO5oA0XUYWnwJ9MlW6iqtIbJFHOKJJCekRjEDAF/b0DqBWzB7+
5kd5ZkF9eeCnWg5uUjAVDje78BOdSmiA+Gj5nE5WLVcBsR/XpOGyTAMVKBJgDEcWIgKkXU+uypes
Skp7yoXrSKY5W/cFiLSrv0G8dwD1yk27bCj6QO7ylOn8Wv9p4IIkUERODsCWDoA1gGULZwMXyA7H
ST14mf6DmsmEVvRJPbhc5D7lDC+0Osf4+1kKa8Uuc6s7a/X9lgwkUHsfy4y7GZ75w/T8Q2/ug2Jo
7vSMkbyzCt15F94GHUcQHq8FdjHqTIYJFcja2JhnZ7NsBviBEG6Td3BgTVIkVPYoOdUCeCpLZCgK
u4qeyi3J25ArwknaPRJ5Y0sMbop1kKEm9W8q2UTOYNpkCZYadQedS/qIvFfcHhpcDq++9Pt4HtiU
+dygYTmKqWCyEaeZaF8dUWpEY7MYbiS92kkxAvt7TFgK17PGOtBuuGk5ePxSElKoMldK4qaU7SLh
vQWDGSAJUqIA62oOI9xPxiOFEdoW1KoOV2z5RwGbQTM4jy2R6fFgoUOPGoX8bd6UEsnIEJNfrYTo
ovDrwxHVTvlbbiH5PoZsm5XJlEqbhhgIgxjLaTcDN9CAuC8da1xQta/OscCt710Wd1qp2Nw60gvU
bnXniFkuigJlNnKysy2x/4x4WUTqzJ3peYmuP7IBPfkg58BRiEM2RE4z0GZRTx7SnCjBZv7A7lS2
LzgYc1l7DQW12Iz2hUDJyr7DC3i2t6pXKOKBW/kMkd/gZIRyPBt7tMYkRuvahtN/k2eL24r0HGAC
lgAIvHjzLW5vkl6B8iyfmYDZjYfdX0/v19RryN/hQ/OIuJfv4opW7tKAaNgIAFvWUqk2Xx6SuaNo
eWDvA+gQghkIpJBScnzd/L5Po+J6PrHylKTWZDccGTuCJ2sDA0cd20mTw3bgW4ASo1mrzY4P6gNE
5chv64afAkphX7wt9X5HlYafIDl0E47CHw0fKmeeyAqK8FV+uuIXppXA8WS342f1Y+SKMZgwR3OE
DAChOKm0StHghKfKj/1bHDeWG9uF0ZXSe+fkPUDrJM+Gex8dJvxzp31cKCsoiqMPs9nnJU8wYIjN
IKZYPH4o91wOXHsYw70aU5kGILT/W9tu4+MRzaK6NMSmo3P/6RCwgGsJn8kGWYMuw38oYYAml0iT
EDhusWuKQM1j3EmhCz2uVK+h0XYw+wXK9TgckyP9mGYq6m1jRE/bVc7RrQ4vLvq6I9/q860AqdZA
YxZuONZSzGc9gEprDgssTifLfAD7fSC53I8qgZ88bSbiTac2u8nR5Q3z3eg/DB7410PbDqToapTL
JXWw9MxqHH/ry+hL5dzLbK4egy085EvkMFW5QeY103EDWTDVO6/6gaIcW+D3c6Kv+DJKUTinmtkP
lbRWLirApbo7wf6Zy8ac0oFmw5e7mitPrZcEQyQhAxZbmvB/3GmBjpFjrnuJObqp1gb+VFbzjaJV
jxEARa3qxXrjcAWNpS2SUoXJmlhn9ByY4Hdq5hSNKNDst/tfIoe/YfOjJNaRQzSuPRn5dUz0Sy2m
2KIUxtoRyxN52ok+0mfmm+8jrUi5fUEMV9Uad6Hs5JsjnMgY31JDHPhsFVutSvU9qfzctmlqtEnE
5YKNZLd9fRBPSbnM87nP97o2yH1GwkXz0o5iACQyArkCegd9u5bP6C+1flBnyHnnG0k4UQOEYPNt
YiggWxZux51RS8G/BVXX1/Vp2eQRD8GUsWlydR4b3mA924UdtGDZZ/KDcbhidADYpcL8fC7mF7Tj
zv8yEaXZdVGJwzQ6hh1ud1wnyU+WYKyBfvpwsjCFhGoUnCyMAaDhhIiDFW9R1GAQOl6B8qyv5Sx9
sL5cPQU9WZjvq5Aow2MpbE+IRfbiFrU+i+P0Yndbe17oMC2QaylyiNJnhFcd4LXCTvpWCMIVECGx
K1K2zedCGHXxU87xQz1gvM2tl1Lth+8Mci7DvYkgX/BTRlVOmk+Wad+A3kNSvDw9YbLR8cxLSlni
1yfP0h3LI6PdbqHPXgDsXGh45wOGbM0VTKvL7Bx+p+Q14KT0L/IQnFQ3kAExghEsy9YGy/vdA5An
1d50jTwO3/w0AtZM4J+n3xwygaCKPye2U8mI7Zmn7O0odcE5k5mNLRTV6mRQgowBCT6h7RErYIWV
5jMMWitQ8DNDuhCsNyzDewP+yqgTSARej3JHvrX5DebK6byd72IbKRJZmd/Mfn3p35FalO31vHFJ
CsRmAk7jBQ/Bpljvs6mbK256KUJYD2Z1OH0V66ANPF6wwSBQK0OI0600rnRFTftB+InlFQIPDmXP
+4QTZM9Amtyxrf6ruyV6KB6t37ZuxhDOYxQxMbRPvXObydoslILQj7mnoy8TxZADl3b+BsTyQRWI
dq1fxPLNTnGGDQZUOSy+poszxxHf5aRtXiZ1YL/bc2s+oWWnYAiql+PJ3FVzvEmCpPDUkaVSN74M
ushRCFvxVREpmjGgMyv5SQFyw13LxHvoS48d0aYks6OyA7yfwOuaz0Imm9hxEZrW/aC58AzUo+VJ
Zhc9X/8LO5Tq3Nhg7XaLl97qhQqFyz6LRTxJKdW5HkMB7UCHOtLN3i9ATGiMuhGbSAFQjh2UbJ1E
wBfQyfA2+We9TGieTuCf9R5bAmpDvvpa3HMU/kkeLWeJgS8E8JYLOj5ChPgYlMZgMYg+ijtw6kmb
NzTH3Zg9MuIM+8Q05XEpB9p32ZOa7TBGnHrgJgBltCLR+nGeLUAzWhIxfaWZ3sqg1PC62Bg42MYs
76GermhAVs8FpN9BYj2x4fFuXV7zjNrgLROV+f7ceTi/e9x0ijD3YYzh9jrNkN5idx0IlQ1Ne5g4
8bbCksBRDc0waUu1YSadkmwQa3ksFtlZGE/qh5eifcJJbZ3LcD5c+PHFoodE7N/NmrjQY5QBfE7Y
7ypWQ61+w8n2ZH37Xc/xXO3FhJli6iENoPbWOsb0d9u6ImIMqScnBcdM+MrXCFSxCcao8f8Aa4vW
MfWlbZ2YZw6n1+adY5QPnXjSoPyALP+NP5Pnm45QUUFu1XxnZ+R1x/KbIE+Wdyl+7vxz9BdACnFI
c5Y2pWqBCtSkqv128UY5WkithCXw9oYgx/b7syNA8awDcKfXZfnd8olREtdacbUwp90wFZZZkGQD
TY+RpZIZ3Qh/4oEiiUCWYK4F4zDsOW+Sd0SYW+ASKW68/DoCr0w/rEfBPe3LPs1XlXa3UBbrwaw7
TbyoNXvGONrYevJiCWzFBaVUBGG2dj0YgFR5Pcbu4qk3TPaeFaWtBJV88uOMK9eyFkk3pr0dF4bZ
VObwKBrqrTOaR/dHpf9CvBZiy0TGX7fG00KoPPvLmZ8b9GO+b6h80Q7cwn5rd1RvKLex+TZBJ52h
ubukARawhU0sEL96GE4bSjOYF16QQtv83FxYgTCCqFP7Erh0fOSCFIqV8QptY37JnmQpx4127tq/
athhasoTU/KvZ2cly5NOo791ij6nY7tdZ/8V7qO7RPkJSzEFqVqpSQdCijCMEnRvCASygvtldAVJ
aN6Z8/TT0KZexah/xuInIjBdzG2eUGF0QKToDGpMIZr9lzRFz2dIKTvhWV70dP9aEvYH7zUEdYaO
WUwMYWwAnn2t4U6Fqj7nsBl3wUYtbMko5GfAFpes9G/wyyI5KXXhqp8TcadSSNsAxJb/pVXx06sg
NHniR9j06RfwuSn25JQIpIba3CRLbQPoMk1mskoxw4WhjYi2cNw+0hD3+CHEWpxixKebwpCAsoWv
yBPY7qx3Jsd71DrQdPceThyn6eKKYhynPy2FDvcmsEEDz0HFEi7A4rFAIKdWHsMkZqlqL/+RydFg
19lYta4zljbHHLLODiWeDXYJmPWIqW/Gl5Rhj3nhD0CF3q2VSrdV8IZrNXtscGxZ0IfPfF1OWgCM
+stB8DkviCFmt5NOEwgcX7vkVuwtmqvBIMxqdXEDkkhNqql7b7hbC9u8iKJPYOhywX9f+1A16wcr
wmF++hUvuKKywK7tdqRdG+wUihrCDR7G88GOO5zlb9W7F5IhumKsRZTIPi+oVfxE/s63sXDBzO2B
ZME3xn6HhrGCzDsGWBNOEMnSpykF7cgPQqGT52dwN0cU466HQkBAE/NJ2kpKdKlVVK0ZddcDvQA6
c/9h7X8GBXH32VVU6pvjjqy0motboOEfPM0P6ehMjWW7D6XpK4Luh4oRdr+1gJ7y3Ka2+OPPlSGr
QNs+l94UKit8XSuhFSpeGAvZbPHxA/rK7mILmgT42teO5ay0dYXMYVgCB+YtE3KtENxDrUgIFxAS
XkABrTszJPTpImupWBtCTemt5GC6gpOkL5YKgDGm4a8uhVy/ZOWK8fO4kRwKVMiR8duF/abLWabP
7dl+Zy/bKXcJ0sKb6ox8ddhbqy6QSPdf1zI5P3Ucz0C6pqA3NFXN35vtFkC96eHzR04J6fQblfZP
fHlm+WA+PMxZeprdiMbCXNFvpdgxFqTGjq0WJ1RCnqGk9tbNBG3BsLe9PcJ+4lFMjmBTa/QbqNfT
XmeyZOi5l3XCvSwoJLxu7oLgqUMhiun9VGzM5KWOIb9aWBCYyqeWXdToy8SR24XGUpdM9vr+7zGS
crNmpM8gfj0kj7RHHIT/0mJtWcjwBSe9pxRxp+fTH4GvpmHHm1LrvxLnpRfC8K5BGRITu/G0zTg7
zjVxp6bHpQVV7rouMJWiGUj+0+oMENjHrOnuN5gjUW8PvQPcQ+5eJ5YnIZed7MHVNAeJDF9MDLVo
jVuWGv/10Hz64PWo0B9s6rh+P6YD2hKdF7SEZph4RXJlpItYzhHhXCett7HtdCGx92+PxfhyHtQJ
ewhTkKWye/AoW8F6XHxpZqlRf+ajy0r6HbkQWaAlax5BuGt8xBcmLIWPdDNB40UZSZpS7E5Y+8PD
KrKuhXFVh3NUB2Y6UmCMwRoyVH353ee43PPj5NrfSQbTphguvScXfemn8pBpIAA31DObha8d2RFA
+0humJIspuvNVvm01YTa6WlChucp7f+Qw2y61inKODiasmfse4Kd/TgBlEOstiJXn99x/AC8Q0f/
KexR/koiDoQ6khCF3NrwZDbFYuu8U3CZwejoRPj4mZdccVQK5NGm9rKo3XFcXPlWusQjCPQtOPsx
BXi7zIiOI/E2S3hP4eXQu+m54Vv6uNAM4cr5oD7BFEcsbH16AjAka/AUmFI8DSIO+vHw1Miz+168
FYpEHQXU89FwAWaZtLzwS7CNXJoIKfrO/gjk24OFCm5vEKYcipIClJkOZg4z91lxmT6w4tNFqZKR
XVy8FEA9C3cNwhE5HNUB+OGmmHOEcLYh8ZLqBPKcBmO9OxEqcsXMOe6D18Z8DsRTENKQZj9X/RDV
xX9dc6+cevP2MX722sPPDZPYZq4mXKMwjnhPwCtZwyEL1uzhmrFhfIPfv5bVt2PZXr6mOEEQD2xL
ne1UR3OqVs9b9/rX+CuWS5Vuv1hYVCklemi8NlwMVqEuyc4poMd0UYiUIxuaDHSQiIszPPworF6x
JlQWlCa1x7bWy/BAisHjxJD1wv1s9bzdaKqr2HEohM8d/4NStL0p22ERUI+XxfQ2z027cHXZNvuN
/WEg9NpTg5S6q3/8ViZydf+lKiJSCF+tS02Gzkw/c4RL/pmU16kCAsKXasKbXmqSCsyQgvlCtrY+
DQoAsgUNFNgGN6rHuX4BEZRHOsua9DaunPkg28PK0BwItlU169IUnUqKIudjlNV+g2Qn/2lQGYfH
KvMiPgCy2bSQ3mqvaZIQRh61sPm6/tHksRD/DVfVCsWstCa3rTkUwnc5yIMy9bW2FAjitELcripx
nkHbUMu1VZJP6Uq3goF55/PFpc4eSXSUK/tx2w/xvG26LFVo8GWPbkQBAP73B7BvlENEx+uKL53m
xYW6y4/Twq7h9vojzB75c1bATye09MRc/0x9wli15zD8eYfF6LFV5E45f/NghHYBRpfEhUytwpyl
AEwIhUVDyw23cNiNg9kt6YzgbI5G+Oe4WmBD/bYQ/pDSQfrc14OIUh+87RZlmtc/Fg8OpJwuV6WR
EMfBvrB3ojFma9NXlRpLkQ/SR0zpJLlW+oGsmjGBFH0U9zrUHrP3P7N4w8E0tzGO/tA+MuUZMcum
eVRTw7KDrTR9g6AOa4haF1ZDccSiHDm8SaJTqMCWIsk1TS1AnmfqFA/+tyfVwgUA3l7dNMhlryy+
hHDfUgAc+uLdi+zZxlTCvOzZGf1SkDPakm38FrgaWpeh6JI2z3NUJuUUguMZYQMdNhfohxqFNPZ1
BuGUAZzaKo0+/VALG7oDDcfx541NNVyEqTh9bItJv0yagXJOhS9A/qmzbUnrk0sYtPVHcyz8VaGJ
mEjWWfXIjA1JKZf1n0qkR9u+c4OJLxgQky634Pn2TqOxL4M4JjbAF9xUfi5ud5gw1l6qv10vk8hU
Vccwlw5YKRIp303YRKUm1SKFHXF77RlA7N2EtOMeQoxLJHmeWwi3HjNaeQAh71UTjkVGeWpCnJRv
bZMTj+k/6pzBm+kHrRWHIYoak9j3aKzZ56XNxySqszXfsVQl77WRsrDe1BajUgEUdv9r34FFzQqV
ntlKVYIhsdu2+cDIyxw7+xEUxIZdt9ZNa0wQVp8oQZ1k0gL7NyCVISpeZefOPivoOjDf25bN7gMj
VaL3yzB0AKlWtdEEkppZkqrU28Ip7kyFJ/IXeFwPGf6AabMMEHKTaYQomElxM1rNtzWHKJpK8arS
HcQ11zQCyUrwTH+jD5E7YllvmcfoW8BC5P5HrMOTCESPQYLlVkRbNuPsTFsPQ7euYLCEyQe7grnv
wN5Sj1nWVXOKG4AEsAekDU08z/gl4JdxyGbFVwwd9QIxfYXymiBF6woCRaW2wQYI1KPk86VliP5f
kGAPlmiIA4fAfobk5F5oljl1b4IgLpjDtdF5YRVnJ9BxSQkDlrpqmK/RjKjFboF6nXYG/OJKlTWK
GqpQooI5tXvOgz3q9tZvqlc6HSuPKtdrJSGAoeSP9fkybB4cIqnBJX6hJOHcwUI+cxO4Pov/MQSi
87wLW7VU1CE8Gxw1sy0ShRAk1Ojx0eAKTPpjX/OQBacTU7rwdej+PjmrzOwjJJwAGZKUDorwWojG
uTzYruUXqV30J8OEPzqc3VfjKij7TwOsgt7rY+X/TDUHJIh4n4seb1noOiRBtTeQThTvJMGsAI2Q
NR94QqfTmJGarQNNDumXYYyar8dHSMpw6XRsMLCZUJAkjfqZA6n5pbVL8xEodwkfaah/Kuc9MuRe
mgY9SNOwN+YktzUVb9xOiAg4dHjyGBMUYJcJfI1Xv3Up/Vw+c2V2kwC6cGMDiYidzYUAlyXkMb4V
3X713qwLwneNAn8vRzCbTW/yHRAiCAhwMBqT7l73Tiu9UI+V8wOBlsWEJpMJgxGpal6Ti3nk58fs
pYTlxjGo3+WQcmtJjYRGxyzODikCfbechDouIaH3kadexkuaJxPtqA8mQxO3vGhwxUffrgQUkapf
jDQr3geD01jV/xOwVz1Vy8IBClEDFaQOBSng2tk7CnbGWoKRNqkDIUfj9CeAZfmvdSeAzVP9A6L5
IRuNKQbJPPOL0RPZl9bGUwYUBtXWHiCxEKUarrhRZeJKH0h//TraNfuvY4dYPuiYygfuc5Smnlze
5KrJyomlgGUTzXNolu9oP0pWd2AYoYuDi6LWPY8CudJ2iJmNamebYxKw9rr7WPdyOOxNATaFeK/m
mEvY1tFxuWP7HEfhqqq2c+2CaLIAFY/hxKXdaI8rV+X6QRnlk0fniek61v5D1aha4SPkNbnuOvCw
q1JC6CC5pYgfKvQztK87eguZAaXTOsv9tQLNLOGIqy7EuF7iemKbhp7duZMtiK3LGjSqViY+aE7I
odlHuT+bEMQexm+mUKddPBIokBjHGTq/GJGL03VDHXj7arjscpAtB06H1vPlTRIOBo+t0t9sREHU
RVoatakyhdl0bRWPhF4VMH+WDZx3EXUDDzNnwMLOn9+sD5bvaiIbyBYRbCozYODdP+F6baGu/sgv
Tc0e8jVK43vKzZpBdBrJBlbJRyUhIlGpA5/rEw/AbGOAiJR5K6LTIPKxaQyxkeul9KeERk8u0Zhz
7G80ISoepVCLeGRICzh2NTU+VpH/IjWKth4Ymbw0vLS/QKM5lnFnS3JnsuM5LOYX0TR5Hh7QPEB1
UPQuwzcvtjoKhEbe+/xoL/7kboRtPtZDwtwg32DXCwYQkbpHccMUINUDEumIFy26cCMWhnhXc6Yp
zCfr3xDiBSFDHeoqNVot0yApGLHc6fMraKS3voit32pZpG2Q0kQKdslU9s2agbkGo/tIxtduSoAm
c/yyl4UzKODSNKXWzLtWzU1hKG61uaCafom1gOyes2qiAG/76kH2WjU42gwoOHSqvj6blq3fGOhH
PGqZL3aOlu3RGTCOnQmOJa+CoLGN6Mt7eznUN5sH07fyrHCmprE+SfhTo4pA1aGOABE1iYneIlc5
wiCF+3obZ82peGzusZgii8qY8BS6t5IaCH00V8NebeQ2Hdmoepf69HDx/EFpEUnEdRI8bf+ltJ3P
+mBvI8lvn6lRIEXH7nzvES2uOB6hDREzaSIMfQRm1ws5KvNaYERWQGXjCccFAZonYq0L12aCyPpu
8sVvfCYI1M3URQv7EK6gzFgt4d6yjKkpFenQ3/6IZEeR73ooqZruHIYSTPO61U8XAbLfBnvUEe2p
VqUht1LWqaJ6Ld3iC6QkmsB+ObpmF4w3DS5GfwDLQ/+CXuFWm0ZaSHHTUWbRxqV33UT3ZPiP5oqe
X9px/DoePNt5SaRABr7N4MxR0FL3mRhQ+/WvKbjqDr1HWgz7FGhUzVK6SFjPV1sEvVB7+RN8VQSH
B0TRcZ6T6P3b3ePcHv+Sj5Jh2wDqTE5N4S8B2YF42NiU45PDg83tFNcuX7jGQA2RSUnZFefq367d
ouhv6tbBaPe7r9vjPAprzsJH34GjqVr7xn5L+aWfQ5UiIGLY+aUpc4ZMHlPobNyR2rX/ok56GKar
1Pk0uuovlTCsHpFMRk7h1ehxA90d1dzzU/+34yimS4ujsv9MK1Jn3BQK1GLLbUitlXEoXoxO/sLO
jjN1bwvMvA5igvOtbx7F+oAYGGHOidWgKTPGu+ILMxVg6z8t5jWjrEICGVwa+u5D2ZnECXlO9MRn
TvZctqugvzeyio9BZ1sn4FE4ih4myTAqC0qw/2UXCZDKGumGRhfBkJTnK6P5jOsp0GXnDpDSTwmE
baKN7EwNog7YrHMXBbpcBd5gUi+QTaEcvSCogxv+rO7jH3/mVW7cgatp+nrbZ2agT0KgC5aGfpM4
LHm1GvQrnczZBE82ekIMi1uAGoA2BKVwIazAp6CaSVqXzCghkZ4JWe5Wf82KcVM03MAH54uz4u2u
7FQj2zPJpTkwNa6HSKiL2PgXaExRImhqL/xW1gBOy3aj5nlpbfLBuupKqOcx8lUr8f5yFUFWX7iQ
GAgAtCirPhey8O1EIjtW3DUbOnSxEzPSa/2ylvdmd1G9mev+dVkoyOeKxZCnFFryKtYoGmLViGpe
ffAz63HpLYKym6eRiewknXFUxvvhrSoY8izymSLO4zXYmykg0s+0gdxdcp8jA+o1rYuGZOLp3JPp
0bIy7awYj7G2xnsy7qWXWFIsR8VYm0uLT2ZJEvxRHe/5h9EEKU5H2ejUSSspgOmbjMzsy5fGklFD
erMs2FU5LaqUZ5VuVbDHom+QvQDFHaiRUTBS/j4ahx+cALAOk8pMf+vYHhTBx+aZCvcdI8Ec1/Km
dyttr5SFL6NL26SG6x8Qe36Nevn+HIsn5wUQhz8XU+7uAuukwVC3t+Pmlrr+p63kcl3A55IP4NPB
0anh0/uNRzmL7skwp0/J+pewrsYtfCBxY67YRiiOXbJyadb695h3nIBUbYWe8hOlQzIM4/Naceur
9n55wLdtvA61UB7rC891vcLxJ4dAQVTYwd66gljFjRTmK1+f97Ko24PISG/Q9xlkZq21wh3WnXmx
I23aTpGQk6Sv53I2fFiR6OLC7imtZ8qRrl9/VZRIrXSpLXu5lhyVEhmTnMF4iP7Vr+eA5GkqApp0
6FK/UEW0YcuXZxDfHlkyz+7Iw1XZLEShgm1sTJFWsGHkhgIlE0MA2p9xL8YZg6TP42iytXITdjdc
rDA16fc+RodfQ7fE9SLdKWiGF7jJzWnsj8EySJ2XBk0AD40jAC2kPKX9mnOZBAHY8/JKCFcM+LOY
oteEmONtetl/UN8GUBsUCa0wS2GmE1zs+RZHsD4Jj6JdZmQRLBcGXS7i0tcWyKmN2tTB/16V4FMn
ebhtLBMk8jhVGKR6qut+l8VGTqbVxM/LKLPG71Ah4qwhnm/TyEMIBmFG8qGgL1+1gxYyJNnZ5J36
CEZwCQGxh31lYgefyH8WM7EwCcmRvOXFWnIaGPjD7XpDBSWQM9umTKbXDUjHmEJ5LOjATXb+LS0U
SDT03k0xqxuORfn1rHiMfhYIHP5bSrj9hPz93zk0HBnyOUEPFODmFm95ALEzXMkONeubsFATHw6f
Q+7s8zstK3Q19SXBrGpcOxCAwbMhle1jwJklVCVQ93UIGTZpk4a7imjapmQXgqEB27E8GdLC2THp
vqTkctLmggyTvnVGu+hax1OSe/8HHhLe4uVS4UnhpcByugE39VjKP+gVHOxoiD4of23YzTPuXuLi
jqXObHlGMoAr/A+lzBe3ttl/nguIlxzin6Rre6bY0PGjxMKLtk6+OAo/VcFYtAsNgTin4KixTVOw
rcRw8o93PTZM2HgO5gjU0TIDiuACNrgjcnUlC29KfLBLoSg/EIbqTquBxD2HLfGq1mALpiIJsh0U
piRlDcZl71mR9JwYPsVW6KVldrIqSpxJC8QoV7U7TjiUWKVwNe1tPIbQuzAmm/ns4ndLefaAvEYX
jBqp8gNk3kSaXoIpOGss2Pol1FCYB2MfjZ1TFhGJJRkVSdvT5g2dAayL6/yPIH2Rlcns7W+q6VwC
CwREjpFRCZSKtome0YbGkIfESghzRpoWCFcPE/TvgOi6CZw7qCZZWSXtzzZIJi7HZaykloGKGkiE
/nOn8LtHrJ629UdgEsPbZy8g9LDMt/D+aUj2uRaGT1/36GlyF2Qf5Nw8/dYiXvu4TrshCOU7pPd0
GPzVBHCr9VVnwe5OCVHxehR1yDUwQOI+uyevjAk87xutGLu0TCqg8mF1yErjGLvvadKjVGno7ay4
GmhfutKrhNYnnvfd/8fX8s5qlG9v8qlDVaJMbpmcrNlbvb9702LVgRod8GlZ4YDYCdj2ZBoEFOc7
g/hIrxYDuZr4AGCzHFN3fR4FFNKfx0ywSxI/Lg+vu5ktAU6EjKTILtTJDqqTgbMuKtGZHxWMN9yQ
yRzVwZwH1PfGSFHiPEq4tyL2sVzMnr5LSTmPsJGKsGVqRhgAQqTdTh6mcNj25dOfEX9RqT1jfCid
sgYxwmgfZQmwtMBAma6Nau2FGslXUNWOyQNcdVLUnzPK9GP2kCt9B2Qe0DJConWDwU2J/HJhWIAC
YbVXQdhTngONqPmmW/cXWTaeL2AryRLyq4vspCd3Yfb5dU6ojYlgJEfi3nYUvlifPsIXD2C9J6rv
/WRrxNjwQ5NbFCSBfdR18kp5nNfevmAipDROZwfM/ywwqUnTAv48WvNsEQoyrPhIOAHcEv2P83Q3
c6NPiY3+Q8URTP/UptxjrtHnCDNgfkqJixr8sHpI5Y/x6LTtBQ2iDP1frb4OGegMwak9s+9iggO4
iuwuoBYzlv/mFNbJ0Z/Ft+dIZ3OJMbwZA/VrpyThf2H/lu4E5MoYqRSzuiUt/LF2M1cwqXQI1jIV
aTdY1vpuFCUCKqc4EQo6rL66bpojt4vTcGUE+vP+7/8n1BFlqFzy2WyauDDqcXJ7CEs+o5Xwj+gw
MIz2nFFFhaz5cnInJLvEN2b1Xn5KDb5U6giuv4Wnb0JxqiW4n4kNzmGcrx9Mc6elMQmscXxtEH7A
vn3FN79CBvaAZQRLyEXbMfyyHIHvqZXPKEwy2DE5QIOH97NmLjNlSXyOHZh32Czj+NODIAjIfCCm
4NByzi8c1BT31fxqgpc7DtSHK8vBMB+ljyH5uocgAQ0jLHAxpkkDlZcWDEqetIpWrk19/t2W+rp7
650aBGyyWfd8eeUoUIaNm038L4vv7PukpkpwHIRvRxf5shxaLC6448Id2xp+KK25bGmrlPMLgc9g
d2+jutuj1jEDTd7eqw/ATu9wY4oHEe1IgU/67Mdr6oUhlD8avOIBYRwpDmxuec2TfRQqOug8LlAU
f0qE0JJb9BCMPVe1C+GkNZcX2xoG/kVED+OjPtn2Mqlf4FpiRfM7mIs3SZNj/DlHssohMogsTZhh
zHRprYwAmPK6r8qWkS002ZMMkqmsUCBMFuNuQbYx4Qo8gZdqoF4uHAFVuy7CjQ4LW2vMSAGfAeBA
H0TrEI+nA1NxeId9gqEFVOYU5ZuJGm6/rKzjA3pFOpfzpOC27c6BINhxF40H2AecLp0yhAvsm3Sj
WYYWo31qA9XFBWzcMZEoqrGZ6cbK3WvuYsSr9ICVKZY1kCSTqfekRvVDuDmAIV6ZXvcoWYjORYGV
PI4icVUNnSZ3mSLszYZ0ibYRNC4iFqaV83nEo5VSsaApg6bJhMShlRDzp8/3FevodsEj1We37Fhy
jHrjFD9bFUOAVJKX8i1OckCYhUkcqsTYvG3VyHYqpzY7kF7ryHqP7b1CVrXAohsu8tQAv44OQxwA
vbX57X1MkTz1hDWVUZc2l5vmtMBiOIeIh3oGO63LFWCh1DRiGQKv6Akybzlc5rGCsJ7YSh1v4B48
PBtLVXfPvOWOTDjNO7unYTnJDWIHeAKaSYvIVYOV87i4Glh6UMlXOtD/gcL0W8mrYFHNabkhsTXu
ZrWPj+OxHBUvftQRxe2Jqc9v9MwEDYXgFRi7/7G8txZqP4KJQCrBwEnYrjTc6tfMXSswvVucnHav
47dV+M7mVlM7eJqUXDonL5PnuxBYv7DHEnTBfnA28tRRFcUQLAcXNry57l71zezpUgwT4kRrY1MN
wrkxgg1X5bbrsfIJhF9Hc63DD4GNckcEiQI0bBZg1ZwvV6RBktHdH4D7+q65AVm1yhFUf7N+gxHz
BoYo9Vlcgufvvhkn9+WCBNizfCaVWmcJ/RACyg4a10V71SxNsy2kuWp/5oqVHPi0zn1dqNLrC0uA
ZNbat03tK8XQlX4dshCcBoh5jjzxC4IJSfZY5ANXr6g2TDn1RHJApBIS1116vTmLyHlkEUPa60+a
tfAGM4bUP1gkNcZDXGSi1q0U9qeF5JF76m3gS81OT4F2LzadU3wugusgcqKGgcBXXzvF4uRIGT6d
33jHnV4+PIslVot7oFnpuLKzRX8bYogUS2v3ZiHBpaMCpYc5Afx2uqIs9dcr5pY6tJ4QGq0h3LlJ
0V/N23orVv9ztUOHA2hjtSL+XHHuKf2/Qo9WRipMY2SRNx3O+rV5UyHz6mC0TGpz28yNoZ3aKmB3
czMeq+RFZM8FSzWKmdz/JGO6M5wFnivvBZqBvmes17qUphgRYcHJkcGn/YurvI3RnDRqtif78wJB
Xh411Odu5rxMBtzgKWzmaipNJ1Q4ZqFnghVeKl3GeNbSfxyqegohc3EsEBRVRCO2WeHBKxgFYvYm
ZBxQBvJyaqtKb7QmmVwJfKmVZbaA00HVVXU0/80QYNOdfFMIZA+1TKNnTlljy9/JxE3Lxp0Tyhac
Tw90329VbAQpd0cxTn3VWKgylf0j9u5dUP5jLCGrwPDSzj/MKswoE6+3DulOwLhKgj+VfKdM63JY
ggN6/+QFHglzl7Cb1Z4hikNb1J/7VPgPp6RJ7xr6UdEI2Rsfa9+36FJ9qZXiIVdT+r7f+DegxzkT
tsrVousuMWE+gwR1ODWM/wfgqKncqptDt8kO1UtSkzw1rkSJ+Ouj/LO+wDmRZcNua2VU1noH7QEP
0rft7yoR13cwpfi7PvdzEFrbY2oJWobOrMZ2mIIj8Er2wCIiniVCpjzoV3fCVYpxpQxate3slMC+
oZEYVPXITwk9JEc4reKdcgv04yx3eFNyM0SjWXJTU9LK0gD4eGjChmdI010fGwvL7N3KKmh/Ipxj
ZeyZfaVAnWP65r1I8Df6QzOUjSWCXgC+FTEYnrFKFj6t8qSbxGY/6dTvfwJy/hnQoNCxxRNmlXR0
wJ4vj/bv7eQ8KlY315nI759VozEPYAD5RFwVp6Tfz570I3CsxkAJW9DzmzGGSwizQkr72JSYAm5M
2KK8UjJraTLVnqSFD0TQM5k9dsvl6ExbPvKsozEkCdIAH5q7grJ++/Jzb8YpJaUCD/AImiupCxx6
Ky8VsjdDWGI1r2Ejpi4iBrp97fV+XRmlJ2pynTMvKEvJMnz6euYPSkwhOYj8/QOezPDX3p/YPfhB
JMvspOR9n01qrvnm1c72lGHdAE96RbqU6PyVtkRrj/tB8F+LLmRfqgy2sZMo0vdaOdrLs+VF3eWx
ZPZKbW63J+pZny4Qar8kUMo7ANh73y1xLSFF8va+kb+aq5rfHf82lD01kTKj0IbfYVDEtcSFmDGT
fKAR1DMlz67ItC4TKueEYYO2eIOB1inSrKelKBSYZr4nlswPqmGNqb0JIV9VE/1raZD8jow4IZO/
6ie+avnTGsYu7o/EUqNEbxu02QVD38LCmPjdMGs68bYnbdnPDA8Ir5uHs3YZxPESqE1q+7KV4T9B
iB7/YcEhAur5vSVEXSorO+46Ia4eoGk6QaXltLpof14Lyj7FTS0KSOPOEs3pLWeRhYHWTd3RU/p7
IXuqTUZtNm1o2n0ov74Hpt1x11lAq0g0g2Fo2nGDJVPOe5rdCkIW0Vwl2zhfl+nOINkdp3BIXpCI
YnzWGe8IUDmNFbDEXdA8gU+04RW241AMHyxZmcWFtZJ+T340URHfHiktkyWybRUC1LcfHeAgXohI
F1T+bszHuzvdidvlMvdoyB9YPNyGo1NKVCMI/rQpL/kpg4BaV/AnGe2VWON7ud3XCetekfXhdfop
7P2sKMMnnQw7wk2ogP6f3iO+T3E5OvgoLbg8Gh7SxeB8v3xZHbmSGkgyB/T2Hu1HbqEDisQII/78
eG9OX4h3mQJ0gMzzR3lD1M2kPlR/0olosKLn7WbG+zJP/tNEjM9DTDceOK4V1ePNWrpAQe0LsLm/
JfLEEgs/V65UaPV1HW60x0EOYf96aXeQLKS9qCDOcJjtq+hv426L8d62fOCHXk3uad1JJpUg17Ec
dfEwOHUVGedx2CSqFYMS3cQTTIt0SKwfQe6r+vMiFFliX80c13c2tpGPhNDh5izeniWdayK9a+cU
8tPJoZ7hNVb73Xm67mF7XlLFyND5vapaPDrsyGsBwVRoNDXVP1ln/13mj5FLyaeJIyC73kJhD7K0
OavJgpy5R5ZGNLQF3+jU/zLAfkh052DBgSLNNm5wU/b/uxisgBiDdwbRUvfkS1yfPQR3SQm4de7i
wt82np262WxmmTXfa+b4uCUAyhvcaxPGdRzRDQT6W9oStC5DvhR2y2xILSg8YM9oRYGc2sAscw/n
I3aaz1zsI7+l7Uv+wFZ0wPWYQzELeHEEXNW0XjuVbjYVIn2JXoUeN2YJGKZK5UxnD+plqJ0jkx56
8FprhW66LUQgAvYlFjF4La19Oy/oGL1bkblv1bGA5FHSqt8N8MZPouvG1Q4t9wZZamKC1G8ux3Me
aYrqnfnjO3g3txMDWP2vP8pxEZ3l5yzbNyN1Mea5zXUp2el8pXNF5Vczz29JZp7lg0b1n5E7FKfC
GRIh/BkE1DXQAS9+Rj8VU0AGgI+QVjlLr4PbTIKMpnm6cB3kFpSshsNorqd+w2aP/lP4R/vjqavz
tROWYVLeoRPsyp96jFYrnYYzjnMbQd28C90mP5mW3HyPZ+aMBotg5QBN6Yu8FanlNL6uMqfoDgSj
MQjSAPqMl+6DHEPF2TKmSPLoBQgU+1OFjUjbHZrpHUp2Dc+9Ni7/+V8f5fv4+EwMJ9es9LF9Jef2
0DIILk0iYYS9bvx4ip5EGV9FHEJSkoNlaS8gPRaxrgH2LG6nnwZ1npoBXWxazdLdrtr3i6qkzx2j
UQ3ap9V75wh6vanc3z5lvzs3UiEP97J1AQ2SGqHA2dwaq34+4CU/OP3GzoE51XBJwFot9dvoLJ5a
kawep458ei5s8nUmlx+rrppYuqGPhqngcVg7mb3CwzY+ZS6Sxr4jqDE0K9PYl9OePSuxp3WorHos
jY4MAX6HQj5yPiy7MT2HbGJUqHPpByk+BsMWFT2WjjB0LIncnJrsyiGIjN0exjYSfZZWNbymiPol
4+2tt29n83IuPCqN0gku7RteFb8pM2b9vrMzD2w5j4u2GeTKM17tbjawXlwkE0/ObEWFfGiJ32EY
Cp3YMUMmyPcVoLoLHd/R1C3KKCQCmRfK3z5n6Rq/+1WilXl2MNf80IupOFzCb7mIflqaX6VEmEur
CrBHpFNw7V34EidNouPePeT/tXYIKQuR4NjcQXhSrx63sSh/eF6kvEs4uf4obZ+ybD2KTtE1+T/L
ANjnvOI6R5fZWMcHXQzMl7OTa67+0yZJyCvqpQP52LgjVgAGHzLWCsjoTB2gaOp/we5z5vI95cu0
AFB0wEVnTFW+g7eJ8SsSMhG3IDRU6k94V0LEPsU9FOcHooi+A3BtY0Vx8WIbUOQulCsJg7qOE0B3
YU1HnxOPWu4nFmytI38sLRN2JjY/rGJn42qDfE8Gc0ME0FQE7iLRqZJwAROzkDpXM0U57JMIbefZ
Yv2jFya3pT9re0p+p37bqbACQ5z3/UAx014kY+nozor3jjeygGBIRMy2OwP+wcu0hpQon6Wk9mlW
JIl/M29jDI65uCGJlHXwbFdtb9r56RT8/mkQF7+6xiivjGUoq2oYr+eovgWxDXYkDkGtPyK8ezUN
t3y1aBtiOsHvCtGTnB4BtSOcpS+rLR8bgnh+rB7lW1VEQF1u5tDrPhIksnBJ/bi8LRII2lE8unoV
3CfvMLrma99d9NrFG4MPE0GtVfeD62Eb6xuzIeJcajc2BB340V50varJuAt8wt1JVW48K1jzYwlO
Xx599Mt48DwzISySTYsi2EvU0EPRemBn2HV+D3qziZZye+qvHjhY6mCoGjoRqNLolCFpsJpHzEAW
Sm1RT4eDh+lJuxWGbyMJktHALEj9dZmhMu/QBhvgg0cICAlbigYLV1AfqZWTKY71L/BFFjAD9D+M
52BlRHG6btBXLsgrAHWR5fG+7NSaR2jAYBMdw4DXkNA31sx6RfTRxoajWxqiq4f4FKyvjC7n2upr
8hmBEPvkR7WDZRcO4SW+YZIePRwtJG6Swp7kv4I//4mWqzB9j3cmOQLBAUp450BfqfQENEtUu+vA
S155AB/PRkZpgxrb8ozKd3n43Y6Bc1vrkTA20+KAdgs5PZC6ZPjeHdtM6vpmmgFC4GwW0BHGia7E
Wi2mQ0jXzZ8JvBwNMpRHTHVhrlx59AB+uWMooSzCZg1B2NAQQtlAL39vnyt8hUoBCSzfmmHsM6rb
qVl4OvIBVUw5w1/0K6e39Jo6HDqh2WaonpQHQqBB+wxnTp7vsjdTtGBW7FloBSlJ6oZC1iBgQ8XR
d1f8dAC8gpO4Ut/ah2wARtVp9cYuv8OIKEt2MNEqF8pGHr6PwzuTP1cTmLSplOA9oxIkfWSKggX0
BuB1w/o+X86mfd/BOFCHihKTQS5w7/qOXf9sW/PUBjLtc2sddJ7FFv/38J/e1DxkjTHYeSRS8Sqq
VECwmOTiCz9ERAUL4doTWPE5ebUSZXlPfzyjeuskR4afCsuzu1RWlRnkVFBz6nmcJi9ksW6HgF/B
mnmEw54ms0owBRgp0rwEM2lyboeoeHb2qqci5jPfkAHgM4uIcIJbNHEmLouh+B+g8OGBQVdzHbei
I9PbjK3fOGbxiJFEowqxg5JIGG93UbStqKdOjBZ6Dh+CBzzK0AV8Jnzzyl54kHgiyvN4Yw7BiWYR
oQ7Ia5MFjFtkjQqNf0eWRN0X2lPqb2ljOa3jMcOYPfbrOKLMLypmVdrrr3vYp1fGvYg88yI+pH0P
lQnCzF/5H8sNuzwUS1ZZIhiGIsja/Zor+lbISXhsfwgHjLMpFN0VgBvuX6NLrFOlAgv9JmMD1y1i
1VncY75K1P5/d1alBLy1xAEUpgb88SRubJ79SJ7oS2Rb5uBUuaOuK6qFDPtcjO8/LtmwYf9l05p9
mf/OV0fYA6Axw9e5xPMqs1N3fWf5LDcD7kXIrrsI5snUJPgXf8FQgYxndxyqSbuhu15DkCpNmZ1r
hvrtFaKVlOD91RzcU5Ji2VK+gjeWMJSSVUegM/CMAoed5z4ppzRGobg5A3sLF5fkUZs8D1xbxRzL
QvKixDlUJzQkAXNVjaVjJSVOC25uLJh4rYL4xwiQlVWPulSDVZLASP22VkKAH0B3Obm+MPEDC28h
kWDFFoOaympfG/9xSnqxYlxGp4rpCB2pMDGqj94BJEKlQVF9rXER3EoHf/LTC0N4HiPGNRmxm3CF
UHiNx4ESF22bZ/Np1rly0d/CybMTynPTAXczR4cEaQ7xe1lNesjnJTKR3HlJGCBAMIFMEQd5HheW
RllL62s1JAoJNkpXHlPQ5y0GLSy/fpWVYeR6ZLWA5TMXCsg5DceolZqB3YCB4NpruNp0FrWVq59t
kszPX16i5AMkJI9Yc++DmCiIlLIaZbMwrc5UvArY3LXXRzH4pOC9zdUVNeKfWRkzPoN2lVRi/HX0
2VS89cGkzNb2apdzFaslT+O5AzsnMnXR5Zxo+gf0m+5WOkVC0HNbFHexAhet/5mzWL1ndb46n5/Z
Ber0MBu9SS+0XiH6uRHoJPD0fG7x3c+OEyQYnrFk+ZyMtu3KBkC8pbG94BHYuuRSyQm4WZODBm33
oecBx3fURgNaK186u96JMenlAIQ06sOEed0MpFKwEw5u5WFfj1PUFvkyx2wXPqDUu50xgXjRx3xb
2tG7tMw1+8J5oUXYFk+bnbrdPFiuxELLIm35sMkf7XrSvSwBBwR+LEj3p3gN3kjtlJobf/Q4XZDL
X7+YskzD0e+8BVe9BQU+emKk9oN7Zw+No2tVEEjx6Hi8jR1Ilni0SLxiwZbMG7WtBBpvC0mWNxIu
8BDIpSQ1VwX2FDwQ/agoKMsQYn6vWRepMVJnr9dIE8WIYGzT5Ew0M5LHW5M3oMrxDpj0iaRqc+Po
mHtnDwcIm8qx+5/KQCSt+kFeVCXHdHaTwqDUF+CzNkCcfaQyIDvs9NJpJxkXCxzTObv/LGMwXzC1
D0SGuJFubd62Fppj4JDR1qwGwlNq3l9R+sDfSTWzLeR7cs9cP/DgkxWd57/cxOCF4BKAaL7d4/KC
fjeclGeSWP/EgGG94j5k/0cKw7vevWrKpCSiXYzJ1OmMm3OboJWzTrUq21YKGFCVkAt4by9AxBZ8
gkuIpHj2b7n0j6G8FviaLEDy0brvCQWK50HeC0QlRhOKBN/Hilb2TGhGz8YFvUqHdcUHblyb9wh2
3eFt1pjXGlsFF/esK529O80raN+t3FdhiuLJWRwdH/6jUMWXaHBecRL472A6WBcAp8MnbaM01zlC
giHvn+XKZ+4QeV26hchnTltm2aGtfYc9CUhzwiLbojCfZJNx32Cc3fofWmmWECg5HWQoBQJ9XQs7
y+xgTduZZ0L6RRm2f849emLOglII/shRWDTEEAAsZoNLHYGaSrT4X3snqdwT3F46qzf3PKrMa8Rq
61fNedxs73ug6naSu7Xiw++blBZReLaawkDJISkpMvpv5+gM4K0LhYqJWOZcoWSfXMWHPG3KxsP8
3cvP7al+x48de0iUrZ9UYzAsPNPmSXOYJmFTMdPLGvLsOfPJrRrG7b0wEZdjDirsfxunEalMkEBD
JM6+bI1wkE7xMnnEYFeV+TwJs7qHE0KIMA6x9AOekdZKSsgz8trl6oLaEomA1fEzfNt5DXbi3v/e
Ozwg++rIXxqVsnRrtvn2MwNHpq/MqNQ/1FcyTOOOvgIz6Sw2ztQSI96o/DXy0G8rHMq/WVcSuDhL
5yRTzBz3O2u7oDwUeyh9HNVniaNv5EDpmQiCaNLMZVH1VW5ctDyfZifcyPcvQMt2Nmumcp1nuPd2
9NizTHVwzeH8BetY7N0hG31Pko/lGyj99xZk3V1DXWoJeT4l37UOqKoDj4NUZaGEkcqBek2HN7Y8
/JV4P/ohuM8WU9dq6PhvfY+04/dZGPQpTdrEYn3ggjiJ4bI6wOuU8iJraQYUoeDWOe/rw2/Noqgp
MBcSwO8kOe54CRrX4C77HOSj0uYnqRbY46QadHyY2MEG2KO+MFms2iRzGkotrng4O+Ywv58OyV5p
gYMPno294pC1BXM53EghEqwFTMYep2avkNSg3ZMpQmNsrAye7QeX++uOZBQ7FBQMC964iFuDJ8P2
A1CykkvOMPHz+6WFI7ranIECBmuE6H7Cm9HOfr/DBLQjBsMqctNEYpHk8ktB4BIUlWdbK+6l1CHW
ww2+UAECUrG3enIoqeeB+b5BBSoGMhkuB8jieOvsJK8nHZeQ65XlHmahmxbCObVAvJApcrEhQxeD
w9zzJcCx+BPDTMBd280ys6Hy1T1eQvk9pDm8INyVnowiIPEGaNTCcRFzfkBXH1Y7v0zJ7ir5snhb
SbJqOz9ltok46XsSkkuTWfpGJeCN5eoJWQJNnSBYdjhqfSoktkD1kyvzqUh9UZg/E9bqoqSDBRt6
CrKgpOqJ/df6YsCIoCBtADh5ifiofMXMh3VYZV8HEVezeZPiQZwHvfshrN2Iv+LMOWIhn0MWvGGW
PAfxvBtEeiatyypcXmYb76wNNZIP3NPz3gAuwOBNGpEewlN5AMCBzOxv8gtMdSoxcnb+11In+p60
P6KcKEs2+gKzXWEOcu3JQ9km11hVg4Y/rpuwh0CNkA8cTSG2i7rFPKLOqAisgpRNuRwf+nOJ6cHO
7945FWRzTEXmN6x/PUqsyTPATn58NCpuHB75byepjwITR4ks+lvgGXLrWDwsOB1IQg3XPAMJksml
BJwZA9ghi/VXKywsMDfhAA14xFrs53e8yGDX0HzbgX0bFYDgcZBbWZVBp+cTqCorciwtb9jLpv2T
woQi7qi+Rr3CA8yGEef9P3ONKsEbuhxZ8l0qjBOimvfGoBN/MHaitxzoAVD5bAFcp4KG7ljdCMUo
38pwNxPLMOSO5Ds1dtEKUmx4luShvTMgoH9zO//MisSPOLyeU2OcxSO403ezXQd0kj6yOosQzyvr
+Gh8Heksx3k4ED2K6AV4LBb4239JpAgLZ/1f7v5RMLQ0G2FQBqcXx5482nQi7XX00Z1eI3a7gKUm
p1fKS5/xWIpwleOwUpjI+Z9P65J2SdsRAy5m94eueKerwVpf4sLOAj+AX0qCYGv9vxPCqX6A7Ptp
C3qAh8W5tmRvOg6WNybyueRqp+cWz4CiLxVSo5rfgEzqhTI7gftpLG/G2M4RlKp923pRUGQN+FPe
M6rJneOfHFWHfrHHDn5YvrBjy55HvVuBLFiufo8MZSUx4HRnwxSaiNLYimKZruAQ/ykKnNPF+xMi
e9TXDZzJH0qciu0yA8s+S5GMYQlOFuXFx4AD6ppVmX6yyXMxCZfLUdQZa1SFMPiExS0/wsJGLKX6
VjQwAZIt8ZqorNxnfYweQbVPd6noIc9o3DErELUD9cUzQpXDqQqlzKE4bpS6MSycj6ZT2/0d1WES
mT7OAfHJPLuoeqPFmFumEjp4sDhp7E2SIxvbgB50FAZNo0cxC1pajWClXDxgoWnyIem1D2UlaU8t
k91jKIZ3884iE6Ga9HxtM2CBUBxa9T0tIwwcfibd0OwSEK6HRmFp1YDUoZMpkfpHZNQeVAgRRGNX
vja7of0C3SBrieMhyUbZfns1FS8ubdBrAx3+Kz+AR2rCpm6Kmz0rVTyphLZCnVntTzqgY0INn9Ug
q5hBpHLSMk9xjgGKU+1K9y/EgX/UJEoNzg2Npq1U4p6SYr0eWRRrZTqVgmAUQC66b5CTepKEnYJK
SseZPy51vcK83eXRoI6CHbrrP4m79fK13JQS982Uqc2GbihEfvOouEWOzoidtPcaK9D/lbIOK1ru
ItorrmgAgyWY6bQlgOK2qd6g1Zn1WDWHN/09mQlFLdCevayL1eOgsT8jzBUZ/fUqld+VQcKsidmX
UWO0n6cDzdCmrG1JpMCIILDijMWH4oLzCQUeocpJylV0BEVUqs4sU39QLQpVqpQeAspLb/gVyksy
Gy5JUjKPF/PfXkUv1ju+gEfeOOatvXdTvMQT0tv5nB50VbVd6s1vf+h+Uhz3PFQXo3LGp1KPuhNK
NCh7D5ehCR64W81QOcavSSXsosQ5vBRBAqIp5p9LVPzxFzwsjXFjjG9mqOAUP3nh1bpV85F0hsHg
E7K6Mz7aj/O2lsyVlKV7hRasN6fVAu9wRNVCTYRjd6jnsAM277aykZ0NncWFqZRzaXDrtk3IrUof
vNvTTH7aDF085GuWPIAbx2q0eQWP0PEsnp+gk+6qW/zIEKeDXGiAvnpRth+/B/zAiI5Xea8j6ZO7
SN+jODYtMVFgrCT2901/tvxd2847cFqhYbgcfhRhf79Jw9SRh9STR9aIldDSSWY5SQW7Obpe6kgm
pnasZWqISt7rHtQWhmflQluajbFopZgWxzjKDg3Eeb69R31mFfvikemMACYcbcfA1dEGi5v9QjqT
ZWAw6oahcknTuUknNS6/yb/H9ojc5MYYNRttoa21bn3a8UVDW0EmwNDOPzWRH76wRceEIMgcuzdX
m0qVsRXp6+nVRcAWlVPU5St0Dj8Uvacf1AdK54/VwH7yEMy+o5GJBz61QDORgo6mouG2kzgAXHZa
d2qCQHPRulrIzAQecguobnkC24EQd1tWQHF13NzrKlgU/6ASIvYrYzW+f+Z8GCsAJxEHv7NGo3iY
E3enXONso7/cvFzKuWRQPZ2C2LCQx/xC6CxoO4FHfPo3TZak40lBL2tH4SRc173DQZaH5M4e06P+
Ubhlld+DLQ/RYDb4EjfW0peVXkF9300YSkADhrBVmgEG8JujP0uzqYGjKvwyymI+wlM5+3KRzn7X
b23uxKZ8CnGAgU46P0FkkhpkVYrT7Z/vhnfuM+RxoW5PDujcYqR+IIxkdUWl0LTg6l9T+Mx6cKN+
/OGq/MaQMRes0LezOtB7wH1UEGLd0k8EIt4XwTVowm3F/s7CCKh/cGxHqzjIIRxX9mpJAkzB1+YL
OH7s4oiRPuq6Se1sMHIjjxAMqTtoHWl+kYq9/bYMEALaTaG8WhxpYRqVRyCxe543O/1lTeclTjZ5
sDr2gj0WZzJTzjwCNmARVpC76ON4EuQQnulgbi8m/906DQXRU6Oi7zhZcC7bttv2xQMEBSq0rMGq
p9aC8Ib3W35E/x6w9kQ36yQCfTLdfKE9aFXyt+VJvZM9OrGnNl46dmbOxCiVbnUk6IEoMUmxUpjS
z3jjM25iyLmrd/GRkXiatuAMYNDC3GMUVq++7WUPgZyJRoX28r2RRGTgqjC9fIIVQAKsSaW1O06p
juiZYOBrAZSPp+GQxrGfwMMLu/fXSi6QgLl7ed4zJP6fglZndeu03qwRr/YB+hEWlYTl+W9nLsIu
CwVBxEvOMdhNpwhjGEwP6PjO90Fs/yzN3enc9g3O3nUaM7kqeK4VM0Fu0y4HKMt4o19FNvxJ4LPS
hzVZk+fUBfaYQTQkqvMqdPyDJkv1TBs7U9YZgxcaqtSTy7cvYhNHGx0F3j41NgXQQ6kUtz0V8gAq
fS+kYxmmOgVtBV/x2Vmz7xJD2N6j/oPuVQc7yY0uKJx7gctDqhapmp8mQ0WPDz9mX3VNkK9xpXsf
IAPq2JePCFVVQw5i1Eb9nJc7RnYIgDl3hWReKcMdB8IMYgxoHQsg9EwMaKK5obAl33Loy30ru3XJ
iaqzOacjpbAUu9jXwK+cUbYbyllANRUuzlREPqR0mL5WRqBYhbKu5I9CFjNSHUFAe/MkKOyLrTy0
wOU+MBTAYcHDFouxqIW4P5jtcPvv+NAa7vpEk++Hy0zl2ILKR7M7sysF8hG+xaba6Qrfu1W+XJn9
9ioY5P3bdDnOECPjQZ+IFqh1rCKRRf9/fCGwHjg2j1AE1kKupWQybBq0A+t7TV4jlaEyxmjrv21Y
ocfQs18bySopHE9onRpEMqZQiYECP7PMxZa+23ys5eam8iDTqCi5Yij6AJHdds/rANhk1E2Jie7E
M607BsJzV5m8kXg/tG6VZFPLmQWJAS8Cld8WU8IWZ6gj3FTQMwpeKhv956XEdwVYs6OjMJTsXDou
/YXYf9MYFWKMKHavXKyUBKYYWY9FkeIiT2MerCVgIGx+EtDf34hMlhaSmPSvTue4KYzhA6e1mSV/
9LrXmf0KSL4Vy1/XQ1uI+ET2Ho3U5xga3ECmW1rOLSKSVqbj03VdCKkURUSQeMnEtXiLOf8j6yH2
l4xY9E13TD5rl8MJBWI0e41TN64asFTqpGgbVLLJKnsHgyOZJaBglsKAAU08U0YMGpoeQvOLPCwm
KjjAVT/TSQEMdDT0TH4PE8b38GD1rGR32JwPfPPkA6JMPuO1nUvAAr+5ps9alR9D2OrhKK1UgpDT
/pxQn+hS7yLdP2vbp+K5bnI2wyqB0QId/gpW4C/X5Vol5YeeFsROq3bzmuCXd+5OJEJMLWCzd0TB
W8WMbG7cERbLpVY28bCz/E8SpGzps8XDtWi0U2YgAIHnrH29k8sHLJQR1kovnUSVq/oydGUEFbi8
hTOndJvSdEALFXjGHJAh7HtWwqEWqRA3KboDT4XbK5qxjkjeDE+dR0xSNkgIq6ldzStPah5k2tge
2h+6ozTXjK6EpeJ+INLtOozdOak5bn0Q7Syb4NQdYWoG9suvX8KeocD+xW6JMT2fEgCrl/Kc8Qm8
9ZZuCvukksjx6ZW+ijDH+v+/jc3sYmMoqOWMCbDryo/gG82ZTEr2kkwa2ui/YdDxZt30e/ugsZu9
LKXMT/UGvNEN0SqLLNmpu9YGxZ2FMQNAH/JgeSXWSdNjPjVt1BRvKWxX4hgpop5HccGg9363BoZ1
JUbqSEHj36Vkj+VirBOUOC2d29+gvS3REandi35PJfzY/j+y4XvLVrvEzLjpQRWmLUgCCfMgi7NU
UaOANUY3x66aLeaVxkbxvCfOf21YcEExGFBXho+5fE4pdw60QRm7X988H96kgn3IpUWCy9GbOVk8
r+qiWOUd5JdSWSTm8dqqFxqlONFQZyz4rsLShySnKzB/vMfmmanM3SGPIQoTkad9ihcx2OtQkHkn
uuwEKo0KXacRax+EvSFUy1mWbc0Rb7z34xzQyaJJ1g8LtrkDOZxHOsYVtkfxH3LNiuo3muwj6sCB
07FZfVePtvDrT/mXJXtOdneGcv5H2vQtQYAeCm4kq5QDlvp5tKT9g72cwBC00Lyy9KFXQYiKJdZM
MNPem6WayypURdMyrg6mTNlSjbahoY1q8+Bx1XkvK1RM1c/4AB5UOCm5/IUAnIm49mZSpw0FQJ+W
iKGPMRu2XUHvA88l34fe0CoFaiBCvCdMeFXMhyzvPI0LYzD0hesnlOgIJHiXFaXRmBKwxLH/EScW
jsm9wMM4KL6/470vfMowmYkU8EI1qqL/bAYrgwVJdzH+TAtVw6MOzUddaZbKOdineoPrYQY2TLCI
fqAxYvv7+wyhdawTrea/48f6QXGfEiugPDUW7ud1uDe8Z6jEYx2SEDIICFbp54902PNn1xItSZH3
BJvfDPKGcJnetDB6UmoLJkxbF1qrGd2MWAybMGCHL68p4VxfOVkNqsYY1jll13t7hFz1TXr89li9
wFbFl/e0n5Xr3e0SxpjJDwjDuQIeoQoxpKoYt2CFo5t2gTeMGIeDmum1dnFzbZRINQpiSgaU36uY
cswX0anHq9PCsmmwTWkvTW9G+grFnu10XdMqzTZbo4ePED6SqvpPcOWMUggmm/Nm/HsGd8Bw+Zh/
wbXuS2IbJBcmGtIVm+TYNNn4Axg3oHaIb3mGEh2UiyaCDfHL4jhJXmBGv33IZNnJLJOjydo5cuRK
T2LC8mymXY/UUj7zgL80y/V41/M7BxllufxJh60+ju6SRRZR2W9A+iqijEHi1nTGLzQD2XE+aqDq
upC8c8LqIWVcPmWvhAJFRml2hlJgmiBWWWbaCDwz6QxeNad1vOlWCImtCZHuU3GN1++FIl2xUwVs
nIEte1yMgU9iT/IgtzBTQEpzXM+bZlP1G2fip/4jtxrU44fd2GJRwV183lsVV5DvdzfqcOKws7mO
drFJGc2jm/SVB45d49JXHTPJXY7QTYtD9ksFk5BLlNyGCMq1sw/QFYwx2yJ/WGlCGypjLPp55OuL
AD342stYHfR+9iFaXkjOWsCIdorrR5Yd1DyLYKLcAyT8AkNmaH+Amy1cHFxd4XgHuk02nl6Cnc5e
z7IFRtuG6N16TvNcoVNSRIRvlGERsiKpTFNmsUJJR1vfSkBN8OCKNjiBRmvkXK3wTRnzRnXMPAiz
5oOvNHi9f3CTTx5Fg55GcrJGRlMwbMIKxGrx1iknZE3kzBvXpXPllFlvduOSASdFoJ1pWBGqawpx
oNOUCgwvv8sub5iy7vtircggBZUy5lYIthdMcQTAiAzBlr3uwFUQdaQpCTe59Jbq7Sx+cc1d7nxR
3nqxk6HjUlLWoN3esf4xgewjjHEXY+IjDzWu7RhsyfGF+4/pN4dH44j8Vux5Nrqou5OTI3EO8Wfo
XVUgRkfpqavTRbCP0VIpkwS3WNJJAhpUaTH+7090Lu1hfAtKWST1iqfSdBcigMr9B9D6jg56aYf9
NCeBp9SxAAgYUCfUp8+5ebpk8B85lqXr6gpqjwi7VYfHKQXVITra7Y+eeIKNBIwSXJADdJ4Zdmne
414kOMn3NwrxMC/kqwygbe5tFzjrRwaqrBgYQxLiUeWjRd0e3dkE53bqI55bvLYngEKoD0YXVDTF
3uwcpP+SoaY+zeRr3juOVs1A9qmbg6/nmexSfKtuwD9Y43oqiEJhVhNnOemJOhkeVrRNjJX31DpJ
HqzMse85N779YvjwkZIXOJvWVhJAwjp3pc18Vjvo9MCxGj08M6EIbNX0kb8Y8HmP+dSg6iVwFvUs
jORaxfMkdqosfTxtk2464S4Jk93ewUHtODkda0CS463nkAqchY4X3heOXp0mGfLyqZqGmTi1CBb4
r2g8qeYcbp6qTNlY6WhZg6x/J7j0fZVyUhodLHPjR+6aclopDDL/YiTmGirAeyt75sH94WLnPwSV
oin6k3AdOOb/uFjwLJUXbmriVHA/DJS/CCnHe+lHPSWIXQNWgFlIODtU0eeWKo7GQyjFTa+e1GN4
aanTC3HhdzmfBcQcw6xFr0Txug0iBa8QhMspIf14FfR461ipGaPDDeH3YLRO1xeyvQEdxffBnaE/
dRgpeH4C43NWXf+qcouLeFgBmZPZOFY0ekspKGxaW2qZWKZCLxLdIRiez2dKYuR8Iv1S0ZUPAxq2
O0lBwFXZM+H/f+u1QK4XPy+o+q3Yk/IO0E9iEYQAjrLGHSbt5Z/TiiF1hQ6STUylhlEnzB3wcJR4
Zs+iZZLTchrSzmZ+lxGjnyha6qG6sXFS3VZwqrDixLHfHfYrDg6Z7eMHwX758bpeSgXq9V39/2Qj
VLt5EfVImylobXy1momIimKlctE66AI9VI/qfzVVNGdqTdcSAmW6Ho2rNBSSHHwdGnwjTtSz9XBs
qSRXczMgrm91fSTBqnsES8Mhlyo2RiLcTPF2br0l5yJXo1U9rnQlb1ShALsqhEWBd4zReQ+wjG+1
l2c0jSkqYQQEBxAf6kGOCIOe16L57KuYqmfifOWox6RaFIutUhgTmfRtcyezv6V8jbCAG4z4KiF/
lYIisS2BV75S53/XdBJjeOVXOPgUHi2bwwFagdmu6NeCU4DsCyOnkW6bLcBNL0AxiSy8upseePJP
g/pPbeRGgeaMdS1F0eAAnzVKqE6AMzkAniwKVxJCCYzYXYpcsaXwWd57AIgc39Ye3xJdDtEXVVl9
of7mgXb9j3xcVBwMbugvOm5RigmKPYzvTIyU6lPQwkLeRFuRcC9ozamI9+CBCZtU41YTy1wNQ9Bi
bq2JxvSUxcAuamt1/zt2qiPZDaZtv35OqZ0pnPiU5yD92n+GjHlztH/dUzC0tpkAFO1h+EwLLXAt
Orb/QR4730TKspB1gl1AYlL3XC3iTIv9LovBzn3BcVi1sZHB/YFdKqm9uCXD/r5+XIwWRm7enuQD
ER8NjT/ISWzg6t9ljnR+E77Zu1PO0z126KqNl2EdbyNlOXIDXVPOTC8BAyOfwYQV2hlSYp1G7Uz5
JnI9nCBlCAxZPZv4DB9C4tJGg2nC1ukKcNwj1lmewLjz/LXoMeqYThYvNJ2wFuA6mEJW/vh5I4GF
MF1KWC7sMpPe4abkepSJZwzguoNxYT2jlD6GHLZiwpvBcHNSV1+NIWG60/luT7iNKAYXtfwBJFbj
LvVTisUq4O/ydIzcGbDxge45fbsNj2K9MSFbCH3ojb77xqEoKl/CFX+08oLLKYCxcGWS2BuiT/EW
SWcwGi8/tnRjIMyC+/BO/mloypXJ3IFghgIiHdkxWbgOGUgwOWQj6zi9t/kCEqx1ltTxjo+CHJvz
9aeNYWyTqAQab3mobA2jlbgXyVBPVfitWnFVNmb4pDSOamruhUi/YP/wugY1pNsF8pavkCy84Ptg
G3k6u0ryfjBGkXi5oUPTF3vRJcLEJbL+BTz0PaEft0bOtDynf4CfB5XbqfFkhvwhatH81E9BjbjQ
M3WAvMO4/EifxYCxEtr+9ixJBhSLbCKDl/ei3wmVQ8LcvssMm/OR8wdY8DumvFWiuoNFAC4vz+b5
GkNEx16M0qO5prcXUml8xCTZy6IvFo06+lfVqfvRWzzltwlTe5VdLduawCtrzRHayHePPIUkx/lk
McYMS3PEA03qUj3mPEyd9M1E2lpfupvwjjP2kfB+25pqPWuodYdspTYj8dV++rZSzPDEb6uiSflt
qcSjo05zykdfE9X+kfytTvlo2sEY9jmVaa/rAu7SmCkOkhmesWqUX0Jor2YG8rdhsBg6YF6aajaS
NmAFCUmNcEih/Y8S/j34lXT9txoP130ZNX/JwbHW1zQDOFxehATM2XXwHGxqP8xX5X1uUUO+oURZ
p1CYQTOLKyOeP0lVWuqDh4RVYO8K0xHn5nNdtgSHJ1w/VFXtGJoWGCo0ZhIPEkT3Guo16ZSg/ALF
zX36sXdnJE9kAc/IomLIsqkxW5iQOQNicuq4eHRJ/oBUjpLSA/dwwnVnBMZZSMIX9Z56ERpdwA7I
HPgaFulD35rvaK63IqgLGTKD+iULQm7JlpXYKPPQ9WXM7qe9CIo7tlnOYnQj0TrEjwj+nWmiWge1
nwDU8+17TGtIipw6qDUOEsfnCXS1WowQVvIOJHw2zQRXIl86swVJP2ETHyZ5AZurbbpuThF8A9PM
sRmb35+ypbrRvC1CgUkrcSoay19y1fUqUwvWX5GXKp1DAnOyL9YJqCzdUiyt8+Ir2TNaJ2RzQrEW
QJU8XrisjnchibupbmESUCqCZNVFfdZlsDvZw6MhfxsS/etETKsz7lbdqz6SgnhsmDzfOMPFxQI7
VzO6AFlEgZTXx+tbaDg8B0YuThLqzgJ3NtOp8gT+oDUTop5bZI0RT+k4HK+R74ghZOYiOODkIu00
265+vugAE/fK37qojQG/U10ncAnGi0r56X3BGtfO8g2MD86tHhAGpMDiN7wOIaVpis/MLSF5EPAG
maWqkDFDwZQrRvFIm7ub/Y7V0tayo3Y/BnfIoxxiwMjGi5WWmW+EWEBKzWZ7jqnbnRCpH7WPL19L
tbEKEEnFU3o6Cm508FUqeyS87OUosG9SwUK8LKgyELgta1V2mtMpwyzK7JWMPaxYJCVjzoOsn/9i
X948TuYUTuLXR1bkiyZnpVb2hAHUhhmMf2+cFnqOKOaPrXUR/+Gs5dArKmN3D4smsURk9EM3qUOG
zu2b0ZXEMTuI/8EWx9mL3WiIhcAu3MyIpE2ABnAIGjFdYLHYN5eLoRIU/haE+ZF1idMq+WJXx+aJ
yVoN4zUZuo2zpamLrqD+sGZcMwAgJ535qeviPX7dBH5AY7IZgf+hWvFYLp88TELvfDGLvoJi+AFb
vJyv6bSJ7vQonnl93dNfziN8W4iOgWAKWoDUqg8o1XLtWWxn9d/awWMyb7A8F5bjO5Xpt2+cSluF
477nWguZBfObEa+mI8zYx0rQyweKaW7xpVy8ZL82SHLgysiaBLpqZKbWgPnIlRc+lqYba5cpHpY4
4RPPDA9/gYORUGD6dTNN3EtH7DLuH2Yi/Xr7zpNHeZr7IjXaPUjL9kBIhICq5bW0rpmSn36cWP4F
A7Nc+eVSvn7uORKiSRE/AmjqAEk9TDlmkPupN+jDef7Aoip7Y5g5vI4+HWSv54zSQYu8dO4hlfNn
2qNiD2cTwEN9TppKRvIMgH4zQ6lHWpWkoQOtwCEepphibkRrqivWo+zbUb5EUUz9y/ITJO5BRVZG
WHA5sz3ht4Guse0xdm2FPT39wDwWtIwStdCVOduoC1CXB2lmF34cyNk8WzkhF5MkgpVVftt10gKJ
AidCjfpH+XQw/eAAigGmyYaKYnCIp4tRUrJfunmWCCBfIL24gU2Grly1Q09D6zVE7RN60bHfL/yj
yVVhXK34blvhJGuu/a2Cclg56CzXBxaMG4nYN00FFSSxPOjfMNTudgMt0ZL/8vzMIpSeWoSpPN5g
2GyLCHnM59nsU1tOYX4XrTbyVEguHRvULptKbRm1/Z41kNk/LUT9b9LGZrYgABFLcCYLPrBq5W3l
EXid7lELBrVNJENkR/3kJGP5kQ5nKg60jOi+RfK6HCExcEzN8z/R5jqnPPgXg4qGFiXRflsU9tz8
fsf5JxDBX1ks07G3283FywD1FnzeulbHBZVBcszkmBR6GbfN0Yb4EKy0FXU0391Di7cYZ1aAw/d8
CFxpaI51HVH5LNN8FfZjtkErEkEqVRJpoj+LczD8AubwSV4KRLqcI6eXdi6GE5jpoVU9EO/SrSMH
g5FtpWG1nB8LDEwNicyl9O3BGpMPrw65BmLjGLdiqh1i+GsitOrc6fc+JQMw00hdFEY7oMDA4zIu
rgEc2MKlcTCiCN9L0In/PhYJgy8cAAbP8Rtou1UlWsI4jFnCozJ4S4T+WNP3AMbftslUZIJ5NDTA
Z7yagBJRwOViR3xPdXGBeffPalPiwznxotAjGQoXCMWMjuYL8r/hzSUsqW+i+lwWNlqrKJK9szuy
E7CeYbBu7AoykYuL/lwJa46mpipLphSJRpWPFIcZyyy5lndVajEIt0qaDB0k+jNPPyrK8JhHUlgV
V9wfexWkE8v8mfLTRgiun3B7e2rQY9LgN2hHBhfD02FgTcFuz5dhNLcWBRZsUxWIf4fq77ExJhYP
/9Ef6IkLvNN9vyRBe6AGxSIijl3Ojwj5C4/FE5v7rbt65wKXwOkt422DhxdHqXoKcy+vWTkBZnyF
y/zQfolFZmJWU8qzodtkSI5RLQjs8VS7yfFjHIWJ2TMdFPv7/Y4xYfLx9zlLBe95Yp3tz9P7EHXJ
du1chUPiBkRWu55uvXe1Iq1C3QNwpp9N+/ikK4KkUgJX2ApKtL6lH8ZN9BzLWjZzvINgunlkjCja
Gz7toFwIaaUrWPr4TEJvaEySWsfLlfshw2zYXKYGorQwmAabvrHxA3lsw0mFhi/kzrXceFfaslum
8ooTXtC+53CeqLjgwTDnn+qbpRVWfmGDzbwMy6sxq/YiZSvAjHnbTOiHi8fDfDwwA5IV061Ps8vy
eEjEJYR3ipIDf1fsAvP0vDKR+ziMTJm/rnzrlhQwtmvF3o0kkBOVKcFh9cjoh8XgY8TSMhSs3S2H
T6EE6A4lCtCTFQAOhz1xrdk9mdhY+DjPnHsUQX7xJ0jtS1nQDagTX36uO8h3QeJeiL1sy9vQBcie
2LxD4XCLSGTMx5cfbMOeLqc1R5dVojBwtrmLqGzWQnDblkH/IUmY3M4awjK9hkjXExq6MZXlnNvv
9+6q/QS+gBWmhyuhoyBCC/yL0cTFzdfnDF5ftNp5FtK1oE4I5TrtgK+yvhv1ABUzq+HNqY8PRcQY
u5SOTIg/+g5CthskDVxgDYSf31mKOwuTCBeoS1X6mR3pJw6frEIuNITvX1yEIiQbcY1otJ6j8c/7
UoXQc3kmJzzZ+/SYmtbBXZXucQJT0sm4GWyDgN4/ouvMAW180SZAEqIJK9BeJXRljWz9iHMzYe75
wZQ/u2nUenr1JZCzomjdCFfidnQQ4hAV7CsKQLj6isEFWQiv4TXmzJ58SUBSd6nMCsSPmkYZ7t7A
Cds2HjsKHhvY5vpTekHEmAlvYIpexeTmYblY9PP2CcswAvJpm0RAGMVg9GmGiGr+1PyEH68L+RNj
V91hDAIgTUPKuoCca2+UJmtkdQbvQjVlQpwbgR8PE+ennnHCbCtvZi7scZMSovAwrqVB3GXgkqiq
ERUnG7EJ4bcsnLkNu331rndjkeF5amuJegzTwAHBaB78lQjG6+7posPwkpipxulUDITcs5Z5Hw+j
KamYiqD3KccaSB5cv4Jsvfw8eCw5yRIi+pPFMRzCPnR2YseOdVSWF+GbVObZbT51p0EP/GtoKxvh
FNaNdt747phHUw3cyhP4yw8nI368dfAIeCidayaeKOEJiSNXAKPFA2HohkK+XsTFFNjzLztCgJpl
0SZbn6Tcf5TxVGZzu5Ij9ImTTzwos/09rBs/xbj0Sc+aIGo8DdE+8shhbRLoN+vzxXt9B1I6g/Kg
WrdlKNq/FwUuZfjFF7pv6yrmUd4gV6YbtO6DyjrTpPyWGiDvfSDWOTTRk/UW5e0dYJCJ8nrgCYan
XixVdPR7jvfg+yHpxSo+CO+KEVVTwUfh7LGYSz7do1bjg7b5BwOkTaAnR0Lt3WHXRY8onnfCF6e/
opkPVMCN+8u3cr2C1a12asd5zzXR+kt4t3z8lDnWqyz6O26rak5onkQxcYajOWihV9hKiflPah3x
J9slFjbqF+RYZ+urguJhjOWT5OrcuyWmpFnpWjs+0tggvy/0uG1tj1tmv5oAPd978FsKMg5IypCm
Iuts4n3bRHuCXyEogJOs2TwY8/LD9xYfQrlrslrTC4JlQuuSemV0jSv7u/LLC4NofRBRPHM/Zfhn
+XJTjSYqffbTojWx6iTwATKLFX4Hut8coylY8Bf+F64QVy0uwsgnVR5ZHTESBJPRh+4JG2vw00qL
Lj2M2OP0tRfEXFd+My+TVeFx06A2zfawg+nWvRcyJz8Jocdty22uvC1P+9nY6zR4QymvFtN/IkZn
dnK4m3J821DYVnL0LmGXc72ZSLErdu73NzcPkie6ftCCzDuw2/DevVYrXe97pNa+5vGlirQRWzMH
bwUmUi1h9HL8lXOi6LhakfcvarS4n8ys1NbA1YGIPcLEuveb3OuA74BMsmxFiO02KCxLhwACUO3q
XKP2FTSNQ3ePzRsYfcUHQf9yr2KNmqxdyjA6lMNPQWwDE34YrH7wKvewwJru3YRt3gonOXYYWGXm
00yALaz5B72zZOzdfNaL7alEiy9RepLH2Qw7p9Lqh4rCLGTdoHvCAwJ3NsY/T9F7b6ofSq/59rOc
Y0WECnq1wt+kHLYygGdFfQfcYw8aYVPndK5b/QXh78G3t58DAXcbgJK8fJzh5ri2lZQI9ZLuAYj8
K/NqECZwugVaCRIeR5aWPsunKmhv6AXweKQy4mMp8O8n7kMKvWuuoogeWyhwTon2134IWebRm1wQ
RXmMs9Zufyk3KMNzbkcgY4cZp5RfSX4gk9wdzYQp/iTUkCF04dKjcQFEUf9AW9o4qpOw02OPtwIv
mBk5pzbnjzuj5CiAxopdJZKUbJu0o9ZDWFdt7qiCMKWEXjbB2+mysSB/o7MldtOmdtOrMkuklUh0
BEy0VEycqDmsiEQbOvE8MzSqBLV1rFJIqVzDeM7BZl/xLGAJwuc5qZ18tkaZ21xGQBb0vaJjsxwG
0y4j5KmHt2NK6Jfq2C7xNLKiVaKNG8IfSWKbP8VigoMv0yDkx2xhhC/uMC1DWS+pkytpvD7AdGxt
FUbX5wbgsNUSm7cMiI/1CoOAdAxbIEbncB66zWTDisAr85Qx4as8OCW3UtMt00fwCX+y0b1K03C9
9dGHzePVU8YSn/KSAUjNGUvCwgy2MuAEl5oSkMLGR10MrCQ/wVqxoplzp2sWRfUObGqYrZqkSlrJ
LQf05+Q6rYvlcTqWNu+kuob957zzQJW2wsC/nlspvIPWcZh5CowxuMt/HiC6MKEG4OQYh512oaga
NkGwISQJEfCK2hHIOxQ0hSMRD1ODbOqlbLl7cSswReasQyQUjPhNYkbo2xPyAYuEVdTPS6svaYm8
9UHO2pvCLMwd/4e/sV5qBcVoIMtPl2BIoiUCQYN4CHmqEYhPSBlufOsCN88sOs69AGVbnYvHj+xI
0Z11NZygagTOKumkT1vvfptcgxLLXvRLd3A2XzMLUjq87ZpztuP2E+TYtpDuffQh+pO101nmO6W0
uMWfLmm1njRW56rrGCNgTIXkU3UchKXPmcy2nOhhPjeR0YUgteIS9Y8XXgPnJMOOsOVCZS6wNJuu
dyA0vQ3gB7w+mPzqDG9pquN3aZ7RBLpNs7JHaIYCFT3O4/cT1HDMRjSaYRSC9Dv0n9z9WYppRI7F
26BAFr7K4W/hRMph0ot2l6VHY5q15j+/Ht2ZR6xbh4H+UUQozvVXiUziFm9JcQKjDdJms5U6DCpN
H2zMyk4PlaLBuopiRQqhM48lPeih/1jEhWvvLlMNsU67qrqw9eqINom5Pla7PLrFYE4U03jkguB9
mqh5/r6i4lBaeby+uf8VmAQIXWHWlBwdniBKWgxRKL1YS/Jtqv2YGpxp+j6iVTu8eexZ14wifHlE
h8YD/LiwX5ouFj6UB+byPIr4rNU+EozVODvZLrZy0tUL+Kicq0JTFFs5zU8TzI5+/+jPqNOJcv+k
6p1188bCCTLjipJdcOgoYr32ZNEzrJ63+Du43NowDLS2pgIIFrAUUQDHLPW/Hbz1ZhvWLgrCZIRd
Sm7KDXzTyWbyMXCc2rgk9TjIVIMddG59DfTmMsWhacMa/g/zaxcG8ervZhw8K2HVqQibNoX4ZlEi
iHK6pgqgTWbyGkdFOQL09eTlgtpJN6HVkd9gCJfeNo4egqO6GQxf6EpDD5XdVUhjFzxzOmEJR0sR
UHkXeBOacNE9phZDTdHl/GpJrnKC7mjbPxMGTzrkU1nqewRNXW2jxG4T1wsMi4qmeXaxFdhDR9MB
oPzE2ylju5lLyT/qFK8Ucj/a8upMm2C7V4InBOikfwfqdlzIMM0BQ/cqk8uregjNa9PiZi6xnL/V
g4mFNffezoI1NtdO1rpDjj3LVKlQIbZfwnBBi0x5IqSc5URnBLTcJSf/n8SLxlf2Ihl3vPCgURgh
foRiEv6bE1IKkGA4fkYTjm31tDImsKxnlE6Ctf8i/PuCHMHAKSRQpEmt9Z3pQEmdnmUU+SBxHw5h
cF8qed35GzvFhfG05dXbccGR6iVi9Wjaf8yfu4Oz2YuTSe+CFiRw+FMnVYDpcL90/R8OhULopHhp
FXd8IZhh8flVDGFpFftx0ye0nN5YrNBxj4rPOETYFF6jnYXS2qBBpzCOYOXYIs3CqfWlHL+vVnk9
/+i0gP95uBp8T3v7u7EJxnj0y2oYhcmqlf0bS6IleuaKqWcJNTiQLlUZf/lZ9okFDJEDwshrSXbK
jzam/5mbtGAE4sRjr8dAzo8pdfJj9pDb/xwg7I1OEAcfYM8swXcHpU7Aif7bA3ow3zj4N8J7o2GE
eHSjA7Cz3fWFb5L1BHlUE1crbTLydoU2ZOwyfbN5YkQf8Y4XKg+V8PVDMLKmxWmmC7QU8CucGKKm
Yb1M5nCFwPenAZfoGYY3YssS7bcRMhlp3HzhbTcG4LhKTQ5rAQOQPwRPXbKtnm1+iBa9hm3094ys
o/N/+yM5xcEJgqL8AORIKfC9+b7+KRiRAgOMDs+Kv3ITeResYFTHCOMCE2l5JIq5O6XNbmFxV79L
NHT9HoY5ezbdqLk46kdlJzsfSsmYgyyx1GsmusTE4qQgU7kx0OpqcXBD7e2granpN/ZBy0eSnGvv
H9yelxWmtrY21mZ9efgIjMdjllTOPqE+PkhPVnM6avHhB/RzjAmaX0PTNIip/jRosPGjko+dLJ4F
2PiBox/a7Uq0N0g10/zQylV5x5HQZSIHdC8/rkwn6epB9qcA/bPzMVhUeYsM3r3/oO2rJ7Z1LaUk
Vyamxq//jqIo6Jy7yzG/Da+YFSA0roXmkDkU3wvM6hQqBAGuow0r/BkRSwFWc4AgPtiEklgqL0DB
hx/6AYuiU9KpTMTPRK4+oR1aqngreONZtY5STm/8OeRhSxMt15JrQHyQ39CyfpKfWfrLuoBurlhX
9Y+F1Zji23mzBJUiFcuT9yzSheukYiL3EFU/Tsu/DgHY+lVqGb2R+Q31LQCs/iD7fpbJ+0dX8FYV
x5lCrTiGwhhPnmbakXbsqnaPOI1wC304WOn/i89THyF/+U4quyCkhs6Gt2YtzKU0LBmXlg9PiVB/
E5k8ZnHuT/OM2ZlFLPdYFswJZkOLfsfRx4xHEEd4SR4gP54qqnMf4Z027lyVsS+gW+9s/oxxOVWR
pN2aXBjMLMpRS8xIwC3GyTiGZ0+rggFzPxL4Vso8T1aJ4AQ6MkHvl05buVhdPWnJKUHk8iUKZ4jc
vT1gDLFgSyGD0cGBjoVNiig104CKByry14bHjhOJWDEm2OWVkMV7T4cQdFd/UQ7aZDCAcgtDCMtQ
vRXaO50VJuJEzUFNEB1gBv+/58DJKQ6g3gweTZehkBgulobNz9Wa+7IPUmq1ircihFqw4x13NfjJ
rXmg5sx8df7lDeptPHudnQLctpb8uutQcsSfkuv4Yi2+in6qfqoC2WT/UzwNaO9KuvqEnlQoMwci
uuhcaI7jBrMjdsl3L4FN/RgkrOiDMdvUrAof5jcNK6Nwg8UVnXmv672jh/3mXkelMIRkClgr8xs9
TkQGyKkKsfmPLOg9qsy0vdu10Ab548CPq492vtE8SkpLI3om7woH5MP0djl05aEUko++zDEZ0pbJ
hpPSU1kAo7UF7EiOBeoOSfdr8nL9u7iHB8BnCt8poxOYNQcUljhmeGlJ7jFQ2u1/7wDKo9HFHgSI
1yTMG45an3HDJAF9Vku1e1dqDH6mbQToSmtSeVGQgcQhYQMNFSs+eUluaPWRlz9FgVbM1/x6x0r2
AkN6pD/OGWUlzSUsFHDmTYvIwbGxG0UW4lHtprzxsA+fPNrEzTQB4H3lShgYufplFtJhYMAh5L/4
pF/qm6xH+AeNGxM02MK6obmGZanL4+8ctp3kNlIBrGXJP3/JPTtDdzfGSXgkYlxd67/uYOdyEVxj
TNRK393jC9Q1Tmoyfrjp4jMDjIyZXQqbJxeq3gWUhyX7xabQwWxBfUn1qS42PsZ9jPpAxEJwQMl6
RqWDl7brqSxuqlJ9NUZ5DA7mVVznhijg1Zz3Dv4x9QkG4mwuHJnfWNhrslnVRN5eg9ZcD5xU1kJ4
49nnqr6ZDOsywiBQmigAhrh7/+kfzDU/w2sheOEQAH9ok9oiEuDvdiIFsPOkYvVRljyo/Y5xew3l
d4rDbYJyXMQwTGB6gGqcHPrq5iSqwhorllokZlP3mZS6hiGRxCQ7vuyYPgAJ90eAxUz2iYtkatmb
+W3p49oCoMtDlsEkJ1Mvxdbi1A0NYzZuG9ssbZyWs8H2Stx9BP//pgFXzR5JQkJx8mjc5DEm0kJ3
BnTjLSYL8dRBtlEqxvzk5CAvDqgky+sgttKOedsCg9Rmpnp33xPd9d5h9UBLguO+AM5u0Mauxugb
N3TzjrQ5H9IxR57xMokgtd5ObkD7A8XpRtsjfGusvAFfAAdU7bfVWn7g6naKaOw/FIChB3Xwn/ku
uVP50JTxPzE06jlp9cOONtQBlbOFXUH5yuQx3tQ6BIV0YBe2dahWXli6a3FqOt9FWVOcyJcTF4uG
5JmHhciyHpIYIh4iYQd7G9XZZ/dtwLxV77YCvfZw0tXXUDJHa+ACwzeAR/UhsQY7+I0f8U6TNBwF
4R300lb0MPVvs9WsgUhpuqpkMWjZRUkAuQT2EQ9aATfVbL9gr2OcoSmDDbgtnOP7PBmj+qd1bnYQ
OCsMB5QZClXZQmVJskEjWx6kNBw23NF2hFQElbi1h7CbBTaSonMeqJON3AwNYYAo+QPRKUosdfkB
3rehNPD5IsNzfX16clpn3nBqZKU8kTgbsYdoU4gYUBTz7fQ9YHkXwdhcNG3UBzPwDUrQh7eQdRAK
B1DzJueDts1l3Cb9t78uVR6WlDQJt71EALACtipKTO6uJVY4XTs5xuZmsRlgGL7804lO5aic9UGH
DDvIi8CHXETcrD8ffj5npwSYPxzdEB615lMMOb8kCX0mWxVxBDHdO45+daUTdmkFw5iWP5j5pVA/
5Xku3vzLF78QwCmrMYwWI2d2E8+IfHsrczZNUjAerLD4+U4JODnur3GtLbrgQvSfTjKVhwqY1e8T
jjzANy+Qzo4A7kJq3BpaLANDdL6m1cBJdkADmpkDAd85kSFkKyum+ZivAuELRoy0hugk3/cx8N2f
e2dBpi5MdwmjUJBg6A368XaKZQ9u3s5uEzydRPJ5Z3UP9KqtdW5aQVNPF9lLmCqmMFkN1W1UKgbr
A7NPcgNpsumdGg9PQRxq2dh06eW7tC20Azxw54QACi7GQCVF8MH6DqXWf5627JMrcfPW8U8N+GOR
owA94MgWH8qZxE9uJiu3HnRbOuY8Tx7sePklsUDLPcnMQ8KwPOLENDZGXTEh4hBaNsQYWBYvkvf3
KjlOtp5tkeK8/xLyg8riAs1Z6R0DmEOh0L6OfRD0PS5NdMi+iEnFx0EJHlFZP/I4ZfxzN8wkKEZ4
goVCm3vgxNq9LvyXEhwhWv7YEt4vBe9UX29mkOSFUvkQWRZU0SU2B8Qx7SAbylflnjCBXyYvdxf2
7tRzj0E0nd33f9mVBA3YjsPnmfWdg+Qq/Q9kJ7THYC8C/2vYe7u+96ffn/HUsmlMBsEVJ4FZUSro
mZjsYebrEsr4FsbMQARsJpCXscMbMxNoxxWUD9CAiW6blj0tXsJ7C7oikgLAzVDD3Vnr4I49XQFX
CJIDpoM52sVn7eWiue6ghy2inlXb7lJ1nMHj/SAhmQZJ/q32mDi7nIwjQyPagDnNY9RNt1f3gq9d
um32hyQhaWwlAU84lTmoQou9cYH5s4kOiWKfraEXZ+281f32hmrEMCnmqFY01lAJt3lD3advAzZY
+slwrRtDxrP0wVao2u9QeGYnAyP7UWsmE+RH1T6QbuYF+Aro2b4kopl0Zqrefftj4rijrjJAp5UL
eMhWT0nVeIB7bhZzAxr1u5Dq2m9R19l8Fp0VHla3CGP7AiRVO5gPETWLkKOp0sjH62Zz/7uvg+nJ
EcX9119H2qqXvDfbNwKUAGIxPEXLFDrRqogh7CPKMlpchIpqMYQYeWy54LvTJPUEYkUV6FsyIV3Y
gfAPR5U8UIjzbE4FXRd6Ne6ygta4SBdRM2r0e70u+c7jHOCJQintLuVmO12o4nMfUcSH8RJErErJ
GoxeudZJc1gxPrvz87gtBbgiXByvcNkDEzny+E4xcQUXb0F4qT1V3f/k4M0KS/ALTZO+pggv4wGT
lBLDyfIxvrD0OsZ7w5N14g/4qY+tWa+2yp/mtUxDrJQ6KFVbRApV9z5UGq4MK6x7rl7Ph0q4vSfs
AbRgOA8YiBaYXOlK+ATQw5NIbxUb83dC4BSrxdNLVyLYn9cLCWNMEA2mavH/bE2DcxipM67Wdz+9
o6SaZIAYVBdlQ7rNlfXIbjwiEcK/YwIl3JksIVknxS3iPISmVZ8m4EjFXfVvb/ObBmAsKZqoNk66
GgeuNSwbhtFypJXLH/5BcKlFIHMtRuO90pUZPlsfRFOySJ8sdJkZzKBSAPwnSt3bztJn/mnm46xT
jO3ISf8PkAh1ZyatsxghASH/OKLVu9O2EUllrcUoOc3VCWEgzVE1aqi3m5vgpZgF8NWsiIzNwZ8L
vBMwnq63LzWr3/OvxumEN0/y7iDrHIFSvNG2M+WLa+qZZTEPV2FtOdpjCYBx9aspTHoSrHuFFA7j
5BWOSoagxvdBQqxz2Lkoq/+ECSN9cs0vus3ku86EQxGIzzGLQrOOqsTNfO/vrHau/HOGQvuJWNRk
OYqz58WaV8sPccQ+NE2sGIMzOFpGSRh/aNI4HD8VGpDcHSuDF+LU9v1Za+h/gH2/3RvELt/+0o8s
pR5xnBPy9ygbYkdX3d/GWJ6NVP44cpO4aCqwWsFsTgJ/UJ50JJvD764RhUQYA5NUxmEHxn0tDL3W
vIdHMFJKQo2nPCVdGrUivgCfc0m7A3FbZ3o1QOCrpXGfpd2O69HEajoaXpX/AXFP+75aPWKmTLCQ
sOBoA+HMBn0XcOysynh7whq40Q6H7FAD21OSHiyylwSUGFr6VE3BCdgoT+xNxS7vETxCyn648ffU
72HtO0loD/jKCzE+zGVfX+Px5Ka2pwJcP1KX/hn41XkqFPtQDIXMvVpBOthTsDhtIabJNjgSVOQ8
c9sRrP+rz+IaLTsqYz0hN8R6PU1W2N+s2HYrh/ecAKx51zGsLATCchzUaIqOn572uIT+kw/0+DGB
I86dG2l7KrJTIkXGpyl1D2o/C/9b8rX5nRkM2zpSmljBtOj3k7/7cuVJ0xX8/Vhf08IFf5H6ZPmD
oWxhHzrJhtYyARej4h5hqaIwF7sRTyQsCi2+ztHWZGao640z0nJ9OShTtm09V+kdQxEnxHfkiYhc
YTPbpZZjwzGQ6cqQcfI0ldEPHFsF5pnQUBQB2r9axXchM8e/6AJ4UUMfmZ8OquDop1lyXrFFkzRW
GZFYpF+rJt0akfi/sJb0dMXWUR+XT5cRE4IQeJoWURf5ewv7lJiK1UAwwpdHbmAztuXPeJUw6hl5
a6E4zYVJZ2Eub7vG3nIXTsJ70AXNB+GD36paze8NnKKPOm4jFduGfppBqikX3175G5n4rJ5VEZfa
nQp9M67PlupRRQWvl5wFcmq/V7PJ2OwJ25UnpDeW9mo3W47C7vTR1Lh8+Yv1cAsAvy7HXYgJTWNM
8DyoavVc6lh9ZRiUuEFi3UIj0zGcXEQkIQBq2T2wvCGeyZJpm09t8CygSvQWggaOdY4IIKE2TfRw
BJEWh2D2rD0iUqZnDv+3+bbL5+3McDbJBweLmKvrdJsOMEehBI6wC3zpty0VKbMQba7sWXEI5GZN
018AAKY+kbwvDRo3LqZChcogdgHL5J1b+YBeasYq1JLaYdg/SdTSDxMmSu04Ei2AYd6y61oIKu4p
guCjus+irWsHdVcQSyVfMRXa3My+fKlU/BGdW4L792v7TzPgGlaJN/hq8LS2+7a2rgU3vwXUgGa1
bS2jjz2q+4YEtf6lwo3u6SRdMTdCfY7HFAmMqb+UJdlCZF/zVtZhj3g8RIKhm/drwFvo0aN79EG+
CNaMXh8au4p/UnKFRD6SpW/E0QcI7eq41tv7PiqeIubAX5TLVjWNeEQxQ/NG21B0CsFKltFYuaAB
tWIgIIRL8aPT9UvyDBvNZA6DCJM6PWJXX5h/xvrrm46sRBLB+XwYepf2ria6hzkXDVWDsvJvbqqB
05alHLilIYhfmmBwn1WO8Yi0V4jxxNn/YSG6nKr57i7wl2V+znQKhFGtObq7yD1Ai/wi/Xf9g+hi
NEVyDhisGaza7JvlWXYumPKNX9j5UJpMzC2puB2pkBVD58nCvmVZhDvMfPohZYASAqGfoGGD1ilr
vaOkY4x2Vb3FLkPlIGsGvXYlnoraf36uT48rtL3lEyYReDVnFTZw/RKw87VXiHF8Q1Gp6jwRDHX4
ZvzteW14mkD6nijoTjQSXcRYjOM9gekOG36xdbUYTSKoVyZmURIjaJQgEDFYGPr9WoJPYDkkw3r1
1i3DYxbuoC+oF8jbhiqST+99UQb/PkxHWxh5H0I3x90AjqNRXXgCI0eLKFFYvLIm/iUGbZ1Y+Sq0
c7Zw6O4Lvyus9s5yUtCfP51skNnEraqG9kUskd4LqjQwuuLEziCVN/q1fWATsOqYTl+vZ8cyu9ll
liLRyx8DEvEcVV1yv2Mc3G60mxNtZmH0RGT21uhDjulPVCFjCYhd/Cznh9sdGhf9n0GhCJkzMK/9
vUNk07PZ3fLVxnm3vA21MsgwpUCuYgDjpZH1RQo7vYPB3QcHEdKRk1MXEtXyfTTCgiFRunYuLvW+
HO2gH4U577YNynxjxJYcIiqV/5AbbnjJv7cFu19GpV+/7hsVRV5ig+3BVlLDRSIztJt3LIWl5A/S
boZ4h0dfDxctbKHAc0BgzR3G27HzeidhYSxUXmyWL+06SEQgoyBc42g6Kx9ftiIdqwWqNHWKAm9N
MJ7z3bbx47EKrAEtcoMdVPDsRmnJ4RXwXUVEorjRR19vyBnNPmJI5eFg+cGAtrdkxFfTLi9sVyc4
5H9dQnkFQqs6nP5mnX3Cp08l8LPzHWCApaBzuxo01Hx9bP3dsileANPf/HEaPLoV3eE4g3zcOwGi
IMzlrRKCb+7ilLXauDAlpcYG5fByeuafE1ZUzBaXeed2DO2QIrOWPojpcsuUBKXuHvCsP0rG1lM+
47cef2winTMPQyjU5Oi4heokG60IlRygFE0kQ6fDWYrqUs/l/M3Xh3rWER/0fqcGaQyiKmoFY6rn
WurIkl4is9ifEJ+iWHOUDRItgpJ53fUZfELr0e52+OQ4A9PfZdmBdAYq4KVHKwAMq08cfSLq8Z/X
sCq7flEx17w+uPx9HEQiegLfikWPqekx+jtAx1AhhiEguq+AgiUP9FgRQUYFMPtgIidNQbRa7B97
B6NuGkbdfmUqc+6/8xNIUWsa3Ta0QYI0sqGNxW0inJMOmLiSIq9oVm3hVi93Eqiyv9LCYzHbyVoq
a3exKqYfCqY5Rl4FeOmh8LVnYdXiHcXMokwmR/M42c8V3DZCOAWwkr1srQLjvbTiBOvdZCemwgRi
KMWCY96RnM8y1VUKd8FIlPE/6jhl+ZmhzDomzyGB9e58/srT74ihNpWpLXU17KPxEXP2Gvh6gun1
uqp1nq6EVWcetYRO11X0//+I63jaRwV9fvrXzc73M/JMISR8Wp5wvZ9UYSJaA+SsjozQjN4nKI/g
nuCjiTDZ7cYscC+fHJjECPlHvZQFeFZmA/GuRpweys9krqNq0717g8WtMq+xAI9IUvazd2bs6lkp
V37Vf6EtCdwKjGIInLKMsqpIMOVK55FBU2P+x7iszJ7x/wXdm5j5Lt+Ov6XF3Hm0KCs8zJPBC0Nc
Dg+oPCwjDvyiZGPsUxeqzsy20V75clBBDNmQq79UUm+jQawcA7g2WUfvxIvgKdMyj0hb1KOTUmkx
BgNWno5Di6EWcugLjD94YouVV0WmRGdRq4sQaU5mvDxOH1D/7QBgBiYPRFgpZcdeIVCWGY4DAHlz
UXoy0gXMXTEc1qkD+sd7vrgkAS1he0ERjl0bJ40VWiCPuUQzUciaZdkN0qBGLzcx7O9T2bGtWHia
xmgX3owpiNfiLJhU2S2lQLqG75Tl0IFINKEsKKNwx96sAnCSqIxg+4m5DDYmes82EqDdUcZMhUcR
Olc+IROkBTXGvMAU8O/0vbL/DzLBanyQCXsAHm4yPBRi0plcjFO50yvUsO1AJi0dzz11OlT0movK
zNx1IcufweUHC9Wg1Df2HT3k3MdESTtFQgFrgGNqwPMD19JVXCvcius1FgGhvJo0DosU/ewCr6ha
vjtw3Jl7IWgoY+G3k1gldHApJPa4eYOjJ5rWeKC3IzOM6Xh/ob+FwBAr9XNa9D+k7QMdNisTWFaY
15u4erfr+Xj12ufaiahrAkEdfa3rXr2wh3BawfvbUB9SB+pkmw3xjVtYqtikUswmwN7N3MuH7IvE
1nXmGVhUy0wKC3apTQnbaufC8Rl6/4Yz7nFEsN+D57yorItH8AFPKxjEePPSTggNX83F2em75++o
QGI+zjD0vRJr8/kgMcLdnVzFSlZ+Zx/Wlo2VRaRtze+1Mr4O8Kfi5nRUhjnnzFSoIOJbxT7TDX9B
dY83eRjG6t5H5G4DhJdBFixkBe7pO5Cw4YWv8fcw84mSDKvfvTuRYIM10kG+fgt8XrV/SpE399pM
TE46gTCXwoSBSGwa42XWkRs+73/Wl5RvHOBALmEKbMzD+oo0EM14Cyz6Cxrq8boeOUbEx/ik0tjI
MCZT282JE3JjcMzhiba/SfWi0TuqPC+NmYgTpObKV6+i8Ej1gLmVkaB2cjTyZlVa8rz2l1JR5TQN
3kDiVMkenxnkCYH6NmoK7Cat6ntedZTuUCDqyV7TWCJslKrbHFjIFSVCrTBnwDGQDv3OkPhuh8jj
IUeDmCyzgHwzwZFVZ/2I1Bva/GmGcuRa3DRgEBDrDb1O0Ky9bE9PrVBs9Y3UQGmCSNvURg1kz8Dt
p/DVLm0KKDUKUAKPFzs6s89CNct1MaMAugY6QOTwzjLsCSDWHr8Y8SgT2YqaSUWm5FsxYc+urrfC
X+ljQcU8gmB6lmiVv6tA0xF7XjAfOQOKNX6SQNafGxXqC7oYJ9eMPKZyPPMbUAKEsDc1gP5NlMhN
JGctwAvG4Y3F5wZ03vmgOBudAUHbKtkPgx6eKi7wHGP9c7Kq325ifi9t+p7+uv+F6698Al0QZ4Dl
7NBi9K4wO9P7WtBqssdlHcVy5kQItp/IdMLgR4pXFDOqEkPpD8sA2ZBID+4c+hFf1TJaF1saihra
Ls4ZOGI6oJkE8jOb5nQBcmf7Gk0t/PXCka3pF4LF//qkOlxxKZUCB13mn/Xk5B8kNXV3GNtBx4qQ
uU4UlA4I613SkUIw+rmY0cnoGDV8kvZXiQjEfVi4jeGdrsiA9bxhQLmCU61Rk0PehE7OlV0GLUYT
kEdyNREisUu87tkmawabzAQ5yc5elIR07alWDqx7DUUtnEUk9Spa1ADT1phbVftBjHqEpdvW7OKN
QdQHqRABxEMajfQSfIk97VdMXpscg3Wbw0aRXx46XJfqfvKz9NSJrxtzSgPCXuPDpVqgCMggxqIN
grM0K0QFcmmqOHf8gc5gPZDEyXsSOcXGMA3BtcF28HQUvGW86sfwd0TmScBeTdWIRQ/zYTgc2pyR
cDVk1/VqqIaOuDKsdjuO/itvBpbFoAl5nJ4OW5fE32TwuYw0NnY2fL49IjhNTbZdUeMQ/tVzFJFc
BllLqLFfsrE4rlcNmWpDpgtMqxyfj84Po7Ej5U90CK3RsBdgJ7412/u9HJ3bkkKC/luv3cD9kJLo
zeNaE/dxDX5IkfwbPD+st+U6Aa8KO6gUbthO2qeqpPwttpon26ORmHmRk72usmo1BJrb6QGqu7hf
CjUq+ertNVeYDCuYoY0YPNKp3rA+sjkohu9yNJCMikFc6kgjapfZxKtEPu1ce9CAwQpY753G9JTT
UZt5kK/jFzcc9zhcPGs5FBwDptnVqJuQ/yVjc8Pgz0Ue3GMvnBvYg3yB9Sx1PM0sd+XUskECI7DZ
HENJkYUXCAblhEEp6GduV+9OdtocFJrdvYJzNQRkbvKWCz6lbxPj38gJcCh0XklGL0JtH05BCJun
ZVJZNTKjmADp71Wdf8wkBVfu7t7ylZBcnRwS3qiNYEFH9d03pC8l/3ofIrHds19mahQ03bltBpmB
ladV+KV86CIac5YhUBcU5EIV3GIEmYJg1NDfSVHcPhKfFF4lgAmSqIZswkZZ+mW9bcH3VaEXLFCl
+SEFJWsgRCd9MWl8n/lXI68O1iEWMsUJtq6pFpCXEi+IFhrMMbTCaKcrd4IVlPxd5rG0LOO8EQty
XVv8Hg2JgacFaTmmaxD+3foJfHYsRlxQCZfmFPE3HwnlmgMM6neHH/mksbsqq0qIkG6NJra4kWLY
g6SFh5QNwNvIkLQquHEr6fcR5uNniqyP/H32GAQk2ihBzikYkRgku+uQ4TLiU34c6ryEid+D3dxo
nZLJ4AQE40EivLG7+oPoHLGngdmcqS1EZjOqawBJvZykLbtcFwLx/eaJRjEsAEdNdo7P6gz2elJT
JdGO2zJ2ZvlfMddlxids8mOfOa7tjFGxgqXeazQgkH59uahSC59HKohiV6qkbKg/PW1q0vApAi2R
Tk3aZzF/g4EyeCRAlAl3DYsTYhquXLEQ0PISxYdoWxoBO1GFpmlcIXx03jWVDfSH6uSPHsIARKcb
486jI2+GQwDvkpjphVtvhaZXStg2leygGaSeAndr/ZbKOUEIlGD/+tWzpplR/UuM/jMi5PxDsJ5e
Pat2PQmhDIhHSPp8nL3Jm0p/Eowhl9bHRBNx9GKwuKvCdrxCDS9v2TmWEZ36aMHtidWa2jotVz+C
gLNsvrtU2iGFJX0Wd7tvXli4JdHkOj0HtMEd3STKVKABV6FKS/DEuqv6hKvPX3h5jUU6U25pIvF7
XJFTiXOBH/jwPWPBXewdMiyiw+chgjPDrQbBNmxo/Lg8qK+YS9aPjNlZPfyavYoaPHX8HXOtepXk
5iBkBdKhT7NT/eIu+2RKvvscAyv36JiM6OxHPw59tcx0jfRk+N3rYjqG33JxSJsO0z/vHuBWqLg/
rh+3oHvvliWQ6SJ1lklO95yuf8z4zdGOC7TQ20l/C3s62STnkIwR4evWvyEJQE6HDR+G7kH6zefi
nOi9gQee7MIRBqPQfa2vABY9+vwmkrvU46moeIYhraITiM/CZhjOAloKK6bXQ2dWj2riIbYdl60C
xbkRTc4+c2dG1e/8A/veWv1icluxUbpP/4HP9mib/Vyoybmy4s5giyfdo7z95aF+yB3XUMOP7tJC
Hog8gRqaFdhXXUrqE0Zq17cM1AUkSckwFcURK0lni7UePTL3A9bDKMXiflkxoAx2xO/uB+0W37Y9
zSIscoZ0cabuYLT0R9JjbO6yEnruIqYnq2UejyzC7AB8bK/1bLNDdMUitX8APsmd0CGLNMXiU1+f
6ghvaS7qSuzzMlLyc/uhzy8KPQT1VaI/EaxTpKMVSviPIe33KA3AFEo2UCvKFJ5Ztxo5XKls1zIo
cra/voi+s2zncUvmqYeAVSEOYegyyY0x672fOPDj4hPxWttEn8BpEydw6WqUc+WqBbu8GTK2zDjA
zLFnlNnTUCEQoErKLsCzWDf7kdlYs1nGRJiHGbU21Ix7o4s5GjVfq2xgQxY8lISJQVT3R6AZrJPu
+djZyYLTpMW1u8OsnUN49hdq0jLaetgQ6qkNLqUA9p3BDrNi8dgut7O3WpSOSmJFKqefjQ7PqJzu
Yd5g3Bp/aPREeJBs/JwX9QDXOYst578sLdUtVTwrc6nN3LTJsVcfaHgYRoM3uCTf6wq1vlq+XOZ1
jJ/O/kNfgJPufMwir81YlHFmxEoFepJ5+WhufUXJTl4h2+28e6Wb4nlSKPdQPqKLE2HErO1UzD0M
2voQZ3hRih79LUWuMJDS/q+j1KRulGXT6HbUAuKMZYCJPdw3M3MFZvuOe3vVcaHdSleA8ypuMKSq
iTUUIpC9XeqbFYsrAQAGHr0b7OFINvdJIelk9X7QOPSsak8sE+GalYv1lSrZNEoP9jGVpG2aGp5K
kf3LqF49W2rn5MILBkB/84nNMmrX2slVVvo81qO+YzK160kWyjqKOLSqhf29aTQdn6g20uoOwmmm
S9MFWr4gkMpSiT7obGVVMte3GHtsk5GPtC0sQMvGl+BbNjC2NNxS5tMcqOZrGwGcX3ZD4Or1flPI
cOERzN9/CMgSlrga2ioUh+55F6x6AxAAjxDsX8aWrZimIQm5O/XoNIqbelzzVIUSiexvs+C8fgm+
MkZncUwbb/1xM0JYPVSQyiE8yvl0bX1xufGMX/ptcknsi1Yav9oqKXHvcFSKnVbnYlQB8ID+/pdh
ozMqerHUhENn1uoyl1ceOrQp75Fpy0Gev9OdlPjSLSh1gGU3VToScig91HL55iqvlEPQggCagcUI
6DgOyyAO8dppCXVSLraEe/Rzp/UIyjN6npGXax477ewRjTTi5Hv1iucqb/s2REjVnRbHekQI55I+
Iwc1aX2wcmxToIejUjQKptk3i7B625s5acfNL8YvhB2edL+6rPlAl5ozZI2eBqOYSIcB5C8Roh1u
ITfdqdSL18GIeRdPEw2tzV+wZvlCLyOj4lA3xcgFIQtTWNLR6E6Ceh4Ax/UGwVcemXID7Bav5kP1
SCd9rxwueKC6tQzL3Mdgd1Bawc9UpQ4M/ailoxmkFWTqB9o5lGnYqVzD6nGFhQveObYfgkPf43k0
DIzlsc22h8xGYLJG9KJdNRXqpubGW0L/SJ73gbQpWHXhhC/oynC4JkjUArmYcR1YnggwNuzC5w1D
eVQyJDQSD6srFB0iGyX/y+79W+D7MVA2lgUt6q1fAC8m1wsJJF2apeeVB+crXZop6V0B4fC63vGd
Gk8nI+V6B5BVuDPig2OzOX6GecTUsnyuoopacQmdd9mQNziGvFJb43DLIm/8ny5Gl0PL9kwtgTs5
d8jALrDmqAVsXpOOB5Ht1hmJFoirrJW/L3r/D5OA5Ch1+iqpM1O6V/h0j0rp1X2m2NEEEroY4snP
iemt05RBpydUjGZzZLTYR5jTFAkSFRbJt9zG8ckMATZ6m4ZGNP2xgNULGVes5J2tg1pg8rk1Pfqk
wQj9HCrbXof7mHeTubJemNX/2hdwTnSpBK9zZab3orB3Hj/kYKp0BwuW0rc8eJudGdzvct1R+pN9
uE0MNLkMpeLqQVhACd+XzQdLCx/1QfpH3j0SJz/liOL+wmBHeQBN7Wsv29/legwz2/N9rDTm8VZD
RwOmz46ASime1x6sL5kMSbsgnIhkBHkik6UiKRauEnut6MQGhI6WrxKqjdw7MAnpv+6v6jBCEKh7
1WzSvjz0IflLpsGzVFhYn6IQF6uqoxHIvoJG79JkgGgxMXQc+sqgsMM316cKVAQjLlPL2ToptQ9h
dum1zchKGQkXIBjD5xiTSbse/EHTBy01gxEpTdXuZTLF5s8syG0NsxQB/N42tIOtELEcHeFCR+Y3
0fEZbVB6tsCv/L0hKJbuIXElOEV4T5Uuq4/U+PygBjngcqQLJUCqLowGQlT1NQ3hyAOJlhVsfreE
IfV9VUtzct9dWa47IiBhfgSFnaTTcTITp9rr3WRJOh68yHYLYyI1BBaYVNvAl7vhXKl5ZtxZOryq
Qk1iK07DQcTyAiemi8rsHge2Ow3beAZhMaUA4PPx/lMHx9g7lh3oAUFCkZuybA0qmTITzja9egF7
yBSe+vC/0sFwTyKVXRry0oqJvy5heEIcZem1pwkT3Ka+Z/4sPKo6l3qdeLgxX/jUFEh3IvCUeQhq
5rfAzyeHRu16LSESpDIsAXY+QpISFb1Oeps7XHp+jLSIFAotvlbdLCQKRmFXhlWNWTvp6bScZIAr
pMmHDMeKaV3xctrHnDQGqHkUmx4naRAFbqavN9ZeETzWdH/TFOZNYotTF66qEnKcO7DCUWuUcOaZ
ZQo2NEnsXl8tPU7Jzk5uICH2co1sQMwCDPWUngMKwsYnhW3L0uDeVtIrMWuWjXpmqXzDxg5WfG76
Q8tfOELJHNvUUMeP9+HFxhGjyGV1iP4qRd6Hw6x2nUhBHQ5zFmkfk3zEu7ISfBJqYM7Zricldhzj
2+mjEHaFotYmYZLuMu8uRNISfHcMJCEpEimFWNEumMI9o0rLgl+VtFMLY/nUDfiXVvaYkJwhLy1O
mj8mAmfRW9ZxGtQdfmx2eFIsu3HA+/XV9MJhi2AOLtJESPWo8Vsayzosyw2357hulG+gMbAILZPt
Kyu7lJHj1ys1ihMhDhp0W3qP2vJMCn0dWAYbbsluBS0vc4dE6icTqICPut2r4D42xYfo/gttPSqR
Cagq1uTXLo5VnDZiQrGu3I8ScoRpSkJvrUWIKgw1A5LXMurAbkqZpQRGdTo8x963Lgby7LPspUk5
+oHtFDBv5M9g4YLTbAjw4HJlxpV4AMjZ1khVA73DPxqXcIoVzE3jIeE0Bl4SYvjIZ9kcRIG4bfJN
Xhv8ooiPu0xWQR7d4hTwhd1DT4K9HVbL38nKKoObaA2aOdS4OJ8djA5wL93w/T9b6ZQ5ONgNpyAp
+ekTQxM/fZdaLCvRf9jkhNi4GBDrc69Y0B/5+uJfmoaQr/T+ZnWJFE7NmZzkP1qpTx17mPrd8M8C
sVdFsibmGA1lAzKJB5PB9V+OKEd1CmVGJDOuTsGynbfXqB35BTBT9hTPLGC8zPpw84V+mH6NSZZw
+FwSgPHYD+BaAV/kldfRENzKC1LHxsxoVPziXDCCcPEdxGZiKOzYSgiLy/GR6Y5cE3hdDD6NF1d5
vld26AbD54wAerz5mrNosCJy/LKON6CNTFpdILowye0A6WdR3rQgHaIjtHUdU4URNd1O/tz8QNZl
P3Wy673v7H5nj+DIg5Sp5aPiMcGU3eGro0XzRnX6bEE6fpUjv/yBQgzCEdOiQaAK1ClEG77vSmpw
HkF1mECFGjprAzZvqfivbFrNOu+r8QX6sTcIZnvK4f62+SUWzrMWsGO5i8GkIrOQEmDzx9/WH4Td
LlWPcbY/UmGc0vkCr5Yy5n5Gq91volPA2ySH4Hb/I3qlnFP6MH0MlYV2YjT6kTnNl/P7H3oTpzg/
Wk04K/PmcdTR08k3ifd3rLsItaXnzpXjwjyQArjCMBK5Se+9pV3Zt8d/Oq59rZpvNJUoMgM6X1OQ
yTEi49qu2Xg7WeMWLzPoJmMNOis0yBVsWcKToV7FAy/nPTHQzgslMM9a395KRkCZ4t0nzbXMgt+o
roY8nMCu6d3XF0Pyn07rNn5wg8DzR44cTTrz6OTCqvAuBmMTOtilkCLCXtXl4AecAje4510IJADA
r6KWPrU4iB5OlWj6MgY9LQChZWB/3CgcrMUtFZzSMu05wUGygg8erAV/KwGI4JqnfUdq+pVRLYF9
DZOjoIE01BhL8mt0lGBSu+nnqQ3c4UUE/lqXrBycbEksaxQ2a9hpn54QmBB7orEPX/MADvfY61B6
lsJe9M6tubh/PCQaD0njSAeXrGFP1UkM3v5veDp4rr/3zbPMBuadTR49vDrpo9iYJl44AB29wYUF
2jCS/0ip2eDePeV24juwJrWbnfAxUk5kkTcFba1r0IUoqDKu9l4sli75c+qu6H3UKDg2ii0AQrnF
ZIPJq720aSWVW/jDv2XjOac0IjohzybNpyc5cElfr8ZuBajjNFZC0q3NT/Q7CDDeSGhhx0JVa9M9
hZAgf1o0I0wD3JoNAMxkbXpojzCqkL2qv4aPqZZRVrMWBB37ybr/kaaWRepHELlL8m6jP0tQzXdr
vy+14uippYUZXjs5SVefu2jnJJ8PVBZ4bkL1r7ZpmHLUn9cOKwr5WpMUbcDfT+8Yi4Pf4vh0FST7
5dH0Lc3tbnjiDni+7fx4Prdt25xLUVcV1AXhtEbBiGu2JhAhT1JFJnf5qKLDEHba/X/Xh8F381od
2QhgkEKZCRcVhddRCTOfP1/4iQXRhU3tbilDhW4PfJFXSSz3lA0tTzJrn4Y4WwqR2hhJuiDMt7qd
9+NekKrGv34nsCEnGOU74uRNnZaYWBwmYR5Cr6VYmhgQ5C89CG2XZbMvHBJBziCynIp6pLvt99bh
0mpUzGyeIUfF+y2hotD1nHzPsvS85gzjaW4X3aIEfpqTpIxGMkL/Usv94ZOvE+6FbbI6iEBEtfVj
GF/bZLj8GxnIZqxpOnxTtqkoUlkECTHHlUXibPfuGYYw6Yaench04OwJx1qvo/YUvyBbpNhVFfx8
wVMXgeHirpCWN8YdxnPYaQ92bb2G0M8siQVLU1yFioLspiEgjudsWeLkl5EyxoM1RCdCqfvIHFTl
eIXHGVc73b6Et2sYT2b+W8jpiwyngo7wLB84WKm77MoNPWYIxzofXE20xpJjGNrze2D069kNe94f
t8CPobH7bcQYx9tJSsUjO84BWp4amSs5k2X2WIufm9sY0O8NoY4PxKMOa3VqfVtIToIpl7g5YMPH
5/lx77z2CPlgWCmVn1RM92+wuL38PMyc9aQRUxPs5F/+f9LG1nogtUq+KWW+14aJQEgzLCj/OoHD
neURG7FqcGzfAJSsNda3DKrUmWXMrygxxtT0/B6nNtYTAH9Rj6wrl+WzFowSRtDV6bRR2oumDgCe
EknvNHiLQkpo7bQLrCzOvC6taQwcn3/goD8FhWeb3ElcM7uW5lAn5BeU4b549A86zvCau7Z68uf5
i4Y1MIEBqxDAftEMBjOQ2YO330vSv6g8QSJWUTR2Ah18ImHh6NpRmb2s4ETjhtRjDTFBlgMli9a5
+GxXHtAYhCdlTD0mVUoo/FJroXECJMm9DsZgBFQWtNfPlrLqVvazBt7hpYit21fvUx6Apgu1Fq6W
rQgq/FCkvTiOvTAkzYe5z4sXCCEDpYVOVMIaGlbzaj+5qxug4xi5DiaXqDBgB8wBxCG9zzEfSjn2
lEAHM6xLkpqRfhM3OujBjJwsCKKmkvfzKOHsw61IR03QFLjUSxZndkmVWGCUMURcpaSOuFlNuKkE
r3GS+3uchqUejKbrc8ekojzIWNs4Cm9RagWtacENYgoE3bJkbv/Lz+XTG9i8sUPU3Cl3xQElqv99
CbrJy4qzQXkR+/a/P5RWYqFSHRnl9/i76w4gjhYN6dsEPk6CR5lWWMkG7LUWXnBKLTFaWHcV4SbQ
9CvYxfiBzZj42PUoHyTZb6hxe0LgBgjCIBmDJGrW9J0LdmWg2Ygew9JPCsTbu2AN3uggixARihkc
hdxKn+JMRUfTNYgxzm2/cb0WQXwqtCSZx8JKxt/rgGyu0i7n8mm0kPxd4vLRO6CP0D9y2FbPLLfn
l6oA0Lrxv07txy8L5abhkHg0ysK4Iib3r/ba+QJ8VHHiMtiJQGNcRnCk3WuGBmlKnHQn2j1GVm0Q
qAJT4xquS7r6No9Yn0uUsXZc8fUepDxzw0S7c7m0T5B6cRGJBuqmRzC+vdMj+P8bpjXHMzywoYnF
+jVyBZiJKvSjztXVyB9y5ERdMT6UNjgLj+3Mru47vgLnc1VeHD9TnjvytHe0jhuVrYBsxXXtfLQv
hpCMaD+hQC37vxhpFQFngVypYSyTcJEl8WfMpTBwzh0jpRWuLi0VUwrGX7wpEfQB9P4zyv9z70SC
B0ZZArcAr79Ywcn1NQBuvFrUGAmAeCfeCDXfYr+lyfAUV4ZMjGrsD8rslaWYgjjCfZZsqZQiQQ3R
LMkM3csWKVW31cOqRbXrEMvdf4E6dAtx0guU9v4FHZszr+zkUbxm8E2NkrOkpknJjm/44qSLe8Nx
w1GMAYmIWP79SevWzV3ejnWktwue9Y5HY4+INR1QefBWUb8POjKE1raJ+JhI5NIOiXFZHTt4ea+U
kMe/weCZMCAGYaDxnQS0iB2Bc/QYPKUT16Pbc3d3SoEdQaXL2STQTSJ9ngPIYXGl1ppcU5PGaxDT
0KQm5jCMf8f7VC1OXL2xejbP9aaLX/CtqqdNjUyla6sFsGe8thw/0K7xQ/svaQWykNH+47C0+fIZ
nHb0wrRSlQ/g+ceGduUUL7LvqmfmwP9BQczjTERWnNV8KCprI0t1NoU9yHVBKviemCBXCzUj116e
ncnYeOj+uaPJ1beUAU/ltQSS/ec7G6fovAIXaKIn9VxWQ53LoG9Lk3HL86FYgTvd3+CwZkj4oLs1
QDDkCnr+P+npq0aD4ZDBYbm8fBtNw7/5grkXMvnE5y8kHrsEjqGr+ez817d+IwCmeNdWezKfSuK6
9NCxXpEs3SJ0UTZq5tbYLSOUi69ePvQOt1rpcXqSIQZ7yL5irMXRpCVO8IvIF7+4BVW9b6qNDAuj
YGF/pJwcakpB50XURvK4LG5RayuV8mSDNmpTFzeav2alcHp8gRJzY57HwTKUlwYv5D13cuxHSR/a
eK2mhgu5P9YRoT26d20ZiuR3+29xR7ilUBEFSdJa4mNCgccT55K/MREswH8kKL+FB8Fs994eQ75u
UKDD0JmbFwdw+5cl3B+agZoA/2sHCbQbRzVo/pxqVXG4O/ooc5fxPegfOlswGfQ/RVwckG9BMOhY
k3ZT3J0J36VPA6WOp9ppDNkK3iJD2yCQMgSPbnqORyBMqVfTmPGEedaBpHQxQYu0v4WVya4SOO6x
jUsQoAp9+DuUWxcLGBIXt3UuR+xohaRwbnNJz3QvQ1UiJeMcFwn3JLkDRyisqqhw0nZ3fVJ78tcv
hFCMoFBOzyd/ssY0fECYu+zUZW/bbuhloZf7QKz3XQ4HhL58Ip751U5EL2AxgLJUu6imDuLUpl44
7brezk8IFYI19T7hXGXgSylYebFNPr6rzDdBjfqv5i3txDOWKA4s29CuES0MRP0WXjHb5YqPS+uM
mTx2Mi2JKlBwI9EkBPjflbiYc82t0PIJ+7CU6fcxjryqsNwIm7b8PQwB6B0Xi+rAC2Okm2gH/vLR
s7JY4J8fU93uXjnyRKCWQ88OGYQgHSZ3BDXICtLAON0s7HRtKGLzTyA4RSKlH6u1sdjmbQcuslP8
O4wZj64l6xip1XGtocOzptVuoHPfrttMxmQkVa7tDZS4AoPZxk1sRjLkTRm1PNr5wYu4rwJW/y8k
6bAxp98T6SXDczasDOLbelqW+9xc7+zGcfakUCIhDUwQwWpy8JqT7UHGeLDvuitaRW+8pTZ2FsRz
j/PJGn5hddjFDkdu0dNrtBNFh+Rzj47/dGAiuvVAzxVdII35+Q/D3P2CQj5gZsLWfsphrB3sp1FZ
Q6LoIl/L5f0ITLTuolTEUZmDTf+QrnlZW03EQUu9PXHBuM/DWDqbos7FjKX6vmklvpsxd4FA8eGd
pbcpg2j036qa0Tzc0faMXGSgjIE0DFrxX754YN1YdTpXZ4w+6VdsflXdsMBmwjUhwamsZiGjkH72
HxV3sJ2TyklH9ZuHQKQWD2JsT/DXiXyyExzdGgdPnBo4oyEPVMrP2hVoalO006NvlSz8sHX8pki+
iTlv3Q3xyspFQPYdlqjtYNJuvfq2wY4k3pcB7/pHHe4sWaWEXvYtq3p2vpebHtiRCHhBLHs7/6fN
WX5BZ1a2zHGSYT8JjZxRx7Hy2TrjU6c6HfKDQcI8Jyc7xgv76hnMe9g/hG+9LCoOtl5hQapYL4Gu
pJbhUQ0jdIKKSTntj55GpMZpEz9KjLZgGlgeNd29gHumndbrNQAmSpQFjJf8dhZz3Mx9Wfjuw4HS
SYmPWnMCWQsjqBYW3+sZbYXimrVBE7myOhLGR32same28skJuHAqBJ+Bhc8PGx64IDO0RB816G/m
llVqiy8c5JAnsLv52HRtlpT8c/qyH9BGmoWo+AEcDH4+xf1Zs55wBS99BDz3aHveJ9ah/KCW4WSk
jY56zADKCGSECqVBNCS6k1+vhja+Mbfj7Bi13S6Z2I7hg2UUYaGfscSVi50QZoypLIW+64KCRksb
fl3Kt42nRltA1sxzDi1xWuOryfVrI2LFCiX/FWd7GBigv2U3Prswh+lN5YBmIv001nQsnTBmonDW
1cvXW5VsfYOPpppgbrLcmBSgyk6Kofo7RP+uvnH1OeynNKm9kdXgL76JSIxdNi1wwyxEAyO8bzcU
HsUnUpHeymZW6HOBPjYSWFfXY+YEZyAXGbfY+6Hu10KgdIef7eyAJa1tU/BXjLplB4NdQTKuCD9f
5RwftLuOWeBsThUnqhbW1/rQKNY0HkydCBso3KqimbXQYE2jLWMOQqq8pm9Jp4+nrp2nu3D/A0xY
Lbk0u52NYcjvgIPoN++gJFZ/CeyHD6WQOW8HIN7Hz4ciy2WHECB2H2uLXMnvts8g8cdzZP5lwT3z
opMuVf5UtrLb63RZ4Jo8szD+98q6KJCZAxn3qSE93PYGwvLYbsAD9/obJ3Z5zOjpT6M+QRgA2TZM
naxlw6GWtqAkmG9b2+shWnNC+1c3OQGXHZaJcYKnCOI9MrIN0cirkGNtFStedT/gS6mTsMg6NJUW
xwwNwFOat1jaRNVkOFksCs3aFUtiXfGbNT5SRFm0bJP8Jh/+NMsknpEiSDHPx7bEz0vLv4YIkHqe
pSR8iOnbvlJai9IbYa2w6VJecb7oZknGj1N9MBT7u7J19cLcyFcqK0/iL9/oRwVyhyvsfWAYnGYP
kygUp1QFn/wHDFaYzdVWIrzBSOsDP9n/ylD3AknZbgLAHt/SMs8skSC3j1gY6ypx3d02QD7sxh21
6nrCQu9Fda2sEGibnAo7oo/+Yn+vhsy7Llj6DKcw/R7uukmjwvRVolOmvqBYpt8wzQSfytVPHX6r
f5CGru4f6hEt+UyUnHDSBDsG6Xbmgxlvrx7IBS9Dh3QriU6Ek5KrF1aJgsotqzO7WdpdW0sXiTQo
Oiv2cjmWx8ycwlFGORB2KD2iQiET6cKg7ibNRPoZeycgnwDrZpbvNpMVXg1fkLaXF0qTZobpRV0u
ZT7hyn9MfT5OWyd16+YTsZaMnRasxgzMXFgl8JCCraw24fYCtdQ7iwYCQOPDlEYXmGc+x2ehqR89
EoazMwjyzrFe5W1hIBDP8lrt+saJinulRNGyNALXrmW1tcmRM7Cg4gzrx47oT9PdPEWKcv4S6bTo
frSs3YPk1oVbPNY6/sq3qa+hI2SBH08XbRz5HSyvvqHrMq1+8VINUOlAjJEAJKWGIH8wuwJLK3BJ
U11GmVzz1gF7aEHaCVr2bRdbH3MbcPBXkOVzUMmqh8UJ8ty2OqCsY+kKO46c76YNbT7lc46tH4i+
RDDxCC8GHPHC0HwwYJludGSyF903BCTvK8yRm5Rjw+X36cmRtYonsq2CKGQzLZLwdlYWsHFQQFuD
PvlgQOVs5Dnm2JIFwkKIY7/5XhHtrZGqxNuvdjy1B3iYjMHnd7O2PvFcJopBQNuQi/Frv4VHQZhW
UJ8qTCNjvVlql4wUT/ZcbWUo7reYHh3d31Pz3Le1S5pFtEmzxsvPUqmcyLgni59raaffg8Ox53dN
bkuCtv+fFy/y4JoL29ebF7g97Av6UIpYtyraHmwdh+ZL+NCHUpaFcDyfeLXrc6y8S9g7XBDN4KBC
qMsql5son5nLhu9QwP4elLATtHbRIzoEyBSz4H/1pN8NVeDzx3TtdbpPGaXuYtkwftJ7aavo5TND
asr77E8MbXI2W2Te942F7n73dwganKrDuOt1VOL6s+g4emXQVEcp3V4vc9kkgXbD+VwyTCv0mogm
AakcqoeXCbRIKn1zk8+g4Lf1Eh5lQwzM7JrchL8eDv6HP/zdNI9+nnQ70as3+ESXNtAq9Mt3E9GW
ueFcrfAg7o1fLM68XQzbe+sMyAMyxXOo1Fn/lZL37R5fm1msjSA3zQCBC8OfH67bAoLXjpxEZztL
0Qp1ti/2vIHEqtmZK39xmzE7OebhZ/oojoTTUAKoVtkzZyI5qDmIt3U9/rKJjyzMl1Py+rLUNMB0
mpp/y5yDSY+9Zp3LiQBUkLz+Q2/CAWSMuyT2fOyVYeFnmpJ26YX0x7wkE6/oXg8wSVS1wEY/dh/t
4h7jQifIyv8oAGumSq3gkDaqfmDtIrcnSPnDnBT3AsejEYH3v5tbgtOJMDBHFKfGT56hxPCkB0LQ
ACf9wAGXL8Vf7o0SRQzDqqFVDi1Et70Xe5GjgL3p3VxFPdSsJzezpVVlbCbdVNHMCAsyMMx1gBE3
D42ZVur08bgx7moYar55kwob/zNHvFC5iZBIUNgrPcALCMmjGHILM2nywWkRd4aTAY5MGmlM/dGq
C9JcSAnfOVSbnaYdj2AU2jJvSpd3POfbOZvprTRCUdSrk280oIHLhb1NMbY/zsIY8KZAVOit6lAx
4t3dne8p9ac3eZrlKNjTx09Ck4ZSx+WglXJxEN3at68zqoGL8CcQapi+99EK7CEZMGzfYLDM+50+
PZz9r6pPNsMiVKqARJOV5XotF/ca6uN+EU0FqnXaH8Sn7l0Kf6SoaxvSWr8A0ElZT2geI0ZjcdDu
dlNX4NRa5Cinh1aF+hJLD1/s5EDZ8JH7Szbr+NPM2lloEtIeorAZp3PLtEXec5GCRjPfB+alXQEE
lACrVaXejkfw6pXG+mJ221T59O1KErGl8csPTgcZa1TZjFgLP6DiwS1ifgcKgCHSv+/2VB3V0LnI
zA867ZORjYUhPLdGzCuZodFzdq186+tj4WXU3EKm9mXCrXao6HO8G34I6BMeh/2ITw26RmzRSFYh
nllEXElcBeiS7AuCG8Dg6VLosf4qXudvx5++KsKYSRdzajPzKSC/rXlQ+HfIpJN8/Yll64+3cY7E
Wmk0c5SffrdQws6BzR0MirWigwMUUZ8HTee7ImpHZACeVUaHVL2KSb2H/As1k1buAG4fVOp2WXH2
yqShi+Q6IciP/l/SbM0EIWUXMpmTKQzmV8g8C69+3277w8DTTQWhw6WbE4XsVVGC4WhhVpys0K9X
IzO9/HqOMld6tpj5RFOOdqYDWmda6VHMElzudXyRaV00/7ShWcs/xUDLMJiqkq4VctRNthHxPDBg
U7FPD9AR4vzDwiaW5KERYSl/VtEJkApZo1i8acRsmardygMz11lw3SU/+4IxifnzTGv0zZRkdM+M
SKAm7sAOZ/VWA+d2haDfWGvxyk4dnsmU6vnGhYJ5PlP9cSVImr6ZECPR3GzGeFYosw0yDSNLkDzE
XnA++qUWGQp4Ejki2Vm426V80ncSFUO7qDsgvMQgdR2M8//dV78rD7zx9emEUKw3vgbZXTwxFIC4
skoBeaNRBgEpiqwhpo+U+59ReFvDp4NmhPtD9a2JXTV52FW9sQxelGb7N6MTMzT0Vlx4H61edGGv
oeOwC42hXDzw7B1SxuuGeUKGVieNpJOCJ4OFHujkZ9tcjXzK8CKlQOrVCbggDkNZcUaYtaiOnrVo
lmER2qV4oeQjhXVxQj4zHmNhXr2CJQzol4sWmh6ok1jt/s7pJroVPke2twPIBNXjVEAwlYFQGmgH
TRT8hzYs0jxVxrJY2nYKlsbxacsPva7Ihha4KwdAP6+kwnZcwH1+O2oMCnmbHn8NchkWDOpQIojE
9WmA19GKL9ONJMJXvbe1s/3dhqOAYHjtuZtCSPGkvWVL4LagkKIzJYFKabIQAI7dia+loLCzjnak
kD+YYUy78d+6cbI0vZOaAbkKvlS3xdloMWnRcbJj8bgK9J7+ldv5Msn1vbmbapAFqXVVzN5G1+3Y
UFPtNB0uu65MtHJu3ZVsGNqpq/sLGQYzCJijVyL/vimTZ0fI/NldZSMbC/46/mI+uqwPvIjuqsPY
oS7FP7OIaWcUWEBDA3I8p3x3zKZ3ILHzYgh8qSSO/tgLh0PGBYBHxK2mIF5BbAOSMmRo7ODmY9/5
fodr7Rbu9YpEL7InqgcXWSdGmf8AjPKRlckuIOSDq6pS7j2QnEwcoGMsZrZUkRwz98HTUwiSAkvb
r9z+2PRoBsGEnt5bKgtxZd1SL4Gt6yS/oyTn1FhWM3fybFQYiOisD3MNMRnavglBF//G70YlhVJs
n28TW2HLP3wtqw/AACvnCPsSFWIIJhBKPu/tk75lYNC7M6NY5dMZm7tHweid9w/kK5+v7YSu0H3V
lCnxeLEV64AkVqqRtEfxt0/FCR6DkSnOU8SszJsO9YvVyspFeMyzddouB8gb4zG3Do5N77K0oFA0
qo2kGnsMhgktDuLXghwVvOhvp4nVcu00LoXg+rciYzaXQe1L8XMkPyD41OCb6EsoCQweJ1Nc7S8t
I9tfxp0qiaa3pwI/vuwJkvCfiUrgQ+rqq0nfrPiLczYH5roT2S/ZZVI2r390v9YhgkLzri/3iqaI
wvF9LXMmO5HJ078EPcTQqVIAxs8rSZ4LrDsvdBxNTP9YiywLsRodRT0yf0RRDm4aeNnE85KW/zhB
xVn/PMV6wc/pQUyCJgUGcTfOIZhe4ixddGr7w+ODYeA26lZif5qdgPO8k7xEhZcZ7CObBA2KttdR
HW+WQZUv8d7h3e7QEhZs1MNIRRKUj2YesoGyTQtIVJPI2YWoDX/2ZALNk6/H/ZLyqIOOBvl9/GWJ
RMyiH5irDuvEriRTck2KBN/kvemdrL8VpmAWWDZ1u1Xk7cYDoZdBgYdmjfsHpg2Mj9suRz3ZuIhh
ZpwSQbs1ZyRNALt/g1NX8q4XpKGxpTSJy8/oCYZhG+/7a6E2hmNcHDshJiV27Oh9El4f2X9woiS1
SXKpA/vM0H7VF2r37am+jsbeFvwV//+RP5sz/K59+EoJDeVBVwBPRxWEhmCfO97eszjfkpbSrsUw
5XfqhLwudfOQv7/ScxTm9S0usJnTz+mKhQfYs5mc4AycalbcLBF4C2QTJ4YQEoaYWtQPvlKDUax8
0PHUjYdLRTWLU1olFvEmb9BtD3XscCbnSx2/tTMOzE/cpklH81/FwZO4UvCm3HoMtgnqK6Doldyq
R4JTJLG15dp3fjl2paQXRLL4yL/j+mWOCqKF//B6mvKmz93wF8CcKmCUFI/viWRoOhzNl7CxEEFN
+y4iMtXMiVSykUqQ/V6R5ZFDYxAd/RYQksCkw9o2NVOgRrXKQ07wBzBXmv2xN5PNVOnyOQ/Xoo+g
awE5BvXa5iHn9bDtJApLOP93bWFGHh9Fzc9bYFslM+r4uyApP9/oH6O+k0PHSVFgOg8B09/Z0WAe
NnN/gu5x7qVcs0XiS08X/4WG6xenJudZPgwB5DwfMDm6ZvP15Oz8YxPbkTbm05pbBiOKnU5j6bdd
a4TPcgX9ZSojvg/S/kmFROLYenC66Jf8qnSgeAZwxjGgoHZeusw/Xy+mtxC8YGvs2vntjvLiBII0
28bnE73xzyfFcC6BKtOpltQVcbIyjSNrrHKYBW70WOG0btKtE8fRFRj1RCahJkRZHQb3iudnSdMS
4K2E18Uvz+dcSDGaFYow4DGupy/HGY8XrFbDOrK9zZ8iNL0JeFzOqeVEzTIHuicj1UEsmigGJscg
HlZQ0w/+cVzaQGIKU64ozFvlHyqdHJJulrqc14bzROYJxg2mFPSbJIJb7AqmaoEVTzJcwIT9Od3r
fBGKZb/7Yg0ul8Py7Jx+ktxOO7t1JeVl0Lwf3LhtG5AXopjmSiSUevL/eJq8wutaA7R6gOmcYIjS
aW0FKAYuFdmRhqEgwYxjhAqyU8VGKZFfnLelYfGkT0Hpvk7cc0/tIeWul8sH+j2nrRvzfmRVFxSC
FgqaFonSn7h0O9HxGAxP1+koMdRba1Kgki0CLkZapYL7cuYZ1nnP3XJw4ZFMAxM/LgfpdH7TXaN1
aSdEfd/UapIM/0WGvYMYbtaPO0G/roBM/l2/MWLN4HoXPHf4C910ippPuaQmz0/KxFzuXo0vM4PL
SfFO1pymVrSjmyzD2nfc82YWS3Sp5B5akfVSIcjOytJE1vEr8Q2/AlSQcaOyoa1D2Nl+Esq/m0MJ
KPN2cZMpVlwr698BVzsp46wyKypHIsWAoou3LGSEDrAZdU6/pKG8rTY3xfjCISZplc9icZfpKBxp
oP/PqdYmE+kiO4d06QUj5aB7eLg38PygUdKWs6gkRLqR1d4aSeaxjh3QIs7rSisKdfYAh6ez2vHC
jPNFW8BPBRQrpgSLzMrT2P6ueTUzKiRlwo8IQUrvjbpr2LpYlfgS/Zix3M5pd/A2TF7sIdY7nzH/
7TcWypeiABYtv5kwvxuEE1zIEUoxY+sCY4uUBzHY+Deec49MHYu6DocgTiEJSF9T185+3eXgkeyd
KgEgfD5tyhyYyLfHY/gEfG5EuN5YGBpiDQ5P5elMVH9jtjeZ4fVd28vnP6gsyeSTjUTMsHSl9u+q
0WzaKUP8GVr/p2yRZ4p/brzl1dXZgxwdz0v1pecAmcXf/oPTsmI8waLtbpd7B7t1K0wn20S8eZ7D
e1nEn5NdPHJ4cuRL2sCVJlTZrcFtfSv26SjgUDukM/Ru16+Sn0AURBNZtDh5dv9RUHalTYq5nEm3
qYiOnMtkjxqUz23GM56EDGwNMPI9Nhx/rug4Yzs/zC9AtDG6car9XHy3z1y4+XMOgYYyPy9EDTcc
Szb/VHdTJ+PSz93Ktx28tyiZ38kPheaOO2JGIKFozS0uyUqDpKuGbRYPaN7d/cKR9eGWTuM4uN2i
kiR5yjt8CpbuiB3tDuPvb9OsCQA6RUuanIEtc/0r6gjRiYsFPmEbeeJNrx4ZFKbl2QPb18m6jgvf
xdR/nAXPWqi3wyKCBxNf0W/hz8woFy+hkxuR5G9jWf1805A0vwW41o9ahav03A5V65gV2ICjZq2c
F5PbqUp79KLkK2jLkr0m6vYNwmFBhnrQdVewhA1Yi1iwZvppER6z32tRbK6pyO64SNgB02JKZUu4
AIvS5z7bh0Xu9DykrApasGoVVGOwPh0nu47nL9djpqG04uGi/plHAxqdcPgwovj2AitcwA6QxU09
Yp8YUbyA32Vdl0EA4WL0W8hVi32xd0FE0Paw8u8Oq4Ore9bJrASiiLrxB307AQbwvUV4bEO6IsNM
aO6ppKja41Iyqv0z13mWMGKcd/LqDM6YdITkf/TPuUf5IUn3KT+5h11KBcuJEqB8TeIvv9PE2yO8
RegR/RFbbRHIr6KACGn8wHSwsTtIZVDw+FtIg5CVt6xP/wf5C73AGNtYd7gZ5kMG+4b/y50hlK62
+bXb9V19RxnvK3/UBiGYAqeiS3G/cOOgREtoJvCZFTHbmembFCMPJ82o+LdfzydZqrdXha4lQIH3
50PvL+MnWe4WlXmF8jcwuz8KBFtihxK92EveU2hp7kJZ6z+rWE5XmnkexuyfjmV7bHmQXiW7V/9g
txXICeuOMOclHVUY9qkISy1fbO0DUeGrij3DWCGEebnvwfnwkwDP7oqs9eMT063j2GJTF/ikSx3N
Wxn41UobsCpPVVRuTzypiza477eHr7YwH95NQeKhLDDQGSei7vb7qd6+njPcYxJBd8eWkn7TDt8j
3BVj2C6UytPQbCorR1V7Xa2rGVfeO4pdh4mbyDxSPnA+2Eam8O2/UcSHPkFEKAfGKSjlD9Rr3OLu
4vqwl9lJ5qA+vrpHia+R9q5JneoPIrVcilWASuBLoFRvhxm3xcix3b71qp6qE+XTDr3KcohSM/M3
xA7lkVfsfMcjRgC+sg7kPk7JUjkt0gWiMyxnfQVXhirOoj+TXCgyt4eHjSOckFFvD7DpTHkHFDmQ
7aaRH0qx1pcDP5Vq8nzXqfdHkBWnAaQcMMLB1qh0ic8reev2WUAKDcMx/kj1RXKv7qx1fga6P8+R
U5VUSUdnXkPWEZznmZIEO1/+RUz2VLfhJwEwFQ2mmkrtIQDiogH+I/8O5YdVl+Circ9Ft44kZOHY
ToFjTk3zQgew5rJNcHjzR6HEfNWWz1fvgI70ASH7in3wdmfpC8zUCe/Amkq2KVOmQt24dOgjqLxv
z15+H/8D8yOdCAik6hEvs8Tb4I9zYGGXoB/kIKQ8WSHcC1FGmGzkFst7OornfZ8DvPWg0otKXr0p
w59oKviaDxv5MzNeW2hm7FzQ585ZQBwomKu+zoSm1n1jmAwvHNqQHFGqkgVxxTHAwni/0NiOYRP3
UUqVq9pEMqBzdQdHIfWTs5h1KWlKwSj+KC9g/5/KN1ntIORn9URLA+rp5LMqfZOalDbMC3yyabaN
f0xOwHJu0LHCYjGFZa4VDcgnvVbKByeyl5vz25jo2KoWfvUZxK0CWquuZAeCVwYjeizuq1gHJBSf
T08posPD3RP0hCG+IlrUyOFRYMZYK0xjJq9fz3O25EvGtIkbuPr1o8obl+FiLKcRiXykOzU6KG8H
/w7JOnC1n6MQHYNIIuaeO970agBynKe1TvNRDIh8il+JHc7sZOL5t5d2tvRlW7r47WCTsChNGLuq
aisDRca32S2+ciQ1iDL5bJ+geCNWF2QxyQdE/WASzBfojaRM4pnqg7586eHsX5CqhvZju2AXBwH2
1AmnZ/kNvonlSPjaB6xphqDEly32xpV7TGmqvlTr6+LVs+J6HR4c8971O64yUZz0BGf0N8OtMIET
ZHzegCzfoabJrPfnIC1jZy/oU+PFjljOXOgsDOQB8uO38lb84fgdMTXW6McY7Wf+n6vLbBZgZKs6
Ok8eXOptqbJe06iB7cODJeUB4NxVelfdA4xRCaS/BmhfM+zM6k3QWoZprqpibIZVaoqmrW6D90wF
pFVhoWqTzAm+KP27Izps80+tSZQFG+GIyOcmv0JzvMRWpHVvj/6wUGgUHWpFoUTQhjESrvd8fjOx
IG4q1kB2KE4DwJAVvy21qGq6l9Kl3EUgdpIjgVJTh8xACSes1daYQ9KWqY+acvMshUKHpFjH/x6e
fPhO91gkWkVXQl3oeDjdorcKD/0TNfrVtQd6GFtLy0YgBdFaCSEjRLW7zzXnjO8v9pzJtjXorpD9
glxnmjkEkyA/ur3rQdE1CFRahjxtHk6Vkkj0ijmAj+dpqw48p8rlrnQM++JsF8LYJ41Y8sgA7o8T
/DOqErza4+luy13H4J53LIYqcSdUfSBM+BrHLtx6j7FiqC1by0GILB2Ir1StVzv1g8P+87/j78BT
uf4e1tBJsnwdBq+XeKOAjVuVzT8JT+wpfY0gJqf68vQQAaTC6ccNTIwa482iA7RcMFzf9kMietFz
aiStVUUTyLl1+YdYWZQjD0vEFTajFuVhY9N1YISmpj/sa5ndu9DtvvPD9ygZAusPBi/TLuaSswB5
jo5JQ+3fESx+1NU5rzo5K9mLblXNN38jUN5Cl7u4Mvp9N+nprwS62H2ZIujmaytHtqjkwTlMzzcE
asGvyyTmnVd2bWmoi3QeV3gtZAKBFXKjIzcaAHFfqGEExBsxXY5CHpv1uQlmPakgI8vhOK9wJW/l
hiCIwzn2NGaauvwutMMfq5By7c7zuKivhEJRF/ssMmH1E4C0ANrGbcuuoSqQSXUuTeJtFPe7BMf3
yJPVaw3m0n+EcRtpcufCgtaxiY/dvxBr8Yg+jCgE9qXdl45X38quRVajrhNCxU4yxAUq+0MkNvhY
aEIHw3aa6ux3drYQBBZISmx1V19MWU7ARTOozMBrUYsicFDWBg1za8cW7hLMSbaQuhLbcQExChx8
2Al9o1q8tcsSWwRCRvNPJY77Up6/wSymEiRv+S4/29GnLKSa0YvxTiVCecfLS5pHWOWw05xmCPNa
WuJn7QsrSpq2rU8Gix/5a+gM2c0tZ2IrHzmHZ5Y+a8mmmF6HFpg4tP7igJUb4N7ap6EWtDNBIsfA
4fFZKwQAQ+8qEleAEZj/oKitzf6OXM6+YmgGLTGEWsic6sQmIThXUxUrH2keZPr13JQDAg7cVGof
bnMSW62PNsbvHyZpU30tBz683umPhrWByifknCMjychT6UO4mtU+tG78WoEd868ptxK7Qkc30t7l
BxGdNFoZRuXqR8l7NDmJlJORgzS5wPO6qb6i9w+2YjggFB9/29O61Dz2QyAxAfowb/IK7oeMhgY8
8NZQnf8dxS4xNdfbvfcHZi9nHAVn7zVGj04smmczWTuFaJuokQkgLq/dQqs+zCG6T1YSyu0hUMWv
KR2gSw8qcRbqwHDVomvmLsuseDTEIwZJCD57DVIu2iwNDLTNCAXtEQzEPJ9B8Wbre9yuwQ9u3zzm
4wvO3y7FLuuRjw2cnmBpKUbNFcFINCLHtDKzuZLVZenwMGsa7cWmP/wukyxev85wOnu3dMcrUz39
BoKde0HaV5DzyMCDi40f4bK3b2DdOHLMl38+BMMrdtE58ToDKAUd291Z/bTLPhgjTXf3MNlREORk
BiSydP7G8uPTv6OBim7XOTQKEh/LuNg34ZtDeDiAnLr6UUDBEHRUkcUsx0NLblmd22gx5/C+BKDs
QihA2rTpkPupEQ34fNDmX1rc+HRDFA2J/5QG9U+KAVhU8DSyxn1Aa/RHCN4DZIbMoATYWhg7Lbp9
jCE/4HLnTEgtsEGyu4go27Ams2k3BQ9gE17Bg2IOoyNLISyM+K0/7eWarSFhd4/AoKOEB2uZdG9d
/ku3KmpCCwrB9zqNSwudmIO8zkM2Uzjm9UUIV2LLwu05ZGrowE2PbI3o/slUZlxDFbEPJjSPR0Z5
hKK+reL7xXgrNp83Pn4TMrKA81+9NniXPFQ6s7jOBHzwcKMmfQtoBJxnLvmBeIvfUshaYG6RKJST
M0YUhpjdxlZgwcpD8eRD4BrAiyBrPF6Ci7KeD7YBSXfs8hLv9yakW9XDsIYQ2VzhSgixrkE7ITOX
f5HNTWAZms6dxfaO2qpi5TxOpk8tBnd9FBoQ4IFwVXdEfM2HyjMqwWCw+1ynxpDM7ZTUSSl//lXr
LHS0VcPmYkqVwzTNtbpfCTWq+BNBZcKXL+3q7E4T3mJlRLuy/DC7XPv6X61dthUqY/IEd8olkMIc
TKEBVIrJMLnX8EMr873BwffApj+Kzu/FYuxDuDCOjPstGVIrK+wEap81pWhS5Im6cxQ1uqUEnt3b
7q1Qt615T/a5niZxvmTsdZDcRX1pyu6hS35smy3lX0DwCKxVx4LbOlZMgfE5HLHJvu8+HYF9vNIa
MFS6iQX8TfDL3V+qDFrLcF6utGEqVERgELg1qKTlnoaHYuAuhkQ472cAP+GGMWLk+mT+Lr/FdRjy
sqgD2fZ2ljRjrQ67zWnTkh2FGLISGco8OvO8EfU6ZYIPaBnL3p8s7n5vm+mehokZ6pYRvXlLRhTK
DKJNaEk5bdK1EUAY3rLxk8iGIXFITAMnX0loxNi4h8Alzd54iAp+DZ4h2flNgUeSPMjpuHM9YQ8/
KufJ3KiLVft+nTuv6qQTf9PXCcOtg86OR5IYE5ln6a+o/4SHl/VD8akWLNcxsvj6aiYYe0wZba0M
bcvP2f9fVGeBodpwiGQbBHH+OoOqGvGsCSXim8LDxiDiM7Dwruh1np5LEM1qpDgBadyW0nomLU4i
EpXeIFpDuTJ5D8SaLLpf4X1ntFFEw3E4b8jqJss6eWTU2QAlJ0CVnrexUeVJT5xkgTYEDmi5D3XS
NVEVLdUgVssT5CD1y/iYxOJpcol62qwJJIuRDq5pNRjSBtlZMiUOVg/hfK/B4f6VyrqAxIyiwnZR
Dj4oSnvrRXt+n4wmVRxT+Jgd+uOxtu2hZamo1+BnRng2d2cbu87ZA/AmvcPQcjJthPCCsTVxw/eJ
Ri3yy3RnlwHcsF00FBKGoruOjFAYqwFTCUjcjnwlvH12ZV5r3fgmH6EyC43IPdzUKJKJtbBnDIsf
PULJX5GY00rl/phyj8dy+JS+a0wgwqLarO0JfpJA0TfZUJeTFE8D1RRg+HGsDOtFuvLRJeacVlBt
F8g6toGG9KSEmHjfhs2k/t7p667hA7yuHpgZQJKP6vfzby7ly5dDeBIRhJ8rF9hpfQIOH7vruyV2
bByJWkg3PmNY8jgQIbRnpGneQhoFXo3ORQAPzpcbzJVBSMLFhqP9l9fetleDPJMtdgOSiymvoUBx
bMCbFGMs/ZndnCBDOp83rYoh2fpQAVtWLJbBQQBOwKh4km0WuT3Q+5ByPA3MfT+UFJkeyo09raXj
fJXpUj8w+7stKICEsyiswAgWUbbMKvl9lR2jK9bnRhOzAo3BIPno+GZLV16V5oq9LcQzntZiuUcK
AxXDJQbDjUMxF+8BRfaT4yz7oRBvhzKOwD03AV99KGEeIuyeIXjW64b/hmTxEYBOTxJFh9+EhKyZ
F6ZsKZGVtrXGVCkNG7NxBxN56Tt12vOGgjLq32cL1uqrMhBe2vEh5SDIapvnHD82KYp5Gyz6RDbA
JPhFo6OxBwIDZEg/YvkkDZzHuarGvmv4DSYwSyfl9yv+BebrAxPU9VboBDmzAHUvI01w1xVdYcFR
mu3l4F+kFBnSFU+cA5aBo3rxN7/8rJ+n4IHQDeP5PFwXJsnYE/DFfUOcY9foLKmkZVceyNC5VSO5
6Oo90Pgws2e3NoSWHyibgPc81R6jBvlup6wOrUcG34e5Fslz1TPT4h+lSZHu8JBSnSQTr+aXK5hJ
vS7n8d5ndYXUL6ob/XERdytKsy8Q2uxb66SgJeG/OEPb80t7Xnj/UJnN8fOCwkObL8dKv/YbZwUG
JQte4JjbTQiOFw/vNZcohgeORdlj0tWB+6AEjfXyjGmxt4UX1uMHCIoNLoJPAsEYcg6ZSvyOATLY
qqhCRH1ypPNHH1UdZSy03JXt5swUwpxmzYVxtx78+INZO+skB7Ew/NZzYz6HQhXvZoiVLFeRptri
jKcmjKs9QeaQMHWixlpJk3vZmeOQaIQ8LLHTnW1HB13DV6yRNxExYKieNER1n1Qt+4ppZc6uCH3o
zJyU2ArsXfUYcuXvAmNJaRSszT+N2Ei8pN0e2/ls1/OcNKCZFQwdithpGOLeQVVlhq5xzUTFjbQu
kqkiU3U/si3zobvkUrAzgqXhtirFhWymFgHWk+CUgY70qJSgBrf6p6qE+fiU72WS31En+44p+hdt
NgGYuH3SrWsiccfPoAB+HaS66sOOSNTeFP1AaPVo6DWXwHFuh8GXCgOD2V1XcSNxNk/EmFXIdULK
SfGsx+SziWrBDNVO5W9Jo8CLInPDU0Y0sdmA0ELIOESxXGXUuKxF8f7s+mYMrgS7G8IPGdPAAvsW
ljE/5GdPQG5mX3HEW2PKbqqyttxipvIBIzwCdWVSO4a0kqrLXUbd72NKfDkO2OVNPnnBalkOBfBC
j0Ky+xDOtkhNyFFKdA8d14fr+x2R3PAeHDWkuR/wEjXK9M6aY/JCSUWwvh4OCwwb7snUKKMnpZgc
JiSGn899Af1gu0gOZLBYM50t/59m/2u6PC1K91Vd0vTun1UxBMUZnw8D6T8xEERhu2KWmnD5uYw6
o6/y/dcsKWxXY4JAKN1+yTLBVrgLGOO6+MD2z/bp+q2J5xRY+TGrbF1N/rHKZVwTsn24QINYld3e
Fsj4/8xnZ36vHKPMcRlapDd0FM5zLQD8MdeC45ZX9w62qHYYlpKI7z3KdbfqkZEePaMlX8i2AH6+
xjnoIclVM0E5V1yN/OG2c33xZRDKJjtCIjkyjdLG0cLSYi6cvidkW5a9uztaQcYDyriv2BWVBti0
+5y8mBeL9ladq4iXthG4vIDuqqRN8Zu3jJc8DTYcFYwbFtp3V3MtnItAy/yyuW+JK0LFZ/xPt390
iDvowTFEV1yLMei/Nowpzbk7Xih2IbabAxhXAW40QRJRZYeZUJXanFh/fg/cqtSXTNV/MGzBm0fM
BQdR1VxWWzBuQg82YdpfYGJZj+Cu+buHWA5+bV95UkmK/DUc6iKgAMVWNZNA927jrA3hiXJ9Erx8
EH/4o4pWfavtZvvcOWuG/qrEs6KUo5vm37TQrccfzVvDCbxSYvX09fXpbNaHridQjphxSg03uEZb
nyLBuCuB7rj8tUXX9m285f9yeeIyYpXkT4qbVmupS8D4NyRpoOrIVQzCeuW6EQSYUqNYNo0iU/ky
Xx9qBqNQHeiy/aRE02uMZfDu1QtqnR6M8Nfb4ogKPHyFr16gb/kMRISKb2sysD/FizdfPqHgCZ1s
Ns6TVUGry8cRfoJarJXreNjoXW+l/iPVcAaZa6w5gxNOuUu3BnlQ/JFuVh2eohMm0PmhvT8A4Ap6
dlXgJ6d1FfS3/irxZXWTxjscYtNk5ZJysodtF9C+EylHbCTZJn8twFxzIzc8FZPP82L5qI/qJMe+
kqjt2ltjDp0ofrV3qxgYudzFGbZOOf8VtsOsunxtUd+KyrudhrAk5hVSE9IFVdpSA3NYNenSz7cL
GFG6mgzoUU1lR0N6SgKcXje2wCjcrCD2Io5md7MyQ6R2dnQjHDJwWsEys78DyDZwmGh2BscXzVKd
qDmGhsnjKcIctFbtUatGUCSxg99vSadno3zW/qOvJHHPPd97hxddRJGCKum7lWty3DvG0BqZFqi1
4xXU3RZ4HFtbd28dEAMbk3vZN3n+PJERerHzX6jSAMEuLjjIsEx9xLio9KR1NsJCbjNI/ovhBpsm
eOS9mk0savVFP0nKKWuiPnI1n9as7obrkuEYge5VLuhkzQF4gj6HyXsMLr2/9qK6TpRPYrAWtL27
K1/Zg/2X3ylKQUKwkP9B7audWYDEVJn7sqgkHDJBQ0WOJuNtNOrZBFokd6+XjlP02NEz061yjpwa
+4m1/sDqbqcUEExHULjDcKRwwZFfEMadTjoQ0I68bwKSruT4GrBadbg8rIymi9oyZcWI8/vNByud
teISp3EU8q0wNleydM8slaAUQp7w4MD2eSI79AcK2vMT1UKDihdWxbuiKCgcps/UWpPBO63QS+/P
ZE2rapMtCK03c3r/jJXG/FX1HUW6nk+nPfsCqguO8IGGCGs0VSO/4dyJ3EeT+bE7bCYHYX5xR1Ze
GKNH20S8oyUBCopZLUqu/d5RjMzOS8fAoGtlxE4IIaiNGjZtDz41ZBhAMkmXglSlR2ktayMLi2gt
hqOcJwXVrR/bKsC5IxFLwMXx9LBSClS6uxF08QCvucagA+wYABYBDvDGPgAbg9jdqhDvwj2zkESb
GkQgQPrBpJGqLHS6cckLWW2H6PLM53T9uUUVcJuW7FUAos/eGffpjK7F6iiNMlZXE305B24as0GB
NifpRsxYeN3jj2yq73okJQVpYKqQE+sym+bABTf/MTClD6yYlaadfEKGHEi39Z2Vn8U6/HWjtez5
l3uWZpPiSO5R4IlrFuF73TKhZ6pxK2XzD0E/OJkakVoTJ2MOaYSPJbdnfBy8utNtPqw28Q7h1d5B
p6GahmuK8GPP/kdSe8AwXAWuSLG7U4FfLK/ZvX+5gcsbQnOZlQ9UD6x3DnDu62iUPxi1PtGaK9oN
pGYDM+U9bYFzEXtWEdIoF9vZqSGHjO2dVTHSVILt1fBy8emcTtYlmxMbZMomtWvGBOnufrOs7Oh6
bLbpem8MYOKaQ4lW4feecHJOWRutqDsro+jrHbgc/CKwIH93koDQTm7MPQV5Zn5Z74tcq/FLKY5k
dHihRIzF5unyin9P6BfUkZz7sIKnM0MBKOVri0xDTjjzxcMyEbcSwfJJnfas8mbuvDRXAvp83fpK
HwMCpQuTgd0LLWH9473PwaZij6a2jkEtCKwy+0jHRKy3WRgDfxJafkLMhqEM3dfaEi0PMluDd3M4
fMvj1jYd8jUGf1RUS3Odbrk6J4vw/X9wkqMRJtc5pSBrrGi4sKA5N58ZckUAa2FNFtXtkzYgMGlq
7J153OaPJkrC9iF87Hj9tr1y2Mi1F9DWhCW8YZiyyLX8rdEIbGy8OBf8roNGTlK2BymFrBzwe9Uo
R5WqlU/6+zV5gcdMpbb7x0z1M9SeDCuBdh1gwWekS/lx1GUytmtKiWlpRFiQ4Bo9Cck3akm83jjJ
7cQRdE1HcwIJjI/zHRVOuQ/VhYQEbS4/gPlO5J2il1D3hB9IkETM8CQiyUE+1XnlAoihPiwP9wSY
Ed7FGwLb7IB39sbyMnxdlDtC5R0lkFQX7/rs0QwDyHIa2ydWOHNOVCxvbZBVKEP77K9MUTRcJbWQ
Q31xh1nhQu5FC78OFCx4b7COKIaGqyjeRXmZCt2kCUrs8ADJWBNcze7B2+lTxYjbhn34RWRVGXSk
SHoIZm/gcVqlrDfb1wMj/MXeMSa3f4BMtJ35mMKDbTQeRlJmKpJqqpAHSPsXgxzM9qq26wETMYsB
u32ldLMyErPMNqkTFBW7N3OTyr2/3ZFybIMfPzXoV/juMW+zg9XWI1aG6z5psExMtAB48x6X22qI
19z5hr4XfKbUCzBeJJf5Iw10qdro8RX47pFJpjqcM9F8FBSl3XHQ8yhaEfT62xdKEPVOkOeoiNlo
aov/uAfEr9rGrMjVufMEoPVQReRn+WRCUt8i4KzHLMNJqJ8fCqUwPIILn+J2ktYx/e13tXFRCm6X
D5yrAgQ1iyawOCaJt74ZacrZsE818OiMxPc8nGc8Izb5Q9b6tgFP5Q9BsIz1XPxaW8QNKF5wWqas
gtUWwQAOSwXml0kit8MDQeWj6tjonb1YS+puIZgERcaHSPKDdMLrNxWXQWDJueilpF/Jfn9YiQ16
vFJIJT/tG1142WsH/3ENSFh9BjbATWxMMlIGiy1RyB99EVkAST/w3zaqTKdL912/gKLmJpjYN+vP
RCz5jJHy94L+r/sxhMV+TFTAM+5IM1oOxPSFwdjVruDcQb3nFOsjk0IFZFahYqVb1SZ5tp6IbDFm
52QTgzRfCel3aQqvnuYXcWQwnXHdfaC6KsLguE20Hm7bqKsOJ6abPoj8H0IQWgjwW/EXe80bIHvo
6XvWBLaVtTCxHROmYDJX5XbjcoOTjksnqBr3CKV3hpEQ7P164OxntjpvFsne5V4EqNVbpmDnVmo0
c1T0Gq85+/qyrLsszGE6sS5cDar4A04fbeyhNanc1VysvVEjsvnOcBELgfUgmMfHOlS9aZMiPDSC
naUOLqDO6KLd/lVBqWnW5pI43EHdAVTB+eY3OGlJhmSw14SZXlfgMIU3iLHY0fZ6+S3R1C4k+1RM
EGMF/rYLEE0j8wwvtIwMF15RAxZNLm/HyXAkiKFufl+MRjYfInnhlvV42eMsYdWsrc+O3lPRJ1w/
NFkh3pIAxdzvL2X+Cq1eODttQIxhg9MwlM25N9vIyJnpoF3+H2699jfa5Lfl8nMTz2WABWNifA4N
9ZTr48vZCB5ntIhJdBl/pWsAiDf7AInePRautLRih+ZOum8uT9Phc4FHUri4+FdS/HLIXAl+vlXU
r+V7UqOag4aRPQm0pEbGlBhg1Svq6vrRUYEETzwCODa9CESdGIZQERXRHBnpkB9fCNfJYd7zRCqf
Htmb8Rn6Uts+3UY2z4R76DcNtoRyCUbQI8m9hunMovCr77sgLXo/Z1xU7Dg5dZajfVUC2FOo0U+z
FpS524B9gSOEQclzxgU8vtsRo0VaxiGzz55JCXiwqvhuhOoR2WIBnmYlBep+eknyaUlVgZAUC8fo
4rdsHUlQECNWIpKrIPu8A78EqVvo/JzLrXJ0ejAfCad3p5PjrJgLquls346mHQWxTRc7HFHQVRq2
UPmGyD5JsDYSx7n6UOvEW1mnYqqjDMsanmL+0/JAeN3k33HUTik3XIeEmEhSMDcifu8CnobzWA8m
qFR1g030vvGJCwWZSrK6YWz6gTtLIkuBdxFERwtgHUa6vfuQgu261ztpx6/sW3EL1CsN6uFWOiHD
gM3p0RkJve1FQ4zLC9+PUZf+Bhx0zcYrJ8fhI1k+ArJpy/wRy/ekpurNWh1gNQtX3agLp3Wlza8e
LpgyjEZ5xRoFHFubvdC3y/UFlfqgIHIS9UiWfRqMvOkm5Px2um/ba1sN0n8hpxXY9xvAO/wBwz7f
wrodz5pqoUFMYtPiRyf3zvSFskFYh97+OikFAyTzd5XeCsoRNNtE++kP9x1KE2VtxDyG6BZ7YxLe
Dq3d5obaneqOaOSqPx8cXrp162arCWiL9i+hFpt4XICJIHy1+nHGwGvYJKez6hgs6XgL2YXQJPH4
30Bxn3/K+TM+XhHSGxnCXWpkSpJhqidEAaN6HRZgIb1dFNjkLcIgv73GkQREiz5tRM6g1M7u9LI8
JeD0HR/ZP0l9gXW9Y8j9xtgh3Cz/njvM3icy6oYqKIfZJP+8ULOhsEhQCDEZXjPNCsks35TqEH3A
+FZ/lo8qtOXcsDtC74jUkQenKQPkmjDLizNFngySahhnRZA1TJK3AHEx81Y/UR74CcF036s3dnU1
REtUffyEqGB5GDS+k+bqlIamWXccUmScS7sL9hg4zzb0hb/S3aaZCo/oSjW9syjHEjzkTJsrjDA9
5TH2213n8fFbqJ5hhmfv7iawr+0bSmuuz9kenePK8/MbHU1DeIgLdORZMsasQEcBWzIIw4Vih5j8
EPOubsnysZwKcfuJsC8ynPQdSMES1bg8NiXLGzaNdS8DDSa1fqIZqX66Xnldhng44Boi1MKNoPC/
RQ9jAfpWFkbIxIzWII10hNK61mgGe28UTlWw0E7mOqja+cPPMxAc3H3mDOz84sj4ZH4y6iAHy3Vi
s63l2kkB6Yeas/S+fxBMgOgqxZcvrbnjTH9IKVL2aw9vcgviLmAXVbv02H+CfgHowfjgoywKssQR
ERfupOQxODV++oM0ZG+K4iUdqRuiXb6QJlteNEI4aO0+JjStwxn2JO2roHSn54dlwtbTCZcZua2T
dHiGDHdbLv2QKr48yNsvcHsgsNsLK/ERHbtoP2bw9OfydTxYUEqMheWBbjftqBEJZEND/K2e+O2x
A3+bY/YJ4wyV60in9qQ8D9OIq6mHrsTFVRPFbuoulwLdxzcenKdfhBjwQNIrofeGG8+97Vhh6GJ8
OcF8RPGNjC0P/qpuZgGJt6l/0K+ZGq2X6vX5sNJpY0xQlez9PiRlD6Qfeg2IyCaDPYirYtjLt20s
yKwoyfJyYbI10hDu+BbpducF4nfUk1N5QAU62v+moqTo1HZC5BhtUY9RJzHK3/8/cWszVOH8D8hf
rI1YBGRtxMCYC8jdEc1S5B+kfvvUH18sHpbRocsFHZ14V2f/Um8v0tNovKn4EUhD/6YzjX+yrT/N
iDBQYTZmGWGbpdDWT2LsKx1jUxdpH35KTFoaBlTfhdlwIg21DA2OWTAr9JUEM2EjrclbvGQlXbOn
2fb7yksgjsMTbd3TsuaeM3Zkb8nwB89sh4vxZy28XB8VcskNkPNWEbIr7E/tHftvOwRUvD9acqF2
sFe3Q6C+X+svRrdegfjPsg5qO7YIIrM4OhdQiGQ/aQJDdOjUWmQkrQGqaK9/nuWxUiTOFCPpbFi2
4YpcSkjmzP9FdVjutHRC0FoXO9phrK39kK8faU4fzwXnYP9WHgI+blD08OpBTtmSsISWEJhTrLr6
1EukbG0eBKz4/F+ytYAZNvpi9ih2C6jcSO4PkWjQ0Pva4vU6MRKRooKK51J52DjBXloysTLhpySa
Xryin7DlPu9QKqPYMCK5wHxjED0l+Z61CM3bIOoy0vFygsTHAUNycG5FS1c2ANjOir5Kh84UdQTA
FUWjSxpZAj0pABr+LHKGsRRrQq/BQSMyaEat7zhJwXhg40r3DTzy2JcQhlkO+TmG+15YdXYi1Ays
vuJGenMZhk0jCRu0fY367lF15ioXgvxsaZvdHoGP/qDAJqAYQdU+h3/VAVOQ/zIz8qT+s4f6id5d
7xzBEYwg6lkN+81akWPeF/f3c3JBEQG+yDLBlYpei1SEVPWMwdCcjjZ3X73OnaUeKfmhSoPvYK6H
YXmygi0lKpGX0v4SinmOwn9vlOenyZVNXRt0lpYQJLfmzF+/pWJuOi8owDtRE/9DnXCNHstfqYxS
V+pxd8Y8f5gH6co+V//kt+o3jOp4rL5jfB5E+h4WCQmjjzkDIzNDVw67rj9i6lpyhk6Gdz1HRy/W
UZ+8KI1kyBFDeJLlAOaE/kci5Nz1fQjS9cmLIcoYyyCy1hj5nXEQLKtPHf3r/uG0K7nW+2YY/0et
4KAPU59xLhoV8MoZbazvZOtwj5IivBtitVQCEmU3ZquhbQX/z9/u2B4ZPKAV63BT4YuKOGfdA1fq
JxamwzBc9tCAuW4X8+0xcoCCYKqrGecMPaIug2nKkGf8SpE3O4xnsx9XoA7zrnODpW0j9J7jJDu9
1xHY1EhmyWJIxkiD4d1B9Dn1fED37CoXH7gtw572ZaO01BQlL5NANXOjb3bTD05kAKc2W3zv0Nmp
TLUwatiEEf0GEtJbxiaW0leNNxiTW21C8/Dpy+KgyAIVcErE93sAYzzgH/y3fytbTLip2amKsf85
Dkot2jthjSvqV3vQGeXNXAxYpChvph/U1q1P2es74c4PeqeoRe68RLz0Rf6MLliK8VnQ6u3FM5wS
7HBZbGyZ+rATz3nLzCAg+W8O+1n7uEXFPyHsZ2Fx/Qnwl6vr2kptyL0+9KlaSutWu6JIgFUdFjAN
O4J8wHx3vqV+VQrC7ZhtkH/lpznA4EqCdXAuO6Tv1AlCglKklfG/8sOKuE8FRPpSQEp2IeyIY5Le
F2naBTRD4uoMWHtlruPIz+/Nzv/SZivomc1xo5/aAFYPXZ/iOBq5gtCq5qwkuskskONdG8/d6nVc
R5b1dFZqYQfUThnr5kHbUV0a4kv9QDjjsNq+jZ1r8aooh6RoGHje9EmAK8WGmeJpOHIOGZHgroNa
opE5wV/UyQmLuOWf/K/azYIMpDT7DN9hJLXqtBca5ips5sAyhmBggSRrFH4axY3vuluDaytYSG/V
qyEHzuXKtVWT0ZsEyN/duBc7B4tocW/aT5u8/qT/TiPgN5f84pUJahrCiGO7eL0ryujFkutBgus7
DyQ4odwu9zLjy4QZaeaFUXTIb8TkbFNI9CwoIeJXuNqRcFQgOmCiqKj9yr1Gnt0PEIWvEfE2ppLx
lKPJt3NCet3kdzgMvymC9hNNgKRWhH7NltpbnNWf9Xwn8e3gO1cydWLaDcnWylQaCDJ9HdceDIR4
mk1lxI+as5t5CbSYX2ET4xw+6ljpqLkiFRNaY98CBQE2kSrnUpIoOegRFiWxOtWv5pFK4bjt7k1W
I3S7zEGQf1kB7gTAMpYqdXJNwbwReWP0FWkmX3Qfw5eofuxDhiFztcqjamJPv1SyWVhsijMBGSeg
GKiNUFDsu+vVpXHeUBOJDL1cK9+8eQ663yMpMmJ12rZkseW5fIVYO89nSIdFLOlGupVadjYAJtWq
yodhArSn2hP3JMnlj2DwZNClENfZTLyGZR4paf0P8DkTUitSHH5s8viCarBokyuT+2IOCn7LhHX/
3BvzzSWDi/uoCI1qf//OgrkdXUM7nZPlvRYDPgWwdXhnBOLet3u1IqQOlxlNwnMDwLXSj2RKS1Im
aPzR4mvXNQV30bb6OwZG/nKxrqA8aLhHhfPboCmjxrJIgrBoCGOc0rXfIPAfij7UcBL5njOtm/VP
epAqwE3yju8zjq0MuwsJTtcT2+6GVJe380rbXIh/hYbGiQwGR15ROawVA0h/v1Gt3rS/0UtiKcfW
EtgUu3GqfN+MXx3cV/bF+S6jXlAVgpO2ZVuJG27R30T8BODEde4caEUIVPXK3GXbZYVxbAT/pXVO
AR3jGPeueTIeQOn7nhd65zyFOTIylzGGd/FK6Qf4U0LtBf/Ij2k9FCbQs7OqUlkmR195xGxj8Lmi
UbL+vHqOYE+5aQR1sTwVq/LvqxDYkEdvN/Bldt5Vj/KaWDTfhu3Ch3VWBTj1U9qf3nOb8c7QFxsI
obWljxAr9aOxlDEb5Zz1HIzZM5xa/qCOjHqodFFdHPMscpdQZDwx5+t6tjzhnOWmC06vTnR7+4hW
TScVFLnQEnzSA9F09vUuPI6j6IjYNqkImyNTGnqwiCI7unpG4OTa9L8q5zXjpvUqtLakCCubHux7
8Dc1Ge3WhDSykDm8xyJ/yRh8Uk+Fbn2yC7azl16F4lGjlMEBazrX+8i5AnLdbiV9xO2Lx4MFxs20
XHCLA4/Fmhq1az18YwfpdAR7ufKSM895UwUHERVaAVATX2NNa4f6g++Fh6pmJvLjI7JaNR6fDKBK
JYgURHEtgrTLTfPavlVoBLeQyDaMc87jtPwD5HIaTVt8Zgu/OVPa+XXHNkqm3q1adJ96UIMddyVV
F+yKq7marfagj18DNijwNQ3p7iazpy0FUou+copclCpJBlp7AQeImCO/9KHg+NlOilXD+ZyvfOFe
3R1HWO/F7HhHD3BMgz2ufLqceywGVG8pdu+63Dj8WGmrg8Lauc2gPKTMcbZ5ifKGv9DCiZktcYLk
oIaU3E16YqCEyER3OryTD5/n/7tV8REElCKN3ZNfapr2MsKfP4hpqKfpdG+Iz7VSg//06aKRApDF
AKTfzVXs+X6Z7muQbw47BDi9wTGtUtADuWBNY/VAKAXP19CEZMfKXrf1tPijfwTKUX/FRWpMcyR8
O+Xka9Gmi7Ncy1oiNaGKmSqVS48f60th8qfw2rVqfmhsmpQ5TWR6y9lqr7MhTRgxVKdj1k0wsZgF
9vyMptC2tmhx6BymtKXV8W8fjCxJntGDWp6c+mk1JvacUro+xmUq8zFP7ayvphJohkHcdS14F63n
vMi81/xW1XdOTfxDGznsVb+HHsSmusz9ZYsqIvvbJS46A3M25PTuLVKGX7dx31taKQBOXonIse8T
WSDWBWTE+FGnreeXP8cshLyXUtuU4iCYapVzDojkhs506rxMuQX8TUV1NHBC8SUdWMPQiZ7RC4g3
1FVOPRWcoo5dUgPTdC9foXbfXhQb2J+eqwiJ6BBsQiA5zEUzBAWYPS2uV4LaFYbPFwIrDdia1mmK
1ba4mPvysLVEpntMBxUqv+OF5EyoKkQXYswpJIhkT1pqDbFr61uiHrX9TM4MNnxoaCvC+qwPW7cK
y+2QoNtk7r2sll1bejgzoR7cNXk09ioHtKRj34u2iy7EFGTaHHT6JFtQeRlHufHi7r/rww0sZIe0
yYYIUvomjU2ZP6KL82BxUTsEqg829gJe5PvmFDc9edBUzEuh7bv5SW+iAwa0/ZZdInaci8qrN9Kw
5+xbKHqrS6T/anKUqqiL9/qlZ+cGU0+oJWficNfIHTD0sXVH1Un2SwSrQD68M89rbBFC6LiJ/cTd
Xs9i11kKD6dhLFKKjDqm1IFHTSkt8sXQ+EY+ecDOi+9Rl/8PNjmetUyujZM0rrwth1Yawe3LKXRE
Wwls8f9q+mAixfgI5Clkw/mgGmrflgi5hE6TpRwEzyRZxDd/DrU0KVpiG0Ex6rIkRZ9VC4EdOa8e
KKb3NRf8Sf6zY3zBvtqmFSibnyfwxmACF1/W4yft08/7/DoUu7660gpxxZZzft5TA9G0we4PHHHP
teCtWJA/dBAtYNyQV8ydQ+pz+VckMoy1PWGEQQaSubmJVahvNNp8caa5Hmx4emlwtO1PzmZIcg2Z
buf9TMfshWPCyt/EWVq3dtFdsJ5qmEY1IFrL6c7mJNP7ZCtmZ3asmMyQw+o7TrCBdBQpxKxUMG/5
MrTXbjLv/QAcdvA2a3r3I6oviUVu87b5R8AL1kV3Ym5vAsJLyNGuhKJE75riLzmrVmQacCkoIaoZ
GvwBtq/Rv0QvP1HqZq6iYNyyYTPOM4nV8/oXqaF55XHfvcRkgqpUHm4xYBW+gqDBLRW0sfuv4W4G
WHmeRJu8MqL1XGKelBxW+NvO+Sm0UVsvRyW/nbgh+6WRxg8fpxw+PvfGwHkGBOmnt193Dfm6BXof
Bjwc8WvtO4fBlroBLf9pb/TrrXaPlAcKLnZU1wPjtSrpzfttKZIWf2HsLaizuEq45Et87TC/yg9C
aRQQbxERPo/PZKm0SeHzo0pO8WRsd643o3P0Tskr2KM+Q/XN6+wN4ejV0IliWTpDw7ROEfYUUfi0
2kc7lGKX8bbhFNd0JHdY2bJ7JPkxeb3D8o58SlaoMpKpna8yAfESz7O4DDhvT4sQbN+rcX+/CheP
O455DJw2Grt65deMenS1U8zQw8UxRry9C60AzftFKllJ71fE+1dcf2de2XUj8yohWGFQGajBMJS9
zm8DHTbSo1PLGWht7eFIdjZV0d3CshaSo0JHA0u+hceDBd46I41RFwRelNbCodnWcQkcW367d3Gn
O5aRJV43w7t1y7VOsj7kOdqBkTw3SMAYtRo6r1xXoDSEEvGfTJzd2scRpuKo76yhRFyNA1bc09ld
KjJKeN2HRgW3cVV+Dbu8+K+ZNKELWhA+ybOCttemc8HkGoiWBm9Y4k34VAC8CNc1IBEne2NnzzFk
tfRFyyKejguH7UP747UqUSIt/RqWSEzk+FpkH7WNvuGbHqD0JsAiuWk08ELn7FnbbBXA5J/ZbNXW
0n8z0EXqpC5oYtctipH2USNwGR+rpfHz4BHP+mOJpjm/tnY6xVMRFcxdKCHczJFYHytXf+qj7PDE
52iYU4GDOp4rSrlHdAt+0D0E5qITLG3qEyre/E/gbltQ3m6Q26yeK/LVoRSVtOqYj2A+nwcLK950
C8LaK3khKDSBC/AVQs4HSOetgtVKDHu1nxLKxIs165D0Pa5o7+lojTUx5GIZSGKhjJGl8H9jdy5e
J0XVeQLZXEBvQpTpSJZ56BkFyc76xJqbT73yNPpMEPLppfUV799nJRgBIEutk05rtOoV4yAA0+4O
0CcjkPodjKGXhikz6mlPKGzRkWqmui1MjSChxVPCigvnGcqzd+onezOS9mY5wpENOutJbwpTN74J
bgPVNGtX1vGNMHN6CEPzGiWW4Zu2TdZTD3Bb1I9xQPb5zFgOeO+cy+IgKmWJ+e/lvDkeudFLNQjm
KynHek3dLaKRwndypFu5TSsqdp3ZSIKo59cjfUGKIgtv7z7hs45v0UB4/wG094RChu5FFCKJ4EAc
164MI1TncDxgS9b2TUcNCXswOWZLyyg01UMUY4zByoIVPPhyNWUhaBMb/hQ9ZVLovpRz96L5MIe3
3JNFFivcUt63HxRxIDFTtNpHZ2sqZfIFsq4yxPzc7DEEKOASxpmnQts3pDujBEO+VyYMn8aLohLF
P3N3p6Yx+HkbCIzYT5yaMZQcabZ0ePJMEdSywJVXBBeb0OQFex52VcamcUO3BmlivOh7iRZdu5Nd
JwHuYj1PgHhD7Qoc8TQo/gCSv7If27ClgaxerU3SYsyCRatJftyJN68ki+6NJZZ3Bu4e2AIRbryo
VkGF+0FH9XeWVc+PlgZk19hdc0qDj6apCyKaUPfo3uHnGne4+0k+PoTqlHPnQtEw2Dpato2Mxesy
ywUYAtk4UVkC5Ohu1X5xcPYk008xQnIt28swe1B9BkdPqEWujxC50cjT2AO9RUSxkxwdV4EH6BQC
eqrofJfiSKQ9sUQ0g+k52t9LrhFbTUU+F8PU+I+/oBl8s5NuYqkazQMUExgWQBH7wbmdQ9S9awkT
3zpElvFuuetuHaq4QtBD4CjQ7jwjsuXvRm4pQVJr+L6XkT0KX8bJfJRFalDw+kP3DkDsRyqIcrfm
m+o4lhKkEcg/DWmZS07uIUCX4iXLMCzJubsddwXnd3sm3PfNyoF1Thv3dyJe9826VrViU+T5T5PZ
NyMmt14FxfXEMaH+uLaRkc8qlBc22CoeBFN7UHYaGS5JVMO2D0KY2O/Am7zHfrLM5050b4R2nbPV
uL38v1smDje8FxSiUeOvW7kfjMVlCLQKdG9494rVZ0pMOR8Vm/yJzoihnqKFC+VNtEwRfjqNkEpX
1mQIrEOGUTCF6R/0kITnM9vaHMfvqDrOh5J/+3h8QsLrW/fEegZQE7FrBmMOMdHHYzUd7+fFusfp
nSAUKE39t2ryosEk9AUn59DdsoF7v17XVwq+QzE76JPgiyeTz5VlHARgejupZOY3KszoWlR1GJV6
dcs5fHUU21TL6oh7PUG8ecMhF3Wwfr82CzdhljQROptKJcGkj2vNA3xRln2jYBfYLBnDOkfiEXPc
wSt5RfISZB/7AzWAK43LKDNOf+xNJLCPp/ZaBkuI5vuoAToxiGaLX5ZzdbYGPemnVje8EgYCpVVE
vCbvu3PaglLUhJcV3TnbXjsYIGa1zcbN8r+vBgR52XAMyMFUdDWdxBtcKf1R+vNhp3Gim6N1Y9r2
o0etdvMaKmymZtV1RsMS/GePbVRWAS9wpkbYgyW68p0LBbYZKREWlC7nsKwOZScSVCZaOjz9kUwq
w1oOShYQX2dmxwxAqP7F30tloAsHdezTamvU6HSU1OjuRHtP+DEAhUvACIy+6xvH6BDci92afXlR
VKDBiYEti88Pnq9tP+unYATDN6oUEMbxsOwlLwK3qeY+8cCnv+1XMClT3v4/mPt3wniUGLti78Tl
kpZg3WV8UEeF2bmrwScnTrI6R16l4Gi+fqnd5ycIiDf4JFXKRnUti9IxbRQoR3Ga5Rqn51m+6a7r
XOpgVIChdQhXQJoAp1PLImbfhQJGUlsg3l0PeodAQccA9EYNhuYO7Patesm1urpmjbevPHiUp4Ls
kvA3pO0oPrABkNyS5b9V+fnfu3J8AcOD3P2vkfFrTZ6gNG0o67DEnlLtSfm4G+1NrkUg+E5pnr46
YclqhKzUOtiMWqLiHj1CxbTUwZxSwPdS6plDRunh/K+G6K3KTRhhDjwogRg3vHTUPEo0vhnZCOwy
PyLkMMkO7DLcNXceDOFDbn788xFqsvPDQJecHl/gXnVNd9kamhn/dt0UagbpDEf+wFmfB64DvJrP
YbpMJEZ895KVzKdpxzYCnEInlThDFCp9wa9c1Tu5b145YhKL/Jk03qX3mEe4moyxfSxfG/gbrpvL
4yraGtkskrC/UbermBoJdvzsGwL8rfJ+q4V95J9KufrDFduyaybVaPL3OFO1DZxCLuIUKPj2SHlv
lx2d0Q/og1uvi9x4QCx1GckENS15ACjvL41zvhHav89vFQu86xbEFtlfrl/I0kYrtUPwNKvwjP9g
axAwSITMpnPkvjYlHKe5bs8UteXE9vcW32hSdmpO5UkL8U2+XH93sbCgz3BImX6q9kPQ4KwU+prp
0aYxvoqR3RVjzNHVra74oVBxMu8Nqlv6WCxjUX4odthmowXPjM/8pPfGUHyE8dA89TtGGD6iflrE
z9WFqgkeTGSRx65Y5ZsLAg4LFNm1DQRIp6+TqGhEEtyjvAHLp+P9cAzRToYfOFh6wr/C+pHdEAWN
0cmo1RLrJ1CIRM1ismzqREpEkBhUDU2ZCKuGynV0TtCekj67Si7UcSt9RzlBCjeEsBsRxx6erav9
+DNu4xjZ/lncEAJmUY4t5zFv3c+Z4J1iW9FYNfwxs68UyidZk/r5WPzhUi38hyHaV8CoQiFUlUw3
kX2JLpLBYY2VVTlIBVdO7dw2yNjzaabv39pvFnmgur0qhF6jU+aOLoo+xzL19mVRdEm+k7vLqpDS
PvF3NzS+VX96r5o5fMXCBVKm64YT9cHSoLxaLDi33W97J+cgdZkhy5qSDAMvsLZdEhRu6gV+Xzie
SeBcRRXSr1vbD9W6eZ5RYrnkNeJzM4x9lDYyaWA4NvZJjHxCfsvRH/r1b9sU8dFHXDUVMTiCvYx2
x4c4u7lcy/jfEqeGSsaDIkerd3dxQ1piYSm9tE8nijwlUK3+6m8bSDhPF9IhFCb3Kje0ElUUnQ0V
urV/5T821svbq16F1Wi0dcYHYxjoZx1QtDZCmspllcrmfvKJbqlscAYQ+h+6KWqTvaMLYFrW+dqF
ULmEm+n6yU/nK5gwgb4GbwUgExbux7/1OqVGlvHg95EzCA/GfU6AUGgK0MXuY5pTj6vdSldUhdBe
F+4Zvsq0xNOMDNStaiqL/szO0uJgO6Q9OM6X7KJDH3nazAE4lR6VmEc+zZKPUR8Xxclfo/ntKM6N
ZMN7CiT+bgWYtvCng7cNHsQbR31yjrCE79byNU7PTagQNgNfC+lPu85ePyBVhGvzRA4Gg5cLCoL5
hR2+CPWyULM7ypnYzZOT7LhDsxoANfw0X8LA5Qv4foerOkVfFK0SCuBeQ4RIpNE4WkXaqPjdKkTd
E+EyifNMxyEol4uDNYOBzQyPoLfTFjv2OjZ5c+jabMUoTYf/RidpQ/b+B2OueDoG7cvFDIm09/Av
r/ksZf5WxIVaFOq1s0a7bX9DmaQKnI0rC6Le6/rwWNocNUxREVPKJl9e7XstsDG1Q58agWotdYsy
G/uxEADuTuAGrvfgHbNnhDx1HONQdlcc9dnCgA5xADBWXp+YyR6PH9mmzLiCn8QtnyJt30dPsIUa
OUcHywDDVRRbrZtbfeSr86aP6avUvYvPMFqYUYxLXdDsleNv22ZzxouU6rkdc9syYNbHOz8GyZhB
WFK6OaCZvekiJPu/n9SOerBczruo0bsN8txtTJQhUt+NbuOvBxLv0iFdaGwyYBmq4cGMXLxXPSpa
JpNL3qa66Hj5iVxnvVq/fXhiXUkcLsAT5dwkNESV4AxoOvANPraS2LPtsXS38RAeGRBXF/ZOuMeF
zPFnpNcTNSoe5UfjwgNDTJcxgyGPbFJAXgOO1bmtiC+K3XXHzelxAb63/UIiO+riLTBMY41hns1U
g5zgojBtBFCFz3nx/rrmi/+b3R2mRc+1gs8cIg2QdxfXD0xltqVfgtGfzNBrkAhNDFGphc7k4BhY
XRnWMUTPgZ5Nw0jX4xK3/M7fJRrZ0JGZpKt1MDDpOg7AhTB4sZNgEj6NXowg1VKmpZMT58/rrw/m
NQfM46Exq58NM3W/Yds+0LsLJon3cffyX41FBwl2VkLK2xhPHAu2PsaNE2docSp+O88lK0TckdEm
KR01X9GTjPedi51+Ze8Nyq/mtYJzYcs75mCCfAzBNcBm5QDEKYSUMOC1dOlaIlFqcB6d9M6vUgge
hM5msgEQizpHD9jjaTWKAJOKPSbHqUmcGZWEVhCvhJ7Di5dw0COEwBFB+98gm4sLyJSwo09/PMQI
i0VPoYEZMhyyu2HcmvK0a50ixYRSaIHp1/pEKeLlrzHQZF5OqRHIMAszhWM47KGylb6z+wibRsjx
1HzP8GqgBt2C84gVITrEQ/BCm4BCSbGZUrb53Qgn0Eco8mY4tmmgRTzegRtu+LHuK0QhNXOENKa0
CcEmc+UD7zPpZDbQYerrh+79rdPufnyKCvdgV0px/EwafbOIR3KCSKjNa21PN03/Pu2Oqt/0C7o4
CoqxPmIqM5WcktpgBHq+D8tZ2XAQLr2kqZoGgP+Tp+uSvMxC+ak3TBaExQAzOUYqE7JGvLgKWUJE
IhBxuQA3FTzcsYL6qUZ3qfBIufvhkfA1zktHOwNKntn0cn4h90/HZB57s5WnNvu4y4aEuG+2VwHH
Cq+a70DU0bD7axzpKgBH77QsfwE3Y2vwKZh7NbsVAInisYePnnGkrgC7vvweubuFX/F4eKlPz5tz
pX9sau0SmgJ6mua9rcOkFNQ1He5+7KQzVbJPguA071Y2EZ8DLWAcOzHwGVuAK1VJQUZz4uUSrAqb
ZkdS2+Fqz7y+LaouEP4czW8gxiozWogd+IlS3O+iyFJR3zFGxp2Hc3kyEkr+Lbmx8RnDZMSUeB72
DVWnDAPk683srO22uYOsGHRwOYjhqPxW6zubkFTi1m+s47tpW2HTfbD4XPsRckC5vyRqvHKrGMeG
U5PP5p8Rkkj3aiuBE9gb6FEzmK7q55PtUsUHLwEPhy7ZJqetuWIwPGD9d69bo+Jok4m1Pd+sPhzE
wNvugNQoz3SOlSivR1Po+hBJoBEohE9G+OtFyq9mMwilAphIGqKmjQZCr4xyH31w8a/HNzNC724I
t0MQOK/wTsjHKiYiulMC3O6ZHwgXq1OFO6GjCvvwRZbSaZuV45KPWiE5+ebXEq8RJVMYlRfAc2KC
w2ePW95KWbTG9M1tsHDR5YPjUWfj2ZXQH6rxf6zUUlATVwxNoH6H+H4Kx6+pbRuPaHflnqKPhRh3
WhxE5Jpho7w05eckQDEKaySJwvupcYdp1RKOX+IR6U0CEszSPsjIQcUfVgaSv32xNOTfZFkch8Os
cIgZ8yYns47IbjAafZQCv2nYwm/Nvh+d4fO1Vg1ateg7qZ11J6dclSJ45ovP2nRfvOG/Y5cUUoxX
s+G/SLvgCZcKFfgWCEzaDjBbmHZGrTMhfjB1V2edr9Fk3PyXo84DFi27qo61+QwGWLZksmfKLMrD
tG1OIzzOYiBWEWs7bcAsL1qd8Qn7E2G2AyGMUn8Sryny6e4mnXwdMjV0b1tX0MQaGH/V2nsaruXl
tica/VA9l8aKGW1MkGJVdKA3vB8zJQClAbJvUknRVtRudva3dMO3ZrrBSlInf9eUBNECu6HT1XXP
AJKxjVRZLC7lCC/KnFmlb/NvaIzt56GS1VoUKqihrwAo3lA9uXMxPk9iy+T//ZchcxGAAD1smubs
ryCxgooVKZ1d4q+Lqf7waDlkAVGwYbFw5Guba9BRT58Ywwc6Lbbi45tICSKOHkj31ZLdRaS39bvz
cod1i/1eHaHLs1Vt2x7vNqlrFMDqC7NnBrRkzdr7ewZCqO7eTZ4dkt+GcfqH6u5a+3G9nB6DtFju
cGR2S4pj3J+iM/7UqB1NSpP22qdNW3SH+30KA+9Iink4Y74xf5mpEt9eiQ/CzR5d+9MdEEOcAZsH
lDF84Z0h2bmvPmwS0E2QBpu35raGb2q81GeO36Tbn7BUBO7HobeHRTxBN/h5ORbfocH/q5XePZ0t
Of588Aj0u4dmQ5qCIfkqWHqDuV4YdyfXO8QE6W1+qUT76bJXpCwcYiV9pZsOhIVcMU3EpfjmwaHW
Jy3Uf/XAFT21Y5zSpDZU4ZCt/ddMbbjfDpl+79lugro8rd//HyDTLHXLqHuYIuza0SqNaOJBndnm
ZJaw1nZZ6CRETVhe7EyQKVjzsy0uU5bVb1j3RtMUcwrMAaBqoz+KHu73GIZyQEQ8F/EXQRIgxDPk
5cZdeKb23JV5zwMihnFi+pBwI8/QgwQtIByrrZ+j9C5VOZSg2svnFm53l3KuKWgb0N/ArL83zcrc
+7LPwxdm6VyCAVsq3pExYsRUhHC6PZlcJ3e3hOaPzc7R/ouinSQKgFqwDMfbEr/bIUtSdQYG+ls0
DoBUvHNjLgv6TYujRzt9A40znZu/D7lr8k1fo7oZ3J3OJyo46nwf0yh/v/8MZKag11VZcO79m12N
mrRoMT/ClE1P/ILZZAnOGOlY8m2w4EeMg5L7VZUomz9TG/i9uGxdC6iH5cWQtKu6Xa35rNKwnWih
AI+Q5DMcsxr2T6ldKFLjEIz2KjNYSoCtMW9urQwx7oY675K1RwxxlnWHl1iGIga7TmNuioY5hXcF
TWzFuEC3noXGjcG5Y29CkVi4N8NLENpN8bqG8ceKU2Qib8X/BlBbch+2riJ5IHQw1xM+rcJfqsZi
f0aeOUOs5Zgz3/VDsGEiChz5e+t9zIbn0NIHgC1yMYufSFC/vLNGACL2c6u7Ao2kGpx/frCnrXIj
mBXHJp9gyGqRUXP6JCrtmoiDoC5keGXsI4DXUQU9RHQbnNm46Plqt0PUPF+64XIM1lpLcN8QglPB
Qywv6tTTmMx8qAFOdOy3ScIsSdfYB95csoX4FeIEzcTIRmIhT2AkTPGhBR7ICHPv7EDS6tLn2mau
lzOcuEZQC/8QeHBw/oMHigP9edrzVqsHR4jQhnlrJI5rn+lG12B6QsPI9FUzsrQbG6Hez7o5xnzY
iOaPQOvy3EPMpXVGhw6TG1mwIRNLkA8oG4paeW5tdmsqEbHgUdMhe1C9+ck8EFeJ4KYAo+b89YxV
RR7gIKkQ9/jJ1ScU6MnGhtcznCcRhRtd19nYwgeNr31TeKKzubEgSwzbECvUHivaEG/JWZKBZ+gs
+4xIlHS2QyARCpHHNT0voSdcTfr5dgHgQID1TOij4y3Ec7SoC4GS4hvHdn2L9dDT/V5Iv471Zq1k
H2I7x49PAB4uXpM92Tf2e1o8WbdpC03BGs3ngjq2+p84bKln49uePBdvil0fAIJCE/ZzCqCR0eEl
I820dAg7AHM8g8yWAHpCIKs0DNUb5JL89sfa85ld0e4KngoiZq+L0txVOv85NJNO2bD+kD749Dcp
ai+1zZcfUW65IQW9PwV8ibea1LHViol19kCYBnw7gBGa5f8xSMqIOrD0j2IDkzXY/SCAeYmExpeC
ypYGuax3hYlG49EOEB4kxXPbDqKeJMwNCkpPOiiAxY/D8X/x4gP1gz6kzMEM66Mhih0xIJZFMYkk
utuwJnIGlydJ8Yj1k+OKoU+QoxvyG1PDAngZ3pRJV9OGb2fvILBS+KKvFntKX+o/uW0o4SHHcCjZ
KMqDfQOu4dY/lW4GSdL/1ivaouHR+QcldnrP6V4pGEpGeYBMAKfYcLHh8pCU9WoODzrSy81+vNSh
ydIDypxp8WzwZnpv5wdXK8U0KY14H8sQDBwNHPNdFTHg48hQe7g1IpvzKg2hkEzOnAcZ1hkskv0n
0V+lz/zprrkiJ+qcJfkRLKpSFmgFPLtkxE8uTtC+/fegTuSDTtTQwcdf56jRX7L2QxD2x8mNLdYc
6Qsp8p7BbcYXsXNXej0IeygzfaZbJv1Rtwr1nAWEy+ai8CXyILD84PIn4+EK53U+u2/BeXBiKtpD
LGAw0NaKdcpZpXQt6m6EfD+3Ry++lG207FCCxgZ6zbI9qyhNWMOHaYgPL7pDuLvR6cIAJWGqJ+XL
o0drLNU6khwlcA/lRreKTI8XKSQLFdlgxwPRasr5mtH9nL5uPHcwqQBAI0A8Aj9LTumas81CR66S
I9FLumvou64Ii+2q4snwDPgYpMjazFP4RZ+sf23QI071BCK+ZLhs8zOgm792u+KZ5lNGgodU904/
P9ysGDAqwFvF3Hs93URqLYB73GXVD9MdYm/ryAa71qCC66kT73CLVzDmF2bWZpryk7BI65BM0TLS
14OcDGupPZNnRLrLlgCCuHUWxJBRPi5iPOCDto5ZLtq1ckOQwK2RImMw3YjF5iTYf0mZ322Q94T1
mwaHgmAJZVSAKz2GLx5BX/zGPmhFQfQYbSpJkPbK46elF4eouasivZkqyfNpcW9jR3vne/3wUtqy
/+1RJkvUVso3K/v9LwUYSxiFttV6zbl+hQ2dw45xUNbuXIopUNAhECFFKpqIzGi0vhg3WcI4G+0L
+VI7MG04TfMAsj0KYXcIHenLl+U1iDuAAjRzl+ZVSxzroCktsUAGyfU5lQbyjpeSM7LnjFSgfo6B
hUumb4eEzdB71otx8Fasz+H+ZW8HqulrRXwyVGxBwjTbfzop2GjjI8Gc/Q/3PTnAo26IdC6etNFc
+NggL9Zsgz3/xI7qiF1aKDdxl2eT3NRoOHBoEBx7tm+WLLZ8TFcuHVeXuRUnNrlVdYNMZqbcIehv
fhiCc9asHVxxkcpkiUHTYpkhgPqvAaNjf2V0d+SLksW+0hPQt24rY50Pgj+S0eN8pICnvGKJHLoA
DYghWd4YZcJVz9TvSt9ukgepRSnF17tC5U1o5F6rZXiHp5sJjrTGA5hnsrerMgoPNHkXuA/yugEt
5OOJXfSf77hdrIlwwz+BJYOqkOQW/PPqB+neNnLlHpo+dTJkoHlvN7CqwxpMbsIPQOxI0U1KgNUw
6gCkgTpwbNdtMKjHK40dyd1Hg92QZM6B5gw8GkP21a47DNZSZ5br8zfCSM3+9o2pMqR4wDfgRI4l
GfhRsthjZde+eKHl/FlF1V63d4NxCcy9hiKkMb22OgowyYH0DbbT9XdsteRn1cHTGG1TS5gQHfOR
D3sifie4FYMiQyd07jNCTDp05UKIWzqbAvQT5T7DBCe4k25bxAsidR842vmZpkKmVAiTEFMOPQ7n
wD0ZacNd7FP8Fc8B9iz+nYsgB8tUGAnvQ+cO/nXwuQCLN3AiQyxDZRAlKsLcROXRY0bp+pbygCOI
/K6YkDFn7aBt5ZSVDEqG2Xl7oxRCCNNB8vo4XNTLeQ8csMo0vy9KDeoHDEjidTuTxdV7le/F5uTP
9A9IrbpKAwYbi4eOtrezg+7GGzf5SIInf3f85hhKJGhMf2sVcwQojHesBgD5INz8DQIWi4L9F6Aw
oZszPndSJPWaRCsgcsrBswAARfixUjX4EZTpA4G6tgWGJ9ZHVQP+XlL3Z7fTBHjg0yGDMDSnHcFN
cvxq6TmUByYDpTN9IvhB/Ul5Y8CoshdF5iuzZW9ZAxDsMYACkeBZOTYbzGTdgqelRJb8TP/hSI1/
LcQtCnKBc6f7PMUf3hjDKiDhn2y3AUCxHqm2zvz1UzGEI1MaqZ7ewpAWHv+9+fn+2SeRz9GGiAGv
led0zE43RxRNhjnYFeFb8AtxSidOjlYXphdZB6bp0IZspVxXIhx7GQlBX/6sqTyTA0thF/zj6uSm
MCpDruMqOZmzif7Y6mDG7Ob0zvOgYtq0LW77KvQ58Wj5W02iGjq0LfmVdpcqJp8ELEA4rg9ux9Zx
udD924ubNLyUiwlTJOn4EzFMKLa50qxPbeTPMJ2fPNfJjnhGTemsnIULbjCaMdFUSiW/7861aaWr
pr/CHgplN/wLJQ6+jYiaIpQLcHPp0NdMGFrZ9PHO+VoJ58z1/2SX6xi6VISZKQ4N4rkIVDuwT1ZD
eRNLXJqpZpRpEnWIAU3dEf53WIAhxGsnHIAQL8w0Hx4okh+EiY14Cihty4BJj73TsiU+qhCJjNqn
0KHgXA+YUf9717fmOu7w1FSBhZz9whN5hlm/q5RQO+1GZcvsbB3hZtO2Qi9PL4GqdnEEdQpA5FEY
0r03naXGsuvmY8Z7Ut2afsp+uj7UEpNpm+f43ijtlJX41NpHMyGcuxFR2BEBh/Jas7yTUocFP8q6
l831p3fN52sK9ZG2kdnt5s6HF1hEig8T5q+3IcO/rjhrhhzAkraqN4GZbbTD1SNgziBXTU4cnK99
yXTyoE2liBi81/xjN5iG9kImz1t4nkr2iA3M0866nTyHg32bpZuuNeeTdgqatuad5+59+VcA1CTu
DTGnRTRSp2SqGQbOVJPRUUBlLChV4p3LjovD8S8z3Hfx1wsuYNh0tGN4A0qCW2ZpRuA+F3XcJL40
cdrkBXBOsrVtP3ZFQDPINpsA6x6Qf3/cYqLieumnUuxwj7VhOW2QjKuXBAs9B2oYJ/IJqq9JqJEO
aeQnibVJoTer/Jz1F2JqDYnhsD+oio6OTNICRUYIzVeoHJ2E4dowajAGmdQTSyDep55MJuhEDIIu
akAuoa6k1Y+upsL5pkXpfrb38Z35/xfOtIj6Jh0p/6coZGtm3shyZxZSkojuAyp0sHGgm9ScQWT+
sQRkAQyhFqcvvjklttTmCvx2e2C0M3bqm1OYl+PVOe6whU/e3a1NeDuaLV1ppr2t8PVM1RQ8o7Ro
AicTyNTXfLtIlqVOdWk4JFrqdZml3ygXLNqsII0Xe2SinzNIXpFxI5Jrr34oL0yI08O/eu4wZdED
E25Bi8+wVzq4NEGYFloXHCu3ONDdCNrJVuqL22BAsQr1E6KKzBhUnRTs864frjDMkMv7Jh6aFVxS
LNkBRvqU4+UhR4CLjs+P2EIoMp0QYnLXzr1iUAAMi0jjCqJ4GvnSD/xbwhqIvIb5eSJulKVsG94Q
R3JEunOP6tN4d+quxZ4vGnQAjtlelGiQUiNhNHLIkV9FoJBXb5a+GIHYRqXd+K3xFo8+UnuGNJEu
GijEQGCSB3KAZQJa6kDyAKZWUE2hM1fqh2dMTcxIqmkX5/jPWUW2p0wU+GL046GUydfQF4SGoxBg
DobU+g8GowVL+KTj+XMJorYO4LXJwHr1YUHNsdxZpvsu7ouAgpFMnUoaXRs/wNms4F1GGFmNaBtA
qHKYKbAoQLJSo4P2SzDmMfeW19U649k2OHQW6XfACToOn9JTMgXvNiq5y0QDTtYqvc/uruwo/HNm
ZGegkg5RbmZkKcb6eQPkAddbPFt4UxyT/8+G+DTWxgDO90f4Q9o+WH1ZAlCbMavczw22NejSQxFE
yzqGSY6XP5t5+zoHqqFomgUAu0EB5xCpPYGiDBmZHJwv9Nkx+ikF6sT7FcUTu5vNgfiALW9SYqfK
yvb/4cHzVVlDmBWV4Fk8pmsbHmkZiNVLDKyxmHbQxKHOUyIgBiORVdsBFj4ISFfYxpeBXyLc/7aH
qzv0vI08g4D9BCOSisoVHBvs27qUhhxOB7J3txW0Bz2+EIROI1regy7T3T5gPsIDUw9h/WomsdHv
R+N1A7pOMGkLrU+lJrw0uDamoI+3pitGiixedgHAlMmognFM0uMKpgpwgdxmR8lBLMKH1lMhkhUG
O0T2GakpGudWvRp3TenOKxoiIeNjCSAahaZ5fkOiPP0Q5rxhDlvU3SZggvwKaAjmKxWurZ1XVTv7
Q+QRg2tBSnAdinlM4t3LEcL8/oOnSasvCZdAM8yUILFJh5MJ5zfh7vdL76xr0BWBypyXBlk+jC3G
PvwwjsZ3DT1UcpR7+WVEr+30uNK75dTVcSBXtfzYmLewDUsoRP47dypTFQhuWLd6FoIYrW6nXIfM
gPsSzChMBFNz/tZWzk2uk1iAIYeKNO4UmZwFVYgTtipqpA7XfT2dYjRLoxlOJNbQys1v4hnPIBZp
wMN3h7uIVRMW4pPV/FMQxVvk/OfiXLlz74DlV3VmvCvmLGqcVOFJfVmjxRjuTiqOrD5B0kGKmc3R
WLflwwEovZKhe73whg4R6qz2uTV+PhJB094CAcE1al2QKl65Guyh5UpwRySCJVuYzAwLoGftKLVW
G85rRfizuWd+/CdNVNXjs7YsLs9DQ42TVn+TEm7hVysfQO/TGoTpY0v8DJn4bkJNL8IioElCeYw7
pv8B8tPgY25iDNRluFJR1TKxFG9huqLvc3199QJjYPQnUGso393BXjNP0p/MSl6Orhlrar5PcynX
qG320JeQrqjyyGsmjZxHxwvxF1c3EysXsepptYco5fhZPQ/P8cXfw4Gcq6BYhpRt5YWo7ncvjX2G
wesDqBjY/hWzpYyCee/NUggyuygH+0kpYolaglW2isKF1l93wGojVCF+oBAay2GHW2ONpbnGSqUq
P44HH5LsroK/BYq0/pezOwv7IEwwJBDz0OJdJwxaqEUbzk2Y5xxn5YslSMZO81UHCkRWZb82yrRC
S82Ct9zvETXcGUqPjVTP3hG4aT+LdtNiuBRaYy5LHYqBIL7bpkT9uIEZQNFqo4/IfAI0fOZjrvBm
zqDKHPz/m6vqbuAagd11XBD5Z47cyo2F/cec0WOYPQHAcUDiCZtfiNNNMkCJyqvU1V05cqgDn86i
tmG5o5aUFXStYop4hT+8OmkhUV5lwwB5vSy17QNxUhdtaPckNL5OhsgYf2gKZw0FO8+GXArBnx0e
uQCDtrJf3GXpQNRn4hZyGZWqDIzJyAChA/aaTCPUgXXxUh8bTyECkvo77BW2Z1gFvUd040Jrkzrc
H3ZPPRrSRtrb2SKP978pPFWYmHoDdW4nGZC7obmRdGGZa8qqlzC4k7VBwvBe+zPLxBGQishRf80g
JLc98h5nwZX4upYcpjArbqtDjUXMQddaBf7lVxxJn1lHd2FwaHxRt++QZCnKPLYf83dbU8d1+WSk
vFcjeS37SNVfnEjkuZyiiFnMUUwLRzLhiDgJZK5GoWpEA2Sub2aQYMESc2/KmVVSscQBa04YfUxY
PqlUfTMGJw8IXf8hs82b//gYMtZImGEZNz3j9nj85r4L5M5omq3aD6VhqpyRBR3zk6Bv/IYvKnxo
P7dheZ/0IhO6Nj2FZPxzHgRlHAlGrNmLkCShF84YMjeaYDwL/o4PAO7+0AzBOadjQX+FYyVdCFtr
ltPacq8qJidE1pYmWaolEcTPORPJ+IXg2hhb+M0t9YKbQDlWxJNkOExySQikIOONcVOSh/pwrqhX
VMoMElmJHBsxOQWCmkiChJxgFDY6bqMZlelX6m020nMQtaL25k+er5YP64QxdnC/6blpCazqWrk8
pEnfzLwmd/NGYE/w1pkOh0w948t1a5BQHWRWftThzLjHyXjCG86YPIEzYmnpU629cb2hnApJMCjS
18Eem9d/UQJSwkAJrE0VM0lp0oI78sGO/k9S7Fw6U9yohqsFmYZwWE0qEPy9UE47+Bwve609mFfa
cfLrEwVrqQKXqqkgIEKx/4+6jzEjK0D+zm7MT2WNNq8YqYCdL4X34XeegdsHxmSRPRRJzxQt9N1t
IJzTpUWeO8ER/DB/RdM5+jjt/huj2RYx+ZeLEgwt6uJn6uy1rDcAW5xsvz6G3jQIz4+RL+dBxl6j
VXKmmPFZxSeXT9XBusZE8mYWKU7FIrlvPrFkZ/IZmmJt7uPZZRStbW7bxcXMr5uNLnaYezaZrYjh
IBgmWWMHgDDD2DakFGIIvfHtCqTfuS0vYsJd0g+MFpE8DBFQaMInBFBjhoLOhLSZ8rFR2Ja6aR1D
h7tAmhEYiHg4cTF9f4icCyWuyVTMfTqBXKw6wDjBlgJ2Sb+G35KtGYTE3BV9lgDYhApgGywaEz2t
+M6NKifR0MfQQhrMxgym8Ov6jglbmRi7II9esOhwM07TvQt6ecnIRVxs4fjeXJGfsL9w4i6sstWF
IZVCXH5GPughgxtu9OeYkv6tKnbaWnFj0zGNo35uB53Rrewz5MM8g8LU2BL+Nb6WLB+a4voVzccq
QhlDno7bStMca80/EZGMB+kZG3IJfiYaxbSRdwJTiGFqxiCOzE+FfKKIikxKtxTcqMWYwj0QBTc+
uGhc7pBEsBCogmBsDGM3LR810FbAe4qwfhlucTdULaCf022HFtH/VMxkYiTtlWfZ1XUTKxKMn3Rf
WM0hvj/rWPC8i6kUkLLI5NGH2eg/G1x01Ia1FprAU1DAAanCrrJU+P2KMdRGecE61nNEgJz+9tWe
acUmcfuzbh4m0zovE7vFgPlqol55ac3G4e6zdXfK+onzia69JhVY5TGH+tzVXZNpXtctW9CvCQFF
ANSpLKNBcjplMDy6bqfCwTwM/uV9W+hMQ6F5Pvz3XfPxUPganzYGrci9qDOC2ZMx3ojWwxfN4b3A
m94UOj+Al8sFXo+CTK59GMp1ffDSaaQnPyy+ATRazoF3B2sba6dB0Gm69MpJIE0U781bKK4r0ZWo
qSyDEc2vW6GFDgM8WJ04lwQNFfv9cODHY22M99//8tP6F36ql1794tUynhIE0RNumgJOPCFHV+9U
yUVzGexcvoDiKZJBnXOxU0i1SBkUl2yBX3CevVEx7/wXFVtTiUSuj3yQitxx8PiWhduCFipP8FH9
ZXgogRU7gTJsSWptRQKZn2npL+Hj2x0LDwPbjCzmBcFPpQ7yPyfrGUDQwFgYr2WP9dobSSmyuwRu
mrTFIShCX6iUeD5goLn4/JgDX67kMOZxuOz8zlOxi4UsZBnD8OXHIKV1wVBVSmFVB/1389/am2bC
R/gGG/vZEbNnGZnC5nOvD2kPO0Mphl8NLF+daEGZUl0dGTSzY+zsVo0SBLXcO+d6/fERfYjFmgWx
bKlxyiXGmO7OlooK2udJGLy2a+kYGL3pkux3FTvKmYrdNDTngE8P5Dwizldvbu2N5KGvnVlOfE9S
/ROOtD+w8yuGMmC/J8gCGZ5vpjkPXNGgb16d4Zk0l9uc1kKh0p88Rfv3we5DtITtIdoZrY0XKKv7
s4wgMWx8HsN2RZSJvMMf7tDdoKfyPwBy1i0U1ee8z5DuMjEMXOkZ8cOLybM0eyKcC0aG7UFPsarx
y5qwPHChguC62ow15gQZ+NQ2VYBV6cnNCBtauGGk8XFbzHRrjknNjJxN7zjzz/3Z9KNEiPtLWHdz
a8T0jBjoXtcvZoHjoavPGgTnI5WNe3RWBF16VOKha4mQ9r/4qGljNpf5nypdB19Q8hQBAWmN6ABu
sJkIasDxpMfORxUddP6pmAqs0mL9ApiVW8TO/tQymOy7VkQ6cxm/VTR2V8XjrCZeG/fTQMvdFSyn
164cStvFXeYC7OiIOV5Vz3zHvFp5F6b/ikRXIj/dFUj6hSMw/qD083zyA4hcGKURsJybFZFRCXai
sMLLLMqLhtloZpjmoTMmBHWpg685i610jiZo9HcsFoLSCkX6E85v+4NeXXUpdUo/O29v3P0lv0pP
mHbHvfD9cpDZryf8lPslr1iNFUM9Vi+ElS3+5wJrrocAMy0qRSPUWxU67W2jn4tirib9a7cK+AVo
v2Q5CEm05pbi31xUaWLjVIdT9ZS0ZXdQZgVrsSM/sYcT5MM16wGR1yplmrgpom6GMp9mUu1cBPNX
Dp0MlhZ5ubnTpvv1U/QaiHVgpwIGiF5BkgzttVMeszHrKQ0b9j4G6OOKqTciNP+Faz9rXMVXRjE1
onKPIMuGt0SyI8GDxDle5NvgLMxL3nzuU42n31ZGOYeGVoT9qlpXg3tQtIKu26tw76Ut8moRyULW
MGxMGXzjtJ0CAQamgslPI1fGSm3bTQfPjhPHeebPIPTJiLVMg+JKcfboyHBKRqqCfDQvOLknJHZr
fTDzkGp5a/KUZT1F+bzjNURtOf55Qz3hBLltr3g/43ovszi0Imv9Rca63a+XSkQf8WYNViWuvxOh
HpmMLFZpZC92JECBHuHWA3MzqLTrlVZMiHyuVmp1dOINOhTefguHua2AAmhWVz8FmxJVfJFhjxHO
jMKx/ofOHFH6IHYcGv1P5lt1/qDLmIMo9yXk4dsfCMxVWT0wAnjheWMrSxNctbvZ4aeB0VstPkwX
FoyQ3FHj4RAnWHQjCxtJ1qfaSeTmwLY02Eu7SIAe8aNEyiKZoKlhEQNqewRMxG34Cr5aMxdZmFtO
zSXJ+e2bqCu11Jc8sZ/tuVIbVYU6wjnT32x3zG8TXInbrR1sKZn/8J6gt4Xk6W1b2puchi+sgGxi
ClQyaLw/HkMzJnUKSkzCStdwzCNUA97SmAPSSPn/hwsmaJKnLxuwX3OivlDYjsp3CQomgwvs1jOG
WpjmrGjknzskh613Km5UZBbbEXVCuB3noH7+IHvDCTjstBuzksrBpSBk3ebxF2M8r4wzBPDkZ/Do
8lSPBorusqJezIq9YysVN9CVLFS1+3Wm8/hBOUxbVbI+6R/WhDttoDa4Pnm+oE2kA9ckuVSP6Cl0
qV6CE0saUI/iS3rlXIaf2uPavAHltmiHIuUdRESdha0Zp5P8OZNGLe/4IYR5PMqeYkzmT7LSq73S
sCyabxsYY4tSBPMPAVzsFsbakmcpB7fzMTc443reeMwaZsJywU60mTPG97WFNmApCI2+RG5/PoEw
5tlLcffgFePPMQyEsTSomn/HipdBij6iEWnVoyGRBuFcwN+TA1n0KaIjD5wvJqPgu1P+b88lYd+B
pXz9P/PIea2I5cdDrzlhKkWjbpUeluJ/L/Tr1yWSTjTRq3GwNfcwutKl/02TNYj4UxgClJR/gV+L
U426phx0JYwbAZMMVyq0tCy7WKfGB2p9Zm4kmlkSZxKz/vzkj8vlAPKum6AKTk9CfEsD5Zt/w9bl
zJErmViI82GGIAVexAy0K13DiRRIm91O9eWv/LX5d5MU9sz6wvWUyQL9TqQZI6P6RvzfmNuolwGA
QmUsyGq5P7ivRWEUHVpr67uWjq/1r+gMEVCyLQH5u2Jp9MMP+8xnDxPeVUevbqbn8GqVS14NvgR8
FskUzY38GIzyLGlAGR00/oQ7IZq50AEnAafEuIBrWmrEDazma97FvFzc62qshdNYqwlf+1/j+cJ6
rP1RHrMuyP6siBcPNspg/4fOfzl7iP5FmnG9aQrEzGHXOgY3gvikfqVyIbnmjnuQdy5HYT/JjCKl
hYX6H+Nn+GSuCRF0YH39U9g2AJUEUmlO74deYQ/aENiGQ1DUS6U+pqTi+3NyrtW9teR8/hTxv8Ig
+ZF2T8E6hJIrES8/rmGn/ZOJd03aUsEKk0ISi3qAgQNdtKl4uNK/0iKHihCj2pfPIZbUsCN/9jaE
F985o+Vjxm0wvkpnkr+q3xTomPWVyAfT/p/CvmQaGB2y41jPj+eUnNLtl29LS37J6HayXTDNBFxR
+EOR10zwBJ2HbjExPI7XXVivAEh7VA4TOAMbgkjH9TQpDgLZqIeecB+KCgpARgJ+MqlKG8W7Op49
FI0HHUh26+bflqF4cAk37gHMB74SqkrOPmetclO/kvZSHeraK9Zwd8pdqaUxEg5JJwI6bCAtXbvn
Ker+grGlVuwe/UZ0r+RbLkdp8Rz3y1RyCIHx4R4tnJvPrFLhShOP2y+4YBYmZhRzL/1uIIiSn6JL
ApLRosojDlp1pioSqEdB3prI0fjJXRK2GkommStafTOLF9ZRisb+xHUpQzYnfiPSHondhQnJCLRo
m/qh0Px40p6GaJ5rJvSHGrKHePLDWxkMklNkPY+/PzoheywYHYZ8JyYjI1Heo5r+5j8bmMYWYeRl
mPxqHjHxGwrq1MwyMogAwuZJjoub/1PzNHcBJNi7HsLva5DqykzsDYeQWx7fO9QRRXs4mweLZFhL
HEPYjWAbg9YS/HXCzfT6tAGLe3hlG7eM5LODtapEVLVWajd9Ubpun+xSFs7Twzxu3jTPitFqOYMd
L5KddZck4qq21+5oOOFqxm30ME74Atg5GLzIG6nilKnKJPADGpGrlzT2g1LQzT8xCx6CqqzQL0lL
M2Dx4LdaOLOPCSnZ5TuAA5mMtRoNPd2aEijJp7uVxL9WDKFuqfxBgvVC247+9lN/2zTUSq2/mN+u
XtyRNTXZSfnNvRDv89LKRlPm2JlszEtuYra7dRumVjA5jO5QuJkE34yGAZBvQrTELlmBpQb1Fyhi
f02nHi/eHR/n8DEXT3NFMX6Jf3FunSmhSk1kXoSMbnQ1qBCP9dj7llpp/8csBFeaquQcje0tI7lo
SVyI6y49AZ0gp+CkXipMiJ9k80Fs+vNfE4HQUpN7JFy5RVUidjCQbrmf21KQo2hlstJlF8ID8AGx
rubs1W5mpmOSyVCSyNJqvjlqHrdvivuvuTXRrl7YKnQbL0onYe+yMToYcPTi1Va1W3AqWDhz5wZd
VcIvlPyopzCUh+11/wI58QJGJHCFipJY2SJVViqLmzfAXDD396boCZg3ZmlQwNOeoIrzULICy92k
aavOCzjv6CBzNg+0B2VM1KDxsE0zEuUcB0Y1RLn1qp3P34FceagWU6X+9+UYtoPYNw4IIJsuCuNH
UfxGoVevP0NWj7RRragBXUkpi5ghtcKkqU03VFSqA6Wjx6Z9GI1SasWG9Y/uLp0GZ99ChjKqKpdB
tUoDiVVniouWGA7AurcakfZCSdgY8RoFMfVmYMVaf/Kcna5dPIn61oMTR93b45Ql8CEPYbREgBe8
IFoxoFFvPRdpl128rjW0Mp8c9RjqcGBiJM5vRoivMObxSe0TuoSsIvFb5QFzDLKyC+5i8wAHVODh
+onmuraxKXULrCMIzlIFxlWSYArNofEsnrMTxqKpgKOJlAA5obepMM1r8pl5NXGEPUgfG6wqXadF
6BO1/gjhGXDQ7rZJ+Pe7PcHLCx378AT4z6hDI4OAMRtm7DLGc0CJz5dPPlvYUYtQyitMj+mw7iBa
DGmBWVhgXS2kyIFRkUByCSaLmcu3tJW8fBL+H4aERcVhJmff+Rc9/jBy5CvKuhYJgJKQHv1iu6i4
5X+3P18XEI+irEHV5Fg0/wlLn4Zxbrgy7hv7exGBveaQocVJUaCddg9YyxoCw4TtX7Qi6fTA43yf
THmLVBuE63Iz15BpikawBdTYpqUnXMKTjC/WWfmERhL6AD5TYq4KxqHdjHSlRhZAEqzQ6sODsTTP
kU3irS8rA88dpTIDHCLR3uShuf3GUI05gcYuArR2jz2C3s9+1WWBuTi946ElBFJmeXNUW0qSkFNw
BdwcvrmyxBk0TY/0Y3Oud2f/K4cqyxGG8mNoJF8t7vtOrE7dgygGfiHmxcl6iAj+sZXhAvrsu91J
fuLPZtpZen5tenKMhr6JrAj6X/iQ0DS+EWrVgj5oOcd1bT/hFttKzr9W04PPKoGRXnfCA5KxJ/oe
A8IW/8XXjUPwnPdYrxbiec54V9Rko1CmXoRG83+uMjxuWzsY7j5zVvWcaU7Eq9MV9dOJzEtlDHwe
IKEAxG4bXVM9JsNCONlDj2QgQKmEB0LQGCw1KAY6BvSP8TU/Ze+bQW6UZ7K/9XQ/IdJzXNA9h58R
40ru7KDXn0URAC7n9PMWd/9XL1V2jyyyEPU3J4khKn7O8YTwF+SfgdE4Xvik09xiKxczyL9bsiTW
ZDaqjxw+wasAxRTVk0G7AB/ZOIq+WIkd0Npi/wCMhVI+zOJ4AGPRnQJT5Nqxdc+FfACUs7HvqckB
/j7i6bc9sbjvShwjNDJQZ09SI66YUtVoxmHFtDOlm4UsmevHpS8ia7SEEQl/VM6LlTD7cDhzjImd
RT5YtR/xIknMSz9zjK8OIUEQIsSlPOv3QtDKkh3Yfk4gaR822OHyCo5oYvd0DE+8UGb4dc/N8oLn
lt+BiIpReEy58OCRkDGL+J0pdHiUEEFndtitMGy5SgSZAxBkPx726f42HnBdvX3m2HOyRRX/nZ09
ZxiG9LLds2ZhaH/5Qwe82VK+IstfE1P3frADgGVikrKCkNSl+b0VhS1s09aCdE7y/zMV/pCD50Es
gHcntZYFBCLJp7RKyOtF+wiUmn3n75lVpW7qs6zXuLPm9sk4zE1IiQSa3sL0Pt1l0LRfClfEsrEm
yscDGiAd2ZYbW77dtpejre8DabTpzyboZv7DuF0m47M65Oing3vq9z5RU9TVJvpkUfJfzIfYzW+N
EAv8wgXE4VCXHK2dzo32MRlt1FdPkrmawf40zbNMvWs2WGHjMuTUFEd1RP9MK+u7Oyj1+u2hPtyn
4pyR7ShxR40xcuCJIwEUjAqKgTyEhiJAwvCEvgKX5AzPtru43tZJdMXahTWZRy/sDN7kjlzK8AZ+
mwFwekAJVm3dOVRQC3JICObzxPtNMVwl9TdNPpQK7/WXnBaQCs3dMPnhBrF1nv1zt8KzN/OL2QHv
6f+rH/tEzkEWx+HCHWlyulHA407wXX9GAE2WDqDZI2oxf51A85Lfh9PCTnoyPqQpDg2EQoC6NB4n
bQ8Z4jmqcaVqAd2LEq/iWjxumooYqrKiFuLDYsEpTQtXZGHbZN3af+Cf5KxhIhjETdL6R0+YNAb7
gIS7pzZVTyPh5C4FV4VWfVwXsDOL/8mFtqNIQH7mHCrYiee2FULLnvpC8FKxlUlCxHLjC9VgYCw9
uF5yqvw6ra5cKK0TkT6KEWlzt6rc9XKcM61jOz3PJ1NLpACAndm+5Fcz4pHg2FmHMmvHiPdMM2Q7
LSQrLISVNQlEseUXl+PJuli/MKN/v+Cf5irXnDsaTvDvknFbm22NT0eR3i8sJf0jk3cGpDilgiPF
Hyjbdh8Qd6pEbkSthyU0rZ9E2BVqcftwTTxII4fPfeAkPcftuJWzFiNsbuThsULiPxTUu22LWVZk
9V9WS3teH5ieX+jzn2ov5NAz5vaBSVP5EbHzalf2Y2k4f08hTJlOldNLC58jKrqdJ9rxy7yDsn5z
ZDFgZ2ySPEEx8PJT/pdQql2afqz3Zr9QaGNHynPGB8htfFzF7YiKZKQlehTu+Po2TLCZm/THPjsJ
uWD0+mmRBatHfSoVenpAPhLvkX+AfYjOvtiRYh/Rupb5Eawyy6XQy1H6BSJQRKy0PygE3RHYKnae
HaeYhsaQFQqaEaDI1MNstdxYWI/okuI+DauJlGibjpFrs7g4ScJEWK65VdlbRlDhxa/zcBn1Br+/
fZJJAJIoDnkwf1mTpLhuwMRr+jG0cIYgIkORFuWFCY7w4NdVDYEipCLl0s/KKghB3MojRX0amMFq
0KmN+SS2nAO1izKu/85BPf6ZUc7qykZMIxaXMVjiL8mpctz8eGJa0yzmiGwO0bbes/xX3bV5ybrx
I2ZCsOHxOABBXWMAjc6h22/fpbeYl972wG8AYjVFb2HJWKdHHFGghbh8UcENUAn7+llhazoXzG1F
BZbDBH7LwGzr8Cg4iN8MnhayyT+p4WmA3vDKkZ5kqVV/O3eelL05nBV5ZZ5IxlnKiFXZXURsxCZO
NJMZ3V0tehY3dpYm6SktLLyFBNGhwZjpj/iGCoXlHDRVwXN4kEHDSdabUvAnv4MYwhWhH36xDtAs
wVBrBgrtCyDT9gC0Nv/5PbvYrWLzD7lQLX26bdtY9k19TtNBhDY/6sGD6PeZpCVAgSozV5pLUlmF
CM079vXgLzaLs6uc1X/QkRzhtzuBLYs/FXc3pi/QDxry0Dco72wTcMiT5v96Bf4Tl8ehQBwImmzK
DWq/DHJuo2Ad1r4UljsGKyDWVERUGG0DyUEXHzsRKZgIqdnfkCLeu49lyqsMSirCT89lrtd8wone
nMrjPnSdBT3W7kVJBXPGu4Kz/5V0sZCQyIIYak8U1guDP+1pwktUHhnzbf0GoaFjeSGE0jbTWhV4
EQ2c3Ee+Fmah5D2YJn0kvzyIVXiPMwgUOEUwREhB28/Hh6EJuYHCsNHqRv+fiZZKRbuY7ULUzTKw
QK8aBDIwBX5EBezZCjKpUnx+YxXQlPZpzLEfe1H6x3AsnWHoQAThiEfbaeNaGCQiSWIrh4cuIuOP
iFOitfHnwvl0yHRT95ZCGCOCTxTS8j+xDrdAsTgsaRo3pZ8QO2azM7oh9urh3NwubT98s9B2ulm6
VQ8syBA2DtME2eBbpuncurMFQmqqwPKkBeKcl39gBvXVU7kKSV/eZk3aAOuMOhfJm7v4Ws1jh9Wh
GYund89KMrtTiLQXpMAt3B9X/wWpSP/JzQbZyTXbBlxdr6S2WY0whId1rfZQWXyg7hmxksgIrF4q
ehVAXT463RPVZGe3SlIMe90unYgHfspnbKcrQZKmg2q5hEua3O2dAU81HWxqkYrLB3AVmwwsyhyg
++NJhlE9GS0lSCH7bQMTI3/e7CYVz9sGzbfJyayGOP3t6zx9QI9TE+rP4s2VWolTQFjikLixYr0e
x2xKEbAAw6a8MSdpUgAXlcDRJzwXpYV5pT28x/aDUCtJLOLlkqeX1LU3D5Wre8Dm4Ury2XJbqx19
XGa2R7UwyXqTDtrF2RY3RGG4Wz69bL7ZCmiEwu9gPhwhAaQnND1qb1P9FDzVKEgwLVJccAr5qdI9
G17GqyFOWeOtCvV08VXJXiqpK/TlnFz8ias/IgRz0IzbGJqkGCTV1Bh+yOW9tu7iY+HhKQ5LC8VK
vJx4F+ZzWhLJXVjeML9hB1jvSkvo8aJ/49U0qfi22QmK8IhZScpLRN45Ou+rlZhisIuB9Gt8b2ap
i/hqO9vFtSM8BzYjxDAiA264U3rBEjdhDbqA5Bv62v62ndo/4cjfQmXRsDk1s1uW2t/TC5rlZWD3
OeQbSMT1SzGokv5YV8XBn7krs/ukmgpMCiQRzt4w7GbGjDkdPlIftCclAyB4/7FLnqetaHz1vQcb
V9EZzfaCh1KdsXceXYH3WFAmRripUx4PD0PBjuLJ9J2ycGsexpgG9qdktpLSnZF8dw9twMBrqMrF
kG2MVtnamxYemsUq5yhqY819jHp25EI5y0ufOInbIvwR6xheEnA4tLyFp0bMhgfw5v/QGjnwJwi4
ebopOdkxaTb2rpgbjikFpJkTb+e7VKebF74w193YZ/c7lqZocpFi2a3mOrxtynCLvjmG1Hwd7tfv
pavrAmAcSA/gg/f7cZBLWpqm8Be00FG9Bv3SD9ysJfo6rN9mIkZ95rPTmxDCD6xO9OzVX9Vex2te
fnC4WSHDRBrLkLrAxq1rn4sDwijEJ4DUMM4PT0gEZF2h1W3UpN756qtsmFaX+7EkikzTLhaMvVjj
MXXPltLuheLR07jpzwRW4/dX4KwnbgpsAVIaNazZGuTggXjIWTnlY+7E4kkUI4ouJ4X24pQS6isf
JUGRt12JdhO4uVvUUKUK1C/vYCkvS6En/iddExyrdWV2geb7AmP14rz1mq/7r7KJKs0Ofoa9SF9r
gm71bLvmP9b0X8n8C0W6aGi1lMV0v37tuI/W6XFy7oo0yjA+UCThULOnTomA7KKgHWrrzNOOERNm
Je48apZACrYdZm7PgG+VaAE1Lv8PiVNj4g/65mG/7wdBwnjGIEneV0JhHjNQBDBH6MIy6nPGWTpt
EfIyU+eHwLZO4a2AO7Jh6xSM33gDtGYMMTWKQJ3GPYuqO1Sd/dCYiCb7x+2fj+5QBmCzpnhZ2y87
3r+vhyO17g9etpwwxUr2NjPDld/0+enhVOlkaGsSkHrtHqJUjZ697t8SRvpxyWY+fW/AHdWoeY9/
2g4itPUOBf83kyjNMyRYjuOI1cTr5bBqefIUlPJqXL5fuByh9h0Du9wH0QLIutRmiEzs12jGBoYb
Dojzd5vmdeZfTvF5dsaBJpWiTBNSa9iTNPsc0a1DLL5fAzLlZNlRdcLWYi7P4gkGB1NyEuiMbb8T
0FQfNs3FE0fxb/kOV5x0rOMEI2RRBbkYz6Ic1kmCFByKC5wYBDe8p6g6Nx275SITq7AHRg4vQILH
sid6n2w8jD4Kob12v3KsWad7uTF7xz3JFTq7EOAOolQl/Hg2yOyrIUmvij2KXpjM0qP3XAM4WJs6
WJs9XFJiJNKRlhjCjSt46HXG1NC2z+rNTjfdw568UkVGKORXXFXcwMyb8KkOuZ+Yw+nv1LWR0MOx
wkzN1IzStw8FC+EuemfKx7F4nzE5n8+mz0GMLsmGfO/SQIH72VL4Jo6P8pkKZ65jsR1LMlWN8Uwg
IB/+DHdxogLdRVo99GrA70NZffpDKhrfaQxE0Ng2F0Coy/YWHu4MdhqVJvQowvl5L+zq2MyIR9bg
qAyC6U/a4neeNfpHn5Dir/Y0IwXkHkR8ppZkMnZgZsZBQKc2oZ9Q+/9DWAJHTOJYozBykIACYQTf
XQdMHgjFgG/phBuGB3o2+OCgSTC00dRX5DMNakAqFw46liCm44enN+rxH5NwzCX3GVzc4sBSQs4E
pFLfat56692r9QtsAANpUnw0oIdFRRVesOOiSy7SNvOfbZhdgIC7dZIEKHXtwv4U6VPd4dkz+FL9
/A0XnVNFzztBAbMu//g0TUjWT2HZ5doUpI1IgujbVXn+OIEHs4D8sRE5q6WpVibrF8i85uiEN3Ep
y7c95iGsc+ihKy0wUp7Fo+h+heQ+9czkIw/e52zYbTmIPTQec7sElKx5lRlyf/LNvr1iDuRbRSFo
734Pk+OvePCFGiOHdEX9Ghn6MS/ifwhIAT7uGqc4RfITepzZ59ob1Vk0IdUIa26/EcVczTth8/8M
W17GhT64zvHKx/k7c5cjnCl3lrjr7Jt3zZyXwCf+fSNpoM0O1xFCHs5Wk3C7uJYn9VsF4FWz31uh
dmdrke2bpR4usJmux9IhAusmVxyfK2KJ03msUgFz9LzyARZ78o/kMxbkIhebiTbNGM3/urDVYa83
przIP/ArukhQzIe4F0IEZLp2TOjCSIZczqwKycWxoR/XjwLmE4ar6mMRCK1/VeL2Qhsjm1sxVzd3
9h4zxFbCR/oHUsYT32Ol7ceC/AsRy2Y90W5hJkkjrKCNTbdWL2myDgLenJB0A1VL3hTsVCgzqc2/
ImQrE24J7Kwv4gURxfjNzIG6I9EXJIfXsk7cmm1yYmR0CqnCm8/dDlt14ywZpUFVKLN0I4OifECU
Yn7ILe1QGVQkBW2wKmNU/nF8VFud/mlaFI//Q0hSgAT7sW8IktxHelzHi8/aOJBZWu1QLTbnxwfp
9eenquZqXbWSv5gFX8GXxoQ+KhWcwqLX2nExrE4yhTmk6fo6a1QvCNHVsr6BiReIBbxqtwYRrR2E
CPtTf4CP36t8MPG58Gu8m9d45eaySUhZmnFlAZIXAs67AZkZ9VYy9Xco/L1498rjsD5TC0p5NHSB
GtbcGaXFUgijlJfsEl12YcP0Zc2fVJC7yLcu7SiaJiB09HWxNBTk40jVnLed4x2QmDZAGwwchM/T
sSVIzHqO7c3pHje/jv+pvSQo9v0egn/BWX19+YKR0Kt4X4g1tukl6+jPW+c+Cf75XLE7Z4667UCT
buKKfBrmv5piiIFLg7tmCaFL9AMGkjEGsUeEpbI2RaCXia/UaDmM/KIcctFGw7ctou4idhj3Bwo3
1/ZlU1uRdSY9wme057xBq803+p+11lH67hcRdynK5sKzdMeRDI05DE2jVt3PG5ryqica6QXyPh63
vNeIrjTAP+O2rNKskZNEM7xHxUduzQ41+rkbtDOxhMaeBZUIWiqd3VOJCh1q/mTIzxMYnTNYAebl
twVUGoP6loznZbzNDmTYsxVjo4PS6HOv9AIMwRiUhSkdSzPSWNq1BpFWhdP3W7l0qaonWQFSqiHs
kbzNYCeNaHTVFAApXB8rYCAtTyB2zYEnJkfGUV9O7pVqXMBDyGDqTUQm15/nwYb62rVniYb0L5lY
KOhwKtl30LhQtTiGRbIwdQoIoNjvL5Oh13LgIG9Nh8DoETcb5XR+/iqQ+qw9l8OCFsOHm6XwaXwT
Xf5fDRaKEmZbvYgAa21gSy5Bs/whc+ilqmAtDdaBI/CzdxypBpbYhtwQq87fetKLsyMnqEXXMdyv
u7jhAm8WI3r3MT5+yqaXaSmh5uvXK8E6B65X16WXZb+lQhKCgBKfBHf3w3sfiJwPdzqfJYFGGgxF
9Cveagcp74yliwhPN8Aw2db804agGJD3vSwLtE/KgJ+KqVegIhxFYV4gHioM34ZfviwRCej/VPQg
c2Ui0K/puSOf5MBcYlZPFfqawN1RpiIsUyRjibvatJcBvSAnDst+JbivFQoV1zMz7DyNq5CHMCq0
bcw/kK6XFCC4T9r6Ka5xYG1rIEU5AoY0ql1Ku/DjZeTn8FU9il1fyolk1O8zaBhNIICNqXGUNGhd
W+yhHhLaK0RSRK4I+MYCWmOrrqMIWjmKbN2gm6IWPWsv30iV1OOGOgwJ9SdwqQzPSh7XTowJPzhl
s4lTPpa92khsEqDX/89oKA1dMguUbcDqj/13lFUqoUVA1BQJECYKWFw1DCgUNrJRQ05jc53/3RRX
2C61t/oSJVcsNDBMycLQtXBR+q9mPTh2PZW6rMFbI/ItwWQ3ofwVP6OQmWWNHg3KaOXDs6F8/tp9
wnIbCIQbsimYVjj9DIJs48PZ6BhmlGxILMlw0HtPic0KlizSxQqMoO/O8fIfrWAGG4/xTAs8QAOJ
dfU4EgBf5gt7dBX9kP4mge14OhZBdcmJk1HiERatHEYfygWR2FUsWixlYwD7Gi6qpH3808JpFYzM
V3znroE3j9qrYtBKuS+IxFlKT2Ypu0C7BYFJua8wtYmrH7wuhKEfJmXlXNwzKtwFQQict/KzRmGT
7f50SmOZUauwE1p52zcv4ppX4j2FqdCcWpQFAF6hENWUTAq8+K4+LvNx7DPzHS4+9LHhpZFmcv5N
glpa5Hy3v6zxa02D4HjY9Ezxo9VP5O+ZGQPdsAN6GBZ3MtXfzA0xcU9+NSOB1QLEp4unJtX5x2CX
tMsk1GH2fncNZuPYmfQTZu/+Kg6gwuxNT6ORRmFUJp5m7AXOOxHkfY4k9CgSiBz0bcKtA8qgj6d+
IPPpU3mNSV7nD/KazCU+RC8y/L4jcn0nPRzfFIjWEr+iF0prXoH5rpml2ezzEDPu4qLcXi8dHweA
TtvPJwwMThAk4QJxzx9mcQs7aA5vdNaR6xEqArv1BQHCPYuYjvQ2PNHf7mr+Ojh3+W7IzcrZFuEY
1jr6nt/IL4zgx2JPHIMArTpVGHBWrrkxpGOb5vbB4SwnPymSrW2oDSuy8b1ITyZkZZpVlwllshc1
3NAOs3Yuyr4tyZjqFCRV7O1ysgb0WZE5ag20hX95yTb6sgLNoUiUGpyIy0SjZa7NN9j0GrBIWVhx
9TA2Vvur8SDhcG65J2dZeMDn3NfW3AF6DQT6R8PGEs1dXePhef1hqm7tRBQeiCXFWxS8eo7bxXfj
RPrvRFb+KBz2ErPVH6Tuuevzf2GMhz780ZfMmnCnjinCwyhKb2183UYhxllKPlXPihAm/4WBOca+
JmC0Nxn+Aa/OUixm2VWfBk3rhvA10JwAn0qG0SuaF+uVPWcnWio7vCgMkHppV7Qh6ZFh2ZAbyx5C
RZcDMfYXlnCu6Q6GXgFGqUEHtrJFliWPwqEklAWmuJoxrBXs1YKnCHb9qqcUM7V8tEnA6jmbZb6m
ygtFLr7Pk1/Mb21alWh1jbrNBbcHCGKEUPyue7Mug4m3CMsjitayLRBvW+uAFlY+fe7lVQDkBFUy
K38CI8DMlRSKzSP4zCj4X0p2G0WO7+n39LgBjzMzrWgk5Jlc9m7VC/NP7OOTs7Yh/kdy7r5T4qzB
ybBzPJZNqxmfdXn2I1RvK6+YlbN3eB+ROTGisymiLjuipNIKB44mq9NARGsndPsPgOMhHQmeAyYA
c/eJo5sGjcvlUPlhaYMXVlGvDW5O8+isWUqhPUJLxrAmaTfdd6egMOU9+4Xd3hAp5EWXW2thscaM
lF3Mws55KWt/h5a3L2kHjkyQn+qBPo85+/pZtvsWeYAdsgC2ijJAhFWqmrZBfW+0deSpsxN3u1Jv
HI65zg3nWoxMjYc30AtmCQT9QiRnFWjMqLNpeR6m03/sQKxJ6EbIAgbRsdujwfk1agAnV/zgNFxd
CqYtFZ4MdCDw5pMiiWsPOC3wytmCrLxFflFUABIBJa1TuXHjh2y1HlRMabLLpEz1FpVk7K1mdFwR
Y+Cd8p8zb6KFJzetK6yH8kVX+rkedMw+tw7trp7VVEV1CouVoq15NirzcUuitm8Pe6WnuMeexqte
HSHSTN44m3WwxXeuaDwDlTQFxFspoIP6cm/HTvBk1ayvzOYrpHrd+Ge1GFASUPQuywqz7kjW+JM/
agaEgeNIiinV/7O/4bTBtoX7ddzcyEsGlcf34EgPTK3Tea+uuuCJNh9B8XuWIz53JaEXU6jEThNP
jGeEywROLRA049CT+GJtg/7TnlAj1CEZhyNc1OfCkl3YmILeCHIo9KGjGbzgnTdYtzRrsl7ST/D3
dUZk2dMqUu4Uuap5qsaqoh23sbjdRyeXVQ9z75L6NORld+h922xPGy08ROzH7p1sAM6P7wckXf/x
dlJ0aUbtT/XwIkzedMZSbGMugerkzbp+L1/avqlHd6X6u880kNi+1W4vFLnG2bzUmTNPcmb6gmdK
Zrfwa2WnCY43Ub5YUvBhudscvjdmr7fGY/ijatbNALHznDUbJQN6fvyiVe1UE8dlzNYJN9T9xtu+
sDYf7JJijjgqa+nadc29Ix2A8udojmwkfoMvBCfJL/8ogOdrofj/wJJjQCp5udvyattK2uEJPH2+
6veJx0o6bjo/aUMoQO+vnulBVvgq7pDE4rLrj6RqViwphcGLpsKDkpclgSJLD4XBaokrEDcGOLjq
NDhO9UCD7ufPoPIoLGiiOlvte9JqxcoRmlgpSejZazTXPt2SkmqQl0D84p2PfgCWJpEmEWaQ+gTL
cDlCQHk7g1xE7MY0Y7yMZJAXBpIneXhYV3bUKThPeAZJwCk0iTkCqGyrIEWTzVwZiAdL7PAU+dTt
1bLh4vR6D7mAi0fqCg1CNd+pYyBtWHrtZtETr9oh5YusbyHsHE8P7WSqjJGFilZKx+7eFnFQ+aer
TbI3SDxM6qq3SouTiY7eMFnCQdqyE/RILwZUJrYE0vpmYczhg/UXcAhAbVKPQthS4p6DghQVpSWn
51RjcfzCGTFGI0cEK8EDMxHCTIBfs92n/6u0PbXaibCW+AQXRte7wzvAkadstVut5hl0l38G7ghk
sJ92PXYtIKa6iq0EWoPlbNuX0RPBR0mwYQUPyhxq5CKCBd3I+CDd5fI2xDciuUlm4r8FYTRMYCPR
CVID2438Zsk5WTKaO6HwFr9vwIVWJKbyvZ+Kw6HbwFILcqLIpEzo0kQkJLA5GbgNYbJNQ9YXxN40
tpXYSJdnwpL+6yWfDfNDrt1guDJ0+gfKN7KQe99Nk6MZu4KNbadb9tdmeOksRdgouaZY7f86EM6T
ibKk4lCBP0kT6WPHSO7WSPBNiVKrVAFEidZXXpCZWT3SMeX0/2/VbC3UGnQCw1yz1+uRZK2QG6gv
Pr1Kj17f11L3VCAV5olgnwETGZsFjUY3y2rPTtF4V45kab50eRTq28H6yYWpKT5mhkbUxmVyr4hI
kFtHJMJ1tr1tdVzS0kpI6zCnJDAoIQIiKVCl1TmX/PFzm55RAmAYEgBNIVMm625z88x3pjqQtyRG
pCQ8wEMhsU6Eof+w7w/xAe5zy4sB18pT+o6UpvcHN39TOcLfSA+u0Djtpiqe8gYn7vtWftBQyYJc
dLcFMp67zSativbIwmq2JXB7eSa4b0GItM7idXU6tMbDuaGpFe8CNtBPTSWIeziI0IkDedIjutcb
hanvakoiCE6wPos+7lc/uog0iV92qMwA7Doqdrd8kgq5elYCw3N3P8pwLaUtqex68pfpXYbCe6k9
WDEDkv41iebx5tVF49Du6kjh/xOeleKHdUwY6YEYWZXIIHwHeE8wqsS2kMovLDyaz+eyL2vmiqFs
+gRIYzd0xzcsp3s4fheuKioJwfjplQ5vVX+2KF6tnt2rAaNoexQ2R0WgrqLC383Qrfg0ZPznH70+
N2ketsAcb+bReqVjq9yhYq6PLKwabN/9WICFA6gRPslQUaOFvyZwUv3eGpsx6PyGdltjLh163ljc
fP7g36Rx0oQdsDxTs7Cjfw0zbwCAd+dhc+N1DzqRDZpHj4EwtwNyiKuxeExpaNYy9wKl0XOMPeTQ
eWQuQXS5uL0nYADD4w+vAqOZ9PW2nCOqMvNbHl7auQlNHbY+GqgUeis8t2LCdSJ1pnkz4BzSOBsl
SS98wChFbkplCJ8HLaHptmVjxi6WnMLsiQqdffAMxpvhlvCRbKZPbLgrm6K4BWLvMtRvspL1GpWM
cM9IPLVx8dt2JLN6z8KC2tkvpafyPBXZua+HGn29/43odbSexwjkolcjUUYW/YLIc0i8ZFB6LBHh
0ndrt2QvdX+XKX+iJRqqcxAgDT/A78wxhvGPguB8HhKVvl4pSYUjJ4eW/W1nHzdAy0Lr2aExKZIY
OrE9EVifcnH8InHj00EJPKGs5EWv8/14rOie8Ury5zi9pvnqvR+XNeAqauM51uFZsyvAbE7QteJD
v+WvxFRV8kg3tU+iYX1x5erTdt+EotG4rL2GUQ0q6qBOTPAXAM51S8x68QKV2r0KIv23d6An6icP
JIPSFRDUaF5KK6ZihV/SYDimtAaP0jd7TpSInlyp4LrAmVpA0eTeB5nc8vAokTOcwqGQ/Kwe5nwc
gkDbLfC8MG2F8g7kwRUZr/4BJ84rFzGD7ODBRCfNCUvlnxscoWzREsxtHZPXGBh5v22o6WjO7uMk
AKm+SbdhML3TCl4akWKPs0nK2skHc6svJkEaWTGrTtWDVeHdbtD7Glhb85CFbvNEjoBUiRRcMqHN
vSi9RgM7P/MGQk3zTIt1QcKGsWKhicR4ReK1d+LHRQRLp9MxxM3eeOytB/2V2Geuyn1cWyb70JXR
PGhUtdxi0rTb1qPlnAtHCpIReQf3kjzm+qmPR/jXESK5RsXWVYrLFfEOPqI3vX0Mqy3HdNYiGCPn
vyzP8wtdhMG7fSAcJEQ2c48kMhuRRpw3Jg5tQhi9W0xnQG9Gs7fCjNYvGovM+3UD1v3EYtdlxRvr
Jn8qUjWej3kiPZCOWcW+xv/7aRoI1iJorJ9J3MzLiFUwcqY9Wvdv/K2T8aVo/sWiNmqlJ2GWg6/P
czZ3ZlVCO8G8Q1+KC1CC6zlluKwzriDELKvNBwPo2NVJhcTqecwgvZcfG8yMYwRTTWpf7nxJ3rK2
W1Gk3hZeoAi9hg4BrljSfOH0shqYSTlEugVfws75rspUSPwDseNh1uj3WKyaxZFZ46snfoD4b97a
g6xbND4YnbIhBq3ze8mcWH7TGnZeuiYI1rdc7ehG9I5mvg32c4jmMx8uqB5bFTwq3Z8IxohPa2ct
9zsCgviu3VORnP6YIDzpJr7JFOCcqjhTJjEYqmlpj807FmtJr5OmlM0Y+mxK6Iu2aogFrZ39tbJs
Til5ZIouIgTLZh8zXzXWwxooH3sXCp4+9CGDnJBNX6bKlyYhSYtpJp2nXPGmvSmjL/NYNL13c9rd
O+asIZgX1ojFibBO05Ioy5wGMysCsYDXc3+p8CEVv2PW4lomuvXw0JSXszepQqeItDHjg0VQ+c5z
rA1NT7pcXQfsZTBDg4CPNPDEV/1hzzqLwZlOp5YZ2X8Atz/LPFny5+HSwrTXCcAg8J99z6zib39I
kwAYu1d1173OQR+i3R2/VNNbeB3QeJm0yYDU5dF6OqypIKPv2eL4ipcaZBFiMG43/KZEVGEjC8r5
YXjpIF8KftORaz7AcJi4TsUgkStmds8+imN5F/k7JARWY4DyKhv+8Nn3cF1nbeeYlckjpAMHmYHP
xqOkhC4VYE/KGp5OpGSV0+7OI8CAJmQ6iJ856O8mRqRE7miEghDJ7omztQUa8JeE488frxqtTPj4
tCIoZgLX3YDJq9zxpLgst1j+vkzcgpiqMzaM8it18kwYmTZ2olfVfZan5VnZ4UtSC3+mrraAhBuw
wzNfPgMs9QZwb8u8FITto1WVd7hQuzV9wq08TxPGOyahgM7IFZjhZANUx9s0q4hPFWeF047H0EQ+
feume7hU6Irm1uTrjVL6438oInI2B3/mtx70nXzn7ggZWI9UJm55U0IGS54V419YEmeceQ5rprtS
xlw7NpAB4G1gFAXApc1C7yi3XdtfsYrWr4KbBCsgswCTmrJG7Tj4F4Uebta7UYjx0XYJomadAoHH
r/JrqRw03fFtsxl0A9o3yrSzvAYehKMjmMXdYAYh6+AbJVto2QBx9WptoLGR6IGglMrSXYBQRa0+
hQ/Sv13WgpFjf1LLZMAUbdv/ffvMcGcvOR3nmhUvzJ92FVteo+xyKfgIht6kqy5ckTk+3EctED/w
QtyWiZY22EK/SjmizpL9xspf7PUHh+dQIiB7I7ouPsn348sLqwCqg5Pdrbwv02z5csEKI8H/tKkb
bbxwRm9vmYTuIotaYdq7PG4QtUGSTkGAf9fKyrvIQfcYDHLa4Tj9b0HxFSwcIvGVI8YyASqVsqqi
VoRt+auk0gwBVcvYBCIIapIX/w9Xme7LzjaCFSOz5FV3a5kkEUoXEnWXKWYomqKen1ADcD9fYQ1z
pDwaWQ97QD3nZb0NEu1pHrL33xHcCPwgIDIGU9yu2A/QA9aklAFXZltq5sV2ldGD4jTslQ0vzwnU
LnY8iOPXjuSx/T5jh7DXxAFvsgyTgqZzc3iySTo+seYt6seZpn2kEWMimkVvCOA6MR/Fcma97vtc
Rb4r9Zjb9/8CGDEpaUYJvY+eUAGHfDqR6huP9wz04zejzT8tehCUmvIjEIfFLl60p5e9U20QrIQg
S4aSXKnvhUIMHt0laL8y2wMhnqcOFA6bgHjiCOoRUXQY+PtgfnGAxRJzweJc3hWYXdaR1Lt98jgF
5UxZr9ctevx4SK4xjBJVz0NqcJxcza5Rfcc7r/nL4/oC6MvkjNEqiKAzEeDy1jMtMN9w7Eie8ivz
qExWy7yr0cb0NLoAhqwvPMzAZzUa3UPfvNcqnTKzo0IKVYYFCY2I7+CyoiVQIy+fH1sSaad69SBJ
Mvc1ccz958D1OwTYMSuKebeyQlS3ja1wdmRPUcf9JK0/v8/Qx+2uzglEfbGncl8Ly4QycNXezTmd
N27QqBJJpBr9pWetnXOaSvZnLCwwhiwLa16W8AjRoOjGicQ48HMDZQCW6oULf/wJjZ1x/Q4K38hM
X7/I/rUjC26FtRZFBoWv5M5Nl0+sVwd4IrjYLDYOss4AliEZxYaXQfdHPreE4uzlETmuD7i71TO9
A6r/9QD8xofWHe2tgsrlGWaQCZFs0AWpG/pO3L6ku6vkMTjqYBx/dDckmHE3B74fbPJpHOGicUzA
p1oLLAkLSDu1Xik+9LIJl80x1DymX+yoRLNKz1uu5di5vATUjANSc+jOSwlkYQ7AF50JstAGklm0
iNhgQXpOx88E32BradLPrjC1XajGUH3AC/EJ+zaXrn5qFKz6EUqVg68FBLq6Xte1wZ/d1ShootrI
eEmj56jWcbm1qpX756tmSQgNAu6b3HABAgLwUKwQMpvpF5Sgh8Je0zkk8ISpegNXgj0AqdF4nayZ
ULqn8MiRupetxRLUx9D4ooz6yBY2TCe1hPYXmfhjM4XaEAavY5sghRkjiMP83CveLfH4HbTrAT7E
3HqSRcW7GM/ML0tJcSxs9HId/zhnqyQOaj/c7fc5Ax1wcOv6/YIELYBbQAwiEh7sWWS3kw6KR+Ql
G3ZpvSwPWjJD27VrCcW3teGMv0YD6liQUOm1zLSg/xA4p3pWDRmnEqbSpZOtJhw7LaAJ5TkNMVNr
QR8xQfZTk0iFAavBU2Cc7pVYU+88DcuRHISp87FVa3mhsK9acMKqjOiPTLjE2lKw1E3W4wkbjHJK
M2mMuqxnh+bDaNMP40ggmYtt5pgHRQ4C3dRcemF+oPwhLWctewL0+7DCWkZ6sjPPjnrJRaiWurO3
DHDxK7fcOir042/Cl7WoiXMU5bxsv6SIFeUdneU0BwogL5nxwc6/wmi7qmzxrxoo8oUOLf6l72rc
vMV5KhJK6YSIyMQyj8KR+AXi0lQ5+DLWn1Anbky3xubK0SXZnzitEpAlEZJ+tyLcQHeiFvlupOaT
rT1F82CPR0PrZ6wlSYssULDk0fib1JNGatvhBQ51M4iIEWYskbYv3A8jEqRoG+Lx4aXkR2AsYPDq
apNWsstoao7jQ1jzGr8OApUr6lLQIEOdWuco+qEPc1QpccfoN2Cj1NvZ65rs1oKFYkTdDD+VLZzW
K++yju9+QIRINEJRwcqi8ykh71iYR2sD8NDby54nR2SCh59Qy7L6Q8oCvA2MnlrrO+Vebr/l1R4c
2t5NKgQwnXLHNAKpYmi+9ZrhSVjm/IUdQfrlJilK+LzIHC32MVNO8cACJE1V9RTJPgVX+ejaEivE
ew2ZHUerhS1li4/rmcXSGlQxXmMmN6/7t1XV3RExo1rTIp09T/4CwGIunm0z5l5Ps2Y3wpagW5ez
yr2UB7QC26gMvptr57WUWNXRTDEEC4+2TzvIiJ99J+44AtsdPwUpfY2yhzNz+d/pUjvjFQVFvhkh
pKGFw9cMnV8W9h6jLYkCObL6pJuR3vfkbhhh4hS/055yvKTxKVnMIUPHTbSlJA7FZHMmZLFT7tOt
hw14uS9xqxoKID4zhvId0VmVVDcodjbz4s8X7ma1QmycJXAUs2M22Q7H2wKVTyL/bh5Vf+z1ubsU
U9n7mc/0wueY+rIREXtapZ9y5s3+Mh75u9nerRuVf+TMHV80o2w20dd1ncdG0+Mdk5UdJ73dDy84
GO/SpqbuEGWDrDih3x8QqWprs5zaN1xHtBtFLgEqFK954jkVQRQwakieYcduTNnXevqxbS9+8h+C
iyHa4m4TnljnnFZwvtUrFW56hJGmECtMQKPkmu+T9PjvDbsIpNv+spnko9MWI5dhuc0ESguBhTrp
rfQiieT5vV1MmPWDwbkA7s2punop5WEYrNvAZ1ty5Xnd7LM3Fc/aehDzGVuEkjOw1vaw/dM4bch3
m4DbhUJ+RSAcKXKa2tXG8oSpa4ze9qflushUKZErEFuPpVMAkgN+UZ0dSN5aFHfhF4jjOiwnMoGO
L4TQue6AFcvnI82M4ViLrbmOQcxO+a7Z3/42jwAUR0fmjGS0/z/79uPH+pQ4NhAxqdzRyNS6O6SR
+w1ETS9FAiCp098Ve8LPInx4hQSLS/QmHrPz+Q7LSWNxcUJbdz3ki3SjYngVP699p2XDaJkhRdCu
SarRW3GbuqZPfRBdoxvHpJ1C7tG1AvweRPtUdzwbg86UK8Y/XrzSM5miYzkb2wAmUITSS38Pq/BN
lFqnvkBqgIT8epq471laZelsV5xShs9qg1Q/n04P2ZYc5+Ufz/pdMvF6KBt2pjuxyKgq6pPZ/+Mq
z4gSCGDPGGzvUEPDsnXqdB6IvSz86frYnyzdxAjaXE3MOK7bghRzA8mmVr2NXOvVFiLHWpgAMJsM
KuNNw7uje5BNEif3U6J604BuwezyZbhVhJuzjETvgvUIermF0qCkW+DO0A+gGV0+wzyUcvgc828k
qD8CujVu5Gketf+QN1C6cuu62V/egXoLUk5iWqKQc+r7PEjSwlPQLWzoDcxCeye17kMbq6ZdKsG9
jgpCHhGOlxGKRIzvcKgB6QahY6lJr0/pWQVTTQ82UcbjkeIcuRBNh6TicYyN6kw9YH1N0AVSh8QP
ZeLiDG18Fof4bK8iscDOHcUqoggj4tVI7i2xNHA0C0vJx5XoSK8NT5fIUA8fII0D649Xb9mih86A
jm+7ol9R6qrmNMQcpt4LvjUEvR2EjT0zpZ5hWxIqenuAK23TOqYImllHvYEcwk9QUn9EjzJG5ew9
e0nYgHg3s8seazAWmpqSm+N5+R7YYMnYfDmeinF8hYW3tlWu4CvixI1fVWI2ilWW3plvHDy3k5ID
VXqbThEzaLCNXfC/I2vvjtvvCI4KahOf8h9UTyfiuQc9jWJ7MpK541pyVruz+xXooGQzR6WcK6nD
DMdsb938c28VjVyM63pkXhyNtCDAt24j5rrPgJGocvAfNRpS5PAm61x3KvjcIModKQNqABuW/mV+
WTlFm7xh76C6eVOv+O4GAlfw4+HHQ5ZI18KpbyntMlnO1J+SF+4TNYv3d4urPefv5IJSn4pl7NCZ
fNP2WZbMKEX34voO5OS8HSK6FJCVN5Y+mgVKDAMDuxARssKUbXqFd6FVhNPmLVXXhX2BxMRGuqC8
gLP51iVKBP1Pw7fA2LlvUD+1s0+xssvqCAVaSSOFggJEtcZyMzFXMPCsSOHXwA6vtrMpOmViCAQI
YZNwjbG5Zdx1X5JkJsBgyQ42BWc02+LSQL+yZ88xplvGSXdZvsVBUP/hiug4XmLmF/gOOcbM0lLi
gaLRUBQaW9FiTtepME3j9apj9/ajjXIzl+L66Te1rjwOEwZ+Vngt4GcKLB5dNusxUR1tjXaHrXSl
+7OZnCepZVzV/G+Dp3+a7FZOmTGDPayIpnK5+I8P2KtC1gEz7w4kY4KSf2/5J9L/jx0lmUqU05oL
PAVZeVSmtbEJpU+HtucoaXAQing4S5gIWXeHtot9vgoJbNiqXqKIfIYAz7hpfZ5etoysF65lade+
yB3K4DPrTS6CzQ99V9KVlOq7G9hFngtJhjfOLrTFpVXzzcOLsM1ZBzGsHQz1Dl5fkv8B9NFrn0hJ
wWXatlOix15k+7EJvEf8HwgN1apGFkOA1C7FC4ZclGxuxZ1ANM8LjEGMqSlhwLWGBnfukNIi2GZm
FU9SQZlTfElER+dbZ70TOJVmFdVR56cUsxtXNcunvcnSPHDfoI6oRW932cHnLD9ZmWjmYCjZH9zu
rojXrYbgyjqz09JBoKduFJqimOjHNl+IdkB738hoch7iqV4OhRk/prLSHtstCRxNXuUDTCDpto6Y
u4367l+ZvRZtbGgBx7tMroyVE/BSFkEKr+vPQbu2yGXc8dJnAsxuNNeG7kWqpkN2jy6iJ6SbQB8x
MWlD9FC7ZotE4i0cDB99SE/9IK3iL5sd9PJTW12jdWTo8s7KlueGSES5x10lonZHsUTTIGlcHaTt
KMzGXYkOkS/fe+aSsRs43d1ztft8NwmvyjsC4NCQcsNvyWBnIBCkze2T2777QKHDQPLIqMAmVyZW
zu2/BKm6iMHOUVdmui1n+tBEM2ms9n4hVi/ngj4TfdSpM5mDadThEcljce5H/lM7HLYpdD6zys2x
N6nVZCFcE/jqG8OqsJjSeZaacBhZdALdgVh0/Fi4iavuIIM+YtMTlHNqYv/Chds3W+K6ZIm1OMnF
Yf7AfxUfTD57mYGgfxk3Bh1M/weh+kWqBXYt+ujgoBRDQDOcTOn7xYwUQITpxCSvkf7Ey9vP3uUx
ILa/yHr/WUPhgkmIVFNAdbENbpI220Ag/BSnAHldVx5grx422hhKQgPK6S460cssn4ylNdY12N3r
UwLtEHPmRxMI2SnLZbBTaKrH8ra1SUAIdvcRTuELJFDrjlpDc5uhiqElCI01vARPdBbgkxWh2wI9
s7H+MRzsnDdtWZa/+hEC5SadVS8TYttNJgDp4aRznuPjuAn/UualVRSvOl/Ml89/XXRexbaFhKFB
PmdL4CcwLQq6UBj+IUASkPGDhO9GE3W9LfVhu1nS76VZlpoDTT43gbSbhhCRwtQ2UpyFucO17/yT
ZSgVyagWkaOWOZcuRiKX/ELOfS8OknPEpcO90tS6p3eN7lVByLqra3XWnhKS0Muee9j0uLA2L94b
jxygsuavZymREWaF41g8gSLta6Sx18oEsaa5tthe0zASxByjePNdkD0B1P/fdnMZE4VT/x9gp5GW
tK57l785z+I3x2m28Yzcq5sqOW0Rl2DFuJRGUEJTdv/5Z/1ahl2fm3EKVPdZh9AGVmSaNtoq5ekK
QhCvrLmfgnWdsWQe4a5G9SsuvA0JUPfiQ3dKPwEuJ6C35woK92Eeob2Gu4E5XU1R6gvnymLSmPnD
yKhI/+kviXDIe4dgWTMuY6vbx6O+25MVTheFbj6JX4Rwd4v+16Opg8dhtKzBLfeEqfgHhYottrwi
Sq8qPjEHnLWJSt2snnORmoAEAz8jeZagPz8pqjkc+FVN+R0YS0l+gEANpjKjeSYhMkPOlPkhqPU9
p5zF9W+75pxUWYrkk/lgvpUpT3J92frryGx+3ZaHdUhcSZuf9T8ClqDyIh/VjfUvxEzeFEIe2Yrw
nJvvClxGz/Fjt6ZiilK5JEj+hWMCcYUP25GXf9qEu3l9SmiuGdCOpqmzA5Cd+v3lhiCHqQtF9l+O
KMgdSWTdZtiRVHGHUIeCKDjO2dH/ncDIUTy6NeikaGYPUbry9HjjQT/vKHQ8aoOJ+xIHLBJr9LT0
3ENenjo9cxP5p1elIby6v9B7epnkMtZBp3KuzyKVmGQ/3GMeS82NLWJEpAu1jaSKH+Suh27XhDvx
AWm/JgaDqt8+RKTZL4gF/Z6zjYeLUTykD1WpjT8iSfVepWU0dITW0MMkbhtFwTBOdWbWpCDTEYDH
sfF5p/O6YUKeesI6gkO7NvXTydpPkSP6coezjV2M64VqAX1zX+dVv5KINPyr/QPQ0YXsNmfenocA
x86i1J1dL7X1IkGiSGxcIxeil1FshINu68+hVzeivFSORItJF4HBD0O6QpM53ScpSNasnV87moyu
bZAxe5A4jNSMIziQt36eUfG4uM34c7zM0Kxollr4+NmbcGfCfsphQpBOKcR0V81SAjRo5TIS+3Dz
3PEiUMX9trpCVpAOONGOZ1BlS1a3AszpClkKP/wCC4UYZ7i4btIvzrY16zZGDKuyBVoeG28gcgEx
3HZVo2/h4w1icf4N+ZEGuMyL+x/QEJVR+Le/oviNxExuX6k9vnOh7nAg7GQnokfBDja5hzBJpgl1
BIbaEr/31O11iCfqVil8A3qotX6360YzErwGOfzTD999XRlw+taiXRNYEbvtACQWIkL0btIM7DCj
oD5LvYHOFKXQCrlkOwcB8WszmbmRZU0j++1FrHUz90cyWQNB+FfnOI7DcUPUOsd7ae0FmQSdRvD9
14eq3l/Lsl7VQlFbEY6U4rjqK3wn89He2TaDuMC93xsHFCTBqaCRTmPrFrf017JW05EE4SaoMOWj
EMT9F7KnqEiRl7KmnKnIhtel3PreV9tJmWCGgtkgfXOMaVxafWAPEuUKYLW2Y7vSBt7EOzOrFEup
cnigaM3Z7a6kDPLsxYDHAwTguCjDZQnilV6bVI3gIWnonGw7F/7QQKFYd9ggxYheNMhXI/Die0zN
tAkhPmIXl3A8baAMpU9jkS3jShROfSYmbIeD2pq1XaqwjCCoPEQ+ZMFR59ax7GpjhyoszApxOafS
WPmOTmYJGTVMk0oHvS8hXj51LKnkK7wk91csNDoapJFavqYhvtMWUVM8UcwwuPmvDpe/0EZdLLbQ
7zdeBLUWwjS5soWhggZerXmMANgmY1VHZHkmBLYrvf8xUsFnDR++xXgWbXH3gIGZ0YaTO09WLLg9
gB7P5XezAekf0z3OwAvyejhN1t8askdy8ABkgQDH2RwNruGrfEzOIF/+sVWD2WHhlL+JsDJUjdTG
iNzDQmGGZK2CkEA7oX45MByHEWbW+I5Wt5mupsm5GgfKXpAQ28uny7fKi5eQEnz5XSIqqoYQLjIQ
Up2rtnX0hGB0vhbhBgBaqqjfwOsrim8qCrOssGLZNLpcqt6BVIRbcVvrOWZ6UkO1KDlEVnBKjjXY
v8FU9XqQJhkHU/tsEiIwaBJOr6lnJoOwP52XyuxCwC9INZbqlEsad1YhpOrQVXLmLtUyoyJLRCMk
S8E/HMG/WWDa8Ey2KZIXEU8p26guEpqXh8hm6yiRtXXwHY1GXsYVxSiGbxg9oGtYbXUeGT/0kRMZ
ZHxviW23IZ9t+LwbLOMQJBedkIBaCywUYx8DsG6LIwFDuxlQ8eJhkkVf2EqGTB2z0+JDVWh2bAP5
27GVedywrQMRV5NvQy/HsSpXa6Md46nAG730vtl/ngL6+pcQVZAfEDbF6mxH/ha1/h/EquUa6qxu
r4nXztr9jZoaUPdee476aPJKj9QW9PR0+9bxPxG5uGUjzTA4hgBHzcCMk6e3Ek4TPTz6nnUKrxAr
OVhFYmDhxXTHoEYZA/DyAamL+ZLH1z+x0ieVrb1EPr7RBZ/ZxhyoYFzpDudp2LyHJn+hx+p8ukAF
VOTTOhbiqI+zJXpl1DYTCpwUFDHj6mU9rrn9pa2SY4f1cIu6FqdXuiRVFM0H+6FzhfjTyg/O/cLX
/AI4hStl+C+xgiX5xeQRht05mbHUDr340rgiCjEVeVjJ2Kf41QYn59C/fjqcdD1SrT+iJyQZV/k4
YvycCvGExmAWu8N+LqTga321bJEPkW9spPnUvaMUsFSJcyORY8kPRs0V97kB5vfPHPTQz9ePSEgg
k+mycFv6v6oLFIr406p9loQvua/vzLzlrCGJDVPriCL/aYR70+n8OUZyJPy6UW8qn5Y0o+mQ8/Ja
GJTnO7So40SEqoPv715mRoqT3BDb1Uh4w1NoVGWKvA85XyrunE7AlefvGTcyJK+yM5XJLxl/J2+W
rN5z2n758ULUmx8+F0LEnVEmYXCfqm8IWnEd/A+e4ClmHqAHfS2lMaBvxZfnJc/kvLRxebsmfPdT
tvM6Pt8TxaHJyyJFSJ85AppjONc0gtVQ71bKbXXLHhx/N9KAFk1fnsQqOAa4p/LisutHSEKT8YUG
IyNn1JQ5LNKUxDNvJymNsElomzwEEAbt8mD25Q4KeWbX7u49S/q97OGBWqued9hql1RlmrkStVCL
am5vdBYHn9reRG+c8HYdAlQSyzzR/SN3EZD1k8noTCJ07cbJl2GA7xmV1EhYxNJ8LyU/BscPPq2Z
nO9YjcYLZTUSwUuJbuGBBMvmzYjbLB5J02JRU83LTLM4U/ftHOfBhwucEUXTHyS17fpTPT2aNszT
amRr/VAEdXwzlutboCLJVlyyTeUPUJkBvvqv89Z/D6U8wwCyeonGaVQVbpfvK/mhdwXW4SZDUrq1
5cxZD3TUrjKmGawqDlE5IP5Fw3sHnEiLz0VK41EkeWksxV6Ig5m9ADgk4wgMzhf6bcuUo50f2H4B
1AvPv/EcPUKBigllNNlM7aZBq0Y9tgeqL4kP3X36ZPt1hCXhg/dwMu33XADoPtFrLCI3XyKJbVo3
KVC2XO3M2sf+44cUyeNZtnzycXzf50f/ajvMB1K7xyj2aRYDdQV2S41THUaTZCP7TvvLHwJpYTX/
08ngQN6CL89GVtBc9zpDmr4hbvwVCU900FAux1P7VZrwb+5qoV0UB/JSmUXap7swOeLqcq8DdJz5
7b5gV8a1VRwwCn+wB9SBgP1aSY8jf2yM2uGGFyDtHJ6K3aJDPE6wWYokc1t++TapXKB6zD9pNsqj
K7aUcJhw1HOUPXr8C+iQLXi3J0HkqeNg+pAByfhjNkrwAhfyFnBUnKVd70CphPr3cdLkom7To4WX
YIlhkU7ABXPESasqH2QCDd7eQ0xodAri/x+9x0RUjSZOf3Z7K6LtOHzuRxw+43c9bAsSCEhXJ5Dz
kDDKZPAoJnN2eo7cjoOORvRsebT2oKN5Iv0RxkDl+IIh3O43MaDpOjViYEdaoE67Buum3MfiQtVv
G2VOZVmzcBibb6UlGeR0KHSY8/E1+pvqg+mNHbEaYIn728fsAPkm8tKzeb78TCwdULGjRf4S+hSe
on/8svrlxFgEgu0gBxOXC/LV0platIa+3wi1wbLQBiR+kc4rorRXorKEv6OPwPvLhnC/Fn27dwrZ
pPzVP+Dll2GcWbLbKx9IjyKb/EEytueFI+w+zssiTliUlmiw0p6zw+DpBo7bCDD7R2+Ks7inHwkv
rCQcblX5zMOzhTDuslayLpu2jFbZAVgsrOQ5+JWvwRkijggjjmDKrOvS/rk5CEfwSMJBdBnKMJcX
VW202MzjUZQasYZlGKBzo9pp/SRSK6JITwvmp9+VDL4RR28a9tQArF51mkYHRNA6+Vg6lZKjYLax
MJulcVT64+9h7sM/Lz7JOC3uTjOiQB7621atsh1NmT+ikm0BL7Qk3AcCkTMJnVltadVmi0kphn+g
QWLjb2ptHT4R8ldcjEGRGErKGWWS+q/9Th13qxQgvvq1RRFWSn1Me2hMe+Ks8gg64VZNrfNFmBZ0
v9DR+1qM8Y0fLONq4ZwUK5BfmBkJgl3tUBB89NwJOQV4NL9gd9hYhyJoS1pThTtfwNu+X7NQlhBf
UpLbs8Kqu5MH9pYo8GcliO7cyzPR9BgMn5a7GHknR6eb/hhsg6XB8mGLu2eQT1HqWgsr4nvsLa1J
ZJWJiHjVO5s+zDEud+4P+UUoayUnCN7nQn2A/7GhE0N9mgdp3vMXMbqc9gfNgHTXTDgqRc0Zz1WV
8uFhIUnSBcOMkoiNa1FdaPjB6fqpSoR4j6c4N8SlgvGNoRMtYBnbTQP0/RECxf5UCdAVjai6N9F8
1Cx6/OnzWiddRPmQ+VME5ZLMSuRtmeAnHxLBZdoG4HSu0UtnBiRyYFwC8JugYs+Rpyag+Fhizml9
iM09Gwu7Sm2sCYxHMia5MuI2kabkcahx0CweTQz368Dbp24RsDSsQwLizjLsm1J+mpXhlIw3B1oC
d+cQPqYsG4P+Teel29LGvxifNCqX8L1GWapGjSbWSIBE4h9Sap/x+hMv/3dhMl4ylG6pDN4cr763
0RsPEQDWg5qPOEGyGle3Tw+1mDxyMVwPiQbJDclJMutxEeQjWsciMdCNTW9PBWJd1x55KgNhzpHO
lv9wXYyvj5dTZH1nsBkRAyBy2CunNpju2yawKXu8S8/877jGixmfckE6jKAHpmeMzD8jhPdvUVmP
Tr1ahrY6eMM3MmiG697UpOiD0sXT1PvSPw/wyghhRMB9c4f4keUR9pu6zIZJ4F/rsqQOdb8Qj3Xn
iI9apFr5rA7oYhEj7CrC2CPZ1GFQk/VyxF2+QjQWz4dUSEsL6Kj5eLXAYWsDAZbXbfO7shAWTRzL
HbQdlGTGcsV83ZjzfZKUo18O4DF+UdtVz+fP8Ev5RVDyV8zzLShj2NBdH5uweFTWjXBvs2YQ1y9E
FNzU76Ccuk27cvC5/5hITtqXBiZYmqWkE4gEb73PDjdqkgP57JOi+mgc1waVorJFOYvSuHP62fcZ
C4Na2k0kYuI77AV2G+3G2NH0gaWGwzvdJ+0KuCzI3em9w2vbn3EsFz/YDIt8dkdt8Y6nqUTGqFg4
2KWdcpIkAhuQATvu7WpSq9GtLCIBsqet/2n3vJNHwRfKFrr7Ie6QBN7cI4kU2iwVxeTMr/YUszcc
gUZCN53E5n/0aR2Bu/zAEQdRrPziO+iJQfABsup8+sD36pfMNiwmJjUm/WC/v9M/4cpy9PkvMWrS
1Vo7edcsVS3801z3iMuZ+YOOcXnIugCa8mxoJeA4jmWxgqax3ouyWnR4aHyQ5wNkrRKMVue4wFBb
3ULG7ACuLIIasdAEUAGIS+JvJYV1ang9Naqt/DDhu4Msb9fK6Q/XPL8U4n1JyZ9Lae5p2xWxVY9n
1z6Y3ly17Wxfz6xT9153jCMsaP3J4egajEd991mfpCrNG7OokRZf6Y62JO+6MHcoN/buYou1W3ER
JOVu2c0v/GtUZsH+qtmLrE7G7s7uWwXz6GlBZtjcEnrTpBmR4NNOorp2XcSW2eAeROwh/TRZIqe6
Knj0vMEK/l19maBQzTIvu5vb2MqjUD8gO1JyzUzDdTYovt0ZgVoT6OprVTGjXb+ivz10lu387oz0
nUnRS83TTq1++nqWRvXtn1U4Du+m4kcnPFigQHxdubklc2KJvN7Vo9fFecEmfuVqtuIm7zuLPF+s
gaB3UQJrmaZdCMIVAUNmq0qpcnjmv3rypNRfjjld/YFyVobhCIWFOBrCaO+E/4tTzaXlVR45HxjU
CvCcLr1htsieg7x0hqsRCNbszGtfjPtpK9aBJe0sq5cjVzsJKIEayvZiyy0PoFbFIiva+iGCIX+R
k7FXrd+r1nuZ92yQ6E/ytr2eUClYQjo2uO2nNy5d2hXdRuFgIXSuP4ivZmbg5ilUrW1waJGBL6Vk
mpG9/COFL9XCzh2PeyRZEDp+9iU/+WtFEY6uJvPiAlKNuU3YvcQ6BTdsv3Sw5bhAHn1Rp9+L3Smx
h3YBYJm1/nG/IgYA9SJPIYs0IyyMZBOJ/XFdDn+l2cwSGn+Qx9Pt47v/hiGw7kIsdMmqBOzV7NKQ
JtM6OGupJ7QKtMI0SuZ2TdnDLW+VZ14AymvTVQ6h5UcoS8CIP3/Gj19Hh33fqGH4iy0G4rFVv03N
JDs4IxvB9K0+tkVPDDP9D7tmMBX8/kMpGp2JuVqEA6FPcWegFTOAVyGZcAy4J5p3NK+6mw8WMIXq
vZ/BABLMlYAvK1T/imvsBAb1ipzrzNamf59sVvVB0/ixr5caiPYyx4IYkNGbJNMhmm/Az297e7TK
1eLqlEc8rBX5YvgLC7rUGOU4F/aCQ+gJiRxo0b8iCj17cqKyhsG4gOG/nhCBGy62WUDNmRNLJd78
/oXseuSxIkp4kFTIfNkEsCmCyj3wdTx6jbcOd225Gy9om7UUv7842VU6hGjsFt+C1M+4Iye3D4Th
hOQ6hWxjv4ykm7uVtW8bFyN5RRfvyN3KMfprX4c1wCGNF/XCkB4jWucC567cVxN6DUo4a57y893W
ecCTFuS1IjUCaFlwuVrpBn2A+lfFuSgmqLhWQ5jI1AcFBW1ZGvxbwLdV6P9sl1Bth5rzN0/0X9dL
6UZS8mP7udnSWbNIfQxILWbkhYDGdBDcwJ9hny7OBiAHlBWpE6oVf4duO2RervOu8fYkYGaqn2va
+W2aG6RCqecy1zvheICS+zNwGcHMi4grLclo2lwEUBf8iAyHTg2UOuSM/CJJl6Nt8+c+jQHF8prG
KeSgaOYBQI23BVsNyKOkD9gqdlRl1vOytFvKGTAueI5GD/PFcgdFnlGyUkb+ldt1FNC/ourfupuj
cCPKpRY54DxJOiuwSabqmYC3h5KB7didKFqFI5RHcJBjECTM8xDrE5zF+hu3kHoToRzUHSI8w9QF
gB+3Uz6QNZ3YHxeRbMUMfszKpzLRoogYyn/OucrhM37mouR0dA27gHHP1l2+T3qyRSFbDyu77Row
oPfff+UrifrNai/4UHcVkYo06Fevpk9zm3Vvx+rV/zj6kl0dfplDb0JneAO5e/Tz9uvE0DK66GuL
B+CgbZIzOJYi28Cq1ANDcN7TuHLun2izwhZkxLMU6fS3XjAia0thekAdLaTyfWEBMnu08ed9f02m
4GOmqBlhmx0Sj/oLEiNfSLbb7p3untu0izB3DekL5pbyfB8QM9k37DhS76SkcJLPKMrKRO+wTiWB
i++8ZQLmDqI8apQURTOeeZjL+qjGpkB6hERaTQV/AcOS9V5+HKbpsu/pvgIU/h5NJQpZCXaf591I
TqtrXTgwA/QqoL83cN/N3JHwIH2i01pJP9eiBb8dpFr4U7NxY5JRshP+f3KyjBds9Y285VqmVsGK
Vy0uE+G+X058FFl7U6MsFFbhlzaaFXDMr5OvOy3JzU2FkGaBdOC71lKSHTobbVYnN/9nvfMJyAOH
SYaYoWJvodm/UmYr98B2cH5QnKTI4UPIrVCMT3dcEe+m+wmgb2s95bAIkXtegpKxwSYRh0xK+UnO
2IlIUnguY+CJNoac9Wp+fXnABETK+eJ/U8MHFBp+MpA3b4xKBM0Ws8EN3lJkHGxe3hK9X33YcERg
cEHFrkMJUPc1INM1ZC3g4/5GkBCReDVJNozgOEbac30DY/GdMBvAfTyzXOr8FFLyLDQZvvMR24m5
8KxTz7rwH+oMU/h7D5cYjkcJsyYeK8DdxR+GG/e6OGDQRLDXt3xNH1+5GEscly5q1n0/JMFKCfjf
FgCcjwoP5Plzq/YRjBAYyTLrBpCWOcdXjXplgbJMWwy/Isu14petL8PllsBcddWSX3mA7kht5tRm
C9sHP9WCvS5K13+nPhnPsGwTFWjfoWmax9JXXvYkFDdonNFBG1ZKsSBrn239esxsrdX9tkd7qy2C
+XqiTlq6s3Z//U1x4kKwTHuRgwLF9MdWaDWuUjLS3fJCXuCL1LL4F0hH3nW0e5ytajFQhvko7Z/k
/9eX6sE+CKveM6gD6OYLqSdnMdqQCLxdDnFO2MzZpTtZHZ/KZifm/5jOhf5tTempfIg1/fsByLvT
rvoYQLYPkTdTOftW1qMU8nwbI+YTkHhga3MMkHhHOQE4vMVlw0lUVTLcSZKLKhlvQplN1FSqSK2R
DG6secevrN4hq9RKqBw2U4k1+D/5Q4Nb/xcZuGhCU7cfEXjFzkR9/zGkHlpPc3XPFA2huflNiptD
+T1wjgNnMhimWwvQn2ZzppisneZzYCaiv5QZG9woHZBLUmOQtmIVhQTT8B8T66jkXXpJyFfBefT/
X25GElLxe7ybN8L/a2soHUlmbtAjVcFMa9/fOngXQphHLKA/2/tH6mWezNklKBSG6+YHjPN66vdz
C4Az6AedmGblDaNqi177az/s6AiKZzYws+BCI2ntbXk4UVkwu+DvQWAqExcDlIbeple/pVhhjcaz
3w0hbTSvFkhI84H1TyWc7KW38SKyYvB3YHYFTq/+5sdrsIESa5vGENHLsHlZcvhED0RF6MpvtxpQ
Sl8xQmKnJJ2/1RfbKldNgvXTBX+i49vJtyfb9I+xgHjIDKkxEiFJVhY1jhkdiOgPCa8OZvUGP1Df
Up8P+qoDeanB24PjFjL1AkOHaOgTqcZ1Re8E73XznUQP4EYoNTpkb4y1EnRue59RgtzGPuqQkZRq
DV8V9ohILvo0lby2YPRl9SfxBGapGSlOmDLZGlGIvO7kRpbuOCDC4OVaxfKyHQtzt/paYVo6TRjR
N6CuqVkaYcyRtMshOLeqg8KgqWt50Ec315QNwVvCJ/wN9iXAevbqCsuyudQraJpt0GlDMFIJVJb8
IIKDFZBbgFlownLfSVTUz3vtZYIKGcCSjYd93b7eK5pm8SgBain5bCu19pDW+UrZxRFA6d4d/Pm5
QkEB3w8ofKJV4zANlCRWtp2vDPicKTdJqpjnO01OJk+VEtaos8UJt9YAQpHH8oYikxa7FKD8mMoH
YPd7PH2ziB5hrAPYkzTFcJon37xLZ9b6D6k0NAOwm0F2dYraBTx1UZ8rrpEgEA1km9g/fzoM/pBc
O2mgLz4uIz2pA88h5BiwwabNUXFgi2fJqKDej5zxrZ9VlnD5icULr0VBqlKkRzx6lYcnM91FY57V
kDW0KCUf9xZ+SQJ7loMAwFxd+qqyWwZWYEyb24QWq1jhI2ciejDdbpTez7n64FHjU9mpA7cN1LZH
6CW9UsOCK61UzyQn43kaSWzkk7T0NrY6AbzrB1i9JOnoNeWNg/XXBvxDuRTdIo5yBtNZwefV4O4J
DZ9zwLvzGV8na419hGi0f2/CjieT02TpHFSpO4AxKAbMLdlCx2aM3FMZ5PXjnyJIhIu2lFGsnUXw
3zT+C+pnNm3jOcdVIdQwBrppkm9UpiINNnH09H7ViYWhv1QFs/8K8h144jQLXh0e+2/DVGQmoWNN
bG6WvAvYUORwS0UUyL7AVcz6OMtW4aAe+iouqNKPEUzo9epsCiREzbztbhadCyFc328S1g6xvib7
hM+qIxzBSKy467GxA/G+9pSFqILUx5/spDNemSyMGV0gOToYvR4eriKq6BUVAhHpnk9+fd14ZhdC
6vu3NzCnNpbbK3iiwFgrHX70OQyFfl2+o+pc9fa93OBGnrUSW6WzkcN1gTdtcjKfrr3d9tyzvQP5
fhrmp4vfQAgcVhovtlIT1NeD3eylQUILkfPrFa2s3e4kB4Ocpz1ZDymNdiWzH4eqWli0vR1MvgQC
d1KOt813wz28B6JLRLhefEsSvGMd+m97Z2L9KfwHcfEEd7FxJgZsGnW0GLd8KSFJ8jedaZYxKfzN
Zmo/MURlQmNrEiOvXtKsUcOA6aWiK24H0+Pt8i0SQIr3VCUY6n3E5sl7HvkPWVa73ld99+9lQN+u
30bZx8gLGyMez/babwFVpiMJW8qneq0MX6B2VXCo16whLe7NgvHA2Mbo6FgUQ7FsEOABY05YmYbF
3xGIgKsBwTMVTFVA+sRyQFw6qb59wQoofH4zYSRQvZ4EvIaq28ebX4VJDJvK7tBJR3JkIXKgAm1Q
DgvwfwgiuFSmlj1qQFFMKHc3LV4G0btmJQLtpqxi2+MyQbLSasmCkixK2oCjjd4I/AgUAITC67uG
3vHFtU15x9ygA0ZOm9EtrcHQdGW/pncU9/bA12V+PRGMRXzWCi6TSbArTIiF7A8ZIaEAkgF06uKY
JmkjYbPh6PKOEYJzSYsF5AnPirpoj3aiAjhUAfxcmuV6YiMI14YmH9WEEc7LkevRIAbDz4gqJ3eQ
8o1ucIOY2jlbK/jfAbRPQ4Jied7rdVSbHmstkJwR3IyQU7fY8tBlocKU8t+/F9z/aLI1pxcjpuRM
f9yz8ZptE6EDSAcYGzLvWs36+P6ZfnzTyuGe4IPrQ4DKxFdsVQgH8UsTWcK/QgpjGw4gowZz9P8h
rzWQoVdrzof7nhLn+2wEFfr5/j00FyKoRj754YUX9zoXUK+pS1JB64ol8nAtbqafOYOCxSB+ShIO
gTTw6IPOmW9zibXTtB6v4rxsW2HYtr7lByGhaMhQDJLX61RGbYG9F2TjkTYtUj5TrSiNpFp+7omk
ZLbNkIeCgxAdlptdXJwYlEkT0BKREhLcUotbGGOMLXo9afjT6gGujzugOLFjUoA+ylFo6JOyMT/I
2li3qF+gSjgvPE+NWEoNSMku0Ggeau9hYtReCL4aXZyxXI+s5On09ow1Jjs7JO1iUlW6arR0Uf+J
b3vMHVrtJ1qh8JsgYyheYVsDDSA6zghAEAEqVtEuKd9t2rmO6BcimaihddK3oPlJuqtA0F3+8Pah
Cvrv14/Mc5RymUP8baJPM9xIBgr0pG/ucTG5fwK7eIRre+CrPDZ7VkIeiVNHV7gue1OiMGSCdsED
Gb6AP+zHLkWuQw/t2bGr5z9mK8iKbtk81hhKYZAUdfp2KerSaZ+M4YhG03SCmwLbf1PvCapCsqUl
msgYd/LxRnluXzt/ndGou+75LUhVyTgqgh+acz4oGg5LjYbeL6SzgzL9PAx7irQds6nZRg6d+6kH
fsI0ioBlMn7b0uAW0FDpZzkYY9R3bPFnCAXNtlI07+76IRqXcM3LLbfTdmuzutcNqP+wcyHvYIJt
7o0FFvEar77I7/9ONj1OhRSpLF8ZbOkasWR/Wp6Wccem+7ZNZqoxnG2R3bP5+Eh6yPs7TNV20cuJ
ZHhl78/Q22ja8qtjaGfohv+ovuFCflTILyNR2d/WOz5kVMOgOSiCtrtk76XxmRJ7ek0QbbqdiDWy
WKmYDlEsG1E5n2uQIPP9+GXYbWgqcFHF6KElvj5FH9Szfr4MVizBeVIjprbO8k7jLOhe0lEZWZSk
XgP+eEcioqyXTj8Rvz414rrp/D232Bsm0pkwaMVE86Ysz/vI5DnHqXDrW8/FzLPfV/Nh8MmIKkIx
qkDquDWUXQ2MKfshl+gEKQeDoaQ3clVK9k1m1yekomDUASpkVZQ5GuWyiE7WoxcEM/CbcH7AGIfq
ZJSCy/duYbWDZwg235PQiWfOXMADAIwhI/h8DYtiOGiPgVcz9/2Q2FQh+PWS0zuBfZK2kJk6TbXt
4ikQrqXl59EyUAQJXjPPZSLJ+z4rUVnEKIJfr4GNqrjjFLOFDVtxWMYH7U7a1IxvKT/Em6Yuao22
j+LitAfl8TD1JdC+vEXu/GHfX/QIGsB7iNtKxfeRuh73zLN+XL2Gz0gINn1SlpTdITYdobrRNfaM
vZXFeYBnhp/tuheVNr1IK8rnWl1vXCAUpfyYhQNGJ6tZpB/nAZz7IZDEHhTxDvz0cEzLp6k/eKpF
yYMBKU3HUpSIb2JlQVjrlJ5GjLaPwQ1m67nU8QfC+4AQamRBOeDvv0B0JUpqo+j66t1y9ycdLZlr
p1f3HhxRpPS7g0YcTK2zr2tgHORSBbhzDDo4Kb4nQWVmEUpiwOX0eMpiyptvHMmTsisZCrzD0EZW
oBuuZbW5tygiWW5BpbYX/ryuYJaQusnq8K5dHetIQakaZCqGyElLW1s/Kt6oDR/aLsVLVhvVIWhi
PHmbtVcdlYpbPm9LNczzFJxgK7a1afFTzdVPcdRjh7ydZk8X682V9THmrVkpzN7TMDWMknRreI+A
UQiFvZpdNo6B9hJZdQhlO2n+ym5OluQI8YlLnINZju7uPaCdPNUijlyJEdEsZJbl6clAKXmae3kD
g3vk1yw9mDJb847LoxfsO3YIXJDmhj/XDMjDHRE8dfh1PzEYsUJkqppjEocdvcI2I2ipxphGC3Fs
gCxuOhm/b8XZLdKODzLxUedTVOQTOfvVhEu4M9t5WbfjevT+oC3WEv2F0TlC/FL6psLtT8RPnB/4
+K0csZUQSyqnW5Wlo5MZrQ30aM0t+EWrPLKBhCuMGFpSdKHsT8kuSWTl/PoLjgV9pJj0Kna0RFgI
dX9q9itp4JTiw8fJFtnnKmy5xPJfjElqwKN+QOted82d0wpuoriOz/LkLziYrUrdY3PFWjMz/CLl
N2oUg/NTITpEME94hLUC/2hA+HaKc+IsvuqtZKMCcif/K1YJ2ut5fQYvQuvVmqX+gUBuAU+crZzl
YTdKtaxTtOMn9ODm5aGqEbASu1ML91tWOjheJV8MtnOFlQdW1qGdIaZFKZCUitpaqEdLov14MqjH
9+YuUCg2G7jO9fnxs6UDZXcQg1eBA5KC//g/nr1T6KrPNI+RNN3NGs9x5coCitzlHSQ9ZRz23+0e
ai7PdySOTtRNOt9E6BympY8+Z7qymtfeHjQeKMU6ZEmYTjbJQp4WCbxxZpm3Ggp+vCkGirJTH484
vV0NiySC6V/c6IXB1+/uTsLk1bni/3OofwFdvHtjEDv0yzXf3IyXFNbPXYj1R4v8j9Y34+gso6Rz
BUe3yh5psHbgf391E5lSI1S/cuq4QMeCvGGNnSNf3gVtDkgGQQMcxVOeKgZqlkSwzlKi8l9Z0t+O
/l1WbkgM9jqWcHUH049kK1O1VTGdhXcynaRj+VUQPEwqm0zccAO8lsqwDSYxsjP/d0IXRK9NRQsz
1Wsl+AEIkEs2LmNHsIkF48xBVoAVFKG2mrzCFyD+9T/29oYYC9Z3XmLfCsO+9oMBmTdcQqsJotjJ
Z3QDCq+1J+i43gcq+j4P69Yn2w5g3p53I8se7R3EQ3j3kd/VmL1fD9Y5UCGSgXv7sIp95Ub5Oqx4
nNtcOU2TloEBujvtzILfMH5OHyCre0Y7KwJ56g/BDwCEbMCgLOyrzGyLcYaepHIxMU+qWVHaVmYA
/MMtq+J5eoqj3GuCBpk0H/aviKJOKtfpHPrnKD/fRzbYplH7xEnenSLy/C+u9Bn8mW1wh07EgVXg
uZIEGmRuP7pdKHSkHdaG+Qj0XS92fGqioYMguvl2laiCvpz6LyUB/KcZYZMFdS5voliP5pVW5pwE
RoXR/5nIw4WNW7vovVXrm2zlYamUCtHM9zwVUcxootIolcPx4CDEpYydzR4/aXbrXGmgv/gFns/F
oig/F7ZxW9vppte1aH35K5mgJU1JcF6Au7YmxzKwjyMpbIqfxP+on7ggqyBmY3xPSZjSiMoyoDoH
cagsHWdRkfdgBszrY6qpYQH9SASXGIHX2V9snYU1dWFc5e3hqCEXMpybHJhoelspxQO6O9xc92EM
vLs3pBDz1qUzKmhz1B6kf7+UIxg8KYNO0PTbhbXI5WUr3ieLt37AFm4wSaf8+X0yXfSEa0x0ebiJ
0xaSFWzIwUH68YmgtD6v7TZSBbG6jYX4+QtA3aqKpuv7N5Yzo3pTKfROhqVFtfPlaOFinmbebgyd
Pj4shRZ4U1JAhCAL1MHY3lqCa8xTWvEbYcLhjU5XmstWrrFdqdYUDqw4A0gNQBFf5ak/IWVJtjlu
1xxu/k1UTsuqz/waFqSTMbjZoXbuusHD7C455UwpOvTmul+Sy/068yzziRddy7bkNamdffoGvE+J
AhTKaMl+zzw51YTb8FEOjSRtJV56INpiQvrjDKl8DZEdihlIdGV5gC5vHUGGVJVwiPEkTgQTJcDZ
ckOuYHXs4f3iMFfT0Zjx+baAjMiERWnRLO51MyDv9lsDdWY77W7ZzLK//RPb3lKtXq6BQP499o3m
ysifJndDFPhEfrBRk5ScISn0pUkm5/xkuQVJThBzr7BXSFFU2Jbpxby0yC6z2WY1SZh2jV9vHW8t
O/1GnYoXi3uI9Q521WXKfMdytQvBiwhnZHSmUV305u3pqlzvY49zZpW8ZbQO+lcEa8KRVaj/F5T4
HC0snEEWgWBwMCSZ2i81altVjl10fzG9vRjaFCTkN1liVRV8em3dQaUj5aCH9gdSJoyet+/s3058
yU13T6lAykJQl1Avb959bCCK3Sx4Xy6iz2HW7xOT4LVSAvu5Qpi7PpiL2p47FLWQ3rI5sMFH0n9v
1y5FsVmayFMMmEKJ/akw2o5BmIW9hgb2hyw/eXJ8uBoaKw8NDt4j46JTYIW3YmtPS07184vKDOPP
G5dGyT1EkhudA9nQHGoTEdpd02E+fwTkVOTIZmSd8wnu5KykieDKpsxjtiB38tjTuhaCtoJE1utw
u2fvQITV9BI6YREXNEZ9UbaH0+mGwciA6gYOh0h/5jJd11jB3SyRFSHLzC45PYTtY8J0FRN9Bq6L
/WQSby4rr6f3h3h5rnk5UhtPb9ecXB84zqXlMGNipi7pJZAwQ/pzBEPt8RR3rjkM5P4L7/teVS9E
60o6XlfycmcZnBnnLAjQ9hNW8dV7o6nszRcW89tNt3Iuokb40EiUBI/WhCeaKFyomZudkkTF/4Gx
VY7I/IQt9juQgq+Ku0qCxBrL82lc55vhBbjIT1c5SfV7OO56CVB4M4vv7RKm4gh++qJ44uLpGPRt
9rN9bjSr2RIyH+5u8qZfGTN/qbxdOviK97L7k46BWG+jv4r6rMw7hgW+YER5oChtcPdH8Hqj/PPV
q2VF7yhK5xqLL7JryDet7+xiZxgMOwJzWj7XFPqqTk13nTJky30LY0JpKauLwBdX/xEglsnjKtNe
8zP/+lLOFpR+pkP1GL44n55Quq1+yx+C40QYd0ft5zKUHuhobbqmJj2Q3W4GiHIs57n0UmquSRpF
aXDIE++fGbNGM7oby0ybRixxCRLYvgbZRHwJ9FGKhbXMxEroDJ5cr7bFvIYMIWIEgtkdLuzpxim+
9V0DurD3h2DWS8YZ6x9JUpTTDNK059kmD2fHfrwzqowcdwcgQo+Zued+N6Q6RQxYRq+tbvRta+Qf
q9UIjuC3akKQ83DNL3/qDPbgFOFyK98EfVKpfaox+orjCwxiT50TcwAdHLruEVt8N9VeZBkr9BfY
O3mEo9GbdD+7UNC0SvKSUMNJro87AKcQvx/kOegsSobJ5bUoQwck0ZBSOD15HGKR2amC2pBVs6s5
8ZLTo9vKQE/GYRQzOXRw8mJWdtDYAFcC2lv8nFItGCijua8TkeB2xqsMam0SO1iERn2B/KArXm5L
4cmlCrW8Q3xvSi3xxZA14EFL0rnTZCB++5tDsJ5+GjmXa2fX8+xSNvznq50Q86rHTZbotwLBqbHJ
Ge7GDDorqsUBK2OIciJN3U2DtjJJXzGZ6qFUf4ubQQO7XhJh8gTzeifydtpuCJGAnS40oOAufTS4
5DUzuiVbOP2WOd8RDFiki8GR3p/RBqaCXEFnKAaYDZ0AevBN0JxSC2c1/ZfIOwc+4VNOj2xISV9j
Pnx/1+LQKVtu/pbhmpioi/VMSZFngOL9zl+jqS+LpsCcU4BJYwd+eCwsTwnTtuxaYdmKNTP1o9Qw
KnckEPhp1bO582GZrXNGefGYXAOCpCNIkrnRCB+gtflldDATXN4rmRFIc3wahocblV3xUKF8znru
FsUK1iR/idt2K52fqJq0jeu4fckH1wPM7OaIx2oaFK2H9ZE7HXLSIEQw7k/hoV5TVkFpX9QuJk3o
VZhVCF+8E5gdzLAfIi3kbnoE6EUnaAyFm5JbzfYCkzMREiE+78VVbm8wp/RclMkWRZ27jLZBT5zX
drNXyriKpJESLJA7OWW/2o3OSdB+UCHohU9oVp3SDN2UbW232wvDd/fC6fQGFG6JjrQSMM60n2Q+
2uYeQjwvErpBxkikAxeu1OY7ZPgb5E1AjkSs0z1ZjkJyq+xmoF61eDN2vgs6gVCltiWWjGWlTuI8
ByG6WPhRmqFalh6heFjYxPq6iBDLz4JX42tMwmqQ+hKkFkeXfxmOxGi5cu8j8ihQB2Rm48m4XUW9
5Jp4TSIcER6Ax/GtpdIev/qbqdQcYUt39mLdIGo1nXkRq5pRM+LU1eBij003qdc4gW8BlcAw9TAn
zbf0fRJREUQZezc0CIUn5Vm1l8UCt9YqtNN6v/2od0ttrV5DKV73ibsN4gGdfTRCq/KNmAM6v9kU
nHNHKkuCtSkJTtWAty6K721Isq8J8z3a4q1VAW9T5Xj4T4ow6G4O13nFmrAwvSz121IXALLpVON1
r2ei2SeRqP3o3PZDvEmFllojbYuUg3nc0DmXC3v4una1bMDfXQeZ8g5xNPN8yBtNUXsGwdDqpNCn
WZRFn0nnpmqEvgM49DHSBh6F1jMjtVp+LBdEEqj30ZabDxfeekqbBZCOXx6zOz3nUVeqUizI0bSc
E63mH4f/554GGCNvyaTmDQm+15PdMeUbJzohp9qrqT35hn619gfHkp4Q69mjhSnWk7LItst0mKSn
W9HRrPSiA/Jcwf3myAJTLIJVt4oqiyOeqB3P+xd1Gk7k5jC6D32Q9EwbWuStxGJY4KagB5PkfZn1
88vzvNDbVSkrzv//91gAJBKrNHYY9s8EkRz1j1uzhInt7SIsNrIxiv1DrPJ6pH+3V3Ck1uzTkQhR
mILRfEYDxVYoRLNf5QmJKQ9+spqYpNaqsKcAzrnc36i+rZ0SRfR9rlbM3sLEeBUCM7KmVlJiEN6I
sLo2HOgsKjC9drOF48MiPyT7QgH3Z/UQsCBq634G5Asjkez5ehzG37P908G0LfxFbtA/W1kd3Vhs
W1cFdx0K7ih9JioDs0zbSwDUPPtCIFyG6l67Oj2doMm7BFMkSJHqGqPWG7qqLnKeoZq46/hKjMW7
LgUsf1zsS7gg3429+7l+MFY4KaM6QY5VCL7Hy587oh81Mi2kl0aoNKlj7y35okPOY9vDmGW9rERA
UfmC5P1rQtcrP5UcGuJw9n9wSTnM/VqDzuiJFGupq5VlpXSjzY5mfbNFN9CSj11xRVdj6bjr1Ttd
s5+SH+cTDZN/uRyaMyw0DAnO71KSjGrDBTtTqKWEtxdm8rf8doH8Cf6jc4rULghlGlzbs5NQQYD2
zWlb5TMne/zH/agXbnDsUCAreh4x0ekbn7g8/uj9Gg4EUw7OURMSxQ03dmV5lWv+v9O8+3hhkh/d
6yH8nSiB+lcEa4Us5bcDKCCOf+lqOwpzBZaSySLz3LbcwNteaPUnyV1ShrP+KwUrskvM8EdB7nL5
UCWgfcHRyU1xd2KhbYsjubXe+FgxVmHQGRJzf7JrjXjFch3lrknBQszF/0OcPnYseO+aubHSFaE0
BDQS3GQp78dGu3ENCCLpt4SXFqQHN0TO/NxICjNiTnUlvwS6N7HLzCh3jlRzmyzRFoh4yVO3mw8O
9HZBZUtmbInOTb/U3HMpZ7dji72hNud+KGj5x58pmNAHR+l2tlpMiHc5GtFbJKEvH7X6eBKWNaWf
0iGglmJ+YS9lnoZhYcC7MHCLI3qCCkEt4Omh2GfOZjK8+g6j2jME6shP6z2BmbevcJCUBdOynjo0
Gsml4fvw4NViURREwpFCsXDtJNaENp/g001PhUqgBsRvyXVvmAw6D2jBql4AjgxoxwOwXDiEpwd2
WBH4K919yhLuk/aASdxkskCmUkVnZ8GvzxZ2ZWM5yFT4X6deuWwmiyAThJp4eukKU2EXV/xyIYTd
Q12VFtHlLmUSkvqD7evywepChK1AkT3kXdexc4xMPXEpx8upc3pAfoJm6lJYVqASqG8WZUB7eZ//
v2YUwRGchRh7d2l/ZTnTLCDjOK9uEIT3R4k1jl8s93gZ7eDyAYHGxQs2kXaMzGNjhJ8sWK1/atlK
GEh2eOU7u6ER1rb90RDIEmdcXbFYWZWY6pKgey8QdkxxT19awcE1zVjbTyU1qbNE8GZZHXqdS2iL
szvYq5UMFImnTkyZP2bpt9Ek6SmurnadiG9g4+8XNVDq6LznpCXBK3D7SWGo2nRt+4KmB+49Ddtf
3nwqFoorxynPmlQDsq4ac4Nq7Z8qIbT1noQ001vo8Z/yN9OSw9BEiYsKZUCIp0ahqj8I5zm0pwSN
0dMwPpNoJM5bcd2u6BTWgUOa61B1n7aMGSHTNfaXDdWPsN2ojuc2fyEXKeLCT5yPrJDlbTfGvwMQ
696s6gjJd48DYn/mdTyy1Y4RuksmPMSdnJ0CwDnLwQUkhrstdxcTJaTzd7yklN0QV0kAKIw+SHAz
uV3iGbtNQ04apC+I8fZ2/fMKK/CLZ2iB+1fXQTST7wNLvme5mChuubsxj0tpLXMUUyJGQYyv3QLa
GaZ/9spVjxXGsEA5OX+QbfHzG8edb2dWIaXkie6lna7yghUapNhhvIPQiUxc9MJOE3xySVADKAi2
QVnPR5fdELudWrkkqPamTfzuc3ljpnbr5y8xzSKy/h9FonUlXhkC9R9vr3Y9Z1Vdivl6mvYFoUZ4
egANcMT2OrpWgC/r7EnVajUFRZI+TKGs1HOCaUZCOF0HVSAIxRZpWegMPbMpVll1v9tV50PVoOt+
GxqbCUnsbiTTCHmNi3JgTlGa4MeH+/O7gMXllhT/xOx6WEwUARWwcx5yrZfG79o9pRjru+TWQAzg
TnYR732hT5mPksL1+TwJR09wrgwDJW4oQdfCsl0CpKvrkv30qfzSVIhh/pHjXaR6F2HcHC3yGmjQ
3AXnBO9JrofTaUkakctKWf8a7ovNK8lzYwUJZFOOoyFYElg9bwYltkLqyD3TWaulwyzcJHPjYmPD
8j+S5OaKnCRPczaiZeKczQMOYDnW2FUmpD/rKNQmY4lPstpxEigzTv84Qud6Em0ZyTlmZpr59w+a
lbqgrCxFIiTkesbvACzETbsvtwJSV2WOYnnv+ePac7a9zygR+I/HT5FpvZrY1/vZCPKOSuEOdU7b
YleuPJ72OAZyMiDssO4mZpxiorCGk9Y3piLaDjMLqIumAx7wFQhXM077NVaiBC5ru2D8FD7rDK0r
pO/bYFw+9//R5X/61mhGsNFw4TPuKuo1P+Of4rW9aDraG5BeeR+AsslM3Y5DLFcLHnHawMqQy/MF
DSkO6autVcCKyzizVIH7S2+rRhGNgdlE0+A7gAIYCvco+6RXlEHQmJKEYU4Z49ckx2PjhyAyzZ3e
59O/BkEhklJeA53XZC10wu+gXOaf3Zk7ARzEUvBQfP6DM6bmWda4VX9900Nr7BfH5fcX3eYb6aCE
J4G2JOzxgsp0157WUBBJMmG7UrYfGzSY0m3jjgl1GTqI9RTUBE3SnKROnU4JoSjGT08jh29uj4cP
TGNSTnKjyUUMrqd9XH3eTzsPYpVLz5w2yME+DMptiA39Fg3frSFHnYSB02C/Ub/VsyCVxA5cIJDU
zP5prHUCS33Tk9qQSFb3ffQOsMqTzQaDngJphm3h/Ki09A0i1U7Jk/O68EgcIqrasUVMyDczuysi
aSCRjzSXxkJw+nUvQhYWVRiQKy/26bG+sDIeCZXIKEOFy9UGgmMi+RBraDCNgLBkaBf15x/pRudB
X0gdWf2ktx9RlcqmWDSsR1NA5bhvWsrLaqt941tCotqpoRStxYA41XsNBi6Fo2qxLTAu5PpmYjNB
ENeqim29OjXD+MZZM6HEhj+9CWXpOrwSAmz2TVTRqaSJu6GJT9ggm291XqB0cxmRRdGMJ4M67/ZO
MXjzqDB4E9wxaZ0YoKxjWT8gKWPoytMT+tIq3NYrX7D2olaYbJI7U2mXJ+OnZz23pehJ1OTn0p8P
RM7as082gwBeJuQq6/PVGYVOGg3mWwUyPlXea+KlcgHIxbrDmHSPQONHDieTr3CbySu0/eU5QRUW
e2aYY2CyuSYg2LAmMEjC7Dka3PW3Ld1SgwmjbNXJ62vvLx4/rxl+rkFMbCH5AGgVD6DtUuk8NUHY
5CDsLgsax913k/afG2C7219ZV3Jp914tNhkZYSkKQlU6UZf9QS5P9EknOphTr+WiNPisrQN+niZK
hYKRrnSGj0riIqCS8AkBeq6GtM80NqK3gYSCZKjz7xN/1bXU9MqXl9tX+Pmd2G2EJ/TcCVCAsfov
WBjDeNH6pmj3Z2191UbW95u0NDasF6jgSgE/Q3OiHBrxSHoCzsTW/khYkMDMfJl6Em8zjOvaJ5ex
F3W2usci5ILnH7VOfdJPclfkKgIi5ulT3Z7tILabuVjYGbHpsiHz7coZpQQnphqUuDtyO13rIrdq
EZ8jMH43Xaz19udFx6Tyd4Z7HhWwxCcspu2897t4f46KeKIaHHHZ46YkLLcRski+lwW7oomIcQCK
HjU3Fy2ElQ6zFPwdXrhWvObZecy5k7DYyk/uGbvbHOi5OFbQxoPM9vFl/ounZhVwEQUBSQ8Mokdv
s9Esqr31rGbOsUQK3cyfpe0GmvSWc7TosjjzAZijHY00dgRcUBx2MpFQVjxs/pIKpEuKLIK34j55
qHj3UtkUtffieC9qRqlFyJ16XDBeHeP065jf9T+zqgRvt6PlAX3L2seiXhf5Evpf3Dmm0q9kVbOk
87tz0DdrIKBy6UzDRriwIQrfnw6bdzC9frKOtI6Q0NLCoRohYZzF7Bb/ZbC+lBjQdIfgu/cwxjRo
6zSuYuAajsETLP9FuIw7MM6OHEuuUSKU7xH3zFrNJJemBwith8mV8GQeM7u0rjXr7fJwvSH/Plm9
VfWI6AXZzt+XVAqmJvWJxGOIzkYVG31/Sq/LXBRdee9A1d6xI5tjK9Y89Izf0tpPnM/PeGkj+61+
Zhc3vfOAIyJ5o2S6qr/kkKdLUz84oaRd4ZoVr3HtIuSXuNuOQ3xK2eDmqG63w4G3QMwBrr5S7V4V
SCZTaJkq98G7WBA8w4zsD0h7qGBaCUcYQSvYh/mR9njpSyZelzj4BbhqVDmiBGhRdyzbWAElYmLk
SYkqCzCTdz8s9r2VekwiIwR5xypYO/qTKPu4Om9hbnyrJA3Q7ksMlHcGjrY+ss+LkmsZ2KVfzkSU
aaHmU0CpHyxBUAfi6aUDtQpm+hzFzb0HhGMoN2zV1c1NOPpEkdBIA0azmiXGX/nOBZ+j7cVcbY+F
MEU3L6dMglOFaeco1UCArCkvFkjkiXx9axRfey1SJSG9KH7XF6o6ZMzDEcR8ckHPfcpoJ6+qW6sk
n2LPLsx47cSL+gUnsZAJ5EyC7lLJX9L5ufO5dmjFAWOGg1QcPX/wzgmwjAENqMbPXeDY5BpPzaXl
lfOgCtVBnmAbDbZPDthY91BXnqsoIG6eDiMcNBd9BrHmLhCv9xSA/YzBRXecHjZCUQRDJFreygMe
Cq9i5GjhASbfIjvHZyp9COsqEFnLBdBg6LT4T5O8ZJyWeDs7xVhZ/pCyytY3NN5wY7NxXgzLeBIE
ab2/Pbx10swxbEsnkYzQjOHNqFmwILGmUimuJXQXfLA0bpYn2IwlyY+REwBctkJ/WyPTG757Q6X+
Z11htnx6aA9wdKuU6G1n57Ynu/leOFcNpaj3baWlcZ2+ZClCFMpK/4BnB6UcEkHg3ELIpRq1uZjv
FYE4H8Xkx7mvVOtRbNoiP9PMqUk/2JqjfRjo+RbRatbvKgLTFkTJnckmHtzlve9fViKo2zUg7H+v
52XuGv5b9+M6LxeStTcIoM8azBVoezjcuWoIPZ8+Bw1xBtq1IGi1pg31jPHzRrmMVpfUgLYUA4nr
ZtdYpRpkb4L0eA1EAwqTTEQVzjR2AtNTsN6MLGXc5grjsC9fJrmFgw489kTzJq/M2PIsB4c3w6Da
luBWdl3fOWrPLyKacWc/x2k6Prz1jtq5k2aSEqIg/BAw5OAiXyov2aEeANuh2GmGJjHScqX/8FkQ
oTGseDa0Wqcbw9icExvxS9bZIsOOlvjO6Dgvy84YVry1M0tn1yeLwb27hgLo7CZr4FSFKeNFmrMX
nDxajAkufaTldcN/g1pyUVF+4apHA4+ukcj2r78ZvZ/Th6TLPREF/7cAsIlCX2nnrpfe4jNcYdmn
0szTYn07x/baRpq9JK/fjcWKFbVzSus9bHctA66O/57Xe0CcsM13iQmamBrKBoi9EyG32kCoxL5C
xBKNN+kYeNmmGE/Qn5twaUTOOq7048V/Pgbtd/81IzGq+Fc5t3aRMbUhvSPY5EnuggFBsvjRgev+
X6fCBn5Yl4ZRIDYar5bk4xBo9wj37Blw9vvw5jK1ugURa8axBV5Dc0Dtl63hYmwI+7IEF6uz+B/l
QtsdwHxiKbJreiFVor9Ev5fDXWOLL51rBfUyadw3slQ1egIMFe3yGmr5+BSBpqs+IWIagG+lcTGU
EMDR5JMq7eoTNHRLbpxBuJPSp5HhG4VGZe5jYqIQ1RkahVeA6QG5TMv7D2VM+pxDn1mwghcQV0f0
cVOcMohdXgvcWEnrG9BRpEfJKKLg0tMSvo4jlXCJcv6ZpVpJ/2yaIDGhO2vyGe8Y/qpNs8S9Y1pG
lZEX+WlhN2rKfdwDXsX/5HhUmT2dqwq+jf5pUFfuaEzyWCxetXupWCkwDI+kKKM5S4E/TDrSVhg2
/1K2wQMjOk4LzNhe5bkPz2t1wgnwjO2elv4rVNKm+orCUlJ2SFR8D24WLOWqj96W8sxwfP4WThZ6
FVBT3fu6P1G0D/Nb2ejTNjKmLTnEkGQNVPwM+Cd6mXcj6oCr6ZaWYlnLhjx3bh9+09o8ndWJTaBs
DZ7XDF2ihU3dzo2P7DTbc7hPn8YO24WUgKkgcxLbdPPkMBPRnDD34DVyld4lbNlONgyzgMI5xQXS
NTleITShNGrskKB4AK42hm2fu3S0vjOrzbgHLE3cPkBhPOvqOukLmWz73VknilAqo6F33T6nyrW9
HxrBzfpjAeSAxn4M89OGVkUMNAAmZijA7z8k2DodsWjLCUeAVEAWraoD7CnhjwdIILHqC3GGprdJ
xzcFWo2GCfCkWrvj1dkMx0JrmdyyVDVdX311/dunaNYEA1ckA0winUgCgIesinfmfebhPbgl848x
9IjzEb4UjJx7ilzfoZE5Z1mfNJyWMesA5BxoWQLaeASu/W3EtwUJjYqZP8QNeU8MCMiLtbXZXMmu
Or6Xjb+DdYw32uTevJpH+vks56I6Do1HOMs0eGlQ+DGRDBEc5OXDu+gjYk1Jzfjnw7qPm+Pry6/J
8Wfl+9QbX9qLpWsTOIor5oTkWGUuzK59B+YWSpygWahtvtqKe1/KApLptoJrgBhPh27QtD+XxwQC
mxHc3Smy8Nx0PcteYTUIdNwow6NF+x6h3CN/gbf5vJi6tsKqozc3O1jk4heRdDnTSxQAnFCRfb34
/gkvlI/DqSHOnGAWnqG/fNAvaCGINILYksqBH3icKaVI59UoY3QdCNApQgrftImM2F7sqykbF44D
0Bmt0+6a/iW4V3MHerKE3Sdo8hR7XOAfzDw5zNF2Ta1cxr54AZ30Dlg6Au0ZKP5RuykdH8IxELyF
in9vnymy4bE9KT6ifnE+gFwmLGnJJY8tV8VbYcI000wEieHC8L5IVYsd+yUvU9GFTmx7GojmKJpn
XuCdyzxR13muwB/CNQ2r8sQb6NUMra1iKHXiaDH6NU4wZEiA5c0hsG2kY9R4Mgej5BVNLrIsddto
bj8x1AnDmkt0s4cxZnMKEdeyHDtO26gQiPPObrnhwS3Fi3mW5lkl1d2+52IHQIYXPAqxqZOf8Uno
/6yTucYoWvdu7wYdF8wI3amp7aM+XF64sxjtL3I3DT0rmyPHPTsKouxL0xuT0TEl9qsH8cEcciT0
7h7qSLe7RCr2QbuvH/Jphf8QFVDMT9tROd6th4BnMwHChn8wVLEXapyxMYHWDhMqZ43L67g/Zm4K
LUucbZPTBylwdOQ8ByIVP1eGJTyUR10WV5u4BmvIJeLa3Wq1Lr7Qg3+Gq8RTTWJh5C66D5DOBAzi
RGq5fYedGtNIVSItZRrqhxMj70uNQ0EBbTBHXkkDSChGwwKPIltPtY8uSqGuytJgU3gUb53YqCWn
CtOrcWK218H81EB3j6M8KJcM24ETvVIjEytF0krYuAee/62hMpzgCaXyc0L5oxsdHgmeFeRWJo/x
asYSnJ8bpXpNPr99xV+V4jn5R02yCggd0OTZ8M32d7bCY6lvEY3wa+vpNgXkcK3R3OmoVwmURiaE
7eydcIU2hlv9Diiszc3dmR00zcDfdeoZDC44HIfwqRdmmIiQwPwr191ao5Z2y08ltvNzKrhfFSCX
Kv9dnzDWviRNTJdOha3h3eFrJo0Y28FTfwjEvxI5GmzW48WKT2rhF9RJhfNKSI27yM9jsREh8FAy
oUpe2aKk/5CeG/1ZsCVOuMB7E7jiVkAImIf0HuZCDjzFL1PW0DM+W8iS3SR4/DINcD6BNIziVJzx
T1L1Jx0XX4fvJcgoncospzLUgTlwEkzyCCx4DuM75AxY0du1cvDbdtE3XPAvBteae3v91Qz2OgPb
2/pa/w3l9CA6Rj8+be2ovM6f2a4JdBk+8Mge80qFrw31c3LwHi9jPJClpd59sGx1DI9VXjqkQyx1
lF5X4imxAAURw/6QLjRp0z27ijDRqRiPdlL7vlqw+ZV/kH7IAWvuovb3PFOdJ4/NotIszbl2ud+a
46GKIvNQTf7OkzepurVjFF3e6TQLw3C4qGCkVRdnZE4m9N62EoLhIC/EYcsoPyk1yO+Jm4dGQCMI
9NUZDkZdqNBXbWY59f02LoZFfnh29cyTn/5LofIq4qF8SRU/W7IXLP+zzW8SC8Xxm/kIbppC3nvy
FibtqjJ3fMTyjv7YWPcPwtgsJNwrPsS24wnNgIjZZ8h0Tw1RinEIwxmPS9Y8MW/XEcP4Pt13/dCA
ttJP6OSFXBECV6G0Logf38RJ3//YOpnOr35QajWIK2bZc4x+AAc1Ov2zOuswtX4BmOyquFZoXZ/+
jHoIF/QnV/et9TxOmUxwOXGW3JZ8E1HkDc1u69ivOnH3hpC+lkhC3fThBbXhDzR8D6W0Aymmk0bl
yuHCZo8LqNRLDypK1PqknycaRdRyCtavArZJEak5kLrVdAs/iyxRmcNjAKgxJofCCSVjbIAiLmhL
cSr86ctfPrKJdocy6qYViy9XH5yUUlI01yK3V1NNBt72NVXR9uAtw7DXar4N7c8Jfy1OGfGGM6qX
T4wp72wyigl5Aryfha8jea+9Qxb+9gGI1UaQCslOqZ/zL8BpnckbFwydNQYNMLTy9iMP3VKKzMOJ
1U4s7f14Vf2r4CPL4xpv7XVqx1qvhlNSpoIQ0VKDAstMSUTjDX2VSZipzHDam245OZ88KMGZicVG
408L1jzfCqcpBHNpe7jhn15SYkYIf2prDV3iLcNsqNwxJw2SDfOvkKEZmXPnU+FDzCpH7bJp0sKC
nY06McwkKwhufCRHeHksJXGlQS06I/ZMFR5P1CtG/OTNd+DmII68pVIe9ZqhGQRETJQzfsOcbzQA
njT4NxlU6R5i2r82G1qBjfr1vSUjcjTaUJchpaNTHL95ilpIsjQpQTghVShkQQ9ZjhekJOKp+B+z
oMWHYnPyN+aINTy80ZZqeK9PwzKQphxp5JT911vD3uRghBavLPxhLpY+fMvtOfuoxEJfKMV4zscJ
gdhvTtoKN4IP2Slqf+xds6Q2WtEoFfdj/SI8myAEU5Zl58iud+cV528RFiUcf4CQ662NSTk1RnkV
oedC6QZKnUi2tJ4nYYreqH1Okv/HC/ss0FieGdr+OajQkh0U890YCve6zDaqWl1sukvM/I+/KhCa
p8y2ljA+bMTRl9aTAMjKBD4Nte0Dk2XhqjcjXrWFEZVQruz/6SGIuaJXpTbUiJSvUlGh2pYmcup9
ZI52kmhZT70kqLrKp4UH24x5JB1zRa0/YW43csTHmDiSHilNsnReLCTaWcufi7tXnrmC9Im75b/N
fl279z2vQo28J5Ac2RXqrFvdgVUQHQkJn05LCGvHBV4d+f/4bvlM36pCYPylDtETrLdWxtjOkFAP
FCnCvIscJqfaAI8+kjHVVpaZ7GuIAX97X7Rf9LciGXoRE/7VJ3DPBiOPAIyNSHPF62PCWtQF7XxA
boead42QUPRCZd1nmZcJx7cGKMWmsU748/T1WiYydUdfRiqH3vDLBrm83WRkimiQfA0UpWaJF8Ue
Xnfn4zYNbMt85RaaFbxqmut8Dc2WcDRxROqSGWRCcShkC7aFPvf5h1hwmvig2H4cE1pIStbRkXLj
BNKnqcQyw9s9UqExAUin+UHQ2KLxnuP5MTOG9i2kBe01Z47dClvjao1khjHyyVZn8iGngPHHiaYg
kbV1fZ7G9Z8m0eyAnDA48iy+47BQ5055zXDsVPDE8YytfjJSb1JPhkQYIhixNI9MPzpUIsQGSrGg
1dG2JavY1ejfAcphsTdUWUJIi2lEEbb7K4vCe34SVF0dMfOgNEMHW9/DbaeRjsaVqT10IhQzstcM
RkCwNUcXgZlVE3xYABGD+hacJ4HC9GbtY3chNrchEJkmjdYsEePbvQ2C2z5qWxWzqa1eRZdZPBlt
YEADbvFHHa9ugykFjhgMdvuOrS7o4qGoIo8gf5a4VkM5DVqeuwpvIcGe8fSbt2AdDH8Y5nhshbWI
L2WIhmBxj5vIl35GT9lhvdyGNYmmGTuoogjCHpUiqvYtURVXho1WuJm9MWveBM/IZZNOjTyt08kX
Z8toKlymctPSPPRfToegBTpslmKrLEeuQ0x+8qyduTKFyqPYtSpsZf18kPOM84qsmnekZA9UEnLm
zAeNIrfm2KkfpYPzRQSRcrSaeru0G9fjTc5LZU7juBoMO1iQcigE/FBl0g5fScEib8raksw0GpuP
Iw7j6fgEoJ7oHVuabJKyG3LSygulOqxBx/hMFu4ptrqlGl5uWnNVpsngv1Jne2YKEMHWIrtw4tLO
yJ2wQV3NalUhHLjVlCb1w7cG1gp782Iy3RPkouHjGcuuDo2+N0qarqRE5EopIndXmkArsoi1njcI
1sBqRA4I0cLYfiF4u6ia4EruSyIdAkk4Zlbxt8lys3+Fin14CrJKbohBdvqidtwhuFa3lZ7DYXKE
SljO0574S43I114f8iyYEgGAVq0HtG1zN4g+Gc/ttWW9S33Sb07W5Ym3ikTQx2NMXr88zF56bXiR
0IXwuNa5jLsOi1iqaI5GaGiuzuky//ibvJXUtwlfk+5i2V4wA3GCxesffKlY2fB8U7IY3P4Itl7y
NXve6mQXNtiv+vG8lOHyT73Bq1WoL6qn21zePjmpSYk8zsdlK65GjkpEQQJXMquPSQd0xX5u+r/f
1ek6kIZJ17DnfvYgUm1QIIQZN/fNtc/50UUX0ePx+wQ4V3AriMLKxFtlMHfBPsm+S3wA/nVaZwet
IvHx57k+oMMOBv1FNOeoAhEaaLe+adYo9lCmKC56WOCH9LWvaNJZadzQvwh98yTZi5tUSSEa+gf/
Yvmn4UeC0rh02uHmQwdFlrIrXxdnX/WeUPtQk4CPzra79Ww4Avigj92EYphYEsvsI8aevekrBO5D
LkMhhyg0Xr1AaFItDFRSAB8eeTw8V7kIuIAN747nTej08nLvosJ2ls90Bi+0RhCO6Mgy5+83gK0z
MPCyQbXyEKsuRGeRfRYG6hi9ZhBoLBKatHNnLr+mzA7T0brvdbQmDVn4lucptiJIFRVsOmrmp2pb
5ot4bm0vo5IZnbNVbhSnoruIKIdHK2NfuDa5de4PjgXYCIuIPtoYRtMQOgiWwCHShWcIAeNeCNCS
yBGA+f91Uc65xfTD7FNk3PbdFLId4GdKO/1b3ONuLhSjt6yTYzwhyNfAGGQN3oJCRrfs/fccL2TK
oOOO6CjS457s2Ky+akPkbeG6Tgs71aCstJNjXROJh8fdWrkFQvjk9wykSjYBgwEwONzhEtGy7FWT
J3CmnwUCGs9dgiZ+YHqlMBIyMdEbKjMvCPrAVTlqnGLJHSRIpma8SmgWEPU2Xvq/hUurRyoKKLCS
6NiwSiXaG8LGmauWWqFHTIoGnzZtT4Z7Z2F6azJJKf3j8wkGkdkw0Ijhrf0kBd5Fgl8TkgK2KFEI
zvwSrOKS7D0lTPk3V13K9EfQajfra7Xc7Q1ZNuSM9hMrIp2tci5gV8Qwdd+gzbusbxxbxi5hiP66
tCcjZaWQFzleDzExNdtU8xNh70gUps1cnDMWjhKRragvBBfc6AUHiwo/VnODERGZA8Td2DU2QZdm
p1ZMDwjr0y4hcKM0pBWO63v9R1G3qx3E+etlH3CpugMruBT6/D6SFFQZ6rTdHi7ivleMXpR2j5+u
8F3P2xETOgOZxfTMSPOxjm26rnrgNJpmcVMlTn3MNenqLobKbtlKUvyUakK/anl+q2+Gp0AFMq9M
l+1Y2h+3q+zo4Glj2ONF0eeIt3gxQGdODFqMx6OBW20YNZnq85ALnnUGNeJ+p0tKqj6tm3fT21ou
wA0X6wGn6+jJ+1YJXe4yyB22yNbtwd4vxS9k/fzeV5E37fQgrl8oFJHW3eFG1a9puyHF0s9Sre0M
j0cAzM6htiaYDdjLnBsY/yZz8hzfx0o+aW0SqP3e3aUEHgnlRUj5l2hzXntLA71gWtuxD9BLFMVU
j6Ehg3K6NVkQ95Htn2D2/wPaeiN7Pj6lLniOIh9KEB81Lm28aZOubG6hQaYwUqexpObLcHUL2AuJ
cpQDBbIcGTiyOWqGKTrUwlJCyuPn27O2h4b70Fu0a+LvafBGb81XeYLWshqUH1O0pYOY/kVq3/0f
ghvmknT+4FOXa1B6+BxYKPin8Z/x8nCP90xdFanqNLRj414BPCdGkxqouw21wG/3ZepQ6l2GVXF8
gmti/wBmUVURhgmlr2DkXT/Nzt2Azjz1cybjyzS22wlab4EUNNRX/mPT9h4M2y4I1iOZaJaYjNLy
bRsD7h/kkup3W7UkgqkHw+kVvPSpcyx5c2Qd6efrLMXzQbK0ATXA87jNC57NwrjIJU+aTvGX1tXf
2y0jAGoKIBM8bnYKiyG6FTdsu7YZ9razv85CgdG0Q60oLNp4nuMzwn6kAvw5Tfr8lWS/w+mXi9Ci
ctAGZpjRgXR5QyZACGIZy3gz6DEYuXu5IC3MAxQRTAwuBZeH3vSacREv+SbDimzvCO5TGhCZVDjh
rYJeaPn8CRmryYJ4UeAzFnfS6vwpbap1MupT7VR9L5tz8jyMXUrPcT5dGsf6655Pmen8oWCdMhiY
DrC8Qn40yX7MEEVq0nECLaF4kl5RGzps0CjYfy8ixqoV+9YLdTKzLzY+7hwDV70hEVctjYUAT+J+
wfX3VzgpigSgiQV2eE1QagA2wvAVZw8NdavcK07e+pZLWfLABpmxoB28NT4GGHVC84f7W2kXKMNF
UnnmGjeK9smn9x8kpL3L8vQBfQkbuQc4nhexx6O3dxaRBiNnHuPrewtHh28aVkBCyTL1Bn3PvMwS
13UD8L+lWu2EJvwDZ9q5Xkq70uxzSrwQG9KQ7QqnaJJcOoHYcn6MkUUhOhYzFCpSSa8cWmDgQoov
LFoThUh5MoUNMHgDytGvPKMXEb4J/pgbpPHiuns+A3XubYGiBLzYB4+3ofxn7CoHMb/6c9jc/eX4
e2xyOi9AF+w3sUqKYOHepy7ua4lhPBtY3XC6lgoMSvjxWgT7aSO6pFAN8waogyZ2dn43O8/nZqnJ
Iz7BhPYfga97fK9oBj8qBQ1Qnjar8K/eHDsuBh6O9G8vd6U50iOmOz9WeNckIbVtFSQ60GFAvkNb
wL8EfjL3Q596bkYbzXX2p2R1DqHBTJ9sy98YuGDX3el4XomkYJWNFrfaDdLI3ySYW2QDI+XRIE2p
czZGsYki8lUpg7YvQnin6waaGnYjjw1v88PmZB0vDYQaWOxnM1Nb7IMijrzQXIyB4IJ7FCAOdqZf
75St03weSRL/8IZ0yDYigOvnCIEDlCEC634sr8FzldimnppdiXBeqreJNuyRuhZpf4xfog7zIdeF
f9uPu7lq+JfxPVnr79+NOC4Ax3rIg5Wm4PzeW6o7FDuDZad1M9ngN3ZSlTZL8AGnjjYGWymvxzWl
Jer1qcNhtF/WMfvuAKtFA9aM7HWZGQKE1NqGk6etn+TNnoGD+/q7gF4qphe7V6uwoubH6+4oWwp4
GHjwHfwGFoJr9l1qi+X3OQXICIwZIlAynqFN12e1GF+BdyVZUsH160QDoEik3vsaeJoAtB5brFMq
YSZl2lyxLF9sfEnUy2guL9YF/kP9batZkysPrmjuYKMJ5tAoBuCVZhCM1ZL/+Y2hBKtL7YwPNxkf
1sXRJyyJ+jCQ/Gbhi6nWYNKKrXUAB2LsNQvKU4pylGFaNq4Fr4FkPL/koflFRoYVBfr95Z/Br/l3
11bqwVdXDyfUqU5nvjAEaSuTRT+FygB+gfll0Gp/0jz3J/pGdiYPi8q7qka/itwy1Q9EOJfnTZ5/
AHDzopSVu7z72teGKiZ7yGILEYuf61P1p7rBtgrk9Rt2KZMd+GivN1cA5jkpu0e1buFY86VHMcoj
7kwFICXfu6JR1W7oBKNnkIe9CJtp9ObbQgit9oqSMak/7WZWhYImasn1FSfwWqzReqviWb/4DNkH
lLMq/j/bLSXtAQFJKA5oGO0z24Ig9SSELnGBpXr+kfEc/AWDBK9MUWR22C2+3N6fQEq/qK92M8Pf
tYQ4ykn54eUXR50PJMr4wZi4rEbm3RLkDbcNRTqkdW6UvZqCPO1m/Px3B+dm+nMV8I8LoSX8RwBe
cnnikVHPH0cnA7+kAqrwVR+2XDq7bKNge6zfkYGpnLXFaJZm+6mj8UG50Z0xfev/VdXTjjvbQ6Qt
D45hf0biE+Iv3yQ09IAV+eC/26ZAiPIljTmIXRo74yLGgJ71eqbbZVGrwGUb1ZxKCOSCRNrzeHVy
BqzGpEJmBXwkGwIDh6X3USFRRFXp5uiFiizfDQWk9pfUzvxKFyVN1qZ/HULnNuWSLiCAeJYfPoM9
Eni8hwFCNuU3eWv3bpLpGQeAijyqSrx7lx7mbEbwc2h6SpGhUaWi+kjIcWaTsNnZ+ogECJ7Se27j
gFGbHLkZ6PTEimpuxmhQq2zNc8TFWYZYwUrlc56cbonIZvqPJJ6tIdCCV4kP+tUAttxDEIUYg5lx
VogvBsVDLMSVCgY9pOXftelomhBKpaH5HEykNhsYNqr11aO+PXfMtXVGgkVqR2vPEJHuqb9Fe/Tr
Elb3N2BmksWNVQGs3f2eBlFcfP1HEy9bKYUGFQDcUkt85//8LydISfhM/UEbVSdFR3zF/LU3YUcm
57wxqnZz5oTIQO9sqlELLDyobCozrH5d+MuUf7rVYk2F2fK0W8RThXv4s9Al6rNSG1y6XLPpldMj
NV5QVij3uJGplGB0n694DEp5vUggXJZ6GB9x3jj4MXVHXzNh9An0CLGKjH94LqeKxee3eFb/zWw/
tq3N35Pa/JBItX3C4mnh+e1avhmwD2t+3d4qcj7uP1R1l60Fc24VBO+e2P4Vsaw4dy7hOSlNX+Xl
Vgtctr5aqIjMsLc1RHTnjkIbIfFZubs/D2Wmut6VRZOLOaQ2PA6dUZ6eM8WqC+PCD8UALtnGV1dy
woz2mmmb0pKfxCxquwEnxZkocnrVBmN7r05cQTuZ3u0jRiwW8pKbRVQtPiloGzj1cxAiV/i5AToz
jUA+/Q3gZEq0adRwGzOZ0DFA9O32J3IWBTtjk01F+XCESRSPjTov7ZCf1abqNlozLHt1oSOfrrT7
ZUDeJB73mraK110o194ngf/kJg5IX9XoYAQF3YQnv44+J3vkRzP+Ov19qrB6PtmdDjduaWu9mUCv
JzPPlisyWfudlmX1ERp24fKZRnm2nuBfpwBrKJiBUk1ibiU10zU5LuGbCvlCF5j8deHBoAAcjgc9
gi3u28vb28oRX1xYgF2kGGHZ+pLBlJFBC/WKb8op69MY2OywaSfPohDVf5v2MGaRuxz8iyFLFOGX
gTkFT7J1ynAl328drXTRZQcy2IZ+Xa0AuYfbVXLtFsv5642roU1mu8aiR3nZZG8nWnqm4ljjVDVL
u5AlNbEnKu4TnHF28wJwTWQS9sc8Qt3tb5BWLuV/S9TlOHVFD5s/dSCHUcjHOElyXT5jRDIFq+Tg
AYP1ZTzBqmIpiRotwq4GmETgM07kW+uAk08vQynYnyCD7658qK+y5zRQjrxAKr5qB3dJetDi8TjD
UA5XSmWcZDWhq7iiK0ceYshp6ZhP+QMz2lBHtoDapQQDx3L1F+wO2UCuvDS0XliWeAJ2VAXctpfj
VTU53y+mw+dPjOLiLjCJ8DRIPWHkfVc4u0nm61mxlajekZmJBK40jFWHgQLrbLFcMqrGdFXF6esx
ftF2wVV9K+mCvqUpF/Y1jIod5aL+NvmqZjGC4KMstb1pPR6OeZzJWOy/EpEFnSmW4L9YTCLgZSMz
h8dbBhkYOO/OVPFkBGLAIxSkZ4nRlNqTS6earr5xmDWLAxam6O4zTICthwGuH3gkWmZ8kb5Xbjtv
uWE+E1vtazNQ8KrfVGl8hDroXmNO3r+QTz8x8VrN0UCE2kUn6ARj4ERjqaFS5aJRB5TnpiUsUjmf
OJju2GfC7U/XiwSF5tyubUoqzxprQcGe7PAkwMug0GBWA/ulUA7czlO+IzxO+rMVOJiUl2lQV+S9
FGbpFQH1zpPBtRcJsctAtP/QE05QeR7JEcgLx6td09dyuk3xddZ+dR3ISVt+BlkN0yyBFCwXBsJP
qp4KPUbjyKOqT87mD30nCodegP4LlHX3JU3nMwpWkijV8UDqEJbnTi/+We5KEO+jA3xVzlXCMY1o
ieowM/q8Y6NJt04oJhSSVCBrq7udKv3CrQ/nPKPge+uHmrZuYDLKywiYdWzkFY2pbVC9EAmpI3Lo
GoTMvyFRZ6UECPj+Dcwol7DVkWiMrnKUuaTMQjNWPLSJ79GiXrkpb6HYJ5qT5/pKYWDpBN9QX2qG
LICoQjFbJSk5tRiOZc/TluXzOqLyNp3eVskAQWnt0D+sRdY49CO06nTXE2B/R2JO3OThoOKFCrpP
7wI8bU+u8541n9/DKXpPBk+ffAmUM1HEAb62SSUObpngSVlfwHC7iMLhBpUdhfZTAVOX4yeShpQA
mcALl0u2Rnh4oebUnvfZZLgkmkPHaw+HXF0ZQXX00Z1fhF8OCD5dH2FM7xJVCDoRYW/TmRpCjDiL
zsl0LbCiJLqaReqGDFF+PwmFA0b1htGWz1Cs7BUUnI5VKcVKrS3ZVYMrjDdMGrI+P3RmfqhtpiEi
EXwc8K2afwJ/32yBLlxYpHoc6Up6aOTtZrYI07t2dd5vCihYjuyIrebD0Em0Mgr6jgswo0tDVAPK
JEtobWQ/oKQh4dySlgVVjRMg/ZI3jEgZ0dO+khZimXr+ZXZFd6ZnDgfnLBa7jKF3E8rREEx/liCU
FDx0qL6r3TcWcb58skhK/cF9JIdxcstN10q7uZeZ/YtCzTT/IWmWtt6XeO9Np61lTgGvSd7ZpSyB
kvRXxRJxWRSRIMvEP7MQ6gXAdjUwroC6cLEaahTAFmJe0hHHvFZiYV+GF5jZxZSJSoGaY0WtLyXl
Lf1pEhtkvWo/oRNvbROUxUvgVoQNlG7wG0TWvyeHcl6Y9kQJZ7v5pZ1b2wSC3mckWKnnXSv11eR1
Tvq2ojPcalpOlAYOQV+0+W8eCAY4XzjFO+fFYGYAVy7yToigAcF8CQT0b3TMzuCIzzGUu6r9jRlW
CYS7eUNpcnqOM2nfKGXwFIVSmpdtJH0bWm4hqJnVv0QTop85/0TMDfStYRgPgrDqNH/D2zxb298v
Lw2VYufv5yYQap//i9Z42UkMd7mPtiflaY8xBVrfr95LgDUuPdK/kyo0A65UtIA9rPjl2A/NIV54
ECqjnSEHFnm14iI8eqTpKBpKdfIxtOuqUv9TMKfmu+KbkoPCQp6HuyKmJ2tnb91xyw5jrmXTX2ZL
E80cxWuY4fhrH9J8h9h9Irfs/utdmO4eU47UU9acim1m3SbSjreJJ/lgvclZaBhipzetGDz+GLEj
ieePY9v2IGPKTjmvYf5phO2mvFS9SzDTfI+DMoVfJt4chV8OKvKWrPvffmmlQj8DGwR2Jr2bCWU+
wrEIp3fnuIHaAzESVNaF6YegjQjh0tMVcfXsIPMhvuVFricC6AFXc03MeT4CP/7MuubQXVy7iSwW
se/g/c+ejBDfGKFgGGpYu3n8uXsLAs+RSDKKLmDZTzf5N8ldFOnsLokCNTjOx5wJnCjv/xmlZwwy
DTC8tdNAVCBCY6kdIDKx8imWZz/IJ29938tIAmOiG0XspFNX21aKWnmQQsmQDvdGDw8p3cfHhcr+
5JJoo7pWJh0ZxdlL8ZswbissWTEpUFRK/ulR6NZUHbh6bHkpa7K015FLVauOfJ6JXBtuZJQHWara
rCirmBoTlZMJ/UuZHfFeHDSkL3Sfu7C1aDoXcHPtArtY92D2nPqZp+rwd3cPSY8fTJguCFaCPWsf
sqQUqAlQ/FvDpVF0DnvfH/6ZFM+wgvDD5pKOqveZYvU+K6pd1PEyAD9z/inLjXXN2lzX3rNf4MBi
BDtK7zszyn/vP0sICrlOc4OEwHBNSQkki5lDE9nJOM6a+K2uBjO1b+KOdOnQ7pdrzg9INY5Htumk
gBijUfMEUnwhxR9xHI9HJoM2A8bD++smYWIMau+IjteodXntiyxHaNHuQZgh46K3zyTJnE2u1uQM
NfIRBCNX3q++2GruNPFXRdoa3pnVpdiiyFzuC8E6IE+SC586G/KhMIsZz4rHD5o3/MlLgvN+URr6
Iyo2NarSQGEfecmmORtJ8Jdoz0FNtroFAFQMz9ooseWfrlz0Je0Fh38XBqMhF34AcXvGCf5s0S11
xvpZRHkNvtNvyB+j33qJ1wEVZGIAd1R2QX95WvxIzZeI2r74oorQi3f2PwMeqYbG6tn7EwFJIlWY
mL7ekOCLHTE5venrdkZMf0CkWxlAlYuuhhMmsgaPCjNIqPOmiquaRqd8FRV2wYAexlPs/UB9yCl6
lBQhaaHiuBYUANuhj74p1tP3GXneZ2Ve1ZotS0svraicLUUfBGUCDppHIMrkgALGCw5U/Mm5Inr5
KEvDomd54FXpqWouz7CNfC62/PLT0HvDf8pHJyjpFIPBAKz0eAdlnnn28T1vq343YjdT6d2ehQc2
xp5imteTzYY+dBg6B8ep8DvNy7G1F2Jljy7Ev/PwnNx84Tiv3eWgT+Nifl/PYqlbWao3kLIyzi1f
RzwsaJOEJqkQvBnCL+GR3efRZ9zAUEu/5flQ9il85n/RitTjFKrjRNqH3+Wo/BiW7qG085B+FHDq
MxPfrN0lFPGEurIvP1h8Or0F4Pl81eifG/QpLunRIYBsNE39KoVMbqoMw6JNMDJP3WpgHnB7fr3x
lRDElomdXABgbX8kK2oKsZ8haDD6ywbtMZB3wHmbJcdvX4rWoBh502Nm3ZKz4U/uyhCLBzEsa1s7
aQ17ODaevEae17G6OlzDdlJsYm8gYzxzpxIHP0JIEsvUHm0dusKHqnIbHn768hlVVy/8Dq4spiKg
mU2PDpRzhZmyzFiG/9bpWzut5SvvfOHL8hp/Lx0qoiqGUHA574maCD63Ieon0VCx80ioydV3wFVm
pVVddDFn2P9CrJHuaWrBd29GBH/8RjYcftczrEO2xiYX+G0UDIfd03i6RriyR6W5xpkV1+BNp8c8
7ffFAR+P0XnvjIarYTt6sN6Mz5S1NbC2O9SQ9mCSAIVVhc2guw8X0FkT2WY7etCuausqqso8hL7A
MnR9fBNtiNo5BJil3RQ5q6NesYrVFDZjHx7YN3jezHXJ3vxMAt5L6qTuPtxhpt3YkpFwLZpztYXD
7E3jaCeLfrejEidaQhireKwu7o5qet7eIgSxmzAdF/WGIDSXvhUHR08l3PlRtESVfgg4WxVFEIA1
jlrRKMq70qZFxscpo7RjhOUsKkysRNVC5Fx19ey2OCk8gYEzE+49h/1IVlBdFCs0xbe23EoI07vq
1lt3RSgfXXJ3dRSJtsCOmJDv7N0fn6lAVRPmqL5Hw/X0hzm2cY0K4+cAty4YOME/tTOaXN7g92g1
wpzQAZVPY2dTnccFI+ZcAho9/xDuL9EZlVgs29LEpBgt2KuCwovK4pqi4flp/XLpwT+Id9QySoJp
IKRCFHxNYLDYUEWwiawkvRjXmsk+fsWpzfpR9IZUDYQJS4bLBp+/F0u892HwfBCWbrUe3b6cRJRX
UkmNUV2ZsW5eSe9P9YgOKxu4R/+GXXe6GSHHd24BBDEkuF4B4HfLDupplylE6fuWSnp+XBuGkhxT
R+QMQHbdi+0/ZyUjrGp/YQBZHXeeU7HqygnAnG9gv3Vj2gkv4PtKP1vfgIkS8m0LEmVBjWRhn1Rd
x2GECCTb2kjNPNRR5dnUujsekqV4fXIv1kfZPqmZecjZ0CPzuz0uliVN8Pbb2JiJkrd0nUVA/42j
XCxWyraFPAjNO7VCa6eFo+SqPpMubT+/rWoVIh+u8DeVUCjt4CmDKYsC38f2LwoEc8TlyJ6A3via
Aj8IzBQBJ5MKtOAbDI57R+WOnYkanHCBgpqZwRIygWtO9GX4HxwFwg81Gtnlgi6bXScMx0av6zIa
y2wgVrv0AXyyBCEri7yuaSkFgEg5DvztkQZE8sP2OyB5KuHvIk2L0HKaQKp6cOrV3Swemg4017PE
xck1DNOrkrWvIUektidTRNlns4ShyD9+ernT6T7X0g53uafje9xhSXNuOf8TtEZWU6O39RTUdknq
lPWCN9h2YGrg9KWbdIisuJIVEdp1EMOaCl9+9aYPlKyjWzf8NbQrm2rUXBy2Ej93NEeEh3AvFNoT
F3eiSatNgOJbhSwpvXQG0DJFPSKw2rhuWKOMXdpC7zCI5F7nUJvxDH1EGqb0FP7TC2vv19l0/Wb7
0s3Li28EbRf3M9jtSyPyGZfz9eLwYtfdzWwfCYUajnqAeCfoy3/cL0RXCIz8YtDidHqjRpNNiYxU
+MruchduUjObaehhJYqB3OkvgAgwaK7DFsniSxLRUE9rkUkOtS2Z8ukaZYAt9+J5krx4yITbsSTC
13TX6hZPnBeTXtlNtk76HTJrjgFqMVNIGL0TrR5fY4LCqetEXILWcpLve7JWuN+b7Z57IegVld1K
8M5UmRvPXrIjB73ro2+3zFMlr5B03NQH1brIkQWv0EPtI74e+1z59AILTqJi1efFCdtTqfBWyzV9
uIwZx1f6myEs3OE0fRnPk6ZV40t90Dujo97qNpekG8KSXNkzhsawMDRFA7RuEikKUBLJLKpgBwTs
Qfg/eCAyLYlp1aZRXHmcEAnH/2ojsRAH4/SnhfPX8OSHnKtyWY7nzs0esP3TJipVK94oTp2slUJQ
xn7ngOP/toCNLFWHYWmacn6QD+aTmrmv/MDseK2MKdUfr56CEwOEHWNvaVKdF9z1OlxHdcfqs76b
m2pVZBI2QyaDh+jrFjrc/mlwio2Wcr3w2S7+cVcRCxETM77/ko8H3QzdDwdPW+yeUiDDPYM3uSgr
vNu8+GJ6Koozil5SGh/qQSPcvXTo0l7qK3KZUFyhQpNnJV4NjQWJz7nyb1C0tckzKvcLw7l9YpHY
AsBne7M+2Uvq/HDWtVTCOSkktmb7OPeKgfygU1+ZCKp1/9vPfzpJZ5sW3JQQQ9MS/fTInVKZaL1v
gYFi7fb5tU7/CEXSNQyAZiGVqVFmR7rdLgxWrGobjSYRtllpDHBxCbKZimljad0+RdvNjCVjxoIL
mnKx01T+ftPr/EGHCAgIoPJmQ2cQVHy1mmdFpRcNjZVg8i3fwZ0Po1kqjLIz14JjvuhTgmGm1BKS
kbbiGP5bbDpbOPx9lXz/9tfi6bmmtbwtRQBEGDCEc1i8oh3fPGIpb/RsGpsc01F2xOoKIbf9Hl5A
zQUib4ZIc/fxzGiydRKxwJjrkRLWx7pXC2UpPL9pOTuqcpVaa25h2iy8IUS2jC0Bo5wUeOCHFK4u
KEt4LaQajTBc1Doomz0xaEpFqNdE4btsdJaHTD1Nk2iAfeEWidxVKDoQfCTbGQKVFimNqqxn+UYF
eQriQ9LOqoWhY9/Q1v7WXmCMTFLrYl+Qalg8cJ96v4yjeATkhCDauxgut6cgFc/NTA/ola68ywmY
w2Fd+4ZkgeuTboqnz4Wo/viWzznwgVKkiqxtYmBNQjiPWKbqqghruodeQ8UbbgtWIRo7D0O56AW7
TbzAk1IkYOeo3yN+VmdR8D7baVKeoQ4UXBSgHx4nHnIsiaIT00UVWNaxmDqHq75OVRWZ5sk9Ch7s
SIJVX3TDx5FO/VR52nbfpLowcPSJW+pVCl/ndHk7A6p2ia+Gfu173oHbTTXN+i1RxVA+cqDXdRH/
7yfy7nH/E1ox9wanjT44N2NTD1ERctJIXDCNY9qEXC7WSbRHQk3INnJspX7vUn9JnqiZ98a79BmH
U8Jz+olCjEIEMZyNVeZUayzc2XK94O/yaGtTIbWf7vOHKNphZrEzxB9DWpFu1g7KvD1cpXhJ7fpr
bmmoExcaGk+fCON7kdetOgiogZux06e53Fo3Ma4/2mhPfV21KFQmou14TkhJunHABi+6ymfPa+80
tAz3YhakEuoNJ63LMVE25/N+pCnwDh9ZG1ndkihHNQPXqBu7kLar6eUkee8NKCtqhL8LM2yvdFza
mRY5Qq2vP9kO68Bt1wf9bTLzFOWd3Gw7frATmwbYJdLlV3ggpXmSKcRlJcfDvMby4751HxaxhQbU
4VgZX2PHyIglHbsR3OLkpjhPS+i0z32g5bw37rubSh8cdNcCIy/uT5DOT2Cmm6FZwZvIXImwqROG
jzoE0kLRzuPZAH5S7L4f2hHNRaKE0Km11regh5JLTwXr1ROQldnXjciVgHvBPmb/xXodFcmKIoIk
xAHXxDKvitb94bF9AznR16KxL58fdxTV93RSf/JvktcqUVk7lsj7XRSlLw6C+pGnwbhHVGrsgbnV
yC3Kz1iOuRziLIsWJcbLF8tgCvQqA6oZPiby9RM8BpA5gMj7Kce4scrRMeObmUa2vkAAXZ56mqS4
er4HFzflDwdPdu7F6MNTZUVb6xu36k2WVwgdrx8s+YmRBFwy2uLEsQZIB4LNBpsulDJ5MoYqyI+r
ZrAKhyofx4f4Z8AfAHekBmZOw7xyHmpTi3XwDDsYW4O2ahO0k14pM343pHC3ogu9MfB8w4AS8sBn
NOGEJDI2jsdyQ1QZlitAa9JnjutYKm1hGPIpJ9FdIiz2zV3qazpWE0CVx5lemV1a0/zyYs07d5fo
KmFMZgB8xR2zAf/pHNegCCrzf0Bgn+wehNhvKig0S458toQvLuZgkytIdasCw1si04xmptSnIahC
+XxWPnm0yTb+uPjQJVV4zC7/BR4pxFDDYF6Pc1NSLxj06f3kUISHnXjks9xiIDibQTZuGaw1xLY2
/FUQ5WHy9efkomB4Q7X62hm1Fe1JS3vaNq0p0APBpFilj6GvUvDnTs/RRIoAZH5kCLN/6oG/pCid
c34qcL9+m0BoqnNlR/JfciUVnRYp33s49KoygEurm/mQaOGkozT5s421MZSW0NxGf2mN+q+4GtRf
fhuAH0Dy27U1db4ea22Xieap8z1BCWPKZPHu8H86AO6K2by0bpxeI6kUPlvUPY3tabg/gQm7oTvb
JLozjy94if5O6+fyA+W/9V1JShLPRS3KYkvWfqGJtgdpAxrD+QdlRDJWdjTFIaQz/Z/dMn6YnPGP
Ja4SmZZfiNfPv8YRjFfMY+zXm8X4tv5WYv4prJ8xENe50EOfcnrh99hKuuWdS037E4oKjzS1DpM1
/F54LnfxbmN5Px5e4tPWLLwGGyk2WhGkAIvlTsX9vmUmET0hZU9TnmOmAPRp2YB1AdEYD9PORLGJ
41jZocderKwI9HocovYOYXmqSpURWAXzizr7Bup0RP//OeTaSihZPEiu9IjngDPu1Bv4uqWJ/IzA
ZFlNqj3ueulOa3FaPJOa4SDUbnn8EvUFc2CVRPJ6rPeG/TVvWSkn7+UGnf2twd26ht9tvBqrmXin
TP8UbfVP2Ve9slF9bRFPjMAH9T8cpOzcz5D37kiVZKCU1BkUZS87V3gCJgiqbVrfMUgreq7gNHWB
ExtzljHkDdnSVg3kyoNETCch8BWh8noF4sL/Ln3jS+cAgJYSC80ds2+NfgCCMFtz3przqC47QcGE
j0F+3sQdV7NZ3KQn9K7p1kKOgeIsxQ3fSXxZqO1CEMaynmkyujw9ouvIPOOXe/J4GtzLBb5gFlbf
6WuYMXJk1z41jDqRo3lzbra99vjYsOja6JfaOmDS819WH6649QBhdw4K8hOd69XLnc0DhNH6YnS7
NJK7SX1kxa64Xq2igfK0E+kmrIAFAfqO/wmwjGtR+ODKzNuxNcQggaeAUjxcu7DEzzFoyzzO2FGV
/uhPc8VJvy4oXJn8Cm1ZphWsqjAnQoZ2b+kKiFIJrvYTNEt47xVxF9pjzfvsmYcWawb5e61I33x0
nZ94acCcg8ugSgzlYx/EMSHeo8Fq4Rl1VfGBsNJwqhSAGMdsp33rxJl7I4KEoJoRiUCxHVUrmTCm
nNztsMj7UoBRYr0HmpHaZ6Ua6hMrwxTSDWoLN6/OkvE5+OU3RsxQhuyRnZtQXejld7I6V2t7hWDF
y8KAxgO6vU5z5pA3a6Iw8qpab7vpbnVT4LWE1d/Q2nxD5Cgk36TXYLzZGddpYrEu0WEL7FecTFnx
WfwF7FI12cr8BVD98dHetvLRKcuX1pioHLy1jaBpJ/V75erJ91gPhRJCw3UXG96R27cPkGsgODg+
rJy5BCrd3aa2FDlD1qkEsW8gySTHZNZZQCkd0C8Mkk6/rCTm18oXMHFI91grHqbk8Nev7tci5WvT
uun4Tgzs99JA4iMRlUN0Glqdz/B+5DvQ78fowNdFzyXFqJt1Hm/7v4lT8dip2nyyWhjopQug0ENC
DHAxkW+VmtjoLOgT97Cush4qv9oaMOLtWxh7TI4Ch7mK5EP3Twy2YOukMibwfE2xsh5AUkOlbZZh
WImhxk/7TwQbCO41D/K3XVwLEG+fVXjNXhdQymLprjehqMle0HA2/CZvBAJtFkNQE/LX57pUBlWB
GhMlv8p0+F+fu4KFwMWQ/83PaassxoYwClv8ZGUpzp15pyIPWZTVisRe2w7ac5l/dygtdRIlPbbP
mgbJk1prFUtKmkXUX6zcAHm0I4XOOEh5mwdoCs118ZakIRCbYbiV/Amv2kwDVbf5GMFWjq8SPuJ1
THAOgRsTDl9Vzxik/VoAwvJnHlE4Pw86MoM4aa40C4mq0C76l9YonAP3u0aNilXgz5deHtXm0niC
xUM92wHG7h/OPzmgzfS3iiNNut/yS23H+yaN5RLJbkfk3MjL7j04uCQCNg7Q3sb/gDn1jYr4rjoO
UhROH7PSh9QvIatV2RW9XutViCYkAe9lgfo6PIDdnvSru+CbSwvQvX9uZg7TRuvHAU8M6GirgO3X
N4Rg8ARxrDxZHkyKJOm/BPiwcpOOS/ObSSoYiScZfl2wkov+XsVutorF3PS4uK5LYzkIlfiTd2zD
347BZTg/gFHnsWS61deDnlBstf9v5REmme6VaSLn3mu6zuzj9jUBLHGQdKq8DNr8Rn1U94ElMDXk
2oLANCSFjWj4UcmOxAE29t8pG8Oe66qH2dFX0DDfF5QtYh7kzCPT4UrDb5Usrro/yJvr1SSTLdmG
jW4j37rB5mzWLYoT3FdX/HBwY5u9cUEugto0nHM4UVzkLAwgRT+AaIyGo1yiFNkoFwKLzLlp+wU7
LsnlJYjI/Sbq+WHR/Ws0XwKsubQpbmInwtbIrqeJ4GZDBjqlGzAjsA0juVex0aR5LclKlbJshMli
8r1i501swmYErkhkwVfAG+5Amcidx+2xTmyXbVrrggKYBhwIoOEGyfUSCY7zrZ5lkGJ1L25X+4Z8
otU3Whu1jn5UREJRF3Q26+qB937vGDiElRFi+abxS1WB55eR2gfdBnpGzhMuzvftP4KORAvZk/bg
75/lZTN/cxuONbCVwkseSjLbu66vBAn9yAtOsDQDUq7N/RWouiUFw/nMBGEMlB5lufRY6pCqEs+v
XfZIaTvSiUCLI9algThkJviKde4NogxRXS+D69xhupVUVB0CYZTxQL2YDCLNrrJRLAxmrd6dpZjC
0z2o7Sz3SGbRAPvGoUPaGYMZr3qRrmKnOBdaxgBU70zEFfgTox7RNe2JEm+nPcBDph1hhpG985Uq
ZFuhPkF4c3Mb141z3jxk3ohcQnRBVo129kWV/u0JCIzh9L4Ab8euq6vVAfzmj4N5fVQK8/vvv9r+
PgvPKYPulOMxsp6MQdHXi/BNNBdS2VoO1qy7506/OG7PW9crGVYTZ8/P+Y37/Zv0aXo2fKdavpo7
DkED2fMvB4UCtS4uBlEsevfCiCnRvwvQhYLQorZv+EpL88Q74cbLU878bwloFy5glEeLvayRddZU
6v2RofHEfUUnPW2ojlmg1f8WoPtqfkSjZNmUjqp70ACIPPhKt5tVeEECGnJMKn8tnPV78/cPpXSR
Q2A8py7qKqMKqtcUr04JgWDAx+HuKf4ELCOqYGVpnv8moLe9yr+8xKUc46eLy4nEU6/LP7oKJC0F
fTXYHbRGBt/AEKVd16r+Mpe+2aTwqI6VVNsaAC8LMrI8eM0sanug+bfx/HJsoAZo9z+OyksioImE
7tgFQOZkH3zPLImnHUKbeC3Zkk1/HdASgchttSzQB+Fxfe/x78QaZW8W53Bs2Z8NeU6fSzz407Le
o6Phb8wLyY1VfMtS12buTn/mrPl6QTHJdR+4EzSOLeM907x2kyP41R1xe/yfQwF/z+UrMqEg5Rc+
isfdln4qRZ/5oeY+Q5OWbaeJb+jGw+tjRtWpGpRYbfuAFOD5XOx/cy/AffDL5DJmEmKEFlpBoHbe
yRB4x9+68dIjdxo8yRP6E+LCrEikkYV/OsKzKVjvlkN1hTcqIbufd3zaPbfWw8hHHnvcMVQ8eEt8
5RXEO+HidtRc9zYkiYZxpM+vRsXnDnui5gUaIAiF46PYzPlHkPXNTKlx+MN2qoja8p0lJXr3f0oZ
YLALm+ikHa/O4nBgn+nhaWazydsP0OLoJbwIgs8OJTKZgB8J8NvEHDtqjyj11vqy0qxjTIjwVy9c
oT1NqgYi/32jf+pvjP0IFGfDJWhnNgz/fMTxF3s6e6CNzaWd4Mv7mEOfNB3+hiUHdd32DoXHfseG
HAD4UGsC3EgEEnYeb6TARLDTzjlpwaTiTb3DxtFRzkoCLyOmY1LzCwz38DFbYnnErGmERsWsjPC/
9u/j6IOa4V4OoQ7W64H1IsgvVqG/ZuBAQ6PE63R0P31uTarwB/zxQ+BoHa6JTe/DIFuwAQDgnhf3
wPDHm69Dkc1bog90j6B30oARrX4jOWZbR4JiCq4rF3Rj9QFOY2l2zCUysgsWXgio9D/I4DtduoC2
sN6kmA3bvcwuzCQBjOyE2TGiv7BLsyJfsiE4Ed92YZcnjQn8GKFthZmEHzbkxTTCCxTqlBMvPy9X
5QXJVEZPUEpOq9pBdr8KAhLdeVt7AUOFi7IdEgT6Yre0/+2l8ES2odJWdLjHBmo5z6bcQCS0SAS4
f2Y6Jenfqn3XuN/k7sGlrkeBZWz0WbLdn4q6n783qT8KPCSBQ/JVVQHomNNVoUBmhZjy8LHwtYNS
GqptXs0cJ0jl1pKg+B7mVp0RvuUKfv8i9PeDbAk0Ev5+AAV9tp3gq3oJYU6tSYqtnMZeQHRZC4AS
bH38DIBpLOpaFotBUIu8NHjNQAmm293bz5djN8diQqHfKuEQCdPdnrMqfaGpjrrLbBzKYiRMefky
K6pbLF9pq53cSAXFcuqW5F6i5vgyaNC3CNwmjcnhOjexGFQdneLglcGPLQTLy8pO3i8eZ0m6nPgw
3w7BWVqO03ZkW3uPUiFELGNheDcG9ViX8NLUm8yWzzJLKUrUPYoyJNiZRgwsYFoZzedWbvS4Sd0i
M3dcT7fjCi6DUlW9RtqExk9Bp88EHhOTCILm7Se/BIsyaCKFLV7XuYe6sJSUbFMGcfdwTIkxxsCM
3Y7HpwHo9i224GcpAUIJiXY1uou7i+ceqqDVajibs4PIvmXGuE4WTiS/1BqaPmXdppwLza0dWBzG
w9cdggid9WMfPAgTXlPVFk8tnzQtYNkz+kK6fSK6KScU3nC9SWvLCiYvVhaVz+FlGT561A2IPw2d
s+ukDfDpxdI0/9FNPhaqia3mOQ7BHP/9V5Zh5LBe8lOS8+sUtiNSh0qm40c9qybkZp8rTDClnR/J
RE5kAQYZ9hlg6SIZpUVkgewo0Di9Bwq2TB2uIEkipofmoaZ6V4bOEuZQClRpLk6WPLxNcs8LxHlP
RhfzM1y2AY9dEOAUl8dqv4QkvYoWtRso53KGemETdKUgiYu8oGjHxXaSxth1m+oHXdCwdnPyuSes
Hq8qIaIQ4/0+wkzelyAHRKQf7cld2wb0ksMclMMnFD0oVc1TOQZ1eMeadxJFa9rlZVZ9GRUGWf8T
BO/ZXaCC7ZLV1bLsiGslnETCcDNFLsxWzayXd2hwVvhTXZtTeg45/UHiXuaTwmUL9Q5vIqGdK/ow
g7XLgIy+GQuTrIxo0iRbKlrsBnCDbLM7xbkv2UQtthSC6M29i7x6cT4PolZKE2+mbPplVcIA4GS4
thoCGFfx5ii+HY3HVMR9AQ9Vm8wFixBJOpBAbwPji6hP/Mm8PYvQKa9wPaNnKTZjhAKrIRaJkAPX
W6oz4myWiGn4we5bkYHxo4WEi7JKLuyODBCvYqqLNx6O6xk7G7VPbWJS59jgYSmOMuB+GVv78xZr
6UDsFx4zNmsHtaFrYsnCRePMEsE5QnvnM8wn+bba//2zXsyQnqM/LA4B3SMruBKDfjZLZSDbPJCQ
CPd6Y33cSYtZVShPWYZfs/GBdtXlQPj0lRrJymBns51lQcqUMmNrBT+UvYi9fCiwvobYehRqo2un
KgrxnOVqjXxDVM5qGxvvAkBNTAv0LfHZXPg7LHdYRqyhapVQs2Su49oiCJetu/B7B/EHBMOIq0gR
AT8jd7Ojx+mFCfoVc9LMEZLsnuFn7Il8uMKvsvBLXiQCsP66Ca9DU17NEuXD8bRmnA4e/JTjFpjQ
kdGOOAhJInyWmUmJR6gdydxVFbAXRLTyr4YIkJkHtMai7fx1/2kj3OjfJHt1KuarkXGYAQhoG6ux
DffHixPF2fR36dIbAnIosLNs5QaMNd+y39ZCgy8XJ5obXuDv2CKF98PN4PiBSZyc97QEoCbIkOsN
QRKUdPWktyBHnYUQmOqpH3E/RjKvLrELgU0Q07o8mtIwuVDF5ZfhcaaukREVeA3wzSpTdAzl8uJW
GQfD+Ipxr1g5SIgO0uI5fYe3Nqt4BNtNIN+3vmNm9snQpA0EIdB8bfcvUK2S093PQ8aXLRmfBCvX
hyFWo4/L3Vmrg051Tm+zdpq0KtV0o/K+X9808wxURNpOCm5wfsptCrmlc5We0yxzD3UMspNbUBp5
KDFMeiGU8gZzWqt9JdxnDGsG9lGBVeqWNIlrfRZCR3ZX/e8KISf3l4Ub015r0r9QiKdwK9Rm8dH9
9xFp12g4gcwINAPzVttGThiHtbptpXMsB9PQCgB/DUp0LIHuvy0FOC18VvXVDBxTViDDp5cxtZKl
NPSmts8zC2fBVJRBpBH9SywoeI+3qL6FqHY1Vg4WSx4GH+Kgvh08MZ+lTjcOUJ3oq5Rn3QgA0ez+
Ltlm1j5HY3OCJPjeYj6i48gYnxm898eBmrS0oIASa1Azc+dpjeSjIJP1nkNMlQR+sw64mYfYjoOC
IpWVX0Qwdcn0Yp3MZC8OrNJezRSHr7e/ILqV8zrqqkxODnnmRgx/GXye7KT5DtWdr3YQd8Q4yVdA
OGB8ORFCMAkx76k/XR06/ptIAafCwAHFdS9x+5yQbg6cQNw55fq4Sxj5JJiDTaGmmZsxnViihd7y
AWkEbkAMjfw0920BHKriulbTw5gykaq77H+QySlDwhrTgWXVyufId+42LMrOmy3VrMJEHtj9vCxO
qqxxvhsrIYHTGm14AkBv6qMwUtXsbquvPcifLosDoSSqV5GjPKx8G6J/j91YkbR0b8uVmGSYSb7A
5UfCpR6tXtSv0rN+OHFv7KL0IdMPdQqL5JcSu/ME0uw5tWu5wwnBpNOR6HvNyFSxakQbAOblgzle
W3pBchfdB9hp8vg92DWms+FErPYwPVeCmX57PrxYnywnVtLcgL+7GikXY/HuoPfcLGd+tR/ttnjD
P0RU0eSnM4PSwiBv7Mun0kCJpJ3eRqFYDbnf7Ilk89xrQ79UTxu3a/mbDxbSe4ANyFMQmEXNAimq
+bQTGCGiKGZS2aQFRTOJONMkPhf4AbM3hMtm4CxaoUbAAlAuTdOC7SzUGZcVbp59yMFuBc5VNWNw
3CiGBuFwMhMmrDlWCdLrjd+eJs9Zs8uAYTzJYulrdn7bN2EoqI5lK9qK9Yw1LuGW7zdQAgSLJk92
x74pNqGSj2TcNwwwfn/Iu5WvV2es6G56yJXR4yUlCQ5H0CBwohly5v+8JR2p7m9Ca10oM+J7g4T+
G2SQCwoI5ZE//M2sVTevxAZRCNxE4fZtXjPlKEfORrBkiNf2YkLDZGpRoiRUjsgpB22TYYQFIiOu
OT+jbGIfHPru0usSVX7I1cXaHrxMU2XVYrzJ2/SmsaRiN+WL/6DBOwGrR1kxBZb3BXnns2PRiX/G
aVaJZa5tJg+PnkIsTUzoJF1BXbPlezLAfGsu+J22w3sJjZo+S3eYv8+VM6HO8xhQ5xscixjcn7f0
zDsf2h0DqnQDsefwFDUuLn6hhf/SyE8/B5SSfduAargPl+9JjPQn7vQL4z8UQ1CkEhxMz9EJOgLF
p2ygvHG6L1oHyZF4HhFD/pcMXGz0LhnEA2MSKlDRB7HqcU9yFynY+KCcLCYc4KsilNFLKYQfBwYg
D/Ne0fiaJ/cSme2ihpqM21CHmUIBlMuRYpwH2HLCGVQg0UDf68KiXJGc+6XkTdHvR91Sw42yY4Bs
LKcn9oSJQ/h0jJ64Rh3EJzMS42VWKANszZSmRoHqpeg5DgVvO/9dP2Xj0Xq3bgyv2LRTfIK3EZqN
0u+TKhbxKNw0lFtv6D4ko7Vn4b9m7GlVTkSBW5+Vk7+L8Vyt0FC2gZMJg5nLaeXXmuxadPnLfcq0
ueBzwn9E4uxGcn+Cf/Mew9uXzUHuCkg2Bci5KISG86th7Ti3pjCtavQZREIefWzj+dS/NOUNee9f
Psri87QucHkblNLXSC/kE8n/nopQjXaVKzqjJAHt0U81LVzDYihpYBb3dEVgzR93RzGZnJGeXrx0
IkDjKPJTcrPBzj+W2Ezp/aJ5JsG404OW5NPmKmGqq1OPEQ4MiGdLuHZhMvv2FEPs5ccU+x8yj19v
GjqIFmteKJcebhITX0VMIn+RZlIBL6JawA6JfIshtslfJeLB92UxrcsFgtRahjgm2nBRi4XD6nH+
Tz8ZK7VTR6xaQIUT0gqWM/gMMh48YS8CkBieSff3DXhcouegyD3h37Jp9xajlS0gUo6ZxcHLcmd2
GX91jrhtBWlEz+FKMlPEaKsI9JFKdb/BgpUQittXk9MxlySsSo04bY1W4zi0TDNaTo/EZmtyNNoh
eUnbdwHx6V2MbLRO8r2oSvO7xzu6AR0He2OLRLRk4bvPZcEvEUcWM+f0kwG+BBgf3LBXXwDQKOLr
iXFNr+2GGA8c9ZYEKGaeb2zI7KeFmq5wt5JT7vi+huhgP5gp1Yz/b/qoiSrt7wQZROg0dNbw8/r9
ER2sD/eAy+ocFidjU+MBYjt0tsb4z6AkJYmxT0CNwr4f5FqR1Vuzi6GDs9dnjs9kuM6MXKE30EdW
C0kpUac2mtyriodTY6WE7t+g8WPS2OhNCCM72qwYcOgHjDpRH+OU5Jh1Mkx+4sYDfasso0644u7y
kPypR3S4FEu1FQdxCsLEX6gJXn59qJ11mfcyU0/iV8o/I1G7rUb7PZKNXWItaO+XnBKGJQfB34Kv
KkOqdfGDbSQEPp9M9DCWfbvypdq59kTD7+LvU5cIONJTSwBL4/srVNHN9aIxkK2YftWEoy0kXqM1
zk3f5brC5f1IofCjbvKDm5syMR/PKjXBVPwCtU5tnQ1fZAh41mIIl5HB2u9om14Cxl0hl1OFYAIc
qogP2oz3U59jXUe233jnaZiA0FNLC7n26FGaVJj8/g8U/vzXZYTnPYQMCHdhBbDcTh0dhNXvPLIK
GhqJzxTZB3RP34xGnz/dcq99pnQlL2Z0VnNICNsN+Fl4NCxq0KjXfjP+hLr0mxZ8VBNfthhRnC7c
w5L/XAjbzHEj5GASMP5nC5OsZRUvHj8TUWyZtNYcXCxRaaM4y0f9ooaIEWMTnM5q8LX6SezBSVWq
J9ciLAsU+uFyEAMgAww3rtqCi9p7SK3EJ/DN5kTtQBmXKnxdIWX4+mGcfhSpjzvTvWckC2FmWG0x
SsupzskJy0bwQTZJTNL2CeADCnhtLLtIzS/JxwS14DeujQomDqlSHmeihOQmhfR6OfLKjfDlAUSN
el2CCh/ji72Igkbkkx6ZJUuKeGDi+PdFk2BXyK6vqNkpqu0BXRYX+beT2DVwK2QpZA6qi217kp/i
+rD3X/nL0e9OyKv2/a69IehMuSQywguBnNMfeVl1GG84ZWnp1jO/orzBHM7xEoo8PczasnuigjhB
O70l5SJ8US26YROF/aCJ2evSWhJFt45pxgHatcv3PJj+MRguOUCly9viCz2ilNiWC2EUaAte55oh
GAajQPfjhQVztRB96mt+5pbvp5wiRLBxS8d8PxuX3M/G+pbnG7kaxlSXxEMG/qZmpiQGVEJufTV8
g2Tgnu0rxck1d+kL6PjPzKRkwooZ45oq8WWAOz+1vGD7inzmgBKfSXGgSxks7pVIt0gskys7N2JM
IgRSOgVtt9+QN51TEJtQq3DDNtQINOOEscTmj3pYvsFfMkdOvjai8l5fSLE8ZByUxYk9GmWfjHx5
TmGtfxA7Q7dzdLYFgYiluS+bhB1doMxgyzc6klq+HiLSQ6xDZ9A7PsyZIMHNJi6jVKu/KlwuUYmS
p9UYBAklSdselo3X6bfbyCfaCuUHTLojOEG8czJesePGmgN/rfCAlkMRYsqrk3PH+xP8mMS+L+TY
tT7j0PoqnjdSE9U3dU4pLIRgaS41072ABcyVyldSKuDVpYMzljGp2EXW3ZU4gtMyfBITU6qd7G4B
7rBnd6Of1Y5QSE/v65Z2VoVPbC060jQ4rgtMv7KURCqvtDwY+3/3EsgLcyCa/AYpZERH4X0o32mS
mtpnCIuOv/GHtBu0AaxZKHUagnoxEkADCjvy4IYiza1KyiZq+8wV50MJaIkiB/BySjnAV7vALmRU
XkyKaMWipfZBSOCgRxAn+u/XbkYSZldaO/PeJwFyR3JF1D36p259y77F6rJpMDzlLWP9Hut1xSvl
q+ePCgt/hGQ5Jy3Z7PAbxflrQMp2S2zyxYeekopDMbKwD02X7nJEpbKq4sc8Wvy6G0nN6dBsoIpS
Bw9e+eVj1f2yrEFAjZrGxAlgoCycGisxGuEr74kHBXEbSiZKdG5ANabf+CCTVXmYIMrc64uXIMTO
pU5li08f+aMlAj71tjfSZLJ5MnVdPEF8AHOoVHiA2ph79bM5SzE3f3CNeulyPFj+1IwVLswC+CoA
gZzuvUTHtsTHXGKHrP+AENVDjZdz+J9K6t9qAI5MiLaQHAKI2bsWmAjMcqv6fPvT1AH8Ido9S4nW
jEjja39c6nK35otKZjxcnSUZGAjRwbMVzo/Qk570TRLH9IYm5tFR+x05yKiajiVoSPhctaFTJuNi
IsL1LDkTaq2v8++Lb0mS96QlnDb6BU6c8Ny6/X+82lIs/eqA5pq8zYK6hm6DbztNZLGffyG57aqS
jWwcEM5XzEaKP6hH9MgTLZhabUn8pqZk1Azf7e8ImQAevX1U+Z1jh2UWlx94Xpj+esrV71rQ9K0r
JyEhrXKcjl8qPKKKr/0Rt/dWqTvbZ+KeKlBNFXpUbUukcqVuC/YjbMBCf7t0gfARAcZM0ZNmoKIi
tVipLKluYi6ynPJUTQrULE6qgwYbgDPL3kw+ZjEqwGELVM7fQD9yrKstcHSYxxXKqRBQJGPVUAEY
xJ2nhc72TllmUkvm+SUWuuGSs682a7pLRLaxSeBukTHqqn0EKwubeK6N1C5FL99c5MS9Iyk57FrQ
0++n21QCo6ulRAfaF2xb3EZISmuMclPsFTBKxSBIkAo/MHGYiyIzmjO3+gUvcHGkhXvEvwgN+fuC
qgwR+8eKJZ6K/WDokNohIDUCj3ZWTqJbLA8fp7d8xD9gaLRsV5QJFCx6lOgnNqI3FvgdYCq6jn9P
E7N3Br8HjzFOTAVn+pQ75IGoUn8QQH5ltRxqFql5CssyK7Sap+pmtc8mZ8Nhj0RT4mdfitzWdpM9
zBgKD4CsMnnUeEcHsqvAf5eMCE1+xuQTw3VLLrT3NuYyaNsnMcrS5tG5o4rv3JLSXYwG9ad2AkdC
2zAWL7J31YQrD7aasjUn/63FxkEp2vnv+uk0na6UZp/uCS9JMsbNpVhLzQ62Vzw2rq5+We8P+0+g
yqwMSSvFV4AK+ySvAMa5IRHxg5zUs4FQcrR0owgJFJwC9qxLsk3p1eQRGeXIAUntvP1uqCbTD3BW
d9gmyiLAN1FYL2TaXOBmCKuXd3p0fSoJmf4rme9ocOOjBqNP4pu6MPKXFXHUqt+ULWUJLmBJJtvA
7KT31QUZr68/9pXsugMauVzopiYNDv0YgFsuKYXNtcVdMpeaCuX9spwz8Eh6sE+jMeH4lw/v9P/N
ZLzjOyWHNM+kmzgjqcfj5sg7fg3yuqfEXitRSMOWcbSnCzJF7pkByVj7juBXej9Ig1K4bOdEojr0
kmbvo4PTtrRbSHdLZj3KsAteFmwR+gyLec3Y/wiHNNCPpuegRc6ZEAFSdz0WiKYzYXkVJVA7ncye
md17F+G0xEzwLgs/9VcHhvzNMfk1fuwiqu52cnLrtwva7TtO6TbpV1s4+K3EGDUBcChoqwwAwpql
vynmcxWD7LkM+zIeFna0LVLzKkDRyMwf+iKErTb8O9BImPthxSG6+7livipvRotRtdmU4URt6qaX
lVkcbj4arTRskzdbWfDVYgTWhwj5xv3crVwnHjljMXtyHr7bHXpba89CwMfN06nThBUhdPvFWp3G
TIWo7hFFrmudRied6/PIlV4EG4ARoM4WPrXvYqhVtAogfCO5EdOhz6J1nPCPrBRHIwFC21fLrDph
Keq3VLStTm3kpKWETqzYXr+2jDPUjc5pELPsofi2Qg+ssazaE1Xuop6fZtlJ0DkBU4DIe1ll4Gzk
iw7I+tmtRZMbF3gYPHIOtcM2VGPix6ZegaGForcJjrN6277PG57U6DqELrC2XtMiPxBJIlyE6yse
ZhkvtJ3D/EklcM3RkbEHfLbVklMmTA1CyGMsaJth9TL3GTraSI9Dj7JUqnD+woLxV/k80QE2vULd
QFCovq8YGeBj3Zx1PrV4+1duhT2FemE0s/h4W3+Fe0TSNlUGxNzafm2qp7Ny5b2dBgDgGTcYIjuK
A+h0w8jM4K+3sWjNZV3+Fvd0GhIJS9JpCjv/BMbnNek6meDFUO4sgDh+hD60q/tejOTWfe5tmiwG
TJ/cwAJ8T6SxdEPvSaDZQOBJa5c22liA2A39q5+FuOE32/fc9eaS7RSqYYX1LOyAtcJQ5IjjWou2
q3oxukoXCrEn3qVrUZ0JFCNfZmVJsMeCRx09gmS63R80xJXT/ysUNMeL6bkoAHf2q5XxOTZWbZC0
MpdBZMvSMz1BZpCfJVM0E0BAnivEz4b95NDJY7naxTizNhwyC3SUwokQLc2ymgZNAyciPlGAUS2w
+mQnuIOZG/kZeal9YANZMcxxXaoZwGo+O2nHhNVj4Sm4esTdE4PMPoRUseVhpWn91V/2n7nRGYQH
xFg57tthzwkAxt4brxmYVhkkGG9sU6/lS5WM5+W39RlGZ1QhhksEo9VAgSr/Xur5QrrwFSg4Q+7O
XQX8laCqivKAm3IZXIIYliyal8pTp4+c5pPu3SiRw40DM/ECMF/oPUy6TRvraiNY9jD3KsU5Cqtf
bP+iPXvDKiT+zGXqQYfISyTbrqBK6PHJvEcpbnDl8hY+0PCwRicwJOPVkyYPyUxO31mw+tZc6VUt
G/bYTefB+IW0xNvhmKqtBuP83io08pY4jUb4ctEsA0evJOhq7AjyIAaEEwUBzTTDwC07zfzKAGer
Q/Cxw3iS1gUfnzmn0ftWVweLupGB2fBuzpUj3GvCrzcVtdZHDAwn1fnX0vnATsn/GtRvIO7luvLm
ewWPdE+ZFUlBFNouFY+fJBEi+bSvzn3lvjD6CjbKVWY/DfJeYK+TXSYzJo69BdbPGbK3kx3tjPVs
kGSlWEz0Smr9vNUjtWNwIUetnqe9/zw/CwQbIMhlRdK6UvEr54cTLaFtuInPawYvr43B4UF/ILAr
romEKORhPlkdhYrrtI1NGwyVGfNBpQaJx+iIJR2ZOrbjmp7LxI00pqBYlaqRMCBNnXiPN5O5xdW/
aAId6QRNi+aHrsDro46u3mCMgYQQcgBObi2umZhSpfuP9XKQ7ekEhHcCiMiqbUxW6NsNMBerYzcK
4ZDvqUmRnnALu4MtGCoO/y/jKNeE5AnUkT2RaP1QMVKdInI5DMhgRgc7fBI07RsFm8ysXZYgFmh9
1hK55NdAAYBKO34y38dlOixLggBfPKWY+nCU2ZTmHpHXsk46bW9rrX/TCNts5NhzKc9kHa/vWNrX
4PtE8hRyOFNDHD0Il6zzH+WrWWKbIBn5upmx0XLnFNMz1z3Hvdue4eRtC6JMhr2ZxXpHyD0hcIXj
ozhmlDmGsIcC6mHF4wbqPX1O380NNVF9k3JvjeckO1tnKbeBnBej5auaw5aCd25PuEMh1bNlWfXq
wHwbTRHT+H6JkWP/3q6raqYd5Sd3agxc9HBzUFqFS2a2HlIVNY0kKMN9siLdpOyfz67j5oypWHc1
GyCt8ihKSet9cMIblcaZ8S35g/JUYqbLNr2gjUeN+PoJOaOm93RooSgYDmPl7avXgQxg7oObt9ww
tZiKbsyBFIJOkCrgtMmFdoJXsM44oDEb48PJ5af4fy7VTJ2cmZpOqNQ1WviyDyVc3R1ajOmrGlvQ
xaBMBmK23NJvPWREs1IyxubkCU4V6LGPxaeEvwaVd4gOPPkdmkpDMOUoE+8pfXpN9QlDXCk746z3
JxlRP22cDCKQwJihAh//YdqKtJ4mLbdVJqYiVItW2aCN5OmqZLuMVkSVKxNqH726izyYTF7w1+fH
m5UryF9qRF9sZ6Eym+iGZJ5zKecbfaneeVxhciDI3ojbG7VO772ATxb+otpj0k4HM0nGrWPzecAn
fqAfduBNruLb9uYSAB8vd9ys+YBihsuPDl926Y3X43bzzsARVwP8+Neow8pqPL/oKIYz/9BqB8po
QPfriu/ZuSGIgBcUciDO5f3g/lP09JTmqf52SiJ8gBHKueraikqNKGPsupsfZR2q3wLm5gLUmehO
Hzx6LuOW4k6pVZ4olKe+Qs0X69Igv/8BMcGt86jVLKiFBps7uRjMiqqls8oBNfbdCijhZOveAqwG
iJfp7jq0xRyjwrTdgLrhzty7as9oLGn7+1XiZqjjftLJTRFLFyD4olpo59jHOGx7UrrGQN3NPN1Q
g/EOQhNk8NVxHQsXfgAFULp6G/SmE+30QZUT7TMfiIMYZ8aZTAThHNip2JbTSGLmE9eCQCnFdi2K
vqjUpgaC1TO4gFw2xIc3AIBER2iZL+27hbzxQgJZnkXvGjA9p/7kE+LiezS7WcYdGcAnfsk1FZtc
Ul5Khfd2UaTGOUf/J1z2r2LUl+inz25DosT9B8VQtJRG6SxjSL7lXFbmS6fkTkOmnSdmdqGvZjR9
i6QUTMtYxUCZiIB1Yj2W/iW4ikznToWADXQhBOiBhmohGDGkzPMPSOPn7zl7FAMoUJcWgzprZkrG
Haap76brPy4ASA0gDmhjL47v7kNwCTiQjYMdxBB+MvqG06v5SY6XIpjp8ixx15GF9LB9xi+4+S4m
FW4/D7o+bNbzUwcv3f/JzvrW3aVbtBp4QeHrRR5qaXaV0CuuU4KcW2mI27KuXj+LA+ir8VNZ/9oB
9GKMkux7MKb+zmTpRBDmbrVZyL66h8YHykC4tqo/ImNM6+n32frNVANWhYE3z7AmDVzPlA6zjWw6
W9RYY2uRjqMeB2oIRqx85wt8uAlp7OcziJaXRO5+zcgVwFvkGLtQoFEueK26A0e7GCzh3L08Q9Ws
J3biVFlPJwxB30oJEUBjZpab70S62U1AZZdmlJAAuvFqpmwMHL1C3eyIYRwKFWT3+Xque5ZLY24P
n8fZJd+dzelOBvTeBfPtWUMEVge1ucCfh/AidOlUYXMyRrk9p0X7FRU96pjK/aMlH9R9VIxaV2QX
zN40JbN7Hd/ZDPqplJPs/7sDT2P121XyOsY/UOoTcyvUOysnfvwVMreVwldB90E8Dt8l186DX4oi
ktoRntUBi4ccfTTmi+Mj6B9tl45s50VbnfATLCpQX2CHMOk27gTYnZXXtTOBAneUONLqAiTm+pfq
p3UDVHIN3IyirpVTfL1e3PSLo+XjE7BDbWkxwmpheFGp9wUaHqkZ3ax5dccuuLnzra32KOsPshFU
mfheaLrC6VBIG1VfTirS8xabnW4qdBSmMIWusr9ewWotRiHK/s0PIEp3fl6+2UJNQjtJMD+EzC5b
mWaoTkubYoaxW6KgdjlHFvrZPxqH2GPw6ZeEgbIgwR86yby4+TVgzAr+LStMh0AnMFPILHHuxa90
2tQXqoMKKJ20sbxpZiSLqckdR7PbeJbkj6AsBE474BleKWPOxd+c0t1syZm0I3dzr6fkBOS+92ku
vv64ZNa/CAuVgwpBnPEWyDi+2DbzQAoblUhJ1O1pEMlyKHYuzYklq3XvFdxq9cPOQj/hvE5OS1/Q
uYThyH/6DrAWVCG7B6+T47mwFH7tbKZG5fa5W3jr6F/vQVHZVgixF3BRQPJW9faK2IIcb96OjjLe
KiFWnZqrExrHEGdJGxZeCbBuDiFy3+4bfQyOX89qh1xgIHVn9bLNKYqePgevgUvAoI8Nf/aGtyZk
9/WL5kybTODA8gqzUNn7xvvM1+qToK2CBSMNcdljrAVEld2fRwBQbs+IEC23+nwkqxYtYc+R28YQ
qEJ1K4cE6/1LXUCETAd+FxGKwaTuTisapT+rD7F8ej2iEM+gbcFWIxZKLvNux2cyiUexMpS+UVI+
oRByLL21plNFMrxNzzNcXojSESjgZShUcVtU2YFR5fTmcxL3n9iaG8s1OUjYv/Uj20DyAHN1iwXU
w0Q1x9LRQskoFAFCNR1fZKF+1IyHqoDB4/Ugv7GqjCTlVwJWR6DPkmh6UgnlE3yFR9feD1C9Ck9D
Sb5ORNLq/0xvCQSYDMryktm0RYoFzIjduOhNRZ4Yh4L05qJqVGN4anWgUlW8IMkKT7BDBdJd2MCW
H34k8UmFsiLJ0ssHeuXRbZWk3qV6j6EbAP+u3X/JuxtC+yBprbE2iaIMmViIT4OCk4NCGZtZVMKW
xF5i7h3kh7dHXaqEbR5rS+a9MxAM7Dk5DMlkqcEH+ufqFXA0sQvWp9Yae1sFY9bB7HKvqxfed6an
TEF36Rw/djXegqItYzdKNdpqh5nKXJ90k3HxOHs6PJ/bbkceQckJ6wjwId+SSPozuzIZhY3Vib89
Kz28BMfIO9oI8BGC28bEb1kSDnXj/QnqdNEcAhBv2G+IMQEqcnbzUtpPQIi8qaNfE1j1VLjZ9Z5+
Y973+svejBLKZO1a5+Wv2ch2zHuq7Z2n0uUndGQ4udLSi0PrlwglBXbiAsUmn7L4hSzdEQ+QzpFg
2B9NoJijkh9M29fJKYwIN1EvBRz1aisoG1Jmej8993zU9unmrR7qT4LUOtQzRTyZeeEmjRse6vun
mKv+3l61VrHaExNGX6SEWnJQRaWvz+/RtLUhKHjkdqn1zCMJAJjw0B7/C+VbJH+J5Vlt6H0cmF7t
V9fWeQ3ZBjQsNkrIbDovYTxZiorozJCUd0ysDLowEGDVNIqLKoBO94GBphkMX7GajJSvZ+LTWL6i
3ukvFIRUsTNbHwP7CSEOJdh1n3E4Mmplth3whQUqXH/Q6wB5TPVeXI2WxkAa4/kvr1aslJ+u5rff
SUjyTEPn7ga31taEjksyYJqvJeRbnKDr0TvBjQ6dJDu8ctNGdOfS9w3VdpOs/O1FYw6mNezRBsRK
KFCmtHTHAPHtl1FdD1QIe5FSCc0l0W7cM/xKjXZKw6IRWsZiV9todqNvbrMUKsGhhQS78yR7rR/V
qB9VvsaBEBaBU3QZOQUtXZMXqBwHMRqGDI09F7fBe7BbE3DSkZF5XaMVI73264I605bIccSBM+y+
W7cHCnas0oGYWGeL0Oz0MxVVmxkmeNEy40GMPdG3ONe5VPdvbH5Q7mYpFhaDDhbZYN1f2QiKZ4Jz
vidDLoL0PS93JDwnUMrT7Yr7uWGIGe5NmUp04ZukIfNrGwGKaizHas+o4l2v7sHPPA4x/+u9dnjW
xLxPCcx0Qq7uH8nBvnAZaG7o3uwIjo4mNCDAAasMsbSq7xmRRUa3DPsYggVzA+2ByaE90tPkr0WR
dH3BIg5bn62D6lKecbWMOQwY0VZadWlTme2ajVUN/dhdjUpFiEd5QW4pzFaDcJJcdJJzqPZXrw+A
SnqS3hTEG9C9MCGzwaOriifLoaQlfsn2+qcXprr4XHxJGHiLXcakgo7nXIz16jkRRZIkjiReJT6k
oI/XCcl0V+yb+Kr29V7jMzbGEqze4d6p4yuYXEHDXC4Ck72kUG6ZCfz8wD1xFwe+J8NFhYcjgiM3
9RdFRhw+Fn8GVJd3GUfg4GIjzSR6+SkeSAMiF4Dz0bE+y/LV8Rk16CT8oF1CFzYJGgwz1FhUaugE
Iq1DUTJ8/DWkzJnkiA8dcWJ90l41NQUFPBxGqr10cmKGyxqyX6M+earaUX034hNoUAMq/X2G1qPu
fycImX7WhQX33ZgzBRNGCiEbP2lcatu78v9PA6SPYOzRdPQyzxnFv2AEmFeqvsvpwp3meZXnbufL
ik658MgOPgS7EeUbDo9EF7SYLY3fN/FQrOwK0EomwXXCFGx718tO85xXayPQ6Rkd+VfYEJ16dJDP
QSDaAdreleAGrWAvT2qmdb555aauCsDxa/Z9Bt600VeyZRlsfN/63eat03pS9pg73UegTcaHb5no
P+eV9muN3BqKxtg1OZ7tk2mTMq7AhLsfk7XZOUXrKbkcN1PBsrCR8VhTws5lg48FB1Jb4kKF6qyo
c7ibJQKlE+qSIIWNyBxyBm70o1khbRxMc0t9aAD0MYtLytHVk7TSQVMjfd6jNUe6cxMgtERhVpE4
rdFhLc4hGCxh+Xem9huUGmfR8ha999eyOky8Zks8ddiBXm9IzVwM0XEgs0qVqs8ku3PKXGe+0Xcq
LHHhI0myVqffzs857CBSiQ/xQU4VE0bSEVZyrTv6gmdJxYHjzS1y0cd3gnwD0XXHtib6dDhoVKiO
genMMm4d2cqntiY8RMxlC9nSjlHvsAL2omclrykCUWdW8n3zD2Eye39BG3WnN+kfU9ZI/+59NKdP
aJhwZrXgYEA6VNXIob2SJWDvJEbbptFWLVieBITvQ/LhFNiQ6wNk0rKg9ftwlxEQW7ZP7EOVT3Vs
hMfcNrG1oJemrsfpT0xerMEXN6ziXiD9TxMgqNF/QL2No7lCv9CP9Kn4tJYJLp3JkJ95ss0eT4lr
5osXbemoq2IvznhpoK8kP01A7oLsmOp33YpzN6Ro0yq2oPTvvwEql8SxsXTiZtjMkV3MQ2VFkM9j
PIZAZxaqZAvZeNMJHex3exrMR04dkbUsY0jEmwwgJXS9rEs8mAFtDSkffCg8Jgd7JTeg1SNj21b4
pxe7lu2H/JWYAjrPGGK1EafPpJV1yltZbZAl2p9KUb+EL139jXStzI7StNa+aP9CRPClbrvh82/t
CKVnycA/nG7TCb4MCY0/dqlBs812TarjYJgmKhU288p/bmZWQsZMwb5QA3mxZRDyDSFjbO1CzA95
+SfjEGzSvnIP3Hvnbwr7dR8s7ufqReSEwIzoHbSpRlPVQMtugPkkljQUjVO5BD8yNP1cuJ5XMinz
OTLngRQ+GMs1i+5JAkl+CGEabus6tDnVXLnzsUNO1fk1P/AYPCivV+snQSDB5YS2hWVAJKKZFJ5O
uMjcFeb5uemlCMJSskxGc5YTNYEjVP3ZbCGlccS/xkJ3MCqemmCjvxD7HoRLslHCgfSitNFEcOrJ
g6tsmkUqxtjw1FCHrBfdzytM+O5Ibbkz52vYloo+1gemhB8yJ0vg+66KzKkofNCV61BO14zoS9ht
ljFUs4nZwoJ6E96MuoeFrgVZI0WrBZL1cKB5IofUeSOvfJRcmH6QcNCcKvoq3yP/P9XUr0qZrG6l
0rYVPkpY+E6i5LLR0JL7HPvdrQ3yGEg9rYSPkFX4QQaAt0j4QZBdxJ/tyoWoXaK4Zf4Djm0b18b1
gqe0w3JYFt0Qnj+aM0cCLUiV0FsdJPXRRaOTfQV+Xp4EQPUtasr5JXiYUCIw77OtOtRj+Onx1MfF
wgYkQHbiQfHFCnBWqULIC2kPHUBr5vVA1SSfj4hhPor84wIxvtC1vwBLsNN+GZqTDml9M38GzvKl
a8DB7zr9/sDvOkaD53OU+oAMX0+HDJeuaGwxGCP60u7S4bLPE4uzRPHSwHVwPaDIB9Mnd4xkee4D
Gnbpx7qZQDHy7ijYN+BWuDOJTTknefzHUgrhkAKakw9jwW4AHYlwOzHsy/uO8SsezUWfhv8Gsd1b
V+sVnQAux9OKt4dMEMFaWnohqXllskTwo2++afVjTCTlZjNNGoaGIicNjOeE1XA3T4yVKjS0EYHR
pp1LIGtm8ziE/t/MB+jJYVeQF3s7kNLyRV0gdHhIqvsvKaLKwiwc+K0uF1hhMnHQeprGpQLVovZ6
6VJKXLmEPP2+zobYNQEhPyGGah7zI40VFqGr7G83xQLM42au8n/NNVISKGIJJVrOOkZ+CvnqnRgw
CzJrkEFEI+p2+xVv2dhQzGVIMW52QrlZLc/ptiyiJgiqEyuYATMsNDBjeJHpRM2LbYUd/J6m6fci
c2l5vjPrZmby0NtZnIUZLEc2CsFOvph0qH6K6i5u+j/ZPATq5BQNFZNtWWtT08NpCGLq37VKSeik
YcQZPcAxZIxp16ffGnhxhgxBhR+Wc5YKXP4sRfELN89EtuUXMXitbj8NzM4gU/dAdvBHJUoZaM0z
P5dIBZGNyuHM3k0JkqGFueDEfQxJY51zLHXjIX0GrDQIcUvPxWH3LEBmqBvZuadmoRnCSqiaswsh
gMeaPxLQBjhF0XLb7ExmsmsdDT8yYjn0Sgw2xKqxcUKo0xs8YTXLrdKc60YlRxhMutnxfT5YfQAv
TGPJXXNnmI3I6ZVkbLRm0/2dA9UEA131Vy2BiuyxpH7JjgMCaoYH9IO3/9xxHS+klyxRmNTI77zU
SKO1vxDEhOJpy8hDAkpNs6NzQI+QdgeHRwJ8KEiUvZKgJIkeupkK5d8V29oMmQzk62XmsyICURug
1atbikVhXENvbT3Jucz4+jH03zRmm8aKHv7/grrFrT7pD1icmriPPynpX2Sue2U/o/N3ASMe1iwR
TG7GkCBiCd4bZtRzyPnhmCzcLW6La7gyN6Hga1bNk6s40JGmEtRbKLkROQ3tm6aqnSbxv9qYBarn
6gKEAGUujd8GnF7J7tTKHBVsm3h2aWgErH5IEOnx6ttO8tf7IlOirLHZu/AJ3Mx6CoKJ9RjESTKE
01vSMg059iAnRAnn1Qpk7z/OPibW1n2YHkOXQFxz1sHGZwBf/nh2iCsNTzIubdFBExnbHk0bPbE5
uETLKrTPOGZIFZRbIPwbIMEb8zQpXFR19MtUL9DjR8fOx7SAyuHJD5zgj+BxUiGxXjqFk/Sp1MM5
13SWSd5wi7qTb1Lwdja3GmgTDhU/HOZzMpBSn7BE6VoB5FtMRcPvy4kdKtcpRB+9dZm8ZC/npS1A
Dyv/X7ta0ThiCxk0eIfap2uKQhg0ilsjtRHmizr1dFIliZKgoy+25IUnG+JzmXTLAW1js0ou6eOx
Zj4yEiZ5EoIZ3NzmqJVWb63gXIh+R2qp03ce5+JGZebevkPYaAxc93C+DEFTt0jA1BGQSoDyFalM
yRF+yl8kvdwvAl3B4NZmbTyxhrUh5GqpdJcUsNZkaaQFDDWFXfNoPpMXs04cjuqljPmWlXbrPkcW
8bTx9AdAux0VV7kM5qJp5mJaI2Imkq5ZY9v9WgFdk9KbuBct3FVlOgNLufcy/4VpP16cMNVU26TL
bHqAjx+lim1tuLjCFHmVlf+cNdDnvNfNu4RVOz582U8HTtZXL/MKdI1jxlbhbdNqYlArFMqkwCVL
YGMAWFQQ8nPHtKahe4uUvLQSgMG6jsPqa3/4wB4q2fhLGL2vDQIxXxVjUrmhRWja3tsjpjjxNWy5
v93kWF47xjcfW5B8msJHxKXLZTPV6vm3RBzw5ovssyQICxkL5YFiPLWozUbgilpcIHTvbU1Xu3Wu
nTGxQYN9kKq4PqlymNsIM/NwkHxmYVOq/Un9Lb68uS2OuCZ3/ImSDxh1GvLgbxRRjB+9Ve+xODOR
uFVKtyyGTv9RCFEBdfvgkzVHBuE5D82VQ4vVrS47spgGN008aoQGH3L7ixAaD6luM7qKxBJZ4pj1
sJtuPGSWfu1jvDzLydUhiRdCTYyT8iXVr7fyHpC2scPA7guCo0YqPAv50sxK0kEpaBh5BdxO/urJ
jHwOng2yNbWKM2BQ4afQV12JPhnJpAkl+kWcDIi8oeCsMKCOwKFoLTtmmBZdq/dekEL/eegbzO3T
bQd4atW5QvjXSJdD+BFvPZyNGYE1pVcHxKZxMYVyxN0rTJD0hSftaQkwMh1MFdw/9t6xRNoKOZu5
D4wOYtyq3OuMRRni3OYOGrgig61mHA9xfHOmnVwzvFhNKLZ1zDhZgTMncQxYe35GEyZzCfcV658Y
CmpJGIQo//1KyxjFxylv+GFMHDFdJrYSn+FZFiQzEpGmDoKBFgiOsVrIWEFty1G6oVYhBocLfqEo
2tNbC35ssDAwMKUSsUKTx42JEzADXwwt8piRQsNp0xGQ7ocvw62qEfNm4hQngB9UsFrgs8w7dO3a
QzCX8Yd8wTHOS9tZPcCJUljt1+d9sy8vmLefisRt636HSL1Sj6pPH+7yZdgEMcRMEqocDxB8STFV
VOFeY4pF9Z1Z4FNxh9qV7GOfYwuISMIo7b0HgqvbXhcnso0GLuT6Tha9BMabAyIQ9BFIdcaa3ejP
AKl448m5zE47hdYPOIOA9K0y5ELLS/Hy9cEdih1nYMvnuQYPr6sJQXJY2PhSC9YN9/haRAewMPEC
NCk/03zCDKraUqxwmFQ/rjek73ow33lQ+xBgLKHOgXv+pM0b1jey8+2XaurRNNNQJY1Id8MWLkrv
/kSYhvm1l6ducztRCXX9Sjg4luzqJwBpLWJ96AFV1HqUJRcqiRXqfAZsoKxcwXnvXBSIirHAQsLE
5uoB46g5DRpHFwu061ATAnd2jXsTcxkwI/QsVe/GFMwLTVriOHs2SiOe0pqdGbnToz/h20D0/QpU
gXb88Wx8aVjD8I6J3IdMKjsnGuJs5W+QGA970qTBY/0MAByPQ8XHvyi9ByasvXCPpREVwwQYCftm
iVt+FGzSdBagw5bTtAZTcqzmb9DSd0pGPgARBXZN3t1x8qKeZ76vThbvHL4KnOk6b2m3eHD3BsSc
re4lWGV2yBLUYXS1JYB7Yaf1TR+C857UEDjmWnGNXHJjlqSHvteUJOW0YrVSiRToyHWX5s3WH3W/
HVTQSYlZpB0WbH+d4KzWfWg6DqLYaKnVMyseS7cJ2oWwna1eMDS9ezcGQryZ2d38U/gt5UkeKxbA
o/fw931F1kNkIA4hPZ4dE9vw+fIPSwqqCu477stKx9ypQsTQeM3Ao6JTBFPWH5oKIuGZXsX6LzNc
0gNOpc6XsrM7lL9iCFZ4tdSyOxZN4ywo635AfV0b2eeT+Fe9xzg3i71VzKxdHR3qjXVOPVT19x31
jVu01DN+B3UMqZsrvfvLoFErrqYTktxdIjqrSctIo2wJ75cbJNViyCMylPf/r0vP9lC3CJRdwn/+
JpKKh+bmeZuvgq5ogDEyJp6vfSG5o2498V6ZcrSoehZOUDZNPLstlG35+dX0PVscYebsGqTsBUQC
KHDF7AXNGHerQeYVB5DrshtWnO/fB98sr0HRqJCkxyM6llnMPuH/DAfZHmK/zvBg46ryMzOQvxW+
bmYyfgEYrniK2M+Wotmkn8DXh8Le57YUVMxVQBA7YlQdmMws3KCz/voGUIh2g30U+1o07KceBkmf
vJ6xymHyEYh71uzha1eDg3Sn1okE+mSw8qtojbJ0QUJHIrWWMJ4R/icafsz6f7WgYFkOqRc+M4bh
HbB0HpJcgRcex9UgY+UJYKyfZ8qSy29OIO2nxvmrQFxU8aV9Dv+GOyuzKfBLKzMbdygZWMiYrJ6N
X1DnBsKJsUBox+tXN12ktfSWmD56BKSWVblVr5vY4AfbT0RISQ6+uzgw+c98fMYpVTBjsP9xaUjg
iDZBnKudc3lKmXMbMXWVcVL6wS9TfXQjKKOzHOtogFvYncyzNAwFdQd+Nk4a76Gk+IGzJIKPGY3w
QWSIv1DGD3SaGxk5HZ07A8opkzxrDG1qjvTuvK4/c4GWzLmFkjnWmfgBPmFNAsERbZZVPRBGrdSK
PvawBj3CKmQGwZuPphmemPY1S8j0POcs8yRNiagMiN4MCNGESOSCD1ev9noOZScu61fA6QW7q9QD
T135nc50PgGQmeBlEhCC01BPF9Cb/nGOE+07mChblaF2+C0+wLEkpOGEvvh+2P0+Wl3kTN0QKO00
bIvqfAxp+aSSh9cWdCFTcKZZsc5Ct7pYjFEDUCSlc6Lujc5L2YfQi/q1Is5X5iHUNCPBzzf8bKsj
OnY5EAYQaxBSZvM1b5GtSqH6pCJiwhnKoStQZT11JsUWoVKWszferEu17QxnYVWsWFwDP8+/N5xW
qiha7xDGNEmA+WWjxSJ6ivvk5ObwIyz90m50FMKA5MT2X9e6K8dW3c/cf+x6G3XpDoXgvUE7ZBjN
PiqRdJZbD1ne6tmrEw9LjMJ5wjh0M8PNE4Trg4NyVp1a1i+gwTdkI4pqgKx9iDELQ/xrDdExyDX/
aDL2V1bRiEogqqyhadxgjq58t5dunx3D6WBCrxkGTqO8n9AfkXSmwCaESibgsmp90hlsLK8RcWOO
5F1K1N51WjHZ+iQGPajiI2dbK5Frmt+2zf8S+9XKFOH2PIpzpOcqnfRSR4tWjWb760BhlOAWeAOw
+uKou6BgR186tOZXzUttr/IfYbZhByzzYtI5woYsk+Jt6mmAuvFdepP4AUGdin4sGyEtZ0rMRh2k
3mc5rgHdbQHhPIYPR4mKtGFDKMScK7q2mOM8oMt1+M80bHe8gyCsJ/v9/dq2PZll6grxTX6iAMW5
ZqaOTywWeQPuNxkWnCbCjSWGabkbxQ7mXNSpGmg9eWblaCV6cI7mU245WMDnN+3xr1XXDv97YiWb
qyCqF6EM2YqgJKOYcDBiOGykOp5tsV9Jk2NQfvZUhhftbbeyahFpbBm2+2zvrUN01p+cWA1rC6UE
NtcUCuKUYRlcCd8gD51PDpUG7IW6MXwGHX6XKQoDKaSifcefIb2U+LqHtWJHByvicO/1QoKOqShi
UikauP8oNWMzr+faugOmyk+VOrvu87uTQqnktiVKY18ddj9yNZl43XrAuWERx99TwgfE1dDXMi1M
4BvdYn3NWe/Yw7vs8Ckyxh85nX2SLsNj0W3EjF6PgQ3aik7REfE6IsiWM35oDz6QWHhPJcv9DPe2
bVOR5IXpQa8yXoimYCle6GC2ZIgWQy0RMbDUF3YdjY6DdzpEMjZ4CNtMD3DrCqs7FCTvJQj23r7/
2JNfnW9REdKEbzwzThr7ob9Ge/Nz3qwoxxF3qjAIwRgqTFkS8Xc5Y+U6oz32fuEASfO/ooOatCC2
YX+0q929ipZAlnqgbqzWKZMEKPf8XT8gtXlgFHBxumpKrVl2QyZvdXhD4YbZ3gg/gXq6eW6u710x
K3b4pQddPYDa9y2YaIKlXBKg2LjsSF0TCT8Bukw2BYRsgeqT2PT3lxg14/9yoPvWw3VyuvmeXVTo
4x4qwGNZcz1PYwE/nK+b/082jaRCJenNIjAQjXb+QP/L2vEine3FE169usQCw/xsIOqqjd7r9OUm
4Cfp2DQZc62dtq/ktN100JgVgLwIQwwUjxE/mOdq4RqHlBWcf6PAJwOwHgb1fmzE7UCaBBE2G3D0
hp4cz51J93ACWV++GAP+npYJeKZ0HomMKyyG+rC6mwDtOXxa6O3p8zcW5UGLL+bWW5DzUDUACgdV
LYPMhIasfoxQ9yABeYJANpgyngb8I8Qw8s7qYvKiu8p17np3vsgxW9doeLVx3yO7yAwG5e1n8e6L
EfLGii4yoAlDbboiytAQlDg5mQU/C+igS4tttHX5bENkEcHuMHBC6H6QwL5iPl77FjoIC+FdYCXG
JZ1al/MZ8deneXZdhEe21mFYidA9pCsBPQJVYi4xF1A8NvIm2vwZfUbJUnE9MSRtOdC7WnE1BFUM
k0xLpuowvRhBbU0kGGbZAhulv/nF3SaYYYUzKQ99KmCSNZbzSc96bxVVorJ6oLRrE+z7DrFdwcdr
zp8kxhn8ETM6DSn21g7GztFrvkQfSXGWmSetyrhWuQ95wz1YR01FsIyWWhryAEi1AziLxRSljuXJ
/k5sELNeo6Jsp0WvCS3WqxFIqvok1GnabtWCwH1nwXNfRanwXHstZ8b1zj5fy2x9QOsWZ5M7OgEF
oqb17mAg+8vn6+KsAZ/dAx8P/IXyoXSNhhZUZD0Lv9NygYTaAZeMh8e2kWrhr9ooDSNPvaPyTEfZ
owZCQQNIGJ7hNY+X4yYkfw4CGB4ZX6ad2kJFSAxGncan4ltNd/IHLFC2L3/ouarCb3DjyrEL8uzP
b3qMFWelKIcFW8NihPg4cdzMd/wUrujEyKhTDw3sMiSQB+evBwaOXc5fGN77SnJtjRiQaDQDchdD
+5f6VZWLJkGUmqtLu41N49Dmpn3S39rqXdCbEtBXRcnbTkEs+h8o1KZM5YhMYf684bnOGUCoUOvk
f0rWuUhsAhFyzQtTDyqpjUwIY9aiPGn/L32tcwG9cW5OurUgFI7ztLCcYEST1+ZMG9QiWONIRbvn
cjNI2Sd0DjUYrIyfSfrVREmHDHq836P760PXvb6H/K6XyYjIxiFRDBYT+K5SO3PNOV+JiSdgKaZ4
U+Z74+RP4/mnUXizr2W6TllHd6bEL1fUppWSadwu6RoiGfbOJb6mVy9zzuuPKHSkGweQyam9LYcg
dw0PRHtojpliiti7h5RULszm1KfxFp9+W+Os8n5V8RrkhM+ZTOrA+965T9VhJSB0Pkxs5L9XFLva
JDkEfXCOZSGrErdkzjjZVSYQne54/tJcVtRwyu12IWIsmIkTDXB2iBdqRAWFh39TlYxrCtWviF3l
UVcycg+2r8CkqUjoT7dr15SrKEpKnU/tJp6HzyJvUu0QtH6Y91+qdIxXjvaCHlX5mTNv/G+EDMoA
q60qUYpjJSPhewzFoi5kg+WIQhI6WXAt6pW3DqG6YtSR/66c/zDJzj7y57slGA0ECcRQ/rfU3o1j
Tcv7CG12POu+rhBuAf2mPEBgRyTuMufSIE3t2j2tU3oTXtC3NFq0yEOcDevrJEcrgOJyAt5OUn0K
eon14hi3CZ2AJBT/qPQsfSHzsoE+SEmcGRGlqfPuQJpIjb+Wwbeh45cyHSOKe6YneVJjvrLesYhs
uSc5l8UmSN37xgsfz6mh07PNgj8Pc9SygCO0Dd5wWiCF9gUADFsiKLnIcqQoW5+U4zpHACrGJFs2
2uFdOSdKb9YLOdTERub0EY+f94A7mDzPl5TQkGb+8o3lSGcjojwXxt2WWT9NHcA4ANOz5fCwjW0J
FGGeA0eyBEo3YKsfvBuKgp4rJqNfeRGmPacTLQnMEnL678F8e03Pns9snljmxhvtVwI+OlZ0LZ4I
BaxyC73QKqRFCaXTkmzsjdbCZIlFWb4So3gt57DmpdtEzB8qVKk72YacbdG3vA2AvrFHI7An/iti
jueF02qY6aU+/X2gYPYtGqLfggoyMJn/EL0RzsWwWljc5CQPV6bTPZcRj40YEGMZDABAuw0Xw5lz
pWSAyPWshdb2d1OiZll5BOgFBQScWs/Z9QEICTB/erySzr1X/6AHW1lFxPH9cRHgF71v+HX8Behl
EA+dYcu6ZQn9OSv7UKyblHA07/lkzeQFixDhebVRCPfbgZRE9bBCaphNpqVnJm+I/wy2AzhrZjgD
DKlUBwLWnZQBnnsXMoRnR2aSGm6xIh1Rb6W4Ip5Pu8YlOPPV2laOCoPragTB62fzZcNOfgormy0N
hnYfbno1mFS4aJPYwWjajM7wuirAJXTYp6nNrrSW/wLr8+YwGv+PtuCYwxJwgU7yK84AywKAQGet
DWZ5D0QJCpc1G7ZrJNpSajt8LITMylhRVl+Zl7VeQOqXMS3Tn35/jFB54+dflxyhvmlzlhPxBFxy
d46BTlcCL/vKFgYPeeZ0l/7Qvw6XB6MggpAgi0nWzOcWHhz9p27iU9GjLl/BtLLbCqC/Y+vY6UfH
Djy/y0WhGMDOdDrgcDOTnkccZwglcpxaQkzyCjikpMvmEQ8AMUsuC5/Ne+rTYtOBXwgomr3qQZDw
8rrdAs+LqqySD7IlbhXlTcguO7O7a5iiTKD7tWuYX8SUMfC2ZYlgDsD2P93mqP5AS6zlRH1vxR+n
csqxZobnMDP6Y287wOfkrSj+negvW2BVHr/kO4z9CLUY6iXm7IwcGhCFExvaEtnJLUTMBO9TtRBw
UMRkpUqh3ziUm4SkSJhFTUUwzUwy8WcfP2hd5m2IJUoyVS+Dnejh3Vg4qQkPC8++Xaxjv2DlG9B7
1SD+yzr6EQiMLAzXAcXbgqBn7sVc1NqJ0Flpjplg+9homTCrh6vdSpSIkSjLZQcjUFclJNnwENZo
04MmfhIRZMDw0R+vmTMmQH4IdqkXwsejz93PRFuwDT1KirzxvG6mqun1goRf0qAuaM40MPhSQcxF
xwxUvnsrICtqXNeGW1eqWhCUlDeIt0qBUkrmDswMMvXxTsjOwkGkEmdKWspDp0ItvJg92QQL6rfA
sjuM2h7q00BcayP9OZQGBNGV4FaS6ayqcUSDIU+TRARI07CWV5IxvliG3+kg3aeKZHacfdFMNGIk
IeqZHOSnMd0szqrjMtYqxG1M8yihT49BQCwkHR/z4+MAvTaHZun8JhGM8qVUMBMoqDGcoqTHrOEf
jWpnlkKlQmuLUmX6pdfeDJusFcm4hoM3cU3qBFr4KmpJndKM85+wDaal2tX6MqbphEfK8f6hyDP6
cmIKjr8tpizJH8IL+Zm4LH1miyxyTUBmxHxp04+FflBla6+toj71e7SCBhsGCWAylrz5nNXg2Gt3
ZBJF0F3u8YmYih2J6uBUF2HlHvS0DighQpXNUuc2vdguGsvc1pJfbrFytCW7mlEWzk0+/+Kmo30g
0x0vALkflTjipvDqcLNAjga9jy1pGfadw/h+cztodk5AX+I5z10o+JNgm5nMnrtD/mZ1eH/QCwGF
EdNLJqO7AyCUt7NpposPtyAqSAZIYNsSAM6ALIPIUrLPlzAOIK3hyqjkU541k3no1fF3lePCtjKQ
/KDnwXJvbv56bW8QxawVcdRU/LP67v9Kja6bdssNYnzmwcoJa7tH6MxIUaLjlh5BIcePBqeKIVWu
PhyCIyZz2gDmYDkHgk01xwwHOxZVrWAMHRXyD90Cwt/xgPpK3wz2KNca2y8VZtIKLPsLdPDsZEhf
RqeqviT40RaYNPO6tBvbAkZ7HVmeB44qW8is35UeKPxl6zPRiFiUx4rmixEiDtGp3quNui6osiX/
YzSMC7YgrKFwUJmSp7A/40JMZtpZ3g71nYw2OilPYF+DPnFiuuPsHhDNDK7ug//3+wdJjI6Bk8N4
8TYwHfKVAk93Mq7tTFnCdcaubPgn2bnN/87tWvstBJkS8A/3obIsawkyx95kkUHoKk8C3L2PclPo
cKTQOWvtKTN1aB0zXH+gxmmd09C0aJ9Wg995iX2MzTu87HPS8vNM3fRCq5Z7D9H+ATL6at+S9iid
Jy0mELZ6hkNk7eEOR5pqnuzJbaruhm5Usasfis+7dAUR1S1YA90lFSvfC9MuyRnWuvOIzcITW3j/
QvSYYEWURbdYFeseJNxm3Wka8Vnc6HWsigrJVWkH5QQjWlfZv5Deh+Pvc4EMJwsefLy08TaBFbWG
+MUCi58pZyL7KNNSHBvgBGX8sG68C9DlAEo6e4X6I45tcLhS2Bgm4SJvy24n0n8H75A7sI7xfbq9
CvkCzd8ZvgSicQwRfQIkEF7TxYnxbV60edImUicQDkEbYnXLXbdGa+Ant4SKs1mrlJN5mju2djdX
t9MbkuGEOPdM/c4hBKsuR1ioE6CAV9FPiT83abrO74SFxWJ9dEbeAso/Q2/sMmc7nwQmOw2WcB8u
1Zq7h/eUexFIYK3UraFvdZwHjwYYhI6ULNcQReKuPrUigFAwcm1ac/qd3TO8GO6ATBWbSvD+Oks6
6SWSx6EFsJyB9mgUbca/SllNWlHGh2zu2hlZofXI/Zq61H2fOdF5SiUrklZZvCN9W32GGCszhCoY
1pilEiAkXrznbhxOhHGRKZoWmcPFTj3XECiNYdgXy7vjPgJmVNPM8C8tQoJwxzWLnCqCUjU5x8iz
oZJ3tzHfbc9M1jtGj4klC5mwo+R+7HN9H5a7qpZla1FXS3U5r6Z6O8MnYX4IPeaLaIq6IDwiRXPn
PPUEa36wiFmHt1lrYuyFhNLAC1VLtelRD5uFXHXu48ys4k0Fx8PqW5DiYtDFn8hmttmMNgA3ua1E
wWO5gsZSMHyPIU/l8bWNcyreqnU6uMLL6ZGRRXOj0Feet3BxWOo0xq1WA/N3xVyjsHRbf9pY9EeO
sPM5Uit2emOfu7qS7z8Bi+BGTUIynF0Gt2ieIBUQBzj0bELLweQDyWz1lK6eLNvcySYvyYp+S1jw
WaV+9FwjTbTItmI43P7ED2zqoN/1H7T0ctVYtcaRC63L3DSBC+64WbPQ1zSJON/aWZxTAkqxg4su
J9X222Cwt+hc6MXRojh+7FOr2/HCFHhqKs3WyU9EJ7nKLrW5X/vWjzWK5c1UACBoDM/Gl8TCujIV
fAH68/hSPasJ45dbWuVJeiO/1CzKNPZ5AL4dlzyrVWMT+59kH9UkQwgRiu/6JjZ/5H9pACdFs0nh
tsrSX+3sArhP23lGEAlbI1nRxLfQAgdQB0hlC9SPjXbHviF6K0/94nVgK1rJZpcXhQFewRfvnm4A
T1IFte/zajBrpaf4jymOLA+Prf8oSky7BJLNOHVOqz+53Vea4i8B5CsWBIXyeZwymu3YSZjNTeRb
TWGhUw/xhq/Zz2FGY1r0Bj+br6oIIyR6ioZbvMs+ostwrvJLsyyQTuZcQCc3niIwjLHWiN69sXsL
QOdNRbTu8ScUHnkDs13ZbSoz8EmfwW6S2bsevsXaGEa1NGcZcOYi3Z3z8WIXCgWP2jwa9vzBqtsn
+5vWEOQwq9OCQt51/X8RZk/TXl1uDvEKZCWMpS8f/ZKRsF3vgXG8wCre4ahZO8K4jO9XnJSg2fcH
qKQwyjaToc0YZV1OUtLYospAk9cZPd/XV7o3cNqlsqI8RYllr385xVyKnF/jrbPsKDRGswAGGvTF
3kgdyiixHEn5moInVEgheREMH61y+7lXiwA5VnX2KX2YO+77+pRuOKqqQXIacn74TxotF32+MBC2
ixaPjRMfzcINOgULr1bFOs2RlCqPrHTEojSxSitEDyaF6q8lLl96SAaXe2PA/c5U+sCTFljAv9aS
WrpEmPpBGGR+dsdDPUEV6t6yYWCV1N1yGV1PcupoVP2xHIu7URl2Eg+cmDIB3ORl/kvwRuAkR66u
Fzu+S8nzd0xTdeXeZOzv+vPrCso4sWmK3tp0VgiO5tqyId+dc734TxInks1zoA6q317GD4tfPgNU
qX4nZMLn5l7/o2BFH135RrZnzT2a5evRiIZWENfGen72P2ym0beYr8dQQPMBU4j4mMz6Bvd3hpRQ
Vofmgp/glxT8eMNEBjtsnCggFYw9Alj9vBVpBiht/oyiwmU+AXIrc/BNR0z50a4Ot1DEh4OoX5/r
vfe0zXG0XTV0K9ktNI+w5bzEH9ahDM+6+LFU4iUPnPmkAvKntwV2l/VR+7wPFH+v01Xf4phi5K79
YzWcS9c0Xv6ayruGfQyA5b+dazJGFUDsR62JV7O2C89yRHFRtvOta1wSAC7GzmFX92bsGHRtm4jR
UCqHhdmINV5epN/3x2iXscJpqiYk5z8P/gyyF/lGUVgegkdpWorCrFU7NaTlP9TBB+RIn6T7x8No
wRj7CpSRhhkg4PNJY2Q8GLA+y+3xK4AJSa+7xbRg2on0wEi3aoDTVte+y8RNvoerc/NXnJWCIZPT
uH7KAhnc6iQkCbCUDOigyR0qiUKPq9dYOC7uJWpo6AS0XNY0h+xiCQ/1q7DOPy0MYgwwKMAsqKRF
idqJZrZE3QJqWX6WTPx4XTha98R4w6A2m2nCi2BE6zATlBIlvd5YWOz3v1Uq+3boBmbHagzsdnwz
dogBmifI338hUScuNFmOjgEGnrrgKOjJa6RDiGd+UvnDcF0eNjXTxiajglE/R8D0uwVWCKrli11k
daEyCV6kKs67yCEij2yZ0T+eK0Ir2R/oZxee9m1HHFEBx54NI4WzbSftZLCMFJ1lPf7TWyzUr5+E
IfebHp+uS0wCrTQUQU/QAYAPE3WuhY/a6mwaeOavTSW4D2y8ck3lvWWJwGsD0n2hLjT7LqaAfNTV
0z007lQr6CPAVNrxLrLaydMaBpZrdhnleFq+HHj4Dpr/1TaVNdsv9l4cdrtatgXbZfi30VJ/oWN3
nXsPqx03253OhEEQMaK6lfmhOnxXIF4UtzF/RrL96ElHEjdjsnCwKEJmiPGuip7qHaHw23HWZXfr
Kk0/yCmr2UYYapulNkgJc573GVpSC03bBBgWsH/lgd1kfupT/l1+j46kqP2WRbXOoi0wBTxxGDxw
O3dQhzWF1Xcv/96vzE+1m87zwAd1ju/pN0mEt8kAAxjP9pYMCHcjNUNzJxG4kjtQGJr9HPf7V3Rg
YlzcMHOk58GfFj/ycyJ139aZjtixN8J71xfFdNK2pQD/DspH+GQ7iCUbDO8gEb7p9rZCykLIXIIz
2cC4xbg60x+TKvvJ5lZqVhCcFhzOq/tNEpoy4ApDZD+FJqVerSNsRz2jZfu+dIplgibOlbiovEmX
nIFqrGBeXopaVSDCvBsqW/gADyFzAg7IgPSr3SEFQqgBN2itPKN62/L1Vn78EGcw0Qk/822KSSBY
4BORlULs4yBHQT+GM75gma6wd8PuFn3zp/77lkA9vkWccjXK5DPFtugCYUfycBbU0XqVjhAv5HuS
ecMyWfoQtkNYLc8cNNTZB7qH7ZyVR90NwwfKbqZW8CVt+iXrcQrA3Ba7wQAcOkdiGoG1iBqCkGE1
nhydbczNnvX4qGCe73+KaZo39QPKwSEdBSVqGinWNR2aqsAcje4en/m9LZlftXoKz4H+IOvziFEC
8v6+QZ0nSdcFHyE/Rx2toeer0qvT/evvwx9AtqTJ1+442A7n7ZqTa2jao6Yk+LEpawXGG8N+OXnB
PEHuYmzcBiHsK4oEZtWYxBSiJGl04CJgGV/X2VH0Ar7SgSAz2voG/JebYNelaozekXzGdDFYNI6m
9e76uxD1lBCfqlXibJfrUWAxsATLX8SPmjqgUJ771YXHb9dKL8g7z5sz9r9+4tkrQ3Z60AYjg+wZ
Zu8cahcmsvEnF60bNussS3v2Iw3bTkaXA/YhwqtjsAeptJuRSwOo9gqKIiuKRWz0+05iKVxcmEdm
oYoVpf4PwuO28UgzDK9aRUNGHSUMCqFN38YGdu8OkmP4IRcuWPcm4Yf8tdxgoI8JDKD5GYNApJv1
p3nluHh/oq6A4OmyfFPKoCQz4EhoLLV2dLZnVU5yQ5InwPgzKaWlEJ8LX2hljtXreWu9ZnE4tvwj
b2lanYLUbrFbUgeYLuw2KHnbOrLW9NIAY/ibB8yXJJ4cIDIaNYPtdsfMZq72VdLrXhFoKzxHnHck
5+qUckMhCr2kEntGH2gDlSVGNEHbNrlRDs1S5UkY/cFX94yIuOFb89W7tDREyTn7+f9HlKN9W7+4
TH1wp2AZXQUI7uXIL4Fq7Tj4NzLkNItsKoEuFGnAfYCvnroAf5jERJjnVB27dqFBj1rTPLgSbwZ0
+D+j7voL56pqhr72PUNKd/DAELq4EhTq8SJml/Ss1q3CcJMLYhapDrKzpenblbfrIlhUUck1TsPK
VhIKcSOUpraociwRhYPOIpUMZGXqBZ3wMl1tk5owJT39sd8YkM8bpBlZwTtF4e7HWUJimV3Etmkc
WiFJSy+Ue6RtG8MN3urzATGUpS5SyqXycpkBHtYVm1JYqJSZ4Y06MJX1R0IXfySUBmgfY2oYkW+B
Ko0gSPC015UxghpFOR8FJIHT0a6tSYjKlz+QCVVybX2bBkSPSw6e+QapmrQNlk4WIQ3rPOXcUR16
ZdJKB0/i2z1QE9gv4/UW/p64IOeVObDx92Nhy9EMwEWc3buhuE1LFI8rvIwommcKKKo/gtV7JMjd
bz0Tv2zdGeMu0k8RHQXZIn2Yeux66K6/oHiK6GYhFJ1wAVFTYsOfJrDDgpANq4MadpCgrm0HNf3S
3E5tJ8HC85E5muvDGpD5CfYIxLibvWKw3vlDcGVUOXd8//k0gB7bm881+K8awiaE60e0wJSq2J8K
jv4j4YcTlpV+SifJ8Uo4a8C5LetBD2n9m80c9Kfnv2QJUUFNDzizR5cA5Kmbr3m5A07VoZQseMM/
STzmjAK8aKob7daUB3KuwJa/AxhlPARnuYKHRonacPDTKpgW4mRtRAhmhPVav+f6PiQ1uONpqJHz
lUHvARACIeMahTEHm2joTIz1OuWL6mu+Vg3snMVJ9CSYxwyJSvo5WE6yNC7pP6EIXJbyX/d/PgLU
qAKawr4cXWYQ9GDFhCqUIKtyvIs1da7lpsitgGAj9RBwa835/ZtiniZsILBXDQ9625aTbW42+80j
A29yf1qoQVwSVCJTagkSF3IvMhyrBgCrr/i2zk4FB8ytWjlh5Jg4aoQg/hLNnFYvZNrCMiUCDIqA
Oc0heSdtcShEgVMYfq4DtI6XkvUoUDMLF/grcE9LD43iF6izuW8NHeygPyZeOAy3t5/Ci5ccZ/1m
p3rlgGoOkaiG1iJca9sjPOJNP9Uq5R3eBWkUOVA5e+E/neThgsOmsXtJFQ4jrlli30XLWk+RNcln
i49ENVAfQelFlS8vOaUd/LwsvgnNiFpOOh90zNFsxdQ9hT7bBCZqbcWnqKPLYEIa8fjMnLCPInLs
8SybhsTdLqBL0gSyYBT6qvimn5GAUZw/dkWKNU6lJdXb+0UXUaCBlIDSvjrnSH8cAVcfXeD3Oqfo
Sk22iFjAn0TctiDY24rcim3mX8mSjwA/K9pDucj7SeHwd69lCcgE8HUPzEiW8AMXRmJ2/GxLPsaE
Qpmh4niyIlloXD8fTaJ0tAogJ/X4W7gqx2t6+I4195QJwPix7/dU6EWlhgw3OJSg3PugEltl7iQF
h2vOe8k7GBSZ4pesBSSa6sS731buK9ZAF+kf0UOADDnjIvTaK0AP1LRXJQ0FmqxplaRHmJJJO6BV
wPAuVerFsiNTz/e1aLsWzAjsXUDSTmYLQbkiPp4/diC7WmrfRiukeWjiJMIkUwL0zhes47NAb9o4
rv6IH4TL2y8pJl/Br1E9ep09xJmXowePT3FfnFHVTDmIuzOJ9KMOZaQR9w3dx5UHDHqCYO6AO03b
qUBWv45KVjBbEN77SMFFw4VijcecJdioQBnGcjCxY2EyQItB+Md/9EtGagceN8uoMrEY/utSZXSE
lwXwdX2vPt2VJl0j9KbQxeMu/a2PV3Svukmr8K0pb0CH2pvXcdLcNRRL07IBe0jwm8+8I43Us8i+
7N0qYl+l1ZLv/PFI0rKFAsssxx5+hK9CJ4qiN8W/SflGYmCt1+p830muOYnM0iDTYN0bDgnaeBlQ
VdWUee5m9/Zdq07WSk0cFYHOF7eBGeTzNDhnEodNAawK1/dHKuvfWk/P25RXuXWZVuPBUJdB0leE
soKOCQfCQNsBni6wvdbuyQQXMy/VYu+p38c/v9Y1KZIlxXSxyugUd5Fg1Sc50VI2H5qgphXQ6U3h
FosVO0SxHg/h2ZkZEYt/Ajak+qL6SOWTo4ZZ1EbBmLFsEP4pWZbplUqwZbAlykBtrB5Kvlac3+eT
KziT/TGMdnay9fWYNO+xFwNhZXbtuTEAQPAJc1oXsT9MWJ2zyINIfis59UcnZLrg7vJlsyiwWyGD
EqGUqmacJnva7w6t7j4xPwgI9dYmJtazIoj5BEhALVpGxPt2HrEIZJsX+LCnctM3FBjCnnWVOXnv
m+IgE2fu6TT3FQoLEGl5gFixw4fyQJthDXu5PN9VmD9489xhneOv2SfWni9lfP7t14BWxDW85wyx
SLaODTnfPJe4DWFFRmBMcU0j/Dh5FHLrbA7raZ99nlOykCCNyHaVdTVwLVp+6sKurp6GaKdgzLby
4kpFs4o4COlia8PIrvO/3GATLBhQKcWcUfDFs0qm0INUF+hK5R942YRhmRgGkpBCCnRlOwIvKoLh
FhkP75o1V8b1knRC6ftow4KKIjee98Ijt2la/N1kEZDlnj0uvk+/GRXE/DM5aPGh743rVeHvgVdX
NVXkcYDJdtUsuEgWC0gZvaKwSMteqEOkQ48FLRuOvCTftOk+y3BEoskKGzNFA15FoqF2duxTvv9S
GKTgG9lC83P5l939ZR5xqPbJCqdBZX+zX0XVH78Q1Kw0d9+CNVFwqKIj2PMaIH8LRQE3smMmQwwx
SsMWfrGfj3zWQ/KQahHm0wOSu7FgXjjQN5cnd8auWztUxEzFQ/1U5vDHKyv9yVvgtPgik5ZR4HUL
iTt7K0uRgc4zydAOWBqXOlOlvr9B/cGDfWIv+m08qyW2cZ/4ztQhvyYVd1ZYzyvpP349wV949SCL
b8AKUrHqt+3J/Trgoqx9YyLYzCAzF5mQt7pc6DOPoteephuTX1aPZEb5GfCetASv34BkfvMr1fOY
NxzazRdV9+i3X+yoNgozVf6zA8hL5QwwRZXIKlhJj/mAI/ZDwQeE2+szNyQaIT5COAilVSb53ZQ5
mRicq7ULJIS+RLdKRIpU/U0O3OLFkIYSCpS4Sge1tJT/F3gCC8zf04O7+8JCdamFT/ASmEHhzX8a
Phhdp3Ji6ZqG1Pvlo7sJPSb3nzSUtHpKQpWvznA5M1MJTJtKpAGidV/F5diYDtt2wEJZ02c68fRS
jhsEgnknbl0Eb2MojL2ACKF+G+LYCf9ZkQlAxYXy1TLGSD9RfdwAM1JH7UIADv5/tbp7bo8d+Kt/
W7clZd0pgeumZ6mOJQfVK2AKfU3E+lGMbPvqx/uE68J2lBjK+aWm/us45HloGpPcCYNyFRxVUrsT
1UdJPT98HtMqpxrZ38Na0lkOz5RQIN+L5r4rD1yEPVC0wMk6ncnQpCrNQ4liVaYmcWZXLShFitDl
4fxjPZD6bN8CSU4+fLKOIozqVgV7ZnlEn1D01rxaVmVe+ERdcjAWg9pv3WKzq9hxw7/OCZ/Es270
DRRVs0dalNIszHpJm19eQYcB53V4b5Dam6y//j/ay/RQdGZbSBMcJWoaW6nAhBEUKQPmrZ2E8K0l
Qw+UUFfvnii+eaC4oog7K4GBw+1I0q2kvb4PTuKYICJXl6WD5pX5EHvIO8zWQhE5l1omV2KgLn2W
T8BlyOBzjBpHnQWkSyXAekDLcRRByB8DQII9LsebpR3FqPrdSyhanmdmC6rKeNsLoABo94NwR3dm
eYaddfkGalJjOeh9KMQ+kg1XMl1/X3bG3wlE8dgn7SMcx/yJ37QiG7LWcPukITx88pOT3khqVPVL
vFfDgg86myHD1S3DjDJ+SEAStNpcginXVBt487gnQy0nO4kTdHRGm7IWqSfCsv3+ZayoFa5+Juxd
MpxH06DemnTllpq12A2w1rZH2jGZ7K9Ly4Yig1ZQXLublyAkXyFsKugjEVGaaZ3wOC1oQ3FXW8FV
M9J22prwp1narL0CYKSe/CvfZCzoA0Dmx3Xkg4FMW7p7pntWdWdD8aaixvTVHzJQXVvWpai+dQQ3
00EUuGADyUInouj+vXm4w34vDeV1xbrTheLQ5gUyuo7aOjE6qCMKgf+RYrAAzHwdlTyqk4kMKAOf
86PmHsruL+zOx66D3oEGFJjL/NGq7m/TrhXzkunevMXmq2b+sA/hCwE2qtNpQXEzrMe0n+kYjM72
xTvShkqTvmP3bOfZHAVDJ/jpreYCfQRD+rW47TsO0/oiFN5NM6IXmQKSW2UXFkZNwblckxLdAly9
7O0PjjwVW6faHQiJZY7AMlnH3stNQzX8jy69T2YaeNPqVFsbymGPqEsBpr3NjcEmJ1AqznEBbz/B
eDMW4XRf89UM5jSaLKt7y6Vl8BlymPGkrfU+XmSe5yF2+W48zniPrFITNA9tn4gQ8hXPvPdJW/n+
bXIxTRcS5Hu9utoNHNHlLaD5mgADjmx75jAg/MG3EDo1nE01AtEy+0fGh1qf45ccG8YLDtaKB18z
b6xOrkuKJSmHkRk42USP9iT1gM28BOxNwwPJl7zY6Y+XC4zQU5KC1ZPc2QpUpQpN5GOtefdXVOXP
ZXgSpiW8w30dQv6cvttpEckaaxsmT/scjNvdbA7G6tgqJn0RO+yEZDW+yiUws7t8axZs/VI9Va4h
emKZveftl/b/Yj3JTRJTgKaj7l39eZ7bdLQstq+EcLwjF5muJKR1ny0Sp/qZPN3T4cM8zjB8AXBh
VP0pyD5iGNNi9u4BsMuVh3ewbpvxrUx1htwjSjR430e5secSPnfrErF8DwgfGNfuA6WixdjFqmpL
ARvOcrb7XsS2keESPU9rQP8j+B5rW3e6v++uaPv0Rdk1ss8yoAOP5YDC3k5XaLC2Oe8jEX232Am+
vm4kZIeMAa+TlRdY9Iw4SuehCWoJOAl15XtekNLQ/9aeYOIjlamrUK6eZ0vQV698N+cK7rZS77t/
ziQkNZv4ksaf58ZdOtZGWHkkMC/bjnd2i7lEMp7gY52807D+mKSeLbqcjDoWqByOJ1ifjVrEHuBW
VZ0aXRIv3cFFxOeQXEFxfmAujS+BDmMZMHUlMG3Ls5C3tZI+0Pg1NtXuZWyhth8Q0xkTjmtYtqF/
uYWA4+Bw7lq4n4b6XGqO+Y3FwVzUdIMjd070RVVupHQSfg3cvodSFkUuZDK9/H0LUd2OJIQwh+JD
6qVt10FhogMwUEJlVP/CwN4h02MSW8+0rCCOTZ/YsCa1P+pJvFwjQcfQp5CXeGlPpwqVxaAvsafH
NpUM25QLaGimmqBfYcAOotjBuML5UQe3O3T6eItcTHYTOfsXjP6oo8la1Y8BCYA9OaOSjjP06duk
7WPJDhTMRWhRE1rz5beS8qi9TANFNfkKmNnRbuDd0TkfNq6Ibr4cnm+qBocnfN9/bp69NSrxNzMl
FYXTmPRJFla0iiWf/wSQ6si/8nWm6p88I8gTB4tME7qa582mLGeQWZuzAQdKdgp09fzoQ+PhpBhQ
Qm1JNpDXSnliiAdncrF2WRH2ruq8wLQ9kzYd9OuGGIc6Rph/fIwxnrzTL5m4+RnV2CZzOMEinNj5
+GNhwS5g4ItdKfELG3C6fawf9wXrAzMruGxuxxFtXEiorbMW55sAkzAP3j0lw/ApioD7EmQjrG7P
NC1DnQrzMYfTU47dphDUlzpsVMRnx5W8OViFqI9rCWyeb6luBpG2KbSLfYamZhWrF1TvfCg2Yrze
lj+3X2WWTw3bfR59KjtVAYliRlr8Is+tz8vXajcpA8ELnWuoWndh0Oou+RJJsBVxUrX3N8RvBI1X
vrAb+CJJl1ARjlmygQyh7jk/0wvoYdkll9zoSOFu+0ViQdFsDYpWSUeaKQE053DwWJKMo7ae/lwd
O/7S/g93aUkLRQvN+5NowdAAR0qzW/mdcw7rOrm4dhrvIMBXU4KeyeKmMCHoe7holbAvb/N3lZ/c
aV9KrPaVhexGVJSPhu5qbO0Bqz/D3YuiAjQmpSCdIUxixMKJ+Bef2ASRe/XrSxy2+7uXt+k5JjFT
VD5L7bWcu1S9q0GKIGQIDHtV08EIKK7Y0NapK/0hfl1wfOHe3D9N+DmKxeBKwpfhp0efy+vw6I9x
eHfUmugEa61nHkLS+B4kySe+lJVqQ8r+K8+X/z45BJrSpFbTL4TDdGXzTbsxlaHgDbXk16trf78a
PzFi+BgvwzZX2n/L67c66ANLj3e9xqTHVW/nv6rpjCF91StypaOoq+CCgyIqQ4SDzwW+jUdsedUN
5TEBiamq9ZqApSt6mWy5z4DaQdEVXCWzo3uYitg1UHU2l9jBfLMlBatQeN9q5YES8foR/F3LVS3Z
Vfbn25DPLRlqrwOd+E/9c0dM/Xk5uKwrDA1ohbZzcUvurjQt8tjm9r4hNDY1L5BTOc7wbs+UcGAT
gpDkXXPauJJnraq7ymccslLIEnS65o94inSmwV3VYoFa2CnYDBx8mWj8nFEu9MbggUYeeA92TN8T
8joJbtaLvhW/abW7mN/jlO3F2JW7FMmJixd7ChWR/OUg2am4gPkUvhwDFfTD2WH95Ztvaaq4a6xN
OsBz5MMQnmcxqU5CwGzjlK6kox8gFFa3yuwluvhvF2yIQyySv5n2n5z594SaR/MLvs5gaa+YAfHT
z/od2AGR8l96OkjmE9ZNtHB4YvzxQ9nVBgQtg1zBJ2pcbCUx8bqBy15DxbEbPLY3DX4U4dXPlVUT
YWTSFdOafeypj6grTGHZxEkPKdb+gtzd3Q4OzaC2Zhfn0t3Zkikpi5Rbm268eXwSAKHbdiifTpXr
C5CHs5Fa/aSMXXpRct6M37z2itr/GTANA+5gbFpOCF0yfSIbr+lG6JmkAmyQKPuDWi8wKBB0WoWI
EiBvw/je6SVOCFFd+XK8qTJOFD7tBahC+QyRYO+DLeKmbcubS/ioD80h/KkeLYwBfFhaga0V5lWG
XtgGLHFcORMg99tjqFz0Y5OZLJbssil8lzDOzc5VUd5Nt//BixD1vNokNNbYv522s/K5ZiXiDKep
QS7qEprneER0xQ9TypUaY77fkRkmC9iA/VUrm+zNahYqz2LGZA5vb1dmtF8Mt6WnsqRwl+oW09pA
+Bf56ZCdDfEGxVAwdCbLT2W9y3TkzWSlfLqNiMxnl/VBswDAt/KiogUPMLdMPTNcV2OA2vsNx9fA
qxJSkoV0CBUe777M5N/voxKM2S5DG+mo9i/VBfyXSZ5xQ7tkHTWy/TKfVWi+osevyRusKBDtOEWv
EbHZZB2922EUsw1vwhTc7tB4HHAjG1Q3J6v0c0/SF+amFBRRQYpeWsZbC1A+wNQsc3jUCKOpv7UI
1jkedS76nqoJ4JduS+YYx497KjSUDnR7wWieyMlzUKyJvxla7EDd0vKUdY8PuVZCAhhb8V7L5BHM
JKZ8A8khcV4HpuSPFvJ2hnYK+hFxzWTvL/oi6DOoP6VOeCetgfASvHeo3yUR9J5cmPX1lRyin7F3
xycr8MezyWJRwqratbPtW+DeBF5q3Wg5D6PIU92H/W2Xuc7PqskqDDF0KxJ/0TmxNI5hVBwPl0MH
O17N/83ARnYwHj8iV7DkGwEjGHz2Ayhm+2PaN0UV+Ybvw0Foqh1cGlGHejG2RraTcPFsoHVsKwg7
Ri8Wq4aJk7tmOC7x41Rp12slKtrB3dNh7Kl3GLM5f/OGw6jDFx+KH7yFkCo7U+qLr+0Ref3EQ26u
myMpXsVkAFXVPBaYYPjM2Wze26vFh8GnX9hfC5BjWzN6rEuoTT+Jole8Y2cBEIRzGzX+AtIcZ3d6
c5PzvKEwqFbHQPycUKHfvwbKMdUS98Kzelf74ZhNyY30p4MMD2Q4O2nB3h+33UaoahKDxqFSrccA
+33Mhkdae+Xb2DJVuK9Ka+LfpaacOnq48v4lpd+tCQhv66IOV0N+A2R6BA3iFMbsmOQYFbMzBr9R
UFz/bBqjDFS23YC8ZQod5O5QvkSyE22gru+oUEJ1AFT0sEjcKYDsDeZ0E4l8I9G362ErKUQnCC4q
hBSwj96qqLCaVsQLDR7WsbJYCgzGRPARrgcpxdzSVbtS1+3B7AAp1r+bwfk3HXIYq/f5OU5a+yg6
EDkpGWtBCGc0Um+SNfJ9Jjy2KuQmQ97BInqRbqPOv4U7/izWf0qC/YThGoBZnHNmkcfZOJ5Yg0PG
0K+UlSecZH5a6ae1gF+R41YAlQIJLo3pxgR5OhMVjk16AZqpR8sAYL3YQG2hIGXqYW4Aw0S0lyBp
3AFZsK2WT18wAabssMXkNkciOPy/HXw7z6LjoMo918X6INF6yAE+bnJxuIQ7LanYe84H5mZ268ut
UmxRfe0AZF6xsUTvQBp7XBmi2wM5CeI2UaDyFk5nklPTxZUQZov92Yj/k4bU3GyqYEbejl5u3o3Z
RDNWYYH0SROVuW7jSna31W5jOtYDA1zjyMzhsgzYf/pJ11Oo4diHePpcwSvEH1seVJTxpT9Bw1mV
tYbRi1xnTg32VRz+AUdfPM5WlseaBMTKzl9nr/rLm+MVNBIrJ0AqWOde33k9B/YrE+xPr4+sLkIe
v74y9PtsnyBQVerzu9t0Wz7HKiQ+CjXcAa55xrmsnKfTK4TMu9XXXpOLxdWq23aUXzbcY6pHGWNY
Paw38YKmnprZZl/jgT9dw1+v72wRAt1ocPu78cFDPkRBRueguQHN96L6ZL046Zl0OJIS58LXQmP0
oonbGwnOR27HLRNv0lj1FrzII73CgmomMp3zgJcznCg34x5jFuMzdCeibc9LTE+FXHLTcpoHj/Od
hQxhLDvYweCpqbUhTN3EyKcWlEI1TqJrYC6f+1Ij+R77Acem7qZeFX67g1dYoqpUq0RDi6J81uiW
C1uxR+49ViSKgcecibRTNzkhP8NPyn3/c71pAmg5QZU2dTKdMdAaL6Kg7slRq+6ncAIc1vFZd6hg
HeAdJ7cjma25wD52E2fDXh1hemuHPi9N2JyzfDpUG4kSHD2rDz5wKlFErjG16lhZfpWvLGRlXa01
tNQiEqmEcFZlf4BGIxpqcXWoqPvdDutqEGB0kgBU/uF2c/efEQBTQZt1YGIfpJuXM+2giRW0CiiQ
mTS+Ye9sY+HBgHbhJkSBokIYm+RGq6kI/9Ma86p+Fu4ugEKzw8bjTIndYU8+51EJzVhwG9o8LurO
xzZUIXe2KsXGRe/Azx5bhNXqxICt2tGoC5OJAVMg/Th3kxpjVbXPl3lFObBdJ0PRzvCWpZVIb8GK
Zplxk/Hus1u6nX8R3nfKN28dV4oT8EMYaUbKDNxDVr9A5Fo6Afm+2GiWTbOp1chOtORf/R3lbBxM
rpg8lxoCxeI2JknUbU8WSFU8Z9VvNh5PNDaX2LfKv6bMV405602pir93OUok5XO3GVj/TuDYvER+
uWO5Oe4WDrBJktpc1CJ6bXlYxCD0SC6BhuhvSl/PnDkZ6vFOzfQLkG8Ujw6vzUp74KDAvPjv8mnC
GkSi9VdGU1fRwwbBoFr7XYRjGLxtfV3iXkwlqOmz5aXFvYqYsWHF6QWgmd6+eoM+412gc2NGxQdR
z/o5Lk2LjySStc2UYAvAlapb6QVkjQ+lNLoAFVl4oEWfqfU02p6LCW0xB6l5gTMWfkAOw9jLA8DP
7NA4p08NVmGxP6Z6fYTcNf+f1HSxjcnzi0GOg00+BIBWgRsI2rNu+Qc3ZHeV42F1VTxQ9aSmc2+n
RucHfoN4XiCTMhQ4PT8wAFJTKs0yc1roq8DWFMsEJISSSoOI8vlNlGdcU8Ksr8arqOCVZUnQxfam
sO7pLNDr7UfYojlYM5T3qay4xf7XRV9PhnF6fTfjd+NnaPljZVU7HJqHT6U+jfe5oKeJO0/ziIS0
Ii/BLnw+grOutZmELgvkfLEGnSfPSBNTW/H+PT3ZifoBatoeClGP9yuOS/97FRxU7/S0wR5tfdKb
DXRFdLe3emW4brtGa7uq9omyxrGSYYfv8vdj8XCa1ZS4rZkBz5UsRIJ33l1EBKrfHF9NOisinujM
c8cS6vbVPgBctDOdlbSJjfJkef8rYUmbLqMa4xPPoRQ7uN9dKGIB+kX7uatlemQvTVlzK97kUkvZ
2ewxV4lgsYsq8txrh4FLzHzOG5hkwMeZbxy/V+hSxhWX8f3/KPmSLr8vZeqcAzvwuDcJ4Kqd+r5L
HDDGCXhCmbKLcrl5V3isyI/QUJ1wMeR3iYMFQbEwQ95C6s/A1CpVn9wgrRLlxnDLrPqCEJ9zOV3G
NlhmcMubpuc3BoC9C53BK7zAvzSPKFMUG8QvbhQeDi3FRhTxXS1p13YKGbuqCdb3aSX+tGrd1GAQ
gh4NWL2rYmvvBc7RTfuZqyyty8fBHgrmwYGigSDftidnL8Rnug4O1k/C5ju0bfLtyzJQK6HK3Wmi
C1Y5/mi/2BqO15QM2qSdziVA9h8wTsx/fcrfooG1lBNBymHbhLsu9/ejY+EhR2b0kolzYIvZKu8I
rA12nfYLXHyLtZ2aj5Vw3XjSHdnHoHoDopYpfHxowZpMcN+7BaBJe5yNUKNHlgyN8t7BMGgB163H
2f4mVDHbU8iZ5i0ybr+LpgYFxT2zhMb9yzQoAYfMNJnrMBQgx3bdHj9hTOW0dTPmMmqYENsOhVU/
j2lz46eUfaDNDbByqAYtv4VacIOFAFQcWHyyVcl41TT12MoHyHo9C+cMoK/2jKahiV6posD1NUvh
sr/uSfL3ciwBHP4WYk5W/Lfu+45PNsDQsCBAFTaUzJdzGsfCsl5YUAJVFp9SLNeOhgU7NWOAFNsA
BeF6eUhI6cXuXAsy7BavSaJK+OQkiW06DAjnQDB2fXgFpj8Cuz64eMzIMKdClVOAisGfqiQ93I1Q
H10/BOp6XBvLAA7k3ly0KxL/D2f9JYg/g9ThPcaP6WOkqxWGGGDTBJ/XfxCjczLfkyeLZJAtac+Y
ukniloQQWC5coywxg8l3eSMS+7o+se7pYQ3+AebE0NELw8nJRV6zAKaokGSYqMaIHC5AULWgLQgw
+gXM6Xg7oF35gvJwvCL0UHEuL1kI6Nz2StdDhO7HhUj0JnfCN8CLGZVV0Tee0pI0Sh8U16YEoQpI
gEzMNrhTj8VQRRRinPK6oRjfhbKQVkXj0BwqNfhvwwxpQPWSNltl5v8oBHu4Dp6uwqWR11HarcvJ
aj0MzFYcY1h+TMc/iS3L3skfGhx57FCQfavDcEGRdYgHjqrgAWgWo8/JLRIzNJTyMGENk3hktjVi
cfaZ9iu500VNCMnHXr3rDGFjwice4lE5ijxew5eduOqP9CFhMZZDxqBZtOQN9SDYQATOLipw1fqf
3REXbyf10J4gY/qdTe8L+AIK+Cyvwz4UcsyIiKFJCrQ/4uYSapY5Fy7FzjUCKgw9hzNS2BIEVNqi
TifVp9ikJeReCN0Sflu18iTeSJOVDTreSu7I3Pr8LEclhvvHEjTKR/BSWWB3TMVuadfzgDnC7AXl
JZtHc15Rb5viDrbp68bfwweklNpJWf67VLrO5Jd8Sv6HBIs3E/WTokF/uFFDNGhIkyTpsAx6lLny
eyyUBhh8B/GjvSw/zfF7c4tQpR+ot8AbcEssRbzuZNDk+g9vsP2jTEh+1Zvequ4LsSfQisYL7FQb
kJ1pUmZ24DFjfVhCYOmhlo4J1/xxoM4XDLQoL31RX13Ur9YPSNOJ4JPVmtz53oOUvYGWXXfQ1R5O
CFiTU6xQnpdIDYY3xltLvNoKeUItn01kZosmpiU2LF2j2AwwDAeEZh2lZsyc+2r7cG/su2j9xsD9
QowR5ka0ysLwaDy6prRmciY1YjNqtNtGN2X/TldRuFS1oa/nzw9DYxakx9hlRbK7RYz3D0kN/f2h
lu03lTiIy/Mlrl17Qrj4DlcxtkMoyqx2pYfEkovz23ADAYksoN6HYExuSd5d/cK2DEB2ZCkRBp4b
C/lfIzkfRUJBQkX8phUCkD1BoU4wW6ekLZbeU3JeHhNrWuciQEhKUCGcV4nEa7PlqDrySTxTPwAr
tzSUAnHpcgA2LuG6LqYY2FuW1HLzKWCvfnQqFloF3JW7lO4thPFS62uIFKr2jyLTTxDe+TemFroM
/qkRovwET5mkJnA8UMmnqH0OVQS0RKR+4/zPXvl7KjR0KqwzDLPhuG6qCOIpocSfCb9Nt912w5MI
/aoDBulUCFon/x798IAf7IdOfEqTTWTeIWdPivhPbmGf2GHkohpx0ltbTyqWcEz9qVGMNVlrqx7E
wL6OaWxE3DDWKHylqlhbMnBSdb5KaWZCo6IxDdXYP/2BJM4mkMokgAEbcdNBintBQbTe95j0vCox
UAkn69iI9FjBgUID137aqyzzbF8JdEtCUS7XFvXg/DUCQ9imoSRBsOdrdXUOUiSCMj3s8wfB5Ref
IRNECEZF7GP2RzyqgQ7ZHRe7QJqAfCi9cUGooC9cn3Gheg83Ox+Qk2h3hnmOagAXMSPE/PLe9Sq7
f/F4zKBGLz6nVJdh5ny6iQqsMblq1G4kxzPcxSJ04JvrwCDfFG7YGPAjQv70/IicS0WGgcu/W2i7
KklxKgg1qvjXPv6QK5oqxfTx5ofEMSQ60dx3dr5I53pgyvnM+6lP3VH1UD4aBP+O8dee7WHpTf4w
dSrDDgDlDVt717tKjTaQMSryp9A/r3rwIo1Qh8ggh5OrZ/roif2ccWnt5RpajzG7mX5DQKeiw1bp
4ekRv7Ftnq7fMWCXQIMjxnjqm18R2UQMZTOY3u7nkXeySIve1wkVg+ubIm/f86ZAHZhb+6x+gMlj
3NmzyoFCquEwJZUksIcSeT6bSCArLmz91+hqx5ZEY+Wj/yuboqwlZpUZHLjPBzw8dzvdvXDA8Hf2
/oSp6+LFILZYP7xLKw0NtIjeypCazW3rIx6y9+AY4UdNwsnX9TGp8Vi9P3SK+90hsB5UOp9klfSy
wOAPmnxQVc40MlR5yFylKnY+PGqPfFqBhx+2I77BCyDWaUBRcBZM2JheNlTe588dJPcFmJzpX8i6
F1gxpWfuFqThNOZnbr8eQmHNr0wIB+xJqu7KM+VZwafjxt+4Zckuh3BtfBz81KNLQAbNxSxt6v9c
uUgmUBcAN+NQiI3Uq2bViY7GZMhEVXIhv2tdhgUnjVKX7Y/LYqBzOX5J7dS/VMTM8xs4HOBY3OKI
YUo1R8vv1/eKEaFAxiHYeLOMYI92d76EvyhaDNYw55cX49YzoXxT3HJmcx45d7RxXZOA257otwsy
X/7a/jz5eo/xLHIqqqwJm58PDtOHL7N/qxGeFj4eHbiaf+B7DICG8qzM2+stgneuuG/bLj5qw9JM
PHq1w4vPqPi2kPyDeP044pei/Uq4q17X0U1jjQeFy0k29K8FFB0rwUTvNLptuPD6XFP5GCB2DRaR
3+Bz0qPTKnDN/4avRUPUj2bvAAyL54Oguynq2Lv3im+zh/gGES32zfKP1h4uBk+AdT46qx3mUPgl
LT1rCe2a1cYO876T4u/DIdpDzu2X/4TJn3rKlskts9bjw9q27qf3ogoapOxiiLH2u+13+IYtBWbi
S7rtkrJMe8h7hVU2evp9vsgu/HsDZ9VLpV40b/XQsGHj3prPyjmZpXcrx+XTI0zQt8plwh3q1iAs
Vx96/3mXuaaz1hell+/G6MDhJWOV/7EU2U0SbCV5no/4D+BvK4uyK/3puihPgUON8Qr6QkvdJytn
PbOonwRjC2wZ2oRcJ/E0VH1sMUcbHhB392n7oic+n/2YYQMyd+lj4AuaOazvTbNtnN8i6oqT5+Xe
zL+KXG3h7IQjYKRTeHzJNOE0boz7kb9sDnIZ4qq/nszMVlBwF7bb3+dKIGMRkoYZSqOzEam91MF8
NB3OwyYPMhXUQnRAoSzNKA63qC5kcN2q+PhN+cHgvzNCuDzwMYyKGdfdOfMBrM1N8fQJOXzTFkAq
e9TG6grjonnbR/7rIOAFL3PNma6S2yS0G3SMxRWcgne6oC+y8JGufIE0HfDcgL4j9Nmhg2IyhV8T
B/ig6EfWwgUUsFs6ikuU7HBAmTBt8oNTkGu07fKSirCVFgvnkwnhKH1YkjudF0hHRjfX5Y3X2t/M
+uRmGRP1lmPs8JoBvAC24BC5I7hwxr6Q832Ni4Dtlwq+2W+OyMbiJpcgptVu0d8gGzwm/MN/nKgj
j5jSDzCCc8ZZuUJdGwdjiFksftlYrdXkC+9d6u6x0JXtSollBMGLaVIvd4AbV17e1JL+ZhFOJz10
Po1UQ7ecqO94qGckCROVY9ccyxWex0iZmlAJ1iEutWDjBqyfPvVJNyE4DEQuJm+A8nClxHyrkU1m
Fbv2zSc5smsGwJl3YT1iooS0cE8WAm/VnRMvkPstmNBeKvu2k+toJ1/6eQgcFCTBEaZS1TXeQHzg
3ZZHOiB0q1DnBOIJNmFdX1lBQONYL+8AnQTlSlaoASLK6e7/U3HuT38tybAT6E3ZEGIHFFcImNVN
9U9GoDxnGkG8PN0kygexP5P8uVkepTpmKkXowxcz0wg7eQr1oiARNo1zGWDI6Hf15iz0N8SqMlcQ
yUmGgjdgO1TNND6HzWBrsWEey0SZU9IF277UHfstguLKc7XeezdJ+EiwUFmRdnkcdpwKjXI3avMF
ryJTkJjGODOU7/jecLnSiMrDAQspA72in1b4OUC5dLOy8FcWnre3a8dKy6k43teLsxiH3xaZv6Ps
uSoFJTK4SJvpITcN2lH7amSy6BbPnAxKzujtZqqCOWwIHPJ/FEUpRGYsr+Fc3AfVimtorv78ScEc
Ly56FbRZo0G7WqVngwo2INlOfqQLiJZ+2+brAEIWkk4P4BxYW5mUetK1q6C86yFYt6gwE8QLHSHW
YX2D8+NGGzi+tLHywDo119QB26ICGxZmItJAov+HXoy7c/GabzRPTV5q2rHSauUDu+VhLUtbJDpE
rkL9m1vQOMRIbO4SWFAx/pF+Gyj5iY7+cmxg+67+sjsTXSIAFLCAySamSPLaPwuhfCl+QAlLVrHq
xQMyXhH47eYca1Y2Q2t5tdggkj26MSeZAJuITuMX/Op3iOySJlR8ylJEcVVoDtEHxhb1CPicV1lR
/3uFmJLzHgpCa5gA6voeD8dc8B7HjFY3szde6TTSuC64rcw/zyslXGUe5n6+Nsy7hUMKdAY88SKA
bXSSP23FSEEfK9aN359yzA/Zy8651kagF2x+XltvbQixbMAe7tk1ffDJu0/NtIBktYaWbNjgssKA
TWjgAojIjwCXqmyP4GyoaRumxEU05rRK/CnW1CadoEsxlbP8D53vUcrZxBGjLVNOsYI+QvSHsPrN
qT5/+XvyDb+iw126NwkOCaW+4zyF4ECYhO6MdXT5gKd98ID4NEYJ07W5f7jVIua9S1sKCoIdUc7o
LoUOCG4/xObcW/iUHvNpAsTGByEhSGh710gjTvqgRHsTzDiuQeuqNCgxM+JGyMbAYQgkLkyc6AeM
MxNDFSfFArBkAiRmR/K7vVkSnfz//vjy2FqjMH3+SUwrm7iY4zrKeyU+Jst6eLXuQkGj3nlbQUq5
InTs4xv03mxLVUyR5MGriKbjWe+qEYmXqPQ8DCqjl942ljcFeNMnavI1AD8IPBpwimbVcIzcyyh/
nsn3yGGYZ9SY5b4pB4tD2XnafFyg+skwDNI4/CtgeJkjSor6MeJgcO2XeZ6UQ8QNuZ1VXfhMeInh
vkjyFczIBMLaJJFwlcNrOURTfUd5fJbHWPJ/w9mWI5MJjooSCrp4DmKsF8Xr+ChBH2BT9tSdFJdY
/fP78YQXfrd0d4c4uJ7+xJFqbPLrfnZUQbuypxEjQvvGiNEXyMS0APdUkHXauC6EHLzPZ18d77gz
yWu2rosQSNdhZBqVNnoP0kN7gkmBmfNmeEc+oJKyhSt08oUFt8EO4cwf4Ioqf/0TjBlK3fTmoL5S
tZbHvq4klyeuLz35qez6GCBIPdi4yvUb+fBX+XGlx05sh0a9SvFuPkUitnEWZIjhcVJYUmweO5MS
L6fS3glsvzmXRJDsj7rN7Sl/FPa7tY0DjyRrbjyxIc20o60A+a9qRuPLUa+Lu9UCMEJVDKQ0atBG
uoxbTJUW4wJBPEBgMZ5WH6Jzxf2DRqriHWIXkpF969CdkbeenvScynWfrL2vNWm3H4PlZSyCkjul
+oGgjvqkiNJmeijS6fr4U6shxim/FF2PxItB3LSZmqBIZVNw4xLsaBc6RtWU+c6aqAV89r8yscJk
4/cOyBxTt2HVj5LzTbITQKYPdiBekrCxW0ui9Z79sG1lh2FYGnDAkZvh6KvlrDpemu4Y/DiQhNZn
MEAs+MfeH9Tpqbp1e2LgxyUbvXlH+vvR8UXPEdmuk8BeeU2cZMTy7/EkktVbDXVXK+9Hanrago8R
DUECEaeZOIA7RbrMcV2jk5Yf2pL/eOGmdfSVN2mDUCT6FmdkMfnUHDPlLFJqAwAG0HgqsId60x5+
MiROcPOxflDLmOeHq+A0/NyhFqUaDI962uG6BX1iKc4jYp/2ZDQTuEnAQOkXdY9EtS+8U8eVeZWL
ZCHNGEUcwVqUdxQzgMalUGUX0uH8OccRCddAKXeidh+r8Cb6Na9CpZ+297yBjBXlvfe69GxOOmpT
1QQNy2ThuBFH8ZzZt5R3Wz8ph0ttp4+xdKSaLaOhhJHB1alxiLQsVsZRvn4ue0VVc9xfbI5zrkIX
wpwNf75Dy6Pf88JcYNerxYXtxphq71MCJ/HnKbk8pQHa4B07y+MKwjbHhyE8l9ffgXgw/jrybbct
na9IRO/zJ33KUQ5H2To+54IhI0RtnfYod4X8ymJy9WSz70sm7cHKVXsq6TR3p0B3236qeN5gE5D3
VHnWQR0445KCh9d1Qnkv2Hx38wDFznFmtftahK9RbEW45C7VYp6IsOUd1I5FG4Pkl0RI6SMFvM8R
Eg1Y+ElWAuvpg3VyTfGnZjlDhXNFTDgfGPxqHei6APgKBWwS/ZFlkdjBRmumtyyftVPF22wNuEdU
nocM9JVBP8Rl9BXkNhC0naKSSdHCEuhvXFvERyRE5+3a0vrpfKTQHMCgtTFWsNiAf5V1lWSVN89m
QRvoFQ5wesL8V4utkFTUUbC5/z4MjoAo5kuLlGj48x/JAefILNo863EWpBC1YhxuIXXWkSGSp+6O
JHzCpjMp5/9OaS3sZA/mmdfCTnNJu+2IaK8un0m9YDNGuNcdd3zCxLTPE+zxb7PvJB4ddWE36WjS
agENpEQ/vk7pbwn4JTsztIgF+cxZnVvUkIoM6TKpik0LaxG3aI5kK4mqJK8TxdBYIuPuyTmKyQvR
jh8xwuuaH+gTKckQwyePcSZePCIzjGWTx8riZX2g4Dv7Z/HQzb1o6cQZVtCEGvmYduR2eigD1bWX
IdLno8yvb49n/qCLG4fI3y6Cd8KketyzUCXDw0DRNAEh+FvIO6C1brZbUmRYjtCvvUL9Olu5dWO0
seQmJDLjGROvyj+ZlrwMNjEYNP9e7axcA9eyvjx7mm40oLP9IdVi2lGapPQdinrRQw2zfb4sMaoU
QAhy5mQX7K8sLn0OvAULOLkNAxzO8xBV4tiuiG++194nQcewXTG/PNcb46acnRDQZacUpe5ovzKH
Kn3v2yPag/U41sO4RhRuji0RUIyy/mC9m9MIYPqNrijmh+UzjpVM0ZW+F4S1AIsLpcEWm8lkl1/M
v6a/RiycvVQaaNa0VCWnGOwDkFd1FpTovBps0mocEDoYiWjEW7NSAxlQ7HWBpeiFvD4tDadH/+Xq
U/6ToH21DZvaE5oSCJXH1j82yArRseMbK2fq2/MfXkrPmn0+HwJ859LzZnEu1yssYiKjaBtro/4Q
3PxcFkvxjbW9H3Eo1Z49iwg+eXO4XZawsh+1uLgpFhPJllDr8BAtewpN9bmebfddVUTcZAOwqU5U
UM8UkUKvWM4eoVGzB+EHSTQbK99KZYIjTlfLvGsnbG1IOq9twGj+8NyYdfE9DubhpDjfeP2jcW57
eMQ8MczrtV1r87qp9ipkCCX19hTc8IwrB94xWgwGLduWxojW4ndrHwyqFbG9yMcTi/JasnYrPW/k
AB0MXnpPRCF7PCIDmC+xlkAbb7kMMF1nHrvAbWE4JpXBgvOGIMR8JoFV69APF8tPnNyxyCgQTe6x
MhW+/K2J7P9oMMurgRyu74FHpWLpIHP7oYHgLJ25DTCKZHJmsYup8NJKF082SpHtu0sVTgQpIViD
08UxjneX2P+iXwQA2VleD1H31YiSH4qix0FrgBODSnSv5bIJ4mVqSzeu5k0HqcC3rlQ0s+gyA3dw
NKJI1ozXbfZN5MpdNL/q+9gCYpWxdIDncdYsQRT4x/AYIbtM/y0RogTmbi2Yo8ov5ehmKiJ4TVGs
Wh6iq58g0slYyE2Vh0cQP604lS7PwsJ3LWaZDKYWeL04LpLVzYCnadtnUeTueDgm2A+WiQPrbSYK
agtjivbj9R5vc/5Frjaa9QnxnC/UMVnj2zrK3JFBG4c/K9ygHuhrmDjZuG2OdJ0dqWRKA1vmAirs
nrSQ+bU8RYHiyTDXkf/c6Y3xSfbj+3GRm+jvh737kkpbIbvwF2l/wcRLmX1o+pnHTM2EqD4y6oiv
sRVaXKBvw7aKqYBj3t/eVv/ZbgXuPWTMwVQVsDVCQ21nw6e2F8zuX1B1Aj0vv+0921bM+B1up/O1
TSa8fRqg//m4tlON/khsD+R9erDlAsILhFE8cSS3LIrExWS4EBj4kxNEusFlOqDdXv/E6JBX8kqa
gy16+ltYGos5iha+7Nmns759P4SA82a+3OIrIBJWJom8HEaJF8mFQJpiwwcpsihP2issYdmyBo2z
bc6ePwrPFr3Vqth+2rwyP29PC6fX7JYUGcVY39+Bk1wNlzN/rwLzRTV7dV4iZXf+RfHMRPEZu/iL
gBadaBGjLxKy/7qUrQ/+q5ZCOGHdxourn277tuLOh/uvwPOLtU7b3kHzBugd0hZ1YW/apPULJVXC
tEnLxgC9UbKbYemAeDyKqAs5yWcYXqjnHF7UL4OSS+Uu5LVX6szsxd9Jn1ha8em/0cB/C8PU62dv
ZLz0lb/7cRSxVUXK2uKa0mJeQ9+lnSwDqL0/MOEs5HY58UnlV2RLx0kNdAPx4ePxXaA1iRjMHGv1
3LUUdKH2Mxyko61icVmV1o88WabQMJdaF6KKjeR6y0yBlxQQ6uJInysunvHDRZRCu3sD7lgwhxYb
Z03nSB+8ABP73JdhoFQ+qx9V6DFKwtNuoVGQx17SXIojQaLL5elXpeWsDUs/Mo5ULVR8CR6JLSJd
lrreAvyfGS6rU6Ge4EUz8NRR5vfSrz9lzr6xsBQe13W8hsm7SYGUAta9c+UuwVNVnDmOhIlkyS7b
pPT/2+Yk+2BwILU1g6nvaAHTrRwilfwb2D/E5SPandvZ+wfmK7Sw3r5NmgiEYUowLZa0rGL8G4wz
rD5SHEJu2p3fk0GekwSfQgSXeUs4MHP8WeJI7nnI7X1WFA71ni1lvnjHTfE+KaKMXLFmHW/Mh9ul
P9pVlAY9Btb/OPf8xFUQHCD5g/W5Ey8vbA63weLLmJjBxlDjakxhSDxV24lvJj583Cf+PZvJEbMU
tGw+DNJoFYJ3AjbHL16izDXGePdgp+bFdbSC6nQj3cI6skR8fNU4MWnJJnYEtWlyEjBxajtHB+zG
SeHp2fxzG4DvmeWDN8xjT8ZwjcaIrIW0zIUhH1mxDsbwpxcnIF5Z3SYsMenFFXcmeB9oNyocXJii
91TpVtJ6vBaPgViiNnETMjAQsbvwFjKKKMEia/CXTU6etKcK13iNcXExjQLcNiGEKkTawRW+wcua
yRYswcS52D8LgpBFjZ27y2TQtzwFHngozsqfn7tW46yxy8PWOxAigGuEGXN5Pkty4jMMqdDAWbLR
RfEkuN7CTjl+yg0qvZdrv4t8tTrZqZ1X12H4A+Gyj6l23AOrLigObVRhNfcF/rdkf3gSXhIIWlvj
8Bou8/Ark+taZjdXW0FIX1yLJgYn2t1K/SHNL6ksAqfwP8kmxig+ycx4txyYSSa509Yz9gZ4rJLY
7a5Jri7s/o9A5LWfOU+sLryvhHq6VZvLeuXEJlWjceTouZcfmYqvjxkWLvazr2s980pOjE3j67BI
nj4a1YJuHruZKV/zNZqYAkuUBxErcb6cuC4j3RSeDsOmJ9xMy8AV3wNkO/GvuXMNMMkdOht4IRtW
5G6CFaUP72Z90B5WfFBMndyZN8E2B6bqM3wy5Rvq944y4W9pR2liZLCV0HU4v9xLEFdmSky2n+U7
6ILZg8APWd4SfvXJKto2JBUKbcfQvneLVNA1P5++aKu3pRQLwxCSQvCz61dUoABKzFY6hm024Fwj
dTtSf7YvaOdVH46fFpWjC5FDhhs26FYDK7Nomt19YngUNV2ZEEqeTlpWcyXJcO1QvrVH5FzrAmfa
noMu7gR/W70j3d0mjPT7B+JaDtnGu4ebLaWaxlHn0Qcn3FUvG76yaNXMuiUJrbl6WED2LGV8FMkm
5OB5/8Rnr6iyJFsH4FTxjwy0fK3bC0M7mP5Nmjn8AeAHFtCsAwEkcEAyX/FwKWpucexgz5l4Jc8r
amiyoQi3Ay82IxLR6fpiMrZ/jS95YgK1tOCzqnmQnxTTIlxvi6O0lpFaTNGXXq6VzEMZjalOTT5j
+BKqmYhHxIQRElEnlsljuO9rJtnSR9vOVqfQI+tHEZYWcT53iHhn4RTkszBi+p2aUl/OgQ2bv3xP
EETj9ZqfnE1KPIG5UH8FnCxUhvq+50NDIDb3tkYIzOd0TjD9hZZfTU9IHlCWN2SOrb67mVAnNipZ
G3njL1HYmoaCshPbIgYc/cyqto2w4XhHwKGB+Fn9DI8ZHyXmPzPY7qJq7FcYt9qLHJHJM3cCYIYx
bUe+5mT9l/NUvg0k2/6tTUx3VP2Mag7xZehmiHhLIUqPYmZZT49zq94Q7ab2XY9Pjgl7/SaYk6+D
D+uzzNpb2S7hSKkakicqym2l/XjPvfgJ4NZXcWbXC+OpDhVc1Am3vyjl8LYUYj5S+um4/tectJ0/
VOwcJ4bg6DjEaZOtd6gKRW8kL+ect1WYfk2Fv2CHYFQQDs31SgLnG+/ZVX0BGVaOLIC4SoQLCkpq
n8Mjv01Pz5AF0Cu4XaiiVgbw74exVl7Eid4zHhevb1c0eyHG0x7bkp4AvWRupYajzB1ARDczbnN2
5WgOraYJ2Bf7zLbO4FJEDeWHzwSXzNVLAcooA95REVVhYG0joDChGMBePn6+5PGWHO2TXz//Ccgu
u63EP6CXxUnmSPtHz3tPJn9JOyfNfU6n0vlAguvkZg4arpdmSp4jlSwsmL0HeiJ3Aqu34EOAipei
OqYRwuKa+CXkjemrIqMYxp6WbxSYYQdk/mW5x53zMOo4aYgwldKhPIFpwcZ7s11m3nxYHgBf4m/b
St+QDmeRfRVdHEhv2t2ixD02V3Tw96ylTl3kc9pZgqcIcNaV9o60spuUUU4Oj9Co79qy5f/6Rkjb
fqzGBY8Et/+v+3iFmmMhG/De8ANV6VFy8spo6dFzK8zHNip/3tkwTKDgi33WvwmiXCnVzF+x8o/2
XO4FJl8NtVQSw9hv6cfkJL5RgMYkOp2+CKCKyNVmc1yHC9AXe1V0t5Anh7KQ34GR3YKgTFCSpNbX
tAP31Bs9jPuAKiQUbIbh8Dfdg6riDWG+4EiSyKwwVFIygShlAMPle8rmFcTzopVnC3qzYcPP7q5v
qshv9tFj615Y5bxhCrhsMYG5sBAxa1NEV5tT5SM1K9bv8BetexafhynP3m2qbda8CKhubHlG4Ai2
1IGJkeZx9zs+i+KxJknAUSLmvx4GRUQ/mst4uTFqxPDr5XrajNCTfyG1Tc6ChEpJJad9mv+emUkx
TKf37g7YI56X6GnhcacP8nKlal7S1DYBK83tD2l8KpqVXoYJXfAy5JrqVUhsLK7G+GofdB4M2Si1
W5oLlhMixgxnQlT78I8QPivw28BPGgyO4tm4robH5dfmcA4YmMsw+SqbUaMgW7PoYnOS6rgRGmfW
c5QFZXKNWJH8NtNZGKSZn2M7/gKp4aRlx/Cc5yKD9Hkyfg84MgpVZZeFzf4HQ2NuRwEQRq5WAAo1
QgT/8/zbb227t4ONwtgFbh+wOvspoCrGyECMekjBITqSnaqFP+lWjyK+gZkePv0cjIPVw+bPXjAH
qoq8GUDpOlLQjCw5nfEqRlbR7ov+fKFvwyofsLfCDR+nf4E6zhNX7XCT0ok/DYQPZkpJXJt7zHas
wejRlQcMCTAO3bm/r6QlJsh4aPQ/SA02DyFByIP15buacxkIMhPl/3ZHwAndxqXO+jnk9PW7mv4c
NUTmtYoOaHkvmhLE6qe66txf0+zjd7BVboCTIeOLZ6d2GXMbxDFd/O5yf+vu3TqAsR/8c0f5gnF6
y/BYzZ86SG/8qToo/4T7qVOcir0L5rkaHgq3lQ1TlkVe2hR6u+E6vry9FOaTGAp/qK5vOj6YHOtE
E0Ie2cMxJbMO7TzvKt3GBAX5I39PuKzplSCfIw5BhaGU3TtYbRrhNd5gmFow0kAVmIvq+O9JPvQK
17RWEbvjzz/ZZa+snysysD35y2RjD4GPtl6E2yLH8NW9N2JWdovOwwNwZ4vfstvHoVKRZ3EwsXwE
LpzTHhwCUyoXo4mhRpfxTMM/VrFqwit3fvA3Fz0IEf4HpzLuPrlV44cHsxlS49FM1VEvhK0Q46qS
/+IHOqNF9M27MiZQMqWxRwUPfJ7eg4TBQhMrjqBL/c+ejhTrEO+DYkOJ5eBBQ/pZYJVeBaU+U1AG
KQ50Yzz0tJliJVBJNuYDC6LGOHQEueme3xYIABZEl/ef4phTis4oQ6+ac9yz2hJBM4QurxmUdrLE
sG0thnKyD1Pobug+sVYmiTtdXopdJU1R9JI2RE+xtfzheQ5FWQ+CcS6TCFCT9ZWKWeMIyrIOBnzq
IcQyf5u1L9Wkz+wJ+Tk46IcEEIYP/2RSDQTuJrpw/eDfnrBsClgsLtPNTNs/OABNKpn+iAmL3yNV
as1z4mvL1vSFSE55OyyXgGeTPopsSpWDd4JR4zq7kyx5aFpkGZh0ItFw0IsaNc/9PoNfmtepD2TV
VDNu/gEO5C2kWk4YoL7Z15g7lo6MlyC6BCiOeh01MmKB2JuPo9cfJMteUUWPfxzORE8VQYabP2Fr
AfU7RmQ4QuoNkSQ+I2cFUFmL4ztstF6pj2xOzlHT+G1GJ4vwxYBtrOoZzHYWfG7KDJfdoZuQzMor
6uFcVJ9fm5LIuTWtPa4xD6/1JRa0eJDYt5gcwT9X5L1IJ0VQwbGu94rJsdHeBIB3JKSXMEXe9Uvh
kqUxqyie0Q4fyMzb38iSSHpo35sDYrB0e3At9Xu+EqCPNkAvY+uF8GTVd+HeVgfv19IczsmzHcw+
Ndtswv8wHIGR2Dzmz8oUrari33pNn8MN6QgcldVa62ru5wsAQ34OCJVzhcvOtJtgRitZ+9VH8Gdg
yxKzKwvPl2ynKSjrda2AHEt+/x2hqsRORzvqj/7a+nj5Pq+QPBAhry3DpL7CqlvQz+pdLZtYel63
KCn0WA2PoLJ2kAt96fB/Jd/7W0wIn92ewGA5Tc1IvbwmFAYjuoLj7QHtZ49kzde9MQIgMbncZjY1
Z8+L551H09Bqjbqbo2Z7jgVWvJsCHObOYdAFBlmOGA7XLDNqyOvk2v+VK7OYg909UyytGaR4ivHX
D3CBv9SZ+Hh93uhPuWsCPgxBSaMQXcrlNUTdyS3rrYVp28iisDzGVXisu83G3LTfoQao4pF3sP7r
2d05vYg+20Y5czTaCmr0EOrgeiFiPDccaMY2TKwed0PjbUCVqrIL/qtXpxluRCkGj7OcJuM9R2EP
YSV9JI0idNXKQ6bTg0ETi0KcjxdsrYvOLvkMyhacPPTV1In/8uEZYbRbAGMsm6lQ8U0pfViit7/y
35LesgEaPQk/F332HBpwPG1iNp7Ac1vqXHn4YC7VWtfSyCkfa8iOgFU+ySHyGC5sE1cUIcgwX1fd
xhSJ7MRoiBN1mJYIBZ3br4040iS/Q7FChMZWD/wCGrQLnNtgoqNlXHq5Oes2iDUkCtRo1YfzulI2
VY2LDPNeOpg3EPc6NR8/WkyFI09Lim4X2+JKMgcqplc6LT0Mm47uvoZbuNKDrjLXURddZt9+pgv8
t02MYBOo9IwN5eCPlEMRO3ADRqGd/UuFO5PghsbBBrrRX5L3E1Z6bAuOVWhEm4giIm1Uk0MhQT1V
GmDpA4UNjsfvk/8hA0doBO0MRRq2g2ILfg3wOBFI/uAzgffzb5SZsnIgqzFLjWnNTgu6uHgsDkqT
237CcLXlkYeFiU3s8Qsm7SukBfl2k8Vi19+EnvkcTrvpUPYXNf4rIfZrdzQ8fMxT3D8s6h2fWnVC
ZSqXU6nFpeRAr5tubOoIoN0VzgLEGVL+sX9F5zlyKbljCCJVC8Vzaii2TH+s6vCp3UHuwcuAttRd
Loty9AvaFLmYCdYKhSORV+l9G3sURU6udn9FqWqxUT6Yruw+uFxfUQmUii7An98XiJx/xtryRXvS
DYXc6hkwbBdku+FvkehwjZr1CcTIN6yWwb9Rb/ftqAMkmxPZDuSjP47hd7i1oESguujXRRwzfHft
jpmqOovwxlSwRR+AX8SPNZSmpcXvKQCUL8Fk7mbyPPRAsO+pTEUaffnQrW7QAyQP7Zo+SoBGGNJX
+eMh/H+A6bKduXyZ/CXMxx4O0gVMOZDUTO1qSQs5OUPO/odmfyU9Z5eELwcwnT7fsL+UWMy1Jsqf
QDXdHrAnU6hXcqmfTLKn8hnAmzlCbjkQuAjOXpYj5I5i0zfBSzONuHmWu+nKv/YMytmvx9ngNMRx
54dJb4aMFqtaMo/ZuYwLWc+xyQimtGaWvjiSL8ezY5wKiDsTiSamMR6p1Wymlfw/JRuh/YVuvCev
FXIJwbtqLgN6xbsZY4HZbFBGwxNVrQeO3DpJ/pKbslCHAaY+UvzWhPQfGCSnlrDP2wvBrvxv0Zq5
vZGyzBukqmztjEL8ipT4+UBM+y4LG/MnQ+MrwcnxouIxEyPDNsUebQbxwPuCLVD9LjW3ahK41kL/
YXbrn79y8P7PhGARPXsAzPwdCXZNNpyHlCDe6KgkSXdcu2zUwCu/3efSuGeYyha2QVTsIp5ysuvH
S4amtNBDlLScQKJuvxr8D5/oTMq+5dLbHqnrg+BvDG0LprgBBTi6ucYCfeZ/c8GQ4v3q5t/gVp8G
WBdaTmMmtB1Hvxtfzv7pK2R1yfK0uaBlShEDCU/4bbC8/DqgYlmCLVqvEt9VbXg2qhHwlwilkOoW
nFBXe8uRXFWl9/VWNeYkuB3AFVKcEf5Txob/U97uYXQ9q0Gk8UKNvuEqlZ8MTx370DJhdqeaxOfR
OK2eqzpmGTUDzcDIuEpB4riygnsqrPwVrR3b3ZSMRLz4Y4927zpdQbX331zdpzWW2kg++ZerND1E
sZGAbCwYr0Nbg0ZTuHFnv5W6M5vhAGIFWKHAeKzthbL3ea/YUljVqha7xT9PY7sry9dnPOH8ZhQM
Zf67US4C53os/+zyKIYdWqljTdkTMe8W1LN5pSPGDkGGAfTRiqREehf0DCGSM/s9RBRuUo69ZrP6
yHLvij29X1sIrd2NHlMVhBb3u2pZfpxT0QkKibCkQFJjY6Wx/RLFCIOqQUyYlROeXDojAUnXCZXN
QtFTwZkbZoDvSd+BaTrMfM7d5YhCAwEgiImyJz/a5w1VeQQs7u+XjD1XRufe1gzUkRH0x1hRzSjM
bFtFDGUYMMs+mS1jtvBvl9arCSJ1TI5eouqv6dkbaEpNbfjI8o9nRYjQGq/O4s5w/vo/aHegc0+9
VIwj0RI9vtmoiYSQ+U/b0EDeDDCogMocncnf3LS/PrNQFVBCE7T+NTe7wcHsRf3eTQxMDqlp8pTX
uNMbLhIBe3BHsH1jFYIQ7XI3bClM2MfNFmGDsgw5Ago5R9TLIcF9+aBYXHfn4hVIsHxhCWiaH+8j
deM4qH35GYolL5Nkt64UnIi2+xiq872u2mcn1tWdktsj7AAeRqwnZ/qCRTOf1vOmuYeLlp2vrxBT
ruTHWdT9WkMMWoMumrHzDC9awlm01z6OQOGAvvsetTwLhU6zZhGAtgLxKUIjW8H5Z8WOXIPV6lcr
SWsiC+chRIisJlnu1m95C5DQ6+hdVc+KDlf5KssyBExlJ9lBS+3D6va/II8xdl7utghyGyu7V1Ji
FoLXEnfRRf6+SbdFS6ATOw1lKrGo00ZYbgsuOk4hAXqkyCgAWtKfkG0A8jK3/CQs1Ot6Xz2ULtx1
+jaP66+bvfpm9FSNzVEMF9EbkLO8w/kStk9f5cX4vj/PxN+cC6tC0/655W7rDi+REGJfFZZoGEDP
hxgXKsFwdTaLNQd7bNxPQxqVAqdbKtZAbY34c29rdZA6eq8vCATFk2n9gayFRnRQ0XCumQ1rxUkO
71KxMS2xfAszcd+qaZ6lGkW0UDqdX0ODp5Cflz61K7HhkDRzNE6MZQb1SeJE7eb0xMGn5Tm1K1S+
h0+BdvdflFKSI7qGrJId05+EVFFAbT1uGNkcyt0fDh/SbBVuGsPn2xrwVI3pKNnghZVSN0fCIhlg
DXNwAwnh9eAl0G+HDwIWP37OmShP2CbYJifqK0nVTH+68uyZ8ycb6T7j/kiGJTQ/KWqxs7+9sOVX
4TWzF9Ol+0BWFdZNIG3LavgDfSd7jsJHh0MqMZuReOaddKPvDoF3wCNHvYK8jMjjEZ+KrDvz16Mg
2nif36+19MxrL2Hle4ytIuCg3FnKw3VRZZ5ea2PBrbEip+V8EIJNoUOj6t9TyRLy3seE0xOlVZXx
4mmm3J8FEMuTJ2ImCmX1sGAQNuhYDp6+9r/vy3AZ011DOaUhWzd6zYmRrOCnd4R+Zxc6Sj2v827d
9X9bk+PiPscplcLFjlNGcYz4Dp1kmtS1+tUl1ExQpUaQY/EeOFdbBgExVXNqpzuG08VL/aFVLTze
tBRDI8AeHK66vMtWfE0xjATlTFkfxvz2oWDXmc1fBn7VXR496n67zf7I2Vs4wVHFhLzZm57XNYM7
esM0a5R+iHMQls++NOnKdju/NZBhiGS/8iOQhYLiWJbVQdYrWq4xBiBW02xv0xATd1XqMYQx319o
gV4krjdMu3/oTZpdHT1X8wHG9IIrdNaJFipgVMWWs85ZBHaAP5ZQ8kfp+NhtcKGWrtq4sOgKSgzY
PrhKRM7SdwkEHipA8fhNfUey5zdyiF0Ef4KpkEcfYKluZBPnpY/YG6PdVdLA03LoZF7i9OxGhyGk
EyUtyJQPAxe/271ssnDjMzf6cK4ZxG9aAf+KdOWxQeluTQxcZ2190BdDtjnBmMj8pWmJqFu0gBXD
3vWXeARtVWbHi14o/O1c2kGbYAGLN7QVaQ24VZrHZuDhbnwxbGnhre2aNUp/EcCrp0ZeuZYawafw
Kr3d2gIC3XBv96eylCjAQP2TeJVyJWu2HpJTHqVX//ak8HXbnZWHH96wA+AMm4fEz/unu+lD5qu8
tyqtYDWYFkgAIWywDZGpf/bWAr/rHslS8fQPJxKGd2W6yRVPcu7xEu60VeBQZOCFHi50ADvpttfp
l5zZ9Vgavn32C+HwWKnwBgNOaYQhQ6585T7ZXkHfYoxEnJboZUweLoCnJPmKVWdXnKyJuVjw08c6
Yi1BN+ptI5G1/1ACM9rUIuO62Ntx1F9CKm3OzNtGLv8Sr4fvNLKycvf5z5wFnTdpt0xTJe/B7EGG
5I82th+2XH+z6brfEUa42/cC5Wt9EHaNxmYjghljTSu516j0i5za3WVqN4UVKaGGnADOnbfiqpBQ
wviaX1iAodhPRxtsaW8KIrTJcNWh0enkvuQC6YA9X0zDDwxKdheb7Pr+1QXo4X4GnD/gvTObBnq1
QzoGKaHPqm4WdrPLkKSlDZo5sijAgWT7xLUzDFE6VclAqMC4I/v8fchn8WeTYRW7CuqSoejcUK16
pjwNRSfQuudvieimVz1fMmHRdmdDyH8s6D1IebauUwom0t2SuicAA6laX3wmNIHtO/Dij1CVF7M9
GvpyrIlnAojLsbHsvEL7V+Kka92dN8T5N5fhCuGGLH8u4D8EOafZTgejyMyh7Ke3bQXTfvlNCGC2
0X+FO1dddXNPQ2JDKGE6WC/nXN4ZvlvMHrv+iRQddXqCmuK1FfdnUUg54xlu7XP/uqM/Bhb3tAKS
UhKOYeW8gILr+2nFHOdeg7AX0MA7i8xDEmYt/yQ4gSp5qhKYHzBzIpj9hGrI37PwUbnl+m/XsBQj
o5vIQuuseNUsQQUmR/Vl4r8oc4KQU67U8+HfR63hXhBbWywtTGn9TA2iCIS88eT0Abpq2IL+PNGx
66PByEDWoFKeKB9XAc4JVX7XhqA0rJk8IenFHKDCmdM4TMzSE0nQNiO0h2FqLvt9RL5UAqPDzDII
xS+bfcvzEYVHkEtbYEPTWotq9whQ0jDc6vtGe/G7Id7a04LnhRfYHjQ8LGbBh80lIL9g1lieHPJw
TFEGUT1Bdy163klUHA6EYlR7hYNFPFghwLEPAqqBDs58rE0pDF7C+srEneVWTk8r/4XWAD/wpEUd
un8STyMkfaChLwAT8BuoG+p4GX02uUv3R71ORdYEw86uQGc3WPMDjTzZBfQgCl3FCljlHgcjxNH9
qHsopmQ7fFLIPsMIYF42QPrRxkTaLQZgmNvQ0Mk7YrtKRUahu/5eobnfBLp/fVxo+IOC28DTs4Pd
kubIWT6jFvJX5uJ7y2ER6pHWDxAaXSxqT5DhBNKDNxn75sox+piU3vA/5zCULlXbIIC785Aew9Pw
Ac9GjdGFVGQKHYRrRxNvFoC37ixvCJbFFmzkXdFjBwbBZceFdBzgmmYhG8gdxDGL+yk2SYUJZIsA
b4qvjE1c7LAV3KcYjT9XcH1/qbZECGY9ldGpKketS+gRx2p+LHRlgttrb6ywdCICCRibRgRlmT5a
8416zBQ6DoZ8EKMFRSmeGvg1zP1JAiMPA9HY16wapEyUPz56OFlA8eDJg6N+34b+uljgvpJab9XE
dmZj5TRngI6/qJxtI91xI7njeOqIecs3nEjL2xT2mjLNZ3dfkIpOj5pzaGZy9LjkA2lV0uzyx0qc
5zOhUAJsTCSr7lPo4+z16VQKr3ewdDb2dgqTVKMKXMJkNr/9C/Ocic+3eSzA6FIHxvVtrLueHlXy
FXmZk7nrRu6EqJjHu21mHnopq5JPwuvFF4se/THg9A7JCdP/uhcfR3LxpARlCC+KwEWpgVdmBiqq
wSVeeR0fzGTGf1qM3dckl5JmQhkt/9cNN4vVRRUYOzP9Q4mrzNwNjejKZD2FWZ96oeVLchwMswtB
0rixOUDr5oq8O87SUtvtdyEeWRGZUTHWvhdiCpuqr0pozL5PjxMi0CYzbsyJii8GnerM0Nd8SpSu
J+3GRyPwmAwWWKLtLeAkrrVpQRPjnaSrTLPt02qbHaEJ9SIKySUH/CgwKvGsskNlXuj7Wy400KtN
D4xR493TNT0nWOgmWsXu/Fvz+yuYLdtosxjV20li86UAPZrKGCJIwh4yg4F83mpsPEcDsfpvLezn
pcgzMoQxx+cY/UWOEHtTFz4eSKutxGhctg8euPi7pyTIEnEFmk9zk5gW2DxLMbEwAyNIfGXL3Om6
yiB0KsV22SnXN8O2BJ84rjeMelz9iQnPp4DAkNwvfnE2McfKHaofvKZ8l3gAEJjMb+WC2NQXCZja
WZZ5AoKR0rS1TqCrh2LiQA3JtLjzCUY8ehUX+6HwOgY99pm8yEPO+P0TYPylT20hBUGBY6KjSiR/
Gtp0Q28ZjruEeB0XlCRpk5ZFdb6pjaf7Oysvb3WXGRS7S74rGUAk9iyhyC+tQGupRqGtBEKRXYXM
r907WGNkx9hp2TCL0ibwmiuvLwAfg61zp3O7oAOh3Yo/lOlJ8DxeGGKNPSr/p1DvpNt16aMg9uDQ
gmYqjlXicc7QiHSSFjSgH6rN4A2MaY3IClUL/2EzlJsdSL/ptCQ60gY9d3Nh1l7xm1jHpPXUIKb5
Wd2Kr0J5KTomW/Ct3MHp/PzeG/18IOY5lslmV72rz8K3UMcTq4AT6vVbcwEmZglC9jn9S5dS/BdM
HXHWbmqYm9KFOQWaC8+SFMPLCi9r7Iglg2Ce4wiNSfrTNum80lSD8O+MprBLs21QM0lf4hl0J2ze
sbY8gLm/yZUuKYlPKaQjz06D48oZmZWxLGy32OD5CDs3MrBdubmrlBuhYa8tauJkRW4fxk3+jzXv
D7N8sn/OW4WLxhx9zDwt7rL/muJGVNJdv9JMBDX6+jCvYXDYk3/z9M/2PBLmdvVK0oNP+Lh7qfHT
TqDAXCxQJGttBojpgZgdJYTXgJqTvkd6YKall2rWSxq/Ufu4ejL90gpmmCo/4r+eFctxkhljxR7D
Gm4vo+k3Jk4PXgDxEzMXXn8yoKkqj4SXC4VcJINsD8aECbKBljHEEybrVy1Uucdwr8gMLXxnEOZw
EV7b+HQ+nJ1ridckTBKvu4qdaALWouQj5Ajx7OUTel6BSth/CThE/oaEY4o1iZBdQleBtqYHrvcR
CTCLvCSBmCbkPwFOg8g10oBn3ZTMqg5rzVnBJA2/jfxdmhZjtmZS1Us6GJtlVj4bAVqjFBTPj5Ik
Ry1M+e5eq7x7Z0qTPM6UY5BheO2rWcVkwoHJdXp452CYqagWYZsIC0kL2Dpn/jUm548/GCyF+q29
NaqdYvvQ8rJEzPeBskKV2BWTQbm4kPrrzFajQtBEmZ12EYufqUPUj9EwipMrvamcwtUsozImhug9
j2cn+w9zsjDBF0sNZPd4zTkCOW1UHp4/EB/+EzUrohwX12uVd+oxhC9kuJ7xjjvYI0uQZqd6VBXT
rduiAm/JeGyy9MbNKTI1PldJdQnXBmPirRhQbyyXgyQocmt/G2wVtPYQ/gT1HFeYpOlDjAr6Ykp6
56dvulMU2U8LXXKRZGFKNtkslT33fFg9e7AkkbSdoZFlzR2qHt+yCxs8zaHRG4oxHwtTDAbBGcgG
iR9MxPp5XQInSp9lSkxVsGSDkavF4rlFl89Opd9i+neyQ35U8KXuux+Qx/J4FprBFmBYAoj2FT61
tm+guiT9BYWyozRMxkLubbkkkFN3421cK55wDpVlB5a43O9clrYPmtfVX9yGSVQ5vDCFVbeKgvM5
cQNPxxgb3hSeIbE/ofUIR9ujFrU+r/z5QoZcJewZngyVdHeU3ZEerHKQ7hGezA79vJSzWKNOlI7k
20pQVxs5lj0IceC9t+nq/tWwIAKlkMmWZJRr+X5BFBbw+W1IvjL1ZM/53qM2v/92MtAgpfUMPymE
TmNmWeYBa2xHPixP4E1hXM4cuLB56cI9Ky1Cip4XybgCk5Z/3SJWre+SwvDPfbgqgtmMRGsENQOc
Wbcg9AgZgFAsCZIEwjHnLPa1QDve+qsnI+wh+SE03tngXYgsZX87ITbiH28EqhHOlgmfy0gMzbX3
X3Qe0eIuTw5416Ex8laBUlWkorxBkl9y3rq2jetMfYMJmDcL7y5eW7SgEbd8oAHL3Fhtltfw8YEx
54Zp5R8ZieBSyYF/wBVvM2q1BBj5JCUklxZGa0JzVZWFTqRIpPfYreCAbFgO1uCT8RwRUkMZuJ8L
ZDvqaefz3Ug632cG61ps5/y0EmsQc4CflBh+iEFqNVAzeotjUw/GCQAnky7FOrh54ashf6OY9RUh
b3enf9kUXN7ohgmjlyGakQwRFVSe9TfAZF3jSxWcrHYTY3bAyta2xQe6yQFLaMVP99uObax48dyY
bsd+Hb0sEFCOw+r1oGXFkldaqWfQSXcmQjJMtSc+7jGfK79v81RgfhXqa3SgZdaMZ1luopIJZn+7
/szaP4qaL5GJJJODD2fwNp26DXpkWMkW3yvxl4ioJbAkp0lPO9JNZSj9ixXNiMXSsuEbOEJHUa9S
E7eep10ZDcX5l0x5QrOUU7LlxmwRErnay/mGf8Ns2jt7TgHk7Mx5/XvGCAnnetWm9Ve3hO087ELQ
YvliCyYoaszkVf0wrBA2L2otxVWjY7SDOZ7tvbepPZUjk+NiLWtZmSNE8m+Lo3ddMiQDlENFG+hB
xTKkTDraLJPqxfcUlspjebfkvsG/ZCijXresIJK+9PuDCKxoQOJXsQAuQOwF+YTZRYyHcyX3xKDx
P5lCTuavbeUR36jKIcNyMUFaQvij2orKVx17Zhm1bzFDTn3rq0yDUAAKe0tP21Ke//z4+mckV9ct
LE31FHDm/d/ZyEEcZu7uwAA8L8iE32+1ujlyT8suEv8Dx/4qgySnT6x8b0dQ2tNWqp9MsRAkT2oL
94Jtg2E3t4Kb/69yTjjSCJ96pxYkTx73zTL53iJRb8DMZu0cxgQ6ltwYGH96azhXPhUIqxOEs3Sk
x13hFwmbaWkc+cDgSpGJ9z7H82syDHbgROu6aWzjssIc6jXywC57RGOS25LFIcBpCb/wQ2naXPh2
p8wxdcwTnmqAnpwqz4K48/nFegL0gVtvonnEl+RAjc3jfrfR383nhqAx8dMXiFmNk2BfqSsqHRc7
gho/HJEsvVl8WTEswZjUFisrKoZ5A0MtcrMl678bldjRHUp9kWbOQDplzp/78a7M6shEXDTG1R7C
Z7eTeklqVK7HvQWK+3iuAEfc8surTB+AKylh5C1WdWbvZj2MXjGz3wPQpF+SvwsLrlPMmBtyKxiK
Rv8a24rO0vt5M1cSggAWf5C4cOBmfLnh7gY2o/CTDiJTJRkfGdOACB7n4BShljaYQe1/L4+ppbFF
QT8bz30VpTUeLV/r2yJP0iLIup5fmdH1Oxkra6MD/GQuvmaWu+vQALatJK3oQy2z+m0K9ekKl9Jj
YyapdIdLKTy1n6Ym+un9naJMo+YtEwlmMCaNC3mFi5N1tN6ZKWz1dWMiq6BqiYEYgzJmk0+UF+Lb
nU4pLeHSEQ18Mvk42OrcPWuiR4QUKcxBbCM7eOQIYDzmP4A8Jhso/i2yeUr75mVGPLaLSIucAv0p
T6rw9X839uk1FUBEbmY2q94QF3CVjibyU1svDJb/GdznZTi1ZeFyeqHUOwF5Gjv34V7+1di8c6Y9
H5b62NBL4ouW9wcsZ2dRoyJgmyhR+Kev97X0nlr+60NaDBNtpiWiZ/pOpPVmX0H3wJJ2itddyFZ2
flRqNvNxpv/uXS6YFEHIQocar7jjU0QbWzK36eVwdmsYp7GEHQKa0CZdv46LTgxKw1V9UZF0CcWT
C1121zc4Vd+sJk4TDnGCL2PBNMgZFL1TYx++kkpAbzNghD4COn0sYOOU4FEho7gxk1EEfyf7ESJR
xGOSoMN/bDUFflxoumV/TdJemMeUmkHts4AaRmSSSWHVwyaWcearRNrcom45vE9tUjkxfdrchmVX
cao/ph4/UrRS4IgcIKAZqqdzQE2OOaRtm7OeuQnsz0S40EUMYJ39w75eWmGMoOQ4pWeqIUIYMUXs
t8V3Jb6zM9XYPXb+uFJRjE1BDRtyJr4w+BJuT5wwUkE0Yj9FnC5b3QKk83eTgr8ic/nuRKvc7uPr
sTWh4wJTe6hFvo2VnsG9NFKeec9vRla5rtUBB36fzIzRaR079PRtQv7M740ZWb62d/9DbfkHRSGb
XwSQ0zOEZAO4zZ4HL1qwe11lRADa/RH3tSEJfiH589U/pBKaoAl4EFVdnI1AT7b+FILbznMWNP93
APHSeZUUTCCbvzLBjflglx25vg5KQ8rjb0EuBgd/oZCpDMnbc5U7rWis4NkpU8ZMWONVXHxW3KC/
rKhsrg4gKkCFVfTsJVH6bDZsTCEp3If5x342xiDZXIVr1MG/Izrergf1W0i4XJ46PEdZmVNeyknK
Gb6Wmi370XHM0Q4RIT4ydVBRC48CstAsM1rJ2oPqkBw9zvV/G3HMOyzuouxJFUXvOfXToUNNWJRE
VY0Mq+SdAfHHatVONZM/crEqI4725EuNJ4OzrWwDEPkY3KqXM7v594AzfkquSl0PSOmFIit39w48
QOCle7Ku4c6yutpCWsZZT7vne3ZVSweLZItLJtSwCB1dbEgKyERF9aCkW/QIyCe6eomD0aHiwUZU
SNpirxJlWEIGMu0P6NAsPFyjBBOFUcsxoZhpNeMoSiX7A/kcvq7gTSUbYQhnjXB5l3TAQvXxm7a5
Rew6+xhqH/bZq2xWrFH1t1i6iSvplIe740aMrBmQSKZH339/St3DGropQ+ZNW4EUbDQnPUcbFG5c
NIW6CZh3LLUa0yWla66KcwB3ihsXE4emERfh8O7SUZv4LtPYCOCaQ1o1ZDzv1CdMOj5+AGl12Nd2
dWc8MJbm6sdcUvMQW5Ymr9T8bxmtHv87TnGF9fJ2hT8gBNSCnLZvxcL+xcj4wgKb6s89s6yKX710
MVTp+RBFvjvkgCgaL7MspKBSdTqLK99Aydwi/lVLbrLWVVFpcwh+3GjjhWFprCf+8NtQtMcsiVY+
IadqMaesGWI8k0gZk+DeiVLgbQ08bVKTVdDi/OLBc1RNjj04r/9L6cPlRbekpkCkm0VbIjHpEFtd
KxFRtEanVfOls4LGby0UPIv1gybGGYdbLM9QFhgphlEg+kXaVhRBZthGPppLD/9vR8Xdpyc+ICcz
yby6du6NBOrViFNbe2l/e+8bGgIOgwVi8GiX+47EynvIHG6Yac25JFuSHtvoanwq2LD3pr4AZ+VJ
lC9Z/TOqs0+EEdT1LXIaTIveHTh0vbLH1zqrPwvw4rZNH8qYUOb/7LvsWHpBdesZ8e4M+LDWqW7+
fSpNHvbWMe2G5ktp6gK4Df9H6mmGJDCTwmACgPwkos6c/chcQyBV7Zx+hXEb/WPuHD3abOqmntKx
ILf8JyIEuR9y+uCAWGjY2K2JVLlJFHDOVgGpDQdiilB5MIUxFQcKQ1YCESzxqcRPsXU8QSq9JWBq
27eHODHWrBUnEZoTeiEVlK0KHNZbZgvb0e5axUmBr7fCb5l6yaA1faXuDYpHvH9pi6aHfZ6NcDVG
N3t/BKmC+k8svLZ3fb+BegXYtr9aCwGKYF3NVke6UXBHe44lbFfHd/vOGfVX6qMJfBwwJC90MXeg
i21a1w+gA438hmt9QluyuMU4KfP7DciUqU+zV4CinqtgHpHwkvy4myJjXl5XSgFWChyAGpAnjhWI
sCeTI/Ym290s8o86ahgQ8WTSJvOti7z8xU60cSvb9r4Ecmk6IUY+odWBGO2hwS8i+X3uer63vr+E
u++Nhea0PmuOctgrAjluc5eBJF25IQ7OknSJRX+isvwE+z1vJPChAzeDTxc8wC5j80eqqnyMxAQa
d93Wm0Ui4+sdkWNNPRUT21aJ7Js/+m6FmNKE88s0X9UmdY5KjakDHYjY6WPGxYMG5489Rj7PqIXL
488jt3B/7JhxuC6p7D3ToWCG+VgN6kH5zE7nCQWBcmAyoed2Q/0MIPEz2GZFgK/L2aqcd/bPkaKM
05pKZ2jpgFlRcnCWktkHZnTXbla+mQWAyDUMBvEGC42p+x+ydE6Y8Ifrz85C8ObX/VbOsiFLcW7z
8eHYVA3cG/WTFuBQEoPvOjxlaBw/Je5K4yJqI/xXAgSW5zdkN0C6WBc5vcGeEpuYqkcTSNzLbd1t
kcm/si9PTkB+AgyyTCmpofgGC8S218k2yZYPL0QJpfkFBhfUEH+vxZ5McOT+jDapo8cVdtrj2cIz
/nQh3o39SwBjGnle4imk9FhlsJmwhl8BV7l+1Cqbg/+4TfV/oO8LXCO7vREGqIkNvIMAyLi8emvz
ATRsFVjNlSqRUB4rHzYm0R53XVMuUEDRxTYeG0DmcSU8Q4MxHLJTEVrCa+Jt5o4d6P/QjMZ1U/CZ
k55kcC6TXii3t6t1Km/Dc7IeX3gwWKGDlYvnUEUh5ku0itBEPKTE2mUnSipqyQVkM8W3Rfhurqmc
M269kITNlxUgsY0TEXhXSgX6H/hxsVvOaAoXPccHhbis94Ho+BoFXJpJyFymPPgzvFGacJywrZMW
6NabWkmblgSxLHHtnjjJR4yPhjpT0EwzdSUmhzlktM/ZEgzM3uf/qebRzPLTxb/bM5rThiUU4y9f
67Grj6LLazSOLHEJSsL2TYVSb5ri0Y6eUteqkrJqfXsUZrikABTp6sC2PYfoNI/nzCl/uik5xKAP
nLiNnLkN9w2sq0f0ZyRzv6/cEpdtE6OyB+dqOOzfbT6MadCq4D6MArnSaeZ41UuB5SZu1TsIGqXM
9RdCClvsrNUI4KBUbp0tEVN7rgK8vewI9kvt62T8OdlKscfMbzfJIABHuYVD+ozmqj5gN7MrGE4E
3wc0NIlWoJ4pcfVvqIB1fFh1jOlrq4ktPPdyDFRAlBGJc8ErbSkPg5+RJ5YTiUVWD5FBnS0zb3Mm
Xxefj/TCDZ50K4uX1PQZRgPzL7M4Kp6hpu65eLKqBfdmC7/e8R0WRj/Wlx0ddXbz9JopefLq6uWB
WeRRYj7/6qx28BH3r/vCLiTDRpzjfLbqXZ1GFPtNPXu/+NWEM52e957coOlpP7ZPbDsf1aKF3nvG
Wr6uGqy08XCDzbvBFmlftTTfaNz4Ore2jahL5apKMgWqHc1wHsMzCMkHwGBu6iY1i7LpAztUUemc
lr1eBbQFhlJbUKj3jJkq2BpgFN4ElD8mie/yYUFmUCJDU7kE7/c5+b9Jf6QYhHfm8ni8v5VkZhzI
IL7uINGTzRjSLZEMIsTKhqu80vW4qHIMlk4CzucKMGTC7JbJhIwU7JgRiU/UAuQ+E0CoaIRQdf4D
H0Rg5gMMmeDtYlLpdGwIKdqOxYo9tkTVxwiVzvP8+0/bQmV6e2ItQ6v5nY7UbSgWC/0b6I5zmvPK
naphHABAj8C6v9wiWcec2WqLm8332AZLLOBepUVC9bUNu8w0k0540e1wf3Mc+WEciKkqrHHgHj0p
JdnQfXeDk1aDNJxtt9nA+fTlb9A1EOAYjDu01zc6MLWzCB4XFwXSZGaYlYllw5TOo389U8KBv9UA
YWNpVWWtgclNL3dSQGg9mi8rOPFQDeSi2FFOn6saG/hIII0bd48/h2MW8LigCVUFgfz126p5BNvA
V5vzy2Q1B3jdGWwa/N4KgNIcLOT9IvFlhiqV9eAM7lBAi8fAHt/w2L0SQmHQiOD0BhtgKqIW205V
08tQmnnS71ac5gdEh2gbys/5+myzJLMkyG7X3q+oEPEB/C9gltvP/ugYmWhRBWWnZZzf7SvsJ6PE
CFoZE84xx1LfDPbxCu20ueduIswQMbwZmnCRU0AWJAGrVxIHr9V0JATGRi6rYGpnvC/MBKJP/Wy1
lAg8cH69eLUzlrFF++ewTB5PoKE2daAR+To31fN4xzIYhWeXCQlilH/GAk1JZ0jXnGHQ9PKBDiae
XFUSKxswy7sMTvMiW20VkDDLd88sSR9RYQYMzwG5rgonajG2ohwLcctcv/HB2PchomchvLzdsn47
B1nc0KvzCBqu/AhrKnIjfUvM7W71kOlgKaRieNV8nIJIGnPPNMdtHczf3Cgfglc8GbqEHjUcY62/
FOSOejiv6GilX7i5JFj63n8AP0AxDPBxKpnE1BLAcdWHrV0uNdXzYgjSz1w4D3HMsnTxdJbxF+bi
zwDdeTmyyxmdeNz3RFE4JdtP4FhNtFs5of4xbsVv9tZGB67XkSC5pRZhdvr9rbd4xppEWoxUKGzH
KNFYHOoqFyJEPIpXIhdrwblZlI9YUZT/04MnGKdXsReJac7foaESYcyv7C99ZT3FWgpS9gILa/IW
MnBIm/XaqaAODboD2SkoCZeA1a0TmN7mw5GClkcEQsOld4t7wIUcJxqEBMaaR52a/EuCs7xBAqp+
3WMSihAESKeeVYa+1zlGXyM6jKzwPuD+KdHxOcHoEmaXz5On6nYWx+pXGLavUYylzY9tKaII4m20
8XO09E7OTgY3VANJc1a4KVJ2EmM849WMdZ+CwL6cvEwzOovI1lHWcBST1dib10GajW+x2D+yDGzY
SgL8NqHkQlQ86jm843XAHlN8z4r0eLDwMye5fdqYCQNqnFcyqdCXgo3RguB8nJCgjcPAXD2lRIgQ
OjNXrIlPut94XvW+q/+N3WNWI3k859e0uGsoICPARhaRTmPKiBkWcl2P6q+xuYCXY2uOtJ6Dbhgs
ZVLtxzdDSDu/Bm07d9rtP6nkIK3YHOqGg4APMNNWjWgGJIUANB5vMUvHlFsU3igAoa9kJ1tH/j8M
47lTGulpvpT2m/Q3unpewjsjHRg8ENopGNTlFm8k3Xko3uH/tL6JqHbZPjtqcyjtgThP7xF1emCk
/dmnthkkUtR10yJ5hkFcOoEjcZI6PHzH+T/9FaHkQ6DQPHvy7I/bOYbfwtyexqaOLk/9ay5tS81t
X5TphVyAhLX5YWP3mifMWTvtuByCzhuCbacPZ67OWgO0xoGpnFIuSnfsw/BRFqs3cONmN7WBqbwb
yLNCgKvpVbvYTD7zRsQFF9EibYY3LwsVsy3BJ91D0ebArFRrp4MAgyz3CF5y0VAuW1JnoJcFZiVP
VJLOI1RKcVJsH4mPY4rJg3ZTpMcxSkedFZPahzkH6NDEIHykAf4vAFEZM2JYE77xme1YGr7OXcaf
EoLd5+OOvIwb76Z4JetNAB/r5lKRsscC2Pt/xGd/mriOXoS2gUnZ0f4fkfO4nSI9bRKhQFCeMb0i
bgGvpSpFW/a8wgB75I+M/vC+4bptY9uZEIrnGYVDw54YNv9p3pPOFkHyxa64gae71JLqwdomVaX0
zXJ+5Q3/VuVZxdXQpSs6s8LrsRcFfr/Fa5KOJQ7TPoeUndiOHQzs5maaJzs64CY+c467FTDU26ZV
YwxaLMTAeoFrX862MeIIukUCCmLcLfOBNRb9p6729X//fcWd1/FBQWdxkw1OIQvGSy+6LOAkmdSB
PSD/LFEbF7cpS0wzO+cWYl+VmU1VMG/42QrxYReNzEUM9P4ChYK1euzZbo9etrTTFRA00b4BATVR
HBk746hOdh8Ulm2Mza91gUojvdtutwYPuVUtxK7oVRiIGZQWEVJbrbTckHMJ5eyc1Xb/lwVrA8tY
n3HBFyYQuUwCuRtAO/6M6Nd+cUebSw1JhBJTr9bSlTGBH14+5vh9e6MtCK7AU1gt/528fGs7/sTA
OuNJ6cJTO8DX4JXzqPE9nj5B2/JJap/hj3N59oL7M/huEMnDul5w9wy4eS0MFPTNIJznLFZLO85j
OsPUOj8kjNSMsbH2/TH7r3nt/Nb9Sqiju2qsRqVN5iSoXWFQfkaTvorC16nomSny+nLDy5L+SMXQ
+X3tA1pj34GiIBzuj152vxSMD/8ok+rH1a55pSwY/Gflg6Eh31ur1E16XrdohbteaCkKgIeN6GTn
afFprL8ycF8tbRrfhyzUQTOzQbdJg7tz0pqGHXUKIFl/XJ+Xy6vs7t2cHIsWYch2t2Yr2yU320Cr
CfLapxbsmjLJO8WCs1f0G1hR1TPNIl9QUqC2l57SNmUVeq+8a9VDqf6Hh5FtSRlKbPfdo0PLGNzq
HjfhLb4gMgB3DkY5idRhVL9HGK5sgc7igu/8KUdlkOgC3ETZ3NYCa7k+33HYlvzwEsHvUgZQVde8
QegReu6AS0ZArSKsxRuKFggN/ejFcFSEi4kQhqsxbfBqg4B9jTdolK/wiOZla9roBc+x8YActCcy
9GXJI3nwbT0q9w0PI/Nbiz/ItI4S14n3Gc0jU603Zu7mq0IVwXnjETk9GoxRsygbYzqM0lgUsjDx
YKcVomZ3YGI3gh3sDF+Q+dAEPy7UMw+bmsZqcZpo7hxvOTlLSsjqY+40J9Da3cn0YivBkC2P9v3b
ZrDkOkvx+NWp2sKEFM1IaAxcn+fveCVfuCLZllSkxjvNIME0VzYv3OoP/N0TJ0gJycix3FE/nwkZ
l7zcN/SVzN+WSah/TzWcA94v4AGZQ3gS1MS0MzHwMyR4AVWlxaFc+jinpSh8ZmPlW+2K0KsTFaog
lGFrAp/zm66nlZq0NQxL6SEzwE7LFaID7Frn8BunC6vkWOCtWNvqaBkAEaVdFGlNo9zqctBhFer+
RTYZCSfSLbGkFijUKbSs8uE4RjQ89z9l4AzUYAErlq7r004MqEGT9wSZ9N9rD6hCMjQyiwfd4ktY
/XWGPrG6Yj05K3my9sdokhEue1hGGpf+MuFjGNEGIs/ykBWPkMX+HW1YhW+dDUp4f63Rp+Ox0OyH
SMKasIGxU7kV3WHXqaeWUsfrnBSkg7HxNkpZeM8vxmQIPp15L7CmqUYdmvI2OsnQJmw3d7PkHw54
aY/7Cp0C+saX0MnN+aiZ5v6vHBkzjbLGzNxGlv9wRoXnpxY9LnMvaIN7pSv6x9MTPVbLXowj7wOP
4xd+u/H2NTB+pGa8xpSehmh3TNse4/kYQZH8iWPFFDVrSEIk/vOEF0H6v2TzUNWTSTihAdR9536X
3zwDrw7PaMrpN4qLRqeASlAVHxGAPnlPNcoTZOObXTAw/oRKJ6EeOGHQZCMySfCtpSx5R7nVJ3qv
NW90wqY8Sx5V/2OuO5z3SQxOo0TwZQ2yl2r6pNaak3SQ18MSYtWFKTT4h9dNUpmmXQTvNwdSdlJe
Gi/UC0WRxHFov7AL9mvF+ysIYOKzXHW8GK4nS0T5sambInalxjMJQn9m/q2NKNT0zmbTTwNFZnPF
KNvUAPol5+OtYJqImD/5QMhkL5iNLCkFD+gZg8ky5FscCI4D9zYAcSCcxoZcSuF2d/ioy2MtWOAf
yWqsKwyFpr0wvYm+PxWIg2dxXyynrzBdEGipwtNEx86vCJkxR1y6Uqu/4GqjRBBE4Y5FlvFp+ksW
G75yOKMIABxKAwfgWPksRB12edkVBaiSpwDIJ6Y20eO2/tFFyo/9ZhYo2PjCOM51WcbcK/r5Xfr2
vbd8GUxa27oIz0z2WxiOFFCfaZmGyyk8FLOIbwYZKDGCsq7JFDNBSEmuo6zynWJrkb9dJ9/Pi+/P
XbO5RAyppjTcLZWQVLsK45Ss+upnM/LPo6hGyQvlSn/lhXBsgHMbtnivdVc2gFn3y7mmNoDearBe
49kWegbkj+C/E1MShKID4QeyNp52VhAYj8n/5B293/6hDn9LJQ3A4mVZzNQySrcFFnTLCDotZsFd
sNp/TfZdcNoQMWMlgP55CkCl/M5gErS05vFZ5jBuF5MHDhMpkVjLBEv3qwwyse5tq3Ad36m/hQO8
RXUCtYMTkVztDLchOp/ykuT85AqTcYYFu83JQml3o301aH8cmdXy4gbf12qxLwbeb8LnqWEhwoe5
WyUuqTVlFZhuV8QerW5cQjpoohkQctivjrh1AtyHUjvtem9G93OS9rNQFTg2DMoJuzJ3haawpAIF
Pmo0Tu/3xZr8/6M6o2m+7VXwDG0QRimt+YDFGVKdWMXwWySqkzn26z4yxV6nljIM6zsd+9WXU0X0
rUe1r8t/9JxFdVG9FaO3hzelA2MPhlQ62mnHiGj0JP5nambxgvqAI/6tH16ygbCWUerDF014QkJ1
hm0jJah3JgxJkqzrHThDBvrrIokR+mSO0nzyD4pQNqOcrILx94IE9R1MyS3ACd1Qk7lxQnVMk/ik
fNAVAe6uPwRb/zGTh4O7KZNAp7mNVHh8I+Oz9CDyhBkoaZSLKMR8S2Chynre1uIEWIxzytmUMHhX
58mzsfiPGPKhZwejfPCa9nk8GDxGuZRriSn/Ufl09HIBFFizHU7EFrPUwQSiHNQThG3kuAJnCjFJ
+GkWfI3PUUDj1TBPOZavKvLDzqeh9pQGlKjTw54WnwvOR6FqrCJZlnCX4rMq3eOR9sVrz57Mj6CS
LAUOCytvZRxcsXl7p7x1Nv8rikxEW87OeS/FDokKmf1yrGU5jC1bMd9to1vNL0S+/hdO+cqSZfxC
xh/pWFoJBJioZ1hjgoqeC+AES8oDyoQiW0DSiUMV6j8D5Y1mlJUmf6U9xy9Q1pf9loVP+F3ihTe2
xFeIuff0BT55PKm6yY+qPWwzvlysUZBIi8aqcd6/8DsQcESEH6MEP2wUBtZ3njsRiHTuDGJ8dugU
F2VsOnYxL2pprUFipnGaWSP0QI63U2YfqwCxPY/hSK/8IN/Leu6vQ5sw5egaAdgvI1TWghei9UGT
wuL6WBi0alkC89bMpiPgG6OLST+56eBW6lSGBY5UpsOzBPUJqCC2KLHpBH/Z1OqzkJMJOzoPlirD
vb1Sf2xhHT/iRbUmPCtJozyrZAX6S2nrLV4kcF8lY2HrNIKS1tcuEvAj1sCtymMx+VptPuNX82O4
ccL2Rq370fJTroBHsXclR3603roxivJUKMSOcPFtbx/nYMNKlA3fkkBDB1G2/2IaxG/1/66i7+8q
HnoKCzOuwvZnLRRbGae1AhfgKQCxFyh5463KGnFvWs53r5HTX12LAPC6dECx5UfTYZxe8V+nxE9d
gx1TcJsCb7IiIpoqz7G8Pwhtu/IGU34gml244CmuaXmnWlHB17MPKXUO0J6hfbsrHMt0+EdtG8w7
K0+Rz6ogeZJ5Y14j5fh8+Odq7qTDWDyYRl007k+BvXFqLKQ5mpIVXKFNEMj+X7R4kbU828IMfA4Y
p2xaPjx5BAFoIq5krN5KxYRQL8uzFEaiGUnMJAZ7Gv9eMgCEE+1L3+X1jUYDAe15l0sUF8amh+0V
VlLsAWC4nKYrttfcdgusxvdNpMoZtaA4C9yXF4Pm+4ntQCXdtv48sGnno1OxJKnhurBXyaU5pF2l
Zk6u0H7Oi1eVzFf31sp3qHQmk+JxHr0fOoB5mSJucnz6T8wUiYCwt73ArwbKqDy4veOsaAg/Sm/r
Rr4/GPMiJ1uAza2n2cWjHKAcw1/VoODtsCg/EAKFh8U7uZbCQi4IL/Yj3Efht3HJqAL5xkRie1Xn
nVfxEaxac9WHzPJwyzAYadULqsgiyKOp1cq1tYrt4c/V4lg4na5mKPdXAjoRf50sZU/wbxASqEfU
DxwrqW4ucosQWs4kAJacwAFifdeQSGoSHA0bRqcYC4kew+HTIPXl/ZGDJUo4dKJPixQ2tfjDnGgg
whA/nXVuuTvZvPew9jrTbX4RYA9yyTLm9Gpg2GhxU4dd2Ype4p3zPp5b4wvhZ4Vdux+JYMu4p/Mh
RxNXIOR+gLn5DsyMGraWnk3pf2Mj00oKE0WboKTNL3htUnQUTPszh0rjbrq91F2YvRqLjLFVL94J
wxO1sQqTKfIqmIm0T2KVervL6qn8Olu5bJi5kTDRI5H3gaT9scOG6PEJQ/VHvlX5AkSdTrshaUCC
bn0n2jOd3xHm50y347WeAclR/QJu9cdwynARTFzuCSikAJwYkK4jRylH4vb0OoSvEdTkSrtktaYl
WcvEJvrE09duKDxoYQu2s3JxPPnPW2ytOEPalca9DJQ2bW3pd2OWDX+HFoOMEPEa5ldWRRnJ3Tsr
YhxQs/IikrsmvIGM2Yg6pXSd5Zxq+mQzLGfJ6pSNCOwu00xV/4SgBk2PjEuDFivr8PXVRAiJX7/0
AFX53y8x1afb/5ELYdaBcapNVstRmudajkSJ2jANsWleSeYsaDDV8P9FFCrsBLrSSR3oKkv4Lgvp
7jK8BDaM1SdJFE7G2lhhKGqNST2Ee5C5sYYEOOn1iklEshFqqoI1f+OJLZbe3wlEm8FkBfRH8GWm
xuhAKqF54bzb237wV9KQsizerXapnp+7zbNzaHV4lZ/Uhgmsz3t/WXcodo4Ln8jr2k+SWyazhsqa
+fQv2b/SJqo9SKTNN8TZn6h/3/SOumvf2wLMzHxZwlg9UQ/nPqpzKG+mPbKNXbGx6N1i1OkRGI6F
TbmvrUhI4NiWZzAJ+TOZMxH7st0PM1+arvdNt0bR0RNnlgYP9BTwT3oswFBTcFgS/rbD6rrk8WZd
iQVIPKiUPPHvHocV2DXNhUGY0/1hWU2YqnBzsFho0SrzsHCZ9ILlRN3qOfFQSp/G5o5nm7Q2fHt2
ZwRJptXBg9cKs2fIbxZdXrbQGUmv3v+itxUmxtAycjS1cJ4C7ShQUcs4fiOqHVi6FwA7SY1lzk7R
y66OQtGrcPDLdN1ZwsgqUQ/sQPtsPRiGiXzyWPqcBw4oSBHnWCUYSzyx9Y94YIAaJ/OmiK1Wso0q
rdTR6shTTqG5fkF475nyLDknbwysUa4wVoYgWCONuBKqgXuu/THc7hSYNVC1KAeA9WRm7TXH25cz
ySqZpK6yzGDLKiPVGT0/pEIa0T4sbQ6oye8wj5p/PT+dM8w00OCYCOrbQWzjAN3mCf5GPM1oShQm
HB8+bHCblws2mutiEB2/9iqYFQeFoCklo4y8t4B8vEeMVgHRZHCUxSIyqSOLcZW0yb6niPozJdTc
4VYmHYHZbZ9qZ/wamRk7gS/w24vIQgIuPYAjQLeYEPW7G5HeXrPjPGtrs6DcjSbLrFAPv9TLiOTp
iVr+OKbLZz/vBwMRfxMInZeb0uktYFfSL0/fs999ZXPZAK1gPVP+OnGF/5K9JWNfvJPlMH/fI+sj
ft+c1oVpYMkhEzGwXTpjCiFFs15HGJSQbmI8Y/l5Rc6ieEtyJ1cQ8zYKPUQeWRlG7Mhz5t4An2+U
PpP5XkMbd70f5txxuAGOQSh7pAjTZY1bIWhaDTU/Khuw/350j/JqL2KEz226q99yusjubtJaNhCy
5rKGa3AArFpGNlqioEQQEQpG8rX8J195fUu6XDaYc/qMd4IOFE1MP66ncMB9Ukd9TQqwp2vcLtbK
KBAcRUsfdvnTOr4lf2HbbEjU1QUytJy736xsCSuIXGgACEQDW1hDAUtKMxwD4BZeGpKjpN4ukSYS
LuqEXfUymF9rn2K8iJ6Y2ioNQao3XG9E2yK/EKFfI3QipyNnQg1zJv/xLssfQFK1woIRqGtQUUTn
s1u6c2b52Yp4CbD6NyKu3M0v+m57O2e/72QnIpGEkKp3sKp3qB8D/+KJx33axqkDYJVCM9TDRWuB
x/FyHbVutYxxb6m/FVjZg1MtpdwK/RkGgkPxJLLWc94lOfVel0nAhNlHfIWynFtQHNux0o8/qGIr
pIcomswFCkG67KxK5pMDyHNtpdVDuMPjuVSydg2yQdhKFxcuRs8v3kmdem6WfpXlKfELEFoyMaYx
PuX2ovDKYKqzmko6onWu5sYxZ+THc2URVeCOW6v8GNs5VqILQ/FIzKKY4/QOYvoeI1VYbkX5Fq1I
Q1iePEGueNQWMRSeDyLZlnG9AF3BFxjow1/6+V04Em6jxDA1eotWozZM+6jFDzp+JBmGlLPHmn5X
3LJ/Jn5vaDyKcqTJXpvF9Lxwdec8UXdf0FSnK0J/jPAPPieu+iV4ESWnaoR02CgLItS8UWSJb7n0
RD4rjPQt4sS0dWI7NmQizw7IjvXs2uji/OXn1abcV2h+oMZ6/e2KCsgdnUteovwryd7v8FhGfcwt
529o+czYnqvvW3HYRWZEG7QnaJl7JXXdEbB9eLh7xYCgaubc1emt6+018RJC+IoK//iqR6qnT/yb
0ye0MU1PqghaX6TEkMiBQCYQAT2E+Pk0axJaEpOUuxipJkh3qZNueBUFI0jyvK42zvwNQYY1z6Rc
0Kt8A1iDtbB1Z2u6+glgcLsjkiB+3qZ6+vVr7fHRDyPKT9ptdovNsw1UUu+TAlYOM9JnaEXxPWDd
5OI7sQwFi6ee/qg21CIcoE5itZ+2yXbupUZm1uijN/2aN0ilOetREMYMiqsA2xdcoBKygh0yrxY8
M8Ce/Vtq4cbRyjlbovsg7uCHdhCwTJPra0XmBGTxXdFbTmX25lnIc7wZkgGkqwoWTR+i1wnoOSxi
e+KvWcuknVpehuYR1S4u/CFcqK/Q5OHWIi0IzKCUBKfaJRW8mFNNYGWvmiv4/D+8ppsWMoonBeJN
jJ7SGmzvE1O/RDCvccfz3sJxAxMg89zQ0KGGktOzBvWhELNFrihjtk6lPvvVx7p+uAthiBXhePFP
CSxC4UNs0YKAYi2ZILkdEOihY3eln1iveRl5FctfhF7DOY+Cn0AXW0ygf2eEHmQiXdxOZzfwTJMf
rwfh/3ZYaer2FTnBcBleiiwLBwRhFy9GKR3EPTqatTwASxbGejnw4vYJP8Zsbkp1cXIHyfak0oSx
Mxf5goQ1XAF0D1VgvB9+nQxRTcaEbDBgQyyHi4P8dIuAAa8d4v8MxO0zXG5h06a9Z6exto87XChD
4wK4Aoe7D6ZF0ZOZtTb6uFxxo2BNfTadnaX9qSq4Ly9jg5VkmrtAOIwK+DRmcn/H4WSESm2bfyGW
OILA8m0vqGWtCz4QLLaHFElSiWB+lgvrqOeu6vYu0BaM2d0JM4OTPFRR8zewiJHoT2wsGuPKKLBn
J+nXi1e0fYMRYXQSxyXe2JPRpf0f8jphewISgetsVfrmZi0qiM5Qv1YRTNZMg98EIrG4bf4L/Ld1
lI5NcCwgnSBCqOfD20z4GvcOeQ/tjrm1hD3WObL0khzJOsQS+4X2lmoknSUTmWIYa1nirGYNwNQq
gwndW9N5/tv6xOI0HTpc0M+miWkZjLvC/FZsLB5OzyCzHiYHQRGK5xiaQpXPyhSz0muP7s/9KmiC
X9HD/EJBAdCQVCVpaRDEBTwM/4iZooijZuqgW8eAmzoLsiecLqrC4N9MBQ6O3KwVNvbKSMIGGtHN
gvRf4vLHKBv09uAWV0cwNMzq9wqIovNhlv2JkNQL0JNhS5lBGicBB/rsLFv9rrLr76ruau94mCkp
4evDnt5H+hwgR0oWVprah75wzo95YN9vL8fdDgD2YNMqY++aguODqNtN1TpD7z8zN9UKLK/F/044
918qzjrQ7D6IDfUKPzNzguxAgvAt8pV5+jk/3w6+4jl4ZiJk+J2kPEytXmVF5K/hmEEXdTyicte4
sCLJuCg5NrIGZFYcOVWgkHKWOtS7P8L742h6QBt4FfmdHmhayDR29/yhq1VoASU2tDLRYDT/MpCy
OtSLptmqu35aRabqNznwrkTe0+uGCrU8+50lGchzPy2IujIxhFONTIUCfkE6Q+i+rPOFcUDuVb11
rEKs7oVBhARdElShEjTmCO/c3Fl4MQlgoMz12A9vJs3uhbF4hJhu4IHnXlI/iF6B8UqZ9uHTt919
HhMABM+GhmSdpGjPryV/ZJSI5UXr5ulRF1+fKzCuTios04Fi4MGknQx1rFGKmz8oUc5isxkAiMki
2I/x/w9TSH0CMl6eSC45K5zdbf+ndXakhhMRsY0eLqo1otjPSZlBp4uPkiF9wHd5EknBwICs33dl
xmzuUQZ0wZRCGm6JEBJAyFU0TYFGzOZAChgZzHKgrVG+kGf5Rlo7CqyLIpHeF6RfcjLbrO+0gMJA
F3hMNKaaDmuVVRBnPlyVibA+tvSRYF47r7JKcddEhXVvoh4N518qcGr+ibqJmnDRgACiUCRCuTkC
XgaJREVP0dRI63pcu4w7/xCGWXLoL0id2soOL/c/IBkPKaFRZXZfD26t4mAke8AMKpSYZyjV6MGW
kzkOT8j0zSh0/dksfb9XjG0ko4fiEHZ2m9E/tN0R+CiO4nPPStaByZy/qLSL+dgyLo1pJVS0TKEj
HrTo/fh0I65XStLpxXMR+WncU4I9I0Vsp0FSBIQBvAYn/j95+L0mrB508llT0JzYGJcgH831jUqe
aKqddD0DGjMfkvaIQScHDzB2oo5DAiwxCJAUq6/dW9zqzBlgAh8R6Dtd3sE0DLviwB1DUXBfB5MD
ue5X+zeSDDtLnEcmsCW8QLM+DXdr2DHG3yuT3L/AWAHZFjasinDxIXWYPo7G/3skkzzEKY8kalo/
OuQPR7NME55IKqwWaMT/Na6bJQVlaAoaoknvksBQMSzNXl3lxnvGLiPOgN7EOGfvJohzB+hP+T33
gHj65RFEXBxMMzLw6Pm+uU40GOGxM5TlIe/B6YKK7I/tXyQtq91qnpeWt37V4FbNQ6F2AaD8kx12
bRVVzZu6ktAwX39QfEmpIUHe2eCAG/FtR15/ys8+3LkXBl9xjrCgK0ry3fHrLp+8luiz1o8njcZp
kY2xpALkTkQyUa5jCC3qEziR8ksAmuvXQdjNlx1S7i6/PCQcMQTBC7gHDxmB6i9HLpsHGjY1GT6J
FAY5N1wqNryaVzWIyO5O5SZT542WPKk2c1oaDPyUaA6mUZGCjmNd6uwp+vfe9nAOZQzqY5Z0R4gK
EmKeYgEoq+F+M3ozk/Qk8begpeXrye3aZcYIHOUDsTKzbrkw8UMkKia9q7nFMQTr2yblYLf0Bw9+
6NVBtE7YhpJ+swHfIQ4+G3XRe6ucsTDAuNnf0xlIYLAOSpRQAIL0h3jiP/ODGUOd/d9Iaip70366
6ABVcR/eoiXjbHof64vOn3IJGMDm07PzZ7PYwtxLnP4I6aX23j6anwQATecyAa1onhOFIJD4mhwH
OJbAZZgz/77FebGvIDTQnLm/IKT9/crP22SpTd4IXnV8n4me4lr1zFotHn0BDVUhw+Je1Ee0HNEy
rmMDv4OUtPbTU64D3UA5AoR1KXJSUvaHP40h9Js3SgL9HkqIRQmzqcU+zW9mo9kwM8+CK1bSgnz7
+PS8b4hr0GIjIOk7Ja0nuiX+0Jla/pTymvkCYHZnAx1pE6hyIEjynYg/h6o4fHY5lO6qWhzBXxWw
BGl6koOvfEhZG6e6D6gjDo222bnP45h63/YZgdVXeBd9ReUo1Drc05tlMOV9rquWFTbYSo9iG0Ju
3+7kN3tIvgD3Kqzpky6Abofb+n02Lf4j7z/1GxJ3X1qkn67OxxbynBPdY9bi1uUhxSbV+hpPOa+B
LoNAuQIOT8qO32zoJlg9/QoCnoEd7vXLpQpWd05S+/KVdg5leBdK4LY6VH3YZsrGle0ulWiM1IAd
jQPc8GwClQGGARESDYLTe7+S57kEygZd9FeZBYzfQ/TjkpuiY0/No7dnKwGYXiBurDvIRyt/4w+F
h+A3kuEZ2tzCfTyPdzztt+81I6kSm9XueTV+dXpca5Knxhj6u1aAzEEL9kmx8i8lisIj97eeCP/B
AxW6jAmBYoq5HmJRs7Cr4g3e21L6U+q/pkZOuFU5D9911M3OTYDqNIdsANOurXJloSrSt9Gl4tjC
H0jd9vKWs2sBxueZ3UcLY2NkeVZQby587ApgHdxXpD18pnjZ/yt6Fpurbl11/xUJKipfttpo4ukz
RlgrQx7XOkARZ2xNJ1gs9FIm+rOjScO6sl30e+wfmu+mSo8QGTztqpEqOd211OioWUB8fSh3st4a
99+dcNyKT/LeaGczu6ikNA/zoP1+HD2gDzRDSll3SbY6/1GG8WIi6TjIDQQK5bn2y17ylzE5JDMz
D7C3FIEtvVKM48HZLfIsEvYVt8VIxUSejgnlEKEfOasu7ehs86fRa2THJqxe6UGyqSyarAS3eg7k
GbQKScKWMRQcW71TzVoMMahSkVCYVwmw0ytV+bMVJ2ruEyBoXewVwJgjdY+o6/Dr8+MUZ+yNLk5i
WBnqDFbTR2+x8/33pzyzYKiPI/tAKhLxhRL8YMc3lLLAbPApLZ6kbbHMknciGVdz4AWlKAXeZOgi
3TnPvF6gm/4tlOZijHcBdLRuxZEwicT+GZjDsWT+IsABBb6NmqdOlXItSt1YP5SbxfbN8SmQeJ3E
GQ5WpyMyB6aKT4sDLRZKlUWw5bT3zs+cdm39DcxHjWYMbruvmuWV0XhF5RbwBW+3wZp20iARkHIP
Mnt0VnuNzc3lIy5wrsuNnm48iDo2L/GyerC7A821OS3cTL0VFEJqI2hzHvOzIggOIuxWc7akoxXS
K+vzJtv2qQRt+uqznwPeiP7PkqsMXIJw2vuxM3bG7WEAuB54+m0RSrKRjRaoYKCJtuEQSshMPg03
dkYlJVIAg16IlOBGBhHmi7m/jHWAbD7wypvKAP+t/n+o+ZHzd5KD3063C5Y4+MmTjTEtuvQU+tAT
/6+XI+EjCQIP4TaOqTjWg/Cu22p9t8ix/L1Pf8RQvdmWy8u6X2wzhI8TcG05yDxs2EMHMPNOusI1
KjqUMN7Dqtdr9sxZQZFx8Ygfp1tc1I+A+mCp+ZHpfpe3aGd/BP0eLdWjbuhv3FS4Yi+ZWyE8++yO
Zqh5T40kvvz9JtRXzmuDb9cD0gIbCPNpgqh6uBq1Qe7gjYRSGdKWa5Rb+g3lfh4xdZaiErvSWshs
FQbyUvtecEXejaFyABlv+jD4zTgbJ5B4LHc3i3scfjAqOel3nTSNKNS6dlnNsNNVuVQza1iyNKr/
GbkXUgi3Hd7zVFA9i9in41olSw2Vh7Uhgc9Zud56ZQL4W/+mOlKFFtkroDHNPg9a0IDGMtnvyaQg
0JUFY/e7uQuLCZa4HRKVABIXzEajJz7mWHEgWuW4Ieoz4rVT81bo1tEWzuwT6yJaFzPmpApK3Ol4
JdLM/OhgZ3LQMfwE3sZFpbFDsDs5Ld+0QccUreuWBF6XcfSfWgMx+s7eRr40eTvuP0nEZC0TzDCv
T6SCg+Ylu1yc4UKiMl+fk8XaVFHSU3J+f3hJ+ZZWZM23K3vQt8vGsufLo4zf/CxxBb0BGK9vq2pd
EHtSc3Iurl/hsl84j9yOe1cBN0uAbjGNeExDKoqniMuvIozIjzZiDuGwksKqAfv7lsLhTvmJZqp+
YjrF11etAC7ztmqzhpo7UnmbBVU3dbC+PxaDyTtXDX+CLlaV59hZyWQtkWFqmHDb97d6AcfQvAtk
8r4ywyZAE/RtkXbgraZUES5TqtOClUF7Nfg91CYBrFzY079Ejs+1swfTrTF52V3g7co+OwaV9qAV
3TuJZzjqVv62Go8sO2Su6ymIfZwpwttXijTUVlrWmqdagFHuVgROVSFM6EeBjQy9TOqn/hUpnsk7
FdZ7In5ISp+L43gov2rncavbJeIcrLgB/dZir/MVYSskitIn4cuZf8UwUDCHmrdQhT7+wxx+WnjU
zavF3dZs8uqlyw2F8A9JbB3vgkkjZgUWAholuPJtMr2xq1VJbKoQr9qM/HCU2bfcQLSfesreXAFP
68SWpzns0FCBGG9g5wEAci4ntaBmDIXeLonjf3XWAweqvWhCRSbhD26K5/S//Ua23mnvmzzciX7r
JlAGblHISzoac2/9waH0zEeWuMnTuD7H2Lmn3TakmF3Uq/J3370bK+j5XPXK4IzhQJK+94XOtGJI
9x1XzRdcvdAOlNFUBPGva7zI5gUCcQtTGSO1SORyCrCAwcPByQkT7H5GuxLs4OntYl1QQAK1hAeI
5AUzkkYepdPmeC3wMRpETZ8ksMWK1s4tfWbBCA6jQMV8TD4zM1JJBwbp1fL64IUDJDUasJGb5jmw
M+8ZMN4CQI4Jxzh4f8Zuqny9fuWAOf5mKp5cvLZVhEWFeFOF9xfyy3Q9FqYecyOTKaejzDn8zjlY
8aLwZ8UCud2rYJVWrpAB9WRIa88fZREOzF9Tsr3CDwul1qVesFOuGykVWN0xtQrf+WeA+LGDgqUe
dv8x1TC7qTqWbo8xAiUfY0Gosr9mTjhYkIu1fcrKCflfzpOS8KdsH238T8Y0TidlCrusMpwAM5sw
ImB7vuQQun9OjlwvRIxQNzgiGd6mfzG8jH+zJ5/Qi4tiKt7H9Q2aXOpvRmVOiHXbSiGrYpbIrIWp
64ydxIefz9tyUIatd2kHPGRQPcbGxLblyswA3tzGvmQXQ4dej27ZU0/O/z+zL2+VecEXHmNJJCpP
hXDpEvQPgy9YP1LmpIAId0rbCxCHAzTnCeYdCgQHscyWym/aI5rMseqKyx0cXce2V43MeTl1NH6C
IFwJRZXHwURfu7n12Y+O3AoPV1p59GixO7+iLNlGtWt5RKHmOP9V3YIaUlaGfd9WzwUvL3kp0hNU
/kvwP5ADOasIxQ+9z3HJ1x5/WolyrDTXCbTK0aMa+GhB5SAFMAaukJalPEGYuO4jwnzvvpX3YmWU
SFJSRl8yu9NcE875+kPMXQTjJZi22R8UT22x9EEszS0FodXr1mWIIxwPh3Ydd/k3LRRuZk8Fi1ln
P9K4cpZ/KrnKjISDI9sZOLbG9IawLSvhPU4C+fbatFP3ufpaDFOq1aJtdwO9EcKT81f+zOqzlCxG
PwgOAVMqpigIXzwrNdlAJvC0KXWskhRQaf/I914s245kVrSthp/JQ0uInxt6+C1tVOvu/ZRIQT7I
hNINAFYXQdx+zPYAhfecj9a5QuTPZJdDXpz948U5KlNc69L9G2tAg1cWhjc2iFjFesSAOqeyPfd5
z37SEX7lCUdeJMtcwX5pwdDm4RwLbyAq+llNk+3XRNbVfTO1H6Ja9gY5/EC9VsWcSBLTskZPxjpY
uBsbOEig9jR0yoBzeBeZ0BPKVVWdAr4lR0FIdE76ZzKfQZchJvb9fnaGdVOFhHZmUN7/4vRplcpV
BAc3qehUu4HXYTKRIVDde57aVwVLsTQ2CupR1pEGsqw5x2+u8uDnIroWdA163Kt89qdGPyIMK3KZ
89lPNawMdlGOq0E3kUvv8P1PUR/XEgpzoScKArQ6z+WhlrKkMN+Pae2r6P2P/jusRRpZ7yT0uOvJ
+xWbY11qbABm6vF7Qz3wl5SrtpIk7+ZuUOgSlTDbkyABjUKMJvPKyTy+zqIaLF6aVNwTh+QYsKz6
Zd9+pXwNd68NV9cOyRI4dV2MRPPvf07NiQdDy/NixEERsXQASXJPWeuwh6kZPWWbobFqQyFCd07R
R5GBz6PR6YrWvOELvmDvqpDWWySLr3/Q7DOD7C0qjVME+Aa/wJhGsVWaX2348diUummr/JZyv7mq
NdbZ+JHxwXFhrd3lw/Mxl6Jl3+a7+lbeaJ/uN95hDLvvh3gj/jGEkxr72+P6AjZxG8gVsx7XHtEZ
YckK7DpkehXQJMnv4iSRB0iH+gM3W/l2aAtYNPujpj6RN8zIIiBnx3TFaOcKOHyfnxY2bVW2x7VT
7PAvd3vYCPiBJU69ZpI3ohX+pr+llj5bDsHomdMKImlPGaqZUEkRwjJmNBX3O8U4ZwTtUOVJ9cnx
IeZ85TT04ODfrYvX4nEYiscueal5LMV6Ls3i3TJLGtGnX9dxpdYVfUNW8R1ksWp3bwiEFcpyIa5Q
GhDr/ZB34MCLp1goMbVCPdhPya1ft5ZRk5vl+f9LT6ToB5HE3wC0RohrK1lkPkKZ35O+KNlhxv4b
2rvObLGbbs6jVrTV3U3I/TxprLTIWhdplSjd73aKUgAvbxxy+ORzR8PwSXYxUalborHjXKiKLJLI
hYKVp7xOvFaaWs6fNnLW2NiU0ccLaLSki4AoeYLordNFhthBDChkSeAw00prSWQQe2yIBvA9G1zo
ZisOIlqKmwuwfbj/Lp3auCWOEgv9MwA6R59kZH5ybpPE2rRtD0Q0pk90f+EvuWtD8McPjATywETg
+H6sMrVcT57VOJpXU6NK8qxB+iWtvd51uhO6AWzpXHo6gGVOVmrUn8tgnZBdP8rfgW26J4X3F16F
yzbNPfQQO5TBByDPp4fbKKdL8D1s+AVG5s9TdrEJkM/NX+S3A+WR8GXOY3vjEOddC1lk3XGW7weM
nzNFuZxt0qFI+KoSh7AD40kJSOnLGcM8pgrSZGVfCeTkV+gybW2XV+OvkinLL/YCN4XfjhByQ9My
U4Nx9Agbr2utmLLajGSKPQuTRhe6jsqYzD6HSGAuuLu86RclQxONri13TfjbGgqJnGfld4FvXugE
GgGz41B/lBKhXhpUX6AA3Pbi+trEhqwD9f/ZVfOzW1FgcCjACDUUrzTxJXskLdHf/hYZ165QmR9x
WLFi9BJd4B65sIfosf8Y6+5iiJl5Si8D1bmqbB2Eho+EX7Xcb4p39UHLTzp4Bs7Qks/XoII004d2
WgpvDxSgG5bROFv+1QPRiLvSgYfxhMrRla7GX05/C40T6vNL65t+YakgTmlWGMEuWYawh5cvSyMb
gyiAf3GVOhom2uPem2kILaf26rbYSChoxfA0oIpenVpqWnC9SaBc7EtJocVt2ykPInFDxZmoEspZ
MA+KeJfAaIWOjSKZt9tw9uRNWqIkX+AC6MmoHcPaP910Lwg0AuGdP2zrAT+/YO8rq6zryNn91laC
k3J0hhBawxWX2DOs14CG2M0Nlzo1+weqxpR6mtRCGsI2E0+1XRWX7ptpRf8e21htu9hMX8uBssA1
fKt3S1CB2uF/O0Xb9zkPJXo6c0+7ASLBoGC6VtQNcv+eqjF1vPyK67wTK7SFO8sXiK9wihnBeWLp
PdF50Unlo7xgOM15TZZD3x8OVRdZfSInovEsl1dYcqfrVSsqE0YFy3EIsfURa2FaUsAQZyEbtrWo
JXTBnr5yIb1SuPrNGwr44n6EPOSS3YA8udDi90I35Ok3J/NjP6DOui2ho/dNg/R12huprjOW3e2k
dGFvnBttXQ8O/B736E7tHDfXBUXEgStX1Q5tiNgPzdJMC05EBYRc/SIQruI67V4zi+kFjH4P4DT2
xwcS50twIXXh7X0dOJbgSilYgzYBBbbSYQ0kTp0V+WM+aTeO3CPP2v4a0GyLLjcJzToOhEblqL0C
OZEapsZexjIKq5SC5SkR59AeIJClStBzsmLshTz1noU33duZ8OV2Ek9uGop4wkboXAhv8Tje1/9D
z7iy4hh8iIIBRnk1iCurIoVLDmR2yAT7KnM+Xq2qVXoPpEdZFJ8AUDQH2yuidavCoiohPlPTi3D6
zzoOem6g5VXFyHmkp+4K+AXgYFro1l5SAOjtQQu6+BvgVV8lAg0q062sYZwZtbaYlVSW4muPVv17
J8l4ZC07yIN1pBIhO3z/jE5BFJ6clU/617DH3jH+ZMYNpOk/E+cxCh0cXvIEmecLevhAc/hOFURm
DjORTOd9jlhMYlOKPgqZGR76CwGFfXT7byMtFWT0v6JtZKkMjE9aMRs8Z2vTKReqy4FdDfvSfN1e
KywiIvSfN4ZCRn7Bsw63lvmklYWrj3PusGmRnwnSfho8myM/1BZQaH9nwKQtBDPWWF0J3yhaSt/H
AFaBsft2VijIqmGKOkoKBh3Vd4TTfT78Xg2BST3ecT+Ga4fIoB8sCguVEiWA0MFSWubL5tYfUgr7
WFM0p1F3vrovoTaImU2H59nmokgw/gpcPJHhR5V+J4gTitLM/8w4YUF+aZK61qpwhBWYN9viAD2K
HowJFq1Upr8P4h+OQCMIbPD/gzfZmYpPk1m+XRXtC8OhquKuR05Leb+8mjNjBl+B7zYnoduTfwFe
5Jf6B4Weti854+XVa90DmuWVoFfXGu/NtHVCKNUH5GG8UIop+hnVra/BfbmDAD0JsbilF+EDMjph
bFswyHCb82wKspweVjmAH9QE+IMzdCjjcCkXG9/+A00VV2b4SfsDyAhMcK2R2lS07ko2BCF7u995
rGSqcIIO9uszTkvPRt8udu61UABHraVeu9VPa1AeJIETrkYYJYrH/BCmJX6cd0W4I8fODZq1hyyg
Eme1LGwG4XA3fwDNwmaajTJcTkAY9y+uSsfTJwpPCQAxlCClU+nENt+aiia3JYCZnUF8QTW1zOaG
qibI3DSnpmxPqzsEo9I79prWT3i+DhSSIeKk7y/5wQQyhxSKcuXCJu8vzOxfRz7Q3vd1y2V8gL3j
0XcjfGkScEwkNCTvKZOUFGM3JIySEwAQ0fDX9OOLwFJV0EXSgU6c9TaY1ENqmMLYZXp64g2y1aYM
ZokbMv2tKhQltmWMr5dXoQM9Zj0eMMplazuKSK8PKPNhjUX6HztJuXGPf+OUp8XFLIlg0MQ7g3EV
i86l73Qqbh1G7neKK9+m9aE2agzHK3YJBUijyrk7s2fwbSAZDHJm06GZ3+IaVEesyXnepaOCmcRE
aq/t3w9yaxUGtqhR1lr3b2LkTCms94QP91q4MOeglR7CuW9nb3yjyTwJofrQj1EWnsWWXhD24Dk4
BQmqnkISps7iApHIktKc8fN7SdAAk2+BE9Onx7zsxTU2pdYmpSvSFRk6GYDC/blU5y+HM1ziwT4p
5ySvTc9zpSfvzkuLl3hyUPYIgv6RGJdQb/Bs3n/4jbEA4Hg/KMUQVt21ZIv2bJ7kNFiKmdq06dSC
VVnlaTMgxcXwBwPOgj9O/fj5M+UQkFaJOl8Kaxljl+DPlnPfhuijIk2i1VfJZtOBQz9oU4bUSGAf
yU8RCegWmmlbJi2r0JFsBqdrBHDoCXE2I5JeBfVp4md0Xmi4sZW3sNrOhWt5kQyH6680tmE5Xaa0
P9eQBtwGfq1EZzAvm7v+swnP88sLEH2zuCCQcTlQ46/LsmjMnVBlEgrwmFgkulbnGpW9VxnA2PO8
PvBD8WUdMAxpJGlE8dXS4gsKza1fs0zlbSGoTZbE4V4QMYSBO7Z5FJbNcVINm4SGfF0f3EuWaqXx
CvUvB73xqtlrP5ZX3YyiPAOWus6wNKp9Y5JPboSBSBC5FbEPK63m40ui2XBQ35j5jkE+2i09YbPO
pJkUWedSJdTxtnpo8h2b0VuTsa0zvQKrY/x49b6f4Ex4Zb0PP1M15EOJPqPl1/7ZdHxRZSIx4h/u
BHr+f/2bOOO7HOnXrsWnIltD/jQPpVy6ReoDJWzlWWRPE39ihkm4zWOdg1Aabl5fFvzlyUd8yoYc
4+DxsXIuwgbdIxB7ovoWWofA6s9cIMq8ZkbvdRHINPw+K+3WeRtcDFBJNE/d9bByeETJSSWj0Vi9
DDH7DypYTfX6/m5KFnXENLWjUsL+DCSEPbtj7et0GUY1aK9KrC+WqXDK6q++urHx5o7yD9Rum6kX
Mtqvy9O/LBtsJldD/My/fUhAdlfQbjrqn+qiM6GBFIuatWj1swwLNXCcz7SyIpVj5Z4m07nmMDjL
cQPcPpui4MnWpHL6KsP1msMMeJbi8DkxX5X8LvKB2pz2mMe3Cj4rkZU+akBuW4fV8haVuGH6rfqs
oqy9qHiEb96VsmXIl1XroxOLtMpL6B37P5Cb6qQr54fE/KAU3iKuUEiQXITGXoox5xNDhD9vcpdX
ytKuM2hAOjV7xqTpwKJQ5RoaWgt7PJ6MvfNt4+8ygeTjJZwQUTZ0t2iBa1381VhB3ElMW8fPAfi/
CFt0yckLCzDcIXK4CqXk0tTYfQcLU3mF0pTV/pyguaGuo4ZAi0pIC51VsT6kmCa9h7cFE71XVs/T
T9blgOFaFaCJLyRcIPOucILYUyPIFNoEnLoPtE1fL2+snYSPbWbsNfkuq5+0ls3ELXzjBjjZjNtu
wQIZqbk7Y+3IwkpjhBTYk+Xdk94oXTpEM9PR5q8y7hcaI4pKbCXR/ios/KFVNXAYdG8rpUg93N+v
vh6YJe6vK6R6RfxDEqOVTHF3SDTKdqHNCQ4NzN2ks3g/vRBD3xEFBNMh+IdYwMtKHETW4G/DXDyx
Ac4bEo+1P+XhfOCiQQzIESXv0oD/tMoSNOhRXv5j2WEOdDRymdO5Ba0loKNWU68RWCSXxNqS+79r
UIZP2TraK0EkBOuXyK57DA3nGJ/0vtnV12ARcgFietm7rhbtAFk7b6TaMfQuieXGF+ABgTn6iUji
tlR2ofD5VUvN5CwMkMNZIyYFk8caXVut03gFm3/cpxyy0RVDEQ/tA5iqXuMQwj4JGgdJUPwDzx3Q
ZFRRlfjmeCW7LiLlFvPWnQOath8EIQp8nnqKTf5r9t9FhfJ9oEDgXbXg5/T3/H3mbaGZr7MqgaJo
uPztN8QErm7KX9msqyaFseXoelADcijCJWZxaqARHqch3FkgaXkguZr4pz6CjiaoHnWQQOCe1kWr
Nmb+eL2YJLZMlnBARZ8Tds+S4s9l5Hmb6lnH/eKKtdNyEMEl5VwKuRZ7XJ4TlaMRCiWp6eEQSB13
xEwv5Rc+JNozj+SIGH2iO1YMYWzJ+63M0ZEFvKleANAj56uM4nyFCOrreUCixS2FSxgjl9qzaoAx
2kH4FgUofSC1wjhtiUWu3Jg9Jq+T36BWzvjtUFUv0Q/D/vjAxzqER2fMJ745YrWga6S+NKF89tbw
BK9rOUm/qIqvWjFIYTI+trVPEwMM24+yqpGWb7syFTuk78Wpwfaz/gEZGXSCUfjI+JMBHw0scZOI
kcRNxORk8s1zTSfpkwc2eiMfqx6/mwOQe9hC00dzkZBPN8595NqGDKc8e9oldXjKQjOGJwhY3Pu9
ewGzMXLyBV64eMh8g+itbD8yWheWzkoEpQo1p0y2hNRWGowcL4WOjxn1kan1FwjLGYId3p5JvfDs
aHWDSNyu5nS1AarMd+B3r7kAk6soO8yRbqa3ikMbWpA+IuMVjJ/p1lZtHTGEomTpGnyCchC+8qqB
T12gzAqAygw6XZp59+QA63vPAk9JIBWB6av8x353DYYrT35qVC1HyNuxrgnQfk6K8G4MdvWzCwjB
pl5Y7oS0X/rUSX8xs1mJVJ3uO1CLET5/GP0G0K2G1J6cnB7DRryFsMuWOeUCO9L9Yz0dG63NphfT
CJwocJ3tb4LcM3NMFtfx7MF74I/c2ls1u18X5gWQJqhgk4inwxVDWYCQRlfVuocB80bT/UtlRerF
oNyocByiXroc4Rs4pw2Ip8dkPLN9PsYj07lPSXX/4V9wpo4YcPEKGmzmIRY05PGY8lgj3MdqrvgV
GRJpSS6b5FYV1o8YtTmwbtWdMt+zbyKJzpo+oR3A/a6UIrLpTF8IvSEpOoNRylkgjzf5iFFpfVmQ
Z43VFFbmPnTneKYEc2aI0rE4DDF8V7b1AET4T18V/8maAxSCPWAJERAp4tUO0Pneh5vSEF8z3B96
hxIIbk6gUaaEvfbIzy1mm1UlB3ZqCFWNEl1gN9MYypCFDodUJ0446v0dGmd1s/V6MqhmR9Rrcal+
A8SikkfByB1K49Kdc4i/COlADqMkNbXDFZPsH4hMMrGqhZ5BBSOl0PrKui8xN9jyQoBF423VAz5h
Oz3KRrvmRn92LV9g3LRDZBUYtA+FaPtW45W3tRM4PFZ+1xB8cAKq/Ba1WmnMwlyIwcea26nfv8lW
YuUA76DLvF7fpI36MNexsguNSV+8SMvwq870OHdvEO8ngD8KLvXY3fc7V4OuyBGwDtuzYdO+oyva
23KHpt3BtNK6at1T/8Wu/qsgIQnIgGKGAyxUB5KEyXfBiI8s4XksFUc6Wxc+G331UIXF9mKgjvjT
YNVEBQJgtZghaOR5IVIL9lmlKWZZ4vC4CvxpvXwCmZ7LQeR8ecEQJLFOc041la8h40Q4Q/KX8w7q
58kXjnHlW5cS1n97s4qGi74SEBWoXHW4FsLKweBPFm33gzOgFN6WlRGwUogd+MenvCQFMixqwivk
Pt6KFgDxt2bkzKek0HLMJ/n55m3+/mGnAg/VbQbj7duFsH6ieo6yn6Ijl7SZ2ZmMoJyVsk4eTSsS
yuqVLSaMXHNrvtIzde5V9QRDi+9+q8u6NxzubueIe4+hwtYL3lsc9QHwgxcVLNLLR8hfASrsJA4W
FGJW7V9DxTfcVwzkQMZMm+TiGjLgMiK5b3FImGKsaIOCs2AKPXG3aE3L6htTjBiylQOi8vL+pq6w
3ZLAMj9GBmjy0ZfMqHVRLd8WoY/KlQdPN70zxhUrIdkgxK3qys2LsLaezr4z3dM+el9tvrRY4KXl
Et/+wsrZMAAX5C8mXUpGYBLacOoTTpNJxaailbyCqBAz2mxCbnkaqtnMs/QPesnQHX+6UKEqSO8t
hMlKPSwBnFed//JUSiWLNse1AIVRWkzXWV4tk0TnG5wG2lFtZfQO2vGXjyzEv7hO2f8T7srKWCdS
rLEa61X6SrVLYsbJLWDedYJDxFz5OarZT6qgx/K4tJNc6CR+lLCiV3TAkaAnCFFNnQ0GbuV2sVBy
sdXXHvRCd3ozUpgXb9qd6hgVYj/LqS6Y7YKn+V4MTYNEhhKo4vMxDD1Bz8GMFlYBW2w/c+12xrKc
s6MNcjwJm3AweCrZ8RE/HjC2xh7NrpCt7dhY0RVt4JMmVGvRPjs2iMcbM9ymtN7dgZVY+6Shqqg7
nMSkua+AxypmYTGahgYZFBltVR1qE4FIncp7wlhTILcUErO82sLjk2qjMsLmw6hnCFqERahcQCyx
ryXlNv65EvuMtio0xxqea0Zwlkf8WsaXsz7Z+1Oh3NaYxCuTcFeFaxXMgGr50G2b/TeJyw88uLHD
qpHsVwgpllF0PQz2YYHk9qQzNJx0Lzvyc/k8L9ivks61ai3E0WVyhwK5Q2r66TQ5OZiKP/6BUa9B
itTZeFj1XfyMbC3sI/OPD8bLQ1MiFuu66iCSs7gOweYcTnDLb+GQ3BSbVQFDnWrSDP1e4pkmvNkl
L91QWptwpPUlV4YAryYRIPmvLtJmjmuI9xnk1gt873JfbJ2ellDcWqfGyt/aXPt9ap2/vbe3orhC
sG3IjLGZCnF1vr5OrsYToGNujI3m45D00H1uxvSRrIdybl3Bas8BWAwgDJNk30RISoisi4FAPELG
/UN+YlEnFUKTs20Hi4+ggHxEcb75ftmc3WCO9vmj0D56gEr2YkDqU0eKdpn6bqx+FQo0XhgHyuh0
8RajXCWoHKqWJ2d1PuvYBgUTQ16JRzDnDAxEjvRnAKnnCC1NHIsIYnYKBgNzmRZHNKQhDYp5BXby
pRUxlB6eJPpfTdZZerOBxzDfwfdpNd3eS+L3RbAJQs9I2AV/ZYT0yZyq2uc4W7a/a+gxmZ6Gv7oR
vwoFlzRLQEoCDQiN3eRVR60CCz/MtpTTgOJJa01qaYM7/F895qZkvQ44yVp2oT21Y98Zd7uBupBu
Q3gZc3ZlA4vROpdcMUXg6i0JeHEiDmYmRb0Gn+WL8+GysScNg9hMErBULuN91FO2TPFqe6VTxxPH
kxLpyhtrCAvga2uVJdiP7xNJ7pyCcebAWKAySCI0TOcE6nAV0bHJMf+wQBkQit43rpU51yxURqwL
9oPG7ZlvhmRixM66snIGW2NkBRyXJiawXCKs/l7+78tJuNYrjtglOayplOCIMnQman0iijR8p9wJ
mHj3NamexMCpZt30qtAB0/9I3H4Z8KiHHx+FZmY606KN/SoNQaiLtwtHs5CxTAQ3QoRQO/kIcJh7
iksZ5ogMIaJvkaVJcJvnwmeSBWdcHTUvLHyoUNlhsn4nZ1MHZ9bR/h/WgJAUm2OZ5VXZdLFp0+Is
lsvgD0GGdYQ2aNXqxVWAuW6rIpOztrw8QQbkSvLyRHeVwGTChopMza6274LcYtRKSuyO1pNoUC9k
eoiF94ePBTiiJRA63jcq3LhC4O8rIvKn7XxSYI3sHbbVW0ZZ4ehOOEfwCIkGbtFL7jM9DArcXKUo
To2L0XUrM9j8oiXocloGULKIxflALjnp4H82kOPTinwpxlTL1b+z1E96TimAL3XGaXPYb6Ydyijv
k0WAjAH3u8txpQnSRG6xM9IA6tOWbKmW6GmGIF/lchfR5G0tG6ytkIYp2QsrQPELhuIBOnqCXYnb
Vex65dHEFim8eCUxkYYqljXzgAnXKpt4V0Lq/PAlC2f+rEkWXttq7uRhbAUMPwMsMhmHrkO6L4u4
WAP8zVzYnKqvN5TnzfpJtRYSF1++nfPLOpYqCjLYRhSDp9bJ2GIE3ZUK19xt0FkV1+KZTUHFOjRX
BxAfrjsnvstQPNz1W8ez5SzsCZUEvb+ELpqy0mD9wt8ZmjxPenHgheALrGsnbIA2a4G5kNLauVrt
SzzPu43tiY2//5sBp/sr+3hbntcWcWaELR48xZ5lgf0UOxFSCWYs7fJP5xglRXAdjzQ93r+Qbx/G
u8RIAVFeebAvP/osw7XcuBEQiALTUvDAMLx2LWsaeVOS9nf9D4H7CzWK048/hS332Q29DP9JWrak
NZu7IoD3AEwjiP4k+NSqQQMm2tn3gOxIYwhOlgsozFpMmdNm6/lcwpejBw8uA9CGMBmGNKHc4eWs
d1NIv/A/gZpg1GvseLDF8eU06ig1HRkieUWWxm0GiBHwxxucTpAaZ2bqPASKlSn+n1s9YGgknz/R
NJpwk0ONAxdT+gevMNGyAb4I/fpe4J3ez6JQuUCUlKdNpGmN6FcQUtKIUbIwH6iKjR3snWymzrFl
iDyzw99iI2lOfEeVh4fj8veOIfo1eApJMHPPpRtw0iyWXe9Rc8sHIpGDy2pBXBfCyrKNJgCbLGom
lHxMMRKEQ2lLPVFbCgmjhnZpfjic7Of4YCwz/oUbFR3I1yviGgR+X62q2OdbaPKeAukRBAZEZetk
PviStSB9kP2xu6ZCdACpMxU8KdjcCcKLiSVOjrDUy9gtpQzxlfSVGt/NL41kpM5YyAc/+NIA2W1b
s1AEAKKpqytPsQUr/lCJFLQDvdj/bjm3WgZ6X+OsceSRDcQk5q0Vk4LrWi9N2+kp0oA2fWmaMb4t
hPWPrgd7dP83+LvRKRtAKSU5zfUzXU8giJcz1fsrfJVNMSbsT7XRt986g6moKQkVnRgmgrVQIj2+
zfz6P4UuVtzvR03NpJ4+EZhjHjnxwOtNiWdgSo1BvkilcZtLpWZBK8m/7UP1Sp1V3FCk8U+HETX+
fs3YTmJGnZy6+Q7+dcSNCj3YbFz5D385fAvLti6FMwkdBwkcnVrjKCM2fsmCaOlQD+d9ns4bp2d4
du/Wpiyz2eL9tvQtdhoP8Oug9pN2ukqWd0vctGO1uuMamdRPbWTC/JI5hMLpW0vOlCVCSPX4M2Dt
j0PtLTb0GDV5xZw+lXunmMjxz0DwNCXxcJn0nPjGaMc3tMRlMTvPqAvMTwP6P2Uf3pj52092PBj+
6R5SiE+6scTQNE10HwAvomy8C3pAiKXZHjW3XYb9dXj/2WQrTOlDv9bwWOhbbFu6PDP4QHW8KwS8
DkEVDkvUo6+TcYPVLFBjAgRB6Vlua7OCM4WWlsteTmmDBOc8h22GY2RLykrpVi+4NKuPm+xKcaQG
ryG3ArqIHZzhXv2JW89MFrwVZfQEsEGPfXq8irvdW5F8hLJHj4PjHmhQ8DQwEK5z0nMTT7i+IAH5
hO9vw+P8BFPc4v296iDgAG+ejgORp595eSTrfwXxgnK2k/+DiLNCmrNK00eBTgzuRUfR8WdAth1j
UUzmk+DNNNngIXOX7d5EhdUbIeJS6BCf/2tNN5fmBO9SiIdGAxcDjh9IhEYMjmDXmbqsgRV9yx1i
IoL+aii2R+3/td4f7H4x3qLbccGx1KkXGphLKWBiUcySzjISXyRBbCqcHLWD44EcrIfrtui8ucz7
7Gmo5/rtgYuYax6tuXc6C/bbd8hG9v4JzryXi6bGXshxUj7e+MSUuO9+9ZnSpUVeScfMmuRgSgIW
m+jHY9RFOPWykyPXlGpJW6XHbqxtLcm6TtupgCozLyT1RuW8kf7gmZVZ7oDJOoU9QkYoTOsmV4E9
zdLisUlRdSG9yrePDbJp4y9Wpqd5iOdrxlP/tTV8cmDcHhkf9lcOy8/ko12hvcnYmdHHhbp1MJZe
pYXK7uyC+Du8wLxpsjb/dpTjuEG2qk7DN+yS+2lPf/eifTGfCSnvTIt4WUVhI7mni8HzhCj5NyvR
MPDhVM8Ulv2YEg8V+zW7gijJwsWbFYZhDZwwob/QDSxtyQJaJR7a4sXDuVtlegGO183xlPPhjHP5
z88sRGlScCa5KFedYXwlk0XnOIHiSTsd6CAJQ26xrkJHHSwcnwhWHXYLT81R49l5nZvNO13jl7Gm
gY1Q/fpAbFE9SVSEKqmEfRZoMsLiuQJybXwNPdMHxla34XdozSLuefj8w/yiIklemvLVriboYB6U
pEYTe2r/v/Dc4mP3lIrzG6z4N0u8085EGi/jiLXDnl9Rsh7BPb9wD3XzvqHWTEqP/S+b8RIUHbm7
fPNew5JYdNcdvPgemItBhAyAvFo/2wVQ0HFHiwVAdGxXOfHeXbkiNs95MRa7/f9HWvknhwigMEmC
FuMMRdFh4aqJymhlXBJ0uGeh+W8MRvFDVWAJsKxcHdB+jE5N2bBgw0l0pm7GnXi4kU60OYhFuLYz
5LTaco6a/rGBYiksjPNvw9SoZPl1KMR+BmVprbUrjUTgzwWY73I1pyuSjrvCp+8uP8M+mvUWlwN2
bwEwBHAEVvqt3BjXm8ucV9LIaOyXExuRymCNXATMMeSN7fa7XvFiYUbaQAQExDJmniMQ573GqtOb
H7Km7AWJ/RQOzIa+h+WParOD2TrIch+LUkw9KpusU+VccpPwexQfqTWpvJ4zTkyO5qUAYc9TTWuc
5F2NlSB9Kr0ZA8FDKpy2PYDpSHFcKX6v3viZqyzn853Bu20Xcz4hNPlJHo8GV5H24X99hR9kUzKS
pIdY+ZWvTb3gUGbs2h3fIli7Ti7XnyNpUNCCz7yhGVy8pAAXdWIwJ+Sv8C/1hPORGgd9iyCMXGsm
K0/qenZ06fCDJqWgHwUXElK/wPlgEZ12U2G/lhBpWVGEPNc81ssEd9XpaJx5fS5aqyIraF6cPESL
Nr8jMnwnHUSxIuXtELydOhO6Sr9uDtWnu9s020IZinYoOPTxB4SoBZsw6yuO85Z/HuvroI4oCpGU
bc5wybUUe0yS+BkA1YPxJjGO+HuUvm4hHvdUD6x+oaSWnnWcQpMEbQhiapc1VHxzQjyDaA1cmY+p
aZCdNlJbJC2mxtzXrnKKLGw/zoCSBVymgwMXKr+1jOqKKkNnGL6F9bHzkmesQimdhgAVOuCGZ9OF
8QCbPOnRioM2Sv/v+7dX6X8xrvFI7Ym6yW2s4KzTaUFB4WDx2quIow0U91V+39fE2+V6SQQNTsdi
cAset5rqiFtTzH4TwJja9qb0wOPuKZbLUfn8JpyY0PfllFkKkPWahUFTfnKQXBA6IQhvDHZYVeVh
WcVUCXM5zB5L8hcdWenJhYbDHL2s+ntUV92swrlQNOXBRJq+s1/UpFPI4L6/Tz3CyFJpDhXjAGOf
PpJ4tXfaYGqFXrS70Ss/xoY5eKLKLxOYECW9ir1flYBRpLSodkcGYuYQRLQWu61bT/k9zuBD0vAy
f5csXizl5Qp0Vhymactj8l3KxLdr3AiMAz7VzHsznFHlA/3ydHvBHLdaK2xtcNUr6F2+qYliEqDB
+4mYyR4BWging84lXsKyXD4Ai8zROoxOgWDBD8dhtx2Q4pXEoAy4fXGIEKOlPbETIOs/mcMdosxN
aLpzkqsVoPYGTTVocD+oybYzmaSGML2UJKSJO5nIGkGpOdBU2G77Qmn+NSyMueQbB88IW0qtpbdj
VYo1yHdo+O7brb1Dztgivowj6wX/fI7pbkeWss3a0FjFhEeYqDXzYlt/9Y1c9N9gF8YpIAyuSOCJ
CLKJSClzeWwpbXCCT+R8xdN0TMuWe/Olcm1O5GyztojJXZZKhOquAW1TjmlNw9RBKmi6wzhkKZQ+
1EWd6TO0HQwvCCta5Yzwx7cJqcTW3m1RRGUlqAjucqs1AKmCSfuC8MQYB/LSen4dhM8ckLARVWtr
cIEAztXPX9ruKrOPQHZF24edsPdP0vFUE7d6jF5ipR7OY1XML8e3o0unEVugNAmB8qanVqGxCDqt
ptudU8C3ujUkt1Cbr3XdVoxjneAtlehDeRgE78bZcWJA9JzZAqh91Ss3le/mMAg090ElB/PiDyuL
Kg14YvafFzjxudKQLyHFKZ287528vwqW3ZVLXCNnF7+hRc8c8u+qHxiNQFl0L7nkIQax5iuwEjZ5
3evBAJaMRcNjClN/agDXaTkEAm+HliY0zEDRdCaMpp8ruYFDv52tJeq93ju7a3HE3hPFGPWebI1b
OKBOaHMsNt0I6f7mLvGLwHDIwnEFpF+8XWbxAWAJ5lUB0wllK4trtixGhimXQVIHRcjPgEqrzmbV
3xSOAYkeQnXCEsewJzDw0MIZfCmoZmUWu5iaAs41lvPRx2ngWJyw2Bze22Ope4M6wVTOL1VmK418
p7FwkiS1HrFXCPVBCL6wnCUdrZwTEJ50g36UxYjs5af3Qw0+XoanTIRM+B716DLJ4y9oI/HMJJr4
dcJ2m198RJyi/2erVzZdWAMtYpjD62ym03bQ9QQGg9EXF2UPpw4D4bD7f0jsL2o40+fW3pRS4hLf
DMIPaidAp1APcRrnCkTU3Teh0mLUOiQEZ/RroHjTjaU63SAISDO5z+ngRp5WMbnc8pF3W3k73CJN
b8kRTjNmLfSugr3ujV7EsaaYwa+J1DUBAwCRPzUGXyuYyIqUTvgpVY5zuWGvUetvLhlvaCy9IUU7
y5BuAKpy8gWBkC8hty9GdacTT9ht/AgOflhPN5HjaWrPKLcYvWjFxMo4CXx2Fv12isOXtUZ1/l8b
mPXQqyxxYdM1SPmCEq3lr/w/d6HAAuuHyeVTAiwEyhKytd9nUj+FJBu0DOMFlBt5Is/VNRX4aDQg
iWu6tFggJcMaN8Ve+qTqnNNPa28C1u30FPvfl9wH6POWEZ0ttwEVMTZHdpZpzgeHBcuNvN/INnb5
ht0qXwtx+1PaVgVjvsSktXp/KyDBYwCm95rUqkgewNCqJX1s9vrL9/3f8QCz6kvSsHGkkRCJVm1j
jIgFshh3pz1NU342FlQ2zE0e4I34mDX0oIj9lGCR91h5YCL838HUNe7YQ9Mp3ycjAmJz4WANKGf5
UcSAQnKSVRcwLSaUwSsxFK56DpVgQvzC+0QIzQd2mwAaim0CRATnPJlT4ck6hJJ8T3Yf3F8GIyrC
K+oFQith3Maq9G+0SOyItLXcIv+CC4dpbS75lLKWBEvLYABHWN/7f8sV+KnArAiNsBhyok8qBJQ1
Et19ig3NKX4EGShgQKDRcxZzjlolvRn6PjHa2P4y/hnRxjTkllObiY8ryZUcLSCrEx6exHP8/jxp
JH/vSEmMe6THWaig1pCstXeauwbnGnvRsGJLNaii4CjCe6ArMvRHHCM3T9zN946Mrfax1ZU2raG6
H6pM2FxbCEhmrVGBXOq9LMjdqwGhkDqvhk889H9SpxwLBotizBJG/aXTshWUXO6ku0d7CCcowuuP
XS7E9n1MxHEGDsPWuUQIj7MYsapj26A2/ZpZR+7G1J5+pW4F5s214JiddGZ1LtHEaBvFjVDn+D6K
tMXoQqHO1ViPhMmC+6zuN71DmAG+qB4x7ygzi4794Ct/E0dl6+YuElxU9N7Av8KFoNnWpavd8daN
sRyRBsTckwcCeKydqTbNGFrjtL2MvwmRzKdkChwXt6/Q9YMHpAb/NVXDpdasCDhlql/QVIRyJIH4
zv7YRxCh1IMb38xM22GUs74/6LiTiWNDMQPdS3mJSZhaeYXLAUAoCKCzCS/Oy5CxAkI89w/lz0Pq
HF/p5PEaAk/TG/D9oTLPtcT5edAhaadGDr2S0Bee7mJa8/9j8ExS3QBqpCqu+DWsqngA6bVJ3Tf2
tsDffozrBE6vv/gDo+D8UuVMpMI+nPzzsIxg/NHyldHaK+KIzIww6hBK8wZagm7mgSOsTehcYzKK
GPCntHQQPw3IiYKXkgFUAx7Up40eGqYT4D48S+epthnPwtLcuiOxXf5JIkOK4RkNNMpIVbZVoVo6
MdWSUwNMCaXp6lf1incegwUdC8s2Zbi7HEQCd+0DtKgeZKcn6gujEQncUq2uJHiSLPqsH4/nyq3z
s2fcJ3toAGYUbQu0SsgIz/DLLNfD3fnN53SivwFF0dAFUX/+OBHu5xksQPUw15h22jp60UOCdSEH
RLXR/rGsIUQ2/lIzkpN7F974LvfW6blkr1hroyF8+uw1bk6mO/QOFf+exLhzNyMs+9tzg/6fjtVK
RRDj8ZoIzZp5iChwvCr6fPV4uCV5AkObLvdgT6mtUDVraLbqPeUVd09bDe46IoO3r36MWJRvxRB8
fnOs7z7pwJ0mmCua7MBrd6i0LRnxr8ZVxSPCKehc4BTVAY1+m8sTu36z/7tmaLHMA8vckRX0oOrw
EcYdMNlzWLH7dLhd5ayE5v33ymQ4cNaP7ucAxs5j3kwxhV2e+t/969tH2Li2jwtfQel8VVm970R1
9hCdG2974OLfXSiNGTr/WPDLM+BZFwrA47HrmNZE/7vZzlg4sXjsIcot+k3l+K3hc/7LDNZARkhV
TcG7MtjgA8CMhmFBb4hszIe2SSYH+u1UBfZMLMY+NKxf1blGMO76qlRrJdmNKhoEkTHQf+l1NoPZ
jEsi/QIzJyW2dgNeCvlAS7j8PIDNNY/+IG8yVIqnE+02JSkPtIgGKM74nkVJwa0XyFggG0xt6pWc
x+WNZmy5uVGuSpqwELZLr9mPfvJ40IZ7t55Rk9j00BEjV9ewTZUSLqFHX54ZE9rJ9eI7ABAs3w9T
7ZntJ71rQAcms7GYcLiNJ7xw4x3VF5O8eDMYVxv5ob6UIbudqvqGB7Giaat/ERiZmk7Lom8F/WGQ
53YH2lwTLPB1y+CaVthkLKdX2AV38eseVouwreH29/uWt5dFcifKkki1GAKLZ3g54AmHeJEEUQh1
cV3ggxyDkQQuj85k4K9EVomeS2G0Wo+qKEBM6bW3NbYt6GQv6alQV6pUnw0SRO6yCstaEb8jHXF0
yH/N6fZcpDxfwyTzjQ3FwGhS47y0mZAZVnECeVFoXzd1QOIDaLLGrPCu1AVsymdcFS5iaba3OGAu
8xEcQl1WG2Np65HesYSZqM9I5YxcFhkDCishE8TzX0goiBwgyCwZCA5UBsfO/cl/KJJShQoKz5eZ
hR35IW0sKLZu9Tv8Qggr95IvZ3hfQxNsvZhI1Eomf0LvcoOqb6jgi2+Hw1SgXzDWmxUhnWa4NBAI
zSiELzjYFOtEJZ/1lZAxAo93N5b3mUfGN+gLdoUxz+YPwwe3Z3eJrXaCP5YqJi0QfrMFU1JpBKDc
yM+Vcq7hVGvRcxX7IyZD4fVCRy+NtHxSwT86p3bFXJ0AIyS2IBWR6fsES3xJW0jILgFfoS5LFXej
aS3KaOxQjYQhP/uEH6LibZjQ0/3tdJ+9wnyS5MZZbH/N3fTLyWgsVsx1f+vjsD2/X3vsC476/Qqp
NS9YuKZ0ZHM7FAvxy9WuqrZJwxKEDMMZcyVAZS+A3UBloZmyI+ImVZz1/NjLo6Go9SBp3IiNl4eL
HSOAdJG48N5cDc4hq7kNibn2tSQDO9V5SP55gzy6KTqa1nGWQTdLItBcqkiqMKEyxel1ni+CSyrw
ZZymgxQcLk/WqVoelYW7GxRetRtyixF6rBws7N05dJ0e8SLpuKSEZsm0l/LLOFD1Xth6l3AuAbPg
gkM5YuzbEBUxpoCy/t1n4cLqbOXezebesrUMahGH5vYa9mr8k5h1J0BJZeL4wY2gVHJA869ZoP/y
OzttU5MdGSQIQ13g5Dt6MCnX7QqN/Kn6T26O5bfsPDYWdWT2iuN0wCVWjekXUKD2uPeVkKLIB/Jb
PZkc3dCXdU37tg0CNCF6r4w0KLqu6Ayjm1QNiiMklQ0B3AVc6aaEkI/UMW4MByfkHNKk3Y60wXjR
qmEkColKpSwVh5XhUiiW3+m4C2ytemGP6wWPAEhL4zxsPvistkf2TBqt/QkKdBSc8N2tHRkj5iI5
bC+1xgl01XiVypr/tFejTIyHRVhw8/LYl1C78laCwGT2hRkrt1PC/WUDdwtVA336oksWAVce5rAA
IqkncMWArzQPFqVWAkni03oGkrhGZhrSheWS4X4Fq12H0xXygKUX/Xz1iL4H+XzDJlY/fwmC5/DS
g8Vb+6Pmz7kliwE0tAUG5KM9P5/67n57wSUWMhHizsrq7chkyudzogVTg2qETWO3IDboFc917wX+
FQki7crsNTBxI+yj02ZaVoNKZUwKkpucxY121NNi+erc9L2tWkcyIoFx/YqMa8HKxquzoFox94vX
YoQdJQwAiHYEYzLa57PC0DWbOayq3gdxeGsZCMjFhubWlJR08DIxkXxhSRkt6RPSoBmo7tUYRaMn
SfUOL0Mp7T3R8RolTfXIWjkMmyRbFpz9VYGvPKm9gio9XWvT5kR2V08d3o58sAu2cyKgBCi/KykR
EIy0AbGxgT8LmUoBISxGa4el24kZ4WGI1/D4WmSYBtIFYYFzVWIaasmzV4JArJScolgdG7sv8p7Z
s8mtdG68to5UtTwQ05epOmfM8rGsMGYmwx0A6C/PC2XX4fGOPmiuUQGj6U2y0k9MB4QRb44ZxBgR
jry1gmQSAxGm/Qzyh5L2EMJdUKfrt9CjLRgAPVPPI5Ed4EQuC0D01A3hTZfGXD9t1pFXFzHKuKwn
9VFuVqp/9qUCUWJrRL/9iFLHjr6QqSq8DWyal6kFRYcd6FNenpSbZxdwWJDvMa5GuXvweZk7vdpz
Nuuhz/RsGEauaN7MdKHRo7VhMUfY/zuwPCBE0qk/W9WGqqYc7OFm+T5zp3v+7HZZ0OP+E/SGa5p5
/Y6GBotKtxIztkrC2aZ/7kwflkk0kEP+JQWiIaANh4KTQOH6LQhGBlLfjN91zFE+HFkoBBs402oc
50t+EslOlv/JerIL0nud2emPRJnH0F1oBCkAP42clSars2ipOz/1R6sz/DSE9/fNg+g8LyzChKpo
qU/zIyyVGZJ0mnjF6nUeCs+XNi5kon1Bnrm9+uykMtADgD61p1RISBLmEC1VEHA2Oa52hl04YLRL
4rqyxhYPbPJQ4lt5VxiA9qmrnPww/gL9aH9teXujXRJ9uFysm2CHobhvIx7uCKOLVmCsitQBgTld
HcyHgGLE2xe92J+ZgbYcVwywd9HYgo1IvaUVdCq4g6z6zz+stwNh78H16+R7eYpyWh+Hb1Vq2n6D
uFYkGyiWo6o194g1wiqk5mpj2f9NVEw9U6lc3YzGnf8S7x0bg2+tLmsKgLDpKn/V0V7xEUkTzmV3
GYoebOcvZsiR7ZasvFZ+5DqVE+ZBmZWdZMMTdqTY9Cg871+xW+dOVu3MjKy+0z9BrF1PdhFyuGoh
Na21qwIMD8mQw1H0fRkzW2hwIOpETjgiSCKXiGe6vW295AQmP9IWvHQQpy/ph5kqya3BRgV7MEvG
AydMSU5MGdEXi3GoycFsPuE5W5FzRe5EbY/4nxdZ2QAuDuVn86mfSjI/+IDcj38CHLA3fXmCCNNO
CuHIq1eItfbQga4OUXfAXhtzeWRumqqESvwpj8ASeehXvNpI35n+0+Gtv0c0/39KGwGEcxhLi/Ay
xcUzAeALiwjfPgzq/fNyssXRI1b0IVQvIiAFQvfR5ae+MFR3jkW8YHtu8ak2Kqoq3+rCylauP7IX
wIzc8pT1HFnWemQYEaxkVhKg8Etely+bVwCKdJrseM9clE3dz+q4tnjb6xws4FSpOHuN1LXYuAtc
/vYu+7H66LC1tJElTfGCe9IlV4x1+WG5zKtwXDlP1wdx+6LOrIfm6xA2BHKhJYBaBl33qy4fOp55
NPNCTgPnPIP2DNpla0y9dQXdaf7sAjyA+lToj+ZgeH77e40v/ODNsqQBm1YgsYtdMuUJLIDHGFJr
cDmVBuYYdzu7zFUh/M/fQ4kNxZvDdgLQrQk7KomgTA3ZU4AW/A1CR4jjeBOK6mP6gRCj1yp3mffw
NbIZZvbxApZK0LcxVVq2f1AAhMQKU5cz3/TzzmSqsxgNQcUFqAaJjbns0bZ3pY2D5wKQ4JSoAVS3
5tSoq3+xaCwLCK9Cn4pIhq3OLeRJNb9QXMMxRl6VMHzTT6hKoDUJNJ8EzJCHxkuJiJkiVEj7NaVf
+wV9AAYwilxcW0iOOVzXt+Njlv3cl8DaQjE2zYmjEeC3EI2MmUZEKXfFySpPO2ZqtPouOFbfhXSQ
Gz45byyg+OJNamNzPg3BMItFUN1a7CaAfnJu8bjiyxQNuE9J7mN48UwvUsvpgdZ+l3XrwcV3N3eR
s0l1xiBtXRYl79cBO3SI4p1P5vp3dx+uDQphmSMhBbWKbSZ+mYWUVvchmPqEU3xajNISVaQNuHiN
vQCq7lCs35Iwle1hMhYNY7qmKZzNwnXHVIa+XDciMgDtqFDNT0J5AiSd+XQ6qmtYH1omdFo/nL+v
DIkG2NeQFzX1Q2L5D1p463KgnyLoUFMoiIkp6jb3hkWOMINHs2ozR8gCWOxdOiurifsj0O6jDCNB
03ciDEE3t9u7R70My1IpY9U2Xknvmw/sqvocJRI50CE54fPD3PnBYLM/YFPDLmpFLmvQ2P9Q+dpN
g+xzqiAQnnVXk8EesgyUJEp57ClXaWPRtLrzFcz8fnuCTAOGEB2TSlvOQMQupSMoGvPTWsqhoc02
CBZ9OWjGT4s9Xi5XWCJ7b4CeQKD5EVFB1OeJGhPZW4/uiVlGzpsVXv+cC2+esZVneYnfoKdfCMgT
3WzZG0l+tbTWkIImBUVBOMeefG+tL8kwdnbis5qLLi0aou+7GgmOOcELc3Kyp7TGbMxDE+b1mOJd
sHhrRB0LAxflo2XRbLel7+g7nZDIteylC1Ux0gAgfI0f//g3ZObpZmtbrXZuPKsUzxbpKjPSNPPx
AIoJPhDpzZ6prw7FCnnLgs1DfLzQ55OjveIzrnighZHpB5pGxCM4LnsykAEVhFQSt4jfR/6ci+X3
IiQw/ItjYvLutekZXu9IkU4VKLpEZJ0ZMff/DOgb+KViECNQXtHMFsSfOr4BUajtcXKIqY5lw2tX
IjXXDP0Ofc5epIReBd9051XpLfCibPjTfCMhZ01Q8ebtv/ddKoaB8xHIQYdLMUxKhH/6o2tXNovQ
ZL+4eCfj8PKDtIxFyrMLt3Gg0/RpSP+ryPPzYbX8zkPXj6/w1Cin9eoi+cTu2UhmPoEwA8vG3dVh
LvgjAoNIAK+tBwu0XE6QqGJ3PC1KceWDNbGN8NIeoqPVUWgl2beSX+HAUsVIos/+ibR2YVuUoeLZ
kxJ/xagONqt+4f5W7cWCW7ZBnNaCtWSPFv7RBs8FKzNMa5W5soyRqczRctWFRH0YaBnHjW9ozxVH
aF/klPwC16udGXF85IMNf9dkc69U/Gtj/5O88n/pSHWsdCCSOw1Wu/fPRT3cbzR0oKWtvA6Gdbh1
Bl4BcDnb/89jxp5K4fQ2CxmMNxcmJG7cQpzssil3UVp20KDxCTUu7kbsNgE2HozWIPI0yMHUFwbW
ELa1WnKe3ylKiglFZvVs+yzqncHRnUzJEjQ5LM5f7vDB2pZlclTZEs3uBc2Vit611DrzkYam4G5R
wH9Ulsx/aInKd82hjdRfcIJGKCc4zxaknUTdeEgcRsK/MKTMtc7Oj7R576aXBSj/YkZQ/RpzX159
rgbd1ZZH0DmDUUHwrAibLh4HtZx9bpZVyb6CnqQYv7vH192NHtJmA8dVd7TCyVj2JIt1297vW+tz
/hfkG2zzwLDmCzBEYuLc8WApkEyhfekl1ZtFrNyktJ5MiRVN7U8GLJREftUEfkdahuOyP7Umc2KE
gf52YenNxzvTAj/iQ8W19clsQuQNH3nfvuLx+iibvlDYHrz2uYc5fZwB9BDqtFjlFI7odiC08WE0
r4Ixi/BRrGN9ylJgUEDyV7+vFYygYYxsNzgc3y+am8g32AoWgbwOdXyy+hS78VKQaVVcriub8S9K
FXhd8Tj0BiHu1p4XspbiRODHBtwLmLbOCbSdYIoLE2F4HIzDaM4GIn2JeBU+r3iG39QDyrB1I7oY
amiECZ3R10L6qDcs8W4NktvRHY0Ft8+euKNa+e0a2cOJj/yuydhn6p686NF8Mk7cJe5NS5Sxu99R
hFY4uyIx363KwpZ8kIBUszZBpQ8qb9zYskfdv62ZmLSNUg4hl0IlZXtIcxz5dbybFU8glRYUHFl5
ICbSdf6y4B1GuOrgv4MLKJGFUE09nWRDK0quhLunfvDdgJkuLTMw7oa9MuXurPXxpJXytZnFYxow
ZvGz6oWYKELItAtWxMQZuTKw1ORnhDzrPWO1Gs5JiC/oFdI+Ts7CP3yruzlQ5OrJsWw8U+6qlf1Z
clJRmntJwOdbNpBtH79A+NJZKqwe66pzHRqAYjoPI0iVpEYg8LdJakx+vm40DcRUdfbykwQya6HW
4SkwxDQ0zjLn9hKPVwydiORN149FYUTR4GrN+pVY8m9Hgv5Eb8thwLbcg1mJdwtRjbe0f9rG1UI6
KjWx2ZVwscED4kd3nYqIhZT7oP7uk/1PVpLqulhUbITS0PmgiU9U7wjv+BsEJDOzfkAJxdFBuhty
9JmkiSIRt6delmG3LFe499JxY4WVwOOm4RtScyMpfocWbwyoiM9Q4jiThtjil72avm4jM+pK3uCY
CM3kGjHNUbijiMZgMTHkSI3y/l/8CcWy3Ros5I3VuG1+VuUt8J6BXJQXJ7POmHe7iuPVo4KmFs3f
My8qUqmqnV/q9/gyg5uVgay+XuKHmdd0jA9Bx3rU458lqTN7H3z52VtvJlK9Dn+RX53HHoKfA0bW
Az6lpgEnYYWYq1gKqlM818/Xx+PnAjmVaoNqIYrv1DhJh7v4Rss05dG4kSJOjZdpeb1cr1IJDV2e
AivMqsHE8Xei4+UBpApBUbCDbhVoEnIdF5cGJCdmPweW1mnxE+9InRuPlORJYRx7Xm6k9cxX0Q4z
cCXLJPEF3QKmotBxtv5yv7ud3M+o7xb57bxUHQZSmsJx8VxWK3xuD2PXgGvNlpbHapXsYXpTPyy6
d2DilymlLEjkVKMbDhAVqHuVPqsQi+gu2KOlOeCAc7do7n4WhM6NOwBTkSI3kkiG9ukREllohd1y
9F0KeVYTqh0uyeaW8GZTXSPTdr6c7oi+Pu4v36bSlkigMd+bHvZ8hg3/0g1kj8JmoeKnnGw5QHUZ
iXTYipTghOCE1t6Vz+qnNraGI6CMWZZ/9ui82Im5ISY8LOUMNT+ZYatm+fNI08QJ70pEvXpRFNg/
sI0Un5kz+ST+qtt00jiGnzpTHn53XB+JGg17RCIiWQFdFlHYh2o61/NcI9nyfHGeqH6kkvKCcK9w
eQ0Ran2xXO6sPoGbcjCJi+Fr+CAKRxfpC6gBEc4M1XYFhHb72XxGgloPIexpogtRao1fGmi5fPg4
3R7S9Rge0X1/LquuliC8pFXjtxaqsLfJEzz2HHFN8MB/pinteYevVVbg7Mg6H+Bs8gLMXLV+aVCS
fSExSfvIm0EkCIl6RnTAWVVMdVJE+oAy1pgXZXADtmOPXOVAXjtL02ppy9YOBuHxtQMnmpweX6/D
vpYZblzgcPhcuUm3DbnJBvxpbshwaOyNb2P+2JinOoMyMTeQw8dWBzB9pcNSX9vIDM1jIIbB6Rc0
stVU57hcqe5CD7yUFrIeR1jumi/o90HrfijqzhmXmeR67Ows493O+jP7jl+ac+7zwZeH3WOXa2/T
qBxhbVu1PqdXF2fgNnURvNKvTvP3bm4xmMEWTMefMFiO3lWNV7lJPHlP0hMNaCAWreYYUqC/2piN
iaiLf9KrudDtOJDqIbbKhP3Zdq67Ti3e2hqopcZUDOHun/UPwX7R5MxFP05xs8MfXom8x5EyAHwZ
mIyvpQQzW8J3Br6AaTvQT3qFEmN+5LYG7wizBfverxvHX5bnFAa2a2sXdiv63fKDuclTo536ocYN
0VfDJsaPdFW7hcnOVZITJnL/GUH+RLUYBOHVuIOkXpF1ZTSZf2noYvvvFOHbiY7ULrUPn8PhOl6L
l+pnmGigTQOOFGMxsWpmGfJwUhUZ1gnMUVi2eNomzWjuD6l5Kra7Y8c8I3b6gaNMw/TbnXFvkK2i
VgTPl0Sw8GEs+L2x5r3qyZgG2Ic3nCP0xRbz8VLmY9ChiB5ioD8C6BnsaEr/YCMizT3QxsQqIqXK
tj5ACeR5D/FI/KIouSq1hzOBF4gGcqnKdXT5x6P5lVbH1o78K9VBJdzl9La/E4b549AYbqHwsrPW
u9ocS9YVACwlp2yoXyF0KpP1RBdeChu/Szh/ZfFi40xoPJ2dhYa65b2sArJxxHAqiuHJKkpO1S+f
ZjtRJ0DIsgfCnS0iFC1e3gF/lUgj4Ic4S3xkHO1t4aD7I9uHJg7s/KT3/zBJ0tkgTDCjjnOAv8wB
4n2Ncc5he/cjrnB+1f9BWm1S5Kv+UYZvi6wEGNodCM88SUw6sdvnZSEjZ7F8CUjeITCc6ewqdpne
uVVjxNyJKXf+2+3d7pTikisFwlWpyTbVE0MzJjqxe2pMedfu8w7SjOHR4jONx8Qj+7S98uhezoJs
TO21nuJXaHqIBEasKxFCYW3TpaE78uEl6wn6me8FI7bvvXXFY6z4eH5s8NhL3IGocxKzPyq6qs4N
cj6Y+G2N71klPM2sEa9qxyl8JryZTfLYETn6JcuZFDXkn2oajWO3X2lQJhyXcFiz+ZUpCGDT3sVX
CTe1qlexe4zSCCkWctOfrOTZ8Fibzd/aJuuuN5MUDr7lLXSa9luiApxhDl5vU31ZsZcUJzXTBrID
UiaticB/9FsgwOAs1RYAYRz+RJrgtaCTr8zJUhMsLhlKKIujrqVJtgVC+uR9uCrIPTA5ktgybo5A
jfI3JNIjjw4YudUm5F/PxZ7PMKb2/DTcndmFS3zD2n4nQ1xgH/wl0E4DxZRaAGIXfPKwIAqpO8dI
DC9A6iKXXAIkPuIE4oGlhMOHkKK2WJnipgZT1KGwe0A0hG33eJjUkM9fXA33myRrXLrPYzie4JYW
mbWUHYIhuRgjskY+J/A+OVooEM8Wl74KNh0VpPJWVp488U+OqioNKnn9gCBxDVv1XugnlGJi9UVB
cQpjNPMOsf/qpffvo1EOVvBDqp7Qpj32PtP70WpbGzJI/2DlOmoMDV65VP5MagLaNyKDQ1F4bptO
4cCmodE3HgJnvgyR5UoLWL6D5HZFhshcZAv5L3J5j8LvT7vgHYTnzpV9bO/Epl9fDCkY3wNbfzjZ
CoWEcZ9xC2DU30mKWIvznDxB7bw1ofZZpZ/C3eXPJGvvJ2m3V9uds0qdV8b0HqORB5SooWnePx2H
4UOCXjuln3nQFIWzvXEh81juC3nFv46i/qSPLhwPwPmHcSpdfdRl/cynmsPoDPVb53B6fUfzcRLz
3cJOdxkvnMaUIcbt3cNjKVG0+tZwHLSBRrTt9K6nwEXFWqNa30lrT8Z1a8d3HB3PDtuoVErkF1c3
CRfjWUXNgUZn+pg/RJg6+/fOCyws6M+VIV4Ig6jiNoAOvinr4oFdvRQJ0IYGAs6IIraVTte6nfY2
wlu9BJTKhRC2v6gh7RZs2gqGwhPv5l6yoXQET2knsa3y0NsYlMrVbG0ta1FR5uPgpL3ugkep6YKv
tvg3JEDMHbbk/MGR41Dr0DrOIk1GKxr7mxiXbpFxjKJje9np8zBm4ovTDctsIqSe0esy4RbF6Wk2
DpyekeshJBxch6TKkfhatnXxHo14pWOThRbLvnOXmbSSWz3eIQ8tZY63ymoGA21EGypd7etXxjNd
ufcipMkjv+6gBd3J83oUSOPQiygAKOC/BSLIlKowgF6/IiMjtuJ8gfhvABu+5slRY4/gkkyXsGqd
k6WaNhHW+H9Ewo6PG+IZv1A533zfLdp2n0+5xSgW+sgwodLfx7E6oMeqcwiXjKYFWNchhq6Xr0Da
VqYsV6wLDIHDmz9aMk9DY9T2euQpE9KC0FoNgEl7YOCWFUveLjbXW10ahELpJbNqexgSXVF3JTej
FqYhzp3+txl+nBjwS7rs+czTzfhGw1VWUqDi4FCX9MtsfDG7oljk8jf2yTxaCNjed8KOWkxlpuju
RSQEQrKiCYgioZ/rjGu8P1qgJIIA2dUu0Kx4wcHRgbdzRP23Bvv1HMqZ8YXZ3El5OEdUUm+kElvK
1MYuMrD2oOtRFLoDD7lndQI+Qa70Rt1DwAJUJW16Y39qSbeLA/+JGzD08rcKbf4Zkqk4XmCeXvj6
XMFxZ3+MyF4NM0fTc95ThNDK0H3ueQoLKUpe8yzsepAo2+a+KkuO3QXFfeNdtBndpTw3EN4oE68H
MdlAvaQYBuUPFYjCE7zvQED43pn+6YsHHVc3mJN6EpxSkiYrN75ukLIrtywgoM3VR1Hh3gnoxW02
3NBeuBswWDSJd0Qfg+1Gwx/bhZQk1fm7csQtXe217EhXpfbZS0szGaUz6vSZ9rGnBLGl7sSkyq8x
53bkqaTd+6kFiGZnId87cc2FQIx8gK4HSUVT7OKkEtb5zYsKczX2oTuDBPOk/SYrs+P20iZmdjtW
/cl80grokWkYhUjY3Zy+zyqkUtbZpkHJSMxizZRH83d9jnULlIOSmouSH9dGjfiC7bZDjQ4l08xx
H5vLI/+20HpciJBcR7WeX3JNQSXmbPQk73X0YEw+TWnFJClVWAlRFQuctJt3j0mmPMfBt8h0CqWY
38kZf0Ied5rkh7jkiQFij6YeCCCFqsIiyeV23JfUrTGhvm01BH4BU77JFBpnpd1aymYNVL6puIE4
dLBAcmSjpaBOvuseb28fmnpEFq1m8v54kOTzHh2r0/F5KNhJPgRwsvP2/AShmmX0tMI5gtYHGwkI
P4sXbqmxL9lVlAAt6CYxY2NwAg/9R+mMGJZ4d7Vyx9Nf17tny5G2hP2DNNCOm6jP0/C0CGqMmTZa
oj5NcW4ajmN9H59uAy+U0lbei7Kgnwyjjc2RijZXjooGSnr/CHMG9VbGLpG7ltOamtUmBDEtYwoZ
nr2SGI43RlutcbqEXGhZR/pd1v0RHFZK8MJU/+W7ktbcbzjdRNp5C6xIDNSoSxCdyGHy5q+IKxL0
2wKNppm9yeEvt7JmZmDj2vrBe7MlRbK8zsScVJQqgdodJUO6E8pSP5557vt5hOeLF+o6hNgde1zZ
L6faRa+06Cy+2YAEKWqB9JAMlBA3Sv8NUZhsW/Zt3HE6YGGP4rPwRVIrQPuECHk8UIAy7VbpKrEj
B5/c9vlfQreLcHuSPwHupYZnn0hZcRk69lcecg1pBmSeJRDg0q27B8An+dLtXZWN3ZSODDYnJ5B9
aPEW+TmLerF6239R1VdViBKMkeG6VvQL12dOwpc4FxGE0RLx2GTf3XOKFSs5+bEoUuJKNOZzp5Xl
R6PWJxV/lPFc9tq2UGRIjeuLbOjBzUTBm2gAx6MeoiW83lxSocoWMnzT1KQLhb9V7sAJP+wwxHCc
uBrxfwOtcMt9K4XfAK0Ia6RbQCXgVgiuXKGRxcgBMsvWyiErY6+DX+2VhEf9um8CoVSqhODr/fsA
CicgmaYhY1rCJptSrt3uFZnewb+4Ea0DztdNWLQlwF2h6+ayhKRqSI0xEENcwIJ+yqhPzht1OL/H
27490U1WE64fsXKSLnn/otIqsfGHBV9dqInHA3O6LGgbhe9T+FckpAy8+d314ZjT+WnZ8tBJFDCr
0zUOOFNEhhbw+6A65li82iEd/HfhPEgnUc6+F6uq02wX0bR5rh6XC16ui0vtSVJlFM6V4TQNXiHP
Dcw05Gl51pe34qAwGB4KXZV4dupRyskqKgjfMD5KbnrXNBvB73zv5hNJRbzS174bQ8XLjS3Di3b2
9V2YoGSLsSf3Doy8YeB8E1bnqGbBOBqjIPu0w3RA4IW6G7Q9VZRBUOVTfoILgQ5QgIdep6hJ0XdI
Q85Dnny1cM5ipX4535cofH9euoEYPGjK9pNYFFQCPNuqwqSg9wdsO9ymgmngQ/fyidl4mmQ+OA3g
yyJBJk7QwOwGFd3dTDHkyEbsaH2uY0RifI9s7dENYfMMtNvlPKwzFNLI89pmeHkxzeVCgIk5GOdy
G0MvXqtp+ZBu0FfwmxmQHJgcBjg35GHlq8j4w/kTn6CJQhxnEspEVzvXXPn6my5ivKwo2g6gmUwM
mQ4dhQB5QcQHE9w7UOFcmDppSm2u2LGaIoANkENaLnvBfbqJEYvOeF5u9JA/3gAa27zqBSOIFLPR
c2+ce4AlwmzYW1THkK0qQz6cXnAwdhfdOHkSQMqCR3HiznIywztORqS+O/ieFxBKzw6RAXtNTNrz
5OC+aftBJi31n3T7YDKxVgBoWh6uzax3s/5Ve9PhWaVlmqW6yVRWY6kntewgHz+OpbA3FYOfPsYO
cvHEPh2tOcO3RLmDSh3sAz6zog7mVV4vZuhrqXcIoq9iLXFHZquXEAaDzz723kes1Eq2mPnnj9jc
RzH1VxghV5CxithzV26Sjcgu9nK3HlQcPYHd2jRFuu8TG5InU49uVYCYDEPQGRqJJK+U0Kr0jw3S
RYI05NO9/CuANf/FgJoru+N0cLwrOuapP6eVO2qMRsGziYHkZWvkgjwUJ/oMi7OAN+vx02EeX/qv
+y50cdrxQPcQbD1y9ZYxDIfAZ7wyGOi6eD44TsHCdHKIy9aWJO+GdkP5Phlk/ko69B9lg8Yx1YeD
W5Sz8AKXvmMLowPbiTN5bV3B1ctYwobnyyDg2fm35eBEv50exRWuT/WIL1noDrF/rILtqcckh/rk
QNFXn2b3x/HXBRM5Z/4F00w2jU0qYvTE9Pjbbk8O3Mnc/5JTNrcsGxfaXj2dfVTo8dszY1v0DQIA
lcF7QVeLQAqIiY6HDEMFjkN3WlhPp/V77rZmzPwfkBOqOnJU0nH4wzGTg92N54WWZnjEuPPIKxY/
9gtTFXR+Mt0OVW1f7yrHB1wAi9ny40I7Th3588BJPzvqPoabg8L5SLsU94NHg1aIyO1hq1axsuSp
YImcSs9tT5SmMT2O00OJKe5DPxk3QjI8cj3tBp8NGRpCnewXE+73sjzSUpXIeYNywEAnDvUB2qJU
oB7hf45YnCpM9NErX7b6aj+iuVVh9o6Y0CmZrciq0JMtsIWrebPIIEd2a0b89KW/R9hbNWOt5zhx
kmj6tUx+RWzlNQpFDlOfxBC83UskaiIQMatcIBaCOeTd0nl84uMxdIT82xE4i8OEzzroPzXR46h0
AdhCq+UJjlLfdJy5je70I5knfr+7pB4MPOQLHKHplwHbxcgvbxOf+yVjo+XI9ohs7eGjgymUocip
iE4d4qQk0xKdI961n+WXCZaTD63uegfhDjO9DiB21EuNrn8dPp2J1iKNvkPzy3Le7qQujF/Lk1Xz
WrFwudGfeHFvqoZk6KANC2YAsVtNgVNlAaoR8j8jSCJ+LBcX7659z+/mmryJ9mt56GZ0vx9PCvwR
z28j0vwigK/mKKY6FUblJbVObY+hQen9xVWB99z7rFqSug+8VyTZXY4xw3s10fW5dyOOtvkwlaRd
7GaGXepRbEZY//u/ltileo9OBFFMmmsBTeggMmav3rtxzJavMVq40l30yDuJZEhP4+nI53FCySqH
yPRFec05qvZxuCSVtWP6FoMhAHRWMydp7uDZaIqpxTVA3V5VMvGCx+xzKTY84nJEAOeDQKnJSbDt
ng0yGzQxGxMPNUUf0NxfXMoh7LVHo3c8aagon4rHv2wtvtoKt6D8WddidwL5N+Uo3xj/SCvSQzMV
FWpceQF8/5h3eURxuqF+VPLLebHZOjBitoUTvodNyNzXgrvcQjehbSdJERKBM0qtVipSrwxQbu3+
Or2Vwii2UiUcRPQTFXkHQGbT3KgQq1SkEgQ9vbo0w6f6x5MoZkcUuEuHbhaa5ncCReaEH8bEEh4R
Y2wQbLZrtKQ/bn6GH0//E4wgMJdOyzcFbwnac/BbEG/KCW7IE2m5qG4HJb8rYx0vnMwIuT3nf45j
rGYSm7gStBq57YaMhBObnAaBNINL06RfkWNYzPgvr2WSroglYjPNiDkq34F+a1P3HPY67HsUrIHL
zZkd6vEbR2BnCufr7r5OwcKLneEBQ4Tq9pCLlK3AvdYnuE/ePBOEFhuyIrNaTSEtMw8nNe1rIB0u
KeDuVlp4wvQN6EgzYRw4CgLPXhStbq1NizyK5SjCXmuLBH1C6NWWmRrd+CQ4YHBwEB4djiFkbfOH
B673JtPzilOdo1iVFWj3ub72ABGs7Znex6uc2Epu00f/7mvtI6DGeIrWOQSEPOb+/esJHTXZpy+B
OXuAo1T5Laf/C2aBjbescy3aPbU0pw484x/IAyhOh6PM7r821j15h5uzuCAvaWaHfDLksHnHS+9M
On/TeTkBm55/x1xJL98r69OpE0jCwtWYCgkpFEtvAuVt69nevuP4hqs60Gzcf52CsN/bnUMWMqTJ
qXtBNfvm6UY+X1NcFS7r6tRz/xvKh2q1nLCu3rWRpbH3VyoNgsUqWZyO2MtOnWEt4UN34Qqj41ue
7BqfA4anAoDpOnPUwLnDG/4oXQUPWkcpAbvZea3q4JkOcNcFOsF9GJ5CjOckQ0T534UQU/NilhX0
UjF8Q7prDUzOO0nCegU0/uVfag//B9J0ue3X4FkR+lE8N7kJfBPDA0R/VQ25n5NZvQ26LSbeIs2b
moGaKJwbqUZjJ8FzCUidIvz/cX2fxJHJUOc33GnH8BQzx+ev7gozmHnFmEk8kxuzFnPhxerv1nXu
snq1+DBnWblXoEzFpd21nr2Rfyi1ZXJf3mCj8+eQZnrmqfgApS3UfASxohvn/OuWJbcbi6Pfmy0s
Wds+ABVKgJRorrA87/GpoPN8OOuiuzmQ940HHM+X3BNgJbvwqEFSHSRFRD02O61lQiWomSN4nymK
5tDtmFQwDfO8qTbU687Jbh500Q6hefozGphoxbxt+P1YnFf0tDGH6YsUqBdBLQ3LGJOdoK6BNuJL
/v6Ppr21zM8NF0RmnD0Lt1UV6u1GCDzoN4+g6aJ2hN7OvUppGfwPRo1Gyj1I3ikI+Y7upDJLsZdh
NRAkxOOHLUk4N1k7NQpX65VuES96Gpr2gBvwEp24qg/4IJ5LSp7qNvOYBiPyMFgf1VPcVeIQ40NR
8ZacIjHW6n3qjvKXhHeglztmTJ4GLxBxRthEPr1bzei27/xYy/Rom57pJ/A/9afIihVr9b3Ma9Mf
moKxEhbGvOni2EpFj2a83elI6iHXSHrcu9Wfb+1n408MufApDWRsamhGMiobt8GTG4O+Uc51tQ/e
RG+fFILlS0cSbpQWTbSc9xZ1J+iFVV8cgR7umVxtFAdLpdYMGZbxVKKRJK0QA6cTaxL8FvV+cLvr
7F5dU2NOF5yp2at2mssx3U19Gj9iFFz0lNNGThrkr6FEmRsvaG1NBpk4qA2mYJrQ5O8e0MoKN9v4
7fwj9Xta0RfzgNb+lzIm1WDMynfA8SPjkJA2/sfvhY8rTaZlzxN0Lh4LjqYlxpJ7oeiOTD+iKhyN
f28w0g3GemxMI/5ZaAOCBb5Z3aalsGPclz888QZESk9ov+OYOzGeCwFvH4/gxXKkMOZesegEHCXX
G9cKn825Kdp8NPQ6AF0Bu6NlaNPI8zgRuKw/k+heTtm0HJCjw0fgHHNr28RdqcEewbPbPaV9X2cK
4Zgso0mfiGlib2zZf4GzmWlNeKbN69C0YEC3u0uYSP0rXqid/15twTqr0/FolTDhFp4e15UzArG9
UwwsD2lupcjZjENlOVbkktykIFgqxJWHvhjjCAaDh1sqHuxGMzXQnQgcbMumOK9c46YERK+Vv5xC
+/qAvciU6oRW80kD/buieNgzLizgMWpEKO4nsvKuYUS9WgG4gHsan8j85EjQubqgVXJCxgtxz28d
KRdBBNqTRFsgS2KiLfk2/SZ5l8+Gh52Ask2C0mDF2K2Zz7KyALa2HhfB4KsXnSM8UliKtuvolMwe
tPP2kYXeCvEnY5Z1JHAqQ1UN+TnvzZFoiWgL0rjZk+ZPFg1Uq+uaYTbQ2VHYtDUXX8Oxc1vaSfe5
/Gd7b5awfvCiHzOYewTJvQccesXHxqGfouKBuVwwd+DbjPgbuhhpwHzeBrqCFRiF941cYIOiQg01
Oa3mK30Ru+l2UntDaZTlMCLuN3vZI1h1Qt8UkmUKQP2Ge1KHoSZuCg8Q3cidUMRAzhCEPMQ/oH9F
xbzNgzQC24X6AP0KSm20OFyBI5A0fVsaLZSStYljXd8Lugt3odsO7sJWWoZ0N3nsCinxOHaLSq5n
hBFWjW6SWIrh2sVauYK5NJT5WvvbNuMi1HCjxSJm2+VyFD4kMjg76ocX61KDGD8fZTUE/LHldeG1
ma7r+h+6JQuhwl2DuXaAxqcK4VzrPT/Js6yrUTfG/gaoZ4wVuw0SZ4wY5NmwKaNBjiIZh7rY6Oe4
Fhx7rUAmL/S5YgmeIV+XOX9NNWjVuY5uUracMTFYaMw2s5aOOmOExHKk4ZZXbiQvCkQGauzbp3mH
MSqXSH/zHTLnAL6hrBGV8G0WnR78HKl0nCiaRanzO3Fvi1mfdXIjQnjmKKaAmJnjP/kQrtMQFxOP
cZ2ttjD9E78OgG0TwTNJI9wSMOzkrHNoynhh+lvNbOf7R1a3Y+lxf+gJuystlZKTZid7of2I4r1k
xx3G1ihU67i0co08WNM1h2I28FtU2BviU5VVb/uqJEgiA5R/9kPQqIpHG3PUkjJOzoahaAC/Q5E6
oauHXFbRnqBWi9NtsI8tGRczpfPssyhFEBXMY793wSGOXzId3cEtfV9D5ssEE5enEJVO75ti3hpX
aSh1fqbE73b/+g7nfd1ao0Xd/1hpHz/c2zCTNHE3fhURCvV+SeGuZ8zLwzzWwOX/1ZMhRU3NYSZw
BAhIB+SZLLGCjr2vcRyFv+Kc5UZVNcAMgasImCYU8wRcYu0GQ7wqv8cdZ/PruNjGQ+zFCOY5nsd6
uEeagnrKGMX94kPFeR23DgFaaXJ6z4alFv8w9YnsXW6e5HfLmuXk6WGAC4j25svfRH8rhDPCdmth
6fcU9oJ++OdPjvaTYsvExLGnUNbatV/VaLhSMU+1stdJndZMvahPjjmiPyEockXXvLjF8YciqWAI
19d/P+w1S4P3z9NTPlxCCspqRXLesNFjI2JHg5Pp9y4a6c2+fuTUaoGL17zvQtVALGx9F4KSlmK+
8q5Xm6cjEmg3hy5QZ3HmMZN3avHBoxhuNboutbFRHecWVhREWoCjtwCk2hUe97rrd9RO5jiUG9rf
xEEk0ISBCdnR6Z4ph0W8IzBVR4DGfrHWQRFh5h2e7+aqa/TRlxVgkkyoEOugv/RKTrLKLq9Bqp6i
EdjvuqDL3r9/D6C5e1B6VH9Tyrk5gS18J0b+BsuIdPx98M2mBBwNvZVFPSyTxKfyqFVUuxU3sGGz
lEmtaER12UTxP0tShJyzZ0akLE9oO0KW+bJbx2DP3pufs0JkQ5qZzhoHMAObv+liII0et86fVRGS
PpCyRailsFsJx/gSdTqZ5+/vFGNBoRIZjPlO6bd5Sh0KZfoOsExAeyg+Cg6K4/qO+Z+RM9aKxJSo
m4gwqtxSrLumFn1tARYo49AIVQqayLGrxiDwsVU3XHfc4IbVqtj02YSJf+l94J68IS3NBHdTaWKH
BOpnosFb9p1GgH3T4TAqRFQRTCVhlqMuxuimYjX6a5Ql9PiFciYRd3vV1ZHmTeckBtsJifl6tp43
aUsXjwHyH62YORuhrO6HBjIdvatjEv8eyxeF6XjHl6p8mBQqxg7BMeB1dmKCRh8c0sE02+R406U6
bcSsneHLF7i+j5whMhEEsGJy8FgaIKg8jpzo5JWLQzq77j1lx04PBonWgKlEQBASUF6tgdOBHuXY
BjQg3QQKLyyKdgYOc6yvyH+Ti0VGJ47SZ3WPTkd5eSMGAoynkmgKArYgsW/f4lQM8YDjEmaSaJqS
Tw4h+GMDevvi74D+uPVXh8haAXGD7wZnMAO7MrW7G6FusKYzCjCJb9D7tr/sj5F3zr/IhpTEp4bN
oRfwFJeRttEdJbjm7O9SGKJVActM4fZipbu1dzt/V5U5prv4zydTEYQ0qJAZSaEsXswmYIPksz6B
Ngkn2FPsPbj4SUAna7czgbg6yJuqAHEy79mPtUaUC8jtTzW8UjXfXoouu28cTLhFOPQlphZ4cSpY
5DDQYObc3TLgpn2rhIO8/ptFon3QXLPNw0be3iYndeqhdL0s0xy6TZGJMSfEAmqpb7UvydXj8uLu
CaIX9pmqIypDQ56IOIE0NKS4dAqSZ2zJw+VHCg3oDlBuOB9+dmOHTIuLGzYULXb+nOBz0a0CrSyu
goHuaq4wmZ7dqeDndEkdeaxeozhlEEPbNqxylasP9o8XgoZBqDj6TlBRIUqb9qyUcWUsG8f027qB
oPaj6MJdaYtC7B7Wuz9+V0+0021Xu092Y/+rpe0m5oJlEm3Dt3mma6CA+4QhwiU8J1BxfGLUbGxy
8AaHQtcS7HT/BKFkoHceIXmUea9NBu1optRzECWzdqeC7MG+qkQMvfyUhp0VgbjkhYiJtD8otTkj
WnaoYMgoq+6ObHbfn7hiCmjUCN/9sYHFogMLeMXa8KeOQsWFkOjDveg7jQGpiAE/PHwRVXnM+PSZ
Gsy28lhY1awE/UU6CW8vqxDCCChtOzM0dqxGYyUgqZS5tCWvOk36Tqy89wdZ0XevD1Bf2jm6+OTA
1sGE4NEXi5fsk/Oc2t8pr9YL7ZolPYucqKnuSTaMVrpX3JsWDMYpdRPGwkmsOJaNIl0DjOo+oyv1
nL22W/OpnI4n7w8F/66atP9u5dmEXjYIZZDylYj5SA8fynIXiOAvbiZYrnokjFG3NIFxJhon7eQs
/LBEOLFAilJm8s6e5Ie8KuTlUBmqZnmCRignbEtPBTnJhvVh9qtxxIXBNbtBbNau6dCIWuazLjMF
YrJHXnZQh84DVACZmwNqqwSYGBFqQnonzNyknzqqIwUYTV0125vTMwIBHs5p969ZlL86F6S6ygH4
MJIKwcH6GX9v66vHaxLCw732oaHJgBZyrI8r2q3Adk51slC9vqIZ5xuFZLiC+dPrHwjW1aUM5FXa
xTAjwdrzgTtDlx3r7P7Yvu8dqK8V33Z12LM2RLHHdgDAiISDPn56D7UtHxugsoqXzkmNtRiNsIA9
6wF881wSsYYjsV5tu9owAkTqIUP8vDT5Y1Yo51Aj8u5p/NEZtQz9as5t9CwQ4RAQj4h2V5Vci0LU
8DAor62s0yyH1BM6Jd9gJk0C7kI/ov4RwMDVvMcOtqNG/Z06/WHaPYqaa4lY+X6Vr6ZNxVhU1Cba
JnDIi3H45I2sX/VFNQVME/wtU0gAxyWC8OVmYEN/GtoyOMh/Lg1JPhnOAA+TwA9xR8QvvOWbOBYK
1kGLo1NoHNK4iupHTM76FOkxj+iBBg7bDjs7pxYFT0OCC9RGHV1F8aXp+MdZLPrs8yFNxesotvDA
BxKsGPOsC1uxfBwbbnM0kOEAcIauhPbce4PMDjTNanQ+xPnEFJ6qSYxkNKC75a7/ETPNC2H5biNm
0cI70BsCfjktAvVrLIbFVVILNRUZ7FlTYhBje/aZr3pSH+Kbv736YhlbDLuV+92svZB6Cp23E7+1
OX6OWxYuf0H/hvASp4L8J116i3XXX6rMc5erWYQGTDyjVwqbClRhVaQlfbPQEgjid2bPsxgicIbp
NjFwVWJJV1lBI+yuMcRWOI3A3iQKOvm16W1v7jhNw8eUk0rgPf9oB3RyCTId6+0BKL8b003NzHNA
2+0AaoBbFvjTLxNPOXYqZmnnvGLcTd9cVU2XkAc6tqPBDZWUdQthPd6i+aYg56p1vuLQB6JR7QSJ
j7sNbDph/otTgPCZSr0LUC4vt5U6hOU6YEofzBehy9KjfbOgEc++JVbJgoGIFAB15O8BP1JY0+za
1UCfa3hUK/ZhlZK6H41NEDKxPXLDzWp0wKb4CUoj7ulX2z3C+WxBgFsBtjv7pTs685V5SvmorKpe
ODzr3O9hXxhNsP5SXSQmPe/dOyf29UlcA1yJrJIyeRFqlK1k2EfEHkPMoXNIrplMqaMA16jdyWDI
C7ibFVBTbTYVa6CqGMR34G3G6lh9U4X8whgV4qQRQUmvb1Al+54Iqr0obVkY9LHrw9F9PD2iHKE2
JCWJJ0etP66BBHCU+D079EAWEl6SB3wRkpeEbv4ub2zR9Duij95G7etr57k2Ml1ckcl6g28fKagy
bIwi4Jkd14jqd7DBN2hWAvFPkw77RFhkjurAADq8zXnuNOjrmjnI9Vh+OnbFdC1WpXjLin058cfk
90b+KQMvXyhYBRBztXZqF00fE1NBoW6bFceMeCWUGyWJhDCxy1pYkAJCOan8pRxeM6K88f3JGpyx
xqjQhyQSDQhU9c4QkUlUsqZBhnyfoZSjI6B4ZWFcz2TjabXg0pqDGEKLaRALzGfCZe4elVGUJpl5
FIQb8LtBFb05/9NcO+j/Mz38UEuit5XiFJaYUu0T98P8+6ZCAVN7GapLGvOKBUlRKGbCKLGeJU+A
ArKk576Uvw+oY0dQRIRirBkAfJ0GxMOaopkRNU8wmaCp2I1T7NyFUpW/k7vrCdggmlt4+RhhQRMt
imHrTbAYLC/g1r2QPJa7qlMFSK9A4yKwhPQ9JyFtaHGM5J0fMuj7a5rcujoZm2E6GbiXxuZ25foz
VfQs21Bwsorc0AV3Tr0myaiN5yw/cl/MMwBKQeGVsJbsO9umyo5rG6MxKx1J/0u7+e80IPWN4Zlo
h7YS3lmljsygvQhs3UFraXAouuycIrsM0EQtz3y4AHPDN9f/IzQG9ftJ3l6U1OrXdxxMC6VwrMp7
34OUI4jnFsqL8GqyZuPUmKXl0M4i9I1PJ34hdaJTKq/LB3yB02S/uBAODV0dkq08DmzOMIyLCtI1
jzO0bQ8FAaF7lTKXWZucwwXnFyG3lOOEh8hBJ9tHyr8PS1TjiLu63XdjHo6f1dsKHvlgOLO8Fkei
0VbM5cmU1s+4WAG17EP1T7TpsCyKlxHl2gBzlLiL+Ql0dqzzFEvNMqorrk/DwhCY4VZ1SMuu/haR
yPM6EPRCuChMp2Nz6LbKXd9uS5pn8ZHks+/2o4hfPVgfXpIXkPsiAm6xdl6SKyMD7V+Fgwz6JGDq
dh7H97I/tshX6bM6a4VEPqM7geWtcjdakZfRMxCgfdNSWWDjYo0lhsraWqeCT6f/TQnRTFG0B/NM
r53eR2wR0c42+4yc8sV901XzvKwNlsFJTjhy8HIWzO9Sma/KSO3qNxNrg3cA6oemP6rwwBDwmR4D
r7NmW6z3N/dtMoV8R+3oyFDShZ/YS7guEJL7e+tF2SrSzKZM+Muy1A93ddQ6ARs6iaEytIovcfml
cA53xdTHvRHYwMga2AspuOgcotNCpGub9G+jb43k1BBhFhKm2l6/NOWE4IXdV262P+shmq2T0ryQ
oNubJka8x+VPXzyUf8ZEoUW+IqkXKh+LaUf1WcIQPq/Z8AGZ2CAXOhqXde0pEU8x7pfmoz9BY5hG
5C9SHAdl6vuUmwJc1PIQ3EopkEbJt/Uh9twb/4iq2XJZC9r+ePgTVbW4N+63vhRtuRWaOrI3a2me
mQ0FN9F+Dub1uRGTBMScTlvOAUOZBxTuPIaExpZ2QF1I6CtL+y6Sdn/QtsBLQf06Azq4G6ANeY0Q
qswcxsbESrLgZVKJg7NISJnktFvNOz+bPSsKcT2yS14hUTERAnafQmFbQs/3N4UgubgtirPahpuz
XusFF+kvqsZYlLnK26gGlTNo8GKntKXq/Cou9TBYzGltu84xWCsYgvqvItSJnxvTm8SVMq2sfQ9S
8URz9LTgZEqs/8snRRGYrFFsbGStd7mLRWGrImJu4ElF7OW3iuOK8dTFyIaMQZkfa79NG+1RS3+9
MexhIrNWlxF5zMc1IYmGvabg1N8IYvVZBnl1VmUfVoCPKi20TJPVBK85uofh8iZObfChpRsO4kFi
amNnH1PgbtSdcDPmK/sW65HPE4qyawzt7FNo2Fo8Egs7GzkcGUthU4ngSvFeIyTKQDr1brOWix/4
4KFZUzdxGZv0EGIJCSi1BZDIsly1iOPTxZE8fr1CBhdLRR5s/Kfqrvw06El3tr8JrlE0D5gzf9Sh
Zh+QfGAOeZQnaajVEz5tXd5dllAoguZfMSXlsNCFvpvodZVxoAvEKkvOkERRRLSuDe1zbo+vRCdX
EFPbUqJHvmVDedvrAxwFYu6IxrnfwTijLYkiHLhT8H4D5PNUOYYz8TWxYA58ACQZbXjOM0WuOOYM
qpIW1EwGnvbMKq6VH1gVEvKsDrjYaYqmJdEZZ0bk0/hLWRcpVAz34OTP1GN3WTGIpQmM5GYNOrIT
dWX75V46282jl+t4DBpJ2qJdtox6YrHmifFqjJR9QjC71N5AjKW02Xz2vJQDKIJJjbL40xC7kLr4
CIej50L0jw4K4S6+k7irlyWDXIU1a8OKMk2TSl++mU3vizyunQNqnXFFNXZ1W+H8lN3wIJbUwCkT
pZG0HtbtNR7dkvVL+I91PdQyLdfw5ogwxZWzJS4WiZEWqIGSHNTWvbwzFM6ZdtFqsYSIos2wAjvl
4CoqYcpq64ZQWkSFo6Cnfx7GoreNVwWvKR+KO30Sn/BleVfFm+x+mqk+ikmNjr3VZPkyz25AqX1v
r5GdGdvuaYevZd2dL9Xjvr4xmDmnEXhapAX8pQtAqTj00QkrHFvNACcxB4wglE2ky15ullWVPAgI
8C3VhkPFQBxG9ulqTtd/G4cYVvljTmQOP4qNFnfFSzremRASSj6zO4qoOwF+DUvTNg0KHZCtmdBZ
rHf8zuAEoXT29eodWbDhoA42EkCEJCKhhSkNkD7Ek8EUiQmePAzJckmh9ZwgK+hQZzKOSeDFIvQA
uVo8hkT/O3Frhg5xUc+zL6zfpibA14p/VGxYLZW3Ly5rUB5xZDT8KsO6fI+C4VZyGFW0Cn2Celun
UrcGbQJJph3lP6NNgefsafpotHo204h8gVRQW8e1ppz7E2RoIGmt+lvM8itSq79VVImLjfhTvhex
PLJcimVW7wdSncXbzLuyVV4QV+F2HqRchIrVJz66S+d+Wipf61lfIzxNCUUP10O+aMY6CREJu7fp
FzcQIt0Q/uJ0G1PKcme3P+036qvQHQIBgPALOxrFYf+s0/HUrzM8Wshvd2c8r0MIcnswujxlU+nw
JJpEthIBCEh4dXgMYzdsW5m+o2boOtXtu8q0K47xVd3qacAF7Pa0TE7TAVBmV0awsP3Tx7F1dUuX
mcIT4OVKnjUkJPqvZXZY/Eh0fzM3rODHoLvL6lF6LwdFt7hXxl2sesNfpBgx+8KJrBKZeFU11q0/
TNmHfVSdEY4sqo9xBo1MQdAi2S7QHswI+wDnHfzvAzqCfFvpek5bCHqPkS0dFu2gfN1Zxs1AmZLw
myfy9jGyjHAkFc6mCh2aQOYJtmcPyf+LFlLyOzISZY7HUUUnHEj4XchtmPq/5BMJpOROCt2ZGbPp
BqOMltqaaeevAuzdo+OsAQPb6ilAE67wCWV68ImORl/Are2NU0QHcczrY3whDc8yTQPJaz87Hzwg
3lQvmNsERW7eIRaeCPPEiQF06f1Hmfnn2oGu4QMNG5NpCHn4cBLPjxbxlIUaRY+z046W1O03ELcV
XtUQYP4aezDkmbMmtby4PoX/oKre6FOJWb6KFjO7nwhYeTnRVInJJL6eVxfb64SM4ToJcpGqC1QU
vGiv1JCDAxqvqCHd1CvJWVzno72w8qhkhiQbGzkkBMp0s1+Wd2ElBfBF258lhfagAUToitkGlv4O
IM7uqIhJy8HjfjkrYV1190tJUbTO/mGBPoreEQrpfdT0sYOorMjUY7rFm9rI5Zbra9od2OAOUxlo
YOQZjz1vVvaSw9vOwisD6df2XFzWc+UmPZ1rkMwBoEfjJxlrrwBUuXCNgeKHY5Lbf1AUh4WBS5ku
ONo9ylSvJ9HXish+fsewWz7oLn/sMmrbNd5bQ3p48QkqRRsijp+Z9fcGDRo4j7ndtyEFIBA6593X
nrAw2wvhef2m0DvUzOPaPQb2tor5jQGMYfD/mqYhlYkp5PC2+Z4BngJ15BaOH0uh0yLRfRNsgqL8
rIsOXPfoXg+zxm6NDn9Q7vP3zSog8pc0IUD0imBn74ClsyamnAPElIVl3qKkETFQDdC5MLTvdzFZ
QXXRO4ReucYa3b6fECXtG3d0qU//SmKJ6NvKwQtv35t0OYC0Yq89N5PVdVqIgUfeOSoMQkYcyMPa
a3mKCNYfuTn6ktIRmffE6GxkPCUgVYi/pjmTw0VdtTsEiDpY+TOALar9jWxnuqBA+Fpted89qGh/
eZAfELmFK7qcV4mWbpttBE5CnckoFxL09jlbHOeGO08vgInj1ssQkFOp1ccjgsL2ibF74lsgoiki
Tp/7J8VHIud/NisBav2E7EaN4IvXIMGmqXWh/KyietGCWV0M/LcUgHYH3V8VFsuOKy7ShhipUD45
ZkAGXq8xy2MR2J3H8kZQAWZR1umXHxAuxlFswyyC3Goz0b/b4cKYKUiragOV2E3I4rr2WkILGi75
lkzkCa4iL57qIZpK+uT9Mh10qXzyuXa3UpkX6Xm0V9UeCdJgjXJMkEAMuoDhu343InHylW1k7Z43
/mfFKHv6gNC/+0htPujmS/yztzYN1L4BElUKKNUeHzQ/WyhZoS/upCX+VsMVxlyTwydY2olh61Gf
uwh/uzivmhwB5C04rzmNeJ0cSEU3vsGLRZVlBR/kDoVzG5oWAWFIy7kUf3Y5muoWlHl3IeJ/dYq+
fz6XSY0o2e8n2mAg0mGI/0SkoMKjFNVvt5fbcNciB/lT/Y8TA8BOpXRxQFuPF3H+/BGZIwzfmKcE
FXccL9ZjpMTsefZaqx43zneZf4tfa/i+FZ4o+/2Qnla+lgJqTALOHTUaP1Lyb8x2XX/RcXE9nRx6
chEzVuuoTXkojq5lYLCd/hOBJVYvzNAWve2fEWS3SaRQlw0V4qbDNyCiOf9j1Nb5fzTqGEcWf6dr
Dx5BwH1qQF1pY5OkTW71u4GXDCAXcrzpQIsrrS0+1JsO2HJ/eMDeaLicthhfSXmDVA8f8fQTeT7a
HBjujyY9AF91hocWMJjwjhQN6o6mvPHeRKlIn13nSknn301CfJC75eZFaMUdPGUCxpbZmQanqBpo
tJjXaP+/tMU4KvRoZBZtiVsU//MujpVUgtyzsv/8EOgDuBoajyfi910OgKCGlrXQJg/P/wqip4hP
XnSV/9zVi6S0xeQcu4KeNmxhEgDRIUEA+aAljT7783biXPI5pbxdAQ8YPg3LenFOT8K0ffGE0vMU
ZeBXF8UzkPT+trgvad6NaXqlVQz1Fi6ApuW4Bc37tTIwLGNfJnM5xtKjGFZxP77mcR5Dh4+to1So
tmgUfSgx5SBWhf5gkynjt110rm9/i+roaH/A3xF9d9inh/JMQjUnK2P1Mp7lFy6sUN8PXE3Et7J9
JUtqx1mSTombezZJBAguGBUyqp2p/5Cld6pI42D5CxbJwDsWSoFSRxH4P4PBnhC/2tdwdJNjOZrh
s11rJ/3ObqE9LHcCo35vQ8C0cCfs6P04ILhFO+ZUT1fp5c5qJ4h7eGXKBETqtS+aEMTptBwHBPHZ
8WfVi4V5rEvpOq/uXbzvsaZVFUmfpbbfpC8pUgdWATpx6MCxuc8l2080rVAnuUnB6Z+VrAcyNKmv
n9+xpSOJSi0Wyrw8jxlQdcRLeEXiHrL66i7NGFEwpCgjm/V23XEVmvkJlBhVgQOxTt3o7LXySbqU
5Ywv0y1OKWAHSt/UdBc3IyZWfWWi9kYBs39ngO6bEP99x/SKsXXEjKVfTISAQS0CsHAhDQorQpNm
yp4zB0e2aiuFumpexV+zy6d9pPfgJaLhs8ka9QJcnCDAbgvYCh8TEk4Fzwu914nHuMvGXDit2mkw
Oltt64h5eK5Q0fLIbDLQUGnBC67Bi50WpUGq7LT2qFrbkD7qVyJA/RHWznyv8qEw1wM699mb6qhi
XTDOOgODlLF3TnlSX/X8P3m0XqMHg+0Vp3XAC9uguz2QZTVfjXv8eJZLDPgukM0JpihUXyxVq0SG
CHAcKA44o+Bec3+GfxB+MG9aJyf3c/KtgUtn3sdFVL1yq+n2osMHABtW21M6V3/z8JVjGPtUoHqV
fK3tFlBMEIutqFF3n2kOtGq3wn5e0iXUlZMiVgqUypTxoKeCa4q0rCc8ctur5osiIpwPY5oxzgJ1
ItceZSuFuFtNExdYGtRCGqFcgFS0iSqDAvvom9peskYIKb/90kRChuvACmB5+Na3OvJAmdts/3X5
WmmWxlX4uZYe2CpD8Lzq70355o5B6f+zs57mt44MoPItPc9Psfw8LusfR8u8PoHkUAGXslCB99zq
WElJlXN/KY8wK1DonEltUopBUOXLSDJlG3Agcr0yPMGP7fxn3xgrAvLvoMbHdzVsCUXJgB7/G317
FXUVZHn87CM9pAibUZINVBcIrfiRb+qYT0V6mZaWEUyJV0BvDgwUgGEAcsEw9nDTE9l/B9BJeQH0
yzqLfmL9sTF3kHb6y48gvLfzBioh176adD7Ev/u/N3fdSMNNbLNapCRzazqFe48xyIsqlYeadSgr
HN/KKUg9dP6HM5K6+DOi9mTA7kkSoNge7d6HRBnxY4V4TAQNLtjIvzHMC1bImjQG+oj3tNVZoHz+
RXvfVlxCFgRxUeszSaG5qor2vIzyW+lBPK0zRO8L6cgo4YaehwXOA/tRnLDyxshp3vx4qCjpKzHZ
2vQRn0nOE5uSmxDOm3grrlOhgdvUNS1dqffOFdsL90OcbZi8519rWQsIpuf6do6sAh5ioJ8d9FUU
TUxF9q45raCXj2kmYuZ/94ElRNkNXdMbwaCBGsGctWBRNoHRkGG5FGWVaYjZRmSDvqEAPb95pIGy
Lk3aCYynqy5peSs/KYcYFEbw1lFYOo0jXuVS+ZG7LSIwMnwccb5I7G8UcTG/jjPS5XGCsJNwcG5/
NqUoAoK6IcR8nt8NvZZvohb8D2aKwtankcxoHbwM6nLPmOPRnHEjBhYjuqF0sgkEJriVJKbu9obR
M0TETL4oPfKgRRP34kyv5MrrpvqdkWIEhiuEWJ8bYjn9586HcfPB65InLPI5YwZQ/lqFBo1nB1qG
ygsaScjHX9novi+v6/YFXzEpVjMoR9wFpFGbj1nRzEHHELpN1914wuIskPOn8JyOz7P9za/pbnsf
vfeGfeEwcSo2ytvy60ntO6lsV3CvxgOoj5A7nY7arNgnVasJ8EFyoqMCdcFRg9KogGobHG86nwBI
8Lszr/npKkhs4KvWj3Xze3qVBWHSiWe6dJJp0zIZUs6iadHPpxce0W/WTuDWXliO6eHyWQ0hwTBr
eZKH1jVgeF7lmifvEdZEfmgeJ0vP5jeHw0pYVKQhWuHFy2jCGmIqEiXBVR5iduhDYRJlokC4uonR
fz/lpsRWj8y7f9hcwjjWPiWe6r3CUNMB4D7+/MG1CFT/okZslUrFRFxlGLY26Tj8P/bB/kV2r8uV
XkMKDKOeBYl0xgXnKhq6jMGq7qBPyJ/II5mNdgMiyh4f7rNat/t2V5noBTXIvcXuRoO05AFWvvPb
urROxodLLqhKm9RVa0fFRd6I+g8M7Y40olB8AG/+ivtH51dDrqXkKJGA6HvgKuQQjlFsBNkO1OhE
OQCN/N0MRFMggakxVJgGSGJ9PDU6zTWvpinOwab6v3ZnXMryDVzXNi//QzTUvJWHz5gK+wccg4ah
9Lz2IwylSBInAoLWkceWJe8lS94v+dksWHbz/Q27JoNYt+UjpXK/TOQsrdlRLUtV0Ahj91pMAG+9
5YD5iFiGfvRPH0GLtnvF7Hx9ZUWP3vHB+GT+e7py92sYI+kt1nrDq0U8vpxo1M3116bxyW6/Q9nr
YN60XssZykFviXkB9tqvaGoaAW6oPV4ApY+iw7YE1sX2KSFs/93GdddilUESkKK/7ahgVSjON6y7
xI+6MhkOkaWBW7sUgjYcepuEGSXgoQFd4JNzMmL3K65OG/U9Swl9MH04viIEYAJBf9wrhKJmAxxg
6gRrCC7IAjmgp7HwUPJKlyuKjYve0suSGznwNSGKQ/r4o2y3W4ahkwvmkEmHB9bnCJKjUFPURaMs
L2u+zyhuuqvAID4RC15S6a8N8F1TwrevhTIWNui+nPQVCghEwBqjMCvbLfQ+exckZ9bPSYFKuAPw
1YKUUPylopK+/sUEPBQR6cQ5FBiWop9oZHHISapDdTHexTW8kYuNaPcm+GbfWy8R258pBcyP0LTJ
/gaX/4DSM9wM6wvfE3baZakCMkL74FJufNt/FmTE8Eu0EEvYAgP+1H/0vIgiWr6yBe6yYRq42PA0
yLMzf23WJNsGWuyl4dqtBtPr0TiJMsl4Nz8P6UhzupB9pm4FEv49CnYmHKpd6uNaHDD9Y5vDuvs3
kuUjm4PCgOH3znHTO4gSSoyAAXLGi/tJjBtAFL2Szyzmzz4FUbKGqjRlwp3LQh4PSQNT0OhYOhnT
iigapJU4sFkZQOiX1NIhM234fK2j0ZuI5ue7LED6J5CC1LRVxN+wB/+plGQvJ90wH12Ken5RtPRH
jcd3KGk1H/DHv7JMRyQ14LVfnSBc6/gODwuanKAEd/S3HUngoos1NMy2Vu7rsQqo2EPhjdTJO7vQ
yNgtzurp+8EAdVXs4k7/nXHLAjetAsq0fC6A9VDapw0USO+7ewUmJNQICmwMYDedZ1skGZboL1DK
p+FBiRX/9/Of/H5fen6oindEuWDUv1CnB7TeUCExnkVEN2045kCvl6psxXP7HSBamubSa1TICJcV
8FZ6Dh0zPTwv2SPIwKdE3UMRnqRJwXieLUnpp+aNDOL7t16N825hxc1yO2lw6lWfLlW9TiQXzy1P
Z3AgVhop8A3t9Xb79MEAy6iQdQaL97xpqnWtifoBz0Y4scNe8k2UyouKTwEjqF20/IZkjVSwuj7m
FWlO8ucf4ymLpzSbuHwO114tthQGAOHLjjg8m7xtA2HZ/vNj3IYhTzG2M+t1SH7c4K3amSzqgTDt
uEPz7wZFQoJr8e83dzfvIz8K/hkm1YwsJH9jaiDNYnrhf+go2+iEgwV9RMrtvLvxSmw2203wkjYP
MifNP/OB7nxxSRJDFpbV/by7RcSqoflmmKgu2R50gCzCX3LLpnBsQndULAJhvh2qPwwgx+cyPLT5
cH7B+RoP6UKp99FpUeOOlawICcGg9dYJBSd6KUKEv0Y76FSvguWqmebwHtDJKQx2n/pKg+7nVvLf
pPdgS1LzJh0JAOVqHOmQlEAT+mtBYUndx8tBCKJOhT6N/N7rO9ir6AamKlTVKsVrQqcgygvhVXTT
lrTTrWzAdzBjG6QFQ8qhjgqpq+AUGZW6kCDKdVeafTu4OycwQCn3OahpXCVSvuMRnHCpmHw3G5rr
7YGLc8seglfF95J6hcQ7qk+KJHrKfJmab38rrT2cIDupiWxJussBwZuKiRoCJRb9SbtFH+C74G1F
pjC9Znc05wsaWhmlVhvk1K4qZzYAMevHEK9SnbUvYYxCVaH9828tnhDkbpj/ZdzxwRnMWj29Q3o5
bDK6Avxw/Yc1AVB9r2Gn6IR35jv8/yx5LcUrzmDW/Yt8XlNmgdwvggpIsKt5wdh/w4C+/ahhLzYO
J7m7e9Yh5UInNU1CTCNDy9B/wgy4VB+kNjOKunxLEIMX7PbFFmpr2wfzboT1EAuEqhwzLRgR58UZ
YXzl6l9mMyC4lqTdHTEyIVPeferjzk0k0zOgPMTiFteNTNmIZosgmrnGvQuVCG+ZwXDWTIJw1Mnw
pzQpzAw40qbESwOdTUyXmk2myIHqFibL3+2Y5+ivNnBNQGonfO/PHEYAk1vf93mLrpJgb6fiD/vc
kjTt2WyvktigCZEblDweMjqg35lRlOEG8a0HAr8m41udGhh7Upn9m4Rt0RzjQzLVTfJqTujl3chi
EYyndB326+CM5VGn1E8H5hhbePULMNESGdEnqEvGauw8s1mMVYWz2GF0apUZIGz6jkA1vkUOe3qL
wPg8f9vSJj0zABuPsiWn0TSi7hmxgjzzldrVkvGgfdYqBAnyzY3uEOlJ84nlCPoiJ4m/zQtv3le0
48scpVHvTPiMhMcFZCJvV6Ck7Ly1ulRBIfwTnonmkMvdxGv9OCKbfWlDv6EyDl7HFu+2YESJL7Gf
NHXMWBbrgqlVKkVZ5KvdiwDs/bR4r1kK0t62X2qqqxIgvh9nZW+jmPLxMtNXzhG3BjkXp8HM8LSI
iE0lxOZndUh0z7uzlbxIesB3T5njl4FTLzPSTJ7Y7YlG2p+uFUCzC1RzqhLUirxzAQqFbcawXLef
h1rabagWAly8EHbcuMow2jN1C3e+0LPSDXWBmXTpD9yB94dX7aY0zurC9ClcoS5l5qsE/F0JaCSF
44LYH1RhZhJX+wX10TyAhI+RZNsHKCCzkcgFZE7/w0QSHD6JFXwzOaH9s9w8oLCxWG09PdMv5YAr
xr7+JPJbUAr0eHYpn+o0iwDYtgpn0w3Xpv73KPMz+1rvM6jX2Yc6TaaHlvtukTBp1kOIpsk8JNdO
DYityrVgazzTisOkAtHI+6r2/RlmwAvnazma3pvBf006maZ3FpWetqT09e93LqrAmk9cXSpN0PT/
FcQ8iXrnABJvGiKQHsQJDGkzcgBA+xbatObGemeX0wda4X6SjpgY2JljyBT/ENejQ0k7l76KCVMM
na8rjVxsa2Iryo/k5bJC8sJTIhGJqfRBsbzUcAWEhIFofccVT+KXUcqqFcGxbMhSWwdznve6z2Ku
Zs7KSDanK++MHILTcTHt1Jyk5xh5M2ZIw4ExyBdWNgLF6ATvZ+Z4+Tizux8mv7pMggL/dN0JuqI6
2HrlZ5LMktOCB9fjzrQZDzHswn86WFePXoLYB8igRr6HNJacWLR6Ck7QIa+r59j1UC9Ms/Sy4DFO
EL4NrqV338KJWY5y0v9LTZJssvmmqfCvr1xcYRohBVGIlkBNAKHRpPQ7MfmaJE0EgwXqw+ury08N
syhY4TSY8mDmne25k419IBf2JUqLegUVeIKfpPx4qSuNriFXQBjAxskYjta8peplPqRIRHlsRKeB
k4TPZ6bzpsXVKGMxB55AaPvj8IC/q6ZdmJrl5HY3LgMAaXYltPTALqL+EBp1pO/nWHZhIAdsTDDH
U30A3hq76lshbkBMSd4ZEtLYtMhyrgWTzkOSYGsnoeSQca0In3HSiBOIH+4I5tc5lvFuN5eyeFSp
vIDEjtcFnOWHvmgzj4DYghtnRuLi4OdqjXvAKAriCQhHQ5ahMCSa2lYLah813YuLHICxZowdg39+
lPzYAG/MND1XA/lltIf2sF1Ux3BagGO35ZOx+EGINktK2E4xBC0IrzoX2P7gjDBa7AmFzyKM7zCb
OVAWLVvuDmza1KPpGnbG/f6HRnsGI1d8+PO4LJ4DG1MNzEd5JZ/3Pc79o5eJYAtzglwmwa9/EO3r
rIrBE/nN8K+tZpmxpHNh/OQkrL/MCm9+QqE/6qSVPMHilHwXfIHY6G9C0BVL+VOqREfMp4OEpegg
EdsDNIZxpNvxf0qCWYIvi/CPU9wsS1ibzSKZZw/v5xofqhTKvkOi8L+2fr/LOPholl46VBgZ9QO/
68+vZNnpFvXkJBtHO3nl3BahJsLKZ84W2Fw/0dlYuNRRPi8EKBinUcJk/R2X6NFvXxCGm2uunfPC
hXz0Xdt+JHUWpng4hnmq7sX8Ue1lRo433sUb6waaC2Z3O/LnQyLOUGH8RmX9vtwmZAM2wn9dX+uH
URQ2JSno0REX8VkzWt3BkFR8alCCZpVsvKoK06raoqKV2x0LvBlxK5AuGmVmYI+96OcuR+27jhIw
ke1FBCNVCTnhHflBGw0veAyfPLt58SXT0ii83wxZ0D8XseDNBPErhsJHjhBZOqG4XHtieprgjqBy
lVuGb6cMKCNVUO691wgBXBgKkoImEaMx63vbSG0fRvX3O5LB4pmOeS/4rGBdxz7ywtXzSmvacpOd
qqKIbP/aut/g0Ut2J+4MDighE+nvyF503Qk3Yj8MHV7A+Htrj4J2OWOKYAIH9sRI8hAZqApLlWR4
mm4pBylFfUj3KC3XHHzloKLz3gv5rKAO74yT3RXwy8aaoSDDiM4r4LQFKeSfgprZ6FD56dq+pMeV
JlWcMZAGmoZQWBZZT4dxo7DwuAnGlJMoyv++uaIgwhND2mt/adCgyPYxefY54kjwsZHTbTl21t2I
v0nQFIo7ZpRm6c6thiYQadOz1j4SoEpZcVIEQvm7T40ztY76qLJA0+DNsh9d0eaCJNd/6ZMom7jr
ChiecPq48vb6VCYlKYbvX/svEoJDJRF+OnOqx2dWplpGrzYLkdOLyQDi/X7Fv/Hgi0fd4bvTybsq
ElmAVQGwbbJkj6WHgc00R/CGWz8JvI0Q3qWesRAJYmSk02XW1t526+O5B7mbbxa/z+l+Sswmcp5q
7nXY5QkVGhiWz2YLVwAnLhTLPPkVylDJkybYLXXfdPK/2AwyYZsHUT2p0TXMh6/MZ56slkOYnmEa
AJUAFP6sfr8LmpeLpqZqHNQevG+znigjEjJtRGkm+Hp0h/zEIh6MHSUliLdbysLQ4Ag47XyQY8cq
teJjdFXOHj5lxjv1Idg/UUgGp9j6IEi3JTEgRZ4yrd+TPuVMPlPgdOC/3CNSAGbJF0Sj1PByXkoB
JopgfMs5UHRF/fWl+cA73hkJQXfS0lrJewkDVFtj9dML3pnd79iImtwxLui3P0Np4PFdI+tbUswt
nIQQA158Fr4+aLzCzy97iUk/Pa6nYuKzZ+4pZBJsd8YOAtjaXrOjnNZO4911YRZHH8p54TGUE7su
pPdA2PpzcT9xGNuS3BcwBTtVM9HKNNOCsrKplk0OwnzOApYvrKezgXJd4wGPpU8/uMx0Zbwdgjz5
2zcRQCyZkM3bGcNzX90duCX8/nDLo7CpyIsTwJRPOrM4MGAPaI/s5B7kbXO1Og/yO/0OMtN+CAeG
KTXf2NLYCF0k9YPvjJCUFyVQX0J+lq4pwawnFEFlvF5fbrwVlTYp6oW8NAQWyRsX3gr59iL+QAzm
SXfb5PWk83DD+alCQGwPZg/t1g61khDtB6BEnvnx3on38c3emYCiyGZ2bpiMn2TXD9ROhVzb7ndQ
nM43c0magfMGUT9Oc6FF43HE55+LWJYmjWStvz9AIg6oiEkT8GbhSmrWX3wxDKlFr8r8WNgEFnSb
nR988U/oSEGnLAuvnszVF3HqazTsZFz4STDNJEHBzevOT/6MsRFp0wvGOJUc5x4U6sIR3zPE6QxR
6lep8dX6FYSztoknEYLEre8lFiscT2nNuQYDPS5paVB+FwymDLmCu+zh/BBeT8KIIiWkidHpcEgk
EU8Rl7XfU92tEWKzfKuyfxoi3DQrvPD0iR8geVJkqsDa34CBQq5aUK2nEkfC6T8NOFs/q1zxfX0w
6I+wnkBnYIkR1opnAQyPxwOLLFQy+CPfCMNcv1OM6mMBm3IFMESzZdvILZaP4P3NnQH3yeCtknBW
f/XfG1RW6NV2JhAum6Hfh+x6jECUJgCtzCOdL5RdOkSz3LozkvWlcLhDG+cfZ2jNGHPuA2mh+Z8Z
Rw3OerAsRGkUGXb2xxGDICRw+tBjVXGchm3E9EWXZp38xWqXyNTP+tkz08prJHJixLK/cu9DAOHO
Bgw4B7yJeGx3LSprOhrwXuaWBDzY0rwWpGUPb/EFd24QUXdfp2ccGExMtQM74UeLsgsUMX5jakV7
l13nDs+YRlIAxk0W5mxezvCM6kGYURMGlUER2aBHSJvKCpnJ4dVeL/JCwJ5ysxJ4PfTPsJT9WXmY
xyi+IkgAUet7WFmuCzPtyoIoFUG3ITemjF8gXgwdHCf15fQYo5HnR+EgbLp3184MrKeH3TAOP5TX
wJxkM4AV1dVrvaQ+UBTHqbhqa0CJRnMVfoedMRrHcCBydSANhZJUlgyaJm7P4BRMM4z0Nl3hbUNo
0l/xvBgFz7FLTz8iI7k5ZMb+OaT6SKaJ2v2hQ/KI//lHaMt2JjvxLeYNIWPuPbftNOvQXqNbHV6B
WkWgwhYG/oKpbSJNtEWbdD++ddIor77oJYoXwq1DaQ4Il06Z9erT0Q2//A3+/2h06/MulWwT1PcB
GOrOpRE3hcHUaTe2q3oKnaMXDJlPUjH/MfqBYNUYFgqspyPFAAatqIOt6NN58k6KAZEi+Gi1tNv4
zkCtJLErUf2/y1U3ed3ZKzjrP0iNYjwhvFWTkreLoN5RTTGopVSFgWx/Y4BG4lb8ygq4zDOzXSJD
cOK3ROPVWqKi8vveD5l6u/iB6H0LUpZ4tbEzKiBvBnPz1FAGz84kKZPzsu0hpPecf1rKDb59PqoI
zhbbeKAgeNNx5BhNgEc+pjj7KecI2GjPWo+OYppNpqW9rfsJiNP0pAeO/ZUJavrMYVbuugluH4pk
tCYoR1M2xyuTjr8shA7j4Wc//W8D4kQEXiZCZ5vjVXO9cYFff0qHWF2noOzTPJacRtMC5fPIxSI/
Um8hEBm7oIEUspxf1DRB0Jv6gJYe7qXb6eWkj/rcGa/3QbGPY6R00FXinIrWMcsW9Wd12YG51QRO
PYcfV0lgMHM13VB4W78vXo2vL4TG68jYx3FS7UGyxg1UwnBm9n8zji3TcDHv2XNo2aM+r2x1RDtV
f3KjW/6sBq1KCuRSgqvhvcoiNxs+Nz3o/fffOq4uWLOaezUE89bAbqsX2ef3Nf03TXHmsrbAxHct
UsC1wY3WiVnpD+phCFQ4X/8gI+yYHCtlKUPPjSPb4Rue3VvyKkRjMQmn579kMlxUTKRH2jOWXVnF
RzvfwZqRIi2+Cmbzl79Te6pQZPtmqRisqtwzGSDkyWOBnTIcAgqhpxdogkLnMmfwurgxBQ49h7ka
Wx9F1WG8+pXVLw1mGh73UMdWq8LyauDVxmZaP1fugTfNAp7XrxIO+ni7txpG82qpeJEAMErTW60F
duTJmaZdGQ0OUgXtm7Cj2AKLBBTDTuDEw1p3FDtRpAgrGW2Tr1SSvpEBbocdSlAIkxAibiP+Ynr1
Wbqhsm5N7LEicXCB2gtgyPlqmVEHYWisnqhfdPgBoToqvFWvHUL4RBd4n6voJ/1lJ/oLE4WZchtP
AThevtHwe6LL00ia5aj6dFjummLBPF2SAKZ4qZjZrdfAep/e85wLJ9s9gwV0JJnsNtb7v4PMko1E
rOMF2rrNt86ZssjNClvo82PHMMl/1jQjwEaY8J2Ot5E4UZ5gfIdnN+uivSyUs//DfeBGK54jdEl8
+FiiAXxovdFzjHNqRIZXsjIVKoAhDJE+0/fD65Nwy84aCFa8Xj2hc1nRRenpWHTVLSQOw+5CWsNS
ek1U2yZlc53Zt3d1EhFRIs79cawtqy7UkQ8ZR55iCfYNB9oM6A8qfWhjHzl43fM5SAIy5UAhQbax
AZuz+T59W+WJmMTz320NGVQqGLomlMw7/sxWke/2iJ7wbeZPe3dqsfvN41zyFVRV/rXboIJkYPK2
DuUg+/BQtRaSGjuyGUdQRMR1cCBOPdDuSpfhhaplJKFqplNjv9hxKyl4Cpp1Ih/XvnBl+A9WFNgs
+rMJVLHjoExFiYrBcnXCf+EU5BPvSEXpPGnj868vaAqU2uHV72M9aNVcmhQzePFLbJ6kkjnDFjCC
AQ8JP+fR00qJWevby0iiawsn8x3jXr763hFgligVlFUGPmqv8dm6cSBbeMOs2lqQrLiYbpmbsMdg
hIeu6W2P6WHe5lif6jdwezbAQJxHGqEm1iW9Ay2t0BoZcIYEwIcv1TT+btcoweKdTowkf1R/gVIi
mcQLkeL2XkH23lBpo1TEjc/GnZZ3M3taGSQXQIcMZ+WReEI3aUGYH31PSEeRxFZZFn4rp8vhBr3j
dLDWt/QuBmVETG215ZivwzzMC8wH26mXNYQiSG3Irmzu74i+w3WZlDHA+zDkrCOf2KFi8nh1av/B
d9tiRZK+a63ovNfx4azDryzJT3U0Un/XtfcIqdzAwDKfj4jizhDIuaErEkgFlKom9wOuLGJ6TJmW
6HSbOG4e8qmkEXlmVsNrckYOQcFTLiBs/oteZgp2tCmnT0f63aMvLFhkZzC77aWT3ssxvhXRwKG0
Ol2vZT1bjNoBhhJEwEnz9BPqqE72BZVG6LkGw3tZ7v6e1D/bHDJ3JkRz5g0UtP8P3/2EbxfurJqp
Md/AjkscI45eT5eZELh4N0YaOG6crjToFF0OZCRo2eXXVBj4lgKzmKQ1c1Xm5HK/oOtJfRDaWaMF
r/PgRCgrPTplkS8O0WABxMyH1adQcztnGe7VmiMI10ijHtBVHE1KPumuNvaFvpmbdcRVblYsHlQl
Zuea83UT92eY/1/haqlvQMil9NNkFcquDOxAULoMHMJ/9qdoPZggO/cpTWTexjefZ1PBXBIFVlRM
2ZwD8EmpsM6W1uknTQN5YQqK8yIcmlVFl4qjaMAyad6TTm9/ZjzJxDLxegYaDVFpmjskK+WF5rML
F9F9uuL8dSdCusj8SU9I7JT7gM4ghcPKh7VPktBJSlrbhx94uDGGzUtV6X8erhuNXC/AxDi2OoVG
8nu2GdAFaF3KCF4nA20B82ewom2PffujrbBdI1M5t7XFcdmlV0mAMSkp9RSIg1WXoeDrdWIM2zOC
6raDOsZwbLWR5JyOaI+gjQ1uPlC8nydlAtuUIxjuvQc8UV9g6pXrnI7CBUkf/jcPY2R3cFZRpyYU
sVCC357l94Bd6i8GInWM5lYnhF3J+6B3gSyI3hpoG3vpRcXKdApW+7uS7IsLWJ5JyGEmU2JpEUFz
km+UzWzP6fa/osUZyCYCaJ56rKfUTpbpUJs1lvKWdyAPatrIi8gsW6kz1WD1ayY4zoevLL1DBoD8
7wIlNIbpUMHUXKm6GWpbrx3i8GWQvG2BSyqlYCzTzdJg/rZ5RjqwJBlDFuJcfyzMHMiZrLhmvLl/
zbmda4zl2mY66x7OwabfEIWZlhvrwkaIABSA+LGM+q1AfXGOjbSNdsTAyuiCSFvtZz4HfDUKAhHV
iLgtleaNZf7JkCOXs9tVEn2T8yf5yYWoQmfPuuRxwKropSTukw7zypmVOtQ6/4pOEhgywr3Bw7RZ
kbOH6RJkrmrukCCSylqJsq/XRW/UqZLSoC7I4JYkyf2VJdoEitC2P0igEhCXlyuEmWiglUU/vVJv
uSgCOq9KpOvSL/0B4IakwTCUedn5tLOFYbwUe0UoQsLuVhGoBu4/t0cvktmgF2sesSlRQxlV3d29
G7+DAxYXKCEcffSA2s4U2sg9Wh23BChtrPOy+3sDEAQln5KCoqNYEPsnnp9P+FNpgvHOYJCkcWLC
woTE0QjyJY1EJ7vbi/JKlxCP84pXY3wt38mcJAq1rhLPElUkMTtxWoO6xsfu1lVqvpDPGvn7Sa6F
Mw1QoEXo7/KaOKh0us6M5nudHstPxSOQG5+W3gFMezUsQvYlfK179HcwBsHfDqEa0/FOwJxwgH5N
dgo/CoyJweLDUNY25y4vclBuoWCiwnXrQLJY+o/tTkp09fFdgHoCb8rVzsyMVwE31Q67ozOXrWwu
C7A/B1efJXTA4ll6UmErplrdd9ppJNWEPRHKRAk8gyF94PZBMFxKSV4CUsHvBWQnD6M1PsPCgDER
Mk8+Phqkb2/aJ+5dAj5ERdADtGatyIFR5ogOgzjo1q5myE5qENjZuXLuXt73yxRnj67F/+BZDeIX
Ri449Mis+JZNvD0xbhZzJVsFOEVZyx1gVhWz/zgDIb1zHwOLt35c+BGrzrlbMbMYUIiYHlwO6Rc+
ZDfev5d+5dy+oxHRLiVxQ2Fyx8dzbNdELHIGWHSng2yeyVsV5VHDEwv4dOMUMEh42xKZO8g8lckZ
bDHdmJBySF0HNhW6ihN9u+9Zq/GCqw6FzTG17tew3SqZxPHzXRcWNDv9NreCs8xHlvnon/B82bRV
79g8ObN4HmoFHenI9PYrjDZtj6yrVT4udA3jp6Mhn6EIvNp3TCLq9cFLLq6jm65Zc4rt3BvMqHPH
YWvax63cjzsHKoBBhBOmuD43DASHF6mVtSImP6z1pO6gTMqVQBz9Go63CnzkXQHh846SRl68IYhZ
5HC8BY3rWbwoLhZ51VYKDzDc2qE0Ad+3EO8F1+ysVLBb2X7Wn8FDnip9nxez69lQZ7C8GeZknfH5
QvurCcV1kaC7h8VLf5Z1s0XC3yZz7PMOV6UOZX9ApLhQ9i9J5J3fP2yK0NXjksvOsoMi0v8lWBFP
Iulv8mUx1uywphUFbUzhberid7Fr/bagz5uCWTOfvAFTm3G+T9jsSS9pS6sRra42UO/KDRb/bSIM
1JxFFRoKmCNceKSgSatTrtMvL35IojjQrUX13+jkjTpAp/2ubvlxJ0vof5Wr5cA5D0k6aHklseWp
GbiDgldy0U1x0MCMwM8GgozNKFAjviG81HJcUcnHDbanftG4/x2zUyFcui+7y1kABa4pR4uPXVnF
xyXIWWQCk6hX1jIiPhcaTdOM42r8SFdLfIP+Oa3uwtgRc78udfxwCBkXhQ8kLYNVV3t1vw9v8Ocs
6GA/juyNtIpM/wsaTmgvsOJ2rDCzeybeuxRQVm4sDYUsWVabQqzJLK2Oz/rALEx7WwT88B1EGD8k
xzOAlKZvyX49xXU6h5TFCceqQPbaaeVARiANMVQvjVk7f5F93yX0q0MXlCAOKgxIUIBSewE05+P8
ZPO0A8wT0q0HWpb44OiMC+L4nAYPnFHh293ypu+s8DNLq2O6eIGB9qrMtbZAI0Wri7EGWx0DNOSJ
Ggzt88k2jhBnXXNnBPJOoj8tOSDzstIEb0fGu1IfmvryE8sAo7ukQAybICH5inqripTEBzsmghbk
infrV7+tLHWBlezS7bgly1Rl++SyCd4kbRukzFUrRNhpGwdvYeGC3nalqn9zPRTIEsk2hxGzDlhX
zdG+Enxvi6pIcaXNIu/tt/onDC3bDBiS/2pPYIFDAVkJXlJQqaB9I1CkIuwjHya4M5KncINk9Ppp
fYrN0clfNz/k55xs8HWOYZZ9ClUV//AibMNcOkpTi1a5uklA0V8FzgsKfVnre+n0fRXVFQCpI/Lo
jxKwvaNlc6Ff+M5tONTqfUy7HCD/nwgM+9HqDgpunOXfuKNdmLRlNi14dsgv7kfXnLgd46BBq2p2
6MGLEvxC4amCjyEZjSZ2Chjaua4ESKFZyKs3l5MpDqp1kPes2G0ielAF9KICElhu43k9sN2UAMDG
s09j/W2o/KM3lLvFf2LiYYqoSL6I3bbCC8lr+I7E+L3b89uIHp13FNN8lEH+s7J1vpMiVxp2rl7e
GYlw/4J/SGdgw7uyDSWZ9mS89wY5fOSYOD7PWOShQwgLP/JPUrpTX5vqtFbl5oq9KFkw8FNCTezi
D2w/p++UWI6yz8R/2Ys3QlFI7IyjkP51vw8RyaThmd2WKEzB65dxzMjC2cYkt5r2pdnfM08mrmMO
lJ1Wo6CA8adtx2MhTSb4CVIErkdUZxIWPtP5QoSPGkCeB7L6ZjiIbl8IrgcW95a7i0Hfs4kj4ByI
ZsKzbm13jVPbHJ6XwAPemlpHl7833RXhes0rmjDrqEgcx7coBQYmCM2b2PW/eEvag9kG9RmjxRze
4Iedf5Z4/4vPEUWPuKUMe/q6pVy0UPhStksajd6JfpvGAzmEijGV2p+EJIcTYbqYpUfzCY7lnKGI
Skwie5xqSnxNswa9MVwV5ZCN8dd0Fqwrd2Dw6qe8TSEyEfIR+j4FKvPTjxSmWr8SwdutTrvI/YqJ
Gs9JM8ZAlVjUjXc1DpVo7RGb0VgWU4oNyRBRMj7zbMAgtK7M5r25kUjMhSqwqXmuygR0gPrByQU8
4z3zrBXf/N2EZiVNQqOsraS1MpUve4fq+V/vEe9zRtYhp1ZDx1ALky3v5ZPt7wAc2YwKbGwWQcnv
S1b1aSMaE2BHgZ5Jn3o78IK1QWN8zVLcutEPfKvnNSyqJx9ZIRQ1ofVLtUjUsqsiiDMW8d11pTdu
Pa2n0FN0lUpAM2Uzr5TSMSvlGkpHr3+fm6prFWxTqsyXxjAlb/3FUMGxXIsRuCplX2aP8TMnP0aH
JqDmtcTNymQ56ffRKzhD2PXxAAygBaxsFEt7aZtXeJpZn0KvAoPuA/kQPF+Nh61VF3iJjYdZmk2W
xhN9rFSExyz8EY9UCbtptxFbZ+M3v8uFc2o6Jfa4YwozOcy5cf+Ch7wy1wnCbFmDyym3wspT3aKQ
spduOzWAquKHSVz8oLIJHU66knyq8as7vq9zmluyoIQSX1S78KjzjMNJ9+mTpbxzN6869gFbFdbE
lOubVu7/acTkUUXoQZniWCrD72IFiImFFZKKzAN8i+NyB5GKnGE6awcPC32aCvd6srwIue8ZNGyc
D+Z3HpU8/neuoYWAQ4vf2RfirHFNk1D+hCcV2ZsgtXpkbaGrZ/n1aDVj7oZTele1siqf/Nz05DOC
vt/+5c/Flm1uFELfqRAz1B7blKjAewZvIfzJm/NBKK6hdwSP9Gv0GeH5bLogzTd//tsHgncwxgD5
5l0pIYeRuPVZxceJHEd52UUdA2WSpk5+A2BcygS73Rhk4Nc5/xcXvEWV8SaygQONp2eGXaewoAM3
9r8KPQZLGbIM/2EBIal4yTixj29ky1BoaVkFOplxFtgeMYCeYMyCMjz7mT4xhRZMq/xapw/uc9TC
Aoa8bM/cMT/JHSiNHlcVFzno+UYXVXoKkKYdlE/IUn+iVNxx93IIPUtML9x1BE3o/QUkSapS7kQ1
lFaqtBoEZNHvtQkYtMBCskRyXUuA96Q6p5XbGqMOzzV7jEbT8F0k2Uev2cpGx2bX8/yW2rk6BhKD
nysveZe2h/o8u+BajRTSI6tlaVEg+gc62wVH8e/xum+iOD5NIaqfFtVvmsJbrfHctHGlqHNJ2Lyl
IVyfDosPDcqIBQ8FsMADHV3igW7vuRBFLUsUO41S/0kfHzHpv+DcDM5ys2X6BLvqjITKYNO05giq
o2HeyGfCG8vDTjqTBMj2c88NHfNxvVYTHMsZvEancFbD1RaXiM615I94aWBXsnJOXgLC2q3mtOdt
bzMh72r5DbmgHtWG+aP0fFwvWiTJjoAg6BKvPP5ilhIvsAatXwST+Ai6/x65GWV7qFH9yZJWzT6i
p3AdFIV3LTklXhCNKjToYEMl4Xz7WyWojFvlfJadzcjsdyI+dX5aPwsf9Vvfysu4xmzjYpfrqgoH
eq55pQ0d+k7x06RCY02vrHpJ+MDnRmwlKzCAZwUvnaJC0ePLXxfB/tQwoF+pc4deAGLid1m2zUja
VOgaw3X/d0NdoqE7CBljdBWTq5jfLhq7LNqZpCR08cYY56b4iv1j1FcmWZgeSyrYiuVg6sRYO0ZL
ifmcnoNXhOtZbYnOHLFSZxNfmVwRYJIO+3MrPPPzggLI2QCbr8fEV2yh7Yown2Dw/KsBP2I/hLJS
mj0Yv0VVLmRGIlKsKMbLO4lRZ8BPG4v4HxPHxTvCsW01jsAzlwcV+b+WHr5uuqjbU3bMMWLqBiSv
NAQ39HsMiBBJGE14UvkTWX0hzi7Vb8NA6L4VvS6GzNeQPhfOaxDfFCyoOyj5oOrOhJ87yKbAHH5z
CwYAaLITebR5dQkpaYBZvJLRPFhLKtyZcwrkTQGO1GGkvQqX0fSHQXsiAfmSdLZBrVnf8QsjLFlg
LKSNJE4j8vYBIuP/6tHiLaKJn3h1ID2ZOCrv0+iJDuHeytz70d/i4LlOzr7eaTFZszRg5fkwj1SR
B7Rvt5RpEORrLK49SzIAi98UsVb8IxZ6j2+pFrA4uFsibE1PL2pI7gC4PL9d2m9ivpI0rE47mK6r
3STbeSVWJOuYq5PPaMLjCmn4uK3uGZzxbBGkgNqDvw+HbPCbk2bPApjeILSNnGGz/ZsjCM7vEJUN
ayMNeQGA3VRe38RS+YfvtQX57RyVhQpYTKCgpfQLk8Tl6cQ1hDp6LyGHJaqBCbc447/ZrKdw4x1D
/n/mTAiJ4eFexOSSGhZzkwJsjQz2kJex+XZztqQZKfQ8XkPDIdtutQq2zxue6QZgiZqTaVZQurbl
Rx+NxSD42ZF4qjKS7aqQK8NW7xGJNjSXMo/f6ng2H2Ty6K7AzIsBNFzRsUab7bRm/jBMgrSGSdZm
aBVqgKdNu8P7z1ql4jpevXZ9LKfEtmSNm9pPKkz2iZ5AVWpv+fX4Ew2IOLxS4s4eSkenyyv7QTof
9M4tvBk3OZSLI6mXurcM1ZkcC8y/gZqJelqeOFEoRVber/1oUCpAefEz/jENT0P6BX7qymiO0vI/
z7aVkh089tyjEBb4eWC+u5yqsE+mNbjmkU/deq4ZBIy+eK9Wt7DlHEXRLX87kKGAbQoymnSRKw/e
ZOW0iJP+nIduGLSXfuwmTloU0DvzmlruEx5rOn2do5GAf9zzgBQUZpAY3DjhpChfuYMDgfXP2tPV
7COO3F2KpC97fM+rb+DBFPegi9wmqhRWeRWiv792cu+8Qhe7/gmR39y6lVj/oXMcvvSGZTJIHepE
Lt7gRJzo96VKGefCblVUlVV8a3Jpt/0FHr454VzTWu77PfQL3hZjTgN+QFG7by7iK8JGCYXIVxkW
AIelJM5Wnf18yUI21UviTQ/uGPu6CQPSr9NG4IpsGViwwH+9e0jk1214T2xFu2A13k41C2f4UQG3
0qpD69RyGvQzUe0bK5h9ofNoIm3zpkwhHnhVCqWqHr15BRtA9IKBzvWgKvSY2AuDcR5QVrOyDAWk
epDsavAe32B0N+82h3DBZiBPDCi/TNaR8tHpnnWQXMudbZvM6mNpEv8/4ZwYzxp+Xvc4wBFMtEFx
wRcaxwH3HQsRX8+RSeF7thx7+6zuMCb+hghlCOhOVnhbjUPScAjp/jfVknhgobVmdTyugb5I2M2m
F5bmSAMY1fYOztwXSc6zWPYJQvXIXvgl3hq7p0OgI6MuUaR3r39QixEr4GQwHjbwrpBscEa+Yhlx
/rlNpqnZKDtK55ohEbwzXgVixeCwpNhBLqPF6uODUpQkUX2BIh+06Aep/BcTXjoLWFFN+Njn5v1K
5AVFWHtGtmNUWOW2a0/KyRLbPp8D3bUusLc5xHdU/fClFzGwa2IfmQGdpV26Xk2jt8IceUizR1Ad
9O3SsSxkZSqIf3bLbZeKIL9vw+dM2Ao69Hfso0gaVAZqYz9XQhbr7tgtwzVLS5iR5PM9LH8LrSaY
VzIsVbPtpYgl/KFee7TtUk87ZeH4Pnk14OtMve5SWJrVM15WZ0roq4RxZfocCO+Cr2ssW4HPw1u6
cb8v5GXemBLFxSIEe/koZByoYL0x9UOO4WKB7z/Ezv5C0uHCKFD2pOqCsuHppyyUudkorAPY67x6
TLVIUyQamB486t/7/GOiNJAiFcTUCw6IncefY0dsc5mevs70y6/taJzmLFHa0A+FKTv9lNSyzMnw
XddQogdJ48WMtpscRJmSTDN5nncc4L3HaviTu87AcaQ78JF7deV6toCNbGOVy9+itJb42m6p8wYh
EUjR/s8HAPZDcjMGoy9tdEQ9aX11ZwH8bZXq94rHOLnoedafj6KbdFGghRnzx4kgmgWP2x/3i38T
jk9puR/TFCd2k3A+tMGLUU5k4HeBV+/KKr/Zx35s9VeOtIZs3cEtUm1dcaSnkZ59+mIjE7Xkrs8V
kZZLGF8wSL8fZfTYZnhSuTxtPhXzn5cg2pxQsLbN8LWAy0Ei/hfaaa468Qp8WutYpCrlqREdNQUh
afijXze95E6/JcGVRZtYbt60JuUW1/XOpF3wxXMc7uiTtSXCLWRjsAiMPrmGzlFscMYF9+zh7z3d
w8MgSa2sprk4RuoigbQ63iiV5hKBRE+yAocf45otkqHR0BtN5te4LWXTrhVlE2ZULSuX0+Zb77PR
ydLujA4Act5bbfRh7q8aQnsOy7c5yznG4FcPtWj0Y2BCRINOnEwZk5KLCnArcDFBWRYY1QX0J5To
Flt3OU1WkV3A0i8XEzMPvvGHhCIPTcCs4dkZeNIXqM7Nis1yM2/AJd743dRqzc/WNi1BQ/Gu3It3
8mKWeRyJ0cAnMcHYD9pcJEXzp13E2/SnxFNKUhb+l6N7d/dhiLQU4jxE6nUWMu3GgYXXuM+OcnYC
hNUtGB8yS/iLctPZseVBXYg7RFfQ/Uuk6HuW/OaGVWXKUp/P8ETLBAggQ5w9lhED/IDQkhxF+MWR
Bjleg9MEX2Hos5XAMjBypeQVZzDBUn6XfxKRrUUP2y3ENAaDHLsVPg/AfpTqSviIMBT9i64ceNa0
PE3rdl+Q8ynpB6cPChk9Nu73TJBnyi7RG7IUkX18Y1H5UWXGIhgNJx2devkRGhFql7QTZZBoNkEu
UsZyqEP9J/ArT8AOJkLZBrtRTvQhGv1iN1UO9mDdHfy59MvTNLlb/zQcEOTCWuD/XMGAJjaga99J
VlR2kJsnriPxXE5vbcHDPT7qacm1/zjeU9vg2Jqa1VykF3qwIdX96pfW4X9e0/IHHXoifXBVnXQa
LM7b0sKuzeAHUDP7rfuXWPLWyaFAqPPe909c5HGLcWc/AYB1r/ymouslBqYORuMUFvKcq3TdDblF
uqqOeJGR+1DUhJkoTY+Ggg2jwWkc09M9k632ebR0fLBE9d4ulkqnfYXAgD4opyz8mhnDi1COpkb1
nus4KhgdlDOgJmjGOBRPnZ9eD0DvbP32LTzlTDhJTaYcg+MacoAvp7XqSnohg5VN9AzsBDqqUYGA
qvdS0MeujAE9yqHrcFwWhzgpku8jqTGRgxvHzU/HhKJJngKf1ucfb1vdeTIHKIsDT9Nkc+3QsxDM
d9ntpWYe1qv1ffzUJtBDXE61WeFUE+qk0HIriipKuXnQHx9cO2mysgM655RTSXSlkxlUb84plwUp
e5T3+JVh6BlbODBr1pkWG2IZ6/ecXYsv/z7jLVJneBz2Pq7nG47ksgNR/JVaAj18/XbwBsq5nUgs
GtcnnRTb4j3q4AURMK/8fYghIGl1N4kCCC7+a83UcW7HqgpBWKyJ50wHMJWNJbtC8y9XcvUhb2EJ
wzbEhLkKesJQWtJJyuxd8p7q1w/BupKJHAwYcnL/QXT8yFf/YaXi+RRPCvRzb9NyyceDdozItoNC
YSFmp6msUSDVtHHctuOydhOipJzdcOkaqQ4bgcritZYqGZFdeb+WDa2K8pxOXywRo+kWtDjyhQZq
7tUqC99qVzc0L60sKxPGNm39GxLVxLEHwKdoxj90ZVxkA3TuE5nXgNyG92GMVxPj/nkkzeygz0yJ
ELfVAhoNzYm7taR47ADVcpTTyX/9e3rdd2ziBw37xrf6rMlK/P4fKBbfvwGFGwvqztj90m9K+f0/
8jLgw/FmXZKnNcwia2a7l16pMNStibSc16s8k8fsPf/+BvIbPfJFsgD/ibacL2zPqA8KjldZedJI
codl64D9ZXtYiptz8f+Xgzxa0LJ3WcMomKCNqO6gjHOnSnWv+IcBqNGjcX6NWJawF/aPLLt1G3SO
7PKLjJkNVR/ctf0e49E3vMj8WvNLBiRXpnr67bPE8z5iyXsTBDpt0J45TXYz9Dw1LgG+z6ThNAvW
b60d/8kkql41l8+oD3AknIfd21ZUd+yCUChNZBHpjLaHOhqYSDqBh/u2SJNfNmqGYq24kbsQ7sVA
u7XXNihuhU4CbQ5dsVgpXdBZYCF4OZjbrV2GH/WXUABWBZHjXKJtxL0mypdFleDv4qen+a5rxqje
vJxn266ZUWqEbmhyqI1Bdar0P/NbhBmDDMv2Gj94e8kUTd+iLeFFKHlvWx/0bcpZyMwTXN6jNJ+Y
t4FeZeM3t1m57JC/Ae4ZDtSw5Fxvp2M9j8+Y6HixbfwK8tEgIaypfMMl9LN658SdPLm/y0/2khD8
lVOMBsyNAWzkE71sAuPtHYsZXfcDrgHGOJ7MMdSA2Ilq+Csc1Yx1xgvVE34rFAUQzOggccYvEARc
+z/pKIXXgW4cjeArgeFwEgjZSgua/bqQ8Arr4cx6l2HePNN5G9CepHITMM5A/d9R8ZUrnQMsi9NU
Dq6hIMXjfXn5SC9jgR01DOgZ+0K34A3M7Z1HJvXKtNHx2a5sBxf8eP2KM/de+rcy97VXyJLtjAPZ
CLRx3y79qz6USj8FN1xKOWvvy6U6XODhgX8pEGExjpl22wWRWBAAAdJ9fCHStZzPZmnuiME+m2RI
z8hzpGaEAgEmBY1agNkNfr5QHgOzNlE2QILRPmSAJi2aMTPT2aow4EbFlW1DfzoXDv6c6in6fYME
7g7x0TI3AB7C8rNC14VI7Y2ZJT/HcIS4u1wI2yLFVodKb0wx7Aau+yZj5+EjU5GCrzR3dmC+fzud
oih+lHCyDvIO/qjqNVNW59g5c9zD3brak8nEHG3dchyWwKV9EqcaWIClDGnt+B6DWWCWpYCoCU65
tny3j2nCditaeDLha51QuDXYy2pZd8NCNZhrHzY1jR6GlSUo8oAyN5EFxYEZPlN/9oOeGw4NnBPu
VxJeK23Vf8uYerl0MStRyiNoa18odzS5wj5k6LHdXUFkAKadYYv+UMhZMa0z2lS4R/zPdDDOVae/
fDKPjRnZQt90QrQcCpZjJXnOiUKAsT9oxQxw2qCemJ97ynvnADICTTMohpRdN6sNiWPk5zNdoHln
5Cxv2jNlVmFgbwuUuQR1mLMh2x4FzfA5IbBmY9JqaHkhh7xRebLTIIA3rnJgGLPidAkHS4ELug9u
RV2nDgYzca2mdidrxmxsX9OoN7E+LT8qF6y5Js+kdYNXYTu4YJiklte+80BkCNHVzD6l3OnpjrHZ
xIHGinO9cADMO//YjCg6Dp37f9YPbMEtvwKPqOsL7rG4QnE3pb0ELJx0ttETSEKbY933nzQxMXD+
LwvfFGpcy8pYaJo9h71XI2+LIzMeiUv3aaisyMMu6Jqp/oX5/kuRdk4w94jkPRbvm7Uz4Lg8bF8D
467arFD82cWNXEI2tvrhh2pPQuLm+n8QHLrftJWoDNXQfQBDHW8bN9eGuNfuSOmN7Mhi7sMb55uN
nySwGzdlb6SL6PvdEIUBIVb2v3BnmxR0SLULerJKvjYPk0VNqtpP/VoS/HxRRaclOssvwK/lznuI
N3GGL22jtfNRVPpbEXa4LFuOWgsjoOjpLMyPS79ehgtFOvIUj7nRBEyTa5ednZYVQp8HH0naoNtn
AwRhS73xRS37oHcbwFSDaquNnu550QHnZC8Apzs/vXvg7ndcKQZP3isjmimxUYo/5K6icT9e4Fmj
SVG/jmbG3aBlUDZqkVF7bL3AhPVs7ZIyDxiZ3ZyrKdK/n6ORevVzE6XmQ6XAo5LS5VXiNLMYKawL
piy5VONGjYYNddjO1HJKBsrr0oMwlonqD/tCwyhWALgRHWJiIw4I2v6ly8wnRrsLafaQyhLg90Nv
XHmv5AuZQ4ESHC7cAx3/jhezaeILG0O95IB9yXqMLf6Qp2j3TL9LB3WUAvLyOa8D9WCYqrhVtBR3
hg413zWqLQI/fiY1Nre0aBsr31Ls5focDvHxuMjogHnfdmXs/kNG4958UZA0Dm4VaTGZBdfSZ7IE
BqFtcq73gy2DcggZT2BT2eOuqLIMUKf3JU5W2Np9mjKfOYjut4Te58uR7KA8Ea8zZAvGn9xh8xdz
E3wmHO0Ptor1wKdq589kIEXWIrqs8AuVCRcLpMbMbU5nhmIO3FKIabPBdt/8rQD3H6hxOzJV4u5G
URqE4+zVUx/DuuY6PXukRw2Ijz/N8oiDszxwCTMYRo/fDAe/tzgVdjYyn2W/ePgqQFMIQuiEv0w7
SvByCBLR9qNxE2976KH6SwY/1faDz/kD5wGwG52/zuinIB1xFlQzOkpcfQGk8OPEDHnWHVQok+7x
Gvcgk+hT6h5xerkOACLvvHvDLU5eMPWN3wPxpvrHac4WoWgvHsWOeoIA7f9/faCz8WIHYXl5RaCm
yOZMyxF0RReOGvh9tJw350Cm4hFMK/4iMcx5LYGJRHJlwKlLslDtzKEeQgdg/k7eBDI9EsFqmS5Q
P0qDtmine81SuHKu1uwlyp+KZ28gObNMtpBsCvO2eq5CmaJ4QLwOXLGU7Z2oBsAKZG9ti7Zqjdw1
ehoRDUQ0f+IednGnKQP17ZuCJuh5HckbwGN229z28G8BErbr2XMBQ5BMVWeHmBEJBD4Ip6BtHShI
eGgwcESaPT5MwUUcx5ixxaUlwOUUllm4Gs9dOGMXPJVVTLE1eo1s5yfpNpstW4ZpDvXr0o4JHfLl
WU9LoMFj9KFRw5hXhRUoSJezQ1mOE+XTYRK736UXaB+Qb+Xsa4ZG5wwdlNcjbYSNwl5OC/2Fn/mw
k1Hq9VQ4Qc6M7Pw/QD4Z5g2OUcV35zxTZi+dYu/NY9GBMNWJvTrHJChxTzy19WVr4UcfNFAsbGyU
OHrrxBFagzEazGR6tQ64o+GvnKaLfpY3Rsmve/jC1M61EUvjIEPChGw4QD2QbVLBJtqKiVCNdAp1
I/rieBundGiXfcZ3sVnZJb7KANagJx4qxDICuPjBZRvZKZu+EBRYBLgWPLThKrzX2A3sHOPSJmLT
sEXqrT8k7bUD6fsXrSI7wCqCHfOjKGLRMFwgXh5KE3uyKu5FdFhJeUuUYXOIhwT+6IT4WLM5alyJ
GCMNk5604NAF7w5sDBWjk37aLSxNG639MmF75noKvJl9u5eigBtaroqxVjZ7w/uL/kzvtYaj0+aL
8NHX69Fnh1Bjg05Vx8oN3PROxqSJ0/6sfbn4en1f/5N3zy5mOiE+ck0sQKcJPbIgaZyLRTfnOAxI
e0OIZImTbq+Saz3tl8B72ZRALd38zlEAttvhYOmjfUZ8Bh0avW7qpMgkdYq9Ii04Q2xgq9gsyYEL
a1n40PaNfBsctFocQoCKH8Dr4FmNwhk08EVJU4az2SwA7D8WvIxMB+qDtn4TzbzmSWHli8v1oDs2
8rrv3MXp8zW3RrrfW7vA7CRaIN4mLQgUoAahqj37ZefFYU6BnyVmXZAOP2wbcnvcSUqLaFimA9Dt
PQKlIOo+DAoS05x5HybEFLeiqqClFp9YUMaLAz4fI+x4FnpoWdoEgAPmOQ7RUclLxvbU3T/6f0Yc
sZC4TVQ1NbjJO9eSSW64XZbxfn14Zd/7Uy5UMvZC62V1cRIjy5mX5tl99eTO10jjHGe/TJb7xipJ
LkUCQqgxnDaCOJvmph/OYUzHPA6ffT9K6PykQg4BdbCqBycs32XA24v8bPmcKGZI6QRDl5QHM4+D
4kCMxeWVyc99HyisnF+iisTddmYMaW9cnnbb2mj3S2F3hU3OKyhFiD6q7DNWeqMfF9qmgNJzSuCs
xDk/iU4+X3thwa6ieUI+NjrnNTE2ry1tAQli787Q8fORIazU8Zslun/GEeTLI7lbrbQq+KORt6Kh
OahdCszmx5rtEbtfChYSgKi6HWu/jq596pG7+xV1h1YolmrCWULJkubeC5N9LTnN21kF/ZH2gPTP
QVTj0N5ksRMnyoAAMvkjudQY3Qz0NUupYBCku9IDcR30+wpzTPL3y3kqCe/8yapFuUY7JJkrl41k
jIl1Fn6vypgcgS24ha/p5drmgy4k6pvLwGm1gid7NQYth2bN28+C18DA2X5E97xWjfstMMMEW5QL
60mhMULbTta/o/HV22umtBhvIjaTMpyEVkbRIzuZa6q0w1r+1hTpVi0IwzAexkiUVbr98CrwcABh
J/sLHE015/RNAgimxDwnO7h2iTUzUKdgfUEo9KeZ2sqBHkR3gmJJTdY8pgrPlZlp5qjggHH5NZJB
2TO+prmB2Wx8MhR8feEwtIyJTzDfmCo0QlGWDfCSM2rNC6ZJoY2/WvZjYfwmOPCAQbReto3BhNfk
taDZkm22QtcRgnvqlYkMIG/xN5ORmudyK9SJw4PVLGSI9iFoppRDVZW9UU+GbQVuqhcpFb7e4zuY
IVwjWzTZHLHnrQD16DigVQdoJG38FoYlKBDcj5ZkPXeJjAUV6lWL1jaO22QkZO7O9LUQefaeFRuJ
/V0f/jUigRXP4UJZnn2f0zTOoZLMAcNxdKR9xpUrkHEQyHc655mNbnxsCPlwgin4d7A5K1KG+ec4
H0Hz50cxZn8R4zwilwC0EoIk31/oAh/UUWYpyjnotMPT8RYQJQznOOZatQ73HA93NGKvBHBfvFvE
Q6Nh2Qn97H+Zzvpfehv1xm+/SpFXh8j/8yFY29R6zZok/NOW7boGBm0sJtRPo+r0Gk/K2Q2zL6nv
0uPzg3RLYJHZq222QpoqRptVPlIJhRV9lFeMSr9pbyuky2UmW3NovPPQn9k60ZM4ljsIs3zSBAX5
JwdoLQAnfXaU0KfSXuwqauXzNYTwy0bzypVrUDWy0+4iBYufLOj+q+csDvmmEB0wxI6bTCQGHdds
iBvRAzQ9YPiAKXf6dmxU39HFG722ZqbDhNdDZjlVG2vFDHkQh1SVTwl3L8iXxjyHyJZMvaYeEBxH
VSh1aOsPHKtPcOvOVorv4HrLuUqllXB/gT6jdy5ZuuyLJOiJG26fHlHKwvKOdhKbhIUYrL7B1JSm
XVsOXYBS7QtDkABJhGOOC/nt/c2OroZ1yf09ll8kLXf3ojsfv9P3Fye11VERBlc6CgNVFfrkA4vS
jmsxpNp57RUvzr9yVHq+UcbluHaV6TTHaJInSQySHJWEcMt5W+jXFXP6l8zlBT8WChgP4RT+1oh2
f7SKTx9tCIHSJJBdY4gn63Lgzr10up731JL1OaOwqow0zLVIi54DH1aNOkfBLUPjbi5jj3PAhU5j
hsDhNL/mDcsljN4ki4eKrwMtYhTpGTFlt/YlNhSkWxf/uUTeplVM/2h9siHuFa+nnr7uFLdhfWOO
6pKgSPPQX3RaJgAmxyBoFBnNJlsomGq44/6/vAAAEuq3MNmDKAHwfxa8n9BCDnqwgSkd7cv7m6tJ
na8e8zTu7V/CZ420vzW0qYRxYjBr+GjOwH3joXhO3OkImmVG4WGkXBg9h3QWX95ekzYst8PP8qDn
3LqMfw3nUEWVGbCKQPZkbmlzZR2zPq93e47kVoAiKG4hAC8KLsVygIBJILTPVvmIPxWap7cqll40
FOe5gmsprZJ4wd7B4rwsZcWKMnAAib5YufEAt9yZV6D5WZfm+z5kBw/TmqOoBLg98ipYOdpYoZm5
2uG5RWx46TyeVrC8dsscU6N3inA0uEHV6D76NmnKR//r5Wnkfk+axyVTeZBMthtpXVPB+p8wzWB4
siqw1sIw9ceB94E5rK42dMG79sYqhDnuNhdaK8D4lwYXD44dmidcQro2aItuI37b+MVGG8D3yS4b
cO8tVP5ynSatPUMi4WzLDSMqbLlhvNXf5zDeGzqUTiPJJe8fP9Gk0swzfCtDy+EJpMDimRFhNUwQ
aegCFxjVYnnTVm9Lcle5WqB8jr3Za+eeb2dOyeRw3JR+YoDjZSTO7G1ltbQhU0RsCjs+I2FHcS3q
4G470CSakFjmaXtQ+r7Xx2SM7s2jbxrrPVEGjqkN4VjBjKywqBC10mey8Bf/RtiA0uQP4nIFE+rM
V8us4LqbSFfjM86PAwL1loNw+J1Z/YuwJaBfXl/feJkEL/Y07bcrhbcet5ez0vzhszSjtrPYppEN
rh5FVPpgfIO3JL/txwlXBBh4oPlvylh3ZDJ55e+nQaoYnYu6M50NkFe9aM72H2KnYnyfwiTo0VV7
T1mfCvBtjWCp0sgnIxpdJEe6CE9mmKkwgdss6SHSWWepBY7S+NthJewrF318E+s0PotEJ+Hl2gmG
CMma5uBvA617AHeeouEzngmIXfQuWtsjaLUTwVRBVI8ZgLCLLBHwVq4Nnrq/pqEVSuQTCuuAu6Wn
HyM/2QFuFbkFUhrKHonuMym4Ha98VG619YNEugU4fHiDIp7QNsFZy9MgJb9mRfEG7/S+SY4/OZsM
sSir7DA/g6uBY4pxGJbtK3rQqz/NgbxAkX8iDrLeqM6J3ivnQy5OtJNwn2RPLV7qHPUULuF3N1oa
vf/nDgN1vAW9NUrkBHRaZhRKB0cD4Wejl3czFxuGvjdDZhgNgHQzq1uzfbVRM2lK8o68rqrTlZGc
ZC7s2ejdUPrOrmg0jXw5/zrBk6DWtPdHBePpOz8MSCJk1jQg4vgG6g9ugh5fv/kmvCmRMJ8fhiJO
vjmXQ7pwca8+9YUL6mFyPQFFOwz4ULmAzhda2fYVac1W2/sj35AEZDrKX7T2MxxtmBozc1W264UQ
EX96u/e8sMDfvoWwL33eNQAM50CP0gyFRsxdmPlRxaAk6onOzYv8JUxCnh0/uQXwRyW0HBRBXcym
78s3odtdAgr+CqWiBftB4ntyvD/qY40AuH0OXjY49X3GJTJ7+fs5awUuPfaaLKuxKaiD4qZGkRCh
9CCxZNUcR875s2El/fAYFpV4R6Mi4zU3Uk1+0yXWT7/PC5ywwGh+22ozNhAaS4ThcvpbslgPq2Z3
+0ZCbFCGQehbknWN7ojiZtq36hKV9grzLsGOmuWPo/v1rnqdSAU/IZusrUCkWFrjDw8dBM+h96BD
gYFVOhYccsS7/5Vpjg32nNDO/BX76pjRD0QRsxuXV/Rsfo6XSDQUCfQFEaGxn+HC/ZmKG7brMP3H
Qqo+8kQvKI67+YTS5nf+J/yicfnaVu81ZxXXy4KNj24v4zWMIQ6yPGU9SyUE6kXo38iH9M/WZ62G
PjCkwh0poksyNbx+5fQyz8i9mo8zeHZeiR52Q4wf/p3CAwLNNi4/p5qpSv86nMguFT0fFOrLWEM1
INGC4yj4IB7DeEuCHGIBDqZObCJPxHoG7mbBcl834QCqXdYW6tJojlcMBw/dhhWFoQBwo+RH1BiS
1SObTYdeNty6LTCtzwhYb+mi5R8CiLM/Vg+KcZoTcdxX4xyIQ5kywSbPA5Uwo4uDwvtt3r7fmq2J
DF3wcY6rCOw48MsSuhmcYcwdOr5U5SAzsssew+cuuBApRTV8TyU591k9oeI3CcObaFDqspMrUEhF
Hj3EvZAP1r18UYVZHRRI2Qe32sagiFQFHawXufokMZcrii8B90eL78zV4T2Jh6eXSmbc2doVQIJF
UqF/0HYnDwWrfDnSPupBJiwo2/k1cP3mYhAImHusej0GwRECBCdmujw6JdBQj2nscm9oB9QpchWB
dq1ojZZ5VIxClriV8nIpdEansdXGnF6BpfAgjRMClznxe8epqxLsJHzONHfbVQsogjTisSGsGnsS
GiIs0Ro5LvMNXwTj4vMm4mEy7YsyakIHe/YyPp8SMnx/n6M4heTLQj8rP+N7jzwT2b2Jxle57xgU
1t7I1PtIOFuryZnpJ9wZOewGnH1nMXFwb7lbgOGHC3Z9MUmuU8pstU0DRgiPq84ixGscQ0twXKut
48HF9sRlkpU6tgnzP4nzy9B5NrCMaVRRXYJcsnFVTWBRf1pUnvPTgNv/dCe4UbUVJnR9XFsQi6gA
Ae0eM8xOIaHeZeYleMa9jKOg0hV+nDcLennwM80qzhCo8rPPFAVJZfanil4yE7XAdAWJZylDkWEN
IBrA3rxwcjdzBYsznu5FJGtcjeHzVZ1Fc9I1ikZUyQT8rvUPzjjof77f0A1aBzxAHUKJ4PK/gV/a
DBJJMI8LtscUXqA+hiBBOsiL8b+278h+ThBtRHyu8fetanD8v8RW/eCd0/9jOpKgE3n9/s6dGqeC
58BgX4u8CEYZsau/P4SY98mfmGNM7sRDQnJVxELrW7MoyR1FGwJ1HyHImBd0VDacu/yzkjwv3268
VisMltZYY8jEGIpXObdIdODtjbUMIXyj3dVlGfYMfoThDuLbnMWskllw+FSBIJDNyszqs6+/mA32
ejCpdEW54FHJQ71U428Jyh4+evZQOD+/X7YWWr+4BvV5at8wJsSUiq2O4bhtF1RcRWdF51L7JOE7
3nKHVBQPRIxwxY1sTk/DqOyJ68ZHnwcboeYBATq76hyoIXl8vMIjVytOlZrjueAuMLrtNiLbK4GB
MHeWbRQ8XJW5xxYlHkDR7DA9AKGnqKlo5crnVH/MY8SOXVzoYxQEg+fFCj09nGB3m3KPeJrY+O//
/GYOllQxmdNAFnyG1YsPOxc55ijBnBkif5Z2nUgo5zwEEiR+FE0h4YKZ4djjtytPuDdqJMP9dfma
Hwbx6BburV4v6Ee5yuteX/9etNvq4u6psHZDNzJr3wroxU9Nkb+4GneYkLxT1wdDGzhnvKpVfnTS
r5nQWfoDHWf7m7nHkM/3Lc+sftYsWKWRpX48B4ggdGKSLyH3wmNi187HcLxAlGWNQ+QxpXbGmLwk
1TqwvzqvWFiEMM2uI6J3Rhq17cOD/LabAgUA95gAUSC34ihqMYYa5PtkLwLbbzsbej4Z666NJoLc
m2H6lHBP/soJdArDAG8M0iit7TcPLi/WGW6hfBfkG3gbf+IY1gw6pSjYFG7IvK80Ganuy2X5jkRN
KVNgbsyxtOn1l3oKcc2vMICIh249nOjzox/vl96ikc/OBfKarq4MzqFPFD6JFvtEdLXdqQltxrZd
c1+Wb+f/lTkErjTqfvgQXfrr2UWRKnMMWpi8yjla1nN6+GOuc3FMOA1+tBOchXfpG0YZJTn3ekGk
yqd2mC4m7wUWpdbgTrqxDKxQi54Jva37ydBiw34g2I18duybDrX9M+9Mzap2awUA6nUrRZEmjkI9
Z1+ILF/pC+PmuoohfwrMZ0bAXVJdCzwtbbe8EuEfxecCCsa/Q8naYOOhAJ+7JKKPEcI/reuu1AHi
wk+Zw8nckttYARwE8IVgS9N9aHEn4ivBEz2pWcVF33TOS9u2mKHGDUL+/xuyv0JJaPqyy6G2ilEk
VUqIY9oIUfnFFJ3rd1VMaKK++SnOK9986FlkgKQQMqE2hKocsoOYFu8kCayGXY1kkxDZa6pTDPm1
7/0e5rWPCjT4qMFQr1/xohF94dIagW8A5kaR75PcstJ0GiEpSFglFn3cIuVK2oaOINfg4N5FgxUl
eVRJt1mCRpxFer944K7+q4fr7T+nx/ULQl5CBpM/GPUWM53GTXvZfGYDhj13Y+cV31muI10yWcxt
zZ9EFpU44treraqwLfg/mOIxg89Ez8fIPTE49BfiI7QP4dmXu4ryD1b87/rQXJ3O7xWZ+Pep07P6
YCTAVyxrhFJ1aBQO1ga9Uyvs+Bqb2ASSW9dOEbhuckL1Wnx9rkbGE0I1Nfqy9S9MwfAZBRwDWZDn
rBiShBxy7mh/zFyEqwk9HSg/2r5uIEcOD69bt+XblOIP4Jf/MaSkqLs+p1kolOFxE+XPgoih+X7W
kYv011do7nBHfx1HQVYPHdaoCe/MJNQR9d69oshoIyIzqgT91egV7IrRGD20Zb+/awVQqnVy+Rim
3VjH8pbW7Al7N7TGrevUcVTZz3rkP1zEuTHBCQ86T1S3lT84q9zTZvahqlF4/CcXc5f0lv9WyMeF
mgFK5ZA/WR2HGda26dHwsmK/ydUW3Of0aj5kAxpvOAS6GSz8zxpVaydkn7CURZGDLZKlavTkVGwu
ZIfWCF+vUocivQo9yFcYuA0hPKnTgkNTe4p+Fgh3wFukuB0fry/1TjhgPmxU6liiSICi5pBbOrJ4
gMk0A7dduqVrgF57sfrWROsF5P00gNejRMBmo91LlT60YRHZQI3aJ38MpzAkR3VuV04UnYbmZR8e
l595TGj01gga8jg3CUfx+rmrn1evunE5W38qd4/CyehtIWTddafP1ZTwES0Zm6t049m7R3KDf+li
kGfv63A4dBdjzr024SPnNiLh4Y4yz2yGkkbTKVAen154cdgK+5X5bRFGjcI9QMCzUVxkMTIM1SKD
2gH0kHzbLIY2lzG71czpbzpWJ+nl35LhFEyASL2NV9/l7q7FRM6Pf7CE7ovm+4GkZKGXieD2+9cj
5TWh4Lkjqr6cpWg7uLdaUqMIcineC2qAMhKy1WhSXPgT+93fyJWd5uFUH0agsWwfvWOfO+Pafm2J
FkaYVOntSnaoi2RILOccPp5SSplbTDzNdwQuoNQYFjxjrHjgFKNlEu3mOPTayBOjbsy6kmbrJxgg
9lRC0mcOmYuRp1EeIhOkSwmHD+Gj6oYt6+D3L+kcPnZtWL4/wjyGi0KRv+1uOwM1sx9wRjSieJll
x2hktloAj4cccliimC3g27BlorcO+JW/UVEYRdb34Z9v9nL/ZTP0Dj1yhhr6rJbbXVHWK4jM3VvN
uF79F0/TPqmmb9jpmKzQugtjA3MhOeAI4I6+hSn+w1FTke58Xa5vCnSbVcWPZNandLiKyVqP+ipz
vg7In2REQ9vSzbw2U51kNfd1Nh+hXdE6MTqz7IXuGWZa/OGVoxjFE8z/27/sDet9tY9iekcCWhgH
GZyxAXd+2jJmnS3kZQKPROBqzxz9TSHWZ4ZuuMjDWFCr1Cgmol1Vie/yhMBPwWjNMxHN1GDApm51
5VKjoVf5u6TyBZS2TSUPZGkH3Ar7AEbfCQlZX3wd7ms4VWr07gXzeeRDEN62TGdxtbMya4dsVICg
5HsNnMZ1O8svkupBMycsm2imcgTlDnFQkIjx9k2l54jr87f2mv3JZz/u+J9w6DqMLvyMoVIqbZUx
TphTZEWSYgvio/8u49EL74EWBeF1OYFlUqwHT2t/FTpHL/467x3/Jbd0qDtq2cnQBex4llRxAORQ
n8pGVThhcqGkD3GpkLGOGNSgHiQSvX9DLEyH64aDMSKAAPNyrOIevW8l8BCyaJA35V055/M0eJfT
kudz/FT4PubSA2U47jngWqBLbmvT8sxautkP00kkukwT4iE+XE0vhHRVJxnWTM69bRUWW5x9Lnih
Ug+ckvg2TG5E+v7qB6DlHDU+kH8siXpFSzBgneAsZ63Cy3DDLak1sQ3HcNlJl03GpoAU4IQ1H+rS
YVhGUKswwW81MO8+eHqUXiRrOi8pRJRCZHdom5QG1itAidxg+5oqnzWXGXPeyCihKuBKaNgwImjK
OkVUEYQb2Uz4o1jNeJ1nQeMlK2cmaxww0nRRVBqOPf1aUBFnkItlA73/6LrI/daXabXeR71p6p8X
3msaJnfs/4YjIKD65HFLjHSfuECFyychtMi2Vy3Ce4oDfCedMIPoMxmvwI0zttnN5TJsLDnmQmPk
gL71AZskXXhouQngIaW10/Kj85dfjzOOoqrp7j2PMuCEG74m6pM29Uk/NvHvOmmMX38wuA3T/vGD
/wTV2x/4Z/MWXmf87jI81KxYU+b2wCbXu9kMCiDJ5R3ksR7qkJK3cxHC1+Nl0Sn1//bsVxyQpUbr
McM40Y2DzcxSsH9gxWFF6npQlUldb9NLVAwEp1NW0pZfkybEXeWtzNpDQrga5AY2lSUh4Dq3BC9e
30gDcm+9/Uhz33SzNHHIoGTiWYJNWojhh1QB7WmG6Q3UHhR/R3O8PLAe5ANCoI48nDvGaDqKZlqj
8zwlSVkNzKNT/QMt33xJHeAyPZTgWqG3s/Pku6LlR75n1Fsq7qdphKbDitN6Ka6nauyM0FLywGVQ
gsqPId9gKNYEfEJeYRXgd6hORbryUvHNdaNK9T1TfpXbhj2W4iuGlU2xc9wYvv8IYpz7DiaNGWgX
w7BNalyTyW3Qb720HIJZZLe70ngunZIAl5eEVYDnLlc8qJ1di4xYg4UFvXjbLaA9zUJxk8tWsTV5
KELzLgpcudu9xmZg3x8VUd7ayee8EI9P60LxaPkBPVM5CGW9SB+6A8I0IuOSZ5w9wR0iydenrhI4
awDdD66Ctq2Yj2VALlXMH8TRkDfqW+g1jgzBVjMgGLAK5XwemGUQ2QBDGAR81x+q+nJJzOTUXxiI
d4C+Xhlu93w3SoYHI6bswV/G9pDd5mhF6V/jxmcbePDoV/KXPPZwZxto2ejc1uPrRfDqrc3lXQ5V
4HbteAeI8fia9DvrBov81+v7DiTF97MyqZPHeyObOjrvDwqZVrQKdGimFRUiSQV74d2LKoXfpR6/
x/ZzGuRU9FaVHfSvhxLv384Sc0yxiV4tUq/CFFwdbABQ8t2hjKrQo7QlrguDaKlAMxKFkhYPdkTH
XPP3cD/dIOJwEQyTaVXdTQFQ5P9I8PpDbZjoHysWR+vSSlSx58oDz/dAXb4G9PGJgWRGw25xvirj
ZQCB/BQo+InXx20sFocOSkwJ3Sr6HgX98bJ5LsRizVRuvbV9xn1Oc5VPVR27x7IB/x5Lic9v0/V5
h8XZF3KPRa526y7vkxGdupZMaB3zwR4Axszhk/2bEwtREd/hfRjPgFm9RFejtHvBiPC14iygvytD
cDsT5TrCVEl6gQCqS7v2gD4C6ptJ08WDPDi4jO5UM1zfMCpAl3XIwVgCpyEn5JPZPbozGlUOAqYY
jHKc4Fvhsl5/xqvIcR++JGh8cXFhDvBbuSfc/4eith1GfgoJS/cms7vn0X32hSYJivWggcYS2ao6
Lz4ocKPqbWKX85oWSCjmg55JpzT42WnfZ5QuMFlm9LedJOLZWdCXjzVPTO3oiU3eF5EisU0ck7o3
JzNMkaks2bxDObtJ/Sey8qxWzEaRWiISFi3dGVBNZymeero3u4zTp9kou2NoZGdai/sYAdlzz2/0
+x8IQF/NBchR93Eq9ImDdYNDVI4gnxd7ofyRDfoifVNvj8Jla1JxRms2POdSaHVBSsQE6hGX8LnC
xlNmF0fYJdvRvghP1tYQnsGBJurh5DNQF4caAhYlFm4LnFSpohX0ZV7CfmvFp7saERIvKkCmrY/V
/aKxHFpIsM57BF1eQVlXedG0nsvNNlszy4Z5bn/eD6wc9RcubJoB5sWkzrMle4INSvKZdOF6M5fS
7labDxPFrMu9YpDdjaVfuj9M96aHlG32utUJFdgxQ80CesupDp5xeqCaY12zWy2UGQHKUOaofrdG
D/BkNwv6m16tXo+dZMocdMVz1YhOfHA17EMBRayjoX5CgUpEkuoD47X8hw9qWN65XOcrMsRMqKx5
OpbL5ovvQLC7lOPBecVoP3oEXzXFm3S9BPiHsxuBZWaogq9vYyqsC4JP2yz6ZFGWDZC8ZBb4evQi
Qbs7YmkxC8n9sC44jo4ca6Vj+jQidW5y51Y/c7avrUyYJX88tpZbxj7vzsw63aoUT2TCxrYaC558
v3uYPkTDuv7jaTB29aVtHtJee3WBdvTXnyVkzJVK7K25tEjQR/7I6DcSty8NWGUZLF75vQ0meeUt
52ghJKrTiWamG0EPQzAnvux7PUrMADiWjOc1XEeIg9MXJ8zPBCeqf7BVl5/d8WIvqx/qdn1qaKiL
5VxC+c4Ndd9RCXOE05E6GasL+FyyF+4VpTBPrKOLkKNlRc9lF8MASTqhx8pwMvO5OlPXVb4BwM+d
cnQeN/HcqceHxn0ivmD2bo78zBRrBKMf1w97H0qPYO2qxbXFadgQhSC8M9KlSO2QIfqTkow6E9IO
ey4J4EzTYCRwLym5Ojt0wDJd00FBLW7rX/a1j8dUhs/wQN7EnVFcRdty3ZPMK/etSakJmq7gwjZD
deLd7pqmq567jvITTBR8AOLLsbgO4B/BQyn0xRpDJCb8bb6o8KVCjX5Sz62EQ+aNqUqpz55Lqjq1
QAjNgTde1/Z3ilm78bh5Kw/BARmB4PCo3HswRVENlzRDz6R7jeei7av01nq4oDkW2b4+jS/c2B+g
6EFiwVH+ZfTxtPi7Z0AhRUQtsN/q6O6+2ur941+XQzYzfBvbvATsmi/b0G2nPfcDiwe9dTY85Xz+
84xCPiSyQgPq9XGeLHl9+l3oXlxpA8zwekXQU1ZT+Gq0VTyMV9cuh5D3dnAtp41QeUMZB35bh1pu
40Fe6iSm78TK2Q1qzU11AZcs5oYJIy6rcstZjqGXUOFwacFMs1zvNfxIukE0aUj+WhVrdlWvOlWV
INnPATooWR8DGstll04hkU0dP0VTWpNiEenZnKqdyNvvX8rVXod0aZbxe4/jX+X+33on8ospgLAg
0b9bdwgLCqZ9FXEB2sPScCDx5no1pP1aoMy2NnmxURFaoRz8Q/nunkD7tQW62SArEny3g4ymKc6F
IH6jlQIWrHNaXhb/ptobYUEmoBRCsl6HfwfFqgJJNL3KUF5+s6D59jUE2tWwzqAe8r2OcsfZEDqS
oYuxfR26KtDqgisWVTtNr8eC0RaWJmNoa6MO6VrFuIA1k0b5NBHDQfQIP1D6EOQjPVooBQ6chI8A
s5xXZI0OBYhoI3TCQymrh/X/FS42Du3T8hglECoBCf1oHMAKCbJom3DTejuXYE2ag0Es8q3RwTbk
oYWAzQdQNa1Rc0SR05I0hlwytXFhZnSifKZcVAp17sn/bnl4k9WOeCvoXe41ccJx4MX0QZ92eAFK
WoXkHaTd2iX/CN+Z70ymW6+irlrN5ylUPWkXprDEVGkiPNUQPS89LLYUTrGLmUnJnYjWep/LtDFr
AUxkW9rPsMJnGDAMfbZEPfU8v/WrSVi9/JvDILgDgSUlP4+1iDr4ousIn93DVuhAk6HhrkbXsqK4
ygKQuVsqgV8quRZQcMrbwl29i83SQZeTrtZ4z7VcCXm+csGJBpfuCoKy/qzD2egbyEimi8gMihje
IxBwXnt1oKudjn83B7o0LErNOZQ3obK6kSC6A6HSRgKfM5tcobhr6MO3PddZExzJbrtkOHwrYnWC
hauEzhTb/tN0PLdnnFJiSLHT7hiTnUZvX5QNc+zWXC5UouxLziMc7OmDq1uA8nGHl6T8rtjBZQS8
OpmqUKdq0cHXnjjvAzg/fZqE3DJF6nZiDO0fgn1gZR2BI5LsgKOUZTYC+ao6RNpGHFhkqWj4Pkkw
SOalF4aewLBjOPoctmTHdh4RDGbQ7j8/qh+TnZVtUa6a9KzhYY7/DG7UE/DeGpLNnIcRrqUGv3tJ
cno4X/8m9mZDvMZzJY6s78lBvnnKuBQefIbADUYVH4tYdCFukFHAWb4Uhw7J7mzcbkGGKvofvUG+
YvRkwMwWV9oST8HbhRipggGd6VFSa6MFhkkdYae7kReRyZgRf/hYlDpmb3LaXlIg3EhxHcbWT4az
4Ap+T2GBzDFNkuadi0wlrshSaLhYDV7DKaNAWJK6VN2EKIm85Jfn47eKhWpvWiGWz/xqvXFSPBeY
9wQXi5u//8oUWKqP/2hUpGdzEYtbK5TL7RHl+whABBgPlZH3hrq2bHN58pL0GDHxpCwc6UUjE1N2
NdI3/CjumeKP6oze7yjldSye3C2nqVcZ8jGK0w0JeaoTldABy+i1tOrZrf5XToiLqRFQaRxyFYTb
xLt0k15bBV80S2jkZv7nlZIbtcE0X4qpsvWYh54Zm1rNE29gU4TFEJwCKrmzs/+hM2jv8u8ylx0N
80I9wZqsQ7D+aDDr74Qscag+FAUr9fOxKIuqSD+Zk0nesUMxvC4gw2TyM/BtfTREOYBgDAghHkQb
1qV2bK7s+PXjaS1gxX2wNGTapMzoLWUWo0+0SaJ12g4Gg3Vlb3uNKX6Ke5ARFTJp/H8t02jf6lcX
ARiWF9cOTLJqzvt0eWqSnUAd5xeFQ0FZE/XTufAufyDq+D9EG5yye4+22EiTyZuq9VojdbMYK0xq
NOQIcfT/S3Bwu70VSq+UqXvi6SUDsbMdjn5uzdP6KmJRGy8PWjvRjY6mDNIMgTJhHn/uonX8RJJU
+Bm9lx2w8X+faX05Ke5dAwXJHYYfZEhHjPNTMAVyv5L7ux1dJa4uasgQnIY4zZoGbc9tV7CI+3fe
smHBrKJpoJZ+17+q02wTiT2AxKuNIeqJx5ZTNT80misuabFVlZRiVM2zYtlf2m5JmMKVT7Jc85eN
Z/znc+7J1d1rwmMLT5sUjsNE00AHJw9pmm/ejpjWqFnAHnZWuNV+tB2LX3RWvKHu64kU+L2/r39I
lIdWwc+DZdc1TzI8pauqJPZ4xFM2RMD9BPTBgNZxgiz4MEVdFsqrrNagkC2juACKWalyXGg/QTQY
VNAHsV1LxHdQO1OLbTlNy9XCZhtRjGtGb5kRG9rb94Rkr874Jh9QWEcukRwnWGsrMp955WJplz6l
9+cxt/XZp7G+qHbJ9CKrikJPiQYcV5umzu0OMs7IQ1mi6pG+qFiDOVYw5yiCcxkQvHZYEiR2DNfO
zjoTkwiytnfS58gPYwycS3HzEAN5xIFGf+nEdHTgJIqfgShzwBHvlUFYDodZprYFWoQGA8i0yVaA
eaf9K+Br+c7wGRHo8Oas/frdaBhiembfwHLpVGyASLzqIxQ+Cl2cCWHyiDQI0dDqlW/+rYwVTqkp
nuKbrPuBuO4y9mR0QkI14IsG5LWaPoSNbmrH8CjQtXQiscw7CahCVpF5sD0kACQKumWZ70vGuc82
QkA2UA7izL/s2tbkdpLop3qdh9rBUqXbXUcFiBQ+1XS9H57OtRA6cHyB7uUocIu+UbJ28HnunG9Q
2xENO01OMIprgTLEeqHnqHu1ph9BzcGZHwDn0xuB/S+kAZ7A+x7LrVs8PhQ0cexfqfNn+1Rvmria
rvyfWem6v4GyNVAuXh6l2BUAz6hOk1Vj8D+mfCKr124vAIMqaNyqUM25iqtbOU55ZzGlMgtKfTU3
xZ2PyFG3uTh9kBoNGYpA1ulmRxBE2CqbRgacmxcxtECx1ZOI/nnKQexqbYzgpzfKeQAaF0w33Ylk
vTY5Xrmv4rvwn+mKvpcbWgKkrWkbf7hEmPKD583rnVp62UkBlFBwDZdxSofG8p1t1bl7WfvMYd/C
0dS+6GrmchfhbnFchGvLe3oO/kF6Qz/1+J98G+yBWztQ1wBUmYReSYc03q0nTIGGzr3ifGCOCIGd
JJDX6UQ/bQ/SfGnOlvBE4t0UHrilWKMkAeReli5ocXhfzXvSrwnOgTd7k6CBtzP5mW51gALfJSsB
+xCPL1IM9blYfpFUKBzihkFwSrz1ET69XLIV9becXoGrbMWThcxU6LqCPbuoGn/pOEJmlFQ5FYUh
BTGNyc+IR09CzbhFobo5mAWVP74uqA9S+8VULchMdKGhmUJ2uea4eUIbvgfT/Bxbmv6zhQUBXYhQ
5ShRqcXFyKPOUqR4ALuIQEjG5aSBwnxl70GJYiaeKvKeYHBd/U/I+gjGPC5E+NP4VQR9dFzeON8S
toaT9wrRcCoAxZJ4QNWLRNr1yZlKVAz/rOSgFpZPQl1A2rROKcsArYmso0U994kTJ2VnflEDiZma
tZRTieC7rIXIo+73bupK6bxCufbwH8iVFtNI3c7ArefatME4YRYR3QlKelbbKqTssoMVXX4wAuB5
chU1CN2eohBgFhSh/teuJpSeQvHxFG5djbnP67s9njyxuBkrtSls8KjQm3dCN9Mx09mShtXnrIs4
/ZeF1leBWQngggq4SxuyqP1A0fICwKj2Q5kQmqVG95c5lYCsSEQtXXARLYAFbsnYl97NHqhYx44D
pESXs4uTMpXwcyq+SQ/gptwKYlS/Zvu/+pP7BdR+40Zv14fzGQDhYUV0chIckvlav071/25QJqMy
1ZUq8uIReRPk3hE3BsOOvaSFSWS9iN5b7oA1ZbD6t8a0GCo7p5i+vIu7noCa4AdknzhKbBuC1fR3
N7s1wS/qxkECa3VwNKSEbp5lyunJsJKQjRc2Bhkb1M+KoJ56VHEgcoz9V9qu1WSMhw+SEL2o2YZx
5btad5/+ka5mhtekKv4HySeyq/9i655KtAF4887/22LEIcTOuFoZwIWufhkzZWb4QVcL+MvUsJUU
5lexQr59rlzVCwaEObiYUaVZD0KFr0/v74XRj+MXhbVKaGjsfhWbySR+U8vvj5XcOU0cRsYX+/uZ
XQoFh7dMQTLwFX1Zey5ULAU7lB7I8Eg0z5rUpzKezQwOmzd0ZbPudTZToteoZ8vDxzoHOSXeblVp
BfGKkWAGGIulLPUAxIykyE29IylNXHecJaJdIKKtXN4JFZPs07zbVd1AdEQs4L+0dVf9c0jKvYHu
5AZlmQV5soV/uDaKuGAc4vpXnjyGuwjiy7R7V24nGeCpb6owKHvxF81QjeX7Qh4/Uo1i30CPFpXt
pTQ+pkgIKnyCUNwOAOPwH1EaqjjNGDRsBeVeD7OnsHM6FKDpUoNsYHihnZ+nFr4QLV3DsIW5+Oe6
Av2FBvfr1Fa/6eNo5YTsDEClseQOTUmMij4/yjMZnKth+JPj0arsk8xxUMSjxxzmPMLpVryjos1v
QN5QH7rqyMHulrvHRuT4Dp8NtcLXXB8a+v4ioqHFmiOg7EIz6cxL0U7TiUh7ZUgqpuL+QHZVyFuC
bb1AVLCY0ZVysoIMUt9DTqv/4w9BhgVg1KC+qijHKWLmegMKAGPWqioDZL2QJ1FX2hHMjesWQLQx
3moFlO5Wyk8v6z12fYhjd54w+4b9Eg/ABJ6cd2SObIsjkNBL9QFd2U2rW/cb+evBcaSsDoShO5Vk
iPnSDOPuxy8LKFNbaXjqM5Dx0xAn98JxPjlvTwkr+EKQgkdiWMQkKoqJh2ESaZM+LBjK5QhCDA06
yTbDX2UbK7ZeTONSXEm/YTkLJFXG06J7dU4arYOh8MO0q1ChmDKaVmYDhmkofZDGMbb+kkLrB/cb
tS6jNMT48Hzk1Ti+2ZLXMlX52UlMn/3tPNhQGRf88t6CNcL0692LNOupdUUVkFiSfJf2gF+sTkv3
SMv8qXAV5RVpQhP4iTnsLEA2lONRoI00wqZDU9bF967Oho0m3aK+cBJFQz0174DhJRp7XYn7GK+8
5hHbi/6OcQ8MsamDxqPSJ0qgnSZOuLpQQSwF0VsJmOjTQ2OiTVeU/HXqRASVNPwMA3KcejUmxqyi
bkUJurgzjmNtXjY3b58lnxKZiHqtwvmk0gihDBD2fbPIEMlWwK3OWTqmPk/q4u3GJlRNPqLhhAc0
RRdlyvoUyEXLRR37pTjqVEQ1P1KuH1wKeZrDQW4xTgtdg4Uu15/xXCxFDtuwDY0JyTNQuf6akSkn
TgW1+IGCwNUCDc8avdptHJW5FQ79bWJfWrVlqd2mDU0WFx/D/SXv2LWbwHsfS7jxSWsx7LCfGfXH
lGUpmV9Dn3mBUPxwxVZ8tt2efCvcgeKgLvPJQV3iZKcwuYUfZdkB+gmDvKnZ6VDLnbR2m39AS6HF
CrtXzYo+gV/f91SA+RK9JOfQGn/xL1Ao6HtslVg6/bRG/KS0oNR8BfCGpaAuo765+5+kTGkv6XAv
1CAJDfXwsYj9Vy1XKTuHoQzdAiUkaBDKmenK8LiUe8+b7EO66SUgRl/1s27CXtOr/93+cqBN1GfZ
N0n8DKmum5uX4Z0x6gYQEFQTI7PVLhdBIdSX2oxNwGjSjYp0p5VqWUc97X5/z09yx4rg+D1aouHT
S2dOTTt9TE3nUYQS4R7zmjjuQEe3F49lUXHobJ+XpPxWBicFSNkeU/13tkKitNsPJVVOcZm9TT1R
ajbfYm5tUAsxKLteHdGx98YL1oB+GdDezNZRJdyOklByGl1iM3RviiEnPEvQOjQoPrEACt4hM8ee
Vpqe7+vQfRBxmOjTXAmLRbgfQi4huZAAUUdEnBW2JOOqzt9azF18rMtrJn+j6bsrH5aLYIPB/hcW
ICIehU6Kjk+QABRKoAUM8Lw3kSrXsFfF8hVzaQB7OY99o0gFIcfPmO6h8Q9vScMbD034znLZE5C7
FlGm6yrjKk+9/Z22ZogiTo5upL6aNu2EPYeI3Q3aRKe1CF9Xo0SCvbj+rh9Wz1DH0fASNL17TqwG
MVwi/IwNYTk/4iXotfqcDg4LpyyUS+PM9r6owBZyGfS73ZskWEpmQjoIs9QaAYfJXuQB0Rv5eNf1
NBu54PcnhidsfAsC8JPpASvf8phSx7WlVZlANkbYsAxpWYdlikCh0iJBs0t7sNwic6yfQOaJSXF5
uBDgT/AFZWg89ngnTwIX/JL0DFStOsyc8coFcR5MHBFyao44U0rATZH8lmbnPbGZbVGAUxaUOlWN
UyfDmPW2M7ntCru7AKK3rSvCWSUPEAV8ctEBrFde+QZ0orQqHaQYneTWZ9KdE2M9tF55rXo1NIdw
y+edqF3/G9+LwNioFgcHpzoIlVmJZzgGiBNpgrIsPTPTm/9TJEld/b4+8fL+BDZolVn9DGmxt+BA
NCeSVK15zJYg/kpm1Bp8DyovNDabdPpwEq8KXoLgFZwdy5H0EAbDgfdu2XZl5eAJyoN/gigafWCQ
nYYvEJE380RfsuGpPtf3X6tai4UeIdT/5mtJ57MLWvWz9p7m3/9+DERE0oIyKTCmE1O988OI8wRg
soi4FeQiovKpRs8f/+XijSIdczkXfNNxS/fkeqq9lGxA004oMZEFPfXkB4nTRaCekBave99abK84
zgNU4AHv6meCnyNtD9/FqmI5lil0tDgADofIKpNqeBwB/E4L1/ooHxmohtiVRYqlhAZ6kxKoZ4D7
Rzn50GmHDul/y8WO/E1NesqW4/cxMTa3J1TeJ7CFB0SElgST/trRdXcXjrWeaCnEWDMpJ1XxJaYL
qKU7IQ0vhuPS2KgFgR++Jk6Eym+UteD2mrihgeitZENkgH+rpazza/ESdOP/HNbiYLmSpjpQU1Je
GxIW8XwNW+V98seGbcSLQxaxo9hZvO54tBkRTb+uIv08HI6brFzbFFnHT70ypJ9UqxmOolQVoloB
AahAe2L+MgeQee7W/puwNMhMM+8M9g3dWb3/cEiT4rQvr48i62H5+JFQ3ttRk8vu1A0LlQbGbjz3
//iTKo9VDsXpYIYlNurgVZ1OqJRPtRiQBZ+0vpA7iVroO0LMui8lwu3DC8XjAK7NmXEDJRgKQm1+
q3j/R5OdLmS7D9SvkogHan63R5nP0D+kGTRZonXjdmNE/Wigualy7jaQoeU93BKmdhs4UG+8pCBO
Ozidh1StIy9ly8n8MgJ6MqpJLF6LdKXZNpTgR20dNoB9UFG2C+SIrLP1yU1y4bnSvstaHHemTl8C
0xStljU9XXWHBd0kSnJfhqSxWLuwRUb+MIAL26sD5tMOkpIm5i7ptaPcaXs+fgZHpyItf+wKG5oL
I7qsLD36fhqN82/U0dFMtR4annzb3jh5z6ThME/HziPxPLhNc7vP+eZt8D4uRIxx1hXMzZZ5cW1N
UtjIfVh0R3dOJ7w2t7Q0NIFdJIABjMg8RwMWHYg4qT9KvcDBqrjqY0C5d0ABoaltsdQkIurEMfSY
phpp3KlJkRzhJpvga3y0TAmyqWeYuvzVH82jaiBrPnJeAAIKVzyczk4sgT4ZAuk2AKFl8rEPoaGi
JA97l2o9UZtLKDgZjKjMrCJIyHf+ZiCISpXqqDzL3nCWX6Mg5rID0gjk9mHa/HH7e1BVyePj5BYe
ii/FxhjWAaN2RFh5LP7aq7D4QSvSfrRM9H8j5U/2amoinWYOZoWF2xGqfiyXRIfisCidGWy7HUxn
+AsqtPuQxiY/0H2FLQIociC/N/VYOIS0JZFMtNoX8Vj2Gj9/Owuz+8o6Ky0RuH3Ig/YGDoU0tOA0
3beDkaeoGNA9XiZOdvnz9s0i+453DN1jqhTDL0XE/ZRTzSCL1BxV6HrIuWqdz7DqL2D62unDeiQz
LDsVhymHb75/76rASC837ap0/t/omXwupRBlVvUXrHP5vFr7/Qv3QXfDeKltiBfQupZP8jWGUnPj
iltZF19VpaSGnGHz1YEfbUV1+1M+os0LbGe85Pdn5gOvpDCBlNMflDPaTbEZNDXsAsxhkaDwrJkn
YD7h2wrqcQaDAwTpDHL4GdqS/R4CflNCQWuM9vi3VLaJWlpyzlioJtYbXcHhh+TJwsoH/WOGIk19
vBpajNuZxnaROdBPrKDslBaxnNO+Dv5ZyyAbubb7ZprQgNshODcKLrAJKjCMv93zUW+Wq+mkUIvw
/+7jihAKgrgn8wuv7+TceL14z56uYSB2iXb+XpV9upgEAay3eJufQO8syiZ4b1G9LNSHpj11bUv9
WVhYM2p6cMBwEjj5xS9jRa+4i6FzFhVA4dP9KbVRwLvv6cqRA2iMHb3zZSlB70JxgEjRS+ihWL5M
crKPzt7EGu/e4Mx4dPNtBoJHNnvuNjmEIxn5jGnQCaGYIFkdVxGdyhHQ6Pk3C7ZewYmlTz0YUuiN
b//UAmmDidKKoByPE4CPVG/atYdFYyrH2UXZ/wXIciMEjCRNzKhqNyFfSud7K4xU6b1iLfRbOyQq
+Ta+4dy1FgGjD+P8BuVN5H7C7BM1J/WmxHxywQGVCQqT02OhBncW8NIVmk1rC/DNYjB7B4Wn/LxX
X+HSlFQnWOYDBkkZDyX9xXochETXsykmo3b8P7PY6NX4iO/961VMYOCLyL4rWucsLWYcciTMoHLi
4pxTHSFSaEiw+NZXmAu9CWoEcllMuSxeax5s4+VZO9VgaKr0AwqKQdtKEPtqQZq1bHc7Zaoc9KYP
4K2CMhnaUq4cNx9lZXXBAk6kMwLiWolxFG3o4/1cJiwfZC+WpuLpb/etKhMB/yXiWH8699D2tgYQ
mSNabXPeDSAc9zy6y4M3Vy1hd5dTLdLo2Gm+VMCLjbMc3xomArMS4l7YJ8FlemPB+pM4F8A9mbny
3rQxkYXk/LQCDeAyRqQqtV1YUpMsgzuPz4TFqENM0kGNYEQE05bORBQHOnvcBLm5npT+7DtUnnmV
CviPqUsN++SE51Hb5MOHIQ47HXLMhZM4I7dO1yIOFHJhFcTv78sHrEGjN9feXJg33Oc91qXTYSqz
a8PHk+qSdnlr5ppLTkSYs8xiRyqV7KunyqEuzJLa+MtOUFCSDa3wK0PSHf4CS9n/ArLjespVWl1O
bqPYfztsLRRqk1ng9WC+nlhHz+Nqsq857ZtNVCSVQ9O1zioHKoZCQcqnW/hTFijbsfV9Fwm9h/m5
h+p4Km4wsEDUT8moVWz8I/SaTMowXE3LQVuB4abomXSQ1kWbrNYRr2z0gApjYJ5mvzdpc6lZYAfq
QhUUtNvBkHOG+z+oPrFGpIgoqm/BuOMVjAnDy5cRrKSbc5jFIQsQ8NyLBTMD3s5bMVjP+5r9gXlW
6iVTYPejTXrmGT9mQeaSkuyeM263Iwya3kUhpDt4bTWKBBRvfckxSTDlx+gqgeaMTtVLnRmHUViF
bvJ145FbzURT1vuPFGry9G64KIGRZwaGirosne2jksnkUbf+WzmLofYKU9mP3OWgElYoCmFDXagy
/juwUrykjnv7VcYoRDmYmTBY01G2T2NZNNeVfN9fHobYge/0BCqwf4MNYYy6Zi9VkDRe+ggKPEpe
1qOaUzqZLxo/kOSDHgjon4DAFJvil30mI+k/Is7JUg8BYwULgxIe5dYBtBa4Y7qHRxew/SOo06YJ
dEn4V0qqI4xzjiiINyXoePLHp23/d5rx48OxSjur37acQrd/AJvFU9v99U2H7PSZgBSgd6LUOCP0
DYq/JBjbe6cri04+G1SvRp0Bj8CXkt6+cjOluTz9r3BKEJQr/2J4nMnuTtDd0jJxQtXKPITABECl
j37h7qp0gRKYLxGIqnqcdG+6TO0/8gFcOKe6kyaOn6E9Zp2g/ifiWoW9JZ9uJv/LDUGya7Ui+CG8
BmX/SJyRZD9/5loZtWZuS4xU+VHX8LbJpZXsa0nLrlg8MkRqxaeMzUCm2GmInBbhvnvg/1g+GySn
UaBgyjun5tJY8Ht4rkrDj/Sn8aEG+q59ld/A1LSgTbwmWTNxgBURT4sqrYGX0VQK6VtTgu0v64zU
PscaHHuQfFba8vGzzrGVtwkUnGH8LATfQFz8XT6rZExcn2o8aEDtdUENhjfaXoudQXfe1c2/7xkN
r7HDY6Q9rPwvdPdnsbhUlhKdbn/eWf8vIEW+Vo+LsNrojnbZC+5IeDJh6FeTyzSldR2L8YAWbcpC
Px7msB7+9o5FUS/UtEURML9GB/TxGjvbxzfUz0Sb1BcPObVmhdXFWAi35M0R703OiZzVH5Le0O4g
z+t0uuHTJpTOp0n7kdR04MIcA2EbZ+0VeNDPt6Xm1CVZIj/mhgZe+pWDwTWh+3YdkcEBA7y1pIMd
TtNwnta7HUI6e7GkFBdyJa9V/3gwYc4iEt7E5y2vTjdaM9+olTNg4sL/FX4j8/SldeudNnaGICGr
FbGFWM7SxHKj8bnAVcIRottEphHDSArP71dnDgw2r01seY8hSl9a/mS9ahlP6OFc3bSI0+yg0nGr
pVrRDahDY8EhrUObjIFhQWAFsQBCn5Tpu+RRtuUBJ0FKrqM9n1nCB/h0ZBhvbfG5kYHDDaLPGQu5
ErmXK+iazwVht6zHir6wfvV9n7eHmK9RjAXTLlSJcgQAVmn9/H/2McvHiK8+nny+gm3DxmvtMAG/
I9G9sHA1DYGSJoyn8aDRcgauEJRNK38PUEIGhYH8HkNimi5gZXKyT5CFmsNiYURSJJeYtOFWZYKz
6LLpV1qrWTARkZtEa3+l/NbN26OPI6o1GZ/ZL0ea1LtRcaRG2syfP/IqNdJ7/Hzvv/nclzyGz+z3
40wSnVWZjExEWHV0MXBIGBHWXZqiJ8y+69Uc0FnIIJosBNLVUFKPHra3AxZogCVS/0Mo3+hPGXtE
oPjfZSnW3YooLaWS9p1IIZG3BHD/fDQ1tugdEE1C+QaFymcjfqH4Et624VXSZa0C7wNGY0rKxOOD
ZedYZw2yttYkr3P75RTOsa7MMftU8KwR/jIbomeNGcg4qqHettkNR1HU4bptNzavanyg1RMKaaZE
Qf0DpXO2lSaC/7TGcr1BRkwMKMtqb79PNP9mS8lD1qN30lfIqplPwfUm8MXoeYsQVYpazuQPuN3Q
oCtAjD+gfq/igDEKhgFRUne+p/6dxbXrr92q84mIQFyu4ddAXqHOTf9dq2R4KN31IlUtJlVaFhYy
zYAH3MAnUGnflKWY8PenJhRPUL1haF8WUclxxyWocBx1ibDTQYkwZCIYrKRr58HOorm+IajaV/2r
5e8vP5zUEkDT2utvn2uK3f4vt3R60fTrbpERPh7s0bxvKJ366M4RS+gbjktqoD4qGb8wo5NKpovO
7YGpsS/eHL5K19OKGA7WiETqo4kVaeEDmYYZT6sKOtZm+0bu+fldCQIkZRt3Wd9MtQY0x/Hc9C7i
oeydNG5O7LIpUQa3gwt0UvF7TBwu2XD6f4KycdM/eiL3MgoKQwPogePr7D+WM5QD7BPnIaP9dPnz
bnsBiH4hnHlrqNnDQUZ9MOkTzQ4sCXRFx4bu7bxbgzYw1MaaIc9hDY4hYGgE05+8rVq08kAVDezM
mDpDD9tJDLdqEG6gTX4ck+9k5+88pYODGF/7ThbaLu36Nt0vBMztSu3RGvXaLVxNQ65sG4pOK8T3
d1Dem4DpfrBiFLGpZvfZcMSGForKwnCdc5416pI/Ahzd2FeBlFu6pHaLm0g/ZSDHaAkxVzg2/pGz
WL4oAB/GyAL9TfTHekog0+8O4SibUARNJjp+VdWzjEIsKdVYCrUQMl+0BH+IfhBqM77bIGxPREo/
xjkMyhUeWGh7DqZ8XqhVasNtxWPBl1cW+B8HV9WZ/csmTbGk+F8kxhiS+OvXwq2XNhctEjQWuWDI
gclViymUWev0qXLNVw2KPMbPEmUpmqOA4pMvh3lIXEaZVMWMQj/YQQhX/EKis+vSQZjiDokcuiDR
jp4ohZr9HfvWPxXkn2Tk+cpkOLMRQf4gSyZG3YMxlWhVwRmiTu9tgxhjYIO0U6+UiSIGL5TCkQbN
G5BuqisiW6DbVfHGv27oXtsE2qXFqxzlL2o0kROFBlqwl2juYa6LnVJIt2doRUCktzNkSA+o2Vd6
MJoGEsh/gsPBagRBss8BuHRIAmgRPV3bkVyAR+zzEr3+nEhrzR7RL40YJ/Dx+YKRAvhsyzE1hxGb
xjPntlQxWik8VQ2evg2x4pYES4DHd1xyRy2bjn2b7pHTyUU1N6/e93tJBwv1EtAQ1uWFHNcKMuI+
ZogF7ArmdhUN1ZBT4RT3A73sRvY/a5Whd3XExadifZNiFm0I2ymK1SLM2q5ocBLeR7V7jbyJ5Q+6
x+/1rGAbgsm/St4R2oVAEjlyUOpxEufTT4dKL2ADFSDBzgsKheXsX+xJiognzO/wIbJ3B3kKrVKG
4I4LbMJNplA10UMEIPdo+jOwry2glWTRZmEPoO5Ejv2qHRUn5T/x08SYxcgdvH8YkfF/e3vjlNDH
QizN3kKXaMgNQo4sNfUc3cxja4VbJAOi2zuxUfJ4N95+0yb+mc/l7pJ7FKyQ6FEdIUGkrXrwICJL
KDkk04yM9dkT/sUYfWAMn6+hRNbWH8FgKFf4w+3uXhu4hxaoUXrT/j4UcKNElcdKtmC8CLecW0gc
RQL4IasLLWS/EZo7ApA7Kar7Tv86WRyCFZ20VnrSE53uBy6M455Cb4HekLogfURd3y2VbOyGjKAt
pw6xupK5w/srNwpFtIQ7pa+U+6ACLEaE27tbE5RfBlDvYTZ+ffQUQ31sVcC/SqdqdYbPtPcv6/qG
Nnfv+sa4/e6ilkJys0ANYuxMnDdxHle6EGroEtFHaB0GSXyXlT7b7mng8w80WSJbqjKMfrAp0gII
b5j2IjLW5NRuzgAlFlYW+cY48MOJ3hkVTg/JmhOEERgICpboc0ELP3qks0yaVgisJRyytJ3f3qp1
fGiFc5rRWy4LLpFXnRGOtSlE7O2KANvda8G7xktYFNr2xTHsg7ZwcpgymUh/R+QlWv1Mtt1zVndu
JpNkpsMy2ovl4c/iVQ52H369r1SMLtftv7TyG3hcx1QJ5dAW5HnaB1kZdSYmHMYwSZVwKweVAyoD
e+DeuwUeCjAx5o1hfaBXUKn2bs7ad+heDFIypuJ6b4Nrrhtfv894+Q5sQlM8sU8C7DM13oZEoxaN
QGrke9zigzZTgUJNHMLgiXKxy7uwVCup9EPNw4mEk3D77G6AmwIA6mm08/phKFZTLtQ7dXYBhdJk
0XRLvFMSLyN8UOk5TNt3TZVKOQFad5ymokXl8tCVJuyM1jbj1InMfcR4pJ8rCrDmjmBlOKVPqAwE
3Z6XKkbGhkJCWfN6d0S2DN8rz8aDqw3U2mjNfhFUvQjOSUnHxNhTd/szbWd47orrJQz45O46ujhx
KApItVJuIWYyV0r+y7JCeu65uk1zs9VNQcffPJ09T5SvuQTEZpccSi36vxZFbb4d4kpLpd8gjKcW
FXT3hJOXJJJ3bsdDKCRRWCW01HMW9zo/qZ1QAHMxMUdkZ2Qbapcs0kSU8rGuLBppfXz5kLWarKX7
ped4K2wUPA7rnvIiY1EFeBv5jmkG/LDNp+wfsG8G/JiT7LrcERDi7221hcyXt39L6/RqmlmXF7+/
fkIoaaMH1Gco3+8sg1hSf+b73P7WEKY4PavgDG8fNqd+QTjFR0rCqftB9K1je7KQM4N1MhJkcRjz
NcrgjDCGZcneMJqP2T+Q7dUO5GiCDREpzYivW5NEQdFcaI6rFoH6FTfPf5LC0lXC0QlcBZYv2i3f
WBD0gW2iah5nP/WO4FdzfJNi3A0WrbK06VZnGmC9JIK5q7d5qFnnV59mrAk5ZmAPlR4IwwjyXoNB
oxrAQc5/ZoNznNGOi/7Osk9TL2DV4vR3kEQ9454HzunVuOMg+3Mj9SlYdUcy+CEtKnMs1pkl9LG0
nCvlJdtL1PyHn3g6PHRsw4NW4QJUdBx2TKzO7aiCNe/jX7Bqg2f0Q9oBAb98BmzzFGUJdgIkWisG
uLDz5Q8EIzNZ7mDv1hoadnX3I/xA0f9C8AM32a2lyFoyJjyvydNcf+FHsXvx+VWRbP89vEV6QjuT
69pmxVeIwKYLwi9VgIoBCzx5mYxVMdOrlXis+M9VXxnGPAh1lLr+TyJq12pRj7ACo40MNmAbZrdQ
bwgvBH+harAB8pD1Ti0STjSzugye6wJF1aEvwJGAKQTAa+zZXIkoIZ6TrzccN/B/hlmMZCHURpzK
wH3IybrJZLW0l3qHN47qQQiqjNaWnGIltJnrZwvip3v5+jYpXkUz9RDw89RVNbGpfoGyaECzfwfa
4/S/bsG5fIcU6pRWvRoiVXNuVcUib8CCqedBxi4V48cHlF0HkPIvY2nvXl7h5wtmEFVyWNS/sJh1
otrCgg08UPmV9PViMsR6Su9ycHQ0b+m/nHpnvqGk8/6YKVSgUtF+8FUraJAtRgdjn3sXKdBowehO
zdA0wPjFnaSgIqQk4Q5KKOu2uGVN/zoJ5pzKl8sx/oHHyfyhyf67TDNon45JMwUrjrdqsYCjAhzY
Hs9CXkQEUFZojGmM0GQ2GRM/RxFNuh7eqCrwCdamgdLqeNEl4QspLdvoq/686ZDi2hwg9NKaB2J+
4cNe3Q1PXyQjlwHIV4YL611DTu6hor/A33Rl6HHme7cHhXfTUdi8M2QfiDIFfc4KswIy6YmxaH1G
wlbPOhsCVsDT2+Jdrjdl4b7DgpicQLQSdwNqmfm+QCe6bEIh3UzFzP4dfEsAL2/GbK0wjm/1BPO4
8UvsUfKk0+lKCgWWSFCiwgmMfU/2MfqmyW8AqcZ/WAnL4XHH3bt709dFrfoiwfAb9ybtvA1MO1Cp
uYFFRQCMcI90tzQkfNiRAZAvGbbTGttfVUZzZdyXtN0+i7nDn+ZQUEmtHGmEOaQZsZg5HOOivMMB
lET4zKBbW/0MIyvF9tUt/QalhT9WyxRx/FlxlS55gjuRZS5sDRdm2Vp4Gxq7/MAwI3KCwTkH6nOh
42ckK2dQBWygQpTyjXCBYilq41gRa5hTuOvtcfiknKfRvjox0voO/wGm9lKBxTry1gmmhsIBIztJ
41AYRTc2Glmvpp2X2IdVVb+Xeamn1nqgBz+8Z6ad9mRIZIlGemv3W5sYJTdjZ8znaE2r4DA8Ljpu
PdrEUZPYq94XcDx23C9yaw67R9uNG8dSYtR+xb5LoMZN6BHARM5x30jRMr6vrj29mk4XnRPLQ6Tk
wdZOOkijEPdT3rdYeyYz/AozfGexypI7y8buBwt/ipXrWk6lmZZBelXyq42sTc8VfJMdt8lFU7/U
A1LNGcc43IMdNKlPnD8nqNxhWNu2gchOa/jKYxUKXAKD0ogfbnVFUa9E7Vkgp6qpF6BQ8x/jea+k
XO6BII7F2XVUQxSzQBH/1UI3TQS4HFB6npFtJ/oEKL9pCmHBynwn1h1ju60SvOirvvOTzxCkK+uq
AwdfSH+zCSn0XaCik1tbi8rBstOE/K+1CvXeSWQt3ycbqW/UIx0Xb2Mz1QUWEQlBOCxwGjY3NGqO
8IDwg14bC1ozqe4krkIfonFLogcTTFJdfaXhgNkr9FtDWKLTTDLgP4VasUGI9jEbv44Slc4HTHDo
QZwgYmxgj8/+/ow7X8QV+wtuJDpyNlUCukelW98ZfzigRdWGGBaYt73ZFSt+Dy18lF4oTlM4AzdO
RJb4tbUJL2UbfaDhWUtxYsYD4JBPKZsAsckA+9ZdIJvMZH7MKam/7AFYrUeN2uzwXeo/9QQ2mvyL
OGS2XYbwRfp342gGJBl190f/lMWFKMKilkcALATdcP6V6kt2/uuLzhT0aqUukvN/wBeEGmmXjS9+
Ppxy04T/GIIL/YOipdHYUllC8ECdDlViUocn99eZ3cwCxnuAQiFeAYs9RJqlPNeRWyHLryFlRZlw
pwCwug/JFfgGN6TdrcsHOV3w/WZSZe+QAl4qTrVPaxrQzoVzcbChQPDPigHG40HShG4ueYpbd+6U
23KIQiJB3RKBabAQNosZ5NVhpBNw1Tdu6q3368ilf6ArNrzREYolhBGBC+0OAmWUoJ7fd2hDRMyk
FqNJpHH5SMIQL3kj53RkvM8C70+7aoU6keTeXHWqk7QhLmKMLjTurm582Nci7R5OR2vzCzNsH00n
B/pV2PHE+dhRz/ezm8FSzxTHOXSi1aSC+RDE8stOZtTISIk9n+DfsIYgmGMAYXzipaH63TaFw7wH
fXnuEA7K2mYgImFJ1T6TehojEc3AShhHviumxMQVO4fbOxJqxLkUge0LyzkyQmOOkRiZFReBgcCb
CxuX/F+xuA1HnukMr2TbYGWzvHbHYKL89vC4JtIUiSo/zlMoQMijch4OJiIsWijO5CwIjpAqA1kd
YJD5DWSYG++ZpEKiuIs5/mR46rOEacArQQLUvgjlE8NTye5nGJiNzgdSTiR+ecZ1yrcG8UsJFanf
AC87p7TEN9b4oqUISf2t/fwHRom46IgpMajiAS6aM3VbTDowmvsjiTnRkG5vPbDx9XChSFwszvKV
FnnLBRJ4IrVd6OUboxP70IrefNbZikS7flJaZAUxkZ/e2o6QwksSQslW9jwRInFs5YQzBfw5UvcN
pOOENY2oQN7nYnwyymKatMbQei07k6uAyZiqM7jjrxPRABgqBR4UKXuVwgGKCbVb01MDJcEsq1u2
4YMh3pTfMCBihTpUtN2RImXsbSK2LgjZ2wmd7YRY8oik4tmuwodbA6RKl0gJDpjNhIacAVWTQBRU
TdGa1xUNNCaBZyLbezBnsfNbmDzbiMXnMnhCdEQpMI8ZaGzA69QoKfC3UQ5BJ8HJnxFNWp4BRNk8
hfg3mIfmXgxuB5Ib4W+H311x54BeWC91+EzTRNxNf+ak32zAmRjmScFUAS3qDXPNfspkrgOQ3nte
Dym9rhjXXsJonyqGnZQs5goW5s+PFjt9XgrYVcp5iZ3MQSJLnh0P8dkY/fJ6n4A8gH+8n2vLmfSE
xl8jQoumS2MQjoiv6N0h70NFHwXAoLxmwtXEr3MX+VUyCbPpg/4VknTRb3q8h+H6IYos7giCV3TS
l8UtIqfXDjZTAVjkLEaHkteIgmxOm4svNgdaPp+1ntnXQ2txiM/QDhY3/IHqC5i+1AnbfndwexzY
wphsQLjhJYWUHcgdOOTRGIPNe+qqnhHAo7QgZtVyfvhl3AXyRFZ8hHqAybUrnsDiDkwr+vOlPhWo
VtOSL3lsAamWXuOI8aKAc0mHBDtqLkOz3rdLQC8scy8M4suEwKEVDLZpqMXTgp31Cnp9JcmTl34r
HDP0mGwhRZrwGHgaUXjLC+AB/A4Q/He1/b85Mp1QJJ7Rm1G27DRddEqJk2aAgt3iANSuZWUUdRaj
6+aMLtdOriDFOtBY1EkGnRzYOnFhCXjPA+EjAux76zkf3b6KL3uhUDQT2G2SMgHROmuVO/PXS7fm
regPs1ZKlPgFaEHiosEkoIvVQ2e+qfXlKfC2o/lSRvOOO2jR5/x/vNp2gNKIOo5ngPcuRPN4qkl4
0IP4Qtl1yqz9a6/vNojgPNsG9a47P4ZmF6+29RCmNs/9rGlM1mX920XZVHpjiDCvURfJleHQGwXW
MGeS10D0kjDnLw+l6AEsg/mGPBfBu2/NK580qqou6CbZALUIXSWKQoaffnWjbdMPh4Q9AUUChNfc
NFO+iPx5aodmykWVQ5tZNLHMQ7M4q9sKRy/Hp0eSVV6pHaGqBB2y7hDCK8fQr8uxvrQW4EkzuAO9
f5twVFThlknbrEqvCTNi9lfP3DHCiWwgVpBPCEWTaUsMEJW7zohBY4OHd8fl35kbcjFOvkFJCOLa
KGG68VIki273fgfFzyUgzcgkv9IOcUH/t3/VaTUsmJUJYFquebuYwIvv8uDJTS48mNwoXHpKEXmL
sKiQHzFC7NLygEwv8Xk0N1QWfJfbi5WFSf1VT6ZN/tc5DTEWcc5RVyfvBr9Vg4WbbLLNAufjzEkI
7+4YL5IleHtL6gbXDBlttAGmXvlaEq43ABMMD98Vk7z+D4h/iG9PULYXp6QRxsVw6mZfy4awuNcM
5sUwRKAD/hf9vHS9THxP/te0pBszHnzlxhWWb1dKPGkirdToahGDZwmxA5Q2EvssIXekNBYd+CxD
AC5hD2MTZqozEu0RfmoIYlutuOA/nxXKZZp02XCjT8eUlRtLl4F9fXLglZSTCKm/3APqRYnnkRnH
djwe044cZkRbyg+lbil0No1i2rZKcVh7XhoCEqhQ2iiJ/2rOJTQRYWC9diufNaAVgkcYz4SmtmCL
AJIHR7WLVlw3GBnAvhz2X6N4JZ+zY6t65Rv6aH7KOMwtfYfmc7jATA+TAeqnSU1dBbtDb4d7IMH+
Y0rG3jnvWKP40F1oyO+tZbs4lSWeoY6bnnax+bonbEZlnBqfvKNfhClZUcQa245JPraZVD2hi65Z
UJtLDpesDn5Ub3f8NriG4RSwghc3yf1I3U6WL2PHr3Rnw/uzxaAXvtZeUPXmO0s0PGOFO8ZKERuy
GogTCghtG9PqdpxM0nvQl4HxZM1DiDTR9YclISKJNv2RlD7V0m13nP0yj8A5qIJATlIn7DTEnAgp
/dGvyMU9/PXcHgTj5A6Ahkn85G4cYbmzc9zyNFAqfgreMyHkrXYbAQQuRFuiR5fUP2NHOHLAT0Eq
UIEB80bykndKU9biN16yd0ewov/mSxfbko3n3GAeBQGjr+STSB+giQGNiYPhBo0C3Zy1J4W0jC7b
39Q2Rvn63xxnOueU0VvDBElVDWlRyfPeZl42Kzn/MQduBJm61wy/O5+qt/TfY86tLsmOnYif3u9e
CIq1KqB0Ma7spU+JqTG/NjcQohS7Gxmws2tYIY8RGPOkWPx/PwWyDlFUuXRKGSFOf9X06Vpf8j2u
2jWfDn6E+374f/D8KK8cbVOTWewYgtfEQSth50AqNRWViojXOVgxBoN/0QEtsHIuUT1Lt6lfY9nu
P0mmIXlEMhvJlNpKdeEggdqKVd5HgnNZG2gjDZb+E85TaWye7HaCVp3owYJBNIH1y/uC96j9xo+e
aTqUDazAtS1m2CTWgENT9Rh7DHjkWIAzrX/iCvrHALK5QY6M7N30R2DCgW7cDBCmLOuLfWPKG0vu
4tpBZNqBsE4S4pT8DtykFqDf57eaTBB7hmiRt4RGIrVpRbtjIzjhnsn0fWNq4TXvnXSNnAvtUkkx
Mmzxt75s3/NUE/DbI92a9AZqMgcsKiNwzkoj6pFFvfXhQEorilUniXX/sb4JFzmoP7Hb6WG06IsU
IMlHnLa6fWSzDmHcIUkEZmeKeGl6tc4J+kJW2Jcq6Qs3syw78TuDnPfiJe1iasOjHEqVav34TrrO
/9bMj+JfeOW36XbQ5+JrFlnsLGSwxweFUtgwkZyYZspn0sCYpqcehE0p4y2KzFdO4W9fsQcm24l0
OlzSqlOPU/A1nvvdtuG1NwhkFN8j2dHUwsZ9emcRGtd6xjtzhi6JQyM0sVDS85xqCYxEn7ztbu5m
xHza3HLeEQHZgUvFlTT+oeRI68ibWwXHuzkQQF+ER4AMq1w642b/8Prp1Q0U/2FHSzqMywKwn8r8
KGqFB6EtOtB5JNblsXvFnT7cKEEbZM4eITpL14tlIynzfLX7RkEpqLR+KMIzFRBHR8XzfTlvyJdV
fJfrbefuuzte87KM+ZYMfiEOqAKbODNjOyEp9NviDrHXX64/AcbgXVPOsMg2mHNkmeK/yC6kN3vw
87nNkbZWMWBFU0wKliPgrX3FO5aIuoJNFS+l/eQLuH07XYg/KRbBnL0Z510B1004cmdufmo9YcpX
Eae46u/tItOWx2ug9wIPPzw/vQPec9ZHPNV3OAPS7LAP9neepDJXWVgreqQuVcQpI5Ave7f8QcrE
R/an+h+rJNbLX5WvN4398Sj3eaXxLRql0IPrOwIfQVUoh57CvqZ9T6ntWCjWrRR7k+oW8KdGjq/n
JXS/CiSsbecCXhhxhRMFT5bapQd1iVSFtZwC29HoI5IvUQ3f47eH/K8XcsM+AczKhOfV4GfZS0Ag
lvMHnis3ANn/WPso63ARYJL3mIuCyShz9jqZtcbiFISicmAxFy/A3Mj0PzFJ9CjLIH9KxmVL+VCD
la0zXdPXTSVzQOumYRkIFmdamuy79wtzVABdSA8wYWv7YmSjM79fErhMYtkpiktaSEEgvXN6n0Ht
1X0XSbY4eqSqEsYcZa6BgPhf7869s9bXHBCx0JqD7j25tQOAqwChMd0V2BX4BLxq0UX966mpa7rw
gkSiNkFUirLv0SrPKz+CMz3G5lCuRBEKETROAMyt1w+bB5OYtgyhIhNU03rmggeHKFeynLROzmIy
uT5R+Mike2Zt3vMp5AGi4mzzOdddlMRoQvMlHrSkmMbqT2apBgMPm4Y8Poibxs466o9OoaCxIUyn
qBavcYslakuw2m1znclHmWOS9I4mZAQ6K4lDPUzRdN6fgTNZ9UXGGwIY+W+873fMVqwjaFUkAzsQ
dCmgeCowDtVeA8xcEznpbrDYTd0J6gUZ+08LjxD/YACD4ioiII1PmSiUBW4lblUFqOsirM9vCG+L
JYe9RVxka2Ddaq3a35Rq5taGyqmLlxZzLlQKjlgXh40JkTOdfALeIxSl6cH02+JvC2U/jGtz+vuo
t2uJq2tpVYOj98mf7PLvaxMtrkmggNGpcd0EWpryOhX7p18Dfx73uVZ7XKB2H7+tSpAFv4OcWejL
2m8lFAdRgqjoGaZw5hlhbuRpQXjTkgpO7oSdT8IcRS2GsEt+55Li+Xwo6G/iNLkXNkCsdkD1Ks71
wB9Oca3jjMPJ0JsqfiokpKfWDaCPhoB4L0w9lsP6VUOLZjBMf+dcyAIHxyIionHFwj35Mey8pQru
tPd2ECmGo7wb/WsaQ/Vpe2pUqSRMeLnnhNOERucvCMXs9nBjMyUbE4A57tsh8H0HpD1ao0WnmqJM
MQ2X/04hk9l7auie47ec/3gsTz8ZwWYih9/laBZqpCAMB4P0TbqjphnIk5MUhD464EE9hdNJKPve
Y/0TdZKmrebcZC5P3EKHa/EsQ5rNPE570QNK8lpvN71oihU1HyqZ3DI5n0rrr6KMapVPUWXP2fQf
AQmz1arT5E4sNsv5BkW6U2c4xZtjjHBjn8b6181Un7PbJQiCmJg+D65iA1T7/EqFk9cy8zYFvlRy
DK3bdj7rOnmTc23tZSMj/R4HNb6lSVatVzr3ECbmKlm/g8EBnTEETwIs0jMoe2X0XJi+kp0/7qEW
W5KnRQAzLJ0REgj4vYF33I4LBnhegkdyfMt1SWZL0tgeEnKWr7J9cyyoWjpgVpCW1qFIuLfVRhZy
WJyImKu0bYQXxpCfG8AVHuovaABTEGwlzNvAN6Wla4kcn+db4RV28aaICd+ENBQzevUHHAEVeOH8
i4Fwn70JsccbR+QiAsptgj378CabGsicCDBzrrzD0PHYZJu5Za6o9iqNiJ7rG+4xs7C3lqHyV9GE
3PxA8moKbre2GiJl7RieMvgjaj5jm249cyU8SRcjEMLQ6YfzA5WsO4j70tOMQDhtYW8qVayKr3Da
AeJwVNBKc6LAm2mwWGoa7FBmpxIJyvU3TNIB29rfwSwpwqhZIxOrgO0lH0aw5dYJPcG1NYg1NZHP
Z5rSyc3baXOvpXdQ2WlRedPoITiLFmVzZaQFS20nbNrhDuowXxBnTmMmF/91XJguVZdo5IELG7Hn
RSgm1MJ/bpsSDIs4uQuhs1pZCM/IvjaEu9J2yBl3CKWH4bJJCSkvoKuf7B53U7MrsXyjyY1RpMMp
jxyQGRWMq11PmGp9QuzKZM9ljWt6E1bl3OPINaYnuGBeUMwUvIGWO7oBGL/MfTMUWB+Ci0yLBtSA
NxEJ2HC5pmFgMiLk4LLrN9yhB4throjtJdSrsv1PNR9ikAj69xdoWDwGBjRVTKmRmkzOx+9ayfeK
Ylb1zwYe8KqmxlNZ0jRkrtpCj2Ux8A3CRyYA9FxK3MyMFA1AymCtTdZzj/UiU+XdHyy95AMbiaT7
da0ORYqn9TyGWiNIeT1DzA550ZZa01h0nkiz5i8qDk3G1Jyb2U/fvPvC1YilrezoJSp8gVgBmc0J
r6PRvPSdR2y9PZFHy+HWD7bHQr3cmxG2BWYG2nI0q3w2UfRxgxK8lPGimlYPhomUQ/khd+sJHUra
pes/2v+4w65/CBlGJ0HmckE9K7fkDxuoIv8/OE5H/dOnmAn7FDHGU7tCqfPvcROVzNrgk7q/BVca
2l4m4SyMBX3QdC9IGMvhaSHQUYxUiiWYxNthU0SRbkHqPgwk/tVy5ABC8duNBfW2vrRRQ0OjJHpA
Z9mPf4ua3YmZF4256N+jyFPHHuiTpuEaBe5Re7uzNYK/1s2AowOZfysBxgVQrU9bPCm33ojSBPej
U2g1C68s+mZMhYNyQZTZC5uq1eh5/BdIuoSva43xhEc3EvxkGIfFa7DeCWl4+HwqiIaB2lfzfPb5
d2u0nMnb26JFFMw1RawooDGbmyX+P8RSjD2QCXv7aRFg5fF/LTD/NlzNeYkIarS+bD6tX9zt12Um
K9eI0Q5ctaH7PnagPfvkhVGEmpl7UqKk/wD5DLreGDEt9knxiIxdx4yzIiXuR3dFiaULnQXAxPV/
ZVtmSBvCWk9WJE8laU630T3TJqHbFiOoSyTfLvvqjGkoLo9LSkMWfC9+MGQuWYflocPKbAqCAdde
xf+EzTw4WT1VsU8RUQ7IFgYLuzRG0Gxc2KuujhpoyMKK9IEbC+63sjm/CV1q4DnMyyIKgHzpuwMV
nyHNP4Npv5m2PezapWMwz0Qz0Jfuw5vurUFf7F/xj17O67Pv6xLCw5FtXX0t2Pj/lXSzTWswsrQl
Gh15XlCc+pl4m00Zp9u02Fhd1/F6H1pL4nKNz3f2/XmXpHwT1M/Uf1MkORpHDBQQQW48xZRO41gk
p8SU4CsFpQjH0tpMqPzTPDqmMjbK43j1g0dhJpJT8PSfUjyF69qhV/Rq9svjo/ZxYpOHFROmBSsq
vJDMSj1Qo6eEqpl29OqdM3pOJ3apZNvR2ZXnKHrYjJqT70vOLzNBu2L6Ie16ZBWrL23QZUEkV5kD
1suFagdwEoi+dJmRAKncx4MyHZ2QD6xIa54F74pqPaJs9acHIxLDlTvvhryt6x4Mw45mdddgC7Gt
3vkhDU7yQJ93OLTOYXhy6nv1gD3IKjoRs2FDaw83r7jydl7yj0EwvPPEXf3xZeMKhA1IefBi5aCG
uq0OE/xNQnyT0JxLAdnv/F7PQXbH3ETTpDHIU27bEqGWbuFvgRXhDmv8pZD4eQdzS9f6Ij9QrU+7
WP+1u/hSSCZbKXF/EEDieX4ptD+S5rZtaIPLJkphrn051/2ioRaSgaFD7A6Xj3BXqThuit5uGZ5H
/1ArdVd1AZvfUU7TyP8L5+nQ+kcNaY1zI4GkxzAnHomqHwFKnqUIkNYz5l2rWPaZPI1GNG7n1fgs
rNVYxhzLitqN3p9b3erRQm9cVojd9vRB3OX+3795o4oAeYu5eiu+jID+Pq/mNo6OLfOvx9IwpUJK
SnFwpPZo2/OLz8hSi3LBWfvBjN6mB3g3NMCMohyOJn7OvzuxhDpl8wqfGNN+wkTMoFie5dAvxiTb
Ox2natEx4Hk8n+h9NJPxLYyCBi/V97EhnW8KuV6DJ3lwOPzXy8duMCyAKJBDd2+GH8HuRu2nTRCo
retM8wml7RhFm8TvMELHeuQKfXY0fs2XZhEzPLuvS191iJXN4f08yc2fxpdB8O8RYJQ1+WAibMD6
X26ah0KWQkZese5c+LHKF0RChW2ZQahS1C8AwhTG8dR0IQ315yc7R0kKS9q/moA8HDldi50ytUdC
xHzz1e83KnBATedr7vtMzh8PiPQaUX/uZSNc1TeMWigmFbkC3gN46n7ztshetqDHK1xxvA+IyPZf
70CXSQlTBV8dS+go0QtUuc3eg4czhSbCADx2g/D1+9PLp+eU1ZE5tAu6Mey+6VVxQdS7qvJIr2Hu
vn4HT3+2h+MFtVB4kbTcFZS2bfKwE8ePsJN0tcmF4JfZDEIoYExuK09qCwUKzDOSrQV/L3BdIjac
bHO1UY/UTl4+eNjy/B8/SS6oSbiKJpH+o8BJmjVULH+n4+bQUS7CtKSOsfK6/SCoAopZmIaugbrU
+15zxXtA+pWaWqlxxoqTKa0uJCXLxjhZFc81LaYegySaZvv/k+PLI03y5TP5cbX7x+zYMJmTPLGN
/3CCne8oncrvy3+liU5BiD+NAFbqH0QSLgbcETAlZi+2u+YGiJHaIA4BYrcaDRABV5Jt5AsFHZWa
g3dYhT9IBKdEfC4JVUp19kOEqrNOTIjSvuEVL08oNJQz5LqIdWt+ffUu03TMmFaYZBQmpydG6w/u
cl9b8cBvwDMQTA0Nv0W59OjthP/+J9aQWRG0G0lhcT5vYueYAl5jmjEYFF/PrOdxTTr688I5HuK3
9IYUuhIC+FTpJ/7/NGoMdP5Z4wI+PdfSV+MzuZOfROqPmQJqjxpEfKDSBfymyDPukimZmETLtKEr
pTe6j6eEhsIGIH7j9vMsFzjM6eDGCCZrrz2G+e2hQeVgu7yit3Oky0uTQD7qj2jPfr90REWdq83n
ArpkN18oVefnZYD9pfwpsv0iz3RWxqwClE3AIC2Z7RaFIxzBB/8W+DPcHqmcpw/t4eFGPzBzE5hf
M+sktXbhWg510u85PneG1fzjExlFBX07HIN5uAhKddOr1zmZh9AeDi5x4a27eYP2UA1L3SAWPdl0
IiXS2SyA8aPiDn27l1ycVoEy5MY3lh1xSgOZZ2pTKhLvYCY6UwoIOBwHvG8HUYdOhbYWcsz8NgZ6
noZoDIILiXvsZTygaX1JyVIvYMdjL6kzuSTpEOVlazfJflJpRA1VXb8Eq+0CUvPPP/jqD7eaIJb1
MdQ1lzJ8Ph9XyxhUGywc027w3AjB/I1+KvxsRQ8nJCMKKic6ovbMlE7N1xqWVanmEEnHJd3fGmyh
DAgTMtKchCdZBhZcgYc2zeCQp/lyuo2jaM/SUTB5anQoRsojfKWiSohK/vc48pR0TeCi3SH+6nDR
OHeYDqfSLU8FBtzGXvy4DkiOyVR4dNel+NoOwXFSWAqN4Rw3k8GwwHnBJBA5Df7hwAE1AvPwAz/p
vmOkHIVVcTm9l2mTqcAw/XMv0HJCHDS1Gq3vgX1lCFy86a+AmurPRqfy0Xr+n27bRFa2HNKQSq7N
O/V0285+nwQhnwONsN+3hpG8JTpQTDrVWh6f5swuOn/RANc0C3rMWjG2CWdb0zd/OjxuojiIT0B1
2TRpT6Dfse6hUMhFWNB8dLOmGvNqnM5yYqgeWbyj9uxt0YUsF286JbyWqf0ifW2ppXRgAG2srAKb
DZJIVgDr9nQVu0/VKdaXk3kf0lNyMZiGmftZWA1Pd05stABZE+b/yDw1gVxx//Dg/9o0DArDbWIZ
ef4DOlDACEeaISF/b1oVf0sQpjTx/z7gcKbnVJfZGaC6DBpgyM/yRoAxkTdXupGosOZocbMv2Ek5
Dv5A6WFSfVWz9QApbcG0sQ6JZR57ebfv+qDTsKM/7WYPZqmlSRU4ZnDQKpMgY31V5UBiHzmrq0rC
YVErGoWW9NRZePfXdRXu2ZybM9vF69tdO5/HRIEszkAOYxyHTt3dQdKUoxeDv4qV8oXb14P+hdbE
KEn6PGmsmlmmHjt3Jv9FGfgaMPqLGxuShDGF+ED6i4ALGgYIsrACsvvT6cOQxcsNWoLDTeSpwuY4
3LZF0DyyN8bJ+N+GuDuLjpxwEDBlLo3TxI8h/aV7DSTjtujp/EgexL1/XxAjcH24CDoKWtCK/pYk
LPv7NW432vagD4CAz87GzJKw/3m0n0kjf8MJ0Csoexk2hmmjzeSyvnpXT9FloGRb6YV4HlWbkCxf
NRp534HZqVk7ijZiwiK1QwGSHnDqTJ3QO6eskbAXDY1iLLo99aBimAaTSsYrvW/E7FLAGpYyLjoD
K29sb2XH99bAHIwee5KCq+JYzWA5a/oNvtge/kDQ/yOtO65kcW189ftlRL02At7LpkI0AtN4D53l
sn9Nq+MgSdXpHOc7u0d7dX1Q1aI6gZywlsO9LlMQOp2OqCdcNw1U4SANQMAN2IrnPonvVsvEwDzm
EQJgKzmyLTHraoVtZqFjR+DH2XY52CCJxA6C0cNi5l1NTZXrxd1y12wdJGZkZ2eUWe3d4t+ZARgt
yyWnNHfZX4wRR5BuLH/c3kDiOdKztiYNbt2JuV8CNGFWyK910sEhLJxFNxJ/bi9UOjqS2Y8BT0j5
qr0A3yAfFwCSEqQhvaak3AXtVh+GZjt1Cu1UKwryRTftXbYtOrBdXxs5stObxPk3FWhK3jnbd1IN
zlyVa0WtbFuU7/0MZQZuaKvAL7W2IitLBXAlAqLxh9eFsg6tOz5MI4CA/xhkJlga63gF8sH+IDim
+LPBxrzSM62EpH1BsDA1+Z12kiq08V7Bdw4r1WqoCXQhhSh8FJjoVwkXYat3n+DJLHJ9GIClg5BJ
HSb0BxLA/TBJYXmBzdmxbrBGkvnNM3wQKFHK0M/OEy8fGpyiV6QTDgnJlEpLz24g+urJzbC3/guS
H5eaUPYiIvQgSgOQmT+jbrgsSLngdOzMHSmCJ7xyH8U+GqGfORk6p1cSo5j+4QH53+sZGwnCd3T/
yGij/mCZURseW6T3xIPvNAHMKyY9l0F26il0GMZlYFxgMxMNHmJgVgd79cHxYQrfIF5+ZAamyHKB
s7x7vQawn7J4IcYT6zpPd/WXyQsnlTdJh1KyHZD0epUDaRS2daZYW34fNNIqxOsAKxw81536zPid
PXYC3kASENdkqs7NmynHrlRf2KvM+2q/hAt4cv1XjwjkIo7JZ3HHUdpKItSAM5fwl82Y2jPwrMeo
Qaq2It0d4V+TswmseZzb/AKwuzNxpFrF+IFEfKbXcoEnQQL6v2KgISSt8W2OiJU0uJVxSfY/8fHY
P7ih9hePX92F0S+yd1KvZt50qgsniMxzbMXqOm9hHgbtxcA46mhfPy+cNhPdxRsg4oaQMfJYnTxc
zBg+rre478eDQX1W82xmWNhcRnUP1FfyxwkiRg+R3MFtTqx5eYhqyH9KqpZNV21DTJJgc2GQlRaK
gHEnj9I4wYC7ENXzl0qfqDwz5Fy9umHronm1PeYfztd15pfLMp/YUMtJdStyU9tVKPtuL608eCIP
IFrVf6XwktJaizqLSXoKllAqEZVtbt7XluPmzNaHHvmioJAIgasSmdBdTMFqS1lK2KIYeNDaC7Uc
rbQauLVXjDGzYmAo4ilMAuyY2TqXsMY0MIDVBB5WuxC85CWfQo/5VAn8RpytguVLOKp7ZIYEZT9x
Lc3aPnCaY5A3G4q5I8hCgwGDd8t2bHl+KhxpjKP/8HTC90IxhyHh+FpIff7kInsBvR+TpSXT3vDH
aSpnLq3bZoTgBJ2NndgnJ63ZbEO60tvTUq0oy8C8HgtMhabW218VwAVSD8rbtbp2qCO9hT032kfH
q3AyMlDcAGhGWYAhOcZbcZBLz7iPcBoYjMmFuXeGL5P+GkOAKQ7s/fBJAif1uY3B7DCY572nx6c9
0WODVM2h/EQtSYSlJaJtYq5mbtkBNYNnNJ56IvAOpdjUqKq4TuhS7zzfkLHpZujJXpTxOITZgou4
Kw7UD2IA99JAlX2CCN59shDyvJ4mlgeryNa0BMzJCwtvI22L9SLTwkXhajWzbm5jCQ5WzlC+Gkzy
43mF+hoyI7YM4ae7hRVIc7GHo5WOoXbVb0yI6d9W+9C6Lbfm7f2zdUYQnZ7N6qBo76A3G9N85K0a
QEq/+qYfmiHj6LeNnazCOGzeY6r8Q7r37fMsR9g3iBENVVywWvP/boeXOlk5oA6joYatZaBxbSz1
4dkX8zFD6tUXl2JNVcr8dHLVFBOpyfXDEvFCVNgHK7z91FRPCBdCu4+xUxOFGpxKYf77S8UvtAqf
Kf02EUaLTTxL80OdPW0GMC2wDMKPCXUmuvOkmHE3/eaVzYQ/W50rL+oT7trCv+6scO41ELQAaPnu
cdDSE49xbA+W1KmC+Ns0TdzKDRvwRYLy17h6apoBbADbGlVntKDmQe+NY3wEWD7vxRxMF8dUBD0N
Mh7SI8bQ+3CrGBkt2SRUvNRSAW1K+GdmFKhZthlY+tn+TnhzfCAUS8y+RqMgB8dV0IAcwL8T4SBo
ED1CoXyJD5HFTaYDQMXQKIgI3hh9gstGDzLYulRQtqCpRAXh2nAktDLAcsH2bY7Wyh4vyetYsk1u
k6pfE1w/OINv+0ofnvp8bACIHybLVf8LX9q9yR3S78m7ejN0fVcres4BxXdtQGj+NF7v8ZEGaL6l
mSGuXLuh/mH99QOfKE9xuzQ9IYKhxWHH31/CjOXqC9k+gyYmzkd3/rYu026xn5bZG/VUtogVy99K
O+BG1ynimJuGaw0TeKtfwKeFiUnVBAt9grcY2CBFvd7X5eCDHD1CcSuDpwvcbb0Lfogk+FmVtl0T
eK5OW3yFSqzdk9bADJtYeHGtXRxmecIFzOmXFZZF51yE+pgCb/0ChnofLVSrxDyITR/hIYMjpOzS
2Vxs9EbTX/V1mjDlkINpneJhEhGkq/GfElYHARysAJ1cQR5ievDZ+Ie6LiAfpErQ7NrXGPBO7C/r
aZ80DcrjWpuPe264uERDagg8f+ToeqtF+Ic/vtkDBsKkAfbD06au9NV9hyvvTRcbllwDTj574Pg8
98V+qsBFZsBigbZFyc3FRUD8W80f05W78PJHJwFZCOsNf8bPv6x4TXbtDE3iVGqXvFL26K7C7VNK
+hXtS6hHJM7S4Dflq59oiXblkseeFipCscNRq0ErPJxj5ULjKh7S+1/PUHLrrRlMXvVhAhsOxN6w
Tag572CwZKN8Ed1h5RpI+63MeV/qG/ez3qIOnsO0i9SztNr0ykQIsAI7vlQv44A3freWHateB8gy
lzXb2c/okA6DmXZb/jnGZtj1DoBwRFkCCTZeoMHZO6Gvp32xTntBe376s9RBScN7OKCaPwQvKkTv
IcCKVK/ZXbqp/Qmyr+quuEOxlM94Tlm65iS8pW1wKgTq6rAaJi2E8y3OgDEdwOxCHSkiz0h/KAJ1
jMkGrf3T5xzna0RSD2SCxU5j6Sxf4TvAtpJnQGlPXFADerksjOXNltqLHRlJLfx/w+Yk6EjdRH2d
0oBLMJcWf8rokCvWX2BEsDO0I2OPTLRJR8aNCIihxl+0z8wn7ohauHXn8Ft7ZIDW695X+rhEBDLM
/DPYawK6yL8sySvfKOUa0c8vAPSJfw38ZU9RbVlgB68KoyFFYxRwi02/1qzhBit7AJR/waGLhOh2
oe04i0MueOv8GP77FgSZLVdjTJXnfaqbP4bmBG1rmklaRSMgYrmg+OWjL7LJH2YWdW3CNijb36Of
faUcamSuTEhzmiUb1LVkn9bve8247/IDhqTAVLaKDGUfaOPKTgC8qRaDDI3AVUN2Ts5FEMN9tU1K
eTt1qMWwmW3qabPAqCVn1nxwuju1fnx+zS+2XF0c4P5q/E5EP3SBKeekpJuTnzjJiWty4nM2mHuW
h/35NjO6/L0tpoCRgaiuTKevTm7lvI+A4bbFxESCLlul73L52VOKEFt8SGuziMTPrL3pKIXXoEl2
0Nk5ZMjxDr9uqdW588qll2WGBj0kW5YHI092RB4dw3UV1k0EY6RSJq0AnnnjG+++SnLPuTKfnc2n
r0OK/IqGoBLdsslU1hiG44Z6eCMB7u6m7m1gN0ITF3fSp1rBNEdGDk1iXcRzT7bFIXDWg/bcv9bq
+SxPgKhm4yXZKDNCTkQDcibYCxKN13RX9fbEYwu8qfZX/xoI8lOzcryFy/CmUwY1LHcBJrooeMXV
LsTbD3qEtvvfmFt3oSfK7XVIEEl7OatlGNTIphIBWeNFW6iJ2gbU2qMpB3JFt7MyLN8lxcst/edN
LpU16Qcz+eRIKThfaxBgTalEi99s98XZPgUn5g3QvM1UUb8P+XgZoefDnuKldYUEr6lMPaiqr6pg
Nb7/zCL8U3P8PurmNZYh67J1X8MPyi4hub8zpYT42PMc9DN46Jd+lfFwHG9V78FluHekSYJF71kj
i6L4/GqbbfDuCdrm+EDJrveKASr0bNbclXtV+qPQBGc6rFTp+oNW5j/a7yy4zEsT5fgqsEGk4+qt
qgmG0trvIKPHvTtl7+qrAKzYsJABjWl+CjkeWCfqf97VRnooUsDCfHAPUvD+vEMJlULpLxIeuma/
8oMxts/EQj4Da3uIg7csxAiuE0UpvD1fdMXVL74bqJgZcLGFpX8IUBEjeCwg7aIJ39qNEzNFeISx
drECclbYK8H9vmfEKxrM+2Tr9RGFugXd/OP/ZdRFtNlo3W7OLU4g6cjMTABXB42i8ejTj/o8olYp
Lxjjft/J8vJR4DC4Z4yYPuRlOW0IwyHadi3SwFmceAD+JPGBsshGZY2hzO4MVgtfKMusWc+D0v8R
cB/lyqTm0D3mznG/BgtxKy2obNyzw3HANAVm0YZfZiMq3A6Tz0aS4/orR3mxA653WaaGOUHHvYXu
4OEVgoBnO+eGh+H/WM07blNVqORVPo1N2u2CdHQfkFt8/AEDEuuU33UySQrFAJ8C0VWudXso8AFG
WBRiNoeFgxx3Vy6HQPV0dOFP+4UT4ubafT63lE3BjZiJua33koGaczJt+dhI3fJHyiT/pmiuPtij
ruRjrXGesMkxzt9gzgI9TPXuzBe4sMHF/40mP/cqznsp1U/Iwb6rJueqJWxIZNutud/57Zb9+7ft
1+k93sOnLEQGLrgB5txACOoeixXN/6SYmuMXuYFSDQWi+uxbkf20tP0WXK9e8kFNGPH8FPcuTgxf
P0R8DVsObLsr5BxT7nQK4G+N1FR5K9ggwgZsgnhDzJuHYWwdEnuz29mihTbV2An+wy/lQtaHReix
vO2Ox/XnaKpQ08eZK335kw+tggAYFnkHi7YvwXzrBMQ2FSCyjJfc0Ib7B7uHPAvfSY3/LHl2Bbyz
QW4a2iNhxs+KN17faxKfnGM25E07/UUbTfhPfn6Hg0xf/+Iwv0/smn+k5NiiBcmKCHXznXzD+0Bw
FzcyEYspoTzeiLGkd7+A2eMC/ALss1tkarbmb4XPiSCqubMKnu+wzyfFZ8NlQTA9cf4XDtvFBWIv
ZK+HWaHXYHOpOAhK7CrJ0DKf24WPAP9dPYOIl13DPkALeWfHvGqQMfQv61uOwsoT8RZrsuRm9QY4
SkBs02nTmgCC4L0e4j24wM8Ci3zfzzS+litTHfBTOOwfJswy8xEoPU1icqAxMJMaRVKTVHgNlBdd
Il2IjFcCzNhNYOewdiC4yZ8AtJ6AsvcyWS2F9tqgE7y5ObxqSOGIRySQEcOpm8QO29TzdFMekMJn
a/I2sohxyYo4z/wWkp5lB8djoSUGfHLbtjz1VqIRUrV7pHfyelh4IRdnePd5FFIHn0kqNAgMmgq4
r548b/Rupj05kNwRKjIdXFfDZPcDK04fiJrUMEXHJtTCNhYRf5cDsZ0LYvIGc3WkRaihMX+mHRGW
JGzUiZNfF8RM5EKCUC7zTF2ObGBvFg86xkk0mFXh6Uj7YWPJlR/W5PmLlfYtDsFQFMptnJXZcmKS
n0oNt1DClJsu7QMjif+n5uADEenywB4wl63MkcqVlKqjDuml2iF/LnsFGOS1qkRXwsSB4bXtMCBN
fvoK/1auapBZR2dry4xTJ5o8RX8o0KO4vbAO4i3CgRBLT2OQJN9/OCE55NYqwc0KKmPI4gx1Yt+y
tZn2zaIDUWK2Oh7o3ujWO4U6rOd4TZoWp7hAWV/m7ZqJkEk8IyfsdaqXsOHrjveEi2hofP2QthWN
+cpQ4mxdXM/wnPjPUVLqlVhDVFsYA/Qt/iPWuUvKz2ni+loL/7l54RXRFpw31IE43rgY7XjhztE3
spI5I0jzhPqe1xYQ7hJ0KoGHKhAQ5SAd6YK3NoSCnDnY44ZAzHbCHZ9tE4hXaDHUDAdNeeTQjRCG
fM8No3hM8O9nNNnnHa44JnyW1UWUkC1ef9vTk61YxpciJYirwg8sgIUUNeQFMLZFj0pnxqoeMJFY
93E0nNPaNuhL9tbT3W1dKGrmxwgUpKc3ItocsjjOzxHGxBdGZBbzMo7y7nSPm/NLTVCbr6/JYVDH
x/S4FUtyat+k5HcbbanX35G9yEqSYgR8YKGrK0uY5n1ImhGab33iLwPqQVS6Dt8U2NcyccVgzQ3q
j8PzAuHL9zt+NTXTFwgsKpvnAwhshwWPbbBncsmKOY+lBKfR5XSGk05FxU9ijXCBrFBRhAxvxKve
DYrDoXfhbXaDHEuLJs9+DvTjUk3SbqkRs3l06Te/DqHL8ZOOQxltDHUxam9NQ784rGXAZ9UB/wVm
1bKm8Y0oWdB9bMjPqw2C0b4uMUz83dBlo2mV2HXIhkexcFi9tROz+AJS820veCe6YgrD2OIfEgrN
XlPWOwJgX3D8jbDkkFdAPKZTbAkhyQpesBRpbeSdVNpuVUHYdnFsDGn1tSc7SUrsRkYwCCxPe/pt
BDo5zSEHH1XMKA7cfTz48UtDJroTKgcThY8agUMI4zwO4Xr8HKw67CBjEI592P1pkNW7JIXDnKLO
vEDFW3R+PuSsslOeawRLFhLtumpfmPmEvlfn5QphrMzo5c2kfjZyhQ41tps7Xme6mYwSZBwP53Bs
a3sQilJr9n9qKFOVOkkc/pJtTCIvfkK55Thb171OSY8Wo5Mw9lHL9MVbxy75ZLAAWnoEpL/a8uJR
WLaT1BDmr2Qqux4YdlZBQsz0OMTdDBnPfGAlHJLgP2jGsqTmsegw5bo1Mh9U9jue1huCakrdwdpz
3/BButiVSFV/lX8x90hGYA+C/nCr1Zp3HDa/bN8rC62MGEX/z9l9EqtGyBQqsIR4o0Hrn5uqXH2E
JViqcsNcthvxTAWQG+sSEIlB6Tq7AJIGkF+UWhrudrPEcs7gvh3SqJzndz1Tjb8ZccL5B8QxkhxK
pF75l8LMx2gh1rHyOst4V/6iI+KfLLif+TAjxTySAvBkx3TEYlj6C09PNhmOmNgb18dGpxnHVsCn
rD70cGrETulHr+x9+RyFPK+3PVZG3/DOzIY2GHRGaA3iBObkKLZD1sIx0gIY/mPUidxGV3X+AbQX
zc1QTx+cer0WyFmj+aez10JyU7O2MK1IgFDLTRa5ENMY/8LE91AXs+sth+MNEeylMrz8mHrmLct5
ImdD0IG2WqZ98eciZKFkdVdqmfyb9vxW/YOARUVW1ogsC1Y1OO3Cdjz4XoU6UOI2sjcYYDKP+1lP
2fhyHqNvIXIOdYnYp8gFScdbt7fIVOlHwqPheaN3sOxLP7i8MeoVitNVAkApQmbh3P+T1Kn0c8TF
7RBh+QltDmQW5g3L15a+cyAZaQaD4/vEq5ruOABel+5xRBlgkLF0ozkBrgnNbruseoRxsYBm+nq+
6M5S/w0ynvVbFQA7UEagIvkR4b2SBsZCKcFXC56LHy3hAhCrHcmxcW0f2JwEW7Wdjbn3SDTUYCAV
LqDXoPTUqMnU8SEZyu7acffQ9EH93FsDcH7eoxKMIr6lWzYOADtwASVDo9xjXDLe3kf5fZo1ZEW3
eFBbwUbCAamn6v0JRKLbBf3vnsIBTMvsRH8Tywr/ccxr0kYnMl82I8plw8hyNkROyUbOKguWCq3c
IGKbWR8lox6h2t4/P5eUwD7fRjl0+zOfTe6Cid93q4MRnSOVEyZyMxAWSrZ4eDC6N72gtGEJqtGO
Ktc+OT+R+pKnUIOmChcv5zNaVjKsICKlWa968IVUt1p1eS2BseRfykgyT7/qA1WoYNknMut/yufx
bSv2lFI35MPZ7duTmc1p29s6M5Rqd7e2J+b/aYWVTXMKeQBU/GKahXZ/mcNBGou2AQ8C0x+sww92
ERJ3GAeRxKLQ4omhSQFsnw+si3l8AGW9ipW3i5uyPkEI9C2/miLJ8xB1snDb7oybGTEGs8msrbWk
0piqxZ+t+a+OKN+uzX5agFMrwUEzGRCLSQR2Fp39Ki9Z6ypGtirIKB2w4y+EvvZHer/W9CkvTQdo
/C7XBpu/nS007g7jXcHPx5s61Y4+rBgmNArwU6jbre58ssrEgI7tTlKiBQTwZNQXGv9lKWBmwKeN
Z9NvSEf/tzGlU/9QBQSY9MFqM9VloapwERvTwduwitm+rs3ub2uF03UyM9gQTFRFyHH89iIthqAG
7oj2OzvfODt7+/zEJ0ez1rSRrJ5qVT+edlXEBPh/bf/dPOadtEMD4Vjl5GCfJrD0xCiWkFUDa1Uq
SJHRkrU7D/sWGXxkcREIkMIAhzWokynFNN5acXvEJDteu/WniIWHQ7WHkx52C3eOr+mO8B0ZotZ4
nzezZNjW6UUw+zRMgTfe/MCLdalhyJBLykdbcX07EGeioGKulIaWlSVLfGxwepUpTsvb8xut47sj
ye7DgpLiL5GiyP8B5wTtlUMvQ+GiM+Yk8b8XINf4r8RN8Y03RFzwJPxa4wJujC4S/cyS6/mMMf8k
mrNVPjIi/nYt9K/kLnzjE91jjEpYmbtmM9XI3xbWJwjlP/Xo/kYk/s0yGl1YAxT0VdBnk+cqjBpH
i9GoFs6nrT9CQcntXoDzLqK8f2LDtllNjWjizIL9AkPeGr7jO4RYFVGe7ownLaOyheBDRwV0Cg75
G/Mf8zCDvz+XhcGg9SzgX4ecWY3Lc5jRiaSG/kA0PapE0pnXoC2CMifzk4q5AiwL9hwSbyBx0gef
IekbhJ5u7U3OpClC4lRUwUyL6DB0AAJt8/Z8G6XGhPBP4738DPp34Ag73UlXIrzz7KJiXLZPkqhI
/IixQvXo5pmKqvUo9uJCRcpWcmFWnX3UVJAXVA0u4UYYKfTmNmvmJ2NM4TUTfy0lEh9bT5p3xvLm
QLyDsPXzYJkPOs35WhgUKWKVzcXvRiiLwdPqBbeQrVo3HNTZmQwTT+vJA6FN7ns4UF3oNBTiwD6q
U9bA1J2OeThsoBSGXsuQFm5tqPf4fGsVx/BsTqIB6t/EdkkfFu0+n+gSJvNkjopS55/IZKwM/RCT
9Voero032IZC0em72wqzeNOMC/G18S7Jg4HGJl4lo5dBXLgykgrKVwttdL0lNykvH5iy2pCV8MIj
vkTpJTyfjkNUkTuAujCC3sMk5+CYv2ij8LfZqe8029bOcjgTTd4J64UX9bkChYQrKd2dwqg6RMyX
eUhHtGdTW8FNKQA46S0CujyFsiG6ak+LgZmlXGYd4oLhWAl86aN75Ve7n4o/z1R1NAx3P5X7Ams8
XuYTGOjTD3EVy76Ape3CVMKxRDbbwv6uPW8VepzIvR79goJc6u9GZoCgQ2fsZj0AkD3ASuKwVQ1y
Gs7AKG0DIvSD1zw3WgS/MV7ANFldf64Zn4vh+lHtS8tNG05x3oWhaulecKkW528e2SSjxZTkmkFo
B5b7OFnPh7unRcu9/TMf2PbS/WdUX3kWm5KJOJ5zPFQr27RMJYkfunT1mtrKJqaiyL1U5uhVUQl0
TnY7V3mNNOMg8Au03KHoRpXWHMHusMcUPz7Ci8+M0Bd2KRUzuPnN0bjBR1LS4ScP/VOFR7m6Wpqt
iq4iW08gN2DUL2oivsTv0gwF0N+IlOkcaEfI2FcE0RIyjHIJ3XvDbntJW8gBWDWEJ2nDZKjz/m/a
L8jlnLVQVmw8pFoq2A+QKuDQuPWPT4kDs1GJeyAvEjnxkzmPgQUR+cAKQj4F0YX3GF5AUkBADENG
eq+V7JUszDzLiIwu97nulyPck6tpetZrIssgV4miCjtBfOLckGhqsqY6LLVQeIVh3JEOZzhUU9cf
8UxpN7WYPE7F3M9dbzhuLWP0rUcCdBC3egx+yHN0b6PR+DLfSEWvsKRLm5LtYWDJ0E8qQX7fDQ2J
RPBakQdWtC/fz18JmzAnaB52t4AUuw+6Bml10EiaLRGZGcJP7z8pUZV0olHIXJSFZ/RS9iE09nwg
0SVmwyNV+Gy0sw9qCupYsu+ZN32whMi40YMlcKZ/vfpmTrfiC+I4VnwO+ixo6Gfg2ld7JhLBPqw5
0iosfNkx9GPBmIn5Tb2XMNsUGJpDms6JXSwAD0yGkZsvkoBr118Yk2HXWt8nql8Aj025KXfTmtSz
Yz8mIlykwDfToxL51fAUc3QDOsScY60ez1fw8T7zjhAkj5c1fUI0DkvBtbvDMhwl18FWfBNiVnPj
U+jFoOoApjbJrvdDPx6a/miODrVAlXJwVADmMES2g1jpBizjsuTsvnhySW1DlBIh7SH+Jf7JIz/p
/BvFpw3PcYE9Xdq1OgtMxsKwzCWh8ek3LHVMFX/Jr9gD9m+OtrqGEnPgc9G00K4Dss0R9DUohG2G
t3eppAN/4vvTUc7ShvhktEHylexS24MmkKe6vURAlyYIn//0FLSoI1SZ7FzNNXVLm0mnXEZmMXCT
vMyevapROBDn+ZREep0LaadX+V5XC5IuVnhEVjAvE/cKGrefknyVZX+7p2B5z4OMWSNC1qzxX7JS
D7QwrSovaF5e4pXp72pMuF0W9VlC2Vrg45zKd8nPkH5IJhSkI3rSEprHjyCmqn85f1WZJDyQrhxc
ucoZ9DCjEALM5/limPfLn0ZI6w9K/5RWJlP3SG7eQ/1xBea/en4SDyhNDXT+owBwPvaAQgZ5+nyJ
ECAWgLTtkvFTVTBfdWMo1gKZ2SxQKdNSvV7Hgs2lEsZm/a8WoGEjywzh5f8NDHh+qQXljfNn6EFS
tG5Dm+EqKFG6qQvviZ6eoHZfOvpAGqMeFEJ6GHpA/8r4/u80M51I5zTO84ekXmnYUZWnHo4/XGuR
JkCh/QkvRpSlbMWoTnj4tmSHJMow8Tswwpb/Ti0FanQdEYrls/JK9HAb2DDm2NfSYREx2Z7b4/Pt
eSxSMrOXKJl4lG0U6Ed6iyIiOSAVWhgDkusHe61G1ha/3Y5jsgqp87/YwdDaiqyb99UfKpTkGW4H
xJfaZY10bn0MYtHaSHo6hrePSIDWkXxnDdV/FDBY8wCVQui4jAZLtUL3yVCcwrgK5bhXtN8+3Lko
dtBQ/SowPx5YZV1iwK8lRyLw35GxscfTeW5nhVmf7HNcSwKeckffFILN8xKe/4SajNsRWgFIosvo
qos+pKy9r1blxn9NtAfDgeymbhGeMccZP9cy5hNJ98axw/TrEdudBfe3C1VNZP6dBlTV/vmKHJT/
tLvvWbe67suScYCNgCSDKP8fS5OY5w3fLSHELI4MApkqy5L7u5MVaEaop9BSw1DRN9PBs1tkP8GM
bO96kEvKD0c2SA+/l5mPv0gwIjC3mrdzOx2cRuOoGAbZEHPZeZ9ONLmYBXU6lf+ulU/P5Dvo0AMG
E7v4srg2DKdbCn1Yg6w4FVWlAwcC4EfnlxY+BQ4Y8KSdnh3n89E634gWjM9Kxrd0J2CU7Xx+7/j+
eoVIRA32vABtLZkUvswdwucZcPl5JeN5bKAE1re/k3rnAYpEKB32r6pQ8LjAMO2D9o+Ao+OhmcsD
TgsUpHqrun0CMGyopVFdEBdxgO+9zCyeT5/a9793TSvYPZ9IA1vOIxKRc75/uH5uZFW4BplZChfq
T6jSa69Pzv/v3Z/DoGhMuF7qcv0ZTQE0p76lOmjhbw0drtJtpFP4FqD0YUj96Wllh7iC62xTDLcP
QMLt4rLxpqrWQ76ACEGPZ135pAKwnDSdb2D8byZ1+eY02YuyvIcV1O2y0tMCbJs5z+sFH2RlZ85f
SgtkOeTzq8qpTpVBw1WpJh5otO1unkgOsXR6kNhy9gTJYKyava7lIeNmBjj6DMdEguGfcvlyXlXN
VCP+TAdl7+HAuUmpSzh+REleE9olZGmMpEucBNEuG4u0egskSQovpLcATK9ej5kKlWlMUNrvj7CV
viuPffYR8TIJTg+9uVPKTw1PkA+KvmDBJ4WA1K2oPtqNDVSED5zS2SwGFsV7oqlBZOhH2214A1sk
D8BlxlJ6Ia3jM3URwXQSUXC1ZrcW/p/m8r3Ah8HSuKVAsc8zGw1Xpj+uIDGIRQnQH/kuUY1HIDnU
Ir3VYKpfp7yYD1+S2qD5U1Y82iwhCBhnNXZJI6V0WhSLIllJnHraDsbYlKw/FHQm6sSuY1bJEjau
Vp18G7TQ24a7OZnGuHhMvzHvpwlwuydfXBdSJOAc/To0AGqeYzXdPi+A6qg7wS5m9awJIIZFbc5F
iQZJKCjK1z6oMi23iK/KAf739FvJuJFUbjqETopyNrrs+v/B1byxeN+LKkeUZ3IyVNyFWFEMpCO2
fNaKBsx8RdYeTL9XWp8BgFp37ZPAkc5/8JvXVjkpDHt37uTZJBfwUAgmrNI9CI3ZZ8Crs5gCp7Wk
fmxjnwGghZuVx4QVRGRmFwLMXAfELuF1magUQ0BYVDStlkch5yjLUpdb/nnp5oJgLcbMK29vDF8T
ILK2l6hyJLReOJlv0isCWFK3Lx7tTYb3qGM46LAz+vqSVmkiUVMzJkbam+hq9kveWWCQ5FK1J5De
UHjkXZSo9UsoOO5G8gMtQTtZegoJulRGb1UR9FPaEhcxuJpC9OKWKrVbmF9d5I99wK3DORwHGBva
ObIcFmLz5xnXv2QlMqV2CvkcWlsGm/fIEwnlCKxIeenmiFl6eza8BWkgYNpxcdUfCo+9HG+z11bJ
DusyzdQPGsAmRW4f5GGGWUmIXjsBbe0oBx1K/Ifm5iftiQ5VTxe4ChxhNJA/ihY6MADZly/OdqPe
LUn6YbfXsbzHMOAIMcKZOsx3BHhs0ghIN/sTF14Nl8AMuW0xL1ArioLHKArhI9SFcf/rLWQF3Os7
dRjiVhj48EzgF1oFJ5peV/fer4lusqrDxmTmNbSVwkUo7IAnCiW3ZWTuCwbw++IA/GDBPz1beDHy
JBZT5sGo3SvgKl1bwdizqGmHZRhnZXs7yPjjov3cS/H+xidwUU67PI77vbeVgYNMNooIEU5MKptW
5FWSFgsKWn0q+CPMljiYwDtsD+YthR5UI++ajzn4E4FSO7zdvjies95wuNfnva9ShFatPOx3PTTC
3Q+nFOmEGnELq8tCaho6p7a5CS4nx3l5Bmv7nIfHUAsqlhfmQD1aTax81495wSWV6pEjygwehuNb
braCR8bba5uyIOWkOZ5UMx6dmYIqC9Id7/Ksu7T6uEuIDrPlFijNEOZ2wSsPCfK10w+luW2Y7W13
ANaa108Ql2HOuzXdCWl758MjWTf/9tqieFXvug34iozBNAxWEEZapDg1g28nYfUGhz0Nu8iRfhXM
EjrJAa+UAeV4cVNvJbm5DzdZz1gDBNF9LFHGoV6C67i25l3Yj0MNizQ9bIGMMv8jqq8YqOmkeZ9t
9XlCBGesQzUCRnucRSFRheHAFhaMHC5uNa0oWslyf5XYScjXkR9i3Ibe881rtGQN/7FIuVTWAl/x
XtvjRBYiu6OY4D6CkZ9ZWK+GY9zWZ/rqKUNOrbLa+DdsbOYFl5I+4GC7KnWm43iiQ7q4+3hU6WrU
jMDLmaNxS6yyPtkLLkLWd7u9Do9qN10K0HHqxW1fYMkAj28VqPu2e6URbB6HvMY7qqUW3kTo5cpw
qQiLyt+2hEl7MWGHMCnecJlUJP6v0rO6m2JslV336lGb6NbRLR5CourdJfY8TpBI3gjg1LDCM2GG
VHcjtSG6ccXSWnsIj2Dw45TA6dFGRkl70FWz5I8Y1GCrBbY9Di1q/vW4y4+XIJfcYofhPCfqbLOW
0Y8EXl0+fwB0VOH5gU7UhMuWVWRe3LgY7WR5IlPtQN9dEayxuZJC3quAz9eZO9DQ1pnrH2V0Jt/y
pNCN3kS6quhQMjlm65rnOva7FsUQHI+Xc3cMwcsfKbcgyBkJN3Zj1abgfyIB+2zF5iEEAKcBq5Wp
gVGUCzPcHymEP76Tk2tbQ6fOIiRKjVbOsIPTFcd7geYOpIIF4dlGdrwTq73rABnhaLan7slQ4PVY
yjI5bDBnAUtXvu3FdLNIFRL7zUvbSWV44rxGnvCyyPLJ/p8Xk0pduyhOUCmtV8AZt4ym+VBUT8kA
+xLyiUAGLd28UjlNZXFFMfKK4l61jgwoRubZsKtww1OcYWbCgiGE5PUy3QNy3n6mLbnlo81NtM2q
tZPuzW8UoUxfV+1aTvsy2e9OD7vqTi9VcG64sXo37CXdbdJ5NOWyt19kI0HOL+SBVkj5mo9aDnQO
nNhfAHjtFIoScW5Q280ws55RxwwoSaT+F72nWDXRL3FtDsxfIXvhTOScHfKG7fbz0AF6QYAzXN6o
gUCUvtXyObBVpMW4Uq7Uz/Y3jz+NyUu8VpA7BcTJ2N++Q5qVIT86SiRVrL0T06oRx7f1Jls/zaWN
+Av/o4bAoKKAAhr6DdqBo8B9DUbioi1daXXhY1s7LI1vtEJUAsMzCb4LFbJc14L0Wtti85l9MOH4
wOU9KB9Yw8BroYsvnQIrTdZVP3oopbi0Qq5En08WzZBN7Q9p0Q3NIPvf+ih/OIyYtbcuMU5YB3xL
mhpgLB1gfBnqr08wZsWxnWWZMJpfTXD7pki2XD2sHQ6LZPlIQ7QDql9E+xqzHI9M3hx+NWc+7kP2
EXoLkJ4ACsOlbs4Z9jF2DsgbZOnWsL3FVICpl4s+r6WEY5olNw15bOf6mev4e3OG60b1ThCd3F98
LT7luib/13ZKHyJJ1NJo+DxUGWPKQiidB/wk+1Cnb2kG+M13a+IPSdmjC13blbO179pEd4ER3Cu2
YuYq+umMHLkg1O636zXVbLmVRoAKVmRxoHNt/HimGjicmtaUd2yPaiZ14aqqNzbW0foD8MtU7jI2
sUhDsYVUU89x6EYqKoUWsCoj8eEgOcezUEgi5oCgb9w7zktot1jX6h4c/ej0moWrucOjwW7fydoG
ayKl00Q+AUo+ZYrdS0DqfBdaTzrp18RmSB5XdIzW98uzAedwVflkJMZ7XVbPbng6s0qWyhn8KEfi
zt7zfaS2vE1MfUIs2hHfUcnDptqWlqMZaUkOIr157MtCVQaVbfTug6evUQroZl1YdpmTvn+evWCP
Q7ini/wznN/BTGoZjYa/ut8/WVTPyhrkRDU6hSK30DLjeEqJqQMTZJtnEhDIBuuCD1NsiFomLu3q
tT503V4aQxILQj8NSRWj9NEtpxhAfqUIOFOxNy4gYqCZzwDbIuDgwnaGmfmqmCkYVnDj1E4oLGrW
ARkaMaVnLUbmT5kz7kk2NbMXp9PoGBkBdOcKUSer4QqkPp4v/1XVwg17d+qPv0TNbWW0/nSIHSpN
YFLP+b+ynenSiJNJRZYRCQoph430g1G4wQblmHBCwF39YB2VOJfHMPk4OAzZro3kiO80ew3krCck
hec9JAdMBG/4RiuJ42Bq9+Vp1MTCwAFF4b8br2T/obKjEtzbT8ZhmXiDYSYtjIiSxPOmM5GnlNsO
Nk85ptk45giaulMksosvOvoc8uOpAT5D3Ub3VUjh2tScW55TEoKwPdxVT3kzH3NL/r8aPqMH6Wv/
i8yK6jnZw8u/5N0DNQ9mMULv4zp7jDNhE5PSmRLhOuq9BO4EwJaDxCAlp9vMWBVBjphSPFGpDKa+
vJKQy0+XFwVkpaMiUX7hZANwodP7v/WDJqv28KayTKNCF3kP/i+0xGkTKVNsaGS3xM/9BKmVUuPE
ugjN/qyyUE0GHvbpX8ZyhIKlye/OSAGMfzfzSXe+sdm8m/fX9vGdR1fqIkY0ZGs/400o6wGnd+UT
EXOHOIv5THK8ZBAXrvGvNg8HFQ2z8ayq1hLJFWN7lrN7MbrPbSjvuCJ/oMOQfDKDBbcdl4eogmUg
jd0A4LFDZ4JaOhmGiKvFCBE/70Z+c5DaW/jCoyFVM5ETGxc1RoZ8gkXPGP7FQtKP8zXYPIMimNtU
Xf9f664NTW01UttqkxBctkkeWa3KWQ6lv2tG7aDu8oBB/MaJe9iA7opnZkV7PMQK8v6tqVkb63TM
MrpCCLGOyx2X0nUdKNjHvRrMnFPTC1+/JfpaoCN92kcF7STQ3By9WMguBMRhrMdpvxnq3czM0N5w
BBye+K+ZpHYR4YgAsg6r23lMnJo6W2wkFpjlegFIFVNP6R8Hgv0V0Qglyfzoig3ZFlWMW4Cab535
ZxgIi/8p0swaOCM6J7W6wmw6tVSTCmPdHJT7fyt9aYQU1aZmJ5HvVYKigGkgT1zuyejUNGXYmMWR
IpN+AIQIPKBlbC870beU+6JRbR4+Qsn8JQ4plz30GFUxg1X6ygBd0br5DYb106vWIj8RLaYuImJ0
9W+l4D+co5l7UvnbwBH+gU88hsOTQdbjrYIp8lfHmnlnLGakXSQE9myZ6T7T7U+mv8DBDpth+uKD
LE7Vd+iLB7h777u9BwtuVLbJG8GaQYT4a1kDQ1vBTSLksWb4Zb+upQio3OOYXEpNWbU95SWXdPCx
EOKffsK7JVRZSKjLD7xs6TsUsZeL7Gge6FatQVqojd1wUHtRnPLXAp79AnjMp91TcCDlglsdX7zk
sjMxLHSmdYDfVAH/w+r2MParQUrZKyHxDlpo7ZjUYOrx6S6+g5XfdbYM0GDGsU/lzNEXM+KqzwT3
KJQmL5bg6bWYblVYI78hsBdSKACjKI671T8bNJsZdF5TPljVN7v+MfKZlQlih2xosENLsGuNYlvo
O1pn0QnGcvGd3XvSfk01fSOMNg4I9dgPf5KAbu/fiw9/5bFscEtM42xpUuueLdM31h+tz6rWYFO1
aoIqn1SEK9uR5+hER6nYaV0TNyBlJrYc2o+sXbXQCX79jVsk6tpz+fzUnoL4hZZK6BQPMbe2j/kL
puYr0Ucb703eV/2ZaABbJ7o5H2dLXjFdYCyG3SsoyXxzJ+RdmilQDZyCai4evAUD6ZDaE/EhaWbb
f9MFmATYD/Ea03tChN59fBfUjblQL9eb7IJBlYGMOQL06LIsRy8qe0uWXVjeMiJyvhZ1lvxrPjIT
VjrC1UWmd/saUuBPAEaQHfztDuU//Su/8fB/uIqJhuICC7V5ZW5CkfyQkx8P1jGd8r726qzsqLvG
6CQDwlBR4IyheffCcEGF2+wB8Xx6OEN4/PXlso/K0Q4Z8FfNc1WVLrmBa3q2VZHbYzKcGJctXRCW
aPFRl1oaW6yPhBKE9Bbm8JQRy4Exo6/H6Hi6LBJA+f7S+SPcCjC5zjjBS0MnIo3yzX0AQ3pVM6qZ
8hyqiNUc8BnCn9cVEwKOJe/Mw6a+4JVTor/5G5bHqYpWFImINPZLEPIoBONP3HQW1YJprx31EtuI
Ami13T0PX9Yy6PADI7c7MYM7+RF5xsux9TcOYZHunIys6MtNW34DfYTcWZrNoz6QXRU6v0mkq7fR
0WoIj+DH7o3Gvh1EDyOt+/ieCpSWej+HSRZGrEb+gPBrygbXxv/Wd7gDuCSFaMyAYdSwZHGF/jpY
27iZxtzySiZGNJWpdo5+40wGJ0EK+1Mh+Z2t30cU5diIRFurGUNijyKLFKM0MxP1P4UC44/BNwgt
EfAvyvTn2w58KKHfRJKBwm5zt9eFUcbcbEuQo0JWBs9+rvktlEjvX6b4bn1dOFbv8Wwdu5BOqCTB
t9aB6F644r1R8KU6zSLoFL+pgA2E++LhrKCZinNV+qU5XlHKC0Cj7InvV0oCbWkoz/BbU4D61Oth
UEaoYL3dwAMrumORaBlymk4WBgzsfmVtn3p+ePa+hN8JUXwtCmE9klaX/HUXe1howQcv/qfL4d+f
INHZHzeYOc5JhU6Uk8o+dT/YWcCPEpmHh3wE1ZeyqYlaixRUv+hY9WUCtCmipWR5t2pCjvL8OTIx
F2wTEO4IS6p5QpLdAUi/JYCstG8QCM2LvnRUdXJDES3Ibtijg9weadhHihFmWQzFw+g9mXpkcbDr
1Un6a8OHgX7JIYFZVhk5S05s/mnu985+1GyOZ1+dE1XRwNocaRbF2DvEuBVCCKviNDw3xGHBMwpc
/6UeQi2LHuMYhaWkv8TUxHZkyvBn1yODbGZGXCD5wwmtoUGYx0dFPEwS3Uh3Uqow1DUccTlIIgUy
piPHhyGvmMlLG/W5VFOepo+UQSU7ATfIrjM6jQYIItWBSKecnz0PwAxXMk0QE/jjLIsLem1sP75V
tD+DAmAHdKDn/W2bru5k2VEYQqe4xA1JxbAl87T3iLmlLosUuf/3A/jL2wkuJ5DpE/vhI6lVa9kR
WXYhhB/r6CLoYaNPGugEJrzydbimUqM/W02HSrnFz5ow8zAWBXgl8b6yArD/Kz5C53s+/pil3wv0
xVFIBT+/nfbhynHMy5l5fMnzHin4hEZ3ITaNiqa1q4L6B4cWYAWszQAnzz1HCxL+h7oDE1KNJbf/
EkI6vCuqRfKm65jIiFq5lP7fmDLxwJLXjjYLLpDNPht161CNqmG9buaWh3nShKAxw4uIxFhwCmz3
cHxWx7Z9Y/FHQunYCcNDVl06cvrSBrZ5XAfdgIFeuY3uJZAbfWLvuim0h/E2OfyHpgExeCU9MIEd
Dh9SyuEGsudjfmR3p4as3k9Mjox6eDrHwJU8mbOvTw4AXtIfg69WfKu+h/HY7jEIqbViHL71IC2z
5QvJfHarPGhsXMYmE6kzuzJ6vqghGnEDLs+HZaGcl7tLksZteH4IzJXn+kdUVoQiCa+C3oz+HzIh
4YFhc2xQn7C3Neq81pLFAB8FjcwwQUG1oECddBy1rHEtKSnfbkz7jY1QZTkDs5m58oqTRaOJ3/ov
ZrpmDeNVNaH04EAIjRGVEyHO1kuQU8mXD04XaZ93i9+cS7u9fWZJAUpRJb9xlSC4vP8IZBXfnMUG
u1n/TpeHwbfRwKoKxWixkpKAymsmmbq2g4AdW6yzH9rKAC47DxmKafX3RkN96GwhrU3ZGREuYSvI
u399+ovY2D3mgM4hzZ5KvV47JCcpnm7CoocbYdq1kdWEjYZ3ZJ7rHvLRGmMEn6G7Ewa62xtw5adF
NuRf2hzCt9IJyXyddfBHWV2iRceXPbpzZbVe/DlowZuV61aahZBWM0VjC5Upj2rZNQkvM+rNCO3o
xN6vw41LJZ1jCISTqEnztu3Pn9Hg5EEwb4aLy8OxkmYYS5Jzq+SpedpHg4bovXRB6/TzuAAkAqdz
sn6wktuBuFI1zn13vaPU3eBioZ/tSUqVNGp9+9UOY0Zv6WGJ82sMWdbstD6AaRQ+Tkr056r4eBjN
mYahGTLgWr3MaL1Z37mIubtuDFMTYNc6T/naU7qlyexBjv6ZPqg55NrUPljhqf+QkZm/w7ikzDV3
Jl4FvzuNIDGCSmmYQ8G+X6uYke01i0q1InfKWzLDp6pynNl6Q3Q1bZ8NLjrL+WUtSJuGdR47kJEU
7IKaz/zIOZnqPiRTFX7OPBfHzWRBvkPBRPdZ+s5Gjb5Q+C2NDCYjPPGLGbQ47od74/F/5Jq6ILO8
UH1IgpShRJrl02xZ+SESdvNlwGUygfHsxmwR7R8CzKIubU3jcXHp9jPgUyCCYmJlSXVFPI8tEwZk
4yfBywHGNXsmagy/xLmBqjhnlAmzY/AO3YDnoSrMqFZB/04lIGjNl/09Fc4Ss9cuToEk0ZXTohKV
AhQMhUCuBztfjaNDJdIlm5S6qjHxFn8FV3uUPNJQ3kGvYhjwQPOdtOgK/iEX1wBqeyku840BPUzL
XQw9KoNK9xKESlnGY4bdMhIbHoqEdd+tdVpwgc/iIMHRFwVn8Sh02RVVJ863ghVSxwNQSmjMrpp7
zM6Kgms74+IA6tkeY/pomgpYknnPmM/HvVI6JGPMuZ72e9QN3jqMPm1BWuDU9awMBRzZli08+SmJ
YfFmgNQk8G1Hz+d7MdGQU+qXwoggPAu3uChGl+cVvAeNAcHavF56c1LLiHUIQ9IYiaifo5kWQa3F
KP1uga5z7dqmflGv53noNfjEW4lYLf7qOxr1/iQPBSpTBTvLl3OFkSQMKepoW6Y8Ywx28pEbrcpc
MpNa+tDeI5HYr/ZKNg2FwnlWFrjkmtVFtfUmzU2n7ass1hH2UCUJFdCc7Ts6lJufvOrYpanrPMIJ
7X2YBV/RpNMBFj+GKRrr5ExChENszhiSJBPnbx5hGP1sPOXAP2UrU5pte/vVm/LIzqcPJwWXKsY1
7yzxx+IbIMr4Fxwlsf6tgjL+uS1c8Eo2KQYM/chskW+ULvhiFhOVlNlHuHsHTMeuE1tNiwgLecFf
gxBqRilqz7uNbiiM0obo5oN3Zzd8S703jJirU0ajbvCDbYDZbFeF9Beic8covLqWLiiFJTlXLeB6
dIS3fqEg17x5YaDSCEtkdofpfTdWGndT8vE85SQefhQNzWBs5I9kzNdngr7hC2aOaLz/ZUCXNqE1
T/Ejq1lpJPhm7c+/VQ3PlF+ICzIsZZCIT9FYx9WpcMNRVb1ZcCKq7rQRQI7Du7pRtX1qWzaQ95jA
SqH4jROg79m0WMMiQfK0nP62fvEDW5sXc3PY/KKhTGQC48VGW8+EPjn2dTFghzWeWpYJmxXM7frA
bwO6fLbZi9b6J57j3PjwJF60DeclVE4ev/NZ1Ssz2LGNz2KfNtByep7QX5sgrXFZvWRSYVAIlTah
CDPrdPaSNYlcszsmhMas5WB8Xk5kOV65m0PcM4Nf+XRjXkzgHDcMWxWS9U0qDRuTRor2i0JBCYzi
yKCahxkP9uxy0qMi1pYy0QvVl1Rss3s/tKkVPbBtDkUuwtT8kT/AIKj+Ic08JvYfD7tGWz+8W/le
4qFN6214Qc/jSNKOB2Mbkfnnalxcyg5YZKLVbomHiSE8FBl9La9z91GWdp6xKIf96yonn7ADXlue
DuWqjzAKlyMG6WVlZYYzMa6R+5KYWVUrE68dPLzfj9VvmLAYI3QIdG8uFYorS51QBHyjfrUc3/54
oVop8H302wMvE76d3RTc8s4Em6+NFLNfUmMPU71n6cvZxNqIoHJli/8VV2e2waRInYh3ExDxKry2
bAl/5+q91XDufPTqLTr1ddMX1XNy1lS8EzW1i/yEh140/AekILEPhafA6pibSeobtYmEVImwlmaQ
I6LxCOxgs3+H6btKCvasYAQVsobEoOOoOSijiPTMXV+JlRoIbSIrE8AnEnsHyeo7WpNiaxDrkQRO
NzYvd6/aS2oAtnyANe60yiJ51pNt8VuQxG74bKjuzKVL96BFIjS1n3IJrr/XvCA+r3HxN81kiJPO
OH//znpL3vtDFgPnaWmFndB+O5FJKztvBPivXjn2Dw5cyNbkWpH5CQ5Yh1c8ja9NOrxMOpYJtEdn
Eyr5Lc9DbBKezKGpxGGbYhFcL1VrjLRWt/Mz74Lq/8n7gja7vBnPkyPSD58q4f7FyJgxLaG9pCIz
j9xjlLg+bNbszxdBq1FLOdBCwBd/zGTds58JM7FX7nHiglF+wEzeUaqJCvy0iP+oRxmDAdklgebT
OnPK5KchOgd5RtTQigP2yfkJuCJgDpYfm/NinPeg5SrR8SivTWsIFbK5HVrhxSZmxPP8KIJWMmFF
axyptboCvg6B41Lkcp52fAG+VTGw8GQy1/b06UEUuhvqZ8vISjU2v6H5kxV2csVWfDGYQ0uyjKfR
/sJR23t8cCbuKpjD3DYjdpMvg/auiTmXKHpUE3wCCoilWYkQINSfwhwljUwbmArR/AFO9elByr8H
4iXV120xxC12VgEdaupZOaixoqW3cwsNgV5HX3b1uSmf2jNHkQ+qrom2IVJ0cxpM6JwrvOBy2xoi
OWzcqEP19NpwLYDbwhbjn2PP2irBbutwWFPUqEA+KKOsdtEa0FkPnaw8eMvkC2D7x+b2vdaFEpJF
TNCpFbD1x8pUq8d4M586puksvJsqpw8mP43+hghuE4K4lu61/O9n04CHGlMDFFKFtJTbDVwITavl
ldK4qS0spnlihf2hWdr84Uj3Gnln/8pg1GtidXEooXU/iNMQIcimh35JsRc+/8RtZju8vWWHoWz2
F9dF7Dk8281ttZ4iKt4j9zNUvxIXte45M8dQTIfnG8h9Bie6AKZUgG7txAJsw/MQ691FzsL4Olcx
Ak/Hy/pCaJD7Na2tCPyPr73LGlQB/4h5KBxczvXQsRaXrXaNPWWVlOWmxRUJCXYxLY6MWOoDPaGE
exBoy8E3EFz9fBmqPg7MiGjKaIqDq5Z77xUdtddrdUoEVxET/d4Q+3QZgAVfvjZlX/rdGwXqiFFh
eeBeENYpBcRllYeqJTzwrp30HHCIQF30269KRyUlLqG4lgXg5O2L8VVm94XE4sqDb4t9WX4DL2pP
TKUKUhhkU2Y4LCTYfd73PfHfqFogYyQOzNRsV8djI4yYvkd4/7TJ5MyP+uupa5e6fn0wSPp/soN0
vRWJzNRXBIEXrAjyqP1vQRl+oNV9HGbR8bgwHw0DCxQtwluzQQvSNO9AG8by7+WiU/eOVo8nxp5X
eXM29yciIfdTohrz3eIA8lJLIrErzv50g9Cuz3+UD7SQNCF+SQ/V2CBYwj000iRlH/kzj6MR8ufJ
nAiuVrV23DZJCn4BcoLO4sLDTpOHWhbF8ocAAo2fLHg8TF4f0rvoyEl33/8OhSQ7aN2nU6kjeOnt
KzdyDdU3RHV3DrTEQIEHuH0J/DMIikS9vwwCXCA4GZPX9iTKRg9TovZH03n1OEdY6HgQ6z9gLe/s
K1IMne87Q1DIGGsJEypmr3iq/pArbsedDIJBA++ySY3WmpwqyrvsDD0X1EoKa2H0iChe8jgZZdSp
dQF4qRfg1Mks6qbiIg9QQbbo7Xo1w5TH5+4BDeNzBnRISUVDfXczFHm/YE2dnDNm4yCeGreVVJRF
PUwX2HjetgUSVgiUYPsnEBGZ7WGiEGF+DniTyD+Bt8rIs5X8+l4UgmMW6kyrXWwpXkQgcLdNgndZ
CHLXtlhLrB2bCQNedcKMUxtSy9GxjnwkUr9L7DBFmtag6v/NW6gmKf5i40us8qEgpdU3rDUR6SKQ
AkhFC8/46/OUgBJUqwub9L2F+seYUMDOU+LYY/pe7w9kmVQ4FAKQS6tT7WTXKAoTxYHEN5fJpZgj
IupGwDbq9m+rWGaNc6T2cmvcdJJir1s1LIQj6izWx1R8Zzrh++jrNrHvviABC5VYNHHt59viyRU0
orQZfKSV2oKWhIAds64vO6LZXtt5lZQSLEet8fNZt7UKOupjgKlsiAUzcYNxqSV9py9CRSyt9nmw
IVoV23+a5yv3n9LFkccE+lB97KLMYj8avCq+b90NkPC6eKVaed3zmrMePSIm39vl6bd0gudzxjvl
/pxVWnm7GmVXXymotQRa578iZ6vgvbzyk089/O4N8Okr+1HtMB1lb17PcVp5kSMXHTmSPZKzXCxb
sUO/s/uzH6AoUIUZ3SiGShrZ0x+CoVYO0EI9Cu64na20b49Ixm0dEJyu0UX93d33Se7FacTXp6QS
SCYS+thKTbqSFyujy7+bnEjEais+CjO5E0T0JTbhMPp4gljeYaZsNA+w79ph96ryziWsZzx/9ckR
8LoTcfv/TjrR+ZRcikJGnh6Z0rz1a+k+prsHCMkdBFwQ9VzdpomeYcfAXtfh51YGDUnyidvmc87C
jLyWFsOwGki8ilBSnTIrjUvV1JxXOyYIY61dlrQgDFsvzRg+VnrFxB56Ola/W/G6kWJTzYl6rhZj
P8IeMZtVctc6WMsc2POjdP3u7Ev3s9c2XvrtwGFIWO+7wgXqzpLCkXuOWzsQ8W+eq9y06+UkBwzv
Rega2p7S/x4zmWMCqfwY5zmAtMsQ256nEgFSIJljE+F8QyxpfIjYcE48lRXi9pOrb+En+YupVHIv
iAAlQv0rIjdVIM1hZj3sy3S/jwKLolUcR/m4r2cjyUnEKg8T+x/ijnZWjaPWeFoKbu9raUv8RFUL
OI4IM8cbDFPisoc75IN/JOpK1OB8yx6rXU2NNCz/mk959EfKJx4ZjPEjHuyrUJOyYMgOyfBnAi7c
O0QoDytQspm7i2HUPyC4N4z5rmztzQXQe4knh3nvDxasBhsIzD/X+/nqWuEHz0CU5MQ7EgxSqZTT
bDfHQTsSMBRAUW7Cx/jEB/IrHEc5gx/iNku6AK9UpixuI9m1Hj/keDvpb9euC4r7VqCijAxP4P56
Gg+KaAXZ3mff8Sfxx0QUYfoTApvFDKL1H9JV/fiRbZr9s9Xse4g/onHkKZ87/Q6fD7Qe1A6EMmtb
YPYviUXhGMrCfP2n4S3WhkTMofKMPAlxaqDjadoVng+nuq7xxp1a3ApzYzJ8ICLWvMq0MDZTqxVL
hQiaGhLPa37lxNeSNGmOXd7lhkff1M9ZzEprACBG3ohMX4JLMbXy+F0R3jRZLL5drXRIJ1ORKXrZ
uJlRGDt7RgwuMuKAJys7VpXqAW3EeUY3Ijqr4t144glHMwPL1KwRWRypqh7+Z1CpZ0uMDQznJ9ye
mcM6/TT+3puLP04d17i9goOPaHSDS1qnHGHBxnq8fdBv6U7MffaHLL0puKeThSCYFbcxp5ISToN1
0FEzI47lYotGT3tEmiYAU52GzzaE6L1RjyfyN/gsHKjT0x3pyP17Jdjuug0yVgTT4x/ltS1Lff7Y
KfOa1+GDvzuFVvl1yKwitteUC90xfEV3h/plmmRyg+cTFz9VSejxhKQsoYifC5ajLWiSjoQK+J67
I8MNz4zNSfNckxn1Qfajk4KbBX37tniOHLdHLQfBZ9s3IvGOMbvE/HWtVEk8Cz0jlkCCa1zwHNHO
SOXatPPZ5GCv8JfLLm4wjvBrWJFiNTm5QsOmlOpukDGYR364VIfnbLJ7Abt/kn40sFrUt6Q4ccBV
a3aRJL+W6yau1+BdRZhhqx1kP5ODWoGEEchtWJ9rqYenH0Tx9sQjtx6hwgvXlcr5yr/bi2jwq2oA
qf9jvEhCJgcwY1UNUjycGHja1i5RDTSaYEKAIRKlnWzXJB2sreZY6J8UxfB4oIpeOs5Vf+LXu3Cw
aC2UCcTMoBq2R5lADh3whp7YVGH+FxQcXe3L1V/XGgJ4eYOY+aUqXykrqGsq7GouirjigiWeuKkF
rHRees73rxajN0J7XLpVAjov66dwKd9X7FfItjF2Z8kVimzQ6gztFDKuP5vNKylc1pWJMk8SEdHC
/i7aTOrjiYlVOvosEAwGo79m2v3WVCnDVqOPyr6JNBfU3dnL4efK/dkib80/RkIYOmUMZ4lPTKSP
7rdKeVHoIYNQ4KcvPP7LMk74UhozZTI634kpwEsZ4VO9+6WEIdcAXjREftKY6T6JozMCMaxDlimi
8Czoyo4PDcu02MX/Rj2DN42TC1svmxETrgoItgu5KrESSH/ADs29crR+Y1oVkSWgGiaoV0zIMFUu
bmq0Gzv9w9acSdUc1iwXkKCvGcCVJHk0UKmutcSC0N7rpOkK4o9KjWT5YS4JdtUCKxU5gIU8CT6y
3cDAfgsbJqPjPtVlIm+PcjQ3GcSqn2r1lOjaCJcfm4zBPnMd/iVeH47MVkFqKgeur6lB4wcCXxWN
KxRGc0pjp1/i5nXsDbI0bAxBz+NiP4AklouSHwfZiSu95E06hlNcEpTY8UBgKFG74sELMYQ4/RPu
+/hHkv3RWnj+rylc+qpbVe6XCA7Jdu0SmCstqC83D0Maz0WsByWMsSciiELsARUB/SJyQk8hbkfT
AfcUXlaxK8Sc2SYmHxuqRK7d1eMo2isJDkc50tYLLqJDw4BW/XfbbRT4ByIl7i3wh6Fn+Bf78+5r
anrxH9z1uWS20zSdX2zdy7q0g3zloQ7u3N7K2srqmGFT6STvVEylssdi9V7g7E55/osaYH/q6NVj
dGyjPyTf/sIW7nWtzQGOBEQ2/tbXKdf/x+npqo1Kwlrp/ZDCZWoo+UeTIDmdlIdkqDMivsunGNVA
zHzsZsTnPF5uKXn9SukvnaWNbJtAp+yOUvhId4OBWGC3zNj6OqUIJqQ04a/Q9rbHtfn83SpKwr87
NkevLzjpu+554+Q1el6JflHJWXOM9Aqkizqkw3jpxpuuMBpJ9MvCynvQb0g7WvFY4qyZnI+G3xpZ
uC8tbpQicYwk0dSU+B0/x/AIGGYptWX0Do91zvVBs+XV7rFvf9U8othT2HOave91Zj3mU2FJ2c2R
0WPa6Bxsr12iM3AMZL6gJo1fFQ6OorEAM+1+7tlOkxqeLxREV+hwkqsQYSr/uZQFOFINFCIUAm4w
gJvVifNjlYUU0zCUKS2UMag/QhoSKCjjLexQNQYJPtgCdAX7kAI3o23HfIbKyng6RxhZkbOrLC2B
u5gL54I3olIpCk1XxtsQDS7wEDVu/pEWu7k7m3dfF2vNqucb/KJ1tKSfLBYHBiWkTUtJRIMdqGoz
I8BeGcWKVDs9R8xs1vRFwtywsp3t3DV3jQ+O1bCsaBZxUiXUryP4uwSOExfJXVu8ruZt1jR1KgTr
0spbyLs33Y7GED5TIXr4MP8qjemrE0zoEBOgL3fLvN7m3M3zCYs7k6a5Hz4fcf1N7z9o9wnXuXR8
AWb4D086uZSPqDWHEB2tysQRQwMysnqGAde/fKeJzOdCWIO7TQXd8f6aKOTCcX9BjFnB/1wHXBv1
2QInNoZAGwgZI58YtKmWnzw34CJU0nLbmPuRDpLPScE2Kv7VitabAKawN4ga4XzVKjDygL01jGsb
DADcqcq9qM4VdYD9oM52Qzlxenumdg7g/rqwQmZZF/2v8oVywMIkWOnOcnMNhGxjnqiQSxmqh4uk
KhpDk0zBpbOU6RHK6y2B53rSrYXNlH4A5pQSsXnQKCpwfSpdku8qotxRhIJYmvCmwNVsLF4kvz8P
3V6y1V2veXCCbEGDBgouEGJC7KHcH20tKYtkDSCDlABbglhmDOf5iVe82bcCiBeXyHH16PrHQMhW
PmPPvNWdxU1Oo4MUJKnTntq5sbG+MBuy7mK2sgY5O4/kDhI01oq3KZPT/u22LlF0BhAVPpVYOsbR
CVFR9x80+8Q+t4o4trCen0/kJjlgM63Dk5Qj3A3zPbOLSjoA8dNJTjwqM6hHNjv6JRTeL5fxokSi
Lj3LEshmxX7ss0MbILxo/rQ7PgXP6lss1LuBguf2/9EwXUV+pzoSjkXqqKrEFEIuz2qdYFC/bDLM
IyvBsRFQsKuXp4AjAgW/RHg222iznd563GLkTU0GQ992BI719LK2DW5JvOL3WyOXvoEjEv8vL93F
Y6kwcPReMBBRcu7eyk5iMpYU+WV021t8rXvokWiDSPu+IRG16AyAg95fo1CGT/sFjiAEvq5+Tod4
xuOYFCcx7nLf8SyJ7+Xo15G4OB/py4UjqeaP4Ls8awjmOETq9jx/F+XbCAu+7RPWnZlqmswyCAWT
junPkEmw3RzO5NbMy3YL0fPelFdAYnSdPLb5GZxWSgK7SUDKC6/myA2hXD4AG+4+KX6rcJ/IqrZD
606wDKIEG0DmrMZmn6U3xtUEi034piCnvT66rUzqEyoH0waQgwUaoKf6+zRNSktMJ+H91AV+VZqt
92EYjpoxGBBeJsu3A072zcT3hBZB+O0AftGMvpjwAtsBbaIUAEOI8JFnwPvMs+SQO7nSBVCHpbmE
ZXlf+MPXcxMPbHckdXr9n1WXF0XzZzFSlO2MTtbg0HGaR8S+2cS66wXTO297dpu3FPBa++OoOSlR
N+1ob85xyslX+7oaPAn31aGzgsuxv3zIwoBJoRP7/LaHAcEGhUl7HGFa2RCTeq/hydwMM94zFKff
LBZ0ZuHfE6yGA1tTGVo18sJ5ib8avlkTvyu79R24o8wnnmrt1FLJ0w0s9Nd886eWy64q0tWF4wup
WeZR5/qYbts2BBssNVDMZsYsh34Goh3S+CeCksGz/lRH4P9KCJlbylbPn/f/RU9dilSC4LZKyn/V
+BZAhnrwbMZCw495Gy1iRP4qNQW4VEbEqhCkaDGAPS9m4rSmXRSKmZCaKKmfxgZPi2zp+DyG5LQ5
08MfcY/rWo63lBcFwrmqFj+6IahMWMER2AGzN2dfXu8CcUxKuhRCBNW7a/Q8VXi5i7XKpdyJ+3fJ
vl/1Rm6YUSSABHfHhd0OML8Ihppk7uBBWB8BsOkuLiyPp0g7pyWaAnWfUg3lyD/1+kh3htFLb/oI
iq0UhzIILuZ8CudLvNLsXWGQlA7P9YJuenJBV+CZx/ZpuJ0Do9nITQgTOYQ2CMG0TKD9N01KNDaN
s70gaHYX3ALKyNx4KOSRQ2TgpHnVYVOEKnXIAzICw+JlxPre976GI3mHYhLHaYPRN9EWCA6oSacw
wAmDOtKW17/1GphQBAwquz5rXTp/jSIIzZ8oL4KSv8AjEGUtJ7VXO7DKyeEvbbIg9H6C6WNHOGFM
hThia/nlhpZcMEmowSzZU0ZfLxHV1Fye9Eigwlxvt5ob5T5MTgwl94UAaiS+lN2gYMtTIGUG+zQQ
LOWrwc8o7c9R8ngs4GOWjeR3EtoZN3Hep1TKWLqM71IB/aPh4EDRmF0fa+CcnIcu6yHU+RiEL59M
N0HKh1+4u7wHWqcm7TgFfN+MbTJUqp4GHjbNMH99k+aPC+qY+iY87DJSUP1bcEGEVvVkyFLERT2k
3NzFI9DPg0dDxbfyUgRGHS/v+6OEGWdTIeuO2a9TiUY7Fsi8n2TkkkpiM+sZfPPpUtNvA0YDIgwB
xraZXQI+zC20PpxVeMYy4EpB1iRup6hdUqRm8FHCKfJ3guUxZKZrFpzEwnbLUG6nOsen09/QwaAC
fVZDpph3mpE9OMpbyQHt+Yq3OrXZAuFzpsgQlJctST443mDIYkCxf/r7DOcL3xnn9sAtPZWJRFME
wiY5GXewcyszXmIs7i7H8L/6y9t/M87IgChTBQzw1WlNLAS/BmNedP4iqydtL698w4k/lX77Q5KK
qeADhC6ejakxYg54W6se/oXYC8prXBIs4zk8qLQQi/tvRb1ljz9RnlVidq7wMPZCxguOyt4BSBM1
bcAaTtwF1/Nd5OUObu73GyMoZupBfGokyQB6aKNh6iaxYGQ1u17jkhwOoV4a4pocdqUW8s0BtJG1
nEginGUiRqdKm3zMSkTN+DuVobh7xJywiigF4JFRv8Qj0rpTD3cAGcUZMbbTX/+sI6u/jKXa9R6o
DAFkvKQQR0++ZUXJI8tfgJjw+R8a1CQfR2TpNuVnB/AMJBrHJudxJw6oZm/T8DfZkNMetio86XRv
DskUAepnF8q5uzrD4qibnEQG8ypRUOI5a4/abQq4C6HtyDcedjyUa9ecrIa/AgBNiPOTBcZv/Fxt
0Yxdd5B4fMTM2OiDD8SNMa+Gz4my2mbeWE80MwKMxp7mk8r19485FYacClY3KFhhRy+GuyeRxtTf
XM+JY1rdu7ZjlreIEDdFXY3WhWC/VnqiejG3dKw+11Ko1yXfiFBJT2VqD/4oavVhFnLaHdol3o2v
qT89O8rlef4uTWuacLifHTcjnY0JLfEtr6Lmjo9sQS7vNsM0gT/WIbcDTGLP2sfhI9EBc10q94wV
RxG5LtsKxLCAfp5D/29OSGOD1GhXyUBEf5gHz0yTDol9Ds/ClHFUHeYzdcXT5vUw8SooIqqA9ECl
6LGfrHNrNL6qQ9WMbGeS3bkkaJ8B02TqYz7WAVW05FUFxASQQy5QhXHAG5oR9+Y5T8f0pcSfMMFu
Tj8QtvWXrtqzs7v8A5cbPFmUcEb34zwZ8n329VqPeE+YYhmYOXTtDk2ifAgyVDvG7Us3/vSU1Ypp
9vfaAI7LZ/dSs/5Cnsf3/FO+/7FhquJqKRcM459mNX2C8PMR/zr5132yttPoGEqPFa/QFEsNrlZr
Tl95wF3bnxZ6prmk7exE/G/gmNvvMFLaHLGEWdUE57kefDmpMTr2mx5GjB1WoFruSf3godLnHR5l
cNfrrb0o/RsWKw5T6NayluFTXW609k937T/SCc3Jx7WvZUJYttg9mPhcdMbGV9OIru3Q7wDolIsp
yUhNYzic0Tu8XPHmJt/YWp9kLW6gXaF7Ckjll1+cmp7N6pmZ1ZSl68QmJy4FDATTc6rf/TgKBfaT
3uVsWkIaZp3AuyX5J8z/oDvl3ApinrflgCf0T5MhGwFg2RzNBB/dr6scwoxGTVtxTNHo6GHBIpWp
Mc2UXCauEFhXDDwfG6rQEfTcancEGTqnZpJeJGOjQd5IV7cYMfjG0EOV+CafWA4KrNCX86UXeiqd
7A5iRCVvIOjDjK1kptYkFIGWaticVrPhJFlC3TNdzEVDNyENDqL9jpkZbw2LoeneJORMwOrBkQwa
5Naqh9oR5418zikSn9hai49m10CEFMCiAEaveqd5G5ZxvQCF8WIikqveK3dXG90RhS36qQzyLLfN
Wx8nO74DeM2QQJwV1FAAX4OMKYMjRKFkFf8WaiFrAGmIpmleAxxV7O5apKVxPNs2xKzIarObMo5I
kekevIhnjdQNVmnaEqw0P5xQ3b5+MJLzqs5Wgyj88Zuehi7/4GR7G/Mb7DP4fwm0ahy63tlDqa0o
LGH/0TYrJ38DobPLcjL8U4yc27HgTxUcTDLXOo7wYTemfHkGxymkBPH0cxlbVkSYKKdDqbT8bAr4
f4TH00Z/MYTTkx701kagCHO3fH5QqE0zy8rGUsvWomRTbxOp47F7Zzhs9igkOS63d8XS1qJ0uDMM
gbY85omsRp8mLsDXVEkJ4qhl/PjyYQrrl4dH7dYl8crJ17xlHUBe9SYzLXl+r+0VE+UvebE2gOK8
RQ/IXC/GgSO2gIQpNRchIK1tcTShAXNcZX9tsEKWsiPHlQ2HDi3cx0oB7tmzqpz8qLxXjf4K5gfA
s2E9UuEPwihfstT0R/cLk6yw8OvJv2jAB8a39rZhV4VRooRvnOw2NxigS79vXaWcbAKxuHjgt+Z7
c7Duqgq1c/wAZ8NhaxcjZ9sZ3mdW0HE8zbzBd5G3SmAfv4XbSUqEJDRGIB5dQMg3/BIz4tdaCg8r
D5x02FWgZ8HEDrRIk/9n+9Z24xtXmDp8Hs+Vwq0CDnFmNaajjSNoVxnCgNUnY7UK4dlNWZ78UbWC
xe6YLrXFNkSIecQn5zcbOjy2qWXOrAaGcdZOjRYNfONFnRo21BgP1eA9QXJqt0OdYdfi9gvAL1I0
fzaoAkmXhtaTfenVy55wPk1LW9wKKPxoyw59xkj2TfsYbodycmV7DQMytBP1H1YjijodASGboc1E
FbeNrodlj9UgEuiYP+DIVBx5oMRY0fa9YVyNnaYu+p3ELxs22kSoJ5/hau8ByVTZBuef0E129q1h
6cxltC5ASL95NxfaaocZeD75PvF/YxMdDRHMb1LnrgB744qfHt4AokZrjq2TamQbi8hYfxyhoYZp
kNXXoA1it/JeO88GT1OJBVZyco5tsf3JI10c6JoRMQARJzayBflbTZWE4SBBvvymyPnfAKNUUfs4
QFkczDhGkd2sTIoXczVMHs7NXTAQP/XlkV8eWDntjsCqT+DPptvmD1/LPOmPCpnsp/ipwF5rkIgr
FbZdE3hHK67cFTY2s6cikAOZlf7DNHd0uV49Tua8/rFyIAWlsNsKSnR4c7TTtjs0cTBqIN6D9d5W
ST0QwJlcA2TrMmDpcK1OWJhKzqvPxyvGeIqgN8a0PLrOCMe2aweotrvWHn03k01Q5kxFXbx0oJxb
44C+SDGkESfMlj2J/lSFob6lalZl7YBoJxAQM5uxDxpkUjlmwcxgypSkk+t6s+VvSkevi9aPUVCu
E+GzSzSLh/NGv9C8bHRJem1bFouABfpOwn7dVGxL/faPACbAWOGeu/3ikfYyF3P6rFDpM6YRsvD8
AcG4H+ORSU0HU9Pt/ZqBHIoROrRiQNzdDP3+UJY2/AEUvf4+GRPhYD8iM3wDyoLNdGsxyAPBIpw/
oeRw2Y68JtGVM6SdT/w5eKmwVtSttVffx4yGH5rPUC7PXGoxDTfxKDVCpw8SSRnBL5/Gi1rbC+BD
8ysiU9U0AD8GIP8Cvk722JfE64+0nLNa+4z6EflyW23yvo4skSsAZ9GIKrS671dG+gvkNNapzkCF
4167fiAGZFqNzjzRSXDsRPQYntyzDeugP/UgSDj12f1xrkyqBkQNBPLgb53csJt+BbUKhxdRkH27
JFhx+jJg5rNmxg+AXwnm2FY+9yTkj/Hldg450QKQRmOzGsjJ5/dbev8ZOlXQTQXREmLIPe0NMwe1
YJDzTWr5B8D8AFNZAjc0unmf7FqynjZDetmSAwtg4udf78w3bL9uAn6WaQWSjwKyr1AmUewYVUUG
uOJA5zLoZ1xOFpwk0tFaanR1eWjOnAypv2q4uVSb1srWv863PRS83qry9wHLEyy7fL+HbwIlDAfi
jECRmv09VmWBejY9h1cjUMfKeZOzMdtirFKvkD4WeAu+QPAy+FF/ZLnKnFUD75nZmsf3YTagGzlU
m7vuS+mMfCZVR+fnRm2joRJpkX36XqTXwTU0VlonHasA/XNRqnzfyEK/NqMr5SD2iz51Th5wpGwW
ltVFpst2lmQdwPc2lPsiaUjQe7ARJFMbz/wSt2bQp/sSfjf1rfU49URdBrvEAfX9iYFk/yyNIKcC
brzOeo8q5kwzd8I9RR8jNN4ej7KtclKFA1657vPgYUUCz7pLzkLFa6qQ/4R/j5OZTZFr9xgNIEjx
UgI94ndpgm8XX+iO1iUfEe1ri/ZLo8xJFey4aXV3ypbloxybyRqizhu5goiGyEMorO3ZrCtwuMP/
QuAH+YActcuVEjN62UO892NYAlh6TWsO3A/JrOcMoyuOmBLziAriarcjwgLN+PVjsD3esjkTxtTI
rcNfOqxhSBnl9w7Kb6WVDJaxnJPWWFah/ImumIHwc8iIBJH1PnHoM0+wpZglMFU4tZNOVHAve8UC
RmQ4qPw39MwBCC6sTiL9/wonw5A9LaqF3xEj0We0pNr4HbEC8Y8exiXXQT8YjHf65MCLjYChAwLs
zBKgLJXOnt1rAIZ9tZq++EMuuJBIvjpLOdRSTTctv7ggSmQbuRQ9h77Aoe+OR3ZQtMM0wybkF/PA
ToNq9rDRSsAx2CItFoE4F3SHGgoNj6zqwRPGSvLXYPmXDU4bvSvDVN4gupSdwkNbFUmn17hpdj5f
1b9ZaFDvieMAbtBCs3eKKjZnN8/rIgjpNbFNFPI/mjqd01uDnE7ZBaJJrfI6/2L09hkSa3J8aq63
O/j1eB5HQTmqZPiOq3yKiupwlIUbtKtHx98hYM2oDgAoP/b+9ImSZux8mAjaWLrZe92nuajxpOHN
rNi6WR4DLMQyb9U+M1ol1cUF/RvWTHFVd+kfmhGk+rFaOrd6i8ggkVrP2isOytM08V5FroTQpBKf
lIAiELGW1o8Ua1YXhlARvwNhNBcp4RJbIyC2VlVMoezlpjCCRUPypU9Fv+wB0jiNRENxmOHivR1e
B2m6skw30TJAZnfmLid5AVVn5uDu3G4AgrFSiOt4Aukw2ymKGJTwiMMUbkp/829jI58NsEFDLYsN
fCI+vaidl25tyJwheku5u5iQWxWLRW2VBqKGnzdJe7fuwLt35uFJUB3eAkVhbIW8lRuB1jXQdQ2Q
JS4suE9i1uopCFiftmWbtcGSmbdFcUe72qIcBfgIaHULk1w09X0nuEAaW9ObcjV+qFOh6NJRiPPr
LNt58ROC9tCpPwCYwo0Go6g4PnJ77UHHpfgnlJPDS8JuRpvsP5yCYbzj851wfDqV4w2FVtF796Yp
CEfoWIqpot3mCCJFe+kYVVtjfO+c4J0Bc9BnMMlwXJQ3ipo9fxhkveka6R+Yv7ur3Bqdlci2FheQ
InRwaP5APMq1UVvU3SqEBwJDQYlEsp5/sM1q6utart3H/8nj81Fq3JVDWmZX8v27g4WWw462efkC
G/LMnIFbnvVcVls9Jkr4r338lFm7THYjFt1Wz32y8Is1v5GhvdPUmoz+EyRXr7R2OEw+9Sb5UYpY
u4duiCIHl7scnIlmuqaOvCpRQDgqggW1NlKIBvqIkHaANTOSsVPpbmKidezLUQa0Hvq5hHw70vIt
Gj5iCYmIZa+1RnyKC6SMdwoatlUz7DTPdk64i6riaNLGmCRjS2HViVFHLMsAcnep1mp8eFJaRnGV
adQCNWc1+RcdF16cA7+w0Ykp3znA67Enkw5mwLzIAEKn4zBsWeRj1IwVEG1f2CapV37DwSvn2M+u
6F6Kh8N68J24xh9Pgi41oYaI2IJBgHRy/Z5WYBhunb3xVucSBt5ezfwrqjhfB8/p6CLKUeKS/ykr
YulKzswNNjqjOT9p4yrmMHaZIGg4jcaYZvv6L7V/GhDfQwC8FXmulOrEqpcWdVY+qu7izdQ9+t2l
PVFFfCuxVsZht/TmIZY7rlERkPu4nOYg+C3VvjHCILPwR/n4VvUcwHKZxo4NaYYwSDnd0ywshCjH
mhEcjeL3zArHr6r0zwIxMrwX5sBnybcOi9cKRsaLaY0BAsCNYhUVYBjf/DrD9bmIXTIy7bGx4yJq
nSVj4C/giRl35ztVMTsdIqZ3WV2fa7ZgEO7cvShiWpE6nvDeFqf7AfhVY8j3RlM5YVFkNy9VHiC/
+2fGW+FzUr3kLD/8xUwZ2YM5BjrbVfrZneKorcCQxUZAapjekvzhBBOseisSMIWY3dJ1bh+SYSGJ
p8EvDETkL4HuMcO6XKUtQ5Ot64QpuKW81IMpB6/xp5+KElKlORpvqo3Ycn7+X1x6idR5ziaIZUf+
n4uLJtGWKRMdeajFJyUwKDfNTedNYUYvk9WJ2V/vPpYcz6cykWc32OSUJxlHkNfto3WbW1xlsRz/
Jh5qjA6TVIPsjTdsLoKU5YKxpU7WuNfpjB7Qd4FC9M/XPK95hqobP0S3xEazGWSKkvi8YvUbYbwU
FWiR0a8MRY4Tja5lO+irZ95GXjXMBclDiVnlul+a9OoMSHvZiGbg+m8DZ5gEjXrMeWU8KM5ZmKru
NJHZsWpE6zt6IfjZQZElo9GDXrKt5+gcVGy6PZiFUwC/LZtYOHxIsGDuSxaLetaVRIp9JynaTV5m
xnXoMgUSDv08isX66fwEAzqgTI+eIzE+yBDrr5hlaFUXfX6yW837cGi7SSYNRRlv809dq2Y4It1X
g9qoxE/8K9h4TSyCxdnb0NurHd7F1BK9A+xEBm+tsXDvyqB3sTiZ2ZsCcS+umDaIaicubET8PiuT
JxaPPdgb3TQrQtIboe+wvDglP8yG8NfbuLzQKquRADKAZkT20RAiU8fVmSPjWaQwBeyImI+SGREY
yfPBYBNuKHj/FcTYtTdUz+qHc6aIEHw9GjQ9VwMLm3Xg3k8gFT4uqbljhcKAlEAvnjkuqA79y+5F
bAcN9fcgGuD7cHrKQnYeeS+HgQ76xi1YF7PXJflT41rZSoITQ7w3RgB6r6+zDkdMFQMhciub1o0H
plzmwyII+OlVkmICNGXgJF7x3DG5jAS+PF/H1pyI5VLUiqK197Jn9ESwJofYEZ1xsXFSwj7WFto9
ZZVY+nCkTYhBkfa2rX1u1nSeblzyXKLJvRIYVS+t8OEjXZmbX8gvfbu4lyzGyog1k4qPmJXK4u7l
FBR/Oueazik3gTm0X0HwHxWDeRILYCnmz45JdH43MG6N5R9BNolcCrLJRkEn4E72N8JBTUtOUlqd
kVSmnP3SoIPpAXBMLfOlALZUEX0SfKL+G4e/h1DK9+DmeNtmxc48C8l2t7NK7Cv5COdyyE8ernav
EXk9h/nawf0k753hZqB+HzCtuPwuT7dRnapDyqfo9ejBj4H0HAAUFAvzjsyej2P9nzn/eiafsf+G
6pMtm3lTX518syzKAwKufINxX+r7YGDPndXDUTYm2qlDdd6X/HGICjMB3ngIu8h605EPua4RWMX/
GP93P8i/SigG5kkaP6ZjfzqHdkzpj+8Yu/ROe9XqvGsHQuGSgMpK2HNoDo7gVV5xbqXdy3HuHd4X
/F81bFxoHb8UpNwFy52i0A5a7Dq2aoTr5vCv3DrZ6H4LR1UKpL8cxOIt3hjNSQQ6WcBLjCmyC3hc
xwiFm1eGB2vMnStQjpmaBER/gxV32vF/j+eYXQbuX/Dk7eph9VFWitFOGbxlHHOdospXRe3e7Roq
mogpUyFKQsN2FqTTtNa2bct+UaAkV0XOSpA8+h6DCavg4sMV9uv/axvdxkXcwS6gDFp6+xYmKSaR
5MnBL548EpYPJY19HD0rlbHsLMYtEqoR9Q18uXL4Idraj9jswWaS+bjnfakx3FfaaUXdYrNV0QDX
DV5OJ+LOBtv9Ry7GahRVdUBt3NsyXD+cjOKKMXnjIzPJwI8ZhUd5ExpfE2kVSMbhJdyStfMAXALf
YQnD4xY68uX0IXqfVmyW+FlgBrerodtnmu7/VzN+2gSIb8YVz7Jl6ahY50tdF0hMF5IdhVvNSQ7X
U+haT1xtj5bvJu7RdjjqXXbinJ3RiKifEy6QZb5kAKYEfe5jZFGBjgj0YZNOMvQ6kwWn4uevxM4r
okZexhqLrp0hEjUgrI38LPrQQk64io9UswQF57/VWPs0ohIGTRVot0SsSn6iFuya+ppWLSQrki2p
jK9qD3Rxi1cZGcjdUSMl0OBu2b6ht/WLEjcLgCxZ8HZCB27FK6ZF52wFU+NJmY/5IND3uYW60kYt
cPLzrzgp8myaENwXS1uZd1p8ukUGL+pEeBxVS2TWD9b5IubuKAAjr2BRO2X9wvfEpIAspekoljDn
onfElzsO2u9uF7eKuleIj4LY85YYoVcJfE3T+wzYDCc1I4aJ2GKFE3fNjwvBx2sUw4QyMFoErCek
fEuzAQq0zHCaZDe5tMDdr2wfF2nv8qvxE2BWhNhrem15UpZZjAE2WPQ/3LN9Sa4eMYsqbBmA5nNQ
5nRy7f6OmOOw47i1XzmaXhG3tbt11YXruz9+69eB3T82Oh9Vxa7C6iRp/pefqYQR37bS3bw3Ui7P
JqG5ENALEjDZloe7Rwihc3Nq4jcJ8Td15dZcx8ZGLUeyHIfda1PEo3BrBwLHurNYIc1uQyEUwISQ
/Fo010prY0x6FHNA7ApnL3DTqMKzw1wgouLS1ohpOWErvzmR/siaEzK7c0w765ec6hwhZc74HfHQ
sDbtjN8KpNN9RpH59nJb3ouunXXbR4nxIDrVYIp2CiFM2/7F0XMfQGe1bzmrA8ay2lwL/uKyeccA
sI2q1DMyDXtk0zskwVpBL2GOhMi8dLFsei+3smIetIDaohDkazdouJOf7CKbpTTpNdEsE7WS1Q++
glClCmjY86aDHCnjDNJYItPfiSQjiJpQ6B1yTdlEzIwMLZTXexwMcJTUEMs2Q4gZ1dokstPvwoe9
U4+WfRNCCjBJpbxjPlmqURQyghZo1HepIh5AZWjq/aSaPyyaoYy+yhhJ0yhCKZ8vUdkzE7k5DcFa
OVWLrwieT0EFn18CJl+9v3zEH7d5NwOAjyJiGK+DeEWkQRbmGjA/anP99zdLLTXL+tlPAIvKsj3r
eMwLc29LmITRri/RvzPVjKNLvIzfZYgkESoxPIy48aFkD/JbwmaQUC8MKeEoPfM9oTAc1zfuUgXt
L+M3Cs+omexIYu4DnT8Miytq4x7Q0SdIwuqtNabyXcY3BnTtYGfvAaDaG2TXr1kCRO2mS3Y3Mrgp
yTQWJcjB8v+hxrbrkFrLDwxA5if9x2QNRAkj0kv9wHKJ7CEJQDS+oB7WGaWI7JXWRo1brtMqAMNW
nhLLjAAVX87YTs7Qzu2kEr19AMd53Je2o9+hSaNeOWhTPhbeduF85q1vQB+bKcRJtT8famVcJqU2
5hL3pqLwUyrHtzLJPSe0xY9XUAsNa3xqNrmAuQrYw15pgJ+UHJHYnq+YOI5wewAYqkUUS+Snu8pn
VdHCG+3TMysOQkjt1iq6VSpEd+vVIgh/T2kXmR5CSZYjhviCIpupFQoYh6m2y310a7j8ApTrtFvP
C0qhXravWDXUYQMSFwPAaRK/qoU4WtGEDHsQPnRY/0zqwPeQJN0OQypgJkVtXftcXbiIcLXoAAkR
u63cEtItBaPSI9gpP4qvqT2A4bTZEpL9EKGO0H+pWeDpPo3tvOySld2cOgvWLSFdIf5a5f942pm0
4h6zmTnJps4+kf6mhtyDHkMUrW29WGUVIxHleaeKYP5iRCjqCt6l1ETpOaP45eCpzmKVETLC9Q+Y
kVOFVaLjntDJ19cH7wLmCzw2ZbficEvjLGaDlN/X5tI+iFsooo8u2q6QbGsKMVuvVgOfgj/8SXQ0
QLoWAufJC1/mzIDM6DQVKH4RYoK7hgjFYeGzglefhzMdNoOqsymW/TU78wH4hpybbGuVjdg5i2HK
+KGIWBgH96sQipUwVL7edFs2nX6hcTtVavaXtgz5yOsLxNo4WyzMsGG34g1TJjcSYre1DrqrG9ez
Sh58JP6KXVEsOb+ZOlBaQF/yyqGKlc3XGGuaca451gcfF2C5rYX/Y2T4F5FxqXGlc1cYYBDOFMhd
4sc5nSkFLawbIIYdM8sCQ9Ov+ZHAwAq3aYwBCz+CbPCJrUsaHsjN0Em+T8GPvSGHQYLeTpWhWWp4
nE7f5y/z6ipq1YHM/RW5ElRx0VuxrRKQerLKLew1m/PWkW3aNA3CF8ddWDI5q7F6w3Yl27DciW44
3oQnlxOo03fP+U1T7cnEBp9DdgzVdvYmIphGxXvr2L0QZBjiAN0l+Ld7lW9QjSmjyjAZkoj3sIq0
6fm+w9hM+EwDK29fbxNSO7L/1HZNBoFUUS5LZyfkwEQXOCJ3+zn0cqdimlRFYvC0yZvPhkNq0pdF
unojQbolK0XE48/kVIk9fJFIzN7/LCEOre/hQMAdMiDorcQCM6+8rqN39rGUzy14BBBJ+pieM6NK
LAkXDzruqzd782RTK9pFcnrFxE2ay6nZvWNHfWjsMxDUcaU64U1bz5GYjMLMpFSXiL1MzRIVPa8Q
Or4bH1wmaZ72NnfSgWrsKi8nycmcBfu2CHQK5UHxSXlozJIAn19vp2EgX+if7In2+aRINE3s3TbZ
pmzRTqKEFGeBV22Be5CloZOI+pz76W0mtipyiWxWd2Jmv0BO4tAZ5Go3duXYxphPKef+huIFRqxJ
1ZI+x+7RkgIoPF/Dt2dED9AmRDJKt47E6HIxuYIs1pomz1llLVERXz1kkv2bbbIZtHqrPZhr1qD2
mk9mcd/o3l9sLsF2lDrXYxI20tcyHTzVDeyM68AeBHBUzfEZxwpxqeDSDDWNqf77xJobm1zCGvzq
hC5guE/USqBGueWPH6c4+lAEOXLyCVoihCAs4QdIAGv0uasF8qTtsg+fOvulk0GqPgLJmLUc6OYM
Sb4kivExhuYIljSwvIs5lC0G5iO9wB2ePJSKhmAeiaSlFGzSS1igZMt0YPbmo2eXi30kWh1KM/Vm
78r5imsoHUM5X11rWj6jy/lzDvx7+8x4VZJeLxPA+sNfmgbsXPl1oAv2N5Mq6y0XZ3lzcPFQWSyV
/3uFSsTgTaCPLlspuArPs4CPvnLzx7lVbz14i+NAz9PHIJ28B3XOlu7pkMivzYVTXsWOEODYJ49x
VU/uSA1tUWHBIPaAIhGjHkrH0woK0EtZkdbzJTl1tSxhQUQzs5hzCYy/Mt2gmUf2svKtxPpc/cO9
R9lyXVCIMe4gfOHn8S+lQQKmmFqoYlNVfdsXgAYE7AeB8PDp/U3ryXK3P1M6sSr92t1Gbjcyw5OY
vJTw5f1XUv1kiEU9STZfdSDz4BWxMig6jx4ws2ihweTEMWCfLFUJ8sEVEC6mG+j0aolNE1U5lIAr
qIbeyOzTwk7NAwSDfo36O3WJ2GRrh9LgM00aoCRpSus8cjWNu+YexU2AgYgNis8EApwfpDKrw7Yn
j0EkjegFRCMsxZjYFPH6lcPrbTJUzT9s6ZrA2bSTm/LDiFrsyGFqKyg1G7e1a6EEd5+mPxfcITYc
tpn0MDy2dDoPvSNplptO67LAp4r9fUm/0kbQg3I+KyCQsLG2LIvDm9OS+4hBpb/HQoJIQr5Cg2hY
paV6fTypkYH264ToZIq8H8NoXwkZxcijkaCcFZ1N+6h3FYsPTmCOZ+m37x6PJipCwunjLIoZmkzf
7NrRKNCNZj3VJOBkPKWb9EfPomZA0erWdDH2YpnMiRWH0Fq/sXxXITBM2F3dRf+GFbfqe6NaSJhE
tNqf7cIb3b/3WjPpNldwOlr7l0CjSZui3y1onB7/Me350j6oXKCCJFgTeU6vOlXifh12J81Ctxko
q1fKcw7ZbNzoqLzF7w43ZCcZlDrPgeVHAMFGtoNPy7GTfR3NnLqMF44vg5RVuxwlYc45m5fiRifz
Vqo+r73KrRiCzvs3qKv1qSe738NDOrKhsp/RTr82aNNAAqV5KFR6dZvGOtQkjl87UgiMkLQzPute
Ptm9JMJVL3Atu4NndTzfHhlobPBJfwwIqxAu/HgOH82cn3tN+bEjx0M1hUVUzy89lgAW7fPqAi1q
5GBViNkYRYUn9XHEImewXpD7aoILXvlLN9yVk6mlpXRj5rAIZzfHpLN0MF0X44v0DwiFMWpCHYtY
2RFIR0PtLAXBQKHr61JcJHK2hdvTRzxc4+2HHYgKG7KC8d6/ArMDMnNVS2WBL0Dv8gSz7ZwGgE95
Qmk8XY/OZ+RM0ikMK4Ok9uzHCeba96BaJMXqXJ7s6m2tnu+JzUkS0VppU1+0M4wbF17zRK0yzr0A
0rOkHkiRqOXHBOFpc4qMmjHC9wJyRFKiR4BRElyrdDev2pacsjnA0P08lyY+8piNKGv/LEebbRYi
j640R/Q0Z65SKXCdCo1Ev47qyftiynQy/M52CpJ//EqC7YiBzQMJ8UdfCZboYFtiJqSBp7ODUoyi
ezuqk8lfZz0bEOGbF5O9zchNet2GoRIzoKyBarFREMSYNa+SKK/gRvb7yWl/vEEmd7VYIg9i7aWt
i/ZjRGp5W6KIPM0QPRirm4A92P14yKIZPFccJ63kzX9MbtaO7RS/Zi3Yz62Xy6K2aNhdFHZMkkSM
YDVOhDMVGQeT50PcuGhqGI5ZvALDpROf37p9ZWVANgT9cY/Hsh0ezCkfsfKeLVgQ4HysZXda1mSe
TDQO3o2zgLucZa09+gjGc5iGJD321I7W9JKiNmSNIdmGuVfvq1JR3qmuMPp+AkcUQ3QieDeZ9XWq
5YGAEf1El67VQr0YHkS6ILmIDQolH0utArr+Y9MNxG7Zyj8Yhd0v5zBg3w79b87Shwc1kHL5XoQo
a54+qrignAv886OjvywvPYMPmNWBgyX1O26yQaChJPG5bF+sTBrwE14GDbsj694fSFqcq4KR3Jwh
6obhmA+WBdGuMmTAi6Fp4iDMs5QHyd1WDXvygo8G/WveutZ6xc+xcfzfbxSQgainfceSrJ71ZSA+
+c3r3yO/CoBpQ4zvsZ11jx2OKd+Xm7OE9FdiIeZJx0gs5bNx3HvvDn2fXD68ZLPwrpt/TUoxx7v/
U9esJDoBZ5scOywIoagAUlSjzAgzUq6QEt5RzEVeDP++ZQRsMscyLI53KWLPIo+71ahTLx3hu5no
LJsh6+mD6Ug3KDxTO+11yddCqTlo82L0Z0N+yb8cfs9f+tTGejqe0XmqZpnrTzNzSuHJ19Ba/o9L
kh6unUIBu6o0H090Bc5VuOBsHpaiWIBk6eU7VTQliYs6HKTWHWGEKt+fYMPcKA+DTcIDg6efi7Xl
8mTUV+3/NmTXaRIBfLNG14oCWShO3vjIs5xZM1WK+Y9NuHMrZgrwcDncwHC0c2WRjSr6OSQrxeJ/
9LMv9YTIKZvnpoOLaTlSqaA0A97y23T3685wIeMdCjsV2iCe3kOQMgXlFg1mB/HQcWU9pnZ2yGHK
hcatmHOToq06FgYD35gURKYQ1ifYIemTJkheaYEAyg11RdXJ+EBAMIOz6CGY5WgJaPSI2R21oS4/
wBhs3+i9XGecgGeqlHbn3jQh0Xm4Bkg75/7sKKweluhTkciXtsLHxx0RFHeopcH2ULLh4AiH7Qn0
HMGz9q+O2mMdwoDc3Oh20rk6I8GWprC/OjL8qLQgmkf8m7mG0RciBa+aCbRAt15rw2wioj4KR9eQ
h1ZskoP7a8r5csyM2KKTkOlMKNOQoqf+0yv3KhHnUi57qOTGzQwzpuQssGoAjxNi1omf8/fdKlsj
7DOnnDv7dUlBnlFqTDXO2qtUqVN6dL1juJ8BT+oVdlUq7y1ks7lnP+ML1d+F8Uxolryd+eHzONNX
bAYG15w94Psy/Y/O6p6LPNoxD2emTCvP+4AIuq1aFkGrYMnX4MvIiiF2pwD6MLVhXYW8/1YwFvAO
guqJ1qg+Zr+NzzpIM8sEf4yWBNNeog9s9vDzVq8Qf3OX4WFtLvqjU11z7nXmtVMdTQXYVEvztXNy
ZhcISDsMb3KN8X1+02e/puafUCSL4zs+oM0MxPM1DNLFcHActsOZ2t9qJZvbtiCCVkGZH8g9Xl5b
qvJki/3tM09VNt/r/N6qhG0UN0VdSvQdwjrWMm24OH4hvUvCYBRTtkaWrYpwiJhhtEDkIZCb73Sn
BEEp60PfXVmHEW4Wd5VisUZAgZX6di1HO8m3LJmFGUKQ46SrBVy+ok4XyG+KFsxh9HgxtRpLQzR9
8Adi57ZJZW8hXXE6QLhIflxHhmFRXZrMj+wDDVVxG/shEKJYSPVD7sZp97XDLRqjF3KEiIxNVqjy
OvzJjB4bjtQ5RSt/B+czDFY4vAjtZP2qMJ0zCfy47GSHs80vODZ1+ooWNu3KBawS7sAf6uy2Z7P7
v0B13sTw1aLUyYZZgxuyTvBroisFs5nQYl/I/Ypj3G7PPesqiNifolYOvt2V8l0oTBzG5rQk+49y
K3uCsrUGKv/gXFYmXoUDmQE2aKdFsiu2Tyt501xJccrVJWkP8CNabvtALn2+Oz0lHhd5VLV8CEAu
vJ1nu7MZdYJvA7X43g15xXFQToEB7E4VizU7ETZEMN/oDpueEWQC+J7x5eocON5DZhJ+yeNlAjje
FofSGsgZy5VW6yuzwRqw3QnV2AEL81zWLdGT1Di/gEDcQNpNj+B7cgBcMaMfpzGTpWbeTyki7JJ9
gvbjPIgv+pQoWWuHMJgvlaUOAKA5srwaLPs59XLtzOoI7uTJkBxg4DQj2dPpA4GkEV9LVu+NG9Vd
z50TRDOwYi7XqZATA7oTFCX52PDqRWI1SJBKhfLe7Rvzp6hmT8uQje3WoLI4vpl75JPSvE73j3dK
MXU5a0I8Y+KEG5q7aSL7wca+OKHTfjwdnEfe6jYbBUFt/J3kOsYcKrhliMQUNmTk2cpSBwAtxIXh
+SrrHUxl7XOJMq7BXPuNXEW5OAthC6HrHip+HnVbnkJM/EYwxHjx5rhc8sWJ9u6Ffn5Bhm35YQGd
MJGkFdiebZzTVun3EdgXfa1FRPhjKYCyovAn4dJAwXfL0KbWQXPlhl54Ek8mgfkFLFI1vEhOqeJk
zoNCI22SPqp8gKc9CVPsSQ9e0aE5d/eTVWBci/VXhCq+tNAVVQWm9VsK3BU4UONT5hfVm8ZhRqQM
QCU1r5zG7c2e2nklM0SXWkhr2nk18yKTaSWbjrcScQSqPRq0K7pJ8oz4WF9WIFyj/qjdaBM3Uw80
iPc0s68c8Tuy7jj60yWCvR33Ux+MWtrrZWAXI6KxpMtEJW4Kpm6NbhPOns2MOW0PuVe/RSzI3HxH
u7nqVd6uqwE4MJWPyt6t6+Dgwh+vy0GXk/V5DR8+wN2QqdWE+Ww05Ycr63P4TsVKFMUtbJPdd3qT
0cpjSDogE1Z1JUk1IEBANfYQi9A4TxRNEMKG0OM00Rpnz0int31+FTsk3AS1Sxq4Q1F5If3aQSvf
iZHtu47yIkp5D4A+NJXuTppsSi67xmJvsf5kzQe/Shu9TeYb7X5BosdmvJKdO2zSgwr2Jg8vjgAf
2bFyVM4/yonb6aKZWRwoIlKzUopdiiNhAGZ0r9LgOn63qr7TeqIl9e1T+ZPk5kA8nFX3Qx8GX4tU
SIVOBSd42I1XeSR60zr33JSeLCChMVHFQ8SGnLaOHosHbPx42FB7jJJoxRo1b3KPkXKCygH3L1nJ
o9cJZMHuBEECnAUD2wAf32EDIALm5L2is6y7e2BDV4lXPOcOrBVPm7NeeGizjXeY+WbFhurbxSdK
ffAq1QnGnecgvtpCgEuTkVg+qB02ohj5Quzylkvsr60ibsMxmmzOVEF9mqwy64Or1121fXwCcagn
ZCWRia/qHToibpFsrc4HyCiGV0I8rbA5EjiNSTMWO0NqL5F8YZpeNjcc8cKHkuwsGDkXv3bpieSO
km21DMG2MXYEJj7paQP4md6DVh4gOKb5F0hdUyUYJ9vCT9DJ3A3bO53wl+yeFi0OWaRJea8gKhGg
dyRqjgFmRbe9S+koTajd2sggDeCG7u6brE+uA7tDShgrL5vSY9lLTz1Uo3fgY5WamoqfiST9gbeg
42Jx4j9HyHPNKQizbsspbvs2NTGQZtvVRD6BB9RCZTwd9r55uGzev4L/8Jq0Kwwl44mUT8ul654g
3LbcrfEjlM9vbn5jwiW9FgKBguM3+ansmngrYuoAQIFWK8RoptNkqQRCVwqXVM0tLc5H+TXAcLpq
EO6UXKEJZLiL8sTVbgDzOAnOfnIZQcEGTspV5B/ygc4Ki7sjVTIP+mdZivtKszfuNOIttsi1zUzp
M4uA+1IczpIo03rUgQGIB+LZJpBq00SAy4rbWLs5qv5LZnGvWHKfd7FS0OrGHm5QMktIBfm6KvX3
tkddECMPUFdSx5kbqvFch1i5IaeOgpuUzB8qutGuL1N4ZvDmuEdy3+X6StqumznbGVmTY2/6CkI8
qjOubEzOD4c09OI43WBmL6ROJsEhIdySS9KRk/eencMVhdNTk9ZDwGLYu6tqjOo5WTioOm0Q1RbR
hlZSHam7xVt+ACWelZ/rB59FPzB3Y9IAzSw3MFw70QbtdcHPhdbeelOb2GzYYTEb8o+YAqelP5Lx
UA+lAeLq7j7+e7Kia7eQoDATI/Wgb7kWUp8u/v/YTOCuFvdBvEBw3Ouq6XK10BUJLJihWhox9KCb
H9859JfbHZgzio3kCYpELG9XGoHbqY69ychqj48ddEenWC++AhC/msKPl1k7fJK2o0lJ/s4DZV5y
eHGCf+mPnHc8weP+R1UmWyvdkIeiiYVTK/rbu8cod1SVvrFwIKsV3+DIcI5Wa8s0Xe0i90SorXKv
AhPY2yttkVoBgRWo+oQGAWXA8xiDkAbbs7FZ2UettupXkOud3v4RNeMbyvYZHUTiPtF4tanyw+Rf
37QDQj9qf1zsZUpIprW0LoZ7K0bfJuvESPBallcaFxam0vMXVftA4rpaAf5OwePpAz0bcDVS4paK
hBdzWpFWpCBbnH4UKVxSM//MWVcgTy8o90GFcpaOi/9zszrVI5NSRp3cVUlVKe/AwsOPuc8L9xvD
VCc7TIcMKJeHJTR34G7dOXRU1JP3h5fjqJlp99p2hD9eIj6NE2I6wn/25aRLF9V1DxCersnvNZyy
LY3HERUHUq+9OJSnbxYJkfVuRC7JafFl4buNyJAlVh/9f9sqT95aZhmmlVERZW1H1+A4HAujnKgM
vTXWmFiLUUALKgUrf5RgeT+gIVWEOcm6RUgNuiJ/TsVxtBH9rf5mGAbhRbsXSl9YXvHaj+AHSSx6
ELOLTzg3fGTSXZuPHZs93Ta1SVsBpd0vwhXTsGipDE/i4WauoxQlF0eTTWGs26+nJEhgCq00H7X9
u/0EFe++QEWhETGCkKXVe2lvXf4gaQX/5UDf8WhaeZMHQatokkKC4anOVh3Plm4jFPanSk8vmlXz
JO3GguJyFs64vZwfPS85ZO1gEIB57TxhhGgT3RUk1AtziaO4iR0vCNguAbYb9HP57LjkqwbnV+/H
QD5bTQfzb1t5zz/YoDnsL+z4quhbFWtycLIoEsJ95MugZuEtHf5tjw+vw6F48R8gtpqVyTZS19G8
ZDPBnDtKzcJIXjlAAlYRbcEJzULH2AaEvdsJOLJLceqpPqXcNgavSXsu/W6Ihc4RTwasCaUwxa4K
e6jORbGiJmtGFGafhQItmnOcLA9c0w/aO+fuf3dYZcXLLy7bKGJjDeEq8WFcpxJ4sGzbLl4YeJGr
wzx35YgCfyOQEuFZtdyDB4IKgrH2q+4GesvYy4TXZq9wEIV1y9pmQUHMyl+Yrc6cZwL8M7bV2key
6oaw5BcVxgBmI4pmvutRSmIVmi5ZhmycL8s2/VbzI2Z+S6DBsk04Bs+nUEdfcvICCkrRX2IW/spW
Ar2mqQ7nAE/qceCc8+1B/98USMKpI5sfIIbksX25+z+IWNyK39p7aLRKNT9pKP8to7d0hijjHTjt
iuEizyv1qFjyOcklI1QAhUVCSl2ETF2o7AElXYAS9OwJu9LBTE3N1t8BhA7vAiqioz5hR++R+2PT
YGdKco9Of+fue6BMT6f1c4gbGhvK0ACyBeJh1okZXcxiwHbbbcAntuI8m+OAiCxjbtauWyMvpfkX
3UhpFOiFqamagEm4jSH74fuAAJXOmJ14ravKj/ghr07LYItS7oi1ClCfexOCUgoLsxua4qz1rzeV
W5MMZY5nGn4Y/X0XDJVYxtto2FVsqFJaGUdcJag3FgTmp8x5p1Xa843n2QyC1Q3oOENCdjMXGhgd
yZvYE3RSDSaZakQ/B8AeRIZFt9dC1BjOGtdFd+mQf0qbNSH1dztzNvvv529FoJPC5GlXZ0B7ehbp
bonWpwGoPYro8V4cr5XERpYZfhRfJSmZY2vE4kWTGs9dtjBZdAAEGXBQ2yRPgyu84qfL8+myD2Zp
AuAJCDAzY/5YTDoO3dtahABGSHJ4px54WQkeF/OZWiJgga0gfDhfpsLAzXwZ6P5+1swm6laWQUQI
0VJ01puc6FE2w6ADBH5+ZewgC88phK1UfaVyvpPchEI6pwhxXOVTGauGD9OZmTsNxzTzwaEzLRT+
M4x4xoQEekvfj7DVYoBwwZOyxwYhFCD/s0oLp8gsK6KbhitdYDaIZxaItQue32PuXY6wn4N2Ovli
XqvC8ZWwhDNbZX8P6jjYQfoIOuWeS4X2wPcvzYiDpr9NcwvBISKXsrKPqW0PP6vbCN7rrTaLUP4r
YFmYSvUGRkhGTLIytnDghvtCNR5dFKK+eyRwDS265chAttz5WNndmvo1NWLfnIxiTivSJJwDHNan
S2LaY0/7jcXxycL/lmw18JLgq8JXm9Sicoaj1qSuRGGxl4dPsY1GdjJaQWioeG86BemwGA4nSQLo
3tRaolYc/OpX8f2qAldbd/OX4wZGQHNMucErYMKDGdRNDOKraPVb2TWNkzQbVOWb/ssC5mJWNUkQ
6xv9S+RjRWFl1rNxemmbXxN8NE0oybYZxad00FCS1KKp5pEl2KLW0Yx1oTbd8fXwx9lGMSCkS/sY
yp+UcTUy0p/n0u7CcVYbYgXPPdLrKRryEWhJHQdewEoTf/c9rx/93kaF3CvZc9c8KBj6a9bPqTqo
lh3ajHB6En2cLHSRGXhs0St5tdcftQkgN7CJ7w5rbn0BS+alXkYP86i3NR1ZFlKdFwzvf1QTpcXm
HkeAAfF2QVXnhljeZEw45o4crbtI1yYENR9ciZbnR60yoRRieai37VD4rg/ytEcSBT1LNoXAafn0
M10U0jqZWZU1JupAEwiHCgCRhQbsZI0ZTrf1FJPCBtK/MQv9C/bqg0ih4uDBsLhCNF3DJINBTDqs
YoqSvFQ7dZwb7FCRucf6iK/FcPWMI1UxPjc9+syJ0X9OzoSd/mTffNLF+auXw55XQl8afzSeoS/T
NlomCB6YLYkA8A3j0gSN1tItiyu3yVDf/PNR0jS9mGKESnGmIlAVNYvW62s+F1Q5Nnlbo1ZMfFpf
8odb3wykG81Jn39RA2zhvlxVxczcD7wNuWq8yvTLN8nYc4v/VWaPt71K0cfoOplpq9J1Kf0JDuaw
jz0cXq5iCqQxNBb0u8QRzOlFncGVf+OemV35zd8mkW26VCbf8W0uMkKKqDPyPMdo4jv387sCidvt
0SSbm0m2DdSGgM5Rx/kI7pnRqpDRopyIahoVx/NNYMgReVKRaCQXtFo4h7IXZBdumo7ivwR06w/o
8asp5ykhqUu+DWS6zP0oScE9sXOzTCY6j2PxeIrD0AQZYGGD9uW2NBDPgtvcHdtVFS/+IN5Ry9K0
OSDqUb7A9m89l/+liQMCxlMhm9xsN34II9lZFD+TCb3nMtPHXIWOMtGOf7E8D+r78R21J+BdCzpL
WAB6ppZRPuHH2Iuv3gqgA9FNbDNnGY+2Azni8NO0AmDGkmCiEY2GPsDvLa3KMP/trDb4yjQkxAAT
Yv0uF0vE4c4Ur0sGRizea4KIwkhPIYEA01bnOFe2CdgzSRdM17v7KYcVbtNcGTt07NEs9TgneesO
todHMmMp9hlc33S1dXnxcD18OIK0h33k8IX42if5L1UoAQDzWeFgBdAJ+Go6sXjjwwBxrOTeVFxG
D6azFgD/zqG54vtLrMXSLKAwsx1dN6dQVrLymd85Uh8vfFDa1BM5XYMwIMhIDY99iDoSlFSMLsaU
RtdMp7ehIKQdcva0rUsZIhbNALgWJ3aWA1x7h4T7F+tS3J1Kdy0XPIPXxmNOXuo28Pj3dRVgVBcn
7/PoGcad5ApV7hfc8A1drX+jm4kr+5Nx5ZLAAGo2djbnSpqrJNGDvCEZatELpvMA5697Gs3zAP8s
VK7dU2rUhiH5roWnUWSC/uBscCC5TIXCUsSQ/wTbdDJrk7E0hGIxQZZQ54lMqcBDBKGv6mhzX7oG
e8wqY2Jv0qcBY8Fitsq/0H2aSt5G6hPlC42FHzNMjslH2H6jkIRV4P8wZWN+dqS4hrka/oABe8f/
6fFlo7uUd4KYfzkzl6ZBILCKaW4KGLbrKee/HkNj1qMGXUIgzewgcvy4OG8dUq6iuV0LahQ7algI
N3cO6kExHZSCnD4cPXQNTuvvLmCfG2uiPQxq7cKNRGdxvFqEHSOXFw7NbPHyN9G4/K17lxB5vmmc
VHyvmIH1QpuRu9RaK4tndkZVjUlYv6/AOaP142qC/bby6eTo5tXGlTMfLvnCEEsjkA9oK2e9fO9E
MPFYdHwKh0NelsJrKZRFE3NP4Bn6UINRVIw1+pifZ7zyHqUqb5DJstBnj+MNj4N1fbK2okawWvV3
LiInWJezonmDqYFZtqakbIQziiG/Wk8CxkQIaoNqI+CUfBeeAwI222ewoaWxd3elS15ToDw4BBuT
ST+Y59mn/VkEMMh/Gq3b5UzSir7KLkYBTkQRyrbyI9Ib3t7v1eksyeoiCraYgVymYzOnK5TGmsxu
8Gfo062uvbvIFSXnGFQ9zppb8TJSDq8IjzlH2ZLLNaro6VT28mktwhi9Xf42HgGggFOeLqcvWa8E
2Z3qcZHBg8j2cr0S2bsRbKT3aWrBVdh/h3ifq8lS7cv6jJGq8LuWdkTq9YuaZgO+nSzFG5xymQq6
CPgUzkY84IWnOMeHju/9pOdhZ+Kfbwrj1x3wtuESFvuFKAmNyPV3F6v02RSFDsQM1ioHHXokNyEs
WYJK42HWlhllvDee/B3uPPxcw9G1dMaUk4g2wou9BGaF1LZ2bycEPQBR2+vUphH7zO6izHTgy5Y0
vg+P5094rpjsDv+L9j16Nb4VnTIq7BlO4DExpdiY+RKUAz5p0P7wp/RpCiGgdYaU1oXWS/XMjl94
74qkoS+sMmXUrBU4bsDOTmnrlQmLhwAxb6FYXnTSB7m8tc7rnj7ZYUGu0Xdh+DDrHI9CNKbhwIi5
6Adg+q6TXSBOb98mcSz9YZM+nSiaKV2HIs6tnkK1hZ9ANNfb6umnrbpeDx6wLMgt6hTJ+ju5TSna
7m4aYpLf7EAm8ts1Hqv/dY2UH+mlgFW6j/KL2sqZ3SC+4iQ5JmmAM3GM3RuYJ16fN+f0GL+yyGCd
lGfJ97zd11JSpQCvpLgJoRqakcAtQEFUBzniSECLZGn0uSHDMpJuJbckUhX/uGTdv5YGXWfh6Mlb
LmmeL8COHAUXW1k3B/0TRtSvp6J9M47hzeL1iPEe31qZnoRF+BWcOJgxUMWbxu+kav+bE/KkrYja
ge8k8MdJmYuVKYuHSVy85MFgzRTEAJuJKXl/5HCmZSdYZ47VAmdlLKH9A7xwyNMourjzofqw1lCm
oL/6lsL64i6ZPCS5mwwqmwKK0oqavQQD1bY7nRuvhehT/nUR5ZqZG64/sK7oTTxFwz1eYQyA+Lqk
128U4MwV/yCneqIa6DMszAzYGzx+zoHTugSASnj3CHCUM8YiMFbbEPT9XIm0/Xf3g6+wZy1KvY+K
Bjr1KxuNdQCdaNCvrr4p5OYR3S6pimlfUPGr+V8zmyDL9SApsiHZnfUMVvsyzXSbHQj8alwLFKc3
Xerz4t/W2DGuKmfX52W+8AhlDICIeypueU7R16VKKCN/aQmaONO9WzS8/Fsz2xpGP9vSmLo6ucwh
L4Wj/Aa+r2GbVP9xEdVuuMrmsy1dij4wiJ6qm/9S+SSuSZLAn1z6Tm5Y5cT/5HJxmMrYWj2IoOHs
nM9u8uEGSo46X/anSN2tqzmMePHKhsXDsHZfsGoYYBReAvseMNqeg1EwayOKqQyeY/9ZdxYDjG/o
5oPlWur3VkNt7cVPqVF+r50Ngqf/yOlIXDVxN/dQ03on5802PN5RfDbxsH/lWQq2pBa8WuqwWpdS
7LS2cNM303F5O/gu0Uojkcm6ZvU1beH+Ppdy2P2+kHnSzabQAKblIjbbxL4VMj730j8Ov4weuGnr
8Fb65Yd/tyTw0oENBj9cc71yP+G4KK6eGw0GX99en8PaCDz8zYZjshEfMyaCUSRrAEB9DsYihYV3
HIdqPo8TmH/CaYYZSPTpSXY3Rj2h3+ck7LGS3HioHXLjrdjyHPAhO7oGbw4S/tI4eE4mCM3fzCql
rEsKdHHFAPjZCmNBhz+2ZHMPgstkhmNh3IgW0zRbV98Hcy5AOggjbuZPRt02C19BvQb5vAOU8zMi
NJFQJAlKVHnjJwEXbHoIcoJUqBC3ZycYhQxOQxjlzy7VUw9kWnU0MzT8DFOub42oJlh41r/Ax9WX
QWkx/cyZ6Bd3xkKMpQJEczPcM6Is5N1jSFKZI7jXEG92wVHsa8srCcNUaSOv4pc/Ns/SpeYn6ZKP
kJeRubDFe+0dHrUn+IqexhyEls6OPbh1q2b31B156ilzeD2WIiiMOt1AZHu4FvF44AEtC2rEKYlm
8j2xFgiHsGB8wn4lV6ldEmxKWo+l2cOmjisfzERHp+L3/aKFIVPwYsT6KpkNv6TFP5tb1b2xB++Z
HAh3Ji3OxbIOnS4n1kMryiqIE0vhGHqR5ThDpoO4ZjdSxhtLUuMM8Btss/yR3Fqb03SusPNCFYRB
JKG5sMVHgTehif8QX4HpUYo+ohRrq6xZS1n1NCM9EeKJhz5FBv4LOsec7/mczgywFlCeP137AwCU
UfrKAPr565Y1xp3XUgRCMrKe7WV9klfsVLOom3E9IYKrPp88er44YSGCPVXJ5PnXmHKnIb1v4oNw
p+3gWRH4svK3BnNVoLLJnTeRMhEYfEhaYHSS0ynOwasrPVyuxvGPiipl38WvHnz5i7H6/lBWMrjD
sb19dm7TRxluvks9Cg4/MKFpNAXHI55BR2mEBgZ/uK4mENXNlaxHqPPxW8EkUuQmNEVBbZdvoojW
NuQpk5EnyUYjbFZBRVDlRFJ4UHJiui15+Z63I+W87OJmFkb7EC1dPzF8BaxIWRXx/D2lZ1GBS/DG
60HTvkV70APQAmv8/PsnzOjmYDIJlPjw/CbtkNl6hROGThEit1OiQ3Y5B9WEl/X6R3BOdSdUDLtZ
MyBWUFwHT5W18EAGXEq3frsKPn1WVr3lN8N62gfo/5WLeIaKnoWRZdIKL5lthS4utRExA3IXao0/
Y+o0mPRjeVuORY1UG8JU8UIrPMG6CFkgPaQiaskdStYnAEdfQarNfwm3e3bxrRyotASZmGzl9lv5
t0OI8UIUEflc+3bKhYQJU6x5dkr77bcvcwNjMbmvFx2xUJ7nXD5Ok88y1NRI8vu/U46fy9antGdp
0q8iMfVwE5F9JD3Z61YyXrPqMKVPEeC1jbXLHC0yJxZwOqcFgtfu1W6IG1x4WOJjcmTLjm/hMpRT
NGXHtGL0uwbe4K5DKGAmAIkglQalL2lSWfUWF85NAv2oEOgnOD4VE8RVNB7W3n6XKrftubfNSQyF
64BNi2QbthYgzYPZOdzUWWAXX//sJPdSOyQa9LQPRVOFdybreQXI+yCZEaGbk1X6H5EDq6zR0kNZ
2toQR80Wwf+7AKPyBe/8BVgSWECFzb5Mrb+JYj41ER+sb5koqldcoZENzG2eezhqu9t3TE6GrEGb
YYUEDSOURKjiZnBHJxYTMSaJNhgAB8mVGXZqfQI8srqpBWQXnKlYe/w3NAyQrf6zfG/pTWd9RNs3
3F2o7Et0HOpriwHBeAAcOZG5HKULf/CZKLaIBeWHruNuyalrvkd1v3yokYVe89mMoXAlnXzMZa4/
etHdccOvOeFhsJEdrJmuHWZO0JwwfoiLkwTmNzp68JR85mLNSMZ+soq2RDUprvVCGacBrhAWRToH
ktA4c+L/Fz7okjCiFwnKNuhVAys0eqyOsetHY2O+Dm7Ti9KA+9Q7FgjdpJIyKuehIH1QnY/YBYoM
28vFQS6UsOrl44jESnfDdZgeMVzsV2q9XMoLAnudHSV6c+4z/KxZsnFi3H3cGOfsnobTEYpFcMdb
CMPsrHlHeQWixMp6TrwURKyce1AswJcFrmjW3VOJ4/drWhuprZj8K3x+JDK9CvyI5VcswBqM22M5
Ik8x+WKZAYoYLfw0tryhGXDS0PyYRFIJunZAbNvl2/8oFMGtb66OmadmbkUyHBvZ/JqEgZnQU5IQ
33WYsU5dditCcVSqFu0spVAwwcapeOvDmUQWTbW+V/P7yG74EwSPR9Pz/NkmPcE0XdqLuIlSUIKP
eOaZ7FjLHwRGSwRiVkgZlqc94QSkBO8y/WLWgO0qrmMhjokSI4zrrEjaOAzC66X1zAtwszDSJXyg
bQJcgJUCUe3B1X7S+j9LOnxiUTFQdPTk3IuRDUdFHsosjx9ACfODddOeyo1jydl4rCSuHZMiTK8k
UMUInzM1MqP8VfTJLPg1luAfTTv5usPYN5EvFDoI3W2/Iny694ps5oxlC+ndqu/kK9ZGoFgnv02m
c0V3GmnpSYZyduepn4zMZQj7hjVINDJybBEqdLyHOciovEQF14w2VeXYDnZuAWakV8hJoqriOlw4
Dm5Ccz22pIUgAoolPVWwhOzRAoMNa+WX4Uxyr06T9riTz77Co5QuL9bDC6Jl91O+rUtJJUv0JfMd
wzQGuzvJ3oY/W6h9XmBmUJ6Hu/SMoWTXGoB4l+7qnVrR0pOF7ENhWiPYkQu3yexDkvPoRP+Etf1r
eS0KpTy/3DmoHKids3zkQqRr9CuC0BxKxoYMr1JG3b1d9cdkfHJdx2WVS6lPgB+vw0no5LBwGYtF
kuM6OFYzcw0Fko51suw3D0Wz+C0UwZBMhRzw1x6cCxdmudamKwvzYlsUHxGxMMD6ArC+sk6+NE8m
WDVLp11s9U332a3u19Hqx+32FG3UuAgAmU280BZgBJhOo8B+1HE9CmAoDayE1WvHVeLmqA4YtKI8
IYL5QF+kY4j2ri0/hjqjJkTsMUTUQvoVtDjGJW0WowL5G3+RrCSmhYw1MKLm41Gvzlyagwoc0EA8
w3za5QAj6OKB3PNLZx+Tg6Q//TvHdXO5qJBrJFSX8QhWLV6aXdnXgYbhC6AQdGhAAFJ2wRvzNK4t
6hpw8SgzttO+LWLwiHqy68F8gHyaopFAxXNh6JyOKw7yNeBRtH/n8mqr0uAcfZC3HCdZ9sIxbgnR
I0QyENnYy7ukn4nuR5H0ef2fzQkZG7HeZTMic6R4P4BXPL2QszmI4PeK33vZOaiaNT6TCDUHHmYW
hLeoT9vWXaxSKI0GvISu2bDS5ev8px7yS69FakyiUt5SzPpO7S0XRaRd8uAKaI1ZG/rRqaxMhRgR
Dbj5P4proM8QUTl8ZdX9dNGXw62AJ+I9byzVaKMzpmirjmfi7YTcW8AV5C358mt8TUFvXn98UDPa
79cYzYduGXPSrZrWfeIVhuBNQUyWhbpqcDD+rKiJonE2/CR3KLJdKO3BrjdBBzfgydJTO4OrfGeT
aiQ+TH2pmZWbZOoObTW2q2niowvW8+VLUODMAZuXdmTe8O3kRN6wH+yEdE5019rmCWPStESlPgEH
bF7WLQ3KEqBcE3WbWQfcpOAqGNS2dTc8rYnx23fxFZK7L2gVehn6Dn6AzKTvelYLYYYv467xuyAr
YykiiXtltwsAWsMpQ9r/s2iOJslPG0zSgS1iu3rHwXnPyS3nz4KT/YlHWRPraR+JVkLIZQbXC6B8
bulonPYJVF7W7WwYHbKmgrORW3qgj9vwt6o9EQAWe7FVF5dx/0ifhc5tWDNhP0nBv0L0QbH5z2h/
aCIfiXtXvJK+QF/vFlxnvvIFiCREtdO7gIyEVtgQtBFQ7x7ezrJO7aQzkeKP3KM4H8H9rj7sXi+/
UrNCRC1PYfS84+PsruSEWbYaXsiPmMOJQyib52o3dj86YhDwQ7xRo4Z8B2g1oCsCJLZ3SegB6ZBO
L8Jy8KKiWDUMD5vUXJ8lU3zftDHreLV6TseviLfxyBvEBQ1J0ZtQR470StGsMYl9Tokq13NaR8bQ
G3Rwh1cXpH/7erKsyVJSU+bFjS2biHx65va3Nwceq5wS+PuV41mIuWnho8mPbz5ZB6FtqpTPhlXV
QnShTasNzsVOEVwY7x/xEiwn7hrHHRn8VUzUXBOjzH9396QpTDsxk3KaNXT4PD0g80USbBxWnQs5
CKhOxU0x12KI6+GDoB3ywBqWqkCV6cBp27bAUfgVvAZP/uxwUiP5+oxdt6VL3xSAz45mN0dtGBSg
myWzVK5cZYZ3VvOT2aUgjr2ow2mHsjVbVS4oyb1m/zxVIfhAIY1McKARQHRxbu4Za3kjgTWxMJBf
cf+iOgouG+VW81K6j0fVuZa70/SMM0H8VgI3XpxDDpxI7LJn8MCZ0qa8cxEPjZA6KsynrNdnrhHx
PyiMeufmpUb+QXWtL74zAWS9ZSi559easOi/B3Xy+XpaYlvp7Co8K/elwEC8ED86R+EHYZqR2gaT
emPUAF6tWMDG5fcyZxV8g2lEYQpdulm59QCIj3vpYi0Wf3XXSEI//p/u++OJmagJOR2EcTULb1zQ
LeDI742I2vUgv7R1exbh/2QcAXDLqQFqsqwoKjDE5lfdeeY3020cmy5GKwRCM3TPwVjhpCrx4DMX
+nqnnovDxtC4SiJ6MOkJEA9gJ3nGE84/ubuVDaCBsAVH0srjzcCDjHLEkDpkqYCuMOyC9s+QixPh
u2HnaFozj+uMD4ER4oltWFnhNuvKte3qKfU32dVM9paMoAMaDr+7Tasf0QMMCfWtMDfQEPKeFJFW
sxeiiwnk4WnAzh1I0sDd///jy3tHS9S2S12wuEt9TYJIzqCPAU3KtTVVZei3zw456TfFJtkSK8ob
JlRrtQutTlw7Qd4ToPZCSgekuiY6gAuAvbfC0LrnrO51CYY8rC9PO4HqQczsN0yaSTTzUimQSlMi
I/20RRi8fpiIZ03XBq7iVC46jLQ5ryNBGX+F7PHjdZOfNXJVcc+1M5yuntryEyprrHPdSFrlfBQg
ldIDxRqIK87kW8CONvm2CUMiffeZMSUeLYLbIOiYe77s6PHZhPxPVu3Z4MkRkbAKYlAag3Ru1Cnz
9tQ/TsNvRodFmVegqlbIjMZGl7GrY1i5pxcP178qzDQsXBWz3iUXWV1jff9lfSonmoTH8TNwxv3E
6EKl/7HIEDURsLluwvdvut06obAg3fU53EggCwTZR5mjKzgvNub/okRUCJRwPlKmluT+vwhjvsQO
/rpivyK2VnPjDityyur41I9s2MAIjf/575EnA9jEJ3BDeeejP/tfFMdwzxlBFuAp2fGOIYfK26o7
Ko3HySeGS85cyD263DNeJnZMr+OU5V1teO4aCLRwGDC+LWRhS+pCElQbe/xa9zTku3Rs7EpAtOs1
RbD41KZoS6VYoHIGyWzAmWuCWomNcOTeCGiuSrFavTxeGWE2J01X2+/isDbnb2NOzMsAf/ixI/2Q
Ys0EHqf9kgg8Au79vQitPoniVPjbabDkFUL5SWOMZNQ36GD/nEQGV4OuCN51F/0yF2sSLEq9G0AB
69xEdYlt2BTm+xqTDBN8X3+i0JwntVtLLPaH/N+B4BkooCR9eiQTqPkFdUoP/s5py32XM7js58JC
D3QwjyoMciT9zVj+aTRv0R94sSNYo1ZG44/qMGP9p7G7VSdqwHtWIKMxyEd/sq6XazEb5c2IFs2X
jzpBrIhLjz2rhuNcQ1NFDQK13RxAF8ItYfqT97Iw6Z4vT+modfJD0FhbyNan7c3w3oFvJjkt6dh8
OVQQHsW76H0pBEotO5s8jYEem5DkA7fuvpxmiXZm7TVN8yKO4BY5WXTErLNJuPo9MTwEOTN8l/6z
W028IigdqgW0my6+KEm/RAN9+CLGXtVh3OhRhC177oZoFeABunLWYHixnTbLYij/Pk5Sv/MUniHD
+8GlYzAn0MNOgBpFY1cfsMrY0th8NC+gQYpthWyB9D9gUb2XaoV5B1FP7Z1EncTkwNUPAwmS3gyq
YMWumm1SbMTd6ogyKCoNjRLgYwUio6oIClELZkXBjoCnzRKCN0nDJPykN3dD+wu0xXc0sc8PdRkE
P5hdDGiep3I5FR5q+6sfnluj46NYltWPr7Vw64/F5bUnSYbNFybSA+YrVY7gnm+FmsDpj8A0fqwC
tJgO6v3AQEdGBufcpKKg4Waxf1yRRvOz4qc1kPjmRkd3sXhkZN0BYwSwEjvwEsOejCjQahYaG1gb
kIk7oOyXF+Krk2b3gRdkyn5/14GaiFgkRYBiKs08enKXOjoto7kKDIxl02ur1y/ebonGk/Bu9J/T
y//Yp/6fzCzH01LKDF2LUt3IpnIb3aHYZBkco2NDplvTFSnSp4YJPCKGHjJPp7Oc+VMszgUk7peW
tXpA47XLZRgVzXpSrXbByXNDhPFnOryaPwFLXkL6qMzIgpbbH2PXLXXu/DUK6N+wmkqT830iCzDT
vof7e0EoNX0IoEarxIdU/el8i8n6bFdUXyN+lCn2cbdxXJsUe/jSCbCw00Gi4ppgw38aqBouor1/
y206jYr+8kwWl7un4Zfal51eEqRcYWrv465dsi66/fcGdFSHrfNdowiD5K278Heks3hollec0PSy
o4Rx8ywNz/v5oYWLOEfrU7LkmL2zL/3jeqr5FCUGU/iLXTBI1M0RimYToHxrllNAw611WJ8n0zff
lL5UiYM3EX0kVmUeSQ8tQWEqsPSDG4nrhI5kQvZCesCz1am82PXNQ63YUT3HLAALpXHiaPp2gq8I
TrthywYZprekPtqT+vsvHOOwlU0YVxS+FGAN7wTHRUMtCCbnnEQHtvmaQmNA7qWTiBDqunXmpa6v
zcGX8WUXRjkSDvC00xLF1XV3/uNPaBXvV3M8OviuGBheBGe3RVBILOeP2wPVr3NzqvdhPFZNmHTZ
U35tx3ezZ/Oj55Qurrx4bg3bjhdukUH4ChxjbwI5GzOIcLlYXZYHW/lzgvNehYClZRbw/b9yc4GY
yBN7v3QO4prnzH9RilHHI7UtrUPO/V1uAqZPtcg9mFbw62NRi9wDDMtxco9mt6ZUtjGvggziHvxf
3SjtaRu4Dd1cMakvNZ+44Eyr5Lu/yzgJGkHo7EzbFTF0g5LUjauDpneEof6tXZps6VKU7PPcz8KP
ZCY3no8UOLbHzNDTPeeIObC65UObd6edDo6tqYKZMZBRiHeMMG8EmLe4hdnA75VaIdkcfWbeXcJr
btfGptqcwHeNPtytO48bno5lVlaJSdS/3x6PHjLy6I5D5JBfT83JldrOK2HQ7YxtOlTWDWAmFt5t
CKdIFaeBPNYcWSsDdfvfIyxKsPTMvent4BqC2/gIRBkexZ8EMmPIGEjhMMledKSfFmTgaWG9K98B
Rydfc61PRM4mNt9JrrpUJlPguEZtkC7H7ybuBjjC+JLxdnWxqOBps0fu7EAtSU4LVAXgFh5WBr6G
XSSDc/MPiqC+s8ZWm+GzujRkABeKh2LOxGFx2c5DPa8yjtAzLE5jP/qzlETkzylnh21bilw/7bUy
WTqWdfDm2BtYq/SdeIwifEf5/0sAqrbYa1FhYCgSQS43/6dCGSh26K2wsuWcpr5Q3wfYHlWcKKhH
p7FwI/89SFtLJftgg/G2mAUKuUQNyqTay6MFUlTXb8RhMWTzf4OwgXeDVuLv0sKMbhw7fejvGY31
yeQXWeNuKcTijY25yVIrcQGXgH23sTf7JBPGaJnr68cRd7hNZDgFbqIHvAEtqRLdnwz0JT8HHLp7
9aO8Xb1J3Be4cjf/Xs0py+k/ENf4HG0bdd4904rPQsVWupEHJfBBCX/Qr43v6eS2symIczdGlfNa
1ubIbja+Ilpk1LjFJNo7GLlc1NPSa+SqfO+mPq3OuCFeODzyJYJMNQAjPtGNAJr76z1t4J362nW6
AM9L4dh9214BX/Iab2ixtwvx+UoMfQkjOGBepOdQeco43NJK4+yAhqk3uq+MIxeUpHeWJ2tQ82SF
59gsiKBhnTfrsx0Om2dViDlBWdXg8JM5YksNeLhHGU48BR+OxQ3xz32vBGv8gV5xViMLqW6yHdAf
mFtusljcLJl9OpGQvsxBgpBxVrd4N8mwmwYmfV8dUCs62p5q7NagtMyhv0LWy8f8q2g2lODC2aVf
j+c8apAHGcshUs792EHt0JXU61mhNL5AJUjJqtaMRDeYJVj/OSDlMYyjHISBdveStPk4R9dmt7xj
uxJwif0j1YEXW+rwYm21jqvfxuDTUZYgwvJmS12zb5LhBCNkf7OpgxHXOzQS86Z9PpTsiTeteGV5
PUNQHGklqEIet4kMjetvb8K9teNsF7A/c/Q6xUXP29M+eKlvZ0iv/HmPG4LGcm8mI5xMFLAdnnRJ
1b5jrayl4gMAQosy9pn0017NLqxclj2R4MOPBlzGa/34EHU2TL8UamPRbYWAQeasiKJVTHW93QE8
uXWl29nzJrR/SOfNwd/KYCRLrCSGXl7jI6wejFziQMqJDDtuXJgA+QuZ3VtyXvxNdEHyT7/3GMAX
2Kooc0gNl5Rk7GEgThoqZl6MZGW8TrrImvdqsbxSuwSKlSlmEFBWC8+vEAPEnG9wCqr2WrRgqZQF
eu52WL3hQ3d8TOEn50+0NiI8LeJGzJZbHxXTtsUyxcik6VcQRQReWECKrXlWjI5iWKRWZUmEVyLb
gLPk1LZrqcfraM57q9qFx8sAtoKwvyD12+iyrOpW6P29aCK+5AIh37PrIg4ofOsJvxHjLMyOMwiT
CtV3GArFlwz19fDE+PzgZ8gGV5OfXf/gBU5xoB4+WzVOx3Dg9XzI8m0sqvWKRQFs818DAYOHXYSP
YQdOcJbzCd/xY/1hqHGYF1+fuVTy/8pi1Dm+fDlt/5ZmrcE2DleUuZVpZJf1cst814423c7paMoB
yKw9X5u+iODo+qQMnqNjFGUgPGZQHVTfuW+66Jn9e5Ohf6kEDao/j8HyzERmHMKMg7+SYw/0NOSH
DAbtazgPpNlaW/E8OW42WYdnUhD7fj8arIsZhy9uLcRUz/NmUuBsMG/1uuF6HZWKZk6aj4u5HRFe
hAoscYMFELOwimHnHSERtpTz8PsBuivLjMUl8QkVyLOcwG34Q3XRJ6olwLrl2mrW5t1WjVKNhQZU
d3YO8Oy7mWDMijUTJ1IGtMNh61ym3Slt7bUt7sQa4Ie/u377KSPtMiGXBnC4mKteh8/48tcF9HEt
tFlbHoYI+4KpWTJX2wqezPL/kPUCza35Ed2IkMh0awWAuXtkW+lgKC13AYz4cmeVYTTEr8g7r4r5
PXQIDfQnocnZBZnUoF7t1HWGFYiHJ8Uw+MGOqzEqdTkg/Pyp8lr/3WfK+EaaGxrdN4/i6RE5YrHC
86As9PbqisaCRt6j0wEO8eLb1DtvDzTwFS2buUqYXoRRPpblhm6vvIVNmJLHzN1miakvPpx0HFT1
47UoJYQptzFSVt6ZuCKDup6CRB8oZRWSh0RB9xB+2LQfGbvbMwxn21INVG8Lz8MXtEhLeMPVkn7f
cjgYsGijKT2J+o+2nUVpUEJbL2oaNEZpRtX1fqhtmhsWlJ53uvWAti7zLSHYR3gbCgJclF0/7pFd
FkNTtLahT+hv7KcpwSxcWyBslZc0cUiq4ssmKsF9uSkg80sj6Z8/bw7r4VbUezZ+oUXCkknNUxub
71g6QdXSTOYcUkmbPsfbdPYEeOqFJSbI2XhY6wB+hRl44Ber1MDD001wgEh8eZkJzTB6XyaoTSTH
Q7DQ9gswHCDD5nQ/f75d62ARSPI5oi6Fre3cv4W+wDCF6YjlShSGAuqPGNTMHMxaTzsAiWv4IKs5
iKXjnkLJR4jHryQWocnU+EEH1aXM1SpCGp1JLTg27zzb+uNCQ7yoGizYY+U2Myo0kOsuvMrG91oq
3pamlZxZkxlye5kKWCTqX/aUkiPJoj29tkJg/a1VjUJEkn7WSpjoSVcXyzzpjliE1ausf0bEXsis
04IJRzZT+DW0a9KO6bB+TvcmB+k1tbwWcV7wWd3OJNUYqXApvV7USwIrOQ/oEks+saRxlqT2pQ3l
7TNlX3pTV+h93oqngxZrlPo8oe5WVOIJMNunNd/zBH5vbLoO71suQlqWnju9gMpQ+Rglh+JomSmI
Q4sh+6hg4mFgmwmu8vJb0kW7fu2EUfbjt7FB0yMmikSwlovxPLA71w/m9CRsZrH7IKm3BZFoDpSW
lz0Toe0RXQXksZ2ZZ+vH4PKN3T9br84e7JTWlSfkSX0v18t4tiLdq1AlLLsGlsaoTi5jsZf6NbgL
wDpq6UzF+WEYTMF/L9jJ4JuNHfPCZ76NDAD4c+8l5gGxIhyj7sBws1QAtgY1fdlVxfsVn0I+Xw0G
EOBKS5Ot3UXnJRfprEfcFY+EbTgevwdhVUqK9rBTG35UigiitYn0CD6t14zbt9lXizQ58WrbLHDw
wtTV2p9opl4I4k+s3eFRom91f4kAUOXE6bD9C5rOX5KX/DrhI8EmSh503ktCalpbQ/7gAHQNdfRI
7TRT6a5GtiCRHwV+5Pk3lnuQHOVb3b0+/8ibLlmlB1dTRDJJs5a9kFSh+5WXgl4RO+VYrj2R+L1A
vqqCHyWNTbX4TkPumxzlMiyP1kfiTybfftZMYU/otPJRKXaG5lbSUK9Ozd35MccLJU7oyrAlctvC
dzdADSgL+LiB/tKDJey0LRIs5k8edomshm5QwLGnTVjYRA2fiOw9kMiwK7UJmTIF/5GlqvDQ4Wae
0v9vsa5NkZw61WeOnvCmloeyj9vGVvYnhKxsvFdPUfA8RIQJ4xWqj9WH5QYZT7f1rlGRW2j3gthb
v7JZGfD4ARUliOmorPfAgIXDhnriIxOspBy+v+H8teB6Gg88czlEwQuJOvfWe1ZfMKk487zmBV/+
8+mX6sTU+kXBs8Kvxz3jbEFXBrLMvqwCyyGwPaovp1s/S1BnT6QJvsUYMQ8hqW6qDYx4H5lagHmy
ppGWu791kYByXOEzb9qxvt9UfdGfF6BfxW6jjmOI7rh5S7xgC3QbQwFeVPyL8Dk9fUUgC4+o7VVm
0WA2CswiguQk5w7+lAsBQIWKJFsDkjMshXxRGI0vJBQCV0T1VT0BKC2/o8+4qq0zwhgaiEsRmVT/
PrRygwwEVgtVXmUR0VOsFIaFg8v4ttd8h5wS+MneZP92L01e1Xj+Qesvs14O+q2DsjrXRmQSTbYm
8KpkLuliJwrsIq/XPFGGud3cD3629trjPzAcoUn5gQyzTA5stUF4w+j9WXgFoCOt8Mdzc10ATf07
Pz139YkkrDvX4NlIyCh38jdt33OhatukVivSR2tOwwRHp9PV2o0AGQ9iZn0dBcqAuYi/yAPOAJL+
P+7/DSl6Y4AXdUGtfOM8RogEhMR37jG4koU75LEWAlzLKxuLF45zXEN5Y8oQeGGDoGYu9xtMx3a2
HLSU3hl2vKWAG3bKw1mMTB8j6xZ0STxmTCsSHZ4FSenvdXbREP5qwQeQ6GvieLA7hfTP8FPWnrfU
D0lHo8lrcbLFmUWwXQ+ZDVxvgovErJlGR8md0Bw9bH73VPkNz+DScO5TyCZr5Msu+XJKFB2HuNOh
D4nKkrtU1rJE9wqC+Qf36MLgr9XUu6031UMy7thcJE9lnLXzIXdXh2fb0+fxC98wTg8Xdz+KCG/z
hbs03rCDEFdWEJLr0y+DsNxpCq6Io7Yh7ULQY35kpuCPopCNVJPlYeTk80U76WPBEsnwA/xEwvib
nPCHDo16DGk6KiMcdymht0UktSsXq4sNbkqzr3MS+VNeK8WAds78mM+fInx5JM6exEbRlgtluEEC
lk60isvtNrz0+5LsIsv6rxHzy2eoE0ZgBt0Y+kfu5CGiApkbS4Xa6DqJ5/EBrg9N5AB9qfPt7wMq
RaShyp4AfoOH61DlfcDDgqrHSLgcEJsWygDUF9L+322D4IySQ32I7uyW86L7urNCoobODKBbYfRk
yQC1qdtTSpFngnJE7LNDieIOBoxMbsHXlLejhu69zZjW6IyHvZ5R1m+cl5LRNC5uX7KvcuRWr/PE
d23TUPp3KaRI/neEtu1jevRQ6ET6/D5kPfk5AA3dhCDisX0qfPqHv43IDvWX34gyUb5OMS3MJeEr
CqR+n/GphJZ4Gw6nNSoqSPICz50flDhEeAwL8ICURf2HWWWtar6y0gMM7NgCwePJUDP0iX9yobM7
YN7I3QeW0yIpWgvWp12FLFqygIItA5zG2AywcgBM+62fge72jDNa17nx0pFLkLynEfD4Pnlvy3Wq
M/2fYlm2rGrIsvPTx6sgt6f7n7kZeLxyRAWqz0KvAMb5fYoWYbpX844Z+ya5veU/qmLxFFi1MwtV
b/Kn0khCAh9jPuMXIFfCqtprIX8B277xh6FtLDC+TFGMir50PaOhtjNdqa2G88BZV9b2W56gD5Uh
EA2MfU13OZC0o+6L8SnmUNluoyBckZth9jIia7HWKvglzQvzDZ+pgYIFGqou/PVi0degu7kkx4oq
xSvDOFINLe5tVMlTcCB+HaAi4/yaSfcOl4oQXj1PEwdgp/Omdz/t3lcRtPUEaRY1+WALBOeJEtWV
II6I50TX/g9SQU7dHiMI5fNU0oEyDq51TCvg6QEcbForTUKAAXk1jfLLEr4ZR0qEYyF9923fnTo0
bIAhJOKJiHjfVbGFDutsiKbJ+vAdgsU6exMJQ0wV/IfQH5ljLdT/VqvEPpa+L+VLcRyXtovzIXQu
uGCDr0xSgGVN7+gpQmC5ZldKVSKhYENIHTQg553svUXTIfXnF0DXDbjRNCn6dEsQPMNxnbnHQ479
h+pt8t9l+ILuU/f+pBmVaKrdqp9Fr/K07MEE5yqCE5dSufpdddoMJ710phbJIESS1A7kjB7ZLRpm
mI2g85L6tz0cX1w9FyDYxi5kOkPXKNwnn3Rno0/oCFaGKTBHaLhS3uuS2Vi+LQpSrsRqlHu4gg5Q
t7udSQ9UfCG5xzJMHrpTu1vmvNEswyFNI+Ji92aZeTVd2rP2GyWoggysH7JRERXCcvwfgXjmAsoC
83kN1+UKdQ4YyGmHzD9KzgWweHtRVrIcPu+1SVES/TvGeyqCjSFEs6f+pwMhBnI8yyw/Pzoy3vrp
ggNN9nKVSqTwxAqLty7HSMGHOXcSdinqcbsdG4W1PzJJQCj17/zKm/HAaFjqP+BfkcUqvaAq4JGb
rGsICywYU5tTqryHjVtcnu7t/P9/BEkkKfTT0LkEcC95w3nq130T6eYVqwvI3FvFa2ua6naUoJfV
IzubteMW1lyuKuR5+wsSlCHTCe8RLHR+5vSxpOWlnTYXqEwlnqBbhQrmZWsb/9C5YVQwjwRlHvYL
5uQbqvcCXIpv/aw6R9QPPFISQIdyxdC3eGCGOBtWowSFU/Y5nLthKWOkRrqWT6Cvcq278aYrp6dV
mYhLrk4fK1tNIUix2NXTMU9+jubgE/qUoHjmRCAWoeLlX1n1wgoXC5hQKkyatZJ7XroXy7KXBPeb
l7xDwVrCfpiqcsgvGvzydbIWym1UZM1oq7dpShWs9EZCKwllPpUzP+sVIiPc9fZn+EivYNtSKP8w
cmtdWIV5TbE1Y5E+3Lq0JdEs0YzoniR+XbEUevkMEVgrE1xWGcyKjucG5l/QNlO3Q6qITLpDUczE
nIVjtW7K64+rLNFZLIBvArJGrQYcXYF4MwgzCMLALLhTfOCWz/aYd4N3CvtcFxKJhsX2Ut4L19zC
GJPjDWmtUgZi6zn8J+or/RuTzhxwSYT3kfAap3XbNlSP6sb8z6ctJrR1lcE3vMc4ZCzObUSz59re
uogp0Ot8gYVyl3p9TJhba1y4X8+QyBVO5dGDWIkYZ89tRjzQp42VdsRfb9mtJLlVa+rYY4eCWwrY
PKlHz4834JPr5uYy/E/0QO/HE8wpusolIlBnEqwtGb9BSYmtR8JOOtq55/IUr1kzalLaPytnVdru
VMy9o+S4B9Rtb99EYBm1WaHGhRG1k7J7hRt8C/FFgrE5mwrVVJtpBOZUwOfdsIcR4+lOObGh+0FH
MzK1q7y7eTxX7Nhw1C8sq129WB9a3fWndptTeNFM+MhSQsLDEVhlXiTY6MUjeWNi57Pdar/4N5fU
XqV7s8n0YkoHvV7qCVHni5lGh8uv/qXznp09OeOXQD4zIWUic3JL+KJFy5mf5T8JdmKVeY88/Wnl
b6SsBts4k6R4FDDYzlZy1fSLeKuyhc1c2VZ5F/AJEmbRI+pUx5PuHEVFgPxBKjZGTDWx1gbhLCpD
/m0KLR2sAyC13BJ3hA07KwBvfhA0xBppyZrHXRFpFTv5yATxTIrrTzqP2iFbrc2b53+V2MsQmoK9
75a6TqJeiEv+i8eYr+0/hjhfq0aQvfWWITSPzwePniaxZ7T/7glQ0kJ6nFRbGTzfadmboQ6SQKUm
Yc4mEweNK5EcLOUQkBm51phlla6ElSrKQQuMlNNMDQD7QtARTrppR9ApmDX0OJn30yJQ/19C0avV
B5va5IsCgywIQ83/oSZNYFJXh30JnA2mCNzAaRuyVQmvy0QUiG7zLk3AMM1cgSQtOt5tb6G1CG0G
DU9WPhOLrfi5u7APQ5j7clhZLHnOL9yWBGxsFNU1uQ9nyqARAIr2Kl/naofpWBJqkwgHW0iHlRTd
k/hHMP26FxPoZ+yRESaDneeNVX5+mj0qqLc31Hqad7SbIDqOv7PEknlih3VX/AHDYT3N2GA+fClO
osNF3KOnlLZ6yyfBwSoQBzyV7wU6Tqe9tyq8jVq4PMnbQFxhlHLf03GVDynGo1QQ0vECz0j1Qx5M
SLB9mN3y3PPdMDx1loao2GPee6ovlx2K6qHPXnpnX1fmludA0NwIVa1zrJZaAhiRRo71ePUqwLIn
52TAeZ1nBTg+AgMpFlz7+ljN+4Pk0thFpgT7M5kFMo0SNmowokb1qN2CDTPZKr5kbef7bjrBNjsM
xq+iOM6u7ZD+sy6ERkB59oR7cokq4aMnclG/ctFPCANIUlSgJV6777FZGMeTvrY21AP0E3AHQ0sP
lbhNUtqL3FLIms+gLTpJttY8+omSCbEa+t/FobrGjfOfqT2ciI5Z7cyJ3yxfqtLvbrsCrb3fG75k
f7UQvKM1/5EOsx4g6Xm1tTCxO6W6s7Fst4Y1L7lepPVqZDZ8+vCci7rAE5OnbBbSdeOQxXH7mFZu
OL6zi4lOaIPGkjZGo0DFW4tzc6gIewhNXg7AkYJRYdvkLpDLAk1n84m6DnrZlmRiWVn6gpuWsBck
UzuAzTQyEOJxGzTZG8o3cHFsWuNEsu9TSERU/ck1p6xfhoZGWMNyBXwdKomO8iCMDosPFEVv8fyW
gL1WvS8JyaynxLWzeU2B+G3ah00AcSs52q6P6/mUvjc0VR1V88za/YZRNVWL5xJW/WM5kLFecyfw
Ul6cJLvanybDpULAbvhQp6yseRRGH5mulBQuYCQCAAX0NNfe7/V/TVStLCFbb72ptrqtkjgDGGyE
fjYQAvwNShht00AawNiKTF/n7myscPKJA91WowHXJ1gv7y6kgbonGiHIAitWiHtQz+5pMZO5d9RT
urjcq/itrUtbT1QVkcsmhKbxxjuKxW2xP+5A4FLQk9yrU7lsXcXt9ia7WgQZvQULWH617LikJER9
8iTX8TrWwBSkp9nIVAH8rrBQwkW31XT8XMpsjPa6FlLku38DUgtz4td1RSixDV5IoijuzD7wpRNK
L60Do3/RzZVBy8YgO7g5wjgdcdtA9FZgnnvVPs+OddNkjoqE6KVEEorPLZd/h1ybR22+zSnt5B7E
Jskc7GMffHFaDJ7fn6SkeKoPQ40u29vQ1emkV3nTpZu23DhS24q3vlhXzJVlM6skQAOV3yM1b73s
XLUAI1sbSeRMDZmOwSJBltB1liI0yyUzMbTRhmDqLqV1Vj477hIJ1XlGR6Xo5QBQOZl4CZjEbqjf
BXhXavcNBUpsaXZFaCefdKHuia1LUn62L2UoxuXFzI2mOQrG5dlJgVjaCVjmA+DIaz8NryI5wvu/
co9QkD7XGTQ+q+5l//LBWur2yWaJWnTPYYZCq7Vpzm9wmTRLWmXIfLSyad41EOxobTtxOd62MTyG
pZnYIFSfHi0DqBjLVUBD+RT4y3mvGuJkcGZu7TcFVGBaHABVIhTf+p/1Wy2Tn4e9rIZiHZbqndmk
1A9CA4Qx8BYp0E4KKKvQLoQ1m0YUTFoa5qroRxAy22kua1weoez4Px+Bp2GcwzleUcRExbmPEaQV
rO9dxhyrua7AoZfmiatHa0LskZoXAk+eYlAZVD7VgDThm4zsrjWfXabkmEoxi5gI4OdIt4QLebeN
8K3ATE3jZf1pabeI0tjHPN45clDJfVGfpB/fNdFkp4W4Jgy3WhL6g6eSjGC4+0/rPIc6ifRZZftG
yEEAWFKMa9Rek0RHj6peG+QsUVxgDIDmCdc67OXfHESGZ116hasBmCLI1ftG4X/9D0HK1dzc8s3/
2Cj9m5/7YqOmZM+XDYYrOWBokANykXsz+nDONu7rPYngXE2e4E2SDlGO9hlnEJDVR1Lr//8FCcEl
qSx3HSoxQcMEEZYTbMFzrAZB8UgAXXbH5al3IgMhFh/CfspkjAt0/ONcvZ32LvboMC/Y9BGz76az
Uv9OiokN1pJ2BE8P4VQ5KzJJwgLEuD/Aq0h2UOaIkgAski0lbgXgL0VcVJEKPpTM3FJIIcCbBR3j
A6VGOfRoyjBe8qbCDQ9ovbZqnNmKeHLj88RYsnREnQr3+IEjlDfj3M5YtNLufdEn77RSjd6zQM3/
LVTNYS6sES9Xqi+tbThTJRhhX51PEgqWjQtCTefGBqkG7kDNX+4mN8aqbPcLYh2i8AMXKwCbFRfD
jTmzuB3AOjp6y+1lTPKTZjZLrEfah96TcD9z590/6AF13cjEpsI/tXFhzzkryCfclXufIGkyF8uH
na9OSmXqgheqmgy+Y5mtvaEE9taFuxJepvGIDEMA3apPRUvcMoqhrnmGy/hscjQjR7PRL8Ks4y1u
36b3ziIS12fFo8W7BLBqH/QLiwwunbC4XkNlsa3Kj/i5TF49fHmOPcxfH7YQqtsIrnfh+Bnr0zKr
zFSEvBGnIqQfj2ndtURj3ZKWeW+yQQ/cMDKFisIcgyjNAaaFsge+Gxg6qEdzdj6NqKMlQnWrOYAq
GQm1PjvXFD5fa7Rfr78+N2DwEGgaLDgda/HoISc9Y9Vj4EyumGFPHBDHpY4ZVO2jgTAT7NQwP+OS
rmGXLzCKrrV3kqQcW2xJcOcmfZ6X0Xp0nrMTRVXnhOegrBo+8WHkeb5wRPJ5Hc0S4ojIrkg5peRf
vdrVVWKVI+sockdivmbodswVKDZBRoSpjq//ehrTUI0thZBPDgSJp1qRQt0ErcNdlDzPRZLJJvtq
lcVjoRIp4qPFXZPr3Z/9whMJaOY1y8KvXnQzDcqqjnkUS3IlPX0yJanAt2nYjRlgvI6UVIIylJLw
WfQANwVOUrt1siTNVz2Vwp8ppVXPJVXBudA8XpTcVa6IHga0Etm42nbaPwrVPg+ri3enJbBUT1pc
nTUmEbD8zJ+BG9lFrnqK7fsVB0Qwx4OUWTMpnj/L2ZMyvqaSwbOJRuV1WEt1sy68Q/LwyuLSbffk
gmp0BJQL6hJDzcPfYt/AxBYHbhHzdi54ghR8qfqPNdZXSFGyDvP6IDQDnRenQ+yvGwlJPz71lu3m
tha8WZHHl9e9GJYPaaW11YAwQMVHQ89FIgb5DOOtEOsq5apTnCKX6gWij7A16f2+gZHhITvzvuCS
RXPdjgteVhZ5RnaBBcrSbEbRwccQE0N44h82K3NRKm9U6hMVMfQg1M8Zy5zGd/K4KUF1WG8r6EKn
vay4Xc0wWKAW+6NDHGXX7gVjdAnkr1oG/93uj6MpSK1zFOSjx0L3SJVNweoANOEp4settD844gEI
6et4Zwuu37Zj1uftYJH7KBaLwXPxzWKxjaEO0XLu+05qpCr5WmTJki/HhmqB/MD/eX9x6VLw2RYs
MssOeNng6Xi4pHTnlp2mm2mXGwWYKuI/3taKzoge9X3w6LTckVPaVYBrPBy+kJwY3te9DisyHTd7
r53FokFrCyfsQ7RZpH766LRGqquNiLizqkR/t8otFCk0CrXEzzeVWJfJK03fD2+ciV84deCN410l
Xbbb3H54Sy29jXk9tAFNULGex6oKmAYnD1otH5BMt9NCmJy7Ww49kjCEVlkwmOY4YrkIdLYTNH9n
yTTbRhvMNROmY7YgI0CKb8Jjq6KjH/Xvh1wlYhyhgSlXp/ZXiHwQmzsRgpV9ZtP6qTMzXI8hj/bR
WH/8rsbjNboYiCMFV4p5nyGY1FmTpphXmptrX39u6h4vOlYQIhIBeRqkVQ0fJV+muG58Gu/EZAIV
2D6iDnommntoDD+84NI3aib/DIINSUpYQgftlJmmDeFBaZ2BsfTKqg/EXuJVNRBd94EYtBsDv+mG
Xf8NJr06r9a/mkCSQNvHCf0RwrqiPem+P7+6sMnVMYn5QpDs9s1BIsvX5lknK77qriwHliGRuChT
13JUSToO+0+11Sceb+gmxfmErgOl29I76yfFwX9aAMuZZFfhOwQHRAQxwD1RkcUZUR7yQp+E3myx
Lv1q0RE6Svk81cEvtRWSRjJjyTSlimC2Izw8s1koC84rEHUfKlZ7IpKnWi4MnIzV3CDL9VsSzyCd
mCNUHdnzlPsf9N0Vd3hl8Dpe0y8uDFb3dbYJfk3ZcR0YXB9KLFd50gTRDR/vAI19yYMP8xXuR91k
NhP3lcmUwhniBoG8uYC/Da4Rb1LhJDmsKjzT+804TENevslDlbHMAYYxmpWvfG1zrlBTfUOqJrU2
/PwGMIxWtINQ/BpSk3IeUMyiFXitFdraKo8H4tYO4vG2Oorj0+HmuHBIese0hrso5iK2islPSMYs
ql0N5uPTLBsdmj0c3XCmxUZSSD94e5wfd41eM5tpvYVmLH3B6OVUfrVWSjvo+K0zxY5NUAh2rTQk
Wn4diK7tKiXA9K4GKN26DmaW4O66DAktiTt59ufbEhexZfXN963FYdXCToalk2deVfXLcG1J9KfU
hVH430EnyollAglB1fQzvMZoCSUecG77EusAeq2K1FJ26VMGdc6k2FryqBeImB/ibeHLhjeQhUX+
ghKt89oIY+j55DHBy3NFh2DzDD3WW6Q74yMJoqM9KNMhE1uD619SjwNsGmvSDNv5+m4+PKaWnghc
V7ndhuke/I+OxgymX7Vdx9iRfSQBoheVDzgdJsGN7WiFiQaauPbAeCJfYsY5FjVgFXKTzDFGlTqq
2oiuVdbYTV8Zink8pRd3+97dLeFDpjwh5rhD7CDIBVHWaU4RcmfG1zGgECm+b+V8wqp8+mLgws5j
NHHQDXHufBsk7ri16oFvqPfAEOAB9KyW5vK7hLNPG9czpGnHV4Gki4sm3fu2hXtKhYnZKWrBT8Nx
eJp6PUgFzJEPLqZKET3e9XY/FKQQYkdNrb/VPjIOwRc/hKKmNPoA86KJ+uUOUaQaGSH9zXxk94+L
GSzDdivAXJYI0cqf20Pf0ZQoPjq8KeMnGBNTSENZBeUNAUsWYGuL2T96QKU5AXpA5FotFvaBNC8S
+2FmsrWpbGyt20MzwQMOAW9d2lxAOqGWVppWEWRCnYA5jtGGt/TYOhEMDHeCIVz580Ud3C55Qcsu
JJbcDIN7pPGQuRdmtcDVYnLQksv941ziTFk4pSlq3zQyTn1ZO3vwsAq+NchqQEaMR5JgdXgRxQCx
5fFFpzYTKGb9WlMv7wIu2+ubVBWNo+Hr9A8mWorIj4fd4n4zMZUIfj4BgunjZWGbGIeOaNDstOiw
I+n56izJ5zAvm13LIBgnOKdopnbnsaH6eJFn6gerSocCYYNCwb0YEjhV27iMLLgIMOecbDC/Nz9e
kID9rziH3IjVcH//DYRPZOsBagZ92YVuDUNj3eimV+K0FS753uBNRrLUEP3/zB3xQkWqF0W3s5dL
qUsjuI10nFrcIf43jRSuq9QalOqjoDmnO6ESjWF0ri90ynetFdufQUJ4USPzs4uckAF3qyUJmTG2
TsO2Yuw/NmtC8fNt6FVPHNBx0f6PE/JfQk+SeYYt/oJbVe0UKVrpYg/CuKyfNRi+6nd9uUh3a1xq
F5UTH5Aj63vnLkqoWOOIpoaB24UdMbgGUa6s8/6wyUViSK7NW6h3+SpLQW2wTNv5aNTIfgWZrqbZ
mev0lkSGZZ4L5Rnl79Fodus1z8lakfYaS2NL3vc6n+7XjzHg/cYy+MGOUhVQhR21ls5SXT5f66YM
9U5J5klJ8FB1b/Yip6hfiBHVCJI7qbCIpnHk9ivbhKSzsTQqkPsVy0bhlKPzYWPv99/hXJH2SkFY
EJYAKAGQkeCtPRZjgVHUzi7Yoe0kl5OlToouAXr0YiT5uQq8jY1a7zPhmeZsJYARH4ZPC4o3/aKm
YiW96T463hdZp37X5UE+t4E6O8/mjkdJp5r7Mi5cq+sfGFrZQjPSuB+d1FSCO+YYchHGvY2g73Jw
+yu1OZrIH6iE/+z4fPc3PSdFrfjizNJ9oPgrgUMLakIwjb6WaqMtxw6JJx/ESuBx4L6QE4cGw8fd
MxWNC2dgvaxTm77szaDGUtMJ4zVz1nnUwMMikbBB+O3L3cIDN3bdNAMLQuKTanwtR0yOKWKWS3G7
ZdP9kTKOKI/YqRR55qn2yQsK+nrwyXfVffkO/AOAHOMVt/zBLgv+s0aJsjcH5KbLP51S8KaggjeV
97uozNtM7jdGZyoQ7Ch/lgYrR7BhT+oBFfn2sBJvwq0NkJ3jxKSZOJjjBBqz+yOINaE7mX1DS7V4
mpevh0BlmeSonP4IZ+85Wazb3IGhtCfog6EfJjGswWs1F5uL2H/LhSJ1qD0+a7o8eRuLZs/Jx80L
D0CSN1lmhIyNmxVXg9GlF5jW5jHO1IJaG8xYSjPgcbbmC2BsCyKYuRwgCCJ7Ct4SnVp50naxASQq
b7mNSLkmbwk/Qb29U1HPGth2r75VPayNy8zad0cqdyt1MZ8xXIcWFgrFB+S9pFM8D2UCofSMLl2I
ywvQVgvNAQUM50jOWj2KdaGFSvIum8aYxASTw87l5GwGPY0XnexZqdUsxERYWNdiYm54G7yNnVSw
eVDNo30Ys8oAPNQk+nUdUwUsxzyvbfL6Kfw0T8tIbvnb4cUm9Tj4DBKB1Yg9kvw0mCpDxnkLHoKU
sl6kUJ+C34tt3UZujhu/mjzq+NqlVpJ1QywJuFlsSDF4S+fRRC8FGkFjRCL3XkZ3CfoLjzTLsZVz
tcrjxvu7PIHSshRDiGjWBd1jWl49utubQ5ww72ANUtc36B0lT9/4o/XbakHv0m6mxZD9Vyl3pZFF
lIhKpJg80JOWmFbSZU0hr8z2xWavyAetakLm8eWI5uFxJgXHSl0O5C6yNuyi/8b3HTlJJ670jwpi
WcIFGbc8ua8NBr6W4Lnp+8wdBvDMCOOG+o+uEyftiXKG048zuzCho6/CIHFuS+AH33ZP1WhHEFsp
6ypOIDj5XWT2ER1Mx1btXHPoy8vtaX76+3vfeA0W6/JT4cGl7g5K5fdp2J5IKurwoNWi+97InofF
hED0pFEYE3ic++bLBdsmNYzjLWBioGEGLNmXxf46gpCSuOtkViBq8j1TKmDafu71tM2aVue1EmrE
onNhVItyQho6r50xyQYxknbsnUzfA3XM99aFQy8bhPw+I9Bb2rhxt+YuzncPg08Cre9dL/KaQyCW
HO438orv94GGfRTcD6jIAKpWu3jDZ3MCnDGHiJKxnBwH1DWyHYuVyG3Sa4o/Z/uBKy7UY19FR+ab
6Tr5zlxHqvINqwAFjR1arBcSj+JVlHHdTHwYr9WThiyBJ933XxWKRI7HroNyS9LHR3mL0qDiVHeF
2jq9NYmyMDQ2IP+DFc22VVVaXnE3akSKSjWL0LVIvOJAVYVsHwv+NF0alsozTqShshzd5Yy+sMmG
oOebDNNkxMBmtjrbeO5EHSihdPaOi6T1BKRxOkEGItd7q2+4zxdI3tejn8p0+VjlyS5cY5ClWGN1
14tVUFrxpN7YgLeV1UDgYUzuZfsSIVJxPU5OdevRBBv/p5K5hnynze5Mmm/nj+nag2e2f8g330zq
Yf0qePLHsWGcvEvMPz+KNOQyJgmxNxynfRoUa8d2JyHNHWjUV3xXmg4/SrrEqEpOlK6sKWUMaCfj
mrwg43d0Dnsv1x/c5E+Z+gv1bQMHUwpmvFxNFhovvB6F9VHPTE6ekGqnMjJl93k4lp6pyrny+hW4
ISoR2dgzEwKSWOEogC0WIKy86Vm896XwHtK02K+KUVaHfdhoHmbkoGjTTIU7J0mp7cJV6fqx3VlT
AoOq97DghGreBGj2NnEyqvG8frooOySSked4JP2gR99uY5nVqShEdkQ/Kb0jO9Fn1bivPUoOIZE9
yx1sQisgzOPi2jkXwb+DzItRc9gr5xepiUbKFRtOxpPn4E+mrhUsZ6hZF102AKUW0oG7AGShR56y
AYpoXBuRyISxauUxLuANwIlaJXYMI0MaZuiX5TSSE6RnBX9kBwK2CYXbGBFOaosgx4EAdK3cHDyO
YrEGDfRxTq5tEPYtEG1XglnzwEbVMRTWmf95+uhkO29Q1kpbGRhvi7ZSOREIraoNN6svtTJI3p8H
6PBF0vy3IFffLyR67Uxx4jg9n9DQdIkeyGi316+LSGoapqButXKkjMhdA6Aemct1xiSEkxk6DlCt
JRs/y+tv/RLObluEpNuylxqDd0mzEK06tmBo3bJapBj/1l9JyzoJNj68WMxpCCYJyj4Jwct0Kaqh
CTCauoz7ZfdEOqflnckgEv6PoSFRLJQCtL9yo4waWPJmhy17Im5drvTta0PiR0cvRF8M/5nz3c0Q
/IirfjmO+jz3S3LD+t1imdNUfPgqPzVf11B1k1RzU+iyXxvmILmzMhEMum/fGKidOC3slfdTuRc2
3aHCy9owy/m48S3Nnoe7Dm17Pw3B1z+b4bmkziZxyBmBKxL7HOLo6Dt3ORqG1bgVVZw96BcXVhdy
JQO3tT+Wdkew/gmaziGiA2iLMHpd5VM7TsKWic8/LW6r5V/QL/1bhcD9y1WheG9FGRWv6IZS0hAn
6VeYdEJi46Nj4ccmVHRmiasEiLDfbozTd1pvGLSepnZXx2ZmTjK9vvB7sSqq8CmHN60LW832HMxd
tH2mPuoHiclNKPFcZFfGtn4LcmhZZ1oCtRzRwHLIghd0sHeQsOwpWB6f9kY98zjWDFS5q+9B4So3
ZQH4k2vl45sOcIV4eB3QtghNYHV+Yhy5WJnJ8QdwN3e08wFcCmxwUg5CBIes8ivhmUUe2Hrlg3Yt
bKaFIR5bNdPUPtdP41OmFEFwkuIViJ/kXdjpgGLBeGQcHa8FVWwqtKeOKYYH07mJhDfKmXIskqDO
XFfo3xepHbxpaDhv2G6U/w/SQfXcPIEW9nQmgDUblxIAr5mAeP9VFW9h/2zd5bth2xZx4xFlvR9N
VazDECmBD5x8o/+GRyEZerURhpUnjlGGXp1zWGvD+JwEDGAnflyyisx6zo9E9vdDLy+tK1lmvHSp
oQ1NrXq4fw2Kd60joS9hoe5NnkOYEPdZ9ss82TkDgv0olHYODRmFcEdBm/V8/ZR1CzW57KDbDdRx
fJptXUVXsET+KI5dBhhompvtcg4FZmO6/7O/TN0km66eYiiB6lpmovMuPL9aGWPawy/78y9k3VSI
heg7/RIbuuVqqy5O7iXZEKDfLX8GzH65z13/HCm+GMJQ9UVdQdPiL2qOn7SW7eHHRrE/TnyYvYtO
6ZjVh42TzVcxiil+GF+2z4asQAULCPVsFROPqxziI2ijAOzMUOweHJfQUaCZ9FZSVB5TihhFFOSC
0qeemRAH74E/Z+vcROtN2BAJUQdwnpWih8MyOIuidgyOo//6fubwlBMKr3YoJMNDv/or9Nlw0WFC
OaiEVSJ0crnM2MKl91IXaqXbC25ok5uudwSzfp/VvQBPoVWG839ZtU3LzqoeoCsGQ7+3JrFq9DIc
FulOYbR39JIMqef3N2HvNAHkjfE74M2Q/YWMJYGkQUdojxjEYoRRq/p5IJtTGbj1Eg+ouJs7tHjD
q8oW42K8NtzkSPJ5m2agAWcFXQdBBFOneBNtHT4UoVJA9STNVUOXGRopWx+206tpVk6zmpWLm9lU
GncTEmB76pbda+/cAkpMjHW8tw168Q3sqB2mclAik67iRd0vCV2RH94T+xXum0Lcm3xcSmGvpmqx
N57c8FA2njAofDQ8/nESj2z03FtkRz1eNrcpFcGES72j5YWBzN1g4nntfkVT80zJm66Rtj9NKUJ8
aIyvCWZ4UOO79RWqwNXhpJVF9K9fBl6ezpJX8M8LL9xyDVVp4ReRUOQXj6iXkTjZzFcgnqTRhMul
OVSoqDV1Ca3LbMIXX7nboqABRIsa8viynN6qZ8WMUJH8nIBG8QUhMXDyH6SRGqcH2pZRUxYsi+zc
CPNNUD6vbj8x+iWZP9lVITyRdMJR1K9TVD9ZA6cCyuegpyWTlYBGV6jbt4Nl1X9lv2SicTkHawrJ
RAnbciAOE044v+eQEPdmm0dAKxXrl6DcxQq6KQPkim90rrAxCeTVskvl0+mwEk8pDd1wzp23QUVm
OGZTcwlspGqlUHFveagUVnyk587r5jc90EsvfC6IqEvyUhMHUjMmW4XfD5KtNNNCFqhfsB9XC5MV
hF5nU9Zs4vHd+XrAii5jnXoaMs8Srum/zoMBItmJ+7IzkgmL9OEhr67EsA4CP5puqTwqGi9CmJ5R
A7Y5u34j9kgrL3nb6OKIG4ZrrtGNZ7rDLzr3g5DuO/zXxwMqZKf99euv8WtE8WoM43s+wuLWWv34
eCnDC294XsXpkSi212T7sJrLfnz/Z30zRbzmNkSZhM5d9NPGNpPDCZ8eumV3QbEluUbGJSz1FeN4
HeA9Uy5DDv+AoOh2kMiLYi23UXI2Zz2VffzLaNX70aNK2+lPUZijpfAvLf759T/fkAg4q22XZRda
vWErBWZ/g9340Zd8MmQ8NzZW8zkSPR3kdQLKrvZ5LXLTMNDR+70pEMc3OFiF4yqJ84KGBXsz6ETQ
DOPDozgqR/syjpJIn4pOgoR19irPtLsnH2DRsfsaYalJFfkSARNxzqtEDlj/+JIUoTN6dT4Z2o8C
1U4BDiTnrSZYoRpCYkagZGvYAmcM8z0B8Fh9i6qFFo3x3IYMjSkzmL5OvVqBjcJtVLQOCZbkt1qu
WEW9yTp9uzhSp77DAkpbIuuGHqzxkFrPdp6VLEsyClmfb0E6A3zxpGFrVLT/yrMFhFtGtR4AF2wg
Ht8pzwKAwMoXwgVOw4ObQpOqspdpBK6w7Uuooka4+lL8DFCHfrgivo/SntaYllJldKW/dHVHIQNY
pcVEV+0yFvRJRU8jBC1h2VjRxISNcaDLINydlHuya1weFeD2NN+xPVd6SmHVSK975uLUCwD1khRp
tNPyel72N4kZev8G2qkkDwUFPYMkt71vOXzNgoW6qe1dXS9WO61DZUz9k/Cw7kg2sRfhRbemie4u
heUy9efS8YHFFEqxJ37DbCFNM/AqBaxi7lnKTp3ReypcATjceyWqi5nSW9XTRxItIQw+zgmMr5sw
7QiCuzfyfpGpAdyO6n+2EFTtDgUXeWZZq005bLFQGH3wDK25id7sS1CLLxjQbewBswUcpUTO/4ZY
svLzp3GQj1poG7yAWddjtuMMrhvezjrYMrhvftfITzluffEF4IXx0ZjgOgUGNzm73Ka7Hjq+jhbE
zMCqWLeOlDbiVlFou4Nd8vSweBWg2L0P2FmnyRHGppArXfGQbbAf2BlER2JF05lSMWS68iom4biD
kVYSX49P94n5xdnQ6RBvneIVoaD5ghLW/+aqpLH2HnCHIlWNkBsX2CN/2XAEdGGXyLoMCwhi6MA/
zgRuZiCcFWwgFsSd/wgTGPBAmnXcdHSzt0CW2s1OwYnzj8a0UDxVDKZK5rukxwwXES9uBCcZn8nx
6x4GAWks8hDhrgb3LmSfBm02koIC8edjxisjER+JnVYZum1oRD/upulgjrugB+WM9buqYlvYCMKA
KTP72OkL6Q/7A1vw9dcgFi67IMpF631ugRKV1zenKsp+tWbaaatvclddUs0xyIQh8zUkm5Ks01Pk
AEhW+xa+Sx/NuVyeUrDMbdPWiJ/UzPm2FPwx+MWuwEK6MLm9YlVlJ99EB03llVaFZfAsGsxBAa1h
w3j6lXvlIkrZP/LBJ/npP6UNlsDO4gMwMupXO0hMT8Cs1PGuzlmF5QdHvrCoFCTs1GME7jsaAWAO
5CD22sUvEP3qpX5dSDmeoqjVzx76vC2n6gvM5Y9/02YK1Fq3ITW9f/Cj1YqOOXXN7nhaCZ0H07xL
ylkJXKae5IPPZGMzmQraIJftm6SCGZaH4nqJFgtgIV5I3vbetTBFacNYMwpoynAMNVh8t8Oe0ris
nZmQuFL4IqrkY+lrDetozAiGA97PCh9336lHByUtpVm6lRuMRcKBMzpyqNrNwxB1KTD/wuOamPjn
obgmugrMOmur8eBJks12ksqqWQ+4fTMSSELXjvEuJVyr2Q6Xcflyez/CSSZSFw33EgtyIRrzpZKV
fRcNe4OdU+LK2VdVY1r8cV9v+m/EeosWFcinCCs7w3hP5+FVJXvrGaunoAWtzWuVzM6rT2JjYLdm
w/qPs+43y1Lh08ufV+h4JWt7IQgLdOLcHL1OfKSGrNGENbs7LUvBh+8kxC33xvfidfIx2UeBbmHc
gL6l3bb/CwWF77YMj/oB0qrUXwGE5KqMJ2OvXv/uBMP7pIal6i6TORdTjDpPQruoKMpHkpfDHy+/
UhyQH+PWxzMT9AVVpMmPOsSYFUdFz9BCfD38RMv6zmEsuUw3mY/Y82nw2V6Cn1aAqdyWJhUgd9Ig
Q+UJFnca5frMGN0IAuSM7d8HaF2MMU7UUBlRGFGekD1d7OaYGK7X7hBtL5th5ztUSwbx5GosOQ99
Ii1kuH0HpVNNxHmd4abCJcWuidmQfvqg8pTXA84tutoM++wVVd+g0TJVfJ3s22RqA/Qu6Octs9uw
+qBxow/3JWkxmLtmwqHE4/ndOFt0dXAGWrlvPR7qCMzJnyjLqgpLj37IvAylLttTwGAaEzn+J1ih
m5MZir9wpuXWo4hIKKf4lposPMvQdq0R8Cpu4mEXeSN0Nt62Qpq2xsBhFwIUnOo8soaIrS4bQ6C4
HJmcuVf4Dgth2CQ1f49FtoeoWvialuIah4/M4rAPWtuTgtvjWXR005m0I92bs1sUrX4pZyOAaEqB
NcJ4fsQL1kT2SJyJNIVTa+DS5h1nqaTjWmnF+ED6a+o9cpo006blUIlMyW/BJehz1Ypfx0mekZMu
PCeFNVU3jHmf+RTlZS4c8zWRUALZ60mdz1xg3HWsQuCuqGT6Hw8pg4YrWi0VhQympexcAiQz9ZuE
n04hIyXSmepFaP44fxNbzNPX/zaCybkrtujvrIb19jepAtaS96WAPYouM7yzdkKoXkCBxmejubwH
DIirugaHiqpsf3W11iGfAe9CfdBh4p9+DOxawiMkRKyToLN1wa0oLcdIh80kbwuUI++uCoifMP+E
xQ3eCiGLeyAcHs7+sAmVDm5khVI1eAwHf+W8VUYb/GhD9RMOEdx/s+uhZXLvEnrH5CHtqTfRqyZu
s7m6rGHXxEXxPkirB83PFlJlRu5iRsI2NkkmcCYdkjjSt2l/8MMXjWvmReF1wdP/0r7ORrE4IRrh
NOtYnYbVWQogAsHfn1h11n23hYUYgL69EQCi4xqOuXw14wG5PYy8NYlesLSimokAp5LN14zrH7Pu
a/XOiX6xwFjuCot8zAayHJxH3MM0BbHuZhXojp51iMPBX6+ewW7xmAXvU1ZsJJDlPHF50C0X4AcW
qdS0hccXYHgrL5bzt7gdittPIGC9XArnBXxOSnLXfmqsG5Hphz4N/hUQJF8Jq1gglAcd8gqDiKIu
V0uAerTJ1mjzM0jrB3b0Ycx67vMTwQEZg/46nEGZv1F7aZFAdQA2Ae3J4rNgBir95A2Iqqkpg/dY
A+JV/OBsxG0lhH67bEoJ5JMoNhNxI+f3j4pmuNYnxeJT0QDwGEMxQD5QREu8KBrdDASIYD4AYcwc
l35ECJLm/e4j5XP12TS5xPppznCAZkJSbICeScku1hqY0MpOkfCsDXuu3HpX+cAYf2U8/Ie/jWX/
UDfrg3eq6bv98K1/ClDYudFgfcYlDk+oilf8udYGyLZYa5crlOF7WppNmHTPUreZqyHzD6zZNdD5
C4w0ijchdiv7/gYfJsl2F7RStTagSSH6SHNo9Fd5ZkfBbvRAKWdB5ofbb2N2469X/Er0La3osF81
7Eeq44m4Q77wHsPlItWaNm3MKHirj+CypYV/n372k2Z+93c9PDsg8VpHqAg6jYUi/1Vpuffe/MRL
rDKjFoubc57y24B5+qLJN6R3E3wmiZ7qIiBEDeR0TbsBhvCdQZe9oPntzq6jDV4vIR/Uxlgf8r8j
jTjRPgIL4OGqt7+DbqUEPS/pYSZjMz84J2xGHo6tk0NSvLh1oKfMrlTDbrozyP0gk4Rs9Fe6ysnw
HOT//PB4q6xB1Uydc2WvH1anB/qdL/WBrVubYg+R1JvxPaIFhwklb+7paI54O0Kr0UzFqyLJceup
tu+RynPCsPKiVHr1GjbP3h3YPx0WT2Xgr3cpIY29YphqMk284/c0cjVoXRdtht1yc3LL0isasKMH
F97AgjZsa8un49eBm66eLFsazgHpU08bKaoMRM9gtTKOyOU4XdPC4vrgo8F5MnnMvqp2jOw07XYU
D9QYwMq4DQQFKYIdhb3ol392qkrbNxtrq6UI7ztV0i9H7ku37UQ1cjij689nG69gaYHaSIyWHJlB
fafzGuoGzpHZwAVGukN5eMABEg+6XQ0CLX8dKwu+p7AwEv5CftmioP8SjqHMtpfjZhHocT7PYyE0
bXSZwzhX0e6BMOOSu7B1B5NUPT1EYHmG3Mut0UGw6GvSoomgwslAjHitAltVPivQ/qs2dV000Zlg
qWiQeAoSjN5xQtPJsk7WntFZIjJr+uhX5SjvX3MBYnwHq+NAEau/xHmd0inMSMOihuCAPMFQDNBx
HB7/0b+TDxe0kvFld6BIEOBdjJAmDPD0bQgTHsUJL8NF2AHYpeH4gxHYC/HPWf1rnx4eJG1gJVIC
zVb1bza3+fzJOPzsgcLGHCuQdDewjKeaPSEXOJwcFLqads23cVAyWZrw+XlLmTgPb6V/vWyPhWp3
LGXpPBm11jo6J3+m9R9hgukbTLA795L9NsrGZAf2K5e7Dg30UJ/Q63nKYgM7dJtrfQZJkBsPNb8G
dGAjhwGr6PCEKVyRogIdTRmYBPuudbJxlcu1y1lOpKANmbUMIIruJklyNgSznuaE0cLCvoAqpfGJ
IgaxIRB0AIZCvO5+uepwEytFe+6VDodOojFEuwRJDGdHcSsQzEx/HSPkgkkTVvL6sp8651PTUUJL
DR5TsbBxrJpjGrrnhwZU+wkgIzNfx3f1vgWCyyrqdsdBWTm7wFDRRgWoYTkbm5qlO3osFaBWfTMh
Y93Uur0bNjsl20V9GCL+8+QDKRbQF3uEpFmrkIyiKvIQGzDlVLxDwtDrl+cl/psQ2hDbqT6l3zRn
W1CTbTjlkpkQprOZU9Xlu1jzEryjWb5lA/BaIy3FO+rfG35ZOGPkhPySZEmHKMVv1Git86RbcVx2
kjLqsDVHYBn5Gk5jcjJi+hywqG+8v1HIBw+4YTK97sOvouU4pYIj7AyYIF4QrPd9k2aRt1Hu3XtQ
YFMeOHW7rW2KVL3ymovYnUZDU4lgrT0Mwa1+uK5BZ1QoqVtsjfzZEE1v0W4fVPoCgtE/UeJTp24T
zdljSl/kFywgiTmXyAOiP2ob46WRWKJFiMVfBQLgV4TZiOCR7zm3/ROJ3iJ2A7KQlJDSrEIA7ji3
cc2L0/VFgStNzBaB5i4tNWGawK11NCjk/KJQGfjuhwr0h7Cjklwgb6NPv4DoUmKfk0Z7VekYTzTT
evf8KVC60ht+TYijApDOUyjYUXNbFuW54sbMj8etQdESwlcdYOcugese9/aqD/pmwgp/guC6/pNN
8WWPzp2XfrmN4qtqU/S9BBkIFb1kOU9x8wki+SK/+n7QFBvfq1K7dDPUug7jxQEiTV2/6aAUdhge
VNsIMJVgFPnfqZrmLoTmBE7avK1sdODtXaPBZuo5NlfkiaFQMWilsf+aXqJvxf0JJIdLm/9srpvW
WVFFqiDv5/s/JI5FhNPc65UeKCEHBmL8/2OQJEqNp/YDFeIZ6+PHXtKnuDAQYdwzp06bGNSrC05L
IXUDmZD2h4M1aXkK3JCDuBMiRTbDNn01OunTb6SSUcBe9IcYf7RI2tB0kbCBfCqRp3l3TRS/+AA8
6GJtlIAyICO+7njGLYCiPvJPHqkYecoleJRP5Pnd0xk+ssxQHEQ64hQcqNXfRTCzDWBb2OxBrudm
UEBLaBvc0PT/jAO8Pw34cRdqMYQmY2aeg4VXupSHFmf4M9nOWTzZ+Mqt7ZwvAp1/6G9aWokTeYvG
I1WiCr4vJKSqiH31myuRF1Ek6lFBdtzDNbl5TDwLKRBr07FB5afwYPdDKkb/zfmksmRv1bqThHEM
9Lw0dG7PfEqAK7Rl/+kqsiHLewPB55hJtBMmBy/3kri+rdIiDwlxi8bCqwfWR0zZXTYbLy8FktPM
hqaDmXdbPXEi6yxdCednyA5SXcnU4cCFFFkkxApE6l2v0bwBJ84Qo/RYrUgQ0WY/vjdQL4vikQ2m
A2fW21IL8u7ItR1Tkwe93w55OHFQYvNMbC+/5XmwUOD76YcwP2bGFFSWDbjWq+jbAp5Fgu3nNlYz
T/+0xMXa/b2T4P11cXY84Wq/pBS2LTGjdeoyNi4q5gDmlV0De518Hs/baYqf15zDhyHG2LlPcFdl
QQ0nM17/zDP56R2LAcCjL4eli4gP78zGo0tksY88w0RGXX+0n3M31yVC1hLujI53UnsOndKOtzma
nsUla5lAez04CBvqgPyqI3QVzV0rj6aJHE62U2j9HE2iHpVTWuHynpMbnyDdQP4bkv2CYhHGyfOI
t8Y/2ZfqZd7P0PbkoGV3zwN5ATSx1TSNtlQPT+NORQ4DQhmDRK5N37QkFYJbF5oGnhW+i5Z5dDlk
pvyrQu5xkOnNioLhyOUN1g3X5qWXb64tS7n1vSlHOdFWuIUI7u+0hXb9K4MiUp4Li5E6aNLRjKON
GZaYH17wQI9wo8zo9ELl5b67VxsfqCmyjo9muGS7ormRUipCdQc56w2dF2sxdBqUDv6Y7heA22mI
UOumomI/shcE99HREk+zzHAdG/z762YJlP7MDhRX5fSJfNDAmbpKa90iWJJvMxCN3qDEWGKKa+N6
zuAvB1gZRSW8EAfHjGakbSysiSHfJc0ODtuiNaROjEEcPLvgNP7NYX2kJY5zm/VAETLjxvVh1h8m
si9zfd32BBvP0bAE23MSk4TT7Eovd32kty5uI1Fypiou+Sm3dYGpEVzisb/VibjKxIJjn1tiPH6T
vNgum+WMHsXcHDSkLBZYL0HctQBzroEqg9UAe9//SE4lMJHLsFHBhMkAu2daCevHYt9ECBtvMH52
axnO7YSuddKMBccqplT1z5QOQphdBHJRKDkE9y1XGaIfxVQmVkgTWhVozO7dGQua5uyG7WaeS4sq
EjClNH4Su2vCLUD+aHCXHsFJ6Gek+GvxhoKVY5wS/3xEZ52Am/DaYryYVBP9eZ9jhJ4TeLi56PmE
JJHoU0dmUN88/adMPvvzvg3kioydwBrpan+Un+9V2PQL/GNSnEbTAVvAF4hywB1hblvOET9yooFV
Zg71aywB5JWUrnoqqcREsMSQCgJ5NnWTSGhKgnAz+QlGj/J7yyfpObk2OwcIywQXr6/ATqQNdvXl
Tc6OzDcPw9oagOVuHHhsnZSRybJRiYlXDQhmOPDOXLcqEIZM4rd9lcFJ9AnciS4fTmd0cOz3FTBH
2BruXozjx7/2T/CjCv9q7y6s2b2jUMpbtyBhp+1Pz2QGFqoGbk7vwIiIhSVRvXgh473pPr3n5NUj
3eBTvEVBSvm1uD6/X7tOtQ6h8EXkUIg1tWpel+xImfIlYFFEKeGe+rXn6jSJirEkxzQx9xPpeNbR
BuPAjdV5yIj5PE7lNn9dyDhKyKGYL1wutWFo4LSoS8T4QAWUTLyelHTAdPiTuYHQ7QjRDhf8ZfRz
J/MeVQVxTCRwtsxEtjUYQWU31X/86K0DqmEUJKm6tA/qA9EHyTT205/JlxjlP2n/GEQ332pOzVnC
/Ivp+sxn+9bAzvJgAjNz21njlA2zF+5+o1d2udA2ZDiLSJd9AjPICiUJCuXXPqizYAdrpMV9O4SZ
8Akt9LKHis3H9HffisWUWTAbpctyoawPKW7HzZ2SWzpzVY0jsklAp+jg6nheS5wMK4u5FjTBf9Cr
fbYBJsaOB8I/auPYMxbp+pdflA+Cj8QvbRs0ovO6ZndK3syTjU+J9jtuaQC8gN0932WpCkwXPsdr
6z7pyBpRhzTkoM/rc868xXfTWv37p+6NOHVvFLBtzn/EWSCjTcZ2DXgG6dUGa0CL3d3rc5gA+0iC
VjVVeZ5SmNDRibIiCrEXwPgSP85ryu2f/h83I9r6hhMN7wkHfYbzTwaBhGHIEAACj+ZJXRPFTavL
R9zaxoAOXO9Hefv7arn+FyaMG6uVBCdkaBZMeqFXb41MNr5iWxD74RPtFtMEx7RgDlonnDgBUvpX
KFWmBrRziFbNs6C86rScWwjlvpznMlRQ3zAQGCywoQfz28Z+mfnYkVJ8cyOmc3RkyQnxbxwagh0A
6e1gQjAaFJPS8yBsyg+fw61JPElDRy8DDdLtoVaAFO80J8LHTNIg3yJYw6mQtSxknHsZcKyeFiX2
UMRg8EuNA3CdXJuAp/kFlhD7mJAE5PCIHMJvm2rzXNsTBZYmgsSufNTv/vByH0PGzr+RbAJIOFoQ
Bn+HvcFSuVKCIT/0z1/2rqr/rvYq22Fy7zXLxFGiqDjMpvsNAmuoKYr/NlpsW1QuAbplWxWuaAW+
uiUM70tj+NBqWrLM9rOCh5z/csXwPGOx0JYsrwF+U5oR5bPFi16mskRnNtynbPlQrogEUw4uV8gj
3KoDhd1HrP6AkW3pxV0JCsxJKNHmdaxQuRmq0ErMxxMQQbhj5sXTVXx+Uxw4yvj+dYytVdCj08X9
WReKmfDrEYWUnzC+jy2ZJJg7VNpYw5LlENNqX80NULu2c2/06+imZUGGxvHy7+344E3bsYEvbsIB
HkGjaw0VzkRGVAwZNDSMflTHt8rci9q5KMo83KhkYdHHHSngoVx5a4iZb7bdlztBvry51OoLTf3N
gN8FFJT/FbJNMHhYMUs032PbLp4Rb7bUe+Qj6L9Ftfcm7BlFpqfkQzSfrTU2VbQtfbd2PwLNeJss
VvmIC94qsCBHhpUMatugrRFTrawOHcbAKQ6OYzP+lW2kUoW+VXxm2AjW8Mq+0eIMqv4XEPIWqSZO
j1LBCulmtBsFyNu57MDQRfBnhC8s/ZRuRSVaA2cuXm6GMK/m1hjDHrPacLEsrImcaqPtKqkTIxxB
pv/7l4bZcs6zvQbpdwG/uTOJ2i10iSyGHRLnPt3rz1r3zOsVQxLQJoux0zZ7hwizo6sZnEvS4EBL
8f6psp0CpIhXr2/OAvAWEnqVqWbmTsjF2UWf+k8dj/HCpStdrBoZFwwebYlGMkYNtoQVmPcW3qA3
TyoDOyjeou0v06PkVy/CcrA7JSBqr82pBpNBMkdrIcTMOIi1o0ig1lKs2JcHliFPEGeYwRx76LCY
9zUfJPYpGedRLuXLlcOoFLGzhr0i+srTfqzKU3uezKnyneQ05SjhpH1nlD3CLGZDgjbg/rqQ1Nnt
rSoq3zWbT65IRw0ZUIr21CxRW/4yrRsiSg4QbwlRLOB/RWMk73ViPg4X46L324KWCjurMuG9cNAW
cF0gFSTwV8tbAlxuYVjMIqdxDrf96umxuQGm21XanKOrtgE0wbHrDqvn1JymOpa/DPQeOtfcWo2A
eT3THbwsZZo5qzjJt2iRZtXT8O0wjBpMgKhoPQkVECmrZUV8qKgpbOm5SKLCwYDyN34er+h2Hmub
74CYgHW1pCU+sJx3J47yfNb6UUoM4diPkKK4qkursLwPxxPkH6aTb/gqRQ5stWYcroi3SHj66467
LfJ2Jkqkvgls6XWkRoJfdR9uo7qwk10FklhgwxPG5ISChoGePtXCpBYclo1fWKZNgbY3By2aLAbT
EoFPshanVn7jo/1FX5YoOk4B7wW72lc4ToklOsgauHWZWC97mEPSFS7y9rHM8PDvplusK7yK+ais
BO70Pg/kWAPGIxz3w+31QIjMIGJGwInX6L2IKUdoK1+KjRFRZLIuuLBblqByudWL8Z5mPesk9wnt
0w5ovRewjfXb6/LR2GEj6fsWRck5C8w6erCWNjbcxvES+0vdqqs+YdGmtiHz7jC87uSAI0zldP4T
T1n7IacKi0ZT9GmwF3puYuJWnWgumuPzXP8DKeXJTajUSNKFsKdgW3SfQ38la2vcbLmK9Oqf1mbR
fyl5ZjeWViCjFeUbrRMet/Oa0ZTy8ZYbprPSOqgbfSCFJ6B1vaDe15l0UzmtqgoAQ/o6nCDUjeow
QBXD6KwvKfphR7l2fK53+71vCd9b/0ouwb1Fva26r2V2IU1sKqvSVGpmuPxUieIPO3AO7ajQH6RP
m5dUzoqXB6ld1Vnr/92dgfmbpO/EDBXu3kep97wdFr6PYGN4WgFFFMfXmL3x0XFXJHGwcqso8/+c
oZ29cEye7y34RVkf91ntUnwz2mn7c10pdq7yqnfCkR+0zarukozY8Lcoo0BEpsGzbgjKTTI091Am
fPqu4JBUJI7d+Ik/ueJm26ayMTrPXpzf7ZX0y/ux3V/xTJ8n0C9PV8Z1f5XZ94aDpIhiwKmjovgy
LdSvwpXPD3GrBdvYHB820pP9YZrMsyNF6cs5H7x2zud80O8g1XhsIjBqf4cI5KpjRyVJ/wlOPbqN
f/vw5Y6Et6Rr8QnrlMaqZRaG8zB8XyOOgzTPNV0SH/2IFqcRWtCq9tC+U2nPSmMywBrQftv4Czzj
ty+5GGdrOMQW9DBeVsO9Ss97Cy6wiJzEFmHkEHOpLeYArCMams7B4NnxN26JbZXfbzKN3HKKdj0L
88cakP3fpHHKV4tUjrHPtvtUrD8BNH4xADwPJdYaJ3mBkB++frNNxZR9PiqO/jIcCd8ZM4J7jAuD
5bCy94yNPM3ApY02VY8/u1bWfkamGjnsLptDgB0+5sX+Ke73VhjCe13fRkWM0rtad/ctzfTsZa2V
ybuu/lSGUv5qHVkz85uGhnMutGWc6QjLN5DA8Zs7sQ1mhrcy6h6doWrkis/Ml5hmYBxAMg2JG/cM
xKD0uSKd4Xet22nw63G0dWX7boOmpBBsMm3ohYoZc3ZO22SMWLMb1nnkUVE+KdjwD4bol77dbEZC
p7AABp6xmJkDA5igFfdODblGE9kfBrgR+1Cr4IcluSbbkJbvzCSzibpTSjInfLylNuWtzhTmT6gQ
lCSYRRcMq4ufRNY8T69p+Kx15uh/bpeF2DG0lYoHx566XGkB3eAxjQf8ws9SCsZUu9aiyBx2tib9
3RX7OzBOUhEUztFq7W0l7OdIf4RaC+HjF7TOoOjLP25+CkLEhPfoTRjf692fXenAfWDkFjj9H7aB
x8krXg3cbNu/sL1hz3E3rfrsrJTI3+DrpSMioaiarkrCqGMWA1L3u7ytFkXRWfDwUenxgO6rOU/T
VRPc78yhrifXxGFi3XbokgqthxSZwbCD5HHFKdHSemkhqg9WwhiSkjUmx7gjBwjhcMGno+lEX1NE
ETBmgLo56lWzDwMDlSfjtzQuJmzerqA8bclgVn+ATgq4C3S/UnAGRoenpYzivjaX2EKOYUinuydi
sgaWRrADDDy4yYZiJVoh5gOzD3tHSatE8vPRRPn1B1uJOL7vqd5gSdLomqPrXq38xR1JhbIRNaBL
d6erchOw4ScKI0/6Diy00CRYsZlhoWLkyZeNIs6XVrKyfHSx8kEaeDOuz+2JfiOGMaVzLIP7DE42
Miq3r8q5Igpn8GxLZ4TSYyy7G3R8AdFJNzSV4NVtyRS1X3ILmyUskAQVjd6Zqo97oZFQq3208q8x
FXm7xrcg/8++jsPoVbtdIRV8ocJnna2eJla9eAcoOnBEr4sE2kMhV8s8Eb6/0heC6sL0wtPShy1X
PjVKvGH4Dy0jLrv4qlI23b0jPfkPhl5kQcuBPOG3LnFcuC3Qa2J5soSTDv7TRLH5hdwFWU+lzcFU
seL3NgcKrF046AlCSXjDH8ncq5s0KNQPKZg+OloqG5bVFhELLraWMes/5YWEUCw8tGjhwfldhdDf
8G5a/odMp+WUtznrwe59KSKAHJ8Fq4H1LYGEL6SciuTaZ6oIhY2ZE2T7rIR02qqQyVBIGew8PO84
nPLsm4IGYA212nm0ljycsl1q1JBQw73mv9Ck7ivyqC+6ncWSk7cizzeZjOx2JQAWvLdfmioUKFdQ
MF1qy2NcncoX2yRlEMNyZQuNtPW/6QQXRF/H00RkbkF9OwOtk0zTvGZ0/YXjhXqigSag++wITP7F
2QoJk4EowEl0aFaBsvYSrocSrUt2wizJLZ60SuFudRF6sqlVUzmrhk77HBvrJJ+ZNYDQKITGC6MP
g92Mj4IGxm5C6gWsxPX+aah07lF2f49NdbVCqCgFJiMEw6lOnbmdqrwnGwrb4rvddoA357+rku3x
63nXkr2f6f+AmF2I7aYRWzFsUo+rqg5Er5OUB4ssvqtYcxLZysYtMD1vluYmnCZIPZo4IIbwG5Pg
2aPwiPt50qSX3bExyB7V8lYR3F5113rywclvEiQZIGqXrJ+wsMR3JlulzY7jC1Ub17FlKZUsQazC
RdnJDZB/EzF4/tsroPJ6QMCrLEPqFAoDti1CLdF7j+bL+72z2J9ouzMLFF7OzHdXOfWZ6Wcgv8+v
zexAU+RwZK1eHVjxtGPNAntSLQr1WtqegMTLrQWybAKuJDD3TezxZRbj5Q+ejrzHMzEo6Eo+VqwR
TGzwgQv6/KMiPv5ijlaWpZWyOgmAOzTLjA0xLwARWTQja0QhSrOYxkb5OsJzh/pKjTIIB5xeX4ZQ
mPCEftoDwiLhJiQ+7Kcv/1vS1dBeV2dxmbK/cQbzgPQZQYoJQqIBQCACfxGAISMFGP5aUA6bVngB
oS336FJJcs9xIh54UryTn2kI3kOw4qaXP6qHlcMpy080d6Bkxq++1/Umn7iWvV1w5tu7eVfk1jbZ
+3xHSEea0FSOYXyzMkOL+ugc3y+yGV5cy6KAYxOZe6Q+rF1dH3GhxjSYfNmEwH6GFlGh63idimyQ
QpajLOG7n80B/uICSCwBZMAvhKrt3TgkEKMrFSLLRwJlrFHGsiHfSYOJPm6QVMJPnbNLwbDSfcLk
1RT4jR4od92MjtpuQvNM1wdB0yJ266SMFjro33TT9pVl48PXgWqvm/sy4cEhDPuQy2OkPB91ztVT
7ft4QrQzhGfVeTKM8EJBRlwhhBvBa/lrSLu0504v/3UBbdu4IArSNSajaJhvj+5jLP2MIfi1xTbs
zy/S9OBUTGhonFr28FPc+p/yerz48dpStKHVGr/qadmMgLtOXYo79ny25/GiO7QK9MficV3L6d5z
4ripOgL/w/BWvxxxJbzdc1co9LJGxLVRFPebrwQ7YegAp9to6JjeDbkJ/PFuXVIo6MXnYreSEKU3
nDRnPbNbgW1YLGc2i2uEuvCsAjQ9T1B6eDXWoZ7gZwtKmZjfB/1V1cq12UaXI4eV2T0rs5Wt1By2
Ox15B+Pgq9Cad6TKoPw/81Z/x7Cjq3/wD8UxKVx/bpr81MmUinWMW6qHczdjnrbc7afr6CV8LVXo
FebdPXBbRDhblbMQpx3ls0c2YBM+6UVx4qwAI8ejXo9leZSNI7QvMYZ3L8AeX3SHvpsFKSEc9v/x
w622HwGcddkmVHrN/Zm4isZBHfClj9oTOfJxQMgoHz5GWCKd3C20RtJLasrKNKflknStFaBte28B
j/6qvaofpGVBfiHqupkb3P/8iWIIiqe1toRZqpk7rU7cBqWvqKS4I9j0i7QQYXxf27oxo1miFKbf
jxG+Crf2oK8AQD0AOv7ijDfdlMgPx7zws8mWrlk+WylXy9ypgJ1q+KH7CxgTIXvRWdKHWdP1Cfb5
/iSg7VFAJtEECYl2OuJvQOIx4wrCmz03t/WvtaWy96KPaceL1VOtBAEFijfzQcZ3WG6zFbN0Ygzb
MsQG65a41NkIwoqN5Xre/btW4oTs8ycgBm4UDjfCrPC7oXc8S4IiqIQIOs/K2LManpyLng0p1rk6
2OAwDgOm25nz7Yy46BVDjSxfbFXWeWXgGqflFpDSmOzqbR+3a7KYTL+MhACTy7wwOBEJCynO6fur
CAfxhfUBwSSMu58M+S/QVPmjqYZRdstW1D+a3OD+ZcUUeBNu19qLcJ6iKUBDlhthgk4o9lFlEeVn
aSBrDJ83NpDmGRngVwGlUxSD7Uf3gHu3/40jJmu9NJQyPp5w91mow+ZQ1YHIQh+HcmtViMqICAgF
caPNgs5CX9bf3t8iMygVvh0YnrSVjm5OX9qLfmDcHrnh5f6Ssj9hYoxpaEvG9RzBGNdEc6Y/YjIU
WtH7CkngvXROak1PdDvQrMKOleX80Q4k942jFhfBzVPwDdXcagX6Ro5tP23Csj5dLDCVaASK11Qx
SlxdLApaKhkFq6UsdhEzzk8Khi9MaNY+8mAUEmH0kcLq2eIbcCJ3gnd65NTq2K482cQUIB1PqTCW
LnkEQHufTp9gz/KbnZKFYTeqAR7QZIRhsXQT9ItPLcbT2qWcRl22mW4xaOMblWrEplogKAtt1M70
ohKHE76uGEujI+88pzcc4npYq4EdgUq8Ut9God5DG9kHHiQLKValK3hzb96OCLonvZosP45YqNgS
RpZVWDykbdvG8otMJu5prtG0Gg0Ox1M0YNWiUbi+U6GZNq4lbqLRrM3M8RdaqsPBR6b9tvXP+538
J5cFRLCnWIh9XNW3Rc9lMTrb8wOCKDrf84uo8TqjMcEWqhX+FpBxdrNaoUWx702bfj/kTAWYHWIh
/q0hTEm+yzrMJfRa6lSBMGoRUeShY3SJtKmYfHvLLlLfIe64z/Bmgn9WYa/E9ztBxaVaL7w+CRln
Y+Qkzp0kcr/YYpkFAbyZCs633wAtAZfZz2K/jVGMdgElE0tWTwoRLwl3BeQIxy9RpRLdvzB1hE+s
IfIxMbaWzSZkjECbqB6EVzyjMPpW+i+UOHytD0dyzhioUIcSGvTpPhvzv7NU7nWR9jvKicnNS2bO
Cq6V4l3GIxSLNq3kEH33NU2DCbISklwcWaWl4GfZIMB1OcrCVqnJDD+hy0h+Y2LxRnIx7ilLQk2X
cuD//9TWCVyJjaQkKj/GI2PWhQFd+nbpyBrOyDeO1UUslRNLgbvhmwiLi22XadQlvxv9877yBYuJ
Yw6/qWMubInH9b+roYvxEVFnGOFNHYzMeIqkYWohVKLrLxVoQL5Zut+xBSh3auuP4aEE8mDTcg/k
52IyOFp5ZYphN88qDxPaSzfIJ1Y1Fp6+x1xLBSEMmXFsV/QGdawmKj9FOmhFVxTnjkOF9sIIWjsy
U7iItEFbQtUmpra6ojsMzlI6+M0gR1TKPfBNENe+03mRE6I4/WQQldcuDlCJD8wQUjCBMKCn5FM2
yWi9TCHsVCPqKoXGOEhb3wIyZMYpWQ9XxhRlPn+342juPAqf1CMJczmLUBTzcHEDV4RuS1TEDxdx
1+GBc8sWur6wOsiMLnLPQptEkMQ/2q/W6eFjetZZ9JRgDoly5XpTBu1NlXUT+9eLHv68eMo70T1/
PUMsZBeJZgc+U6Igququ29p8N1EuYGZ1o01BZCjLggEej8FhiW0J427o3aHucqw7OmmgoZAm9qbk
q3Zq2c8InjYaPE/40aYoSMvxQK/jWtlwgZnX8wPcd4UZnWzZuBAyjcfxBhpqjPqGgOu72PyC+Wwb
nU1/rzCl1MyrmEIzHkZspkHVvhRyGaoKi/Nh/oU2d9OSoKqwJqo9r5avP7Dqg1aB2XaT1a655Fel
qW8696EzovS1NpsgxmhgnarMaWsdUL1jcuvWbebYh54eZdi4NUiXNwIKXrc1b83RiebwtietYoS4
Tr5jLpbqSFhrUHt5VFSySPVn9BSmsbsEBi6eONkzdgEBWhl9cdThWVXEpSrHOEaV9R2FyC2MJVNq
z1+FGVqfacKtxsRvaLwGVjHaQmH6umW7G2fCHVlLocIdbgpOKVKGwRPM7TlAUskCEceZEiLkF1+F
2hChWJd0ax05igGecWVmuAng/IHfII7gN97OiZ3/tyJ+LTpmBcG67sI0delwREv6jhtI6mgpT5kL
oPcpO4c2BNftXqDLWeGTlhkbED7RQXn3qh+mAgY5LQIVpCEVbIAcucidqYdsFET0Gngo3KnyLx+v
laqo3fAg0nn+3AAVjpimI/n4dYjDDkY3VxXRcRmDVCuIoyGBFBx1mnzirxMVvO/ICXhcUbLXm0Fl
1LMiu97RRreeBGKwjfM0zhxFnTrcV0aM2K8yZ2R9CSmFiaJ4NDqi2aj7E43NrBafE9Zj5PqeeMuP
twQQ5xCbM1X8LBfyA9rCuwcljzweeTm4ass4MYinqv5+RagzmOMlmQ8CZYQxPYPr5UsjCB6ey25m
XZRvSnCo4sMs8JYIQgBhQPXl5SINrrd+DYFPgQ7tnkTQMp1Q9BYgi0u0MUnVFnSdHJGGIIFBEqlf
aXbxcr5M5zDEntX42DjP4AV+NUHAvgTP+wFkqEQzRHbaB2hdnvVvCwUMl33fHlXVs6BQcxIDP2ms
bZDpKTkdQFoS6ypBSdBWxh8Y4WNK9BccgKIq1UOaW/P7xWmlclvpErf6pQmMXwRRdO9I2stIgL5i
4/1EX3qJ6nxTBKDlBf4eZfBGr+RaOgxCEZNbG8MThJklvYvrBmoQpySRjAvxervpZQOANMa8sL7y
/SzdmSuUpz6sl7z/wkkyrmI9zcGYIbzw5Z+/ehTeRLjJ8B9eH3gOb1s07VmCK6b6K4hPcFT5Esrc
gJleBnFUbK83O4vTaGZ+zmpQlnIzIZxoNOAeTv5Hw6bzjbLSGs++iOCQOBUiNqpxdwPQdZJdopm6
YeO15NwWMX32adMEpaxDydscDag7ZLYz1XLZA16/f9dwS1WvPlhQ7iMeckTO4FptFbWdV0KWE4I1
LWFZCJXXxqbCDSio7kmvxOFgBwc/sKDbG8ojvr4oKqoCVGAYewYqIleAWM4MXGx8wCIhVcOKlx8a
aokhsvLdMfjrRVoFREow7pYL6OX3kmpq1+fGOmhmwFM5UooPKDNtBeRkLnYZ27hvb4ZkTowFcWea
1HbehIgIQvYAq+IEniZX+E+fDwEbzLS1l9ZlobwQC9RB9aD6cjboE9+qihvG/V5d6XIfmZPrR6sj
YhPg71RqZZZh9dMCyOhQm6iwXZqDkfkEmalwxftcbEIx3c+a3mwfhRBMX7HB32AgLRCsjtTtQZ7w
uwevTLFEqjSA2SSAufemBMWpZ2/5cx6MJT7noaocY7XavDZ8nVps2KWszljEbKhqY3Oi8eeigcau
SH6qNlguVKfEEgHfyWN5rH1+HO6n8vJG1mQYoSjSFlL6UWORyac8ZqtqvZBafnTER3B3RQm1gjVw
eOgk/5KSdV7uo1r0U8WpUxs74lALG6Dux7yd8OycNJZ4gcNbSXd/2xsvWZIxMUR0EqDgONiAt2or
uXEe203oTfrlGB3p+0ZHpdDHUnHOldcPBivt8cMR2rPGGUsWYlz8JKThz67u/lQcwULfg+w42yH1
BHrWXaeP9Ah1lL1AYGOOJUzTEERF3aw6sPwTWidbW0GETtBxJcLwBGFMv7yBUtaD8JXLWyuVzXBp
S5aOJ808g+wuiBoVjgTEi/f4GP5ctkdxXjpQc85wCdgvFiARj0nWt+BsE9wwKoSGz8XYCQl5xyql
GHUYpoEK9cwc/s6TYdugXssNA3dTQtke+l6juWEbfgRwgYT16z/TKAW2MumPmd2TH1CBOS1KjvOZ
mU95UGrbQD6ErCKD+iZYfG3gBfsQGlbyUsbZEv2BZd/jvmQJOORNtpofGbnNol0fqIOSmO283DaD
Fu39PMjoH1YnKJCwMcZN0sBZQ2QSWOrVxU+AdfDHSuJBjb/lWjcDqPuXC5VGXWzMFEizKUm8bf0A
cbwv3w3OZMrN+H1lVVDsCGyYoMO4oVsvLN0zYWmFZgiImW0GOZf9nPmgoeQRabgQqF72/9HQ/t7u
YBRJ7uuF5wAWZqtP3KDHa7gXNp+0N+OiBswuIHq7/leNFXyl9hfp14X/zxFWUK8VYWD37fLhZpnc
LJMUwiWjUAwL5WsrsvhVlGawz0OcHiyOYHtpA6xz9ubIww8eP1InJLR7xus66jZHe1rDE7rG8iEb
v6Sw/mjmu47AUphZM4C29f36U+HNknpHee4JgMkoJqKHLNvZGG/zANA9UbxuvHhMk2116Rumv1li
MTp1CHbkhhBYX0f1g0oKP9WmFkr0dIh/72L4oI6aaEsSumQQIuLSbzoMstO22L6ttF9ffRIjn42H
vAtqxXY+vHv5k4J9ZyKwKGjaz8I1DgRen3Hf3EDKpF06GVzVtZBPig7/qB+rz2rkfjKcv3gbt/J0
Any9JekOgL3nATNrn8l11qDykWPBZpWYI0BVcvsIQS0V+ybAbBGg80y+LwsEgrfwfpR3+5uurIiM
xHUOj/rWuSMSN9qOqFbH5UyonJr9qepPstwWyzXoZKkhHzg0BjbIfddydLar2LrjjaZhpc1NwhJV
2vrOb+lSFFweZnlehsynuzAcjeMSQ3f4bEUTl3XX+THzx3J5Yzy/jvltjpNONZvb5J3U50e8r4rW
Rk2qaKKcn3jDnkgi/wXaNJqo3SF5MWs5QzLoCIqxInb85FxxNGRIk9CG+Czm5Bkl68wSybbWXlxV
c4SIVFerSk5RXRy7PkrocJyFvmEa3AaS8GNpSdX4ieHDTno1c7H+PcLFGpt9x3TraYanLLEV2B2x
zlsx5m7vXeaXK3ESi5EBIfRQkbXrL9Xjv5CdYOv/7G489idg98tOGfChO7lGuXX9f8i/woDYe0V1
vh6SDSxeNcOJKeVCaaGjXqQrboQxX8tDgcv2tCazomhSRJ9/UHZceVc53UpfwjyDqatSRBl1Jz6q
s1ccyj3L/IlCBfVQBkscTZh09WS4tj1dieAKwfcbA069b9Ua3+e5U2b4idoOLC3Dj9HJ4RaT8XW2
F6UvAf9iFBmdZGVwgU9kAzdMtULgcPbNPw7qzEkGj1hAnpxAcVULm7QTba9omtffvVP8NHNpT917
Jr9LO4xlXVMCAHYYFnxwgvPhBR2KkLXFF0cK4VBTigu2l0QU/lsSZqSEIzE27Qq3PBwH97JIWK6w
Ny+2NCFPBAb66qfr9YUItDzbnf0kaMKbya/W7L5LZuZhOJjlvAbdLTkY7vz+VCVq1zMT0cW9sxuv
svxp6Pn3jyQ+fGSm0xzlSvPbauXFJ/wkDYnTyVZlM9rYu8q4oYT4gbHMy0jX36lVytSOwqYW3C6C
z09gpIB3LYCbD/GFmxsQH9VhOcTYFPaj3LdUI8Z2REqRpfTkfuWzQ9MK41PCL8glxrQpo0YlbRhV
e/QT6VlF0VXmcLciNsblgMlhEVbGbX5VfANaCaT0kQkKGqtXcOqinhUm9M/GFozg4ciw3N7yoAnL
sT0Z+uob5pmoGKHFrqkC84oqf2QGw2GC6yQnKNZ9/AsozXZbdjKhlzt6iHyG3ZN35IFwZyp8Kem9
3NSBO53vKbfV7OgqEnaLMYn8YV5dz23M3c/xO8TWuu6Iy1Y+rXOZB4cBgAf4WST5j+H45Rnk4hjh
vIFqVeJ3u3M07rs897uxvLQs0V6prenwbHGVhOUiKb85KDQT6mGDv8jQ4VjjEO5LnFQwegKURz8T
EWbgVx3448GUGfrYAMKp69XXkOoxhEYlNIQto742MyR5NWqDhdtWtAa43DlJKidNz3FBMFHe9bc8
WZ8whSc7JmqkPTkqtnng7nMo1yHzVtkETwumFSEp42q1pujaFWgwv4QQI3nOlBlPPt2/vsc5Q7jT
xeQujTphtVjtWbzv/YDGHQ/4atakvTBOuPydjP4vQkblHpg0skPIyrnfWiZcN5hMCNMHhn3nIK13
AeufeSSzPc+FouZfr+SrQWlYlDPBZ++rarico4+zqYWEkPd7hCHUlFiVYNFgPBD4bKejv/GIiSpT
OOmDilYFz9RpPL0VXPillIJphMzQXLzpxbnmPCOJau7YYZ7Z8lcYdTbvpueRCv5+Bb87kF7U2EBn
HLsTIiZD6fp84G7BpmY0QDGJp3PvryrUPFxBMCsjuQVZWKrkjdRlyJN2gPbLm9syLwb8pkwqAypU
WEXPHP06ACXOumB91CeKn7vTG4q87IojWAGi9/gCQy0drwR2lCXnGtWsw2xmtsfUCGvFT2z3sgMw
EMaKN17xtrUcyhICmdkyl0gyMxZb3WQAR38PVs1sNVP1mKlSB7fgLpDa/0JC/pug09+ZG8ei0SXo
8hiGD5C9Q/MwCVJfKsXE+yjLM6TEGVhkNfqusYbTfRLHS7FK40FznnLbsTLi09gDyIqqCM1VHsxF
sTODyzin9dtvEcK05TpVasxeiLnvjfmPeawT+tsuerJj0Cf2rxXYuRS2nxwzy1wkrf7XahIGbPQ8
lbAeD5smp47KLv/bmVzDgaXrZstPvlyGBtR2GySfXxvp0XgjCqs5Qv/IsOYBzsX74cYG+z8FiCx0
h9a9rYp3x5/Z2XfpJ24kKkGOQ6X8adEU4h/YznMX1Ik69vok8a3IqOenjrXvrjyNyPOYzArQ8zAK
kuJorJ0I/cRtU4GWKRchT4yxkzGm2pds2kK3lQMBPyJSW1VOGCNHY/7B2HxoDyY4/J9sKUp8t2/y
PhtXRBzLbY8oKd4vqpF5hh94C0s/d7pC9ltwbYUodRYbxXCs1tqneWbOgMAJtP3BqXQj6Kk6Eqpu
DkSoyoeLaNp5pUGd8OBgrI7n8voO6Ap2m79eQI+I9XROWHDoYO45h72E8TKpE8gZDoqkxf2ks7yR
pckwOQZwdsawES3oqZPlEcw97D5BYzneyNoEOUjxsLIibisIH82eWgSX8bsG2WMtaW38nfvx/hDW
ZHUdFZ6NWLnQw3Msq+c5ZpcgHcv23eXwm9ZSR+7ob1xQ1cqb/kWFLmDtVt8blf7CZ9mWMrIHHwIR
v+tA6DHkzZses28MlFJStUrvlqDtSX0cM3YllbIO7SHfJGn/sjLapdUXRpABZ3Ph4OM3z3XEXUUc
Cd9jt/l4MN0nZo3HAisipXpXGngA0SISp4RCS2btMpLl0Zkk8r8AU081ErXWjUbX4mO6WG6qmIiv
cACGLq+6A4OqOhNdVEtsGV6qEwvZh5Vt/0Y7XLtcJdXLXqmQLs+Iz7Th7SyuVB5VxP8AJALAwlTk
UAbxPe4WlwGj2WDhebCrDsJuWIdb9hrR1Kro8nQQy+whfuTvZ8CyUMKkoEej6Bar7y//jhCmu8G8
Dr7loUgcTzAp6d5HB9V2MLNtTZhwfngZISjihuEnfrfCNxiua22VRTzFalFMYk4o0jKI3RInIfYO
EQp20sCOu2jFiNQqez5bqyoVRmLiaIzor9D3ONL9+y2R7vzBjecwVZ29XxSEjjID1zPcY46UWooZ
38uh19RwTpfsbbSyfb8bMw81GNElWRPe0r2Y51DynkFRlhWu0mzvo+dgSqYEN1JfpP+KTzLcXDO5
M9fBR3pC1+Fe7glpJ3kDG6LJbKdb5sngT+dVcR7NbMsifOLYv6urkxHzlg0haTv8aYlYLvtGZRi1
rrZiaY+5idGRkBwLhmwSlAiiImteP5XdaEOAj6QHmzMK76PhUxAZbWfhRQWxnk4nPHTqIDUVSSmN
Gay1tHKJR+/yITVbTQDSXpiOPf9aYW0yjGdvWebRaUVlUADIwg5TX4t0Xv7YlCwDAU5T65SHwcWL
R5b5Vmkf4+/hMaaTX/HTJ6FHTdAsaZB1aooqt5O2h0wfg6DADcs4pIL1W5kLmENEJMndDmARJ3Di
2wOKvJyITYFfsqj1AmC+MioejWM/ufOsEjDKElf3HwPtUXFjllW5uddZcRHDxqNw7hznm6wI769E
J5zwb05nGNCn9T034Xr68Xd0S9INKa+5BpJbyYQmTrKMaBY4S9PSoqwRxg0TnzAR+XU9Wj/1Fxhc
1RxQiNcuz1gwjih97rZITYLwL2REQQT0Dff5Y8VhpOHvuvMoVYz8xAGzaYhCvfTWfuqOqabiSzqS
0rO5O+tVldgzcqOomJfGHgZGqAYyPxqPchQBIvltMdeJWgHeI8R61+l2zZ3pr02CFnaSb7IdZAvJ
ZYaJuwg9Dtft3TEpp9d2uJPj+OmFKIB6XU910LJu54YHN2sdLqMyxVgAcMOO9CiDgbj1n2EyYWV2
F7K8Yp8lde4JUDwCDvIOR1DjyqUXkmCxhUqNFcMITyoDvyDlssu6DQBSXxNKC5dLjBoIaksBECF0
YQVoeflRxn6MombpIz6o5m3is9oC4vRSUSV+vlZfxeTOvKUABiJTLqewSZcw3gVb+QfeVlcLfHEy
GoNVKvIyq7h34/x0yPMLdJnSI8L8Hvb++s9cWoQi+6vW3AIVkONdz1cH7qKTgtT/ureYUrAeFiVH
3DN+x7eqcQC1E1/A/g/ixnhLRoY0fFNjBi5HLlIPcS5hbVZBBCDG/2RFpqH8gtWrOeUzQyu7XjlM
y2mA7EN+jeAF08RzMf77TIqOsJLjcYqxqoTPRjz/+GNu5OtHfSurOQzN9CY6HiJTpnc/bwlMktGG
OLunF4RlV9VpHa1uZWRY3SQvp0BHDcoiKZHHzR2wRNu0Jy9f7NodX/Ae31JPxamAgpl2IlPd4ZFJ
8tLEuXdC2B9SH9XyA+1RnLlRjEtlnkIn38BF/GmH8eMs01L1mjkhLPI87lgd30aiutyGhh3SwMDw
m+0X0hOFsiccBRepeT4UGT1eEMMgbgco0BS0Qz5lRon5nX2zbHX28/L0RYxgNDu54cLLTmPONadO
UJDcGBTeBv9vR9nuwjZWeH2XWc1Nd+OW0zTPn9wRrXJER6fEbVakQtJAqCN+kj3OpItBn0tjLWjk
Q0BrlfJw4tsHS0WyY8cA1FhIuOm6o0s/7EkaRZf1lQkkTSx43jpAbzLQYfiwwxVmWTpXHbOU1b7O
Ac14YRNb5Oe+CpdAxyNaf7LbDGH0O7OuQ6S7z5D8fh4Q8Kq4KOg0u6TAT9IEZHPRVPNAQLOEbgUF
eVd7MXBGc5XMH5NbgzPedHCBCxEBMmRHQiiWbTe9BJ0qajDzczjxWAKKL0DdC+oPXOXYmZk277lu
DdCHuxjVL0or020ylDR3x5g4yQXYUL13V0HfKQHYvOQ60qm6OU/Zw6oJ1SQX7vyxVvk/VN0wXvkP
8AdHJ+WBeiHJsCHNbtAwPdu5IKRuXkBmqLuCf9YM0W3scFUMqPV2TV7ATrvsYfq9iXhEtYv1D06/
C+JKj+sTR1ygCEDcbtRrYu4uQu5SM1p4lVAOp65l3PAHdkyQc5r6+iDTr+DllsmaVZ7jLlaXcHLB
oZo5SNThmDtGdEVAhI0UaFNNouSggeWc9jmHlgZtKlkDjB+DBZTVOSQa9/8lW0V6JaiTkJ+26++W
Pv+UZxf0LM377BYpMo9VJ0elWcLvxnUydtoVrsgZfix0ZCGq5jraALGF4tIUs52o5sAfhbPd4OLI
AC7Mfeool4PEXgN84meWkgrrPUZYX/OrP+sGRDQf+RvlANP7+TjeruLqXIGgBSEHutoRlVttUr75
hnehybhwnX3d4RSa8NqnuFbsZ3AIlcf9i8T/ugien0Sw4Xa6qKbuS4LPrwOlAqDi49sQKVyI+XcV
LyTaPXc6wYaOsgCWQH0XR/BM0P8JmeT5mxAjXpjnahM0qMSbkZ+L2J3rWRMck2MVEaKgX4uD1rsq
sfEM1tUiJ4lw5KyOtgQTwN1ceTAyvwCLDsfU+ipR4Tb3ai4eOUTI0aQafKA36hBdVflL/8qZfJ1l
4ejUka4wmPTM2rx3fSiqjebD6ihSstlNCTvl6lh2PTmnFOYrdWwPSwLElpqOiVfbXOMlmWOP6Rgs
4BeMHj9iQm0iVfYLHXa1ZXYxeY2fN1InI7fBZuj02J7+x0XSQN4WeMS2Cug/wVHn0ZfEpNBJZS/+
GdierLFiFLuEPb+gaSs9/Kj0XiGnkcz9xv9lbkS0MzBsQCHNLBoCnappHNkCzyB2OnmITvDY6mGV
sDDN6fSILrgA88qz05chQKm0DDlPJcC5mP28Zn5fRwBGdCu7vXmr635SIAszv5B9bYn2YOByzS3z
dpPqQsrnsfPXaVs2h8PmrFpUeQbWej8NEiLf32gJw85Z18lKwvn4MBF7sq3ld0pV/Qevqlevgjj3
HJ832keho77LKLMNS5DUFSYfvHGYLUHDAztq5OO8HMADo/Zv/r8GGbJnCo8DDgEKR/uMJcehUxKa
mmf397kOq49JFsqOexLtMt7SvUzMKQHK+N2Bmb/JlndRNtxmJ2N6+NBs4V+6zwyHl40QF8UOykVz
qfh1v3I4MITQy6hjJfjg5T5Le1AiaGEpFXHm6UnrA2VQAO7YnxaSiRM/W7QGEHM+j+6pH2Q+RSu0
/9IcAipZv+I521OlDLmsC5E2MwkRi57uA+uaCZd8n+An4OG4eM3hdm3C8UL8Nqn7LAOwEQwSap1k
mS35zqdLxCNo+cECizw0jygDiYzYUhmu37iTraXodNfHTcL3gTfrgiC6iRiCnEaEUtuoPvOmt2k0
roJNwAnWDuXIQ+aoxwfonqgkbpElSwEnwvwDJXFFcl0XgIjNjOgwEkYpfxipYRkFjsXHSUEVZeBr
oTpxh7kuG1tCtbI80fN3R3TIVt6IRlrpk9CX9czwqUSIiMB0fZHG2L3a8/AtNne8qGHvIOKBMhy8
mg6PC6taZ9fLh/4QyIea3O6MCasfUk7xijg/fjsD8vsKfD/pgus49VV52GjBxhNOE7CJGAdpwspq
6REUl94cYchUR3WfkbPgS6v4SvvUnpT32yhZBuF8AD7nUPBeUbuL2nQgHe2EaUGtOyv5P/EKAgJV
sDV3jrXL4EojmjWhHDN8+Isy4so3uLmPig+DLnBMvq4oKYJAk1zhm5HWB/FD/l5Z99aUQ/3XPM36
EpRmrxHTGKNk8wXPOhZ4G5Bpa6WIOZMSgiEMiEsHLYFWb+BI2Qdeq1R71/H1hhBbL5QHpuh09h/K
SrBjkBgwJ0VDinzmxpxwDRSivkT3TR0uNTeAQkwoour8znymgNxjZxhdjYMcAnj3mV35CjaGK0+2
GbBfIF+SJX+IKu9enUBMPIA1YC5cT969aH9Wd8W5IWIo5R1OQcTH9XZLrYKWN/FWJllzkDXlhtjY
lq16oPr4CLEZKl1bpbCZ7Jr9PCy2ApJywqcBuDrTWy6JjVbJhme6cgpg4HiFlizpwLiP7coOvjsf
XdGBkvPqRbZYlYtDiNlBF2w/LpjCYyUz1xamPFhaGHCqskcW8wqnC/CXIDXi6apzzqccqGkV36XK
Mny5O0ku//diywv0H0LU9IjhOVWaZLuM+Nd6Ijsgl+NQDVI9zOmr9tLiXCtFjKeJmxfvL73B4emb
C5z0044b3e+2zVtkNbhjQBks8Hb+qr4OqJBVC4BlkhBwS4wumK8uHhj9QgCARV/BMWVNo5Bke98b
03G9wNqZo+FlP2/26tSx3U2v91q7o2rUMKKSk/kLUiATkfH8DixlMNpyXVt6XYkJBrB569+4PdJJ
feDH7sdZWhnOfeUiW21/OhTyAYgqIcOlBz4qQXevDpKMIjSiQihVCfFfaK0N7jhfdTNRaxsYKvhQ
k+raBkkHQq4jEDJHayEG6KaxgXe456Zx3M9Ba6N6RVRzUD1nadYG9LIi1Q+rl/PU51uiqz0Q3kHi
9s107sfE3Wge8/uvy7BdmwR46uhkwDD4X0p32iGbaE7Q2IPNqf3s6zmzpmGsdr4+QdIJ2HK7mWox
mcnI3TJRfQHMGaCWnfA0b1sfHu9CI74xf9tOF1zE6q2aOpH+hPl2Z1HVzrFr9HEE77BjPcolZ5WY
z2jnwIgc8kQm/XcaQ3jrjxYs/jD2S8OaoTBHzxIRcxJ5JMApnJbPDlKu20NJ58RSfAVJy5eHKKPU
o9nPhOjDSrjEe+ZjpVyOjPArUnFalSOPsor7xrlTelf3qMYxEVpit4/And5E1ZIMbhtuHPjc+/vN
1zUhiIHhZ2tEn15F6b9205DcIEJjXbW1ugk4d1J0Y6ZPKly2Zr+aJH1BfmxGUvvCDV6HmGJmSl8x
6leS3afo3r3Oz14wc/PdvtFTqqvESKHA80Eda0571mdBYveDrsrPGIrRMjmwQ070ZzUdJkrAT296
+UK6pO05bh7VMT4lojC4KrDMrEuj3lwXvL0/jTOEPJ4LiYzlPPwOjRJ3iM/dkW4P+8Mds/0fNVqD
L8tAtZh87oShEGLkmX87p8LFfq540MsRp7gvQeZ1TPPGes8i4YlLe4wjpKYK9QflcwTBemMI8BjU
b1JcBv5g49udEVlGibIt0YyisbbqwSpVi/hInbb5OrVT5HX8lhCdY1h2qBjmY+0T3YVHCuu4GfLJ
KNqKYqh/p7r3GbEGigiytrxhgSwuQqwzPI6rdszpnZ2CwGqhtrecWcp6LPDXP5hHiu/Ikk7TePJc
ku3JlyYywedr9bzis7Mmdjs1xDYAtzaCEf7N/yxZb3Tj2V6d6XX82e9PzzyNJy0ZZcSxE5+LlKsy
/aX4SQjC4pinZ/W2kZ+0jiIpOKmsgnV6+cbylxoixTZH0BeQh7NcCXz0nzVZwmWYo45urBm5ezns
Wxj5qPO/veWvSSPkIN8YnFZM5gv6NztY+KaGotMCa388Vsm28zphFY3fEVEZ5atfPZInMtiIlkid
oKI5L/k2+ZKMxCFF9ErOkiT1Pm3IkNAQdj1qCGH6OLX8Ef0OTzB4SWLD3t6X+v8Q6XHZpr0VOvsY
PynC7oXKECEwdiBwJe9dY0i5zvK7GZqTke7WWxCDTHp2hyL+OOjvKtV9Ek/4wj2v7miebVG/IVK6
PYUDPoHKUaDrhY6Q0ZJfqXyv3nOcmDV30X8rGBEipRCkEb15p6dYoyq3U3ONlQ0dvMQUD2Rt9XQx
eWkMO570xZrtFqKSyu5ZEpyZCsuzNDUZ44rie6mqE0p/QUvEJU7EfAZL7cWKQHkpKtefuUKOcfvj
Jg79vzdOkWdOXm/kUGi4kqpKYUnZa4SdFjLk+r+sPTX8R+kdz1ipyIlhbKCai60wDF6AOYFy+KtO
7p/5GdKc8FJAgJnXGlunXqB9GCsKSx5dE18YzHfyp2rM0CSN5ykNFDVkrWkVBZyMBeshQJw0nmb0
o67qmqgN4eHka+xBAJQMoKV5agzXiiQ+JGwrfumqFJPid3943ftaFJmWespxTjBB5KlLI/5BnNsO
JJnmMm7T7yE4/w6rLwxVmZKDUqHLkpFHrvcUKcTDadIPl3pvdeodVvE02s+FC+C+9gE1riyUvhQw
Y80kNVoRZm9rY8NgmKskTGXahYrxD9ApFd6UE/GHohAtZ8ufa2y1k7YVBtpyELPgWxeNlOwo3lA9
AsZKCorsk927FRNi6gP/G+nN4r22gZ/CNKStXPneNxAB5+LGwVaPIHXUlLtlvfpUvC2NvakRG4/D
HK+GkOeWb6/RNiavwGBnAYu4qJbqVBemgAXSePLdbk78DXJqSaVnpvqhgVYZgVfwNUPS6gQjjtaf
xgJLHmToxdb81jj9Q2vJpgbj7cZmsja+PvaCGBYFboMiDWtz7YSxfvt6uX0ydyfmdQiaboDoe8tH
pUFM1mEg40oCjPkOrsgSRUooRzt2GWScGTD/QQ/aBil/IZZjtZABoqQ5yvFcRHI9Ku8epfNOi9sv
78MvKRMcHm9WpXVp4eCRM+YTTgn9RlvhxghYbs18cX5Sigee1SCywqbucVjgErwP8nVNu31ZmpBW
3ztjf5Hu/t02ChrYjUFjhXkj9XMVeeGCrYC70+gtl6PuTc7+T1bXrdzWjJws1aM93E4l7ElH4ZCA
n7tDuWqhFdOtxensPVVkuJqqj4kUJ10HR13MEwrBliktHhRcSpdAXxrFsD6huTn/EeUe9vAIxXoW
9MId3Q1YUPAd61EtxmOT/NrlU1OLBEqO7bonIMo/MiiTTulp/y5y3zM+UacCQf3rHyNHCZnr8RRy
vulW02Tyq077vDmeXUorg/MPfHNmPtYgHsOM8pcEiKyJmPopkWJyom58juARBf26UMZctTwCa9mJ
7y4SQmH45eR9dhIIQTkjMpc699XPWXzL29uOy07aW8OF6NkDk7DjUHzhicjKvAjQbOjJR1CO0zNB
O5R6IO4sexsfKT2hGd+CDH1LTgRAQOZRTbtaUMYd68M01dPI2v9XPXHhW4tXKv89QzFHvnSrdTuC
nTxQZpjovhNrPck40BQvwlnGIZovcDCns8mEG2Ibiu4nfkzDFlntcfcyc2CZaiAo55frZ2Xpusk4
lcnXtbzv1BMIXmhrfuZZyBYLXlFVX2kJ88D21e7eGvx9tR5G6v3pSl1ujr3AvFF7jKCMM1lHhcq0
xIGrbIM8g+YzxTVg+/NfQxrUbxdVr2gtvW1fGZHTrBcNUM9gkb7ElMz4wtXFDW0wCmEvngaaPXCh
26sY4h2ArpAroZhSCSdx/+14WfhSMbF5Pi77Uqq/sTCwmlraphQlGi4j3S4qLO0huR5WvP0f1/kJ
kpBJw6SzTJpMVTBmbrPljquzKe3VuqZ6OvaEjqiQc2s5COrewglKmEMpSjzzCmg9zX5VOAiXEULy
4zh+3kkZlkl5Bx5/NBpm7osMvf8qC6rza/KtGBLtNdDoZnv2vUd8G+n3hQ3c/I4ydw65/z1CIGDl
D4n5hbtvkccRUhSCM7dyRG+mti1Km8kYhKnDgSKBcw3ch0By59j/Jo2HuBVqJj5obKjO2h+uTqd+
jP+pt0N5l91gFzQqNDo83nQ7wS09BHedDdYBTit2yvbOKfyN4U2oYKYzSis1H85c4E2BhYAdAkcU
7406hVG/KH5MXrndNLm4YgBJUwGdIyYQC5xerrrA7Ze+2Tb+RyQWERzRH/JfTpxsycrJN7E1f/fv
qFWXAuwh/KyXSf6ifUE50NevnRKS0beucjVzpeFxjIC5GTIGDI2w7kkYO33l5ktedusBG+TvTCfT
ZLsZ06KinnDBZEwcuEgnoBjd6AV8rwMjo4/0iL8l37TEM273YroK/Zdd2NvD26/nKO1EjHBB1UPJ
lE+1T3N2deHqgGq0AZ4OFC0x6Xo/6yp5kqAQSj4JFx/CdXBqCoqLfVtaiAEPl4825gnliipxcUwZ
f0UOMcbqPC5PwZdfZJossxa92/IDDtvqhkswgr3KpUmZUz9l/aImiMui58qbN67TwVyYzT5jjDxO
LDc86Iv27rRMi8JxoW3IALt41TNXO7f3KvS65V41zjuy8PcHtDHCxfE+kt1awrYzNnWSvvyJ9IWi
QZLFV9v5GRKSM5o8Z0peZfk0U4F4D9j3VHwdC2rXo0nq3DYJhI0x5C+q8tpGqeOiLrAHkRqnziOG
ylUs41Kqb4MjxNBjXl/+a6s0aDdFuHjyLb61O3O1ZDH+FCdcV1O2t6NjTFlCEz36CR2dIgkR6r6L
7yxLKdIXEiCWQm/g83FF48cwDLnB0Km/92VMV8xvFKt7VQ1njems5uHdXF/WKj2HJTM2BFncDBpb
tSGpxOUnQKvBMRRcvnuwJNXaUi8ZWJbMxc1Z4ajn86ojMQTVlEiuoyAbAp/iUnaLShk2JPDHRLhM
2waMZPzg3/t+474NN3kKZ+WU5VLnolaszIzxsUlKcfR4/s9fmJRn9q1zq55IFd4Ae8Ivd7f25n/I
kxQTJBpdQ56z8IMe/881cZKH9sN0PXCbpeYv4oGZyqPC8LnYqxrVJTsBI41De3Wm7GaBQ8/BZ1hY
O928pFZo0pF0wZHwGkUdm/VMzmxFFPp2Gty7WPJvpNzB74x4+BLr5G+EC18O4beljTqwNcPOApNG
kIedgTOMdA5nYtoE6L7pxlilIz5ll+mEzcD4lzWqiyPqp9izlgsTuWZ3F0rB+YKjUlJMkhKJ7Dbc
k17fHDxZ4Zb4fPgmj362woheLfLQtZvNRJC9VGt3Kl/yEF7oBAItU/I1DCaiENCxJEFVVCw1LY+Q
LVZArDXreJ3vxyG65SfPgf8obinjfcNTbx4VbBhgZijvLdbl29JVQOEvguB6/e9jS5CN1FrlZugy
4BZar8kjDRxczcLZ6XNFJQqwt1MZVVmBqTjvLfIzHtnXV1UL0bpX01TWCLbJ0BLEM/5uUO8Ny2Ui
hOLrbvifgbJu17JSGv2U8OyFE7IxeZ2LvoD1qM4MguPIEiBfFAmMpxnej6KA2cFjdHY5SMQfc1RD
YblW6XNcHqkUGTFy+2toGZpHNUbv9nt/nxKqJ+OzvgUhY2rlxtXm4XWMdtVGeS4VT849QQeF1wLR
vcYJBTGDwnPFk1xgHWg818yrJlleakabvM+Uu+O2GFdePYrCeK2zdVc0dq9XNftOywGymCnuDDZL
4txK107zc+WD4yZSQijKdf70P4frcQQMxuiRVDaByXVAE+tH7uVeNCj4/4qsPqFDD5qFCl/N6rov
TfcPIOTrqiNXp6disHzmsn8hYCWEuzefKsT9nnRCXHPj2OgejhZlDHPAiyj3JQo8V4QyUYyMqqTh
24rcSpF40GY+kcXypyi4gFMUBmAaijKftzhKG/4y9xL03g0DzCieasmVLSt0esYjiJgbcCj9lBVD
H17/oysT0hKeih8N6z0eNnG47CvzjA/l7pYnhV4EqP2N0dilexb7jZ1xY+diox2HeBsdTkb/ZFkI
aDhWRgwpgS/5yWeqaBMRGw7ayLyv7jKiGdCmKFCdgDwByMk1jNc80kV0n0iDByNS4hgHapzsV8vh
YeswPH//kRfIsHmJxKlUCgOl+DDQfaJxp277db2X/N7sgG6hf7wr7vwpk03ivl5TjM4GJ0v5Hq3n
k6RjxSEPD4RYEn0aYetMvVFI874ZIxFTx0kTXvlCfiI+8dU5Tw+OiESWa5X0eaLyPgUK1lIFLkP2
MZKkpA8JjVMkHo3SAqsJpQJFqomJYa5lBUXgZHaQ8M1AAkjt3oa9HPABbALUK0/mivRqaCGIchvW
xWfjPBTC7Hiqj3LQkAhar+k4VRyE2PYspiWNTtVqCyuHREfF/VUB8MYNa9QZVw/bwJuXRD+WUX7s
/Y5Cl6uaDQDJGD15ys3qKEmf+s24sh/zUvrwfceOHGtx4r4NBDKu0q9Ya99D/IXu3zfXsZlkX3B/
sYFX1MqxzyUAPpMD1Oiqr+d6xbkz+JcjIkDtnJNn6PXc015R0cMGSa2281K0TwsA6SYY/N2pMv+W
eNx6+H36q/KMoMrApIGiPAlNQ0A4HzuC2ABP2n5w0t6e76jRN0dtlAANcE7Pe+kqvjqlpERQwpSv
/L/03fhhzjWl2F2qUHLp4CQLeiXW3Y0+7AIOdf739Cdm5XtfW9vZKYCTtypeRxsFtOlUyVi6dxyo
s6J8sCQpYXEU5LU3htfNX2d3eiKPj2GCL6PW4n9GDmTd14GlElWwO18WGGOi7ZOJ1N8IDmIH0C19
hFh+8uCCN/yIuLoZZRHBTb4vjHZrpmrKv6qg99F/SNRkABUcY2FHeaFb/+sPGniaqArnDLxp1I+d
ztxqu3I+aKpx60L5DuYbDHPD/f6/KPh7+M1DOcGJ1cxxn716kDT44CSl52grNi4Fe7jFei54/Alu
cagb8aeMm443HzgbKUyTwkc0xxdDQjiiBgMebV5qEq2EuG6sEjMgvdAqOg/ilH/UWAwi8pxehO8d
vYikgNr/e+NjZmJTuDgl8SZDKxmlqMfxWwJNlJSR2fQNnegrNe2n8f6w1lIH6kGSHcUgcaA687En
A/Y1udTQ9znX0ihS2RLjvKMTuvHdgKoEQGa0lN+cOFY4AHNaJOi3np38zmJ7EDLSUu0ct0ozBXQH
GID/Ni0sZ2PUJJp6nEXxs2TMiNlrrZm5K6Es3v4mtf4ntI6PimLjPQj0q5dip994FwxD0o8OpHOS
BEZNjIWshJwjeDrBWPaPhOrvnNCPBrHlb3r+Ok33pHfMPdp6+GYTb37jLvzIsePWVqmdnGuSesbt
UbxGHgF1RoByX0xlzo1Vdofp1nqi1VrNxDhEs6TohchXm096XadZOsVbPMri53U6m9juhi4ERZrY
VQfIRBYUiYynYHbEv2LbFBGVoz0k/5i2RhkhZdbn9EPlZ2tjPKQeHY9o9lNOZ1XWdXybgRXTaPO0
FoUiFYZSF+4QrUMUtZ4Ac8LciyBrTA94YNRjpIsAcBDrsSQ7NVrXhiPYnOm2r1V7numhyoTpJLuJ
2Lol6c9xliQ+DAsUOtlZo5mphagbBmwK+wfgpamh8SqheGlwRiibQ/0TIx+gyMOLpg8mvuHIHmT8
qLOMjLh+Kqoe49ZaJg6k2oPpk26OlWfN3CbHSTQw25eyTHkSYW0v3AxuYB13joY2xoYhVNYou/tN
QHUmca1kDsyoXo2/xXbWQ2joW21/bmyf6LhSgJ+dFlcq5cZ9WLaCCZypl0bU18nrv33HdNJx3u0t
ax/Qt3y22lCmR3sVv/U/BrzxKNRNysNO/G34aTeis2vYHjlWSqH5jmT5lYF5pJfZhXpDJb7Djd3v
pKgbQagb62rM2UNUBbBm8++UGUTiGN8Bl4B6FwEDnu+j8Hhv8V7ZWluU2PQ8A+PVE1nnkS5rRZ0g
Wf8EhHEyvw74GZ1wxscu6PFNQnl+6o21bhweCnDhRkvdTcYRsGqKUk8g/8irm8RR76AvCkMKzaf9
aMlYMCLesjEgnLI5drLbivTFy6NYHcJXKD2KU3gvLeMH7eH/IRuiS5ZmqkGxcrGij53jlj1UIQYj
KwgVlhgQzD7rOZXYwWfM1/t3hY6WgBuc8NwQTMlFNrmX41airkeNxPFdo5kAB6TfzhJ3MxLIJh8z
Z+7wnBw71lQjejPtz6IrES8uh++Tt8VFYHdctL34gHDQYUDjgzJkfMaCWtWwEppAQIfVff+XeBt+
TxcWzD0Umwp3zD7EJSb0yn9kSVpk8no/IDGCQas7UAETKzqKU6XgPfZ0m6uQmQcimkbcRhep2mZT
lrLiemRMLJm88k2tEaju6Y25/44vYyuy6Qv+JPW889oyR5x9I0SqzsjX7qXqy3201AOQwAEjdtgn
Ucv/dntuAv+T9wm5WuEdlKGbNLh4Q7+1adbeULiTzV2eK/XCBMq1Ea/xuNGLMijKsnpVHiYXyk/v
3C4ur7bEtBy+Fdupk5jOAMPruflRwH9OdJlINYzc5eIVEo723J4IeDlxzeu73YJTQuk0tgHbFCBa
MBieB7jXWxZwfK4d/rDLKF6Sg3nXXZcqas9WWbz3oAouxlEDcdJYjBhbq+2NmafWNlQLPMp4GJmU
GMHN5OELhp+eZvNIyY4LU/H/guXQSpWuFWkwUIOucze0y+TVL5K6DCAQGBodRMCZA+iA7NGK6nXn
vTLExurI3ZDprcOsqRJ6dEnx8Ep8CwNtauSOu0qxl21hx+giScbCNdohgx+4ZXciOXxAeUWIrwi9
YdznXCVt6zxi6XhBWEKQZW1PDYcHtXn7R6yG+Xdv0vAqFnTiSHXPNWw6YjmEEE+RtvdZZqx/QxCH
k8/cjroNUrIpzzuLdGby3blhyPimBs/LwyiP4q8HuSZqvSBuiL1kaS4Ayai8G0yvwgCVHzSC8l5e
e+h2/lXiCTSKb8I8eH+xKW7sMvyzm3hP36nbrK49pOdn+FYWMIN0DHhIjG7zXZaWI/RIYllmvXPa
nWMuaBUzVwUf+J7332E0AqwM2Wv7pwyC3Y2+hn8OklriDMnEUFzvEup5Cfhcd16O/EhsBpLAOcNT
2t8LJS3xeuMaAXEoCCmAMng+qwZWPCi4nqJJsV4YVB7NoZaU0XHi6Spt6lVqUiiaGeH0m3GNnLdV
HuNjbkosJzEgAT/kKYbh50m/bir2wk8WC01Wkc91OxOBWcQpjXfP438yIG86YF5avDdt8nVejIDk
swmXxL7Qm1hjPY+4pSA+0JG2ltoOPm9U5BJce3g6PWrXEWDGPel4kLs7w1c9CVauAWQx1f6+DjoL
aFJi/JVyUOx+/f1JmGcJulcCAfj9/6RsPrCePLyftZIbBXe2uUSRBM1JFAMSaRoG6m3kAKl/cawN
NdscR7aunXci7Fvg5z/1Wda6OYAdi91S1uoNoWwKnS7al/M8KIEAMBaYfkCn0Lo1GiXatETfQ4HB
KeD+IFF8Be+4j3wbDq/zj40q4l+16MnJto4/LcsIdAZ4GTUOq/gz3eOAWQ3IFlZLeTFbtfPqaOex
2LpLU/VWaqPqvR1Pahut5dq0vXSHSWgtuoYLjXhVx2wYfcXkLyHFmePsUJrkmWjvoJ58vyvwzxAV
sRtETZJv6polWjNn7GBJCYUDr1XeO6F1+mc6mIz76QpMbjCEGG94djO4FmpvyW2jr4Cv9yLUydET
stv2M5impFAOl0A1HtHHOOeBVrNp8R0hZEAHbYIEiV297sBL6Nth1jJEgFMsHo2i5OHJ2HvNQSbR
f8jby1PFqr202ltIriyT7BFYSBoe524ckzPfJAT6LFCc3HI1GY2rdlkkNZU2Pk/sNi4YswMq9W+R
UzUB1O/xX7q641j/rOGnFk0MJv/pbb5IGWE0ZCDFc4JFlGn1CQmjf+oVRpS3kID6y5k97GSDKYm7
+gR9P4/RKZG7pC1SX2owwrXWycdA6jdvisJCWGF7q1uDBr+r4kWAE5sjgRu4RhUHG02rfRIhK0kJ
in+BqoYJT1/A+7Gw01CzTgC/EfT/+1Q5xfC/pPQPmGzqdHLmVZLeAx5aEj9VyBW5aorF6tB1y3US
z2/l9156lUd8ZA7oG4nNHoJc1iKDewX6mL92Eu2GJ99vCgZZnIGb4T2KOz2V3p2/lsXJaz+V5HO1
lA0FZNT8uG28qOQdlWTSCiy9bn54meW9ykl1dVMKenpbRr6HP2EcMilF3yTSBpprF739i5UtWKRl
57azkxqRrKcN9OmvpHHCPaLPHQSPkU6gbv0RlbJOUEQgVkcDuYKzp+H4Yho70kmSKTbX7vwlJ9vy
3sgUwsCeU6yvFyrMgAmGGuTn1knMr8tJ5i5P+mxLhIvaD0Pki3sjGbqku4eHNMvUB7AMqvDaJ0MV
fnbnMCuOwf741Jr3VM6PsVU4mIbUeobnb91B22ZMqQoASJN4Wrhv7IM/16bv/Akf//joH05VHrTZ
gj0kRY9DYweQXxspk/wrhAQpGFjqGXdw3+umF/e37piq/HDMSIxEF68OWmBTbR478yPINWV7/IBu
dOGHW2ijQahUJTCC9QMoOyZytSRhGRDsJbDGkhgjwQJVWKQokKetz1c6RuWE3bhEYZ0ssks88u/p
xjltsXCUz34pjllAt3588UORt+P+uyzVKluNR1w+4mmbR7/vP8v4MAFQzgFPDNTKuTiVfBnFEJqi
dpT7el/4PEmSI3ubb6qdEkzIWElue3pEWasuBRW425/Pst92PVUKUc7+gqJCwkOSs3lqR+cKGMd/
mpaEbpVDU44UJiGEAppe8PbIxonJkeSs74RqXJU3hZsdsRD3VRFc6cOYNJYTr1DbhS16PrRLIbgo
osqqi9QJRkpaEOCew6rswFLZTLafPmcsjAxGggvv+FpGKugeNsihFnN0cmZ8lx2eXwP+PgDEEQb1
IkDsGHXNVNdJxRMMwDQzln+m2cULYfa7NyEaRxcb4mHWOuZ9sARNRFD/GKLsqkvATbbrmh+Ava3y
Zq9uYwvSemow2cz9pLzEYuB22pEfcKcgivLvqX0tGasH6B4vtpdLWB5hAUA1myPSlesX5dxe/TUY
SeFdJjSPAgwztlytUYLYIosQzukJ8008YkU89Ff7CEcAAoXPT+RMqbKdH/vtPPNrKgWBw4lT2+pi
8400J+nEmwenEDRU5dXFxOci06VED+endj3zA+jX2+7vAxNNmLUMvTPkLCCz5pLduDn7z6a/dQ4u
xgyn7VfVO+RuAUjBUYHCGwPw5sERuMCcbqNh3ivEGZ6wLh7uHE5tsVKv1E3+S+M7zuYWKDEiNIaL
FQhwwbV/qeUrwFbPdM3KcCXoF5aRNXcWnr1+VG7jN72JRVCS1SGacuuOgGWiCbbiUnfk/uEpuHBa
SjPBv33TJGLH76rhAtXPw3OuTi3fG6Avna8UC45P1k7vi+pBvQEyXhkBCMmpuyIfG9y1MPzWeksB
A2BcZ5wr/xJwJSKR1LDhFymJeJwLB9fv8N84jUAlHL6SEln0kZvhZmgK57jsUJqCjsayrKzMgO4n
6MDMNK7L8fZ9Dzs1bd60dQRfRUfd2sguHXzGkt0ZPpWeKOPhHupTJ7mtLUKt4mPsNL5Cn3UXpW+F
5OI7AWZv6wXhO+RzBVyKejXWJ2Ty3z42OsnRaoBrb+LVatDI2e3JJ+Zbe7HRK12Z3DNBaDOlKQU/
r+Luh8u+Qg/jIICGir9bWKHysiW2hmWz4quhvQWJgq9UxJe0KTxB3O9weKUAPn5imh5Rfp0z9C4e
WwQ0HjdzWEcTfRV5varHMvUwlyWHHv4D+2vJa1d+jDNtz7bH709TmOiP/nt4vIhIDKsKt8ErBaok
6Nw5jOdK2GgzmI1XroMIK4/r5rHHzwriiBktw6Dq/Vx4C3KVVl/ZWRK3OBAUrSZp1m0HYMe+z6n6
OH8H39TbuBberqwDFz0x+LbUEVUIwVb1dVAeOoumrsKA1USXOtCKyXU3CaqSmZULwfITAzT8N6Zt
Dh/KjJZ8q0Hr77gt9eDLhyD3Jb9VhffUxnLDMLdptCtUcnDHnmuw049Dx5Lbo5n8eAvLiFqV7YEW
vtftlEenPTIOtUdIQz7/FjW70WS7Vi5mgVMHuePezBguKFb0PmZiZZKHmn3BUIi8ZcDPHKRlin8D
7uDbjmdocZbio3qtCVcEl1649WVLAVSEVZc9epI55MDlFhWTrFc9zTvC+EVs+wSfBnTIgvhj339T
C/Uf4t+4IKagsjzEfapiLIvePZXRnCrYYzOTOKLpqFGZAMIrW4ucdbTuzuRCkmQOeeQgxx+zMiQT
/9t9EFyR4UVGC2CsH1+7NnV+xNXAIdg0tMsD9DyLPnl2ybfYJidLb5BbvS2b8+2kp9VoJkpHxvm5
vQaI5V5iiP0EbddDeI7pIR3L1fr05NFPbci4ug/jj++dLj3jJxbJ6wZVuCQiIBIj5DcJ9UhDsef7
1LRdc3+ovyIlU59ynhvZ+QfLdlQUJaHIG2sWH4//CXpycVoZiopGsIcBCeiMN51aaDTYNcml9XVE
lLcw1j2bDTAkH4MP7OBoVejOi4pmCsKGoKf+YCLqE+bdZXitAyziN8J21f4WXV0KF9X4cPCScxC8
+epM4qqiYoprNE+6N9XDl6LEM2Rqzd9yqJHYsESJ/2JUOsiwr6eleEwfrLCe3xNaEIOD6PmpP1IR
hrXGF7ujdcEoQEEHJvZ+tySJqCvwMya5soKEhXgOfoM7hOspbpp5v8XDu7yQalRykqLTDFXK8/UR
NKfvhTWbtnXa4jRJnMMa266CwS29DnywegjOKq61O7prhm4jVVK1PxjyMK9yyuHg+ZbcsDYDMFhW
tNRfOu/kDH3pYOGx7MMf8DPoowGyc+jr1Er4eEqRTjVLBj8rfCb4v1LuoM5PmUW2FnKz5E7KYQbA
LrG/n+kNdiLfNDGJ5oJzSQs5/zqffZiz9qyILYugZoEjxqYT9oaRQhfLXa+v9fKgcVG7TISHH+c9
f6GwHjMRfFTf617q3YeqaTNyEWeAtzLybAjeeGHXuxxseYQTNhoPnSzfhHYzE1erFiZW+DoZQQ5a
9EHbnHdbif9XgZQxBTS95mLe62RMEsZtsLeFF93e2GbHqZDxYmVmpzUJ/k5MS8vHQlrEprvtqKNk
L0vhAIGayO7hSYVp0Joywv4adoPNil3Ke+7kIaY5RtumxOju5OOK61H5cyPyYqUlYmjOiFgMWsnR
eg5wbg7ZS2i6mHWJvpWtlr1NLyi/+tQQDE+Pyp+Ng5+Z5olfdRt7afv9Yviy47RrlkHKdmvHAZW0
FFQc96iPd/JxMwXRAgFKSKh5N1VmBtZqSnHLf95b/OLiQ80Q8XPE49tWZoUgnpo20T8MWcB2Jerq
q2h49odsoPLGgsm9kdDMuBoFPJsi5L4vvwuwZW9e/4AxCDLreW1Chs176sC72P6GTkJyNh1W1gLo
OF9TpzIh68xVClXeM+2iRs4briIkRaRQCW8cb+ChX5v1WWncryrNdemKZLhrR7zpzua9DgvU2+f7
SUdhGyRKlUdET+BrUwYj+hIS4jCdw4Oa2wCBBjfPHhblWwOSnVZRn3m10tl+jRXXrT3c8wVGyiWu
RJ/Zx4Rt2hHR9dhmadSw3xu90ahXnznNWdphQQDc2Jl8WQ3zQEyWlttiPsDJOqNFtQQMke4zAJpO
Xj/QpL//E3lMFqqxW6GQr14Q0J7CtNeXGO74FGGZqkZXVvfQPnBWVvcX46/dn8mOWDm8oQ+Z8WW7
PnV1Ml3nQzwbR5PjvmLgpjZ38cM7ZgVZcNRWH6E2Id0PD/lu8PvT38AtH+UeqjOrMkHI2v2mtuwZ
VmNtKZxbw+3W3huw5mcMUXZdcIJACevrcIymNQSF1c01vqcVfmWbO4ORngl4LVWzb3FMQhnhwj2A
es8cs8qYDf66nUvJKiFryto88E9+TrCAvJuIGXqvg/WoGIUUpEhTj1jUDJYy50VSL5ZoSZqOoUMS
8SbnyxNqRHYkjiMUMshKwDNOQKTSGwqDag5yABhzv/FZ5fuUGcZotYOl+wd+3y7aygO9evuWshmS
o4oGWlAGbG8hhBGwE5/t2xpgAthPxmJtExqN3GYoIhiVfKDpuU3JKCkJAAbFjq1DGHA1sWyHLUXG
nLByD1Rt4WRB9fhhxdZVy3UHbQzpUk/rCbwL0wkG6ogRherLuChV/vJO92RzHIwa4S2eDMJIJzPM
SC4DzIhR/yricylH9v0gN0Ngu9z+mmCkO43jiNa53WYlvJ1qODS709m2BjRTnUyjoNpuFbz7Z34n
EBLADQ9XWZ60K3goBOjLuF37fbCsWqQozhzN24h+lnQ6tykAVXXKtGllA9UYT48qh4AHkrJYZVsE
m442uMrKveaoeSlY5c8NDaI/YCxvsZw1geOygtI20RK/T+y68h/RifeiNJjgL6Jw1aKw/MpabqDw
TBvx0/9BY85pbYJCrbipDisC8fx0RnOtDJKy/xbTZn4xzd+u+bOt5lqukBpIliKPuMFvvip8Qo8y
Ye5XW5y6dZnG3dvh9qwad7pkpCj/KnkpnXfJ/VqNdN66mwmKRzguuKZ4FAuQUmrxRAx4kfbMYwf0
u2ZMvnFK7EKMRltUTq0cia58rjFqUvyRjPiW5nHn2ZYhp4zC5jSwKz6YXYISWAKsFK4psdpFQXy5
fQ9ixH7DrVoeM7ZPrOWyDO5r6f7/5DTxOQZFjlxQpCx18qJWyh7QdNZAY4m15B5MkQgytGxpg0Rv
CVqgWCFeuvWBXoO1/gZQhp5afAEHMkoh084VMDz+mgMxkZy4n+O0VMsjTlHDwdOP/jFMRKj+WFC/
SkcpV4nvqS+cIrQkrYpnJprU7TWt5MrcO9+q7JUMs96anV6MGwO17D7NdUXKpl8pEoywpNWLO39N
diRtkWdQ81WAxoKR8O6gcvP+1zaDaiPK+JxoieczKVb99j6LF0aO8ZJHbtKWJz7Xg8qJA1jQ6F2w
H1goyn9c97yQL0ANqq1s7NKjS+Jvo4jJtgM20fhVM2myf4X/arbepvRUTcdHzCLL35ZBGsrTGAwq
dQH61ls/X5hnQw0cXY3x0lfbsBR5knKvHba6xMRmyVsI2u35qThzE0BItiaUNZu7iNP0mTTEZjCu
20Dx4dLc1Tg2+SBn4Ruuvgl0wzYOsSBxIrLk9Wpy5ysVOIUGD064eyanM3d3pn58JyoTN85qnpTv
3gZPS3JFTwNvYyHbjsK8KZf18maUHCfIOOQ2spOW9F2C3dbG2anWz5lU5yQvN6JgEEJyfPJtLB+1
zqGCa9SVy/gBstcskhrD+Sm5IEffh1q2NccBd73iel6+Qpofp4a1537VJ1BzPIaA/2QwlLrdGnBV
6jDZU7XNZR2QVB8AqiUxg27uqR43PvXr706ELmi+Xg7bgMITnllgz3vfre1P6CHq2RGnsKydxEwW
gP8QiMDh5PKQZIULRUR15P7o4wW9QLVIrpeNq3kPhlb8lV42WKSkaJAnAneyIJqOzYlCjyoLFWWQ
kC3dtdcVeO2abmKqorLbv9o6VSXjcvSCC/WY9sJWGV0+317t3ZsMTC11REK5r/BhVYaneGP4xAB/
NIpIEcBCyjw5jupRlOQIWSx790cQpRW+B1E/0cDz2rjDGsNIZvcgYm1d4tloacL/PMGp/Ny6/501
Of3IzwzLcL//mSjQSB0sNlDmUkD/pOx6T8s6RevpT2rtAThKQd0BkiO8xzMB58caubM9guwdue26
tQp9ACNnkFCJX9gz+V2YyhVK2RhgKCX0lHr0+T12hceKI37dIQf61LbKp6Jaf/0h1vQ3u8EhgPEC
t15Au7tLv250Wi+Bciibqc7cB/tN83bcbWXNCPUyhOArM3B02Rvp9TbNvsThKgzwfiBlqUZy3w1b
yUkvNHoShKA8VgIjNz3rbWJK6J6Tsm1NRW2+2zfOffvRV8/tQ5o6O/8Vvqg7Kc9CraRdaZugOVJq
MJCL9/rseLTfg6xdAB8tlzidgmCP//IHfNDJK+d9NYKmvkkzE9wBvQ0LaaXYFj//uEZqutKMS8mW
O6DZ1SN7PboElKOaiG9Fim2p4j3YBh5aIlAKMel/4BfAKBzOqypZZykHf4WUGmKFvaCpB8Zz2KCx
fD2mP0JXZsqR7419pVyiiauhK1LVinO4MqOb+uY9wzBcYZtj0srwd9Wm0VrLg5O6z1pD6XJ1nh/i
KX5LpRd0dFP77DqNW2SqQKASYBuR1XTkSPiy+89BFyr3LfzEr4BXaw/jbh61ooBzp+SEg87n+CDZ
EMyMdbWuDrGClS5Oa2Xc9Gom/hzvFxn9BtuTmCXNooDPmUP3vKHh6/9cBNOUJh3StcfrEo6IyW9f
0lzITnp/LHVEdS6toDKXUqoxoYj4AYIIzel4FSYF9pNBoHJ4bPO1fZHfymKBVF6XviFqGenf7qud
V6rK7XCaS8S4I8ybdhk0beV4SBn6xBObWlVbzsqCIzSpL/aYSl01wQVdtlhZ7UW9Tb2F4LkZUBsY
RxuUZejBseHWXPPm75MG/EaWFXRti4kc6c+zcQLEXkMK/y0KVdKqbSvR0qacNAKwvBqxfgARbl/7
ZUYjsBthH4gO6xfI41TKd3zuGRXpE1qh6Ng0k7l9q+eEzyZYgnR5qmTVqhlFP4uwmT9hbYF9EZTF
J/O6EhtDxJ+Y7cdal/Q4guv9ZmCfgkJbFUK493a/W6ZlYiS5mqfI6OzPw1/8mFbfInW3rHY7KCK0
fwFckTKjaSkieaxM4vjdmrY+1PTsg9KqxoRcT6+8yV2j360KrkMaFw/s3+r3J3moHlktfXMGjIZw
GLFts19WOgWrOXo4RdAtojzmqqJOFUjC1Zonez4Jl7RhqXxaXMS4/xSBlJa37805BQACtHP7JRx+
4HGKyl4U5lZQBH/BVe6z9ul/YUuhkMtQvJsv5QAA9AIpYEmyYD19LE8Mn9Fx4daMfZWbBJefj3KL
khB9V2i1VdcIo5gBj4hm0SNCvqJvJnC2k2u41RrH+q5zhyr4cmi6zrOQdAw5MaNuDccKmjGXSCJk
PxuocLgKD8ruaPSumwWFhhsd1Wa9LTREcTifq5qLQFlw6yNCyyXoWb0rX+7afPVOtnA1Z4V/cvfH
PDSQbTT4nkJdzJVfNjjmsDN3OqV2Jpgbm3PgSVxpOcquhfapp4r6sd3gmgbyk33ouY9bYmwh2oPA
9t2InagEBBRvOFwle2MdL17DMRqGjvDvFrF0udU0lw00s92EBqoy4SJjyPns/oy+lH46r1Tb4/mw
GdCJk3QwgbX/77Hi5HNkUps0g4/3u6ZnqBiFZfAAaZQYIt0kcJVIEQi3DHmB38LuiWQYCa0Ocm9B
7DrHHejaT1FTjW/oM5zrzhZy7DTL7oakPwU+J5EmHEDh9UShs/HkY3hFmkgOKeXmvraprMgoXhps
lKcL1ZNEUGyMWGCxrctCzRXiZl+q/Vj7m2o4JCxnH01/OQpN4yj36sDokvzjs/015zuDG8fA5Qfh
ZIwwTobpq2vvPS5wQHDBPAqkkmaGJSCts46VBMUEAqJfGU5u4gHxmv3bE30gQ7k9ctlqZy4snN8y
czX0SKGLPD8bVtFDbpUedPMGwqizl8ujK0OcrKnEb2PvRwooml6vRHHlfc3RqkZlclOfIueHpAV9
NJLy5VsUHQyYOrGAXGb1DUG8dYEfetp9wcRxlFxxRUAYPJYY4YlxLyMd0279dcJXaaQa2URPFC7g
GUQCqg54DqG1rgWUNqV2X3uOYZrqnQ24lEbevEwgmJHcFVCLcON/ylH2GpTaWIo3eTYRbrZLXbCl
dT1zZtWIAU50ujSSXn+e4g2u7g0wUl4amQdotrnWKkL2icVb4yE3HmNBzLzroucmZjCsrIXvkcp7
t4DJIyvVhXPEQW3iUpABVlfenQcTKYeIwiti3U20w5jC9P2Fw2/32vMtvjuwL7vfAlbx1cdPswDm
UPcONflzNm2xY5FzyyNxkIb350awufwOX0AqL30GgIauWqveaEgzt4CY5qal7DZNb4OWJKf2L3se
Xh/YmRbi9IcD2me/eC4EWh2LNsMpzMLFREXbL5ZfAVwa23k2PblfLxd0Xqo/VwtwyjQCWOTEfIvW
rjFohinZD3vpZ8fKfAw/rL1y5PvAGXKWlgPJN/LAKMnBQzL0cDpktbwuyWdSXJ7wa1umHjps085V
IkuNcIu650LJN0wBhQ5ra66i7W27aPTUGwgMysogS7r/N5JSxYxVUYoX4mbYuD/QInRThnvZFknN
NRwtN04bVVmh4CjALUH4exesQwlM64SZpv+Dp6tA+IZgDd0covwGh82a+H8qJbyzZTYSZqgUUG+2
NcxumiLWHCy+/fNrRnm22qj+gVPISqj2rsdPbeoerJDMddQvBLc2f1biJHP/72J1eE46jc7eQAgh
wA1h8OFJVkxKoTiz5erk3WFdGtYC6SfKo4b6c/hRyHhOApPqRW/4Vkt0AKtw3K5UIjriPSL7psS6
nHY+3Zl2jrKDYnVTJ5HHuY4aGtkqUDpGCYeB5KFg+ogCt8HKfNYh+RgletK5I+ElP2JZne2kt/CC
fm+ZqpflGJt6WzHDN5PI4A5Lq4RMQ5ds9L136vukb8LLh1zA3rNX6Pf8NMijj6UDoov/okk48pFU
2J9tCaORjcik3M9GZLwupavtnarcKzT0P7S02ykybaMvh2yrEPG8OZMFiJ3OTVUGyuxhf6h40GIF
Dpy+2JyMeA1FT45+3z7CSQrXfPFBsWsRYIw2J3KbLGvAHUWzH720vaa9ZvWDkN0XrWdAufmZF8nx
F9xgB3ndLvs8l6MXAhpQCuWd3FoEcFggWhs1dH9son9+6Fxex79IMW38AbUoav/tSXgn9PrCAAKu
hffyZQrMMQa6PFIwVnIkXf4VUnZ6nQSjxMmZM5ApbmUeleigitgNkPyq/bDzIDSR+U9ec9CJK/Hz
QX28Yx1zmjRj9zY1BThF0dcPpu6q6aR4HocVhUmf5Q8jjC8DgNf+5I3JxxNQAecAaviPDKE+bVCZ
xPR7ju6ZffwxYI60CvT1JS6IGHptCV60jc14V0LRMZ7NePVZ/DNBqAYEMScaOFSiVClt8WhVLmpb
cM3PfmYwglVkH0jptNSOKpomUnwajjfuS2OxsXzfm9oT/NURIQcFpOtUhdMo0NmjfegpX3aKXg2H
b3tIzjr5zC47/ec3XBey9IFM9VuAiA6njb092WQggEw6iyxwr9I2eY69NTrPxZEAKUYiLLSfBhqL
XmIuJQvXlBDzYBgPvZ4u+EZBNJJcUB+HzY+L2Pp9F2vDlwoqilJyLiVunXNQAm2SMnQakQYBBXvE
81iqGPz5tLrEECObgxsnDlb84zKxV3gbj2pbu4etRAESbgeiIRJSc0I62KP6jJvW/pNb+nH4b47x
RjjuS4hySVGtZaApS51bweQzMsrVPGaDl1Rrt5vg0TX0AuuMRoOZaBidasUt0qULVZjC+G0PtkH+
aRhst5PxW/UKd78oPPxTPIc9Wma/A6gnpmxN5GK/GEzsrT4vh3+rN8WqNdMScOayoDwa3cr0ZT8D
Kv984Li0a+F9pBr4TZUpEYhOaorOLj3CP1pcCXjs+SzJx50TwDPRD7vVQiWhGG1fuNkq+8DJefTd
YhYMuchr7Y7TAcg2tKLi5DoACpZFMvWXlxZd4VPx9IebUes2WjvCWKTcZwnjtKz8RHqEqVPS20Dr
o2nHvOwnCmOa/40jJgeiJE+UexwestDbZWpFUS+sR+ke/ujxwaFAeXs3nwFbQzoxQvoD82zOlYIi
ysmGXA8opGU1Nv9JfCxQ+vRQ/a2weayHY7qWMvwT49jQwV1Oni6GL0fOdGr3m2z07eqlBjhJ1A6O
f/dlywhP8KvgeBk8b4bOONI0M0g+9t9fXoseU47iwr1ZHwCh9MjORdx5vGxTYWH092ti+rRTWvw8
06jiFJWVJ2v6oXhn/naB1/wHLxac/mmkblJA6MMMCKIaY1vqyVLAP1LLnkS4Nhnn86RbOg1Hyc7N
IUgU5MkGFfxoUqq85OC2jcmJO5cYy9MgjAKowkcJos7zi3zeG5QMIwy9yV0xBc/BWpK7buSLmDmK
AqR5yWz12j1R0TfBJOssiLVQdAcRz0xjhxSQKe7W5qKn8AzCKws2rxC+Zja5l0bVrElfjesl57t8
9NshRD1n2xc8mHvxpMeodWjkyZmNPguVnI06Tw9ZNuiwpOBACOqCzSvNf1BSdzoCagGDMJ3YK1lX
6M6O5jCtrsPjfALiNYtzvaK7EtdsACUqs0sfpGbSQr4BLhG5xQPn1/PX+Ey2E4TkmpxwDj6Wq5hi
rg559HwMXLWTFXPkCACDvH0pZZyuxmAtRZn0gW3eEoJhef6BPl6BoYIEavrziWKPLFBdyNlOnN27
AtWbiAsyfCA0ai1RjYxC1uOccBiWfHPsO933SD0UcbvYxxxalyXysYccZ0yNU+J4XAIMsZAQ5ic8
h0lHV1RL19g4SgY8TY4Hu66M34z4T0R9T//I1VtSlFlo1CX+tvgmyVojljxKVpM6kJ3VAw5YR3r5
0JJpUBTZCKSJ8GOOwdw3lvNNWW+Kedp8UrSOOfCeHeU/2y5JKrt3L/I5v5Ul/1/9WwkVula9WycT
st+Fj3vJ/pNqWniEtBrbq8ib9kf0Gpgqi+H8Zlfu/4uuPu/R9kBykNYfDVEwjQLynZnGcMLKylH5
bb9roCprfHQteot1gUjDxIGZEaHNfnOfD26r0HNfl0fEZh0uoMMr8i4cku/0geoZDbR1tDU5pNLV
wxU/0rrpGjrqqVcQ9D/SXqIIsVa9NSyYOsuhqTe5HfICnmmSo5+l7shdo98F2YNoSsyc0pVIujjk
5w87wy2c8btANQMy4YA/YywZ6//uT+c5HukTJ5o6w7QnsgsXiLxdcvtDxb30bvsoG7KpLqc+bD5g
Cd6ljYCR8e0a6UXVxhLjNhYy+VBmtKV+QVl/tMexbF/8AnZVjFAx9k5iBtfoZh8ShgXc7CZvI0o6
DyKN6YC44+edf2w4J0BAXAXdGD49nRw6BHC3xIJmSShpCt36LT3p+fqeVXz3s4JZz4O3HXa/dAuu
+/L7q3tesjrpGWhX5u20bWwRUkn4z+dQW3ZQKnFZ3ZMcUoYKyWISSuF1ToRoBpPfLjHz05fIk9M9
SbmyxxBiaG4jMNx4YGUMP72F6f1DDKhGuHz8m4Ls1awlVzOsTRTKT8houoqn1EGJnylyhWxc3yPl
bxLQGwDVwsisKG964r7FkroX0IrY+1szBB2X5Pv8O9htSh+eCVKMx3V40BgejKW1SKBVyWuqLMVS
LDo/bLP0M34aPsKhxM+4FEH4E5XhhqEm4Em4smFQVJmjdrvykiV3ybxVW+cVgqyAym+BaTW3UaMG
/gYn5SiqAPf+2zGg91CyGVgnf51n9o7/Wsc4BGdsBIynRGf2ps+5OEp61sKWaA6Ky8wEbbOcpfIW
hVriJvqyfL4gUz8jzG2tSO0ajTHhY1sQrLVPvrS2Ft+13c+2cKTq4QfWMt5D3azzHkdHmGQKp/DF
qbbjblOKoUHLFb7FnYXPUaM6BeKDDA77FAKcI+1//76zcd1d5MR2dAs6nRL456jGbqYC+EnJRVnu
ytY0e84GksZO4s5CAz7t4uZxP4DO5RcbLFS8AcunXIXgTrpkuP849Sid+U5AdxpylhjV+RuWexfn
1IBeOB1zPVxPDkh3Wu0w8UdQWQMgR7CJrWQjFUNxKFf7lK8a8uiqKXBOrZotwGTzo5pkg+uCIwf7
/7r2DSA6c5N07qnn7Ln3Mth2KKTVyH9C8TVgzlXYkAxk+IS5LHCB3Wll0QFnzL7KBfiysvYECVGn
tol8gpTJFT/SgV447dl8PrrGmEIsMI7uj1pIW94d41imUjeyeI4orYxVrKYJ1p8c0mvPlZiejOqb
kwpZY/Nq870ShVdGpcKM5Vv0d/3zUWmHAgETKJk1Ut1UxLlzI7E/zDng2UaM7D58LXTMTrxLpYND
kWqyIMJUANO4fnjnS3neFkL80b15ueiNQt9eVi1VUZe6zCJWO8PkH5Un1IWq7IQd0KAvHwSRzdy7
g0Jw7suH7uQU75swbQZLi7qxlcgsAI4LKaMAo7C8FWb2yA+LydPiIMYK2C3k3F3PKAtcPETt7GXk
wMT6OMpbUJSF//lpw5Tf9md7PMi2QSRY3oXQBMp3/f4qaznEH1BUtj2yrtZ70wJgrk6Dil/I8+M5
aTLwu2ZMp/dzBDPGZRYH7oS9fOiNkw73k9rKIXGE28iPd/vnJgj6rVSyY1VaWM9lk0/MU03usYi3
QAsxkAdNVLQaNJoJVVvuQ3KsxCPssImn0uYQ6GkUGBQiVcvUzEBSLnNszbMitXw38eJa/tVY/mWR
EshFERXRjqgWeFv30Zq45mEl1dPbVQf0lBBpIgC4jhkdpWtGryca04equNUgNKP9PYFdNo0M/yhb
S9V1zIOjy1SJdYdqcIqU5y3n2wlG4cejtcAZhJPnZMaAgRSDef43hJuFsdGpGY2akj184POh6DsL
KDVez6qE9i4SQPieZGcaFcePESkDED8Y4eyFKj9avGRYtmb7vTtrOBIzoJO4InQbXSl0KImolFCl
AWF1GHTmdW7drul/eAAz6HIHeUds2MoPNx68QqkT9FSNRKtjMfgtPMKGdKpAci5ZsNzhm7vni55/
IoLskrlul/CWMXExR9g224D6JyCEqTTzt084FwHilaCfP+kCezW3rx5hbQ9sGowOfhbfJF85WLaf
eUzzj6gqhspdtqiW5rvP+lSnLpShXGVZq9VaK7zuyMHA1T7ZXbHiWp4sDZ0EQUZwTGCK9vPxtfqf
9XCraieBeQXNVXMQt1/RiD+c+RIpD5yQv9Ik2usmmioU/9N6xRqLXtAiC9CR3PRxYZ+9VmA9Xh5V
pVgGknTAJ/qNm/MiytWr++FOnKs2+RKgEZdOdMZCbTf8LkIUZ/HTYNVCJh9Wb95wEuOYp29Ur2wh
sZWbctp5JWb5ReIX5V2fhQn00Xm9MyKJjKP8JifpmfAbgUdMnqOexxosib6qvfW7nzmvKBhOTZ2Y
hcRRmPWvnwLow5Oq6WWHQWi2hLQKHi+Xg2kWqj80qGhr6lSIu8x3d5aHl3HRcsB7YZIdC2fqGIIz
gzJW53WMAyvJG9S8s4SXz4XTVCXLloe/Zp6f1nSrDSWIhsgfA144sQSNnCai10WsED+x/AQrzWuk
sbXevEC7ySWPNgcw4AVbPoWJTe+KvyF1QdQBRSC2WSL0oD8kswptqAurswJNeNAInKb4zKeNX4oP
KOU+g/q7nXuxT7Sgyq+l8Uf++e//d5zT1T6b6kBMu5SFMyOET+PrG+pzCDuHeVZD/VLkIaJbumv7
Yr5L7JgdHFileOsTpaznR7xEHkTc9DmLbPS9z18lBVvcP3DKA08vklaKzk1DS1OevrIOtAVV7sbG
lA81OleSho5XIYIrpoC8sdUHsPiNc+K+B9IfMst4fywDrHL65uYyOxJ/VGOuNpa5wHBSlwI0EuCa
TAnYpwYzkFbh1/bWMPXZsJXBzGMa2bjDLWd/XGTsCk4jm2X13ass+6auLZrKMlWY23oRjXFsjH8r
r/ZekQwCpR3W5Wk77710cDjwO5lhOvvFnI858/s8fe213pAesPf5jNQWLnjv+eP1LsS0Vs9F9vy5
iosXgo43UZt/Eql7GsdE5tv4NlXb43Mlo86AAiRaudLpNGV7Rl0hQJsyVDGwdRgw15plyfS9Sm8p
xdPIf87wFGk/e1El2evjmoVJxrz4n+Yu2ZWGniLCBt+rMV8JtTZJ6qCi+VHMkhAjmrMyVB+SE2O0
yoFfvimgLUQYbZq+XsiEa37qrhqp0miHteF24RtXsMvTSUCct1YMyuZf42dV4TvVd304f+ohBfAk
Vkd1sk/v3c4QSOUAAZjoXYyMy4onNV6HZASND55/qiEOyOAnm/PmENIHnugb4PLtFb1aVJa0rpkE
i0N/KhSrXa8ZRg5pwsMuxSmJ4MYlDuexhvUvYAMAdbNR2hnW78rRO6mQkYb9POG7Au6klodg6VZr
ZK+QPIA8omzbYe+fhFQhAeMzBrujwnAMdbOYQuY1+AUH7q/HJ9glF/p7zj1SSq7wvvyR/F/Eqe6b
WcPqiCNAVaa5LFImtm4VY80AuVgJXtZ3geBKvnbsLqcnH6iN7qF2qlvVlGYERhcuc+7Nu16ti4DH
mA2gvNKPZH5HQmQzCqKOHECVa9DYUfDPSL7wtEVWGF4fXIhlr/acPtwCM0nB+lHeK0ZssYANzUfx
fI+z3XUDhyyEjNe+bCqIOntgOMZt6jieoINbG3ePn9waPC86X0I+1c50YZNv3hZT01R46ov/HXlb
d1ihlugdaa0ripmhsv5UFvY/CohVNb0AhFDqRpcrYfV+CMKvFMJMHBadmPHkdVYQtwXCHG6fzL2W
5mMSpv/bfytzAqqrd5MTHe73bWt2k94L57/0PxBZ8hCITOwqrA2OrItmMUwNb3pM77OLYF0+VrWJ
gYIztUL9kC4n0lDfWgAOBUINvYaBQltiBbNAkohbunTI9bwqE4UsRHG5RtAqjQxbx+jNeahoDCPu
Sq+BePBp3ZhF10md1lPljmvuF79zru1LS0Ch7ESi1uKsNmz7mkkQBiVGEWL6jzZtiu6EOUdU1i5+
iQ0Aesw4+mT4XKGUTCGRTL0Hn9oMdhrEjVKl+LyHuPPvE0BKWAI1ILK/u4Hk6uJzZLGiSSS4VmBD
jDRSHnAkoynjLgro36XFRK4Qa+UCYDdSJlpR7M8/5CSpITRlvVWAYFNYQXJJqdB48YK3jyWQCl7a
YEOTADAmngcK9YBRa0qPY7CdHbdG381hHSiKNp2FORBOToOQupbL7kS6r1fxaT49mJuTZEaO3SdS
MnDHfFfhz8n4THVfJ/6QGiQDfiJQsDs6XNQ75QiDEg5gkkEDHy/LkMDWQ/BLKQ4a1/x5gxQEqcLv
jyTaVRTcknXoj/nqiHcnj+Q9oq/mJsWG0/794YZ6wufIAToO1W5ebIcExCK3zIby1ospJrm2liLm
eca+hI2V4W7HeTHnzaF86u/pync7TwNqg72T5PNQSJ4yp9Y4g9A18j+Mb5a9HEpA6lkWS05smpa2
L3J0nH3/RLC10nnSh4zeAoZxNh4RqAUXAgNgqHj0ZyAP6QXG18Z114bzKtNk6acoeWJYQ19HmhND
u3bZx0E2lkZpnGZn9Hvu+7WTUfzEkdbpTlZSY/NBt6d5XYVRIcDBgwbUhakn2U2wU0ipHzxb7Ffq
IUKgAKA6h19SLxXXgQTUMmbkTv75/0/8y66WdXeumP093OCmyu0SHpL0Kv/3mExoSd9m8HrCE1FB
EaF0i7lD2kWC6T4VUlhQAKgKdT7GaemTfB39vElO16jiWpZf3bOsjcVr4J2+7KtUVXmSrXBzDP9B
UwzKwxlhiKH9pfoCW5YTt1biIYpZqa7IqsJdyA2KmcB0isMbVXX+mOZqazgM5EZp13YV8mmgh3Pk
jpm7rUvEdcMNJk1uBH1H/0cIqy1f0saUIBZI7dDKmxVcXlRhzsHb3fTJmGXSb0EP4hO1nVJNMo+V
kwHEYtYDiFx4xbIWQpc0/DapdwcuN7j372d2vElQPeuBOkQum7ty4RjeTdmRAKLeyYt8po7DlydK
k5ET8JtD6gxwIu9gVDd6whcrCTYy1O40XqcpT/s5hnBUW7fYxhTNVc7X/vAOivjJnVUQiDcxKZvX
Ih/wBd+K8oQdAiKOF25725weS4uaKVhGlJ6XN81LJyLOfIWo8kLFStzcMBrudmuaySlxc6FFqORb
WNxHCkrrcpPL6pSIuqI6iFgiKRTXUxyWwZEfdylOoTAL3o0+Wlnp1LwtpEg21nTU201f3tn7QYxr
cOZdqmR9y1wN0JRWPzFRl2sMV0iplBDTgbzEx6R1nlAl+4aCGUK8+P8rdYXyKXciUyQaocHyUQLi
Efwk+eT39mYMIKdB3ehc7WZpUd1BOSKQ5B9bqI7zeBvtkf+LxFnFOwgRqdSpNm/ijHCh3RHqV6Db
TUZYnvFsM2oI4cy98gfaAP84psgDJUfKwp6kjFoEaXKpTsJV2trf/q8UF98Y1DV8RfiJHi1OEyLA
cpXdhlagqHQK5opo2ehG9m51ajZrdch7J+HVZkKfP8r5JuRTx5FBI3ci+XA9rwu43uTk6V9IkG1F
/rNU6Xtk/KP6DmlSrLjd370G90qgaWDWpoIW1UwIeG4IjzOcTI+IV9dpN/qvQEtCUWDrygH9pg/k
zLlUIrdVlUju3q5HukXuVut/LHXIs+pmUciyDhvcKbMe3QyeEQsBKQc/xCJCIFSyTo4I5sSBFmc5
dNkXcYJDRZ1sr46XYDprF5PI0SYNug0de+hpsvZjTEVK1sVt2a4HM3sv1T48WsPZ1AbtKBNMNzMi
UiNJdxFJN0c90/Ux8mm2lX6ROV3gazcvNV9OfdoF7vQHsaGfbZtA+HXc4rvJ9QrVBW5mSOKwh2Ro
/KRh2JaugnmVX5pC/anyy35YOSLqCTNql37vLtEKNwHFCWC/XEPuzVSOY7xcvCVqs5YU+LgsGJpb
cmvq01JIxdfIVoMMOp39jnwDcxavBGu9SRm2GidhLF3FvngTiC6cf5r5m93E6rnv2qg0TI8678f5
lkUgoJ8GGrpmcNyif/pnnDHBK7H4Xm4wdmA6cn2wkpcCTfYzX0xpksy95mFOeGY3MGf3W5gipGI0
R0o1ck5pT0gejP9++eQapdMKnEY1upak4H3+KWgzZfNr2lCDgwk31HeS1ytrdYBVlBXZqxOiKLak
AJQorgpiMFVduDonZYB99pC0e7WKg6OlVm4Q1e0PT9ueC3X+oIMhAAHpGOAPO4EBR7h3h0oxuNNC
ArFqtBlgZxfVYfpIO4Xfq6qglFNZ4QRMchuFIcr8NutY7voFA5dpXnq0DAzlObMfU5WXZBRybs0Q
K7HCtMf1HGS0xUh+7zNZfySrrlmPP+jAoNAOICOii8RpI/ituiqjgI5ARTD/1F4s2S2yFuVLmRz0
mB0OTXsdVB8oi9Lhjhtss53dbun002NUOE/NgYHowCNFBeeawZBiBnACzDbPgVE2FLK3HU6BFymU
gz0f6QAWFtnHSAjeFmqU3a0qfud5HIQQn9O1wK9ADb9FEwNXy+fY2jk/b+KHl5go46qSk6PZ9HLL
VZfUvNrXVSeaVQHsOkHFNzNaUJcFI4k2sAIKyhVApyJ2fl1/Yitutf9NE4mUJfn/1F5IsljA33C3
t0VskR1cOh3EJImnQ6MQ3OD22ZATeYP3vMD1X3wAkBcCbewwKp7Y5OPHnqYooNbtdguJdch867Ko
ekGDa+BD8R84Y9px6+YYTR3AJtdXn41/4qK19ydyrlrFCqODk7kpK3UGsxjzaGSqKwVqgQjQl543
3tixksp3HrRFGYQN0RnPXjyh5AfXsgQGMGBdFhzHr7Hucea8hhgLCDi5+9fHP8c6QwfieJAe2BHT
pjxdOnPM/t3EtE7aeew3LfOWTkSqU9qLs4B1hgEUU1xuzZZbkFzu+zfrBZo8B+Ew04Dh9q/nQ1Tp
dIg2Wh8JhSmYGUae7rEt+9g3dpUfc6hbDJivXTk5gZx2xSuK1B2UJZcR1woyq9qxyLo7cMdPmsFi
xsznQPa7Xa3MpDDSdqF/3zBmgUdSCIi/bfS7e6LIpsSsk0JdpcY38a4uoLGSYlxgqg/bHImsrYte
fWtyMMiI4MGAjpWP2PhVhUDEAo2lXg0W8PrPpUNlQBuysBSu+2i2uLdba/G3oQqwLIiXkkKOQik1
Kk4p0+8Bbb7tPcWf0CFlyvvUCVumfqtm27fWZ3EfBBWkraCKN3zuQFJsJGaMBzxeH+YqOeOTmntt
jc7nPYYyIgMWEMXkvOi9xxkm5WSeQMlGpGEpXIw8lHM4P9QK5G06mBelwn4S2Ec+gyhnEHkzydHg
stFuaGgc6XrBY4bq7hZhEG3R3ScXYqkCP3zBmunnBVhLqFW+VhpnMMaWVwwEN8r2xXNwySd14k0y
jOVLDVwHYev/R56xaFK9+YHS5hz4Ixy9PkrJnCUa82apZcvFhcISAqpEPFJTEOXK3llB53iw1nNZ
f/wnNetgawp8n/YIs3DDwWIiu/TGZYbJU/Ax1Iad1pB2wwioWyFsM2/KFRPH5xiwgZTF2SeCOD/y
963GlJwx8kOsnL7owmzegabYjCWDstCJvZ5I/5Ewg6bR80HKCJMu29YdQGmB/nGFmRSv+ZDa6qte
T0IWijfIYvHNExqTAZO4PRiOQJ/7Xj0p59eUMb+V9JcobFRdAS7QXLmZ9YBbOJo9oy9Iaoi9rd3J
9ggtCd6W/o1HVTODeCw4KucoMEHf14e3FL9HhQLj7i/5Tvau1hLDyGS09Ul3TTzTeEx4TENu6RRO
hewYONwoDpzvsGi9zk4g2Swt4Y7hblpXB7jxFsSj30G8wd/gQI73wtsPvfKNDKsAPVeH6KsUsRVy
R+J/CTL75UG8rkSJ932kVUimy97StyjExdqWo5Kx0vupHR5NRihqsjQjnSL4NmavQj+u1k88629S
Pwk+7LwkG3ZqGunOwjWC47SzpawHYfUETrW8mXKzjtGfHAvngku0ChgRR1crlq4/dfhHSROH7nwZ
6tcMi+Er11qQyxXnzgVnReLFS5/eiwUb966vyCvDkAsrZthedZDeNrUw7rtnkBeXBPrvI67Wj6Bt
i5aeHCSy9IzAGw2ltp3mSLrxRH/q36Co5sBVD8BkXFtrdpbGwLJwm1M1TnZ5i6/jjuCJta6NhEQJ
iYIEqsJzGdIRE3ea3XkiteIsUi9nXHMFIY+wOy2PKnTs7l7cuKQ3kZoZ17PfbKleIlgGQzHhn419
5v3uDCCbxj6/L4x1GB+Q43ReY2SrvDpVGkmSqDIpp0TFmcMzjJOK+7y6EdchTzoEn2gYYuu2Ntpq
v8SXKyT1Q7e8FOJ6FtUSiwiOkepINvKVQE+1klTeBxUTpp5oNGKrEsfu2WmJcImUR+IquKVD9p9T
edDNkLMlmZ3OJnQT8wkbLVeiTz6vLBDDojDCV7AdI1IwRDwEpvPsaTwU96fiTHopUncf0QMNy0Ub
Y+vK/O2t/K52XBzGBZdU8wTfKBiyKB0gIkkaEXHz58UTQFiOYitVITdGI3G42r3C2rXnNF6aHdw+
g7qjYXMKhz/8BCBFrwDX+4WdyQSEwWPdEP2GjVXsraCW1KmzXKCjCW32VBqhOsh7GbBmDH8thtyn
w3wJ1as++2w/cd4LpV7J8uMUTjwph9EdE1K5wI49DT1oZcNIr5MEvVabJI4y9GyceM7fY7dA+3Z4
uBgUZLnYaLMfHstN9hPAiWJuzi3FhEyUKnMqNjCd2sbPzzltH2jJzch6iCPzGTy69Mki1XMuT1bX
VOMM5SsRnq9sxwj1VqB+01uWHHgul7I7JnGLkIjlitLVr7/HFksFTdTqgh1mMnzCliB2s51fopgv
UDZ6YivVqauSmr6u8t+Z8ygIptAQuuubdsKf0+ktbe6BIn90GM6wm2I1unSH60milEMtDOKnGyWB
1j92B3BiLB6MDmsJHy+sM2msFMLTY7z/GRgpHj812TCPYLi1AWnA7Sp1o+c1w/Nl15MnV7YVdsGJ
Dj6Mo4fQi7Y67ikm8CneLyPAmdpqPBSF76cyUGDuLx264Cp3nPvIaiFSZ9f8a3OSQn5ZRv4s8G66
QR43CGEzpds+wajHaOtj+anVPwItfxAIXA7HFHqBlDMNdzYzQtoospFUdjlbADqpQ8TsTXj6eB8S
2YV9ZYQWAweba2aqXMtcvQrvnteipVZpXfierG+4dJU5xPrq5tgCmIr8spg8FsVn/zGxiNmKItHC
jgd10uVImVcUIkoZcfb3E8r4OifjGpp8Ppe+jwuore3tw5jTDQ1CZsfCcj7EMafy3nOvO9gjM7gA
qa0wEgEWTu6GKHMXbC8xJ4l/fNHhnTvGVElpAqTjQ36NcD2FSZfroB+fpcAthQGzpEe06fpfhsh2
jXy2HPqnDc5jh646wGk9wTJl81HaSNfpl68hNOaoMugp7xldVjaQA2vA4D/htJarPcdMfZYFnV68
bKf3WpWHf19UKcrftviETAozAb6GK9LNI9k5QK11Hv64pub0Q9Cav+NQD1Tmrl4vHZBuxG7ZeIJR
Eg7cDQcS4Ae86pC3BaDkes7i/D1nYTPnukxfNCewwkvUzzmnyFM3QCqnUA+qe02NHiwfbks6XFba
nsv/8rrS4G35voxb+Pqp/DYuC/anptZaGVqQA4mtxcPWtXDKfi4mPflru1Rvq3R5SXCPHhY2rfjL
lXRDacDOqApXzq/5oIwMD39hK4f+Bd16DmILUogbJP+NL4Cf7rHahpK7nsq0GveFmlgxLkaWwt9M
unb6srHdqn80uRAhdcLpoUeQzEgp1+4U9+X8GSDJ+1ZwBWk+tylrfFMdgc5QK0pV6vBNHQrRxWvD
GN/w9m2s2YTHoCxcD7x9zq6xzpfTDNpbPVs9WgECPBvFhEYYIWJA4WAi7gJ4C+Ks9sBDQe6GQRHn
5gsZlmKvEQQs1qJOK2Ppr1yh4uqBBk+n5alteayDI6kBFPESDjcTe3QYxSxw19StItgyn2WGp5EP
5hikZ4fVH+RpjHdl5VmMvCVjf1NfEJZMhvKpcojr3IpCplCvX3mjgeG3BAANb/djYYhJ+OG+zoN1
baf0m5kQTjptGWQPVutwDxvBxFvuNjQffvdd+ImsDu+vImEDle8IPuFAUABPcbyRtEnhAwStyBxL
M+Z2jPvz76GqULmJNvP3WCD/n9j205bU7FmxYbA43cmO0W093ymWXyEvEVpmNEZ24lK4kq3KeMuU
pOQ3dlG6amv48pnScW33tmMUZ7300M3MNYMfHucyfg31SNOy6lYkcqx4v/63ffWcOFaTZytaPXG6
Q8XYTM79jlBChaA7RMkLhwy4ZoKc0gviQy3Mvx1CagQ7/yGfiQdyaomp3FWWCmfVPYRZsJCeXXgK
4QA2/ABmA2bXNvmjApGfLm67bm8CUWvBcw5mWRPWvfpn9bA7kcf159OT02IOlagwkMybTSnkG0ON
s5vzNAwZ4V9P4GekDNdMLvDD83X4SryocXMkCm6PwaHzQoA2svp29GukigyUXgJrOb6meY2DAzvD
92GboE5SNrm7131i3QlHxvWOqagoS2NWGHRkFpDzRbSFAq6tJ0B9T4OYCPVSA8AzutEIDxovrsjl
tyU+kyuuP28gr0EpHHYEZP0SFu+EcwxkMY3t/t2URGO6o6woJ83SUnJouY5qLJgtNjABkSGtKuik
u3j8/qK5PFzJVKmmAlQ+FmMaziDru79OX9+WEczd9cKyO1AIIELKHSNmpZQnQqya+ZQP9mgBir4i
IygJchcSq08J8Ce13mfmonb87bsloiJrZB9azYfbpMfHL+fm0D5WDD07rOxYrJkY+krRHKG1A7KF
T7MG6XNYW+iRZ8Shvk7SkcnoPJrFC5jZBK99VRfVA7SZGzZuY1FMo0CVo9F0z2bigDMDr3sOddAZ
5u3SXK7t5W/J3EUvyDshXrRzlsQBpXLswYM8AMZT4fytUUa/9fM57SwmiE+92qqp7Avj4PR0aDP/
1YMdRkCYg9lUWE/RoWcbrHnn0sM37hDU1ZEir5wqow1OHXMiUgHeCJqXQdpK2XdPNhHg/EYQcFQB
hja4frBEKGml/OR7ZEKBtDKNTLen+4Mf+zI/ZS8GSeszJjY2eJAfLheiWBwlbSUR+Derd8DoGYHY
cs387q5VHF7J0xQYUoM592qjOmcbXNTZCPYMrNc/KLBUeWkZrJ+p70feXaPkSOZleh1XjDbJ4mnU
YdDZ9C/k17Yq6VTKSrmj1TfuFV0zU+yRkkpuJZQr09tue2RBMDa7YCc/B3E5PbARZ2ThNNrdPpBQ
aXD5qHDnowt4eV/o93WspLaS+CDp2Fha4BdvLKLKYQJXlFoNMZd2Y6g3Slus2zkMKnG8YSqFIiDU
8GSxoZj7RTbNUShukOWJo69ntaYWRI2M7gNKniZq/yWEumZwBbWNQC+mt98fpT4Hca6M4pU7muLK
urnyhSp99tHkyaTfsHiA8vmMXgb6LkNPr2vyPcfGa30dPfEbzdDIX3kbVBUS6bNLef+xw1NvUIbH
3nwYqA3EFXWCj0ew6iOwiVUpF/UWsSmTxHsDQkGE8TJJFNjykeicE9bdZSQZiYLM5z5tkvPmamNG
SplDnvkYpUGTUPBydWmHsTfkDSHFqJjKXcSEwkY/wvgGXQbbUV5rkNsFzHPDGexEdhn6vleaEtX0
DWCWKU6P6hNGFwovrj97Z6gnFuRGq2nVs6Sgnr/5XU3Ljx7dQWI+iKuN6bDfMGaVzAs97ohp+Gr/
ejeMA0VX9TUeBnlghhqmDAEyFI/Mj8R6gUIBJ6jd7d5Kg9uoudaO39x26JwsLg2LW+QKlXUiExbN
k/qrGgH6z+GxnltFTpLW0KvxGMMfPeTBZqoHLUX1EvmvaKotOsPSxGz7cUAW4TP1r7Yz0BUOxdKS
DeqirjVwVyqKVcKKWIjVDlliE8WXItPkMTvX7/yhATnNcvjkrdj5af5TkkAo2R75IqdtJ4KNw5Bp
q3G4ttxY9PG+dFagfKc75P5suWKV3glwRWv8ChSJPmOQ+XxYi+aDo2DSPASHhx1TZBIHme//xx+X
h4A5k2xmmHhHWS1Joug+fiQ1lv5Sy5VQNiFf1jtJAO8smIeIAdtY2c0/0pwBUO0rBTMJ11rSSXyG
OS8f19s10TxqVEKkFUjQhJzU/+ZuLzEKCpraA2fmpdY6kcBQjaFaFoFBUjsbN2d4qdvw6RVZeDKd
mRLBdgfnSFmtbpOYqdJoxQQRVE8TVrvKL1m5w7OlEJ+lvjIcaBK5lKcQnuhvdYYHty6B2gbYP6Zf
5mauXchb9ld4nS0GQ+Gx7jJocNriWDPCEA3bkwRLIvs8VVoTFasMW+q4JkIs4VfhHqBbrbBTDHJ6
rL8jorOEJP6ZnSaPHbWvRi5wejyQrS4IxIdRJWPq/IgiaFLPUbEwBWNa11ZFNp6n7H2yKpD7BxZ5
HZD48jIfjYXKy14kBolztfiQ9Kjv24UplAo+hjIETdgQl/GOLNUuntJm4hEdQ+Y8Z353tA0oqWQn
1BtDEg453R5QxiWpZi1DEQ2wAnm7L5nNjeh7gIDLSvR7LA3ODex2+0fgWqAOWRWrtkzXzeB7AGos
s756ssWZ9I/Xw3bc1Wf5ffFfVaNb6AxQncIAoOYefCdlKe/yyWe6pes4K5excOmvDMv37WBXHOZv
TS5NwLG8BkETgCuN2ZtSH66KLkjuP+BEiSNd+XxTo03gw2fPZtjqDgHm7FNQcMk6C3RpWaKPhd/s
kQt5TTR8RxbDIptPeyoIuKjgaL5lqUENP05XBQ5JBf0qPKNCnG3uiY6jWjDEJnNLFTwzDNlEo2Yq
BMTWiWCHGh9H4s9xRfbTw/XyUKo73e0Yrh11QvZ7VpvPEPo2X1iKazpJG4J7aG9Gana7fB2/lLBn
AjImYL/JqtsWKrLo/ha3TZy4oqo1P8J7PIQGW5Fi2Q0jqg6WGJQz3cs2ye2rIUhLC8dQpAC8IPwH
fnn6FPL6T/JdvTL/Peu/zJxCsnIWEQ7OkgeNgl8dGo0X1bpd0K4vODsKqCpFwreSttoJM1LEGC6u
nDatstP8NJ9+06prEDVqYWgdvW7h7cQdHZV0k1Uo42Rpc/X1n/PDXK+/TgAWA8PIVqrgkdAcDRRy
dpDquchzM/qcKGgF4YspV3QRLeEgapwaOU0ieMqHXw2KW91s7EyjHNWjwiFLlLAYQjUEchnPKrVZ
/0qxLathh8T58c3uy2NqGMb1mZvIe1mi5PjP7Wm8e5j6VVrZ/8FlWGWaKNa/QhFPt5IMCjqGJqYD
vOD6CQwQvb8CcB97iWsLgk6LyIISZ+OxGtrZ//9cAG+cN6zgkLZTsTruXemfOt2OqAnUZZmXgJEt
PL8H9EOdsJpv6PbJRBTJv73xwvKNqZ/jS0P/bfhkm4wn+OLhUYWlQ/2ok+1lXczLUOL8Ys7QKAjy
mugcKaxFXBXVOz0wfasAbPh4251dZHNUHFjavugw6wVnRzu/AVeS19KkdS4TXG9czS46QfotDSxM
E8Rib44IJD5yAPMMcdDcYcaio38Yw2UpXdMSynQiDr43DJXFRD7ucrIDs4LmK/ThuF0WloM/CAff
YA6vb4HDvYlDXONaO2XM5svOJl7h0dSzsY6i9JG070SIP1+9fdcCrU1SOrmBlFaijsKvyItdbONF
VGu0eXDI0nZ0Nkxd/sV57OwYkWW8CwkQ68prmBLScn/fZJ072TwhJOdRw4ypmpIOJTwU+Cs7gk7A
AKBAdMi/Kw82pbZBASAPSLiooxslUfSjiGDXGvQLcMyY9Fipwqhum9naipEiIEq9PGetKfJjBJBx
U7qL3tfHPgc1HNS+A2INlwvyqL573Ci/aomNDSeXfQZ9jHet4IL7OPnRK07GdWf3dosf9kSF/Okc
2+ZIlD+9bLKboUvd85ahPoH1Yv54RIEWJGfiB/bWwVWJfZEhOyQ/sZPlYjy5+6TOP6oIIfYWu904
50zIPfvHm3D//L9s+C5QWw24cte6Mw+/LFZ41Gntmh7OGzoIXtLZtoKE6ExkCvZq4CrHL2D6Qke6
l1v91G+boMiI0vK5F+5BVv0LOVNm/EP/oLYdAKjvSwJ7cAZpJbFvQ4UXHm/GICyofat/LTXtqe9v
1M/QG8X0SJDyGt1smbiNaqdtT94ou9F95I/73oxDgYknU6n3X4kLPBkFmAjXFphDiISpIRcPYArV
T0v/JRCvJEjLa8LK8mSxF2B1RIMSxMpq3MlINn3SvMwaqz5pJ8OAs9pGXr8on8Ec1hIsbxTO+hnt
oXOv29Uk9fFnuvXED7NBaquVBCCtgwr0qstLnni49gLOvt/E0F+pLdGFUCXRRqYv/7RmtB4/2vYY
/8angC2jOPyVJx1bFN4yInR7rsblaw39QeiRitqEUMtCg1nQUmuDyp2ImBIVu/AxLy4Yh73nU10Z
gGGvQdMXa+nBOm+a/Q5U55cqAwDU8NXy7+hNZKTjHeef7wMXzdhfdiUQR2iHKbV0zj73KV9JIAc0
o+is7T9yPcL8m7rLC6Jjp4S0cOA/btYdaymxYlQMx0VK2Rb0ka6jYiF6J1HsbRuUpX9A1Quer0N7
ZWIFsdZG8mLZOjggKH7/2aCAP0nn383/4MX0DnvFKMmH/HqOItWm9aJqxbm+MSPGaxMuxfPT/yMu
pzXJ5kI1wy8h44omwNVzLjp9BOzUdXXxFN4A+MJ/0YLqwWRS9VU8yaau/V5UXLkQOBZa7TS7mg5D
3u2uEDw0PsenEg35HjLGBTsxYBSBeWjoxfUroq3yyO93R+RlPlqX+1HwKtAZCOKaeZtqKIGnaY0S
2G/izM4OMTvEsKLAxw2/w0gJ6BMXLpsbEy+OfKqU4mi1/frsK9l+ptKSVibdhETC92AlNtV4Xvxh
NdX18G0GmduY1NSbBgrj4evryqILLSRzzqqUPtnUXKY0i5QnOdMN84CPqJCoie7VFJZ3JwrSSaOj
emG64tsbQ3SqPda3robI3gC0XKRsOIMHCu1tRtY+SUd4oBwh/kMeXI5h+E4cSYS5RkKxM/7tdNd2
kWd3aIf6J7jvUcNm+ItBZVKv9Gt1IVFnjxAgmjfTRaAGS78GZeZHApkKXM2x5cvJd3H5suqdFz28
Inazk3gkjzgFJQcEabTY8kLXeARnIffc8XEJxmOjAIad4GOQIeRGtP9d81ucuBXD3Fs0UP7e5cu5
LKbno+80yMf3evYhxxIZzGvSQwKHNhAMcSEbH0BYmVHIN65jfLlNh5HyhMoNOPpxT9+tZ2/RRELN
Me6KFaKHxzCFf3URWFI6co8dkwhk3LImP4CZ4J4yel40lR45sK0NIBv1809Lm2xRn5LFXIYHQDa8
pYJkVmuDtjJbBaFna5MOxAtd8yw+BV3XV9HaUnMdd4pvGL4oC4193cqDd2agOI1TusrGpl0x71sS
ysBbMt4Y99C+BH2OyLUbHuKSIKs+Se2i4dUXQi8NS3H40OlBRQBrwPNum+G72usKyf96geAX1S/3
KGtHe4RDPj9N+2o2M6KNijZYIBMG1Eje8btDFnOc1SR7SA3pMAUu2CO5yFMssL7eOtLd4uTWKXG1
tl2N/KFHijnpVHhhJYQrYZIiaijamrcJrPIAFyxi9Bxfg/Vs10xX5t5hwcliTk9rEzejULdchO8B
vmyeArWYri/j1ljNi8JShaKDefPtytpFIjVh7A8xDlqihOQ8eBfr4QFGgFvmh369YouLx1n61rk/
4piu+3roex/P/ryNYvKG1Ct97XNQq/UE20jrRskSQLi9ZRD7IZV17xPkFPMiSQX+klYXU5Jiaot5
15uQTJKLR+HNic1iie/Vtt7bU9kceWml13fb4bYBz9385k0Lhou8DYJiiJDpo3SnRChAq6vhg3Ak
4+WoqMoGIMHNspnMb+kqvyaotRTw/03UlJrlfYOjaqBP2nMPBf6nxVyzWJGriehgMwnVgFLgy+IG
tipM4jQf9IHQT4+H73BfjlvYXfJr8jmqXIHzQAXaQNlMB2ou0aMg5NTV9XDWzvLPS6aYom/I+nuL
7CNutPYiCy+owH4ptJG+efTTMunnKuH9INa6B7gaGPcLhaC4tayuxrcL+QENDHPyA2wOTZogznhY
UXkmURywbPNXYOoOvfBaAmDpPaVkeKGWAtpS6Xga3U2tiUVQXuMtiIMJ2ehJA/VNaY3RxwLkRVEF
eQYlI78eCIRLSdGSOCSjXttx6+6rrqJdjb7ioJ4NDt3KWtcfS7NEwt1XdlL8cwaWkqIPQZqCM9gk
gyNYn63J6i0q5jnylFhJO/3yLoCLsvx8kfD9kO/+AL6LvNQOcq6z3CzsO1rWNmsZCRVBBXkJgEVU
qZd85kGI9K3BbpQkELLG+RQchCxlb11HCGdWNG1DLh8GAYbhtLXkciHyp4GTeYF9IeJwRAGmLqF/
UV2sZccWwWbLOJ2pscus7zpEFaDSRrmWxTJ8E3Z2ULK8XsFoIyz2OsGNoCkNrFux5bfmqEUb/6mx
QP9kyLQTEe7TueCckqsoubhJ1sMEa07AH8Cxpbq2rizTQB4kdT48lqJAWTftTDSfty4E6pm/Cav/
/dKSBm1u2jMgiNeXgp1oeNE4HOPFMrKSMiwCMmDcvpj9zayXvHpOGfkfPLVPi5dMO7adO2CR4SZO
TIyCKALcCa+kXLxXrbH3LqJGQiYiyF9Sqjctj4m6W+m6fpR1gCz4wiAtcVBJweQOy12xhXVuk6sc
Zh1+g9N9Ye9mESlw/66XDSTCykXxMw7J+B6N/Dmv7Dt+HRDSLpC9Y1Xeiu4TQxBuO1FhHaR3QgLp
eWhvvJ1ztESmg5smcfACHCrTdxm3m3gIu1GUIOrzbep+l5n+vnsI5T3/xuTISevzo1A7eaTNA0sP
l7HBEuCKr5Ny1EJ3pMBP4kMJPmqQO8s66i1X6na+JL6B4Mdyr4PGmPYq0hbRydrQixQmlS7jEi++
vrHNHHozAQpC7IzKTNtPK/KbLoelzAbGagb2agCj4njdsqWRhrYtBdNORiVJwGBs4w+noq31JjGA
ZpgyIVe0A9Yde4igXqpbKq4qpXynthy3mjA8biYIPto+xG2up4xN/wVcSE0KQbv9JJ3VXBGObTXw
PlBm/mRx+hQDBSeX1p0SlGM013dMtEIaEGY64X/jwoef/48JNR1ATNrX1j3hpdRlMFkF7XxttRdX
UwI7+hRHa7NQkaeGYbmG95KcvFFyIfttE0WBHwMZ2tC/KaaF971u0TcB3TIjIkH+DHNB3nRatVRx
csyVSHTHjocB2yED/6suONUn5qS8a+BCVTD07vJMqdZqjgqidulr8gRaMuxuuyyMnV8EcGB9xF+k
+E/sWJkCY/sqpWXi8YpqZnL8rfxgUs7P02ICOmqgR6O8a1GrI5udO41NqzIRk77xvrwXwnmMOJFe
j32RvjS6O28RgB44WXjM/UA/p7lioUj7sMUIHUS4hHQCJ4/7JMC/KpkM49cBB42V9F5BGefgg1TH
MtKLJ1yfHandTGKwvztO49HZMXnk5KA5T8id53vaY3hd3AncImTnoi5KyQFwhP7ljWnFYj3jXMRy
res34tchRNCBBvWrdSPPbZmjUrgBtDTK4ku5r74mWQJVBaLFtAZZ3fHpiMYQUlTURLftVoqz3/fj
0FtYIttmPPMNQ2MGaYfjEBCQmmBofzCd+bR2KiXM7bzE6NwDJKlhz5OPXf2x4yY/32aU6EOZ/6Ig
T5hKlBaAFao6x0iDsczN1tUK3ejWSd6e/QEcMIb8IRm8qaXwGaj8Hb5qPHMaLB7Q31HU0zRY7Jw/
v3Ei0en2y3g9rK00wDgQRnN+Wv53t6UjdD5LokE3Z5OIYn3Wm6SLiUEt1AiVkjOwjCqwQEOfaod8
4y+PQnhdHH9wQdEp+Xi5sTjjJ3r4EgHbTv/RMCj0u+l3izk9w4qhbGybHkOnOmY6x7pF7jLdPJkf
LnHM8BjErlFiLf0NpBelCDtMatnW2dm9+X5tMG/AYZs8khFEG2ovB9V5BiDi5zAZcw2HNuDxbWVi
etFKR+KxVZ5tyV55lD/lWSfmt0yD+HdchKyUka1JDAewKc+1jLf4teOtKpuWrR65eyU59RU2RmCH
bsWzvpsWjWkZc8MoBWzSupXAiSDCXJSc7mYZ5i9gnx0s6waEwTFX+psD+I4QQy465IIe0zMeZtSL
ngqQ3uTY3Lcno9SEu+UU7WTuHYViIAUO4ASWv6w0bxaz0m4Dj7cYK1A/Kc3pmsZmskqHRaus8nRy
CjX+LyXehlu2JHkWKaDeJFywAnR8Yycvtd0LCFFcVG2I9CCSBk6FOqtsrA6M/A8Q9cHjxwqIrpep
DwL+SyksKOOePN3VrMW9cH27ZizseJrbqX/JHcZ1rG3vijWCqynb7RmiVhHvp1pP1bWisfRIPEJP
fJK7INl60VBBCxCSXhzWZ1aNtBYp0EJX22gjtEbrU7Aobx30zZjy8tTg49H3i41mT4jPGHrmbuU8
4ZtGwAKllwjZA0PiZgiojhsBs5cAZhu/OM/d/VB3fJ6yxigUjnl/mtUONtfx13AK3AnSTClBVRdg
4UrDlqomCRH7iy2YTqukFmQo2GABibYcCgT9Mt7QXdBtCXRXnxD8Aw1N6eiVfzHnJUuopdHBLGGg
5TS7EPvm9ZKnkn1wa06Yi3IiHx03KBYnFalSfD3p4VhWggDMfp+GongS5wueMY4CUf6LrYisYnUH
vNchygPRH550T4lN/wcY55pSdaQMzZvXkMjhHHF0L+b5eSg+b5OxwRM/HDiT7AMQZd3yVx2JzOUA
OY5BVcdhibZevqH+SUVoDWGdtGuLyPYsSb5PFuw1kAo693mk/LEPgRhm9OY9MTwaDu2hVi6UG2D4
5Gvu2YUB0wXjihnNIpxVFwEhroEZieTJ2Xqb9hheMVJYLvujNAbqkKXTewUbPcm34JJYTPGZgkl9
k5/uj2NVKvsUJ322UDG3NRszMXxOSnipovfUJRXByjnIl6fLaE/RwAgtNo76/bRevT6tMb+itJ4x
13A+Yw7T0EFaD1+w6QprQzwGqN+VHhifwt1DBuhKZAvBbu3eDdsj6JNHyBeOZFudvipajGNP1xZ/
JIkqR8tp2O0p7s/SACj2mtObyq94HqJVAaGoMqnt6ejaqrLyqv8uly6uZ7ZEoBmfLBvrwzA4uPrS
tRDbHFI6KwhcqYixqldgWBgNbXJJlfvjKlB/0Na7BCADMKQar3r/lnlIOgci5WEcKps9i41Euf8X
ukXieIMabzM58Yts24lryeLJt2eEqLVLaza2uVJ8ILX8avzNUzZ+QyBqNT3K1b6MLZPmUsQhGhY3
Z6g8uQiz1moo0JhMGTpX32gqzxRELPgZbmcfQDrR6O7MTw/ZDwcR/CwiibqWZmbKZBXBVHjlc13g
SnR5Ru1Wj8SAg4s+F1DkVDjc9GbxNILCQhStQDJj8VZIIfcDvm0fyrjp6RRDUkZdFDI0epIUzRMa
V969qcL1cGXNnFXnBueIMJ7lcOGjQ9SshjbHpcNZbzIRtIY1Ym2bELZIr4PwCW8K50WZGduFEywU
EGxtUDw5kNM7KECbhZTSsR+h57O/gz+R1c5Yv7TDsOL3rfveJ9JEYg0W5FlS5Lp9T3FwQmfost4I
NjyYPl9OIeDMozRqnqiugN8JfijzJY3lSxo9LI5geK4Q6UFqZt8x01Rzr5Ec0nBMYTn/KT75UqS4
1hh/SIQcFWavlG5CNqpSOzl4L3nvznGmC0ubamaPUyTgL0GZKMmD1fJ0ojI5eDBVI7l/ko6mzkRo
hJ20fCv33n2t+6tqbZvz2nIQao5NT3bdjwD6u8lRxBHYk5LXLRoS7i5r51iYt4W1qxVJ0wtlbjp4
vQ2eeBQqI7QKLwAAcrvnRZ303UO6W1RyaHdnOyADE0//OjO+DUiHXALuxn9DyERUmLqqGOM0zMgC
H43yvRHiOVhvSQ+0v8MqD6IF3EbuWAYQH+2pS1g/RImTIWyHvgzqHv4yPVP5HGhRewarttSF7G3x
x+5DXmC57M2ZBwtx9DGBJGEBEnRE42FhdNOHsJUm1AKiqZN/Q9dQCHJPnekI/4pKb1JQQdA3qO+t
69I9XN0yZ2Gw+BVlzAvYb53LGzRFByzx+4zC9Xe68AHc4DwwtPzqwpAKsOQ2zRluB2rkv0Hp5Car
kzGZJdcRKAcito/sSbfivbi2UUSSH7225tB9D2u2691qTcGfCAR8wS0O0OOPDPwYn5VtJ7XbsDbl
keFJ1XzI09t1uHpBdg5w597sM80If/v22oJvxTfwoRJc/800PO24dYwKuBS+23l54qRYbrYv/ezQ
MPEjElEVtIrikjO+9zAwrm8X/b+KZr6Wk6pDzlnxFQjxp6smAPyGvwDcANNxctF20EndCpGGQZSQ
EGKOk2gIpiZG5WWanks1w6vtPYWUvhRuqazY06Xy6cDl6qt0Ntr4qt//bMzPBw+o+BZJ/BdLwdNr
Bkqou6LGpL+Imyarxj6cMDeS7IT90ZoyUtJXc2IpRV0dO5/PDONx0/uoIX3CW6B5vO9Sv2Dn07gX
P63jDSoftcLct8ZLcwTxwCKZfzNnJMwKiPkSIdb5HdlyJzxJT7LRMR8oUmTOAHgk8irCDNlaZavI
T3ef+uM2/pbTa7YUwvPYlb/Xom1mc0fzOOIo+d7TtZrBcY8vZWLq+in9JwhPkV7Nyn9vdUX8q6SN
X/Go6USvXWCBt7/9CUH27k/Ql2zJElbrSNJO4778pjsISUc6fjqyyYoferdpYnJPutHIHJ9PgCzn
z8bn3ctLBOQvFE9C10E1Y6g78BXeQLNJi1x5h42pp8akFQjoixWwzrlsObV4zwd+CZESFha/WrKa
dq/iM961ytgOduEWLJpfA7NIJ/ssKhEC2vff+Zwi39pHf7MsJjeIgJFtUr8Xbmdgsg9bVxHU7YsG
oFKu8dwpAh2zHlxKcJCborw+mBjLDNXOdXzm9lQN8GSSvSINExjRzJz0c2vlDIZfO1yZipgxmjg+
XvsObp23c+DVuatMbBN5QFILary/o3/Cbgul1Ge7O8lgFSJmMO4rF6tUw/bAbevBUzV2id+q06d9
uhAyYDmSsIkcPdU2iitY3Mj/JZ1Cwn9zZSQ8aYieWRF5ni5FDlKADcbmBI3jakTdN7hyQrgSbaqy
3/Geb/7IOWdamokSanAeyJwTOGEvjfLUYvzBCwZKmt1O5EQP0hxIT5Em4XK92Sd2YZvj9ut1znYJ
5YHTPa1WC1NVQkbuP9JHqEULbYkKSWg49Hz9ezwwjEMBBbyzVZ3vD9jOSZolYaGt/iCvpesR+XIk
j9oq3T0gOodRtxu0uhWY1fqA6Bfwd7HcoCkjhH/O3lJWzXzSa10jLmltDouZdk01ehiRVfFc3H9e
Eex9OIaclbji2g89PT2iG0XG65uyELQEBojYCEouZWJMRu/Tanydbkia4W8AsejhB/v7MF1nj4W4
CJJtRLGyKkZ72yo6afOMv4qhHtsVkysPOEEUQ1eEUFdCGILQEAMrJPD2llEe761H/C5uJQj5qbSG
kOuM8z0J0XC/kTl+HaLxPBEPq92/f4jZEWMWW6+ib3zlouVKJ6hu0AWK+a7PoTnPgOBMaYmHV7cq
Ae3C/cAfZgtRvyVl339iTCCzbQbT0R/qIux7BJWpuvCQMqnu5fE2NI3yxKMLmnm7y+SByT/E59y6
+15QqxehLyqL8c3GEpBXPwg1NJrkv/DjoDwENhChf7aUwLucBEiXxXJfJQPqvIycTkqlA9cJihJK
38ZNMcGeZU8q0hYGaXHTIYLcU7ezmbwacAfQ6vX/uYMipq6DcBFtHOpm+3/eFKSS4XQFGrbWnCST
LD70RGJcoWVEjG18VOq4GQaQSpvS7Io+TXDJaa672GwnYLqHN60e6wmkL+lC4h7EyjF02apAJZSR
5SjVNnn3jHSB93VXib84/wg+huCmNI7gQcdiwlO64J+eC7MK4M1j22ZjMCN98zYnhqWYI0Om1y0Z
7DK9Aq7NSLqfc9qYkk4O62cAJGX8wJGd8SKqaMTe+cTHe+2SA5cxLhLWHV1LwLuU1zjLpgLcMha0
ZghFyf94HubKTUaOJQ81gWvqO6Xtd0cjw3s3wMDWxAPyrcvuAKFWXnmQEsOv4zQKzzCCPs3WN7TQ
z/OZCanbmz+DHLYsL/J8Uawh4X/63ZnZmzkxZqn5S/tIRZDEQPZDAhC89BPYialR4DCxSIMfjW6X
yjOhh0p5kkUamlyu9vTK9ewuJ6L/HwXqhMSwH8kcC1lvHXZdJPPyQcN2U+Z4HhZxseFTtBulDFjn
GS2CjLfmIt5ca825sa7OUt+k4QDctB4zr5szV/mDnqhuYf7y6puPpEikOxuzZ7E72NRa1+yh4YXF
DizACcZZ8AQeG3x6zU3DnFeqlNVvx2i3ngwv9PEkoMECaI8VBmTWjf9hNhEPUXBFbpTvC3iMpK4O
uyvz9MYChsEoeJnXvza9yw6CStCTI2gHyBUeXTC18yDkVETxJwuf6p6pfIhC+TluKJfz79ey1/rr
KL+mokusYvsLZH/N8wmf7aNgF0YDz4YPpG0QEaiiG9ZgFHL2SswQbEch0LuicazpurV0vG0OOY18
7bxuuaZL0UgAU+jQKKEeYxkF83kpoNV6HIeSazpJTDfnrDVeW5FvRX2cDzyq8zK1Mbb9sNDN5q5F
BSh0EmYGhD/y3a003skrX6nV4ZrEyIZPvDll812sbEnQZ1lzCA0bixKDRZwCKM56o4zNVBtd59qe
GaBKxK+hhDRbKNsii9oA06lUni8e67+YYbK65HirOF6Xw6JxQo2fu3r0XKScsAO6XzGxjcrdMUI0
9QG4UJbdgfZpO4S/FRNo6uGwg+sjMbQuog4RYKfDe6St4G9F9nN6sbNZnpUcgLQF8/C7mOSk4Bxz
maMFRZyB5GsBp53eFCcWE+P7QKEBVeEFPmjI6qCbwvLATB6sfRwH1T0fHOgfha2x421I5SKTn91/
4yhccQ6a2Wq32gZJN9eWOalg1C9gDNw8NMPM3UJLu0uhCiyelXNZmZ5PA+xaJuoI7Z5OkKkpubFK
MOMxLoMDGfTiC5gIZ3d1KD18uu3fSUciaje7AEPxuIe3rnFGfSx8JOxa0gibDMeuLrzs5J7uDL8b
h3x3F2dDUEjVA0YT+oD+F8TYQq89Ml4dRhbNfH4NqeU1iEXpDlwQSnSwerPyccLE5vq7pzNM3slT
lbxjM+ikQuUh/Bk6+7gsvwHrrIkRn0vwD4ZwfboyfG8bldtA8EuP5JTF+vUhvZ0bqPQP3O6jf4rJ
Sv4g3Pwz02WoOMVeZvdDXc8oSt+X8ZFyUv6JSZbOOGnBvwAqYDJ5XSChte6R59B8jX0Q4PeHMcQA
NWy3UXHBy2oEeDun9VdZfCUINKDWdB7xV+ViAgDKXtjCiI/h6cM8+Mg6XHiP9aRnlRLQ/+/Je+F8
K5GkX921zPbkJIyJtXb4GJL0KbSNtYpbdJ+k6lbFtkExGdkvoM8r6U+ejkzWHMBHzg/Ix6F37J97
owhX+LSw6HoqCkfYNbddQRHFbufU8Wngl541sFciv7A+GWKjOWx/+/H9sHiMrfCzH3ClP/FKULP/
Ul1JpvoevFF0zSvECOOvaMRsIE+jnMQGk9hfO9Jt3aYd2LQmxg9UJRKSg8NU2mQUSY57g4TwZgB/
h+xVL0ZJuBufrNEF/T9jMVRvyGhHgTb35L9jS+NiZq+jtE4TVxbDXgLfqXLu+Mmas4xnm7OdfSvu
yVGZ+nvJfXAwcCBlxfV7zPjyLWU2lqry2bzS7U8F0ylNnVC2/pzEnyadoVk8bFhdyawly7o1QGrf
B2vfeTD980gSgd+pob0tjkVOMyuWunDm5Jyy2isXYLJfEuEIu6JW4L05ZScYUps05hY6nctRti63
/n4HdHIu6msH1w/+1Xp0NgTIv5NGjZqI+1SMIg6loqTjPBNUbT15puvDupIGNqQ+5Rn26kkOI0Pu
wnnmhuMDiKfch5T7JJ4ZWQhu5COgKLlWeMLpmAE5ns1K5P8WbyRuEb05SrSjKm6EjycgFFlLYLrB
OVDxbHQPFw3zQQmU51nBV2s9NaoUBG3KYCYQAoMNnup+1Gf7oV4vdIM5Lpo6sQzLuvwlntkOjhJ4
BZ8T4GL8cF7yZXNPxdhpGAIETtAsbXoFqpp1tc9D/6A+/euk9kSY50EjZlL7wN9nIJbtQ0NrdIOR
0eBj2T6Y8tOTQLK8+qQL5UvA+e9BZrVQmV13mI06OVT+Wa4mOs7mXp4CfZ5uwL6hPqh5A3DBLhai
SN3EQGaEjb+7lun4YJA74qtUajWcOoYw4TJM+c/b6OP0LmROkeTzrN8tTrQpNHKrRydZ4Vi6CGVC
dRKrm14pfPV2pgWWqx9p+fWkGhCv1sNhaPLTm59xZyCTFAzOYjowE+dX2lLCbNRlQfpX7PbflUkN
CZ1AJh3pbvs03cS/xIAeuTnTG8H7sdF9oGEmgwhBasZhEIxi72baMAxqTj8MBAIGSilURcOLRRF6
inR5L22dQJH2vhCNDVCMulkXQM1+F2jTVzNBjA41vBFwde073ayXfJ2nSB7kiKqNZ/htHy+3/fgU
i1UyawExeHknKKxGCJWNfVIO6s31eHwuUumBv0cB8T8ALymeIM8TFlhPOzjlXhp8dXao9vdR6Lry
Gap7JzRLJvUpRKxZaMn3mdG3ch0XzHYQXAMS4TTOOOZhg3pkIXmnCW007wRODsklErD3Zh/EPpns
SzOod95LzJgC8s8ts5jg0rX70mDagj029dO5bZgUr87L1QWl2MBdBDy+wX51HUWlWN2ThlqPH01g
xZu1RPQpttdxfEi5duj+WYiIwt6ueKmsXNM2iQ0jT7D4k1NZko7nRzzJetYskczJ88/kOu7QEMLo
GclahPLC+3vKr04+8CXWjIf+xzHWGw4pbtag8L+lhR6DbTkTspYFG4VLSZB9quA3GCG/8hEnHxxf
WPCv7thf3BndfQj1ryh5JFyL5P3khK9s0/n6eYVZR9lcAaFOZ89xGtTyUzlAriDuHKpGGZSR+bva
DAYphjdcMr1zFbK0ZaerAG4L+f/JdkgIPVuwmz891vCiknTcpeZrwPAoSul50Kzje0xD259yAoBf
1D7SBG9CEr1HEoGIUHsPBV4mr4O0AdcxQGOcnBFJAsDxUAyqGGLyaX52pm5Y3P8POfK11q6qDtnU
iUn9p2f3PL8znv9apyk430QQR5hlYPY0KkjEl2Vm0id2QwMU7LsXMRhQ9DdfGWVNidW6Jvgy4haq
Zb/SQx8blvIpUr4rTPWQFGIZQWXapcXMhCtshIZbuttFiKSw7sQg59nRQtT6Pgu2sV2yjWAWw26X
lQwjjj5MqvOl/zaDCoVBiNl1HG3XQdMSK2SjMTbBWsRJy8AYjF55PAZq1vHteHni9OkTelA49Zya
3puQBxK0zNurCFND/o9mmNzkO85cFUs084DXlW0XLKg3Zw0MbRbek2Bfa+YIMh7vnnaejvXGh7AP
BAB9RN2mgD5oclDLmGel3iMw3mvkGQ7vABBTG46nSSKdaVDPBqf7L5/EkQ4a9/7KFG3aJgOxzor1
cZoc9XN8RVW4QVZ/dJMeDx0k5vbwKO/XAR8Ff85O469PFiX3eif/x2ZmthIsavyaU8iBN/XKdDoT
4OZ8Z6KIFhmcoaypHDttu2DQCYYjaDS6EHIZXmIyueA2cExgELB9lyM3RLELPswOnCQg+/ZJV+Ds
26gTo7OHO0eS2IYUR+TdclrEdrBPzzPiy9uTeZ85BDyR1coXutZm30c5Otj+CvBmUf56KoaowT+6
spmANY3v1+gGggUKqmbLGrTzVbpY3JrcXJPPNNU+h3Ug7ngeclWTj7M5fRmMDe07EmqhLqnsT02Y
ws9BjW7wa0pcwET0S6rJXNSGg75jTffquFlCthtx3/cP3QWEuUmcTiHuISq2HhFwW+LxZdojoIFa
o3MGZIUVjV2FaaJJGseqq1E0xXCrFEunf+fxKNDg50pqIcfGWzBJFK3DE+Sa5dVwrlyeUdP8rZLc
0otN1QeQbAbru4j5IwF9FT9EqgJpvfFL+v9UQvyohLj/QPqAVC6mfdXgDsTr445cEwrt9q2wZ5iU
roMOcYao90Ic0c/RFzjs0LuvGa2ntVp5xUiFmp3gEUtfw8d7VhtTS/6XugS0UQEB27YET+sV/5iY
alyC2tcxigH73miYF52AP9gzF+jz5fn0TvLe1XhSJ3NAHaQz6ZFMRGTP0lpU7/F4WVVdbInfPJS/
9ubIdhyHbxDl8rQRMbanNYP0RFT2zOWkmxV3dqimWkeZTcuY4J182nfNNBQLGtkWpDQGlZpO1Uk5
0QGPbcAglNYyMAzvrY0P0lfFfg0x2VbtBUIEfvVwr5jU3PU305ws01fsi9mlfaiYCDLV6b5E9rrB
dvbhtyY5C6r22777s09e9VTp0K3lWhbuukfqM0kTpAw3eznQCZmKuBPyBYwPGuz3qaPr1UdXhYzi
GroxVn6xIti+8yrOsNqtsdvbT/a57dviK+Ulyq8x8QW9ZN/WNHXdq10A9atwuDjEdvYmXmWaI0wB
sCd5wNeTzbA8GaCJBdg+DB02LNcZZdv3s45o2GzWUcOgqWgajcwhRESnVnxS1P5UPKM6g4C+oL0o
uvnzG+FyhbEh/rRgh5FuEtogZIpTt/CtsmvlTXadEukdDEsFmRMTvp8dDGhDnvQOVBZomq2ZB2Bh
FdENB5YK4c4cZUNDMK9ZsXTT8h56J7/XPwy8eTTQOYhJoESnn7p9alnYNPYx5SmiB7GHKj+JSJWi
b6ytk4zV1xyODnG1kmBmFjOuS1aCTPJZ7gg6WYJGKSAMruK2io4Qfl6WLEEYLlN3sI+QCh8y3Z0y
ilewiG8ctc4zEkq2c+CAT6FW7B1zBVu1Kk4jp4CJ4r/txHZ4Wxwe42BXv67jg902HiDNhyzKJJH/
30M+t6V55qET6w7ksWgNDM62AIeJkp/DCqL0pIp9viVxaASPK4oEzfalPOqqmUJuuyqOGX+hk6IK
LulhIFMcsHHcjF74A9oqCekwDU+1LXVA1e4+vRducTfODDBgagP7suF251PBTPaQDQfzfazqCI6a
BAgTtP79o2YZq9gfndPJ2rkm7vD3l3Frt/uzPZWBItiIHehfkTx0NcuY8j9/DpryAVLAoUn8qix/
nQhtoIYTV4hZjYT0xrp7mu2GAPpBoGFFph5gOHyqDfRZSscatqCwhy8QMg8Q6gnmA5HEzk+czZZF
g/9PC7vEQjkWnxg+lTmO+/7Tux3cFv4fwx5Xee0ma11XhMhFpw8OWUlDhFa79Ezu4hrY2ux4M2dG
oIQ7ydM2LCypzXFOAMrAXL7FPalnM/EYIa96vvD3mVY/++UgidV49zUACABEwToLRCPSJ7U8tjtZ
L1sicSEPLMC7eIn7i7u8lNY5/0NR19P6fgdQqAIaSOtKhHYVnBH9EI7e5Ns8UIIsoVCrPHdW1Eoy
kB9OkMtmYmWLyl7yjUb9NFVY0Z3DEiS5aMpUNEcTtVsPA9516BqRWG0CZbCBWzWaSvU+KDnwqNH/
S385U7+mqQqpas8AFKahHokkjEYLQPUMVXzWQ+MQedtw9eK3UXuvAQ2/VRfIdqIEg4hExBfLZenz
5Fe9YxG3Lsh+Y3eMhKVnHztBw8zY7upGBT8IfEP/8OHEOeq1+LixXCXyUJNKsksEQwkKRYUVSvf4
aDoR6N56owzb9E4g8qzBVpBrhHkjQiG/0Uwjnttro0EUUZtcC6R9qYHqIkhGgQkG5CSFRJ5xvQJl
HD8ZleQXGgu0fPUBefsYIIrt12UDeVODpiHhe3Q6eL1tvadY/0VpwNmpUpBe4dX7ONWWWqcCnHHk
L49c07UL4cOzGhJ0DdedY+jthuxgiXk8u/kcePkq+J7+DDrzEj1YHPy/DemF1lQ0cipMGg14M08s
vjkW3UiEkH26vbvSex04fgHthSfSClW9kZ0a31pGOvPnHZnJrP01t4f0XmTfSoPc7BP2SiWa0o04
8FtsDT37g27h24SinS0KNrfocN1zfV3vKgC8tqAaau457aMQehXcT650nkSd9U4RkKygKhjXMlsj
5IGvHOVlO178YfJFTpq186h1NDl+hF6vX+gAQX0OgjKco0Q73ib+xQyoo8xuvZDUjZJ16ch7j4Rc
PcROKbax85Ony7O/txnu9YKvkHRrQkf61VnnA9FfoXy3E9SOZF8ZVnNCIHLlWDVDPpyviEQAMtFn
Dm+ANk9N2tRESEKmAtIdLELl4P5AkvFqtDKhdQzcHnoBZQ64GpgkWeK3NueG1tCtvTbKYyVUgxQ8
DMfxMQ86pepfMJ9rBX5OrFAi/BtV9Sbwy9pHYEc1PbUYm2kVnlmsv2O0GmRwtZRgePi0AQkS62Kz
/CLUtpc0aE9L0Is+0+a5jDW79uklLDpy8pNBwqUbRJ4yX5vPOU3zl8HKIbSPrYfd8tybSkS+GoBu
Ku6LML08koMU/3r/bDTHH8oLjAQxLwwFhnPWYtl2D7zxX/dr70EYFwdNEYEMvu2yXj0tHT1/9k0V
gqN4d8qN/lWtjXuDP6tN/YORXmJpr0J+BTc2lBq4xagdos2NpMomN9ybUcKkzNfXwDJdZW/Q6i+N
ae70sOD85UR+BcwcnkMEAr8cVsiUrTci59yA7rysoqaEUZ7M6fN38og4sv1Hjgr/7yQd6h8nbogB
9qi7NxCUVeRr4qRJeWFAeYksm5+xn1PRCiGRzJ8Y1YlNyEe6B1+mVJ/VBqV9LhbMqlpzrByASMyA
1JmgWXQak3YFHVRjyGP3JWGlgotiK33YbogacS60L9HTCs9aKBibvbYK6OpwDSz1pBc53iW1s1RZ
niZaLXaBqXtzBxvYQ9zaxyueaPkowV5R1q7hOwM7jCdaN/88w05EAax+xlldnFkV1+djOjcGHerl
AprkDzwB1R5sGs6ZPjUbaneNz4OGPQR965qCKoNgFA4ObpjMZggqH7pOHjH3ZCHNS8Y3O7MWhrEu
vL0ydJWJ16rtkJ25/NrC8OBKCF3WIvnCJ2BWuMbeQVrWtasP97hx+F9V4K8DwtzIp9fH0/9dsZ9Y
dlrEdYo/F+h4pCpFQ3jwrtAhmR0zwgutwCdwhwhKhw0se5fntUke4hCLYL7Psa6kpBunvA8565Ta
cOXcIn2/W600eMzN2LZuDGI0rrA66dRlF5PjISPnZqvs+/cf802wXRFxGN2Ei7Ayzic74oAsZ9ob
U02f4fZt0XLXo9svbh3y9rAPTWtAbXwdg/ADmA8lUSdCMV5jMvr5sNbruEZZl1yEqEmQM1QMk6qX
R/rC1Yn3iNlJNCSy+nTMboRpp8yg9LWwoAE/+m/CEwWE7ww8RBoziLYTKMqSZFUr1Y9aaoNsghbl
cib6egccPlAB8S0fyb74klVH9ocOzu6OOL74Pb9bvLasFHzTXExTiDvfd+8MdvR9XZB2arRB5Jqw
2oI4zbrtIIQUL14lKSWU3ZA1sVuqbPCbnqgYxLbiaimWAhxiWi4bZE3WC4Dp7UX/KX0oKTRKwDTr
dnYqSFLLWm7MR2Qz+Yjkl94xSPklj5ewCwjq5aKOBsvn5UeUiti3ez/UBM90CucrWtYHuDtGjN0J
E1jOg19Wjw6nnlcd+GjEADLxPi5eeVsbQJarKBuiTf+xIpx2an4FSHMRzazQnFK0DQZfnJX8qJZ7
9JhiEmEbDRy4X51xMoW2Wl188Q5/tcfrSSGLmVrys3+53cMHsqLB4+vcYJYs09zJEcS5g5DIBzmd
2pf+gzSJhV7TFJ/TEVleoktS4suQ21PLhXyaaCKOa7oa8HRk6hcTZW14ajWDv9AhsCFWRe3YJS/F
DPNQD62Wol8y1fG5yhBCb1LLegHSnO8k4j4FHRFx/eDhvuWKKM51ZHFZ7ekB7oqZleGm1jEkv+Ql
Z0oVBSojIf0DCLJhhxm5ntZ61UPi7Zq/S0mzWy8QLnOKsK1zkaVfIeZcGTm7ZSHLZjBfkSmn9/mz
Q7E5a0bx7kvj3Aunx9wtWOxf3C/g83lL8sMo0eNYVc9U0mBNEqtBsT3WrPjKuqTdqmlfZMgEqDft
yooF5WQWQKW1nlM1IVjZFb+rwxHAa9fU146+ko8aLMNizRIpHYahMwp0I9l/66kkcfbAn2mxqvYM
YQwbGx/V+4Q1yNJ5A+hMPd3ZxLkglsZALz3Pu0GsUtBAWvAqAQj6iexZtWj70FU/zVw18m7OSCfq
wrvvYupHbrBk6USY/cajncI5L+RGkqbZhQkbU1J7gU5++miBOezxeEmDra0vJlCdNcRpcN7AIl/Q
SiJH4IsKlzf58NW3UYXediAFdcipobp8f3Q1AVnWZBK0XO8RU4E7WefwfWla4ycrltislCrQVUvn
DzPiUEFqpi+DfjubF6kgfTlglkGlqYUpPPIsR7KoSQbl6p3yDMQw+AfMMV0ZoSV/ADzYbINHNUfS
QVjIgvGj1/9kLbgZRsTEbjLUXq8U5oMGpV1iFOFv+4Ls/VIezsDr+4PhGz85Pz0rn83TctWFwr6e
omWAS5Po6RdNTyNXuf9HbGRZLFDYJNZpyIuaLeEBAz1sO/bglQIAlWOwYi/CFkjMVRrEA1Nl0OHJ
FzV0BMxsz9HlbpRPHTDlVZljWVdDxvcFVYdUEQPdo6TMuUsY97OHRoSLERxiW/hNlTFACbD3hVim
wRKpHWiPthFYM7zV8tf5yPbWTJfMIDN/KDUOB1UxHLfcChqYy7/THDRGmBcjY4zl0Bt8hiS1Zzoq
wEbs8zInSMwu8ENOCGo663g84bWaMm8O2WDiBEHfBBLJqnjh5sZ2knVaFe2k7ZI4lDYL5ws3DUit
oqHIYKnFAVbjJhvVhzWeGTupjHU5nBzOfvNcn/z1uQADOtCxpMw9cViHNf5FtUjsxz3gpECC86Xn
08gJKCjnFtoNKjr8U9ZwrcWHX+0Tmt/kIp7N6tBHkiu6Qdhfnts9D27kUdg+wuM6joNKK8ukCR7J
h40oEmbAcftLuAYSyVG7lAJL0uzn9noBIJ5qB5ZwlYI5BqozkezO/WG1Vbeo+YaZjlACERtagRKx
dCzQX/99Kn+VEStYh86SfStcV3kkiNrJNClnVqefQND1V9rfbCnVRYIZ7FT585S/yxLq8JlnWQGS
YjHooks7+au/rQvdlNs7otw5xDKd5CAkNx2ukR6Rjc3biNjG/meQdrsdkMjZpe1BEEwVpTZJAXaU
BlzEKzghW40EtYzpBn0QRo6MlqALm0L8I3PJ3xu8Drbg6zgZRLJUxCSzYqciuW7ElKOsuVuuhQVX
7lP0vFVQAKpUkCcn41dNBPkSZSK+DM/hWPR924f7THuX+n7iZb80z7Ytdoxt/z2IVi6C1UhAVTjx
RPu/H+CEYVHZl9bEnr86K8X6cjaj4j4PrhpwHXS5s1U0h9B683JQ2lDoFY7wIQIKVffdFKlbxodF
AL/rG2RfFSsAdpUSSseHZ+xXHdnZxuPIIy+G6T/OSW6T+w1VVcy3MUWZl6Imw56NV43Fr8pTPLLt
8Y2FIobEQknmsXkRsCZktsZQA/PhLW35RYq+nahD+VCPxz2wCE9/CnWK1GOeJt0Mwuewqr2/lJ6H
CJosonQ2s24O6emgeV+eRo2t3+y1K8+0MRi+uXL7ixrTgVI6Or08s0505XcMxJg21yfOo6kFeTSB
Pe2YjIxm2LJc8ptxFNVpDZBMrzRHjSIuIuRQz/2rXw4pqzg7tmxDAQuCsKnGZwhP7ej5HzXvIjqz
r6YUyoiD6pix3reMyLvwugLJ+qDf68gAoME5RhkUM55/QAon6CRQkfQ2H+tfibhW8Am81Gkz1b4e
hysfnhvZ1yq5nAweOLqXQ16ULmFqMLbCdLQI3gv27OzPu3YLHmQyGTrB3HeMqnZ1mQeJS+lRZzwd
1zY2u2t78lfcip83dFySi2TOSccZbQ+agck9/6u/HDpofLZTrfAG6jEmb9aoDbO/8mcfay3TrqJp
qFbmjpoWJisu+B7HYpuv8fWm1qkhQgq/SXe3za7TVDe7GtvnHmsBZEqKGqyUUwuMEnyB7z8VpcSF
CBnpHULtvV5QxrND5oWwEqoIG2D2qys/1JD53LTbcwqDNH/vP+EWT9sgPCtXYq0or3ws1RtKh1sh
00eqeXCFSewJivvwWIwkZB8+GTVbI4njxKMzsjkT/oPRqWm5/Pfm4PAcILJFao6Nw2oXvQIa8ue3
BgZtG+Si30P0hbRdWsgGh3cPYbzlW7ZR/mr2l8VHL/YiTiUP98cHNVy/E05fTfsdB4vjVNgVvcEf
f8TSpKyxXV9e1Kak/OQ3JQo8X0kVsYJKl7sXzVHMFXEKSudUFSCQgxCHtB9PnHdgKQt1pd6uNwSr
Wo7x+U6lrPbYBXsTkD4sFL8ht2aGYlwG8uwZhxzzSUf03f38mGkoHb/EaL6oEPCJyUd+SrlOFoVc
ywC8Cr+sWsmLP86m+VrVTrC/4YHqA7KyZhTHQpmZKVDSRgEkKrL0MRs/latbA/bXFap12uv6ELSC
JeomMRXSf7ZzahTUII9vvNKD0/BjLCoGmAwlLLNAhcd7K+Or/xcxcdNBJmbsXhXorZPptNpeKPQy
6JyzN3pmte2c5Fpbp9DFtmJgo97iJzdvMNmX1Gk19iNZUAqpYxTgyjBYgBkUn5IzNw22JUAtOr6N
7qhllTrF8ubwzEQ8GNXIlLqdbM/Km/rinCzZUFeZYDp6mq3oQTuxzaR9/oZwinMglTkTtaFgZKjE
/Ig3floWWIMErWiKGAooZr2T7mP97OChaltg1vHI0uu1LN7HfdjU5bZ9JewyoAZ5nlFA61XyALSV
LfFtybC7OqwIzsXsCu9flKAJexs91jo58bdXNMToYhlOZfHacscH4VKgRfIm2/aVj/ovO/TCbrZ4
0liHLuJ7Zc6dIQ3sIJGGZTd152YRkfMS8SIqGjsjn3mtW2hFTmt37tqvUaF9Sk6x6WG/1q5+b0pU
J/en7/7e2Nj7ImIY0z7hAVfat8Rm0ZNDILSIek/QdFzSfsbcXPP2+dO3EexfXbvCJX9TgqHWTqAw
Chae/lEjI8fGtWadgT7qkJL5TeyGOgAhrsRCNBPL9P3fhx1lM2s6OCpXvRbkVarwBdF3EDGhLR6+
9JDp5Jic7+1Ix/NY9PqlngLjSLkmGUCOYWaJT1DJjSwMFfZ7e3kUKSkgRNAOPZL1c1W7hkMAgDoL
pkwORxxOXkxdbifAPW7ykv+YQzLnAPBDk/to6gSrbI8rPuNrx3JGXKpRFwkCdZVZTnPui3U/L+Tu
AmvSWwRSNWlddQ0XmKhcTNnvrY5ImF7pO5Kmqi91JXTjuj17vpQudwV/oa2gzfiY9XIMG+SFbjkD
ljbpmGz7WcWZDciOsda8pMSRKO52w0nr87Wlsvj0XlZMW2iI6GgZIXPbrvxYMufZJWRPLuE8zxT6
fyFftEaLWr2ecJ7I6foc2AL37g7w2bUOAP99G4eglTj/GlcKilfQH1lVaZQSj8WGeURFCaamZDsw
6btuXdFSyutg/aRFb9lycfk4McHHZPKWmvWOFrQJj8nF6+m0d2MyeT/jlx2Vqu0/cCQZsirWq4RH
0TF+OUQ7gsoSw8c5wq2xzH7moTiP5vO43Z24q48gQ+gW6rBowNtT8z9tu1L0C5dS+jdizxKjokC2
SM77iLrrKQoQp1fKvEbkVVpGSPRvT7fp9jmCFWYa1RuHYDN3E80GoUbQRwoOo2So0DY+y+u+Qllr
6kmrG2jUev7YnE+MrWUIiyyZ/QlXkwck8Rf8gHyndD+CRZhuhj3ntfGpFdHCaH7lUZffOFiXSuwL
SkXN6/GHFG4xS1vWlTDKy+AiRWi0vuSaV4DhaYuzBzKpf3YOAAWyDW8bIu86i4CzbDv8/T7urN63
E6Q/PlXIJI/JYeiL8ahKu9lhQR3reS3DaCcB1SqMAXz2wpCeeYf9IrTwBSRhEUysJ5eQNJQRbIQP
1HvQ/TOmsZk9+QAJOIxExm5VnHxrqnjyDGzKorqwjL/ys/sVd72PloX3pfnt+DHyQALD79fCtjc5
qwEX8J90AKh4L0QD3POwH5a4Plrwlgn5ymThU+Cv2F0RRLU2y0pSazkLbYTFrAxNNQnJ/T0ZRN0S
vMjDqXmi8n3yMBlHadM6wvVHYSMITBLH3YcCP3HGDUDrT502faLIXcZyduOuU3FPpzMm2CIf38io
nhHM6hdVdxycGF0qk9M/o4FP0mQzgx3juETKlt6joj0n0Gq3XXQk2ygws7yTpd70iR3mVBu7VWIS
383JWANgKTfG7aNruBn8S4gyqlWxbrYy1BnOH1a4ck5fEENEnKOduGj/CwnLrP4E2c0rVj5OgO/r
atkLaQ7WrkdqRc0PDl34o4sjV9W9kkvs5C7GLcQMLvZs0Lxc/O07g+0t/KTeQM7sxf+ED6H9/z3J
OJl96ckIWWM/BszXMqzuL9Lah5M0AZ4oPS21+xUoqOVeJKwZPkiVaumv4nrsTILuW0evFju/vYkR
lF577JYGJl9hskZcvTVrlD/xOZgUgqxGOenGYl7n/ltk4uPMOU8FnK7V7j4coEqeBiGSsWgzjNSj
iOEv0Np3t1SJvFzxqo3FiZXH/OCqtTMoc87cZ2jgleXpTvzoEi9pTujK2998dT8PQZUYv8d9pqVO
EC8xh3uCF7xupnuoQVbU5S1EtCzp6LElMQHrlYPV9PX8WFQn8TfsBZURuep/227D0Ku8p9OV0mID
FAD2d0QmS84oWmF6i400u9vhQJ6OCYChFg74tgyNpeQZzeHAA0z1cyzVWSxCkeM95ejXtdvtr03H
jkC9MlLtBD9co8m32IatZIuHOb0bhWEpUmiqJu/SRe1NE294YLXBvSubycF43ikim1YxypwC/uLZ
EhClRQWjbRxbuXIBLmRHhrAfXtMrx3WUOJgQsquVqRQkFT/CPXdRJCyqBWWCWl5aEDiq8OdUcjd2
mol2u+C+Xk/sSgk7jLxyftpfVrtfRpUjw9rLUAq0AnIFv3+CAQ+jcfRf4bD53jPAqpoYt5JvwgSx
ehjcTd2XORVZBLmZznx4QYIvKdH0QVODPeRb8PqktWcbSm896lWrzRQl+fqWicysvdo1nxcJvyMW
mCwpr7twe8cH7zCBr40C0YAVF5SqjMomIjufFG8e1qqr4CIX68Z8lcfpo5l4Z12+ObI9Bu43iBIp
3BdHwJovORe+aK647edDaIr+vshKWfSlTQyuRuIDnD2ZozTsIIB17yoxte1W5tV3SGp5N+mF1Ly1
C/J9dlgUF4CUiqdwz8MIfGYs1HICjotWpb0p3INtPuvI5UHjZCVO2K2kB0WYU5UZcbdq1AgP2k2q
2Sj1UvTw1xWSYX57nW6c7rUygVAqXI5WiBefAix05Eu46QBlb+TRuGD9Bb6zHp841L3FzjZuGMld
unfdocjmLkfQcoeEmimCmihjRXMgLPWInFxVNQ/cKWKXFwvUGly5iIUNToxrKxGGS1onOs2md5zs
FdMPRKr1T61vbZpyFdLpNN/UT0S8ScOA03rC4HlWFBUTBiVifazIweYw0wGr6CR0r8ZSUlSag7K4
zer6tXSAZnFMW9z3d4uh8jX9LuzJVVeG+/w3LV0RtTFwNZXk4lA7hWpsCMmRZzXVt6XoHtaB63Gk
guM/2xvCLCpAgCL1MoMdH9FkG1UI1pArow7443CT1V6ZsMgNdHJoT505ZZ6/wDHpzuF8WLQODkzA
yNAn5gvUc0dIJcWPvD6sD/ycp9k683sb4yuEXTOgao0d+xTJtU+Y34TO0DM9rsNRGstHGg/UNi6c
MJgcrcLoLO6ri02DLmLMGk71Q5h75e5xmQIW5eQDu2kJG8JTCK//SCkGCR1Frs7GjOpu7TjRzf9W
FaEpbu76La2egFcvvRwPg+ZQnZX5QNGRy+PVFxjoK0oVIdsgZs2lJtf1l2GjuDfLf+tij0R9dnnC
PehUWyPUdS7/2RU4yRprezkS2cID3pe6EqLJaiDsOCT4+hjbWkY9gzuEK+BFWeJngyVUqWBYSARD
AiDh1lraDw43+9RRZVvMrXCcb+f50m4IRtZPeb7E/pSuY5dVwKm65yU9EXKl5PJhty73qauf7nlE
R1RCWWMd/mIL+Lgu2VU4wUm89kpbXA6wxvKp/fBbVKcfoyYidUy7XcJTjnBSdnj68SHcKMR2bli3
e1igXUyGu6MsBxOD0emCevb0XeqOp4uD4dikB6g9pCarGfs+XGTTTcfa5F4rprG+AlandXOtuFtR
15fQzY3MzVmodp7D1EJ9r55985RG96vN0utmWU8VIf+ONlG7PGQt+ocC2qkhxbsAUGvJt5ZPEMKK
aynYxY4JlE2FkeebKt7e1TJSRyLfBqHVVkLNxtOaiN+ta8+FX7bHdT0zK5JwDDOmt7biFsKMQK2V
zXb3PSZ3ldwN9y9VZr3pzdhA21LcOGCgqhXXvEZY5qtmW8AYBFG7OcF9AtlgWXxEmTAoqpC1EnAP
9SUu9PQIY3J9T9nFWPR0QCjbMtFO0+JNnRvdM4C9imJs+YYwBtXpLZZvzGyPJ8OC2yfC8M1U9Uql
+jTX95mSpWsRNrG2XChbqjGKbpGD31nkyuy9NPodV2PTZEcmf6QVo496RogTLv2HJEA5ZiRjH12m
TCY3L8fSPDop3UZnlY1iJuTXPLkFFoSK7b8QJizychKtjLjUU40O1FFRPP6JM9++y6/HNLTHYjkh
FhQDa/Mgs13r3nhljF4gkt+JRGgvr7kyKX+ECBzprPO20knD+KFzFg2ur4JUA5Jat9ba+knQDaCz
4DRaeWc6jt/uzqJ+rID+N/5mmTDZWZUD29JHjmLwK8CqqLPUlWqSIEWS/Qtwp1jxoiPzMWkpOE70
Yjss+fQtb7Jc4xhq/LZ6A/ZBkqN/6Qrph2P+2a+zDZVDVYiNGi/f0xHsPGqYxM6yD7SEvu46gQTt
c5Lfof8hnHOMn6lLvJOUgDT3em5yR/q8pHYEKnKYVaLr/Czf2yitrtCbQY1SRF7iWKCnYaNtRSGt
TOUl0+LiOH04b/0VUBQo97uks3IFkWxCLkC5PYJshQ0NCkedJeUYahUFQBSzMmM2WeiVznxKkWv/
y09EUd5VEO7ua+u+QliCLR69Rtl4VB+igPC68Wa+i3Wr3kaJP+idvuyQl4kU/5VGAHy4wvzN1rtB
Yyn538oqUrr48IWsV/cjWjBvEop7qTZt4iWX7FdMgPeq3ZYlRNH6LLsv/jRBw4S4dmK2+txlKzmi
5ALBwaDggLyPcPeOzXEDFeknKc/oV3CKlHHPgIlB1cirZ5KHvGzQ+xtJVc24Pmhgrz1cc9eVCmE/
ulYBZmQDOCd9nplXk8NWt0kJT+jr688JwvZdkqpU0HOgVaJJn12b9BIuAuG7yLI0vNlOnrESN2RG
yv5oXqhuimJq7gbraSwxCT7Df7VM3SN70cru+LhjQmcETe723GgTLiA7NkwNLKuQoiQRYUWL7mSY
U64iBuiO+0TqdxHygVQV7yRyc3S3BJJ+E0ZrZKHR3Rrefv+A+m6+xbuFw8u+lRKpSh2BQsf0BfSb
CCTxbbz/NvYyK1c6MH5/CtvBo2hoB6200iD0VbQ3IToN3/uQiQKlsM9O7kLnMeoVlb8ini0i6atY
/npVlwjJzu4Rg0nqAoHHbDaTqzSNrmBo8rFtfh7vvK3EyZY3hG25l2GeZO4QQJegYQn1a7zZcN04
HUwUdymqbgJPTLS7q3mdsDqm7vLxfp6KOWtjGoEE9jsFUHGMq/u6L3pp7Am9YG+kVhdNILQBkqdj
5n6IeloRzWO9E6K+w0/cQadLIGZEDr0Kk0RIQ39cuVQqUr+rstMgyI2pks3kz3/KWpJHwGbCgFR9
jiWFM9cskc89zI/1HKuziGc4wG6kxhu3BsCHPFd0CIzitAynJz7a+m7rMKRMT6QLClPPUUu+oS/X
IQKvOQ5O0qeTjydbQwq7U9t2WhBq1eVXKp7djzW4cOl50uQ8zNC5H8fgx+azhCVmO57icx2VTOLG
jlIveZUxh3y0NVW/diGXn9S3XX+ssI07lfYQI2dodAvAHKce4FOKCo/4s6ociUfDYW4lBXPovao2
g04WHwKAz1i4/b15BDFKi8p+U+iUs5amGIb7M9zUM4VXgoFk5ZM0fB7+dC75GOgx8DtdH2H/+FfD
uMVORiwK6i5WfUAQ2QmvwMu5nWVArhCXE9l3ayDYMkYW/7Z16V5z9dAVpcqvLbJ1Fdim5aqkj1EP
nQ1Ex6XPB58Dr1rP3X4HyhgOvoJ33Du3WM/vvOSZa6OARKrdJ2knNqQrld2kxVRtIk8jyIimwonl
AjPn+uI2sUEL7L/+MDjmhYmmWeB+X2eEN1FP0HUTvLvSkaMhUllJORBnQRf0DhCoE8PM21GKN+/P
yO6MOx02+iRoasohRFDQCwzhst6ERj/lsdOujLD+0rqthyzDIEE+AeWPVCOTeQ+8P9bchtHQtutB
kN6AnciAV69LNSIh7lPCBSr1Z+EeYQiAkVVK17y0Uz8jQf31c2GMshVDf8naQ9ucS6xN4DYhSHLc
Oaqy14ZeIroWOMzVHUmIhzBBPJFtE17F0BdlvSfDaZHbGAWoCCuMDArY88UHhiIKcvZ7QFrxdS8r
FiezpyJNNT+1jXCXoQ3h5shnI9+XsvHxSpDwhiSkGnQw82WovWOCCU/D1IEJZMoIY2EqXCZwrDFL
zChHpPoaB5PiA3EfnC0BfGVqTKjexR1KEfSPo0Xo7N5/tn7+yXnYs49rud2YDtiFjEga0w3SM440
391l+A+XwecY7+LzTfYzJJ6demKxVrqv+DywRn629F4WyVsUSduI3QI3QX1L65g8kfZjhwm5zf6L
SBIO080mnUad1jKVgTxLP/Ju4wCBL8Zg+0+WRI4tX9alxJ76JJ5mSKojAWxWamvN0Tmttwc+i3xa
EgeKNi3QbhlLaoECQ2Uj1sI0id7DDGuGIrGJfCtGbOSHY+z7DituXqXO+ubOKEQpYmcY4ZQfnHb1
0SmSr3CnSToh7ciaQI8ipMYvIooj4veVdMLyFNEnH+PlYE6n2UvHdcSamjEzbzfyezLmcw/alCAc
OyggOtlvncMFhRLK5XQa7zfnUDqiKXRQoFEcIbJSFIvBHe4n1PF6wRa86Q1y2VJODp+g7pRcu6WT
znVrs/iJTH+hTutDi2K26/P+tHz6wykEYi9UXXy+x33mrk6X2Vk/HzyANdlbWY1VoK3xp/N43S5g
N0K9YSHrQeYodePJp0+oD8GeEJ8J4XRY5GtbJ+1Gd/dgP63RdAf5pNJ6uX+4f4BhwGksOUpG57S/
54sxtdBxaPqJ+xGZAt57nCIzOhz7lJwQ5arn3sUZ41Jav5M5Y7RMQ4OwBvOAeSfq9BBiHQV+Xw6D
gtcCeuPp8wGIG/aR2yOMOG5kZ/8oe6LeZJrY/ED9bh70ieq4ieKQ0re3poeDT766JvXw86naNPYG
hrt0JqhkAiWyKdGYFHGaOctFnSYfFmh6VAlK/AYdf9HUrFrSCYcAE1EY7InapI4nLYzgOIl2TAc3
W7IBNlVhPuaIq2LCxwWINp5HzgeKW0IN4ChUNHOLhb+tfI6FAJyZRJs5UE8KzeCH8Jl+ALSimrMz
Lsp2dWV1NJvnvqM6blXBZr4FhHjv6gry4iLM0HzVGP/BYUDzN49y1pONf+IAu5WOrSa+5yfGsAKl
S7YJJiSsBJlLBgAAB4mkWSvBx04Tp3eL7bSCOCToFeDocTHgYPiTLZmg1Uoe+LshUd/SPKJVDaWi
ALxHV6uBrCkfvx8HfgiPu63A/jLhezxFqEqdCmSNu0QDoeJOq3vXJxgRhIDaL16tzbuE90Syt9bv
1OFDbpJ0acvlzAynQJcAsxAWtNXtJLjvKM2a/EY8IB8FHvm7nGfHRf073dyNcmvw8Xtvma7hXeTL
cAqPb772lFaL12jMxtZFOvx0Won+tm2OWNFl3edAEo+Li+XJUt5ND69pg8Y17tAGyhJ/9VbMrr5B
bu9W6KxsvIPXXXmsjLcjT+wFbLohkUjo3gU/HYxAqnMMPIrQobcmpHuYlfvrAGsejNjVwYluE4Gi
NIvXT9FN3xWEHh1uUbZz4HiBoUvdN16kRT96++mDGbpr+3+MB0+aRWxde0+bFmOtR945tjUxqEP7
GdYf/+ez88ECoNDOOrbbKGZSCEjDH1mGkELWk67wldHX/zC7fg3Dd/MU0yPJgjb51utdt74gg36P
gi4fnsQtHTgRCaDzoFlEZZvpH20hxU+rQLSFd/nm8c7+PbviPHi+JMfTotVtiihylqhG53dSpORS
xjp6iZNNKOfI1njHfq+5sdOxqMm2ZaRX5LcEVfyMjbdpxumwD90Nobf8Cv5HR1iW4+7N4DJmBsBp
FkM0QuUlRMXA0npuQkUYx+tyKmuptb849RHEqYA1SHZmuKke7t783qoBPlJJ8V+2gODmlWLCPtsw
Xf0uOO8x4x4h4SWriktZv0uCYgbJMdhT9Z9BR/5JdJwmDsoVEyj8ei4YEWfQKH0OvVpIdP8ztEZA
RsN+Yn7XOYUdlrojgioBFdq1wtR11ReGLFIOjAELWPWrdhPtsYpJZ9JXL7qYLTQdI+N6A878UpTz
gRBiTkWGvs/j4dGzMzbDxmbVUTcAj5wC9n2hnuahfnHemub7ypca3PHLEmIQVkhUr7s7VTHwZ7UB
N1GqDZa6FoMua3m8M/Zd+fyD5e7hI4n0D2FhOgZjgKxRwdrkvbFCp2SP8fRAaQitq/xqJZ4BjPGU
0Gg9zbPNd2mm5UNDzmZ5EHQhO/0dxAdCZinmBvGf6nB8aptVkHrrb7Fo5KCyUICC7ad24XAWtF2U
+omwHWs8CDtqB3okpAkNp0N++rztkyeqXYcNQLyp9HWEjlCNWSfGDAcq2vs2V0DE5IMKhTAth9tZ
8hTQsqzxmlVDmgxt0g3xm9ZFWWG8M33vrVvE3rhePLH5ZHWHEhNWfZFmX5MWm+4iWKAj4zmedikw
RmcjXvnDDWmq3GsvwCv02WvJ0DRQLVXFRFcA5CXXuIRCCHrA90XGHODjxunTSUxR+Ss5ag6h/Qfg
menlfeZLdYYaE/q6tk0UVy5iuWPmyWUGuVRPrHC9H0OH+dZEhi22r00a7hoXMuvTeLuQclxIJAbr
Utaofi1yKBnKNgMifTvgmBFxm8XmCTv65sPzNDclnrTL/vZaznRBJrMh7Mk+YDMj2uCYY/qdgdkR
LrFhWYYA3bQl7SRHyFTQ6OwZ+vbSSrXT3H0ivskui0G/sg7K5OrHfbHy0ia+vi/8DgxzlJJv3hoz
eQspgMMbG1/omd+ZnxTjXZDTvsegsHPiD3AqJj0vV63hqkTkGEdcTe1n2+x3JDngQnxr+/wMTiS7
PR3dQ+qL3vLMVAJwiwuMwuHiEwQ79CJNdXnMFuRvhIRzX8WuYG62kBPnDrnzDRD+tTL+WcBmL7yx
O3/xhbDd0r009e0xOM8zO8sOsO9ShI3IuvNuebjUE5iE+lKtIoEQDHXPhgvSK5wvkEit6WFtJgw5
nOtFI7qkHhDlkbgnjIYtnrR/WTr99B9JECZl5/rzdWm59d1EdbvTjLZuMtzlV1LwnI4JOX+5Q9PC
bhw625QgonGVuTUzYRbziYQAGoWIIklhd+Z4syz3UZdrkC85lc1zDmTeJRHaeG4g1LrehpH8+cYr
0ayJ7nSCa9Dn90mHvsZnfTyObMD+8GugEb+KNlKwr3sqGrDBGpDnDh81ozmKRbQUET1M+U3QMGSB
T34vBvq5ZcJAoWdHeFvEkjeCMNL6n9c7Gzmwg+Jj2mFk2u+y04d9Y0zHnDmLUxwLLeUko4SOAE+Z
/t8tzl/Z7LwaZTF/mR3dhaRAgYxjhqFngKrJeHyXb+51gAwjuFG46eFwDqsr4kkCv7TIyMsddkbH
xKUo9LQWGmGDBS9qRgwc41DNehX+AK8wTxyjceGKJzpjal2XKzAsk3Sb6Lo/4iyk/YyOsJQMYmb8
d9f8KE0t1UzouqL2GU5CT0giqS9EYxy+s6uwiNybxxVT67VE9XP1SIGjTEFaSZU3zd9kA+7dLWDH
7v9TE+u50pD+Bo9MmpgSfzMsVOiiAoCcYvfZCyZotJeElqcL5FY+LACKWT+/6iOEE+on4Yet929M
v6sKSJe+7aM1QBu5RFldNUYknfLpVGZG6iU1Mw7YVgFnYieCjFPuIUnLZvsWwH9gH8xZOKhi1pTu
93bMR+q8YZ1vF9B6OT0JFrUUO5a8mM7sD3BqCBIeP6DR1jkxTyQuMwPXME3nPThp/B5l61lQ+qbC
KN0AfV0YIViB2cG9D5vfrXOkNtfuMJJyh8qiT+y7yt2zxKR42pHHVgW1Lw6fJaq6aFJNBS9iLzOV
Woq5rJhklW0W/olyh9Q59nYKV9wR8EoTvK1hGxXcZtev4IBs9y0ToScn0Gyc+YV9uwaYlmUYCIEH
K4MdY7rxk+gns+jDT6ubVbhW/vj5qBxzs/JScmoPEpuwUege2YGjPZQXA/kcqKr3VocNT9A54cT/
lFkcMiGIRMaWTJruVM+z5S6PrCZcgEOiQbFirwBzQNUxXD79LUx16hP3lz6n5kB014yxYgXsd5zw
AZN4InTRRN5uQeGdWEJlyRK0M7AWz/0Rz8WF7YfoDkVgpFxyuA0PJiQ0jddHIjoOQ/jkae3sWHux
lxVwRPviq7oQMhkVkVdvlJqOAgoxNN5wfZJIKMfN44g0kreBDGK7i6D5852mvmiBzNBsJLcV68cY
augQlaFgzXQqTXPzfvY6M8JA5Mi3og029SZOSXoKQF+8gxByzd7LPpSKXyAQ3vclZ8w2joKprFWO
6HJzF6RADiTRBxfFeM8tH8A0deUU6X/ynH4Pbtl9DCP1LC4LLZSVyIqMzT697sfJ0Xg3q2y/Auox
h7f7HrKDWI6q2TS9HSd2cpJiVjlKgxvVaY8dG1A7QvRSTsBMOKwUqPo2IqEn9iwByYX8RKp1J9w/
Qt6SzW6c3LD4x54wxNHtizXR5NLldMKiisBinzExDtkF1MMtRX0yN56NRrsQBJ3AWxOjlKrn48WL
mgFb2mljuAwLhWkYKyKENxvc7UPBab7gmg6driAIT+hltQq2s6aeF4aNGo3+/6AnpFPndX6NJVnO
tUTpsGEOu+siljzI7WUm7MVjAw5kstaFKKJJzS7obEY1VHSja9X5IGljdkBitmFXNYai5ZqOoBbv
wethU+j7lFi/VvWZ2BSIbP+QYoPnCug41YVOxZ2qxDJqRR4yzsr1RRvVEwDgLOIx0wDnsA9Db9mJ
mMNpDsApw77lfx1vu7yhFycSefNKHrqrmFY2ESsAbE9mLHUqnuLaPOYUgzgjbb8m2iyEQ0VDLvpj
HKpWtNMn4tjNR/SmQ5w5BEDahOWYHLJXfKlfzSMLc+1nDmDTWxMyTLOENPTGaGj+vsDWBDPSVudt
BVLgjmrG72cconac0FA3F7JtwPwQmhc3HPALz7t1eA8gmSYjfXpJ+e2OvthSpDzpARBrRAeUDbU2
ZrwFoOVFVp9pUcrzhwvML+3BdqHVykuyEoHxzAJ0RcAZXJS+XIlsMqkr0d3n0PtrSqQ+TqVNO8Oh
Lmvqf8dvi2XVlOv2jsCvOGm/yWj3D+Kt3vKrtMSuszUrwkS22gmt0D54uG+3A6g2J5xAT65ILitB
VPVWhUovgxNnKXV+UuPFDLXsBa1z9RhJ86WmdL8W6PHEmhfHKZKFPI68/Bu3lSUtwJhP1oltSQDt
nhcXsk9yHBwcbi26KsC5SJEO7iuje9xHXBtYwoJPivXu7taCEwlM0g6RvquZkYadxrIzsQnmKcr5
YzCEzGRhhpptSo3duMIYmU8x4rysorMyN3+svviiI2j9yLk6xYawzfJZ5f92zGp2rfpEg4sLA1P6
5xLiKmK57BpoExrKU+224Ln60Igu0q5mI5TOtKFSRXzVcSW5S7RIjtKHEwY+KYsPo4jCagF/iMx6
99UTdcGJRduXQyN4UPKvwu/RNCNMV5lCzUGRqUuVDko1v8qglSFRRxhfPl99DxoZ5s6X0HkaO3Zz
pUtBGZij0P8XYhoojc+GZyRUG8xwNJ8mvSATZ7hWfRnIx3b64FIObXg+B28eD3LhBxR4WLt3J8KM
rgQdzUJuogrghZk690L2vHZWaD2BT9J3etI/rVjJbaqKQ4T/vEJ2jJ3uxfiFOypP7LLPvUYJ3Wap
nIo4Ur+v2TvilUPvCZxz4qzvxw/nglUQGk20axJryCkh2Qn5jypcZWAlqb2cmrd7EmUzwsM9V17/
3ZgSVDYgiqWCURDhJgRvMCSbCEUTSzCptSQ2BSleAneDrLdNfBNc5UcNkYje0JCvf4s9gR15/uao
Eetxma2lyk//8ukebKiLGsCyqeOtlmD/TmhSR3cZ6HfWc3ljLnpBpfGCLq7csJSpf6fW8QUc4x7O
aE6ZouNwkohSO4QpmFFu9PsDtnpzPf/MrJoc8vUhmBw3hW9FKDqPXW0YZm5oyaAlreQ5f6pS1GLv
hsC8qj8feOlJstZEFy8KsxhcNbswZpf3Ti9YjTdiziTNovzPtIvz6oyeGulxbkSuyWD1DlolbSeo
9kKxy8NsWvOKSTv3WtXaaqRqWP4R4w+atu/6SAtu343aw4ss0YqBi1ZilZxoDJ/E7sODJRWTyZco
3spzlXA+e7gG/9nz/o51zjERAWP6YoPtvYkE5UWiEQAthz4JS0LDZ5mZB098WJzQyXqoU8QI6k22
ceFa2HFiyXmQoYlNxZUYNAhFvZ2XzHhLBo0UMwmm0dCWTOizTwPrlGX8BSaor7b1+zpjfkItZTvV
EF3H2VefwGq5HzaLliEq3sVVIEt5XXObzt0y5wI3mExw7Gohx1U6sPx8oF88uEBNKJmvmcHQzrXU
jir6vp6gVRYIYVy5k+hKnOHVH8Nf18dEPpaHJcHWnVJmlDLXlBjZ+btWRYOctVnzxV6tpDCjc2bs
+UQCm9tmKinBcO0030s2IzajxcIs7IQQJ9RPPxKFyx5KPrnkxKCxADmo4WVb3F6LoIhuaii4vDKp
rG8dULlnDLaNRvh6n4veT7RU+m9Va98jVTrnKmH1ZRRUsVkY2Fmi4Mc9JC+QxJmaWivSMQWjsS0P
w6VxnY2BtBznrkImxphWhAJuQMYMunLrlJOplTnxYwlY5Yril20gzlye69SzBPWKbzvn27jdeJoy
7OBWiQLzgdsM0xce8RoGKpRk3wXviibWFLx3na9jHyRk9XL1Nxd1E/mzab4cOwa2QFJwhvXYtZrP
LTOFknMBCxQOqo45VMWiDaM2HjZE8nCraWWVn7tg2rDu62+shesJiORHJu/Kr6FX6XgcjsUzBTdk
JjiyVuAMe+yYKQqPBCWBiZj4iAk6cd25L8whvgnlMuDPokRZeVOrb7oPzIcwODXdexl52waXh+r5
gFW6DuUEG44P4s9PrIKSQwqRiQ8fe/l9SQ/CtTb9eYP7l6kDXHq/HeBhVkqgs1Gal/GXO7Ol/dTm
rZSbKo4mAxmN+7bs/5kSg+6Fpg3gOpEqEYsmkBzt5xZYqx6A86BGqLVD1eHhr0MZ1ML+iKgJ1rve
hLlpV1uyaBR80WuBJdLg7qkbXJkKnNHLWBd1LcNWIX32Hof1Y0pMJJzzsNV4auJqj+2On9SpH4Kj
1TiPKB4Cf0v0hEewSwiwB/PgICoUOWEuyrThHaILh6L1FYMT19UJYaRRe1FskcYfF+TcDxHNYUhw
PJknGfkG5OOI74HPZud0EGbTY14Pa9z1ivjHIdL7uAlH+mSDpXm2v+MXa2oPriRJNChnjhxADQuv
vkFu+go/UR6g4MJA65XWpcmY0uhkwZutWvuVbiN+k0k2GRso1eFWqIv4Mpa155OjcdGpO8t36N77
R2rGHly44qo5J3seGy6rBgbyAVEr7dtEYMAnREflBESrBare1ZCkQtSLBZ3cE/1Bv+24ssSYHOno
eL2MKQE2Uwg3MfVmySKZZcCbffEC1E/7sGC6zxEW5P22elnigXI4Le0QtBND1Ub+W80rGZZXlIsY
c4oyRx1xNWIQD+5Wkh8rZK2b1HdOmpRRpPMIoFWGUeUbaBaNv79oJQN/r7EEfIteJntpMX893OYK
NiLH88tpautFg+n4dNfLwZbsxMuFMzWB8Xe/JNjbC0o4YUu9tAOO6xCnMMjF+f8VWXGpferbhxiE
pZBLgw71gtGZ0q7TYac9WEsET03D3VzYtiIBTLXO791799Ew9j8ibGygPQm/VncLzG5GImtaG3LN
1fPjK5BMk7OwYaSGgCeDDvXnDIsScphdP0nRvGKVG6UQWY54oxXxY4W9CAI+ShditchobTvDhNX8
8rvBRBbjavZWX+lOgAfItYpQBeTXuG3tdMktu3v163cMCaaopv5u3TRrduVwBYKhYHhBOSbXY3g2
EC362wdN0kuXVyPTleKhBbOfSeBihK1BPuhe/K7BdvvwEYO7s+2Y03pS/V3gMiAjvaoOqv6mM7tf
oL74FxqkO1824kWPWsFxWanSuqZDUFhmJ7oYpgkGR0wGnE2nQKYZO6BhlQuqPK95tHbw0qy68Sn2
v/Y/GP6ubaixCFsL8AMO5iEE0qMVrs1aBOgRJ45YOB5aZM6X3dLyC0M++pm3opyhtm/UFHjV+tu0
A8NtMpZILmrrnxnnd+I+8UTSJC79NMP22uJWssvhGrIuJB27jYJNO7ur4FLrC/xt1XyeBOH9mGt5
njmpsY3K+1BNhz1AvpPv8CioYPBUWZMslFhnCq9fdxs5uV/TijTgoO83xEuq7aUM7M9WNFsDJpCv
LXGzSszPbH2DyAHpvX5ga7G2rHtqxDda/1meI0XJrNCoJhuhuVmiFlui6R04iN8YwqIsKNlEqtV/
UjL2TqAZoegi4sMq0ISDjd1nQosEBm+fZgvo7ouRNWK1FlwnyOEmWMxG/9w5O2t45Vu2mDruPd98
uBoMXsAzxmMRUmWPcb6raf+3Ai52hnDaFxdj/rxC6h1QDaBSw4/q10RxCFI87cNrZQLt2BUDl2dJ
C38++cj2F/vH/jUODlyWZJ347IwP1yGzpF2Fb5TO3y0BzGGOwdk5EBi6boozBNuVjhLyuZY0dETF
Cw8kIlpn/ALklOYKYyt32R4LRTF/qqgyGsqW/0YTPcM2nfTqLqmVuBB3v1yR6nqTsf0Oea4j6+cO
xggXm8OCB90xfxrDrwG+i+ChTV/jYwecF7G1rlPwyV2PwH//AfN0q2cIrn5/y6IBvikKGmnIf/LC
obYZPjt5YRmvLzHRWn80mLVJUuufwp9gVn4I4DYl1Q7SkPg+WF00sH0yRvW42+lQVqW6m17SBn9q
Bpzk8/4m4wHFu6REqjE44v28uDXlO71LBkATUbFgRP6nqjUHJSQkZ5kUM7m/IdX5WwyDJLNDHo1d
HOM/9EZDZum0fVrk7+lViLj70YJO0IPyjLr86aprNZKqw+zkB1DZM7wDifQfoL7QufgxVycKkeDp
ZTj/u8PRGgm27nCmo6lF1ntVeg+EbsDGCIdTUWKhsTQ4Ubex3JqNjWRUMDRleSf3t+t1Yeszf6+7
f1bTxoZOV2clGz6Yc9IVBUhkmPq0O0oDrPy98hjf1wGlm6NRbTOjNPl41Kz9T2k9kupsRYkQiwFE
0bYrZItJtazAVpIGe7Orv3p5pouxVqEPbsDC+ikdVS/PQuTOsWiPgi+nEm1Hk5a4MvVpdM4a5oht
8HeE+GT4Kgfuw9Xjn1zbY5/+ruteA7y+3wmYMRk3/uVpP5iBELU23SFQE7yCz9Nw3btVmbSWah+G
79sJ2q+SV5mf+1d5xy51GPx0L7UIkKRbxZJ7eaYZLsMOa4YapQdDyyEkVIdOHMc8GLRSdFxPJx6X
6doLbp3kmcP5etBkIgl0FCgO2UbUrvxeTNX4ewgl1p7a+IJ9S3bJIKyxTQbu4dcXdPIcDxfYUl4w
+S6dOj8ZyA210sLhvSyz0B/rgW27fcux+rd74Fsb2V2Ji1dCb96mNAbHkL6qFDiKDKoCeamasz01
ptDfbrN24SJdReJHMcf1+Qm2g9e/r1pwFaWha/w932Fafc/nXfgtbbEzVR5WMVUUJ4wO/+BxFndr
Ypy/AR5/+RDVgXbX2D7o99LmPKtzL5kClzS6uNOnfk620XjAfd8JpOZzs/fMK+jiMuHtugZuDSAR
gcp2H/nVyOEhui3TzQWRY5wuAyNaWg885VvVSIVVZttSdcgA09i35Ji/Whj0Jj/miGqXeJCH/Azh
BDlS0YlQq15IATdQ88QsvRhhdD1q35rsgz08BxCD1VqSgbZwr/J1j/liB/IhophnsCq+HQRY7R25
gcrGnMPr4wegiBEaajqUTdCXrdEQEriA6aektaUUzb0san+wt3089E2eAw9b0wO3aPhkYfrbN4Be
DWTJ7hEoBv0x5FW8MyQC7opjVm60HRepqgiL4p2Flbp7UkAR5ugwhobn7lERJyoth5B4PUT+ZPSR
b/T1/W6GX2nOlUQAnW61OvD4qN/USCmkNZ8nKhLbhoOx4/QWMzxc2zeTwxl1FsRd6i408QLUTPmv
qAH2ghfwPuU1mBoKlGg5cNd5rE3TI8tzHSEVClAgAjgb5KZSlRJjvoT4JouM/4m5ey67YEcxZenn
pC6XKhsQpZyNHRb1uqxNndcdLJ+tVkWyWflZsYLr4gxMWF6lWV02JlUzcwrCOLs42dVCFRlYvQru
DAPPfYzAP6Zr8l9OVIjmp09s+EZ/xXKqLxGO4RtmEnbPvMW3iGkAeSdv50TUnRYPW04hD+9LOIqS
UAvmWuc1FHnJVe6dgJ+omZ6J8Hvt7mzFBc6/FLCHpH7YFHiwXxZfs5AUGj99ftTiKdzQMk3ydgeo
TAu5VIQjXj+BpfedLZs06bpbjLXWAEu9Kzg/6vQXYsOwuc+Pd0SEypqzBBQaj+qAyHzf+iizLJvR
rIRNQbjuVuBjzdpouyrfi/Zckcn9W1MvLsu82xPFvblw+I6Jl4lr2cdNe9PsKn2I9XNAwbPMMEte
OCeHCYaX0cZ0P+J+vPgL/AQXk70l/siL3t5628QSC0SLqE2MWvunrYQrkpXpSxM1+/OhT0YKR1iW
CrPPywDu+djJRGYjBN81lnbv4C4yutd2VlZGNh7nIqBIOAFVH6NIt3XTXH8FNa+5Jz3DSUZ2XEq7
siFQo5ygmfvWd9TK/LIh4uazgu+KtUZiXjA97jOb9geZldJWUHh4vOC1gU0UENCFzBdsKoWh457W
3ZFQeUQZMu/+IsuBC7vNQJ4SQu9RJdIDHWQFG689ksZgRSsxy+2jv3uzA8C2Ougi8atLySW7STwh
zmRJAMwjL38UtA0QcME1F3om2pj6bVmP2AMEEwwLiLro6gb8VqZT2lJqMWt2hWlvqvd39guC3uka
ZLEfiXGGIe2kojsTgIcfD5CzrSDlHxIajBc6wpUvB/iHVG90NLFnpbKP+BcCAeKzdI2gcl+fNMaW
xuyGKWRQb78IHbqYxkO03Xmrh9WenCmnpbq6vLsTyc2nUYpw+rWLs7GG7xTauCiLkmXAnAJ2GEJo
eeHO6sMF/DWBxDVhi10KBgnSHfrXW+Xd8e8aO/o7a40PN7gygfEjrpyD5OqOfTtSUPAUPGUQUkVS
bdNDpKTyv3kl6hDv7OPvwJA5M8G1UvnGg1diGkeHdJ009JjigstxRnJBrGdbEoAm3/Wq2rqL9Xsg
lMAKLBzjn2vwR/xoqOcZbWHx0clKRPxKY3YdSpnj5xqEsl2NgFoB2qXJdShzaYz+0ppX/Q/KjCOF
Go2moroj/tm++RcSMJBWzgxUP2oInWX950lMLRpYw+03Z0hP1Bcw+J8zhoaUI46vIYgP7Kda/b7W
Ex/OXHvVd8co7kY1aNXnX72/fSsYdovEbDd+v1lE4mYxCIb0VAEST0o4vsHjXRnuFuArzgRzqfLu
JHgETrG1X5OsIYkYGUR4dwxZe+R5vXfETyF1tG3/ndk6h9jUzbyz9O/t04g6wOA0wOa+Dl4v2dkb
BhcdZtemYsed0/jbToyXPrVgs8DyBzIRMLMBpczJZPpmFC62TUT9GZG6q/ImZym2j2DJqYfzApYS
tvcf7DFXQGkNuUHaohzQ7hASQ43RP38hxKmOVHjK8z13LyYz7nndpfZJuONM8hq8ZcVJjLBabUvL
u+peUKQp9qoridUoT3F+ztF06F/+6TLFUhWtdnXPJ1BMCmx9k+w3RZVUX7BRek9BkRGCOJ/o6TPT
m0O3GIJ1vsd5bl81Z+Z18bVQkp/kqBrscft89y+q0i9Mf/2cB3l9YPxJwXkj9Oq6PwAdzBNofmn+
jyf3dx5FlaPV7DEYAZE6uwDpf8obPMEqc9tq6Uxr7m4GJtPJBo9a20w8ba7aM7CvXJrFdkuFISrw
p1Yt/yiCnYydiPC7BSK27PZNEx8Y0MrN/REFNMHEKPmWRP3AK99Gcx/prUlwNAdkd2LKUDJ5Pc7X
W28jYIDMG0Zk+cq37dBfGZzHd4eaGiLJYWw5alnKN/KXKT5sfzQ/JJe3wDm3Idt1n5PinYYSM4dR
JX1kQephL1eniAet9OBOD+ichstnYDSacCFyeE1oFq6dCi3poLuy+oJ6tHcFdABkuqZBKagC4EGa
Y+vHjTQrFiEOpUwRInWUpNsg6hWgULMNqxm4AbUm57DC/23BbWjm0RfU38iXRq6MndWDBI0gKt5C
xrkcwJmsEmP27xLmG+tilcudkKqKU369gxtvIPmdNZLyAErlGbqXD2yjq4UDeuGearyDbJU4rgLZ
HwRiSTAKQcU06eJEnkp9lBeMNeDjGIP2URg70izmrGTv0468uyXhyMDo5fzgYNEHXSYpEHoFt1Sw
E4OdleI3sqcSYsNIFbp44CknY/V0mYlfvvWFTD2OlQrWAm0/VSufod3EIvDXpirWrfbV+9o2jmW+
E5qSLQxPWMKgBdjJura2Pl33dBW2vYh2cbYfDwJ1AbbPivxHWKSF6FCY236CElZues2pTXvjULLi
DDq2sMl1zrXC3THsPutH8tVaS3cu/B+MDGpcc6q2Cb0mBByDBhrcfYaYRk1N/hXPUsMdRjNNltr+
Uwy7bBOHZyBruT9Zx9WluNC3KMRXRzzrlWRrq/W1GxaNfh9siJt0vwYUUdfUE+YU+rVN89Ms/SCy
hD7sheerV/ywXM6S2KZpnEfAWF8zK0hL1fSaYglrX65UQEWdsxRydZILrhYpzG0QzeKSK0hNQbly
685olHnGJCDwICbQJtDlD+Jo+nigf5mlQc5SXEzVxsMKHdNeDnAAicrkf/2DD9oHO9SBXeQxK3gD
Zanr9WRp0yIZXjpGHo6YcmVmZ/fQGuO9U7gLajGEmbFTumdT25V4CyfG56rZfdM4XoFBAwfXGky3
5JekdGHQYs0Vqg/bdVfjBn04TLXrCkSRfEzvai47uL896f1KRg7iFCa+FzAvFLqVFbQhqWte2+w7
9jMQwXjLoWF96vBgeZQY5ebV51DvFYsBKu7nCx+R1dsXriZ5cZ8DlBFkH9seyMBTUNbeei6XzsDT
RtgXPPXl/J7UiI2Q6pSPcylGjlzBx8H0zOhhjNHaJZWwzVMbMPQa/S/b/FIVbTIdNsbrjB2b1mP6
cZuXT0G1+YMN2V+GW1ShaBbsm1Ep/SxUbJInPjjfDw8WIQOM/JauAqZ0KttEWfF1Gj16nfI/ghco
aFU0E/AEqrAL3JyNAVtt+YD21J/e1w35Ke3xILQh9CU8qFnW0nnHVMad6z/BV+mTxH5WIfkieYWn
xupC8Hq46r8p+SsJpse0FlSSF9PQcQBg5qf2GmN9xuu7OtSCzMqAE5Rr+g6wuPh3ng46g14smkYu
KJwOuR/t0ys+6s+lJ3xy76j4x24OuESXYdIaCfqHHqoBAixX9V2QLVr3ntxOH7zndlEFF4XDe8kp
nm2cuE8iqP8E4LCz8Fw7SFBU9WjbHtDtdz6dGhYGxsguMuzOLQ/rOedBa321Be0/YZzJ+35A7eoK
kGwCEkOrmxaEbRRjPCGSQ/MwCBbKQP63+LDIeucnDxAjqdidt1qil40vXIv273adWi+tQRu8W8M+
3P9UsrNUn3P2H9/ortzdnhwg0ier/3iHOYmHnzmFThTiU2Aa6eCjbpHz7v03057wdZ/7AVCjGXT8
mUF9m5Kb+4ImcWR+8Rob9qwgxtMSSQMsIQWB+UX/AWBbGzECXuTbli+HekaBMOcT1X68gziFl7R8
IAO8vuCvX4TvpuTypg70o8Ek7yvOoVGslgA/ExKWObwrYWipsUyqK4iMYHuRY50jJkg8wPgaIO7M
ywwApp60FLQKoNIZc2BN8nD2qj46VFrwiZTDxoPhToh0gwDnAvC3k2PuTjuG+kWkwdCz/47Xv0ss
m6Z5A8j4vApi55lh66CXXdg5q7vLLC/0lZoq/0HrTwIx0dCW2Z4Zitc3w6pEwiErQZD2vawlXAf3
PNATDTmHb94VCMHqSDBcKQCxTu70a5q2o4Oqda8kNC9Qc6cuqbiS9vn5927VO6lvr0MEpkHzRH4j
OWVt2Gw+kxOafu7UVodWW3ddTz3etLMccayTItO/XuZTqf6VEkuVQxnTMjN4jN5g0XS6VDtEO+3/
1DVQIGvXNsyMJgo+1Uwe98qGEcwQmM8yguKuuiJwVxjFi5SwF9o7IIbKO5ruzHxGgbw/r05pN8P7
XPe5gFAxj+O/pgbVtga6NfuPVfEGF4oYlCsuvS1mtmZ3A97CoRpIRL75lGDuKNqk6nDCvQsALl4J
c1Pcu9mw/YGdf7K57lxc0Od2MHgOkjbscoJWivieji7WDEffJAN+gPHytTu73AXbVmXxW10tElSt
LZcHSLCR3vDGwW9QnPX/3aSrZPdLCkNqvTlcMOPnx8mYJxScDAd04TNr5vqyJsdpQRKski56UXq6
FA35d2UQ54WtdT53STstWTPUM+Z8RfNV3/c+XNrnI6maPCujwtYI7YuZ8MzOf/cEukCzNGELMvdS
lKzwUVFq4hcSrFMD/h7Lm0YL5Srcm9ZUSJixnj5KfOkIsOY9jwqgNvOzc+BsDfd7Iv7hG5u5pMQk
oto3T45TdzhwYF0NEuS0ZVlVO+hB+nLlF9ro8TMLvJexa5UJd1SC43jEetiLty+w/Gp1bUWGvuRd
1gLinQuK0jC31DsZGLGHjxJUpXUgxgr/QNw9msqSCrJEq+qDgJDuSJMV4nQrGqi8uSYUbWYgmpWr
eGggCGVCLUnj3WCxp+06sTnTHDR5JqkCE645qiaWTturI8DaWU0rkS2HrZSn3Hp3WraM6EcqNM0z
WAea3vIyZcSTh4FEca9fy5736dru4OkZLcY2oHiPceJTlui3E6zF6onSbx//p5x/cW0KmgNXKKNV
3Dlddklwd3L15L0lR/xCbrGK17zK4y43z2jQfBwZVE96PAIYe3eFk0T0ALMD2qNS0UMvFNb7I/8Q
f+nQQP7yQ7E43Kg3wt4Cb886Xq4yDCxZdVILHUI7XF2gY2lSeIjGW4yJ1JiHb/oGoO2QWG9Nu2yz
h9ijPptpaG+4lSKoKxZSgpkFadEVDkbjPrrPkNNytvk8jU4r8PgEcbdKiIT/9TnY7t3NiUGS4w8A
z221xd5aSu1R3oSrlYM0xmeZg6Szk1c77qtYRoKZ5Dgnlr/lTZwgBOSQ+tDdQsnnGsTb2WI67Q7w
lwsAfV9Jb1eedo7JLE3ZLQXgCrmS0wPmaUp6tHmUeGQRHG8lvH5crjilYAmCZBJEXzn6wrz/kNpq
7olJDjB/1gBcJn4RY317wd5pYwnVjxF/zTMlOO/32lvHVHSDQgIeI+xJ3Rm6rwzzieqIN7+5cyaf
/YiWl1rshW1HsrAd/alf8H+EaP84lwO1Zs7ujfafJfJ/4Vzykh4Fn9Q8nKgUNx9UxIrod/bHNYI2
TJ1i+TRcWADKC0Hc3wp4Qd2k1EAxBLd9fWkLN+EQpmuyXqrObG6WxNXOJ2jS+weX5P//w7AwAqzg
DT3z5Vsg5iA9vZLfdnJ/PR1LlmLCUgTCUVJi/HM+M5hUhFEntWIC0s7rwC2MjuJM1LiqcRqbkZDL
wwo/Rs7tKqUhS6+Os1QDw8WgBZZR4KqIQfp7oUwGWLobVNxGiIhzwQSBKgjViX9Yn5HeT8ONRiYv
56nOLUx3hGGmO+aTqB1apvm7Z49tPgdcScJnT9l5QVBOSZqNSsHW3Bg50brmVScSgWq1jV9m82mi
3X4BceL2M8JGKDpQQDKfjk6hzeOFKYYe6ZLue/5ndjZx5km1U9U7vqHKmNIKAtyRGWqjRdzS87xF
wJkqwTLxHwBJBe4KZj4VzyA1uiJKYOMGSgOqv+T80GJnXUpjIbX35w1cAqCMJ1ne0+1WngvwkkeE
1G5baPpRuQTCogsTRgpT+KiwaEF8uB1YfHMbQdHf3FsZtFgOO/02hw4cAj2mRf6NTIpqvw9SfID2
KXq94DNNFpv2Zl3E/O9eG3M1a2hZe62J3SCLKNSkGIfnnnyBdL02af8gYJagG/DNqljIuFVxlOJN
8dsHdMGPEQylVgGKyqm/0lKog5KkuGSheglKBq4+s1umZD+MYK4u/MhDiOTfP0Bj4zslqwGvM/uN
wcqtkYf97V5H86ZUaAhBaX4P8fdQqrh8a6dJqdtoRYqbKB69PlAxsjAUeKbuNyGj7Xj2VPDCNnF5
EOe3xUnv5o++BBXhnT2E/XOdbsFI5z3nWjx1Tm86HO4JRd3CJ39GFzA9piCAqKsC3hILr3VQhe3j
JNZ8L/NhVqccJQFyF6NBcWWOtuHXbhL8YdL9qVDO0c//F1Ym2Emf7I/KQdY1KcRvTnNtjmWvPaYN
8fMMZ+Gvh9zvf6BKXXEkije2FHODsDyCxHya6dyPL6gfMrNq5crvG7eorKvHtop2b1edueh9lRu6
MyT9MAMbonv2IxPwPk9EsfgDIYaJtuhNWbEsM4KPwPTltzZcbCkD73cZIfmfx3Z7qdVT2JMYJGNB
zPqg6JqB98IFXlA88T6c6SEXf/X3PnRojaors5fFrr3WVjbyjga0iQcYpD6ZaOG7xoJp0F7g544v
8mkziT+e+J97ZK1aTGtnB20T1TJz7JLUthPJs+2p/ZZzEXAbrL5HEBTghCRls4HhZ+9guDbaLdkj
55N0Klg1k59DNvzjRXxmMm54UD/xycZYqQec1WadB6UivxEUWY4vQHyBDqwqJmcyBJiDeEyGMbtQ
pcSsCKgzmdUj5qICpj6dS9fPOmJBYTwT7dwBtyRGmzI/T/EHrA9wTDlmRTBAG5iDWG0rVT9GZRqP
E6QeLGmlLpYP0eca2UbGXOchZxsfByTeDm1BEA+6N+/6j6o1Lwl7u5U+OMB2U+ZNVyGcu30DIYVF
2yOTEbH0avwD6F02Vp0lGI9WsMmoejD24Arz4PtNvkV3R8KYHzEcdSjmpux4ekF/LOwIrhRx2zVE
iHYLHmgZx4WHtnFQpF+ZzJqU6reJyP4i0slmF94g4pvdv8FwGOEspes+NeJW7w2WgOA1pItzFYQj
Z2x3lVzsW39tTwGhEybA2Sg1aSSvvtaNQYtzfLr/FPo/FLDI1RY9HV1IE9UOULg3+VZZA2h89VFz
/z+J+Ma5yntITo5NqBUVlP0TbzKgG/WDmFsq7/VLYG09l2Hp2uCrsTHKT95oWaOe+8IMnviS8PeB
mnGNPYHjfFKTnk6FKVoDmec+qG3F6Ldhs/6M4N9kRkRaTuyespPgAIOoRQ3yWKMjfL6cbbxnzS2Q
mEHUvugDsOyZT6gkS9/cUFc/Izg1v1Pgkmcux++4TUx1u2uYnXvZXfzR1ILts1ae3go9SLFhPck4
joNILQ3+NvknMWdM39B2SCT0x6+sQfIN67wojTIM6qjFImHjQyjMaM56NP8x28QEWRRMJysX1leh
rZL8MJ7AeCZrCxkHTV4dpPwVmcW9bimX+JtwGJ7ek/GmcdkCf7RmeEKv5Wi1jXxTd8JMg94UORhO
7dN9NMwRlRWmcJWU70qd/bzEHf0bXlIenOVpvmC0wK53ROoS8eVpqbiZSo24N1ZltRJNXXP9iIzZ
06Fw97N2AzGJy+mZZAxjEB4HVxerkPtQHEfhVGqgUODFa3DBAVY0fbCynb/V7EsuCReg8N2k1zIG
tl/fe4fl2wP/UuBRAZWWY+SHfB84St0emAHPk5KIejeYXA3entPJP4vNt5x8wVj9kCiO1mAHrRJz
JNKbRkshyH5ml82Hkqk+hukxBRzIdY/mEaV/b2iskvw7ZMqByXjLjdzFlpmIKNNjSwTSTwjxsxN3
GowYDLdOklDK8UO6ueiVH2IVcLvh0o4QNhrnUuUR0IpWI4AYyqPVJubVOyKd8GpRIMwzqTqA7o7o
3cXLiK0aNoXLEl1J8uandlEMk+Q9oIHcMLOLANrFdEGpERdniNvzLhUoJiyFSTALTBA2gbqFV3rp
NrA29Iwm3KZdnA70OBAdHvDx4F8Ts0oZL2AdO9oC7DvVK0CU2/k6qI+LfPEv0GAHussst0Y5Eknp
nX2skALf2C2XTe6rPKo2ybSVczfRwI+k4nCsZNdQdP2ZhFBn1lCX/u9bjaSZuRJy/nRbZKy5j9ty
R6vk/DARY0kGdFw1Q7nT74bS5agXfQmZ5G4xcbekjXIPTcFDgpdiQrCkd0uhfPPVONWJ4crEulnQ
Rb+53+baL5OhSSRi9HMI7ccKA+yEkzLzRjE87OCD0VLO+yhqVsuIrov2+8L+5LzEztfP6IrE3rpx
7BCLfwuic3+0GueNl0ukY9Ess4DWalyo8T7xjOxDsHKcTBwxqgis7cY2YERK66oC0TeibtJxSFAU
J66WI7EXHMLva4L6U3UXSG/+W6Mbc7yClaNvK/vFuYuB03XVYysx8Aq92BmYD2aQu355NmFlpMCi
I9hNPSkkIBgPv6wnxY60tHzc4mG8JLAy7V1g3fJkq+Y7XIQrUW7SweJaV/J/Bcb2hAaEoW1NeHjX
Nra/dE5kW4BZzO80uhZERVO+iOl5rnvTux0tGyJN8xHn6wys5ZZMsag/o++eX4K8L086NNuafEP8
n+YZUhAoj1TCNWkrdWIZXi1uXwkBbKXr89njLW7vE1pHjyaED6Z7VjOBN7bLX6PAImxnxEsFUvIs
2AQCfSpLAHyTIMIyZyopWTs5R6S2jowzUBixPihv3YXJErhgbc0sd9ODSpc1dUx0ZHm6vmQZMQ8j
ovFGJVRN/PSqDROlLaSN05T6afgpn+swKgmBaq0QGmLeqKaJH2dV4PnH/zZYomdOw6RdS4IW4gOk
C1U4zNRszXhoCqk3aiMTgV3Mof4wY+2ZlvFctKDmbmzyH5qEiR3yMohuhr+4xyU/MZS1mYNuXzvc
i8E2BENmY1CtTD6ZQuafDnvZHBRkiiNV6L+e7EzA0Q1PmGRTp8a9zjTp7Bj1E3Tbw+lma1Ws99je
TmNh6m8E23EGfvjlexGZRXw0qXib2WVRRdiL3bZKAnbzPdaT0nJxrp0Mw6/wcfOjJKSp1mnnXElM
lKL13g1zu7jgwln3F1CLI1LaDcJl+YoqoMipDgz/XOKfdn2BU4Oo6kgXPnymFmlavA+TBXi4bgP1
ekowgCQrCR+4Zt35qDbkm18xij/MS01jR/Kg8EbnusqTKiE1fNvAbJ7r6kyK+9/vnm0vU7tvlIan
xeCLp15oxO9CX4d8mZVOBwadFUT8+Hsbdi1YFC6uKjEiIBVKfjPsTo9lPNOiv/2ismAD5gg4G1Ps
YwPES3xbx6vqtq6Ane0sjqdCrSC4UXD8x0NDOp0mWofsaeIqaWDaksQyC6lHgSukHOWXHDDbaMYH
Hkobaxtxu1Wn9ItoIb2IaL43eWvouUHkAguRxsdJLYpSaDhgyrlZ34j/MlOQ1o/SYL9ky4HKPU6k
ilOPQcRPPZ/W40lq1jswlD78muLW4/Ck44+ZPCxYpFq02y5/0/ohsdX19ikxZzyHxIEdbf+yn5wI
QGVuBHYZtvvTUaS3TKeMWd3dtwP5/fRmuMpLxTNMI2fDyMC33orB4VNFRhv+OwY5D+cLfZkUi/hT
POETRc/PiPzcLN2lwBd/MDSCFozSmiUfUEPSPmyFWatffJx+idM9Ck2pP4KF1FjQwb5W+bTUe5R0
DSdTmjP4d0BN3id4GJS5S/vSJbHxS9ViSLHjsc46rc1UdR4j7NUOAMabk5c+PWYx02KzuRjjP8L0
RV8FuP5rrbr4RbBJseI91NsvksIhUiRazNSIbJb0iun5M9yRzz9AEa1P+lpk4fkikojHTBq+p87K
ZwpCwnhjfRHpt8LJMXdFXs7zxDrHOeBx1yHdy9DZ4vOTpnjQQO+nEd6CPp+/ZaVHv6EJUAwtsHLM
MWyabzrUxfQOVS2IhkaRRSBEHGM2i0QqYhdTHtXLeEKTNpLRum61b/NRuNHw0KhN+0FRWFcHMJZz
5WaL0tscTcjK2xbydFo7IdT0WTGUqEuXAxdAuf44YUZ9v1UH4LejhNOsC5N1QM//YkU8XGcWtS5o
iotKVYdFGo6OUvhL0x2xjQGFPx9KYtr0VHLx2KDV8ih91Pw5tM/nKnBw9ASwQY1nlXu0HmbD6drs
mEZTs62Zpao9qwi2vY56x5gkmyhPGnV3E/SKrYGlceD3HSkfMir2YP+qgEpqkbkHu7OPogkzzeBP
chuClnWd+1dNbvf7eRaSOdV2Bmpp7JONE1hdWTDLekn8/wX71a7OVWW8rwqu/w0GW9eqk+qojPAR
aFcceFm2TYO6Yjb7V2VS+zdhgf+RBXsdA8u70ontux7kDkmQmyrTg83U8qXXY66tUqKFboBJslGC
RKnJKLGVGO413tbJ1gXcwnHXb9Emc4cJhBDXvqcU8xcgqwvp2ePmHDUemsMGBiQ7zhE3cQmT/wHe
k/hk7le6cwhIjdyy4jvENHFEz6qnMk0u/kIHEFFuEmT73qdpr9sgouDFXGDbM+sj3HN493iByzy6
4Mp8wSUL+CUbzUBGg2zUt05huHJdMufe7IeQTq3FvRu0t09AymO83dG35yH0HpAnhhhvEu7lG5RQ
uAalLROge3muMTR5XMVJkuWbnSAJB8P4DU1/shOJCjGLxke0EU7RFCTm4cPkOPvCEE4Vw8Yx0i9t
VWIN/1H+vwXTJ6mftU0rp28Tzj3AIPqHwzSdx17nhdJ0ZK5CnQPJbHqDtdBkCPyokJM/7MeYs8i6
vbBGz4uChAQ9R8p46GtkyEOz26Io43lz9wU2BuUXvaUYD8ePs6W9SAMCiDL62FSMHzneihCivpPK
g+1+yQ6eoj0H8HZ5DNp2tliXHmcJ4GyBkY1oSUZrD3Ww9kfFQcjOpI+izukjY83TXX1LSN8VYGOZ
ZnZbRG9OkP+wzVnvxaO1xtTz/xXk3qP/xATL9A/9aDhfOvlOHGN0Fy/TitT+KwWEuZZCykfTJWM3
AThIfamLVPLHWNfDvXE7JTnDw8dAjfkeYAZD99KbZCtdAFietfFH4fwdyNAwnvZ8bBjkyB3c5Nwb
a4aqKkXtZf11SZ3F/yWnRqXp8p3nargIm4D5MJWD99HEIwq6oymll1F8Za7bmsASs+YAYwOIPaeT
A81mAIMScTszyBDqFHMjM6tKZ8ujTguyXmReYb0OeUyyRYROrt6d9TK3TzJXVBc0aEnqJ+j9EkNk
4TJtHUMAmrh7uk+DXyBy6MoOdkHtDngCqjGqR7AvmggrcbBWelHfIVjPR8+WkBtcWNE91QvRCNSt
V3GLbzd3YuZQQwWltv465lL0mnHBlubwx1drh+9vKNwkW0GIvD97V4box98w+obsbrbKaLUZw0y/
EQ7Xbss5PG/AySqyIP/Czu903IL9rfnpShhYGjCe94uKjOBnEkhra2C/hr8zJL/QAPWF1Z9p7o/Z
m1LvoGP1+DuHjQCZNnHU/iN7rAC+BQAbQjBsJY17YPFr50TSeNeUIkQ5wOtxQTtvL3OpBwm+QgFg
mbiDDPnBTrhJJJs6ulz/Iwn5OmFYF6GJPFiZWwsPC8E07ITSgCz7uzRPQcvvVdbk/kZ7U68PcieL
JC3F/7hgvxBC6G6vNItSL/glZbuv98c26Gw6fKxHAdTEOgKqJvN6RfxMSMddpEAyzp3/zfsHWhj8
c6S8VKvpzTV5mu1+02WprrjJ1LpYKH23DPuykFl+qfzaTHmSf5MUCjF9sukUeLpp6jJjYvkrLxXV
L9PLVYHW45n05MFqNWfrUK6YqAuhclfkGcxOQpN71mFWZbZytfh+8TmJkwlldREU6rbZqdY8t0K4
H6I9mDtrDih0mxs1stoSGVBQPaS38HlcKgz02Nh4OmEJnn2FqBqY91Xw1U/tVyTzwjsiF/H4F6SI
uIbVU7svAgvEqPZ9WAnOvTu8l7AAuC7i3sCsG5AZLHnEuAQQb38u2IdZljXR8p49flqX8K9cLVmk
aabOIexMzS04ohvsQTBKpDA7PNOyP078ZnyKNSRnE6blx2iNiDFlcK24K8OYrx3/CnXz6fp7Obt5
yq7lte1p69hRLw5LinY7OZoeaxa5NBBHxqI/zumWyJwwSJv8R6e+dG0k3IpHM1ofNaiXzHhvg2H3
0wDio7OJImGeLiTyTO+5ATp9O+qmvBCm9IcT0uN3hyW0jUXQjrEvMzr5rB+zjER6LWQOyzOh/zj0
Hey2mAjfHO0mnrH8wE0OC/H+ovb7gwbGI/wVAU6vj+t6KIZLxewsae1FecjwSD/B3pUzPnEgY9t8
7bk32ssAzmRY8KimBMQk80pq5VQXQwrg2NZGXj5RBUs9ekwg1G41u5JdB9Ovfouc5g+xdljHjhgP
AfMHIaF7SnE+yklC9aijXavIVM9Pg0Yml0ZR1HAokPmVHfri4Ame+UdC3L0wF36bJZtMJ5T//D4d
p/2mkvmfTFNA6MfFLY6cSaq+j+S/ZVrOQ1QB0Z7xo4oEUtpIwVvffClytpW77IolCX6LrqB2mvje
CDx4+3aqKtG9/xslBd531kZnO/5DU2OW0mT7r0dCRwXRGwfkzkUQq62B8ta6pti8fw0EycvTPM4N
i7iGEDP+eGZHIS7BjGeqj0bxrpFNNMf0M6trhTHnwx8/Ktx42Tk/A+nOIP3F3uGReTBFVTHx+fdA
Hn0xDsXaPgwJWHuUx5HBwsNWkuvm//d5nSKBuhj8NbECnsjHX05NCPftkMjJLaI61fUAFciqmFDP
OjPbYQhJzd3yOOOCRoIYpBHU1uMRDxkUD/npgerEdbykh+ZiBZs6ZjYkW5R8eAsu4RJj7Nuyp/p/
AiiGDZdF8Uvypu6YvFPer8dmOwNHoPyiUJWG3yyKGvWSQWqbnhOyr42XdesjnGIxvjg1gjsjz2lE
281iKuOGVvtMEbglqUrSvqkGmvOpVyvEBv3vmybXlq1Q3DaiwYn4pONZ3aayUkXV7x/A2M5Sb4TA
0kkbQv/dzpx6Lg1mgC/en99JFUZCEmmTxc/BVo64x3UCD+07xKMNtaZErBAJbGZ1oySyh+4ZTeY8
DM4LoYABqeLdEa04N1t9HEwKyEqPPsckYnRFV/7aVm9/S7LKBH/Exn0r7GATRvYIw3AriH3W5t5/
UktcKC61ZZFllomxE5ZCj6hLxnzxgjjhCV47BJzXBZtIQRWVdXuV2oZ2N3f45lxVKm9DysUS+eX1
0/SjX/adS9wRUcx6mwKcFPaNwcfFgUYS2kiJbUsWk+UzT4Wc+Hisu+zKyumSU1fTXnLbhHdvcKo0
IwxXxmYV8TTaDtvjLTuYLCdT8Tjdbo8+rbtU8KLQVjfMnvLHetAn6g90DgieWgScfE7NIPObnNC+
RAej69U9AkVgy7DZw61oTwnqBZu0kTCsIlb6TlvCMVkwEZQsT1MnG2edLf1C368MD8VcVGpZFiPH
orU4gMXtA5leGUaBT4UFP4btzslSf4jnwEzQeTPC77MeJWGNTCX5EvZscZjbnVU1LnNP35DjiVXN
J1KzhGX+kVQW1+BpgYr5Y2u2XZVkkN1G4b3BY3Yy+Onkrxif2Picz9hqBSB50yGs09fGVXk1blyX
AEtYkCMV02/NkM1JY9nPSR3vj3pWhyv47cVmCMWt59UAAqal/2AcO82SKQRdiHah3ib8QpdnYtwE
ui1o84vb4w9XS+5lZSofrogdm+kImXBGRzrq2GTdygP1vM0RtbHGZC4r7IM0bPD4uKqu1r4Esq16
q5F6HqCdSdSYrqGZ5cfV3KjO3cqis7qJmGZ2dtKQl1vSof7jAlBPMD0rCgbpi3/WgnAyH/TvbIAN
XwKw3hMd9lvksaECXn3qY8Dfo4WkIps8qHC1KSTSsiJ1pjCy7b+Vum+oTQAEBC45WIA4si9pB40s
sYJRIe9l7qkPBFnqkin2Tn4icwKfxP5awRRomXl2ibrlgRNVxh7pxIH+3d5jOcCX1xfYAz8XJi4P
BGJ0gIlgXpI2GzxpPgDg+viaUewdlFcTY6nCQ1YGsniIcSdTz97hx3ivfaw7yQ4jH4j0zp7Kj37s
pvlJvfCDR4kWpK1Tg93ll/hcioNfVEM0kDB3sbcN1ximANp57T7UZ+fkvBu/BdA0np3w4GltElNH
Msgi02rdoZJ3u8JHv9erJkzAvKhNWDZ2NXVXiMuJixoXp2KJzY6PwdKuzGiImLRNV52S9ihjatpu
e2sParb88IOiCdsZVmKW8KC10FF5LpCRFx9IUA2C4E/+CsOOrXBFlKIB3Ovhtd+Nw1YLEIr/L3/d
cHor01gAZgWOWi3QkuafgCFWp9BYCq8Y/rHqN18UL+7vzOTuKIu2taCqBCEh/XC8oHpyM3x/CwPh
JA3uLAHVj/hO9KLdyEuHJkFJbn3h5nHFmgYRivzYqVE2T+ZWbgjS2Fx849F696gkXe0KZJcDIU+p
RGvUG8dqqZBD//s4LD6paIqdHH4+gOphxqDrvUcGPjFrX2+OoZ1KD8XDJvfhvzmwj0DcuGkN4/zx
9MZd9sT4dHPCzNLc6a4kapNM7NctmpmAEhAh2rHnGFcNMtlkzLqs73agvHGa9pfh4xCv6PVIIpur
47bGsw5YW3+D5DwQhpHU5NDsMLpCPvdaLu98F/xf+cLAQNtk98qS5Lha6dwHO3E1gCioGWoGqLwT
WdWBOjbiTeYizr/ysgHV4f0seg1y0KDoO1iOcDo6bZomkhMnBjAeT+XjMCPue0eGptBHrEjiuKOc
tk0U6D/lFIcfqwDT7yctzjq/qyeFOzvd9bilE1y08dolnCTV/AY3uiQAPADB0COYudjBgLdmOmxK
yZDOSgqj+VgSA6N27KhdONCXyeprTzVB+3N+uMVQ6/1ubL5a5dhh5XGz+def3LQ+ldnJZpiXDsMd
0E17FSgBKNBB+RykgA0mBTs3d9hsTJByvQGPKIV4kfmvTZ40QJGvPvh4ssGTnDRf2ZDDCeQborHn
Gb1g0ozvzXv3PWL1OOyJoaTb9Xsd2u49QwONAjR8JGXPmlXthOmb3mvPWl1peWLWm1ESXPw6G9pl
0yCVA8v0pFQHLBpJmHQ2fBwuVEEBK6vHXIiMP/YGV2MCg/RgGrieZC8yOovyL07k9jfhoBWd4n/J
kkev5dN8CLiOnFujUG6wTKmb5f8peqwJctPT/yDGAkyVT6VzPdMaHMUl1fKhzovfZ4iMIFXt85kX
J0m7toB/UN3PxmYkzBi4axzvo5MdPdY/FzIamvD/1fJMfS13LeRqHbuIcBvRRMxe9db/uXN+UJgJ
3NqGRJHYir+LtSwTIZP+A7a4ruAZ0BK0k8VtYT39whpJaQ9UvPN039LQ6HE/ekJlkB/RHJS2tSaM
evYY75s9yfloBM3ebzbM4CzKSEfLYsp32T+Q9R7nh5EqmdsrOO5Bsw+tN+thdjtY2FbbgQt89hry
IDGfYmDxiLkHAGLGlTjmYemWjaAQ9dyY/H5AnM5TvSxt9RX2n5iCD5zbH0w7UpaX9A6NoO1pfd50
CgeptmSI6QQuaagjsogSjb0GPvg0FtZiBYaOSMAcCMuWamzrgMAD5sEN3V8FekJGdJcaUVSeHmiA
OG/3BcNCo3TyW1pM6oTc9NfwipF/MBb5MjQje58zS4oRxDaI7N/s9eKfdW64IAGEdP6ye2CRvvzZ
q5zNrYgL9bUtztf8v4DYqkPUK9CxwyhhIsmnL6gG19GTY/4z4BUf/Fmou8Ia43CqfxXMo1vu1Cyl
gPcLkDJWZYaUJ+CA2Lj6mYNOxY6045CmPe9iNlkOf8POpvyzP8YJRa1vnQX7QoYtPirbTKj1Bn3s
tfyKmi8VlA1n1mFkVp+gp9UPcoGQI4N5LaId+/gSrS6iauPxRpQ51iOrZTslXVp/CyI3lHDLfuwC
jIWqHq3Or8aODLo+Z97wqO2LWP8o8kyFiRLuUR0+EMQEh4ZpoL9PcId9tZnfYv2Rf7xz/NsMxMVZ
IHU2PVhYdb17NFllwfSbBWFuRZnNab1nxJTE95E6pyT2sti52rgN++D/NwR2Wp/HdDg4KYEeIDh7
s71aVhskOafqXuQXlqnoS4/YnUvahDP/9TndOdhbA6HXx4yyXcH63jTIoAqj9rrw3aTbVsemQMls
BvdDB2YrioJtTmQ0SjFd9zm6XyZegVxR4JJikiWTlU6dW3131WNBlYQ/mREql2gWIolyL4U9OANX
1Q+7xWsYsUqX6qdEta3fCB3URDKzzW/8VdK9SIDbvx+qgR9Z/l1L+JJ8s/732drWrrU84WLlHYi8
gw3nmxoi0QtX6gERSKG3Sq+Lfsf839Dbdces2UgmzIV/L6ke8vno54mO8kVu8vZm4adfKxU5/Gn+
HqtrAU2mzR6gkyZ+bnTHzGmf/u6lTFEtvjTXoyY+77sI4iOhGgd1sMi2ranSLwT0Cx+PD2dfdCNr
uw3G4mYRZsInCRtQPerxZzWrHx9kkJxfpLFlPOcGgVbJHi7cfiO2xVH1dcM3SYwusetJ/vz0wMgF
WH+KF36ZKo3yiqs6O8C0H6SwkrtEJ2PHnOxLA9F1yfIheA4QgkfZfFT8JOG1K/wKFgTOJsyT2Mde
F7iIr8vqsgBGtrn8+nwEgCvYN+QvgWq60SkGdEdRWieP1Jqp2uCqgHn3Tbub7sX2dCcOsniEh+Xr
kmEZzGq0OJPkQ5A7F8ev7TxRTIDKiBZbsS3P/MvNrlJwVcxCW3/KkWIwwcRuTcbeJgMLM/SxCqj1
yQHq5Gub8bNhwy8RMyfFeW/4zSdqM1p2YDkILz5jC+V7DLbpVbFSrBOvbEcx9mV9YQgBaMuc3DNM
u3xnt126aDVsKltRYX7MYsaa69c67QwOAIiWW5Up1yMVmmhfP/oMZ7KllW/9BVpvFf/pQH9iI7ya
wOwK7HOquRXfzPpkIWXggNeDiH5dGAPNon4/iMZ9RkZznMp3RjytJPk7e2brKzI8oWuYZllIKWJP
l5efRYz6GVOtnly9W7YCFckNOGf+VllWxS2t5gOJX5pt2MF0pr0xPYU+OQyoSeVuH4X1smZy5Z+1
GTLGIcH5Zl6MwQ2pLdfpJcaJn816AyZlDzZKK0eSYrql8y3O026Zflux44ZDcdOv3G0bas+fc5d0
7+2O3PPeqgX+cxUyF0OBNxQdHtc/XehkmBB6l10Vs0m5tvyYLIinRjMyJwdkp2YLYR49Z3YFnm7o
jGC+L7XO5B4AUvIcBXrMOjtJ1PYYOmpeyn7p5I5E9S8bLvJo2fDLe9BynrOtzbebmEijIHL3raMQ
jzLba7odBflEvSzBM6wY2Jy7oZhb2U2BMicRbmJDJtMwtm2WRWdrZNULjSrqjWOCfti47b5yXU0C
cNz/Wile1LJ40r88naYXqE1UK5ahZWHnnPoboc66uXdyvCUzZZDp8s9uFBx+L8mt92kxbRjC4ssf
Z4Xf8sF78m+6cTmDqaGD+A8Nm4aiGF7FFZmm/xAQllQgVIQxIE+t/Fw5SXv07TiKqqtkbKyHLRXu
WVxUMZBmOkjF82iF+VQgY6hevNvVAsj9NOuRL+q0H7zHX6o1heJQ65msCkeYFPUliSDPdfVPFV5E
DxyInxvivQ4SwOkVyEkSFvBmDruxwWB3P7w8kQO7J+zTq8wJVEQ7ue0wOa5yaa4jzZ2IEUZMu5Fv
Pe1fb/ciFypnbZvZjT/5L/ygCo2k/UCmH8NKfMxB91CTsi1hz1pRrrSKMe+CW4EVO//sbvkySD+h
uUibk+RSctNqyIYTiZ6BK09igPQuNTQP1K4MZHRuNXslIjGbD3fnIAfCwqQgVLy1xCeM1+iN0Yak
KI0JAWVl5n/OIEDWbiR/UAQhlev2iEvOlVBc2Na8Pa0bj4ytEQYtz84AbIYwQn5TuzWpkYI0vFg3
dklZfPVPoiwk1ft27wIYWlmjmDG2I5QlrW31RY/bu5JW7iuLpvS7947ZgFp0QgltWLgjKDRryIer
vQEBxZC3e9KSK4+gV8ppsO19E2vXtYf+2dYkcY6DpgCIJwZ5XRe01h2kkISijY1meQ3a/c8+/SQR
eTxWZSkCfqwCE1kkLGM29BJ/7OPDy2Ruc2HgxAAMHNTz75MJZoTNDF+zyCNxLhJ44Qfo5hyIImJR
o6qtXLJWuEL3DDnuNft5ru/lLm6TT0O/rvFIasPhIUQJ5a7xf1yHR4gSXPS2pATHffYcYcCpU0BE
om7xi+XktowVZg+3gFLLPl5urOxwDfgISt0HX/PckvAAea2hZ5TpUH1dWgy4FtXBGcpvOEE3S3Ay
BHhK6bdqgn4kCQdU8dHQ8aFYtxYTWBfFEGCCo4ur2UmPdhkSR+uM4o/do3/MGgCUP/EncFDnpxPI
OXniTm1ff/pCUd0ssCyto3GgDhHTrMNzsDK0DYi7qUBY5uBSfapS7mIbcDiHc4q+rzNi6OBzDGdw
a3t5TMz0CMghQmjv/gadw5V9q7DgRDWWtNq43oHUmwuN4rjdo3dkZ/RirMFwhusdxYiATvYzsxFv
Lduvay2tbBf5cVyxQxlsT1O0cNU+ZqDkj2yRxV1CN54NSFVdzX++f5xZBLNCzRuYqjfcjmIEEs1F
FdCWy3AZLLAguUjJTeal8y5omeQ11S7lD3PYJU8fVD0yrfoDxcAP5gI4pOICHtFiyfR3Aux2lUZU
0oB8urB6NFkUCIbEXwU29hW4OFKYsHKA2ydUr+1geZfBej/ZDX4DbnWt7TqDY+ltbjmYNvkAhECT
eE/dabzBwDOCzC1cNs1oidS7jtBpQzhjSKq1ZesFWL9CKCgeh8s25MSTUpa/AdM6uT/BIE2bmqKB
F9Jj+QEaDiWPDrzVZ7xbujkXGQPoZOEMliihp3keAcRMsURx/lKHT1CA4RVvcafyvmxU34NB9T47
ubl7w3wLTtf7nkemBmPE6r6KMJLmApqE1sg2EgyNd/3m9njKv/Svsfqw0Cy/jWh9loyCGDQjzUp3
RuhtmIgs3fdKDVPtikBMz0O8ViIX+fhOADA1Dd+oQf+Z2HAp4pCbfUQfUbdDq2YV0PUI0S/Hj0jS
3ng5X0xLMKxeWhVqf8zlCg3LIuyMlA54jwJK9DfpqkeVasos50SxIf53XhhsRgsk9ET87oIB9+x8
8mxdg/uWkFxtePtMvnYhHhgkjZ4A/BSQqvnJbRS2A3OY6jdzUenzStiUqJQw4ym2WUeplZYB6tLX
w96yuLmvKW3zEy27B0rbAb/yef4SGtZzYI8x9vyRx9Fn116TeHRHNg35nkKR/X03XSSvFalBgl15
xZMCwWxqiZ9BeVNH5L999QN+MuzGdAolxw9rq8pnHgRGBsMWL1BIubPbrNerUFuZ1wBepWlGbaAp
OxSocP9GxqGDV9WO0DMhu+zZ9yowQzSYeCdT+k/q8RA66i4Y45xK4KQb3Ca/7uuFFmEl7A1/fIVD
lgi2+31Ng6Tu3PSKxw1ZUOLaftuM6Kp+0uRr2hMwEvRt7JMMM7bOh2qGt0NqVBwlxSE6WgJ59h/m
iGI+NPwIwVmnz7oOWWNVDgeNaeIaGhi5z3dwMBB2hSlL699XJ2QpMwF5d18CMEjLPPkdGK/bXo8d
jydFUbiINM/tQtjdWQnhiEH742UQ0+5BS+IGTkKLVn0jWy3UIbRqTtSxqgTve4tcSvS5BYBksS00
ZVGiRANdw2o/jCM4wqniFeffSHGdgREpL7QSLBjx0VSwgDJyZAT8c1Zcu5BZFTuwun63rlvxd3w9
zLMfuZUo/mtJokmEOZQ2aYX7IByWog3xaM7lP8C492mbFNvHD7HHtr4BnW03YxsimdMQnmxlnXvl
mYAfn+jQDwc+8WEhrWxe6dLBYiQG+zMtSWqfltfDbnl0lTRwl6YgbU0fvs3SArEL3BhD45gT+nL2
t+/cysJ3tyCqaKzkvZ6kiTszV9UXLc4rLFQ7EyHE+PwZ63mViEE+szQG7B0ZDjoo04R6MB0quRsd
Xyra2t2mBNxOSv9RndMe/DCRohSc+rW5fBueWX1bvkgIY7LIFhhXKeKrDeVbZXevyA6DkwPr8w18
5775ZbSdfUVfHBJdXDqf6o26pGEvERdfc5DwHD+0JcV0U+g3Fe4MSTagCzKO1626eLmmQQ70RKs7
5TQHZbnOi2CWO31VgqX+buVc/HbyZnh8AApTvW9aIhhhxrzvPHF35AfFqTGW/GuO4YiZp9ANRApy
nXaHqdW4+DqHHVVqna4apPdRuL7PbWN4WQ/UVA/+U3IL77bPZtvjDwQBwx9ijP0qDpDWHIobFrED
EcqQjGbUurbBcwvdIN97vpY8n1uIlBm/66KvdpGamEs2tX+pvkYTWavf/1sd7w39b+NgxMHgSYIN
9zuy2oF7tavQVoNu3A+oZr+F8ZTGzrq2dNJqS04wtV7fLczZeD6KTt2Yi8Ukm+JAE/K8huSseX8o
DLcLAQ90rKqanzlS9gUVZy4D9dPHbIi6VHNbyGpTmk6QJU/7wYEbLpyyXyklC4Za8bM0B0rPug7y
hqluuubxrzKkMic5Jf4HdQ+zkRB5LHU32GQn/5mgztWhGXwcBAWNVTE2WE2ydS+SHy03Tf+HX1Fm
Ccr7hAvF+QF1OMWqkU9KrbWLKnxsTRB+hr5v97+s9nYgfEF6mLzrGldJ9zMnfaXtAoZ9FaapQ0+V
ZA2drTKHhGd7p5La0nUYzWFmTof1PXJd2XVLBTqSF37ZDZRJflbfH7xxNqAom9C4eEilPt1IvU99
7BmtTV0YUIK1auLtnJ/TjsfSeGQpp/f7KN7gaRTA3rB2NWwbj+wLpuB/vHxSzdick2ehMr1EEmvZ
IxxMoFDbNEK2hg16gws1Vr2T+GmX8w6KE74vZ3OsR47jjO9ah/TmDD98Dyt9xoYPFG4odWJJwF7I
2ydJZGiKdxNrBqUZDYsecxP1HKKltxIv8wH+2ylvPiKqDDxQdV71e7fjw1+IPnEw/TCwkjB0+tIY
xjEEmtR5rFTqTX+uFZcBBXUEwtni5bOrzTXo/GhShbq0uhYoDeMnL2dZK9Jg/kRfAiaYWTRtyt/K
nSlee6FhRcju9KUNEvRwZNNzeC8WkTYN/qV+nldUBw1hNj5t56Cv2JJgznqLJTBEcIySo5wZstPs
LBChRN8k9Euetqf34BPsL/4Xht5gdlOAEV/Ndp0ISWun6zXLaqdmtHCNhV4yUOMFzQivLZciAl75
uV3KoLSCxe3kvn6pnPY7S8U0q3w+mxlWuuyfPnEVJh2FApXMVstKhHhH8ddH3g0Kf1Q03Ngs4aVD
9KpvqiNAEhamH+SLUtCd/CPGnp//46f4iSnqtSW7aFolLAgS66G+4sknfxH2wVSPwtrVRWa2IonS
TmeKGE2WwqMLkO/B5Ou7ytzbG8xjqQW8buYbvV4bAGBjCEScQtPA/Oe6e67wYxgx6rGfKgRgXzzX
XiKIIEq7AoAqORGE07YE34Mxxiy5AHH4+d4c1xemRb80j2tnHQckXTxpJ0iP/U60GNjJqITy4yqD
H4SSZ5ObhCeNKYsTHFnpdznmDeMzBJROn+VIjadGgjNyvLwaBoyaT944KoGQzg1vmZcMp0hmEl4u
kxIX4efnmfD07fiSovKdmNw1M+YQuBE2CnwRZ3vcVehs37Lg1BPzDUZ3EnaFs5xqWD7+wOc4ICQq
m4CmoLFNWgxVG6EiWcLsN0d+eDhgG440uEqApgd4/jk36NZQlfry5Hj/jdTeSXu084C4j/BWRy/5
WBgIpNDMqFRCllNmfVTJ/01eYhU5jJXYbYMtLdKGSnoJTe+9JpIq3LAT5RY9ONC++1KmWcusptwR
TQkRESPaqf1Sr8Or1dUd+1qEClRGUhJN4KksgqTB6JWH+q+zhlW1AabR4xjVZTJPMGcWMAPP8UVT
DimvHsy6yzBDP0BIBZ7HYXbsMSgZcKOWEOLdCzMNvEno8ndpfBgKah4FPaP2wFPoXW1aD5E8hIoH
K5OG9x1j/+h3jrwsPAbbPgFk1pCA0NB2spwXzqzLh6FiEMhYIIJXRdvPefqH6AJ3nemetp/zoCun
J6UZxFw3bj3O3DZsRtyyMN9OpZTOaTsnutLbNBw3hkYz96VnWOmbgdelUAgXA3GkCYEYPMHiICMV
qrZcIeN/GHurI9BZXMovBxm+CQ0oJfkcZkn+/vxwSs4zeT3eOCTMVtB+NLSoZ3p36wzGX13hM40h
ODrCK8zvQU0EgxO56QnflQnCAtI5SL8mm+RJf8GjTxjkmUxJX6f8CxAtD5V8E2CiwFXXjejMhhyD
cYTWjw7lwnMvwjpFuKeMVJ9kcNPUslHt7XJmQFmTNQaKjYFQXfUVg08VfXg04Uf5eon8og6N4dRf
CDxsFT8j5SDQR8DrlF5W6g55QYiJgSh6Zpk6wkmaS1yK81Dtmmv7tTgQYa84+hMJ/U957DbypjVr
1uU9jyd8aglt8bNAi3ymrcWCTjY5kZvi8HM3zAHbNqRZiWD43X0V6cXKUBRgQjVd0+H+uQCB1YCn
5jrkPaVOsVj3iu9/6pnuAQX5/G1ZDouydRwCfGZimtiTxYuSTDB3LFbSnbQhqGYti48f5li40eS9
EKHQS4sgz+z0ogL4L00hIHFR05OubxztbRnEko4S6njBv3b5ObYY9Cv5hWPSJFd1Ch8T4qvTla/j
StJEyFHO5ONu3L3Gu1s8wtRoT2Bcr0RDtg9o+NEHv9sdIMR2/QomPj+C4TZSneSuGk1TSjsKQDLE
86r0NO8oCdiyljGIpiDoo4bnLrgp1QxF4JOtwlhlmCv8ICZgCs8rMJWioJgGu71fdj8hUv6RRlLJ
yDzP9sMY9c+hI15/1hrWBxf+5J0PWSnM8rZ0GzWvBOBh7WXc5tfy5u4ynmSflaxns65Q88r3hp3p
qiP0FZdUoE06t26ypEtvyd32ZvQKHHVYZkAEY+HzRoiMIrhjKLO2FJWJmOgtGULS/jhFwTU7wRax
SakXwBmdqprIsiE7x1E03ZOp5QT/V0LKH9d18tTFhs7pObpta4gmv/nmSpv0iU25JlxMAqiXEmxb
5XJesmB/eDmeddEEjAd8A3DyaeFaAqRz8KYF8C7RLxGeDfweyeK9a0gxyk5ryfEYKRYmS/tF3rl6
qVMYROMo6lPnFlabQIQUAZ6UznyYs1iqPV2LxMTL97N1AJhyPtiU5FlCQ2l8Z5e+rYmLa3cAP1Q3
UoPQOn0uf0RVPcRJpaR5FNImZIK2x5GrJLdiaYn7Fe/bBsucLVHsIT7ifXw2HEsxolrVSp52WPPx
H314aGSx4xmLdismhEVTFL0Oj66qVjVUASDf+zHuj4W9sAeUo4+1UGGh2PCZfpPnZY1AVL8nbBO1
7KHhaFAtY1TbWwRhZtzIlDgxJrZjmWW4zSVh42N9Q9Y3CzkUIQMD0BFtkk6PT+pxDxFpbMR//9cY
F4wNhcdQM7/j0uW3guT6zL1VigM6ZW3VYkzfY025m2CB9/MC6dnsymV3qp+Wh/wxUMCeYSCqSyFa
oKuGPxHhzX70/4ICDIv2UFD/cItNGRA6f40XiEWgRR6mYfekPQaVb9Om9yS150YO3yFWQ0qAkx60
xHdhZ9+eXKV4UHFlswkOOkGGvCyf/sF66R4EybFyB0TKPEArn6QSJoCbSGxOtQ6v4uxB65NeBE7F
sdFp9YUd+A2mUFpdwYBfkv5QQV3LTIc1uR6YkJ/Ah2BEUYSVQI6ab9dkIrT5eMELKbZOIxq3E3yv
pXUORmRD+/ObJUXCLC/JboO607u4EBvZuyVZnUlcyj98FXHvvAvYIi8XkPXgrkdD9BXnncit+bpi
qa4Y9u/TPSxx4G/nvh4leNe9furBPE8kyRcXbLTUDDjP0Td4K3tpmQlsEmsX0to2qqJAsKT4qyyK
kowSpHARSFZtz09wJfNQXV63XGQelv2WbhGaftpXUrR5XoTDy9mQlORsnjVTbfa5JPSw0Cb8o4ml
GpG852Sz/WHPqawkdUXs5NBGA7JBF8BESM9G++a2+wE78Q1VO7aO8QWXufIs2J7RgnRKFdJJYiLE
tSJ17o4Nx1WLSTCNCJcj8gzOBx1YIJpJrtt1smURcvyMZrEhpbIx7VZGutUwVl/0sOJTgAqacTpW
2CarQVzfbwl3EG+zhhbO+v9bGWwbngF0U5ec5c22vvdkl/6AQIDlnKRYffbJFSVTA6sWSL1nZoox
ffegPcyG6krcInhRGHHsF//W0QKWj8JD2UYuZVbIK7mECxC7lIYtteyG1VEKZI4s0ALCX+ip53Wg
LKCsZkxkeQdMNROQ0gom/iPiLBFlRHWvbp0H2lCOqfp5Jjq+a8aCpc91KgwwomiWOqfpdG41WH+h
oqxQItUvRXGQW9npHj6m8ZG4BtjIn68RfQn+bytEfWxGeEEh2p82b/J9nVpJqzHsB5RJqJna/ckh
rzl1XdjFdqciloyPiGPKaS7Lvmw0tR/Z3hDpnVw/hhhMFEpWpi+zMlMmO2Xp9lMr5OEbv243vyaR
JkLsWhg3vOTvxakt1Ttsx6qZ9ZvFyXawyu6C0H2HtNZkGsCqOfMAc3vogCfEfKC90GMNMgT8y17Z
6zavrWKbnLXZwWsFtqD7FHpIT40n8dikmr6Y/1kC40SOkgVd79qSvrMHhbWUZqkfQZ1EHwVn6fhv
7KFDVuCvPUmYP4eRMcZ5RCJ6efU9T1SSVRfyVcHZ14z6wIHCO2FbG4BnYSXc+9qP8wZ1VqM7O9N8
8xLlsgwnfOo4gr4BGiu8tjE3IJJoOB3qF0Ub8xOjMw1Nji+m+B8enlKLs8Hc08I2HMMbvNsEV4hp
9JvXdndtPeEGUqFTX62Tan14FCso8olr3uVC0Kst6TxgQx7+fe1665Rs+fvVT1tJ2k1mwZ4EwyDQ
sNxnCTXxVFVBWfs3V+LZdsZmcgWVbm1vZNxSvxVjlEGBLLZe7TvurN0R7k2uxb4kK8SHfw+rOtCK
ZDA+bPdQ9WWmJ+79/LJIO139S77KmWjFK6jt3QNPR8R5/bZGc3Dk79cCgbwQDx9oLpppBmUb/z6I
p6HcEuXnmHKYXr7ngyXcy18WtePUNGQvn/oUH05U4OMOMDL2BQm8HNPQb3rRUtuVpom8XjULnDqv
h/53rr0B/VdePBwS1+jaugAzt5/NRRrKfAaPzT+mf/K6Edg2YJg4LIJwskH6MIxGEwsZQ3eAFyRN
cECpZL7/XJlON6f1+xB6trEUwqSOnYwXnVQ2GGROzQkrpzELNhQiotrLAIrQVULhAtpml7VnzApn
Grd+NqcRDCKWuGdfkVNwZbWw96rLVcHSgzjZJhLnQF+5nRQrVqca2c8p5IXPBXz0/ArsZhxoCO77
G07uTwOY+VtyHrKJLDjx+XiO4Mk8h/SiO98vgDSxjVEtgSJFNxn7bQuGhxUbxH/BhPkEVrChJAp6
y+OTnRP9q3ihnVQtOypaWyKQgOvzTgW+M0cndYgCcJmiRmSTJMoos7uuGL14+OwGrDgWx17ZYAgU
Xi8rOhicIxx3l3RH9AwM5OMMj/zDOpaVVBy3vIxMS46yUoaPH1vkKUiAf1aWLFEW6cvizjy6kLOM
chQhjyQKA3u0kMAE0A7tg2UnChuSa4CLi1aMC9u1RP65K4CcxgvV6FrfIeg4kKqzoXLSV4WJjsy4
z5bJMGNjpCULdJ7B1ICcpvE7QWEGGZPiHoFi7bm1culIaXTX9kVKbT5Bw2+yjS0pa0VCaNsM+b+/
KagJ2RuAuY+0ifmln6h3YxXI0f7dycvY2Acjp4qhOunmIc2idHz/VoQ5rfzZBJnWqzLBOebIFH6S
HiabidwHQZhEnRROJ30Kcn7vs73vGyYF8wInvRetGbZ5Mf+c4LL93WNkYIucDR1zGXKUsRWcpRTS
KF7+CevQ2bv8+flujW+rSwT5oQEYrWUJS6LLQQGXzsCZzTMtcj6S74SGFCA+wLIDmJNQBjEjujNB
g+rffuUM9hpCjh7SWlasTH3NsKJ9BTeD7qReJ0o4wqsZ7EfSIJomteArTIvS7JJ0EbzS7PeOi/tq
LPSQOgu/SYJCA6Hmsl1X5OM8pCHj7+saq88qDyQ0Q/UBOOft+ngSmN8G4K7M0A3OU/Pm2+b3mQTv
0t2jwIRAe8GMvhco3WszLISpTxjAX71DtyQ3y+oR3ROadm+ee+8J+ChdBhSLsPaP5xS9kx0eDu57
e7LkbaM0gJJh2rXbKVi48G8cj6Jb3T4fzE6VlNPTnAx6GTn4L7RPGefJkkelrWARS2AjzfC5Xc7z
MRuBbRKq1d3r3THjChHY/4Yl6dTzZ8OCfwwzAmEf238YtVULvVX/56L9jFOX/pPeHwvojRgTQy/y
Ku+wWxuZCV6vwNLl0KZlI1vDXwQ+MQDhKdFlSiaROFBLxDX39PoPlrvyVCAI9UJ2tUh8nYw1rGQw
pDNEx2Qai4UWHyuqNzrkXDyrKq5OVFPJVTMy7ma+Yu4oUsk+6ap0V5sIZRC01/ivmC7DzqCJPVUQ
/+S+VtHMu4e/q3i22X19x0Y5oxJ03a9y6gpdplM90ZJFMykG9G2yzyvI6jeDfdZvpqy3WlPsIRIb
oIS+oygphcqy9RdvBizDbs3uHD6QOQQtjp1Nim9b2Mn9Wbt2lnNl/NPXs8FqPB5k2fK1wRXJvuQN
iYsLn8cmQtDF2oVMBydImnNQAMiYJzgMkBldA5Y+w3K913NqguZpZ+Y8LAad7DmJL2fiCGlPstHk
TJZuKEFLLfM5+NYws9Gd0985e3rHcjReeG5yTJdwvS1hm1N5tsyxXGv7wh+yN1ZHvukqvmHo8QuL
RlwuRoLocswVtuKxEMJkWX3JvUC8REbGjCaT8mQxpr27A12NQo4lraVZd6h/nJtFE5Xhi6x3QQnK
zJy9EXF2PirDubhRi/lXW7WDCrYA7qYUeyvQqxcXdkA1XsQd0tM3XhHoHFfmaXaHVc1wOIr9FYh+
fFdJ+2Mh65j4GvbcmjNbT4riRWs3XKe0x4NuXyE+pBrNPh3sM8Jj8ezEh25AX8rM9zqhDjST4EwS
CbqBOAMTM3vkx2Qtovtgtvh/BqZ2qkDaKRhjZ9OvOpnUEkyRrxnxFebd7JK+KqMssmtHwmalybQ2
5sLV5zepvY/F/0iIgldnkZpt67QVcvwVPYSQ7a9CIaTZ7WDdJfDjEWjOXcGNIy4GgWE+oz4FaFc7
LbcKxFmsrrlBV3VC6qQWh5BNp3989qwBCvLbK/YKC8pu40XEWdrR4/G33hiUryHoxNX5Nw1Z/7VD
yTbvPAfrJvN0Y/jg09ZYMo9wgOYxHzWIeFTQCvg/p2SeLx1AuYOn+V6WRdyU4c2QC/Z7zSDZbGY9
MW8VpPZzImGEtknHe3OLyo5VkR3agO0HfL56OKg3jadBy8xj2fTQBYQ7S1VKimZQbkxTLj1yPrgL
cAGoW8C4dlBjPVOUCYeRJTJlH0yekkPq1nhYddMyNalCWUT7CqYjzRAQGfssU7D1aiDIIXeI2Egd
2mq41rw5IXXYmjLJoaHhRTG4hQzRLRJjIq02bF4yRLFhFGW5V38mWQKPpE2DnJRADvClI88Drl3d
G1SVVDXZs4qeaZkjG2gNx9eN3ynOAOln+qJYflfUZQXAUhqlsiL0G2PcqIO/YJhSdm5nAPyvHHvh
g3txCsCdrJTUiU9aOnQtTfjPr+ne9a8qif5E30aMXFNhnjAt2Df2txgiqRlUEzwakK7J7hryks2i
htQKlff/zUt8/XzFHToIaVCJM8j7iKssGMMQUd3D0f9YgcKkElirJokc473qtGntqbSP4pG7SlV8
8elnOfiW7qYaygh8VuzZbwtv7vkEP7GsMCLZdVq4T9sR6046m/n02HIv6Cc7QRb2UV77w7+zlI4G
3MiCFAuc435HQSViHUOUh7RndIwOEEfniAngE89Jxml1d8A+pxZQlVEAjmX8Ol0RZlWI/CdBcXsR
/A4rYnSdWRS9r4I7Jld1zkjX1I1U+3f5NvuWrweh7kFwZMryKY7R2cxFpkIgYVN9jFZqheZKJ2Ce
DsKdspf3YHswuo10qJVBJnpm3g3IjsDXtWO4dHyBaFHFcfrNKsoBCOYP1UOV9nLgG/LVPhBHoEoW
4jqUIWjpNQmNzG2iM8m4PVlotcX7K+TRPZHkV8XkeRIp6lIC5OTgwsWvLqVDlqqnsLMstQ4pzy3L
3UelX97zAjxW9Ovkjz1NU52dnQ6OrpKhF0VsoXpYEElS3jJafVtAPWhI3qyl7jlPTrMVwda6KWxj
nQ19XL8I5jAjGqA46raUi494pET12xRugmuzeRjjS9twzLNqIPlPmLXAyL86vy3tgUfJqSOEMkCj
HNf0ym4C9JshNqh4EGcWDUHm4Ccs/GucW0inQ5TRLvyX6n2qd5l99so9Iwe5XkJEWu/GwXvSi2lk
JqNNe8pLt7ueHKCK9i2gyY1xDh5kNjH6VF/g7TyKsKVIlVy/tcIUhMrmdvYGDGpDtf14DHey4J5g
i0bRvQBIaSpdDCVGtQFQ9H5f4bPoOuXuoEXGeUq3gz4hWi29PeKeO7Mz1uCkT/LI4ZN50jMQvVRN
Vn1cGNbJ7rr/dWwg2RyG5gttO8cuousmzzhbEZ2of+GShL6ZaN5qRVRO0i2AZ6i/Ku82TqZoo5MK
f44+DvI7wyTQR+f7ER6Y/pu3lT51lLlxoHLwd8igKmsgN3HaMEqJqGK5cTqxklZ1celOwBvBAml6
AacWvuCgiOHDFkxUAVyLFILnYFBy5aL3Ald8UhVGd0K6+5kNI1LcuovpJqMpuhOXRbzqtDja3gbG
//udDvDZraTWlDa0dhpVHdDsZICGPWlQEQDkYj4JBMFomRKQXkRv6jBTF4Hd6xALPadn2w0RnhAR
cfV9iUxP/X1vybz/YgughtEvwOjYAhrvGTEuyLrxXwfX4KsyOQtp4VUAAZSBkyyx4b0752gZ1yjP
ms6e8E4ndTPCB1dnAOI5mNimhrWex4rXKfG/4ncAFEc6gIZ1Bz6w8dvQyiho0fnlvRkz4g/fnm9F
hsLn4lUCpTMoTwEitxdUkpW12iiNxdFfWwVunj4joR47aq2pyvwI8GukcMtlCG3YqR/1Sfaoe+tY
bChhffi3wFEmo04EZwxk6iboKZeUYJ74ZCZMQsRpQnORtnF1w8R4FonvdBCk9zROOZumuUBm0T3R
Z+rL68mlJu9s3NW31jvG5ek4kCc6gvTGOmo4bhnCB7m4/VH5nFpa551WdVFhrSPsrz5/MDEEw7q2
Fg/td9Zo43L8oL+FRnVK1WKcr8igYy8Qi5h7QX9NS4MRCXw5KZA3DXjsyU26cV1f61qO8RvvjY4+
6zNRFYuWfXHME0e+seEU49KhTPPj95756KwnLPnPtPWOUK/eg/v16xBbfaErY8LYpVCCP/vw9Tmn
V4+PIoNxhICOdmKgAJK/Ks3mKY4WfwXklz2T4EZgQVzEio8WwmVFrmQ5bfPYQUx3Isxqq3BlEAsM
NzJp19mWAEhb5Apr5v0DTiLLmeqGxC5GqE/TwZReAgorbzWEmvPDJ7/HHws3KTFiZstaM/r4nwap
xdfP7qYrY9vE2oGPe8m2+5a2/p1ZnFNLExbbE805NekI/2yHwcq7c/YavCt2zBWcDXmv3VsSZa+G
1+04T6jkzDhnNcSXYGEPj3Xz5c/Hcww30kYp8XctptSdDbrqzAO/zn9SvJawcecncYIx+JjXQG4Q
9NB3gJI6v2Rz1BpHB126vv6A4fHkGTkFL8RaX7+ISkuu0Q9IrpwGN4ekq1NHEh60JVCqjOAmWq4r
6uGimU+pORgGobYubDuJikivauGaZZAlxPzWs/HXXO48mtpqJTtPyjidF4UZmgN+CKcK3V123pi5
zKcLN/mO8q1aylT1Td9yD3GUVqRxcXGQPf0Acia71aBA+xROh49FB9lm+pkZiVMgo54BdZWXldb0
iJb5dre6/LGXuEEhmFjMAj3OnZXqWmrKXKHBQLXsPG8ybLZWfCVpcbPCjO+UpqhuGzJfSZaidelM
Myykdc5GKdoVxL02BfXjO5TYwdHqOc4UfLjxlM0FXR5NJm5JZtGg5NZDmEFOpyUAMyFDPzZD6R4+
XqK41x8hxtx6i0k5SJFGrVD52LeZtn17Nec9iOYaT6F8ojruSqjHkqOFkyY0MkkJZ5Bvq0stXlPs
SWVLFyl9eWTMu+DKMh/t4+GwVQgQWuzWepTMycDwqi9vrapM3rhK2s63SUcWPV5UCzBlXZ4F+pSw
g6BewwhPyB65z3Fsc7MXaZj050PuEElyO2wU3F/uik3yNh6S5WcJxdwjdWxLvMyVykx6Z2WnGtsw
+G9l/oZOZRnWviSIHQJBsQruE4+topAwVyOfzVMrg6qs3upgCoxihpAO7BsihCStzPdWdiO6/slI
A8pwLfW46FPNgD4FBNguiPcTH/bM+Vhrl64RyyX06KiUQpautrT8GtB3SbllHtJT2cCxNMkTWyaQ
ugL19DtJ2DR65O3fDI3eyvVGqqjLpDaeAzycPK06U4R8jrWOrB+hTSLQ0UYO5td3TYa6Y7zjBM7B
ogDH1W/2Pg5hWMlxCdIbpIGGgdLyXYYH9yKlR73MX9j4Hpk67BFNkSccQu+1NAMt10I3igwbO4r9
PQ30Lt20P9HMmehB9L+mvSy3hccmCm1+cXHMe4BIenI7R8qBAC3ek/FAehjxXRZLVBylY/iwcQ01
9Fwe2MyufCok1+5qQRdykXyMeYtRA6hYNs9j7MjjWIK9WBEjBxUN6Wxm3fMzOJGJYYuMwkDurjwB
vaXXL+2npWZiOahn/BMNS6D7bgoKJqaRlfpG2HjPkQsfXwwGABou0/wSfLEW4rPkI4YVcy2bQFNW
CHvan7IiuqS9x9OdFAZL5vR+YSUybADQFRNvXyaDpt4g6s/OIHMy7KlF7vGd3wYH3CeZBM0eFAx/
jN5vd37/+5uF27p9CRBJKkkwcQLv/8gJ0Gl5yKYEJ/kgFFe+AEUBH6ql6eOb8hMDLEpylIKnC17Q
Ey56OHSdVGT7iQD5EVzp7V3oNejT0ro3hz/8rvbpy6VHAnmcSihdtF20D2378vsIw72zkhj5quxQ
ciW8FO93IaDkjBDNd10rZm7Af50FNb+rf6p6W6vJElAaDJjIfrraE//FB+mPhxq8w6UYoMttEyHB
NCnxEBLgd72qCrPWyG9Up758pq87+fuCfrkSGNdBfUNip5Zhhv4FIlWwop6Tu+WOhB1ca0KC8Nhn
PBP2NgKKTb+MO//lu0o7PGeGk8AdKfsFMFn6EYc8yTxxdr34zciF71tX7ynl1Y5GOoFdL8PQN40s
qI90hTLHjRb+a8JsC5b8hGpERldwot53rRXVMSaBIs3WEaqs5R6IWr/o0frPm1VeCyKtFePhNxRm
TUDQvbPdS9KFYrdu3Uaa05ooYf+sfUxBHtKIBDwcBI2Ig+BG/U/wSYS54LYtjPJu50GkfBbv4VL/
OD++zjvqyLxB2NTjt0CjDi5nisfXyO1BPz+W3iR0ydsknPhw5SSGGEpJpWq4YRTAJ4FDuEy/q+Xc
1dw6/0e3py/Bpo+6D+0L85GKLVckCHNN5vVURHX8oyhmK95uW2uh2f0BK6Bkhh8GF4jUtxz3K5mq
1idGusjcGiNK5CzwYgbvwdtdYAYbSc4FvzB/XTDn367N2w7ftefitPawbgR49TQu5Uj05pYowqGl
QSlqywLrqEHUSDGx4BvYfFybXodfSlxJhGc95AOOSI+SyO1RrcKz/GFsgn/IIcbeqrO6wRucI0uk
RJyrlI3IGeCf6P83jrG/NwNcYJrJesr3EWucCNIZdHvrwb02A5r+oNndrjj5oAkXTrrI0CtO9eyu
/RFCEmaVsd4+1KpjhTMK/TsBkuq+a7Q2hM0yfzPk/nduafIeTJT652wZtALZ25sBATir+YzatQw8
iwMsxYXB4h2pDzqVbgeZhzqBsKWgWsbr0diOIpnE2nkSOOdhSVg+ja4B1w+D1PmN/yqj0p/FuN5a
CQ5AiT2etOrnep3bvZ7viHmb4k0JOyZk5Scj3BO9DXhK13mJxHXW/2IyAuIsEmKfN9KzuarOl/W3
KrZySsBJHbG0tH/8XbSqTY6BJhM3WugiSFOYPRjT0zCIr8Es07cKXzBn4bgquYbEzBp1T/9reWlW
38SMxhJXBJU3loO0BsvDlXTrl1jqgsl7S/fO6CjS3XllIHd7ErpGbDlRbNeSfh/Vw6L2PGuuwetg
Ee/UZB2tEkCxXTF3JJ8YsRjUjguzgiHdwwWdJt20UB8hophFTDYtxvdO+YpfvrLR0e230ZdbYHw1
ndnb0oiGRJdVlagiasrUpAu36Uya0HgbQvV+Gpi6nmrv2oVJVIcVkPLWMCbnYIP9PT4pd4sRTU2u
NMtx2SyLKruLp0vbGiRBrNhwT/RcwASHbVjt1MDIlFe0CZIoHufHEePC4+a6VzzsXIuOg9xtlCP4
8bo4yVy8R5GwxtLgS+tKt7lvi/Q5yRU8+EB8wmJb4E3igLh6qONdGPj1sfJijDdeJTtJ0Cim91yb
Lwa48d/EsoIExw+UefMBAPT45bL0Em6Esnm9UZBnkBmXFkYDu9nekkJM2hFxbFRhLsH8piCzZpgy
be0pM+ozMdMi+Cz/28ZJ87YSYWydGHTJmXe+WV8hRWGWREyhigxK1uhlMnGIoODVGL/0LqgkF7WP
7+Q5vS+vhFOj48jgobWOS8d1mhF9P5uJ5LRXprCglBBDyM3NTEoIbJnU68N5PhowKWCfcNgu01zw
uJ5RkzevMRECzdijlW/VZBJE5XXb6L1He2MGrE/dwNowJWlv4SA9LqlBg1A2IvZx5UTLpPmJ6Bm+
CduYAqSZAf46EbFDXKXpWcQjaAYfcQLyHCj5WT0RIKpmdmGUHixCNq0PQf4Jih+q0VQoxAn7xYxu
8vhgRKPfcF06ZJmeKomdBgVBj/IMZ1yutW2vO6LFOnm1HCcwXynCC0zyvcUfZGqKcrtomPO5hw5N
Sp/a8wwCetUIGyq+4J1eGIgIeTTkwbqDrRQosRetoMkZUv4yob7Glznrnp0wayzACITRTjYypwan
FZxbCGyTNExh72p62v4ie8AaMa2IeF7gHPrsULGvdD3aYe8cuQ3dbVW2uzkKdusgI4rxe9GHPAqM
ptPa3l+7rljWYtjQNPP8sWCeGacae0aRwzGF0d1hLgIW5zm2LO9hWkrvoE64iPsBs6En+zFPKr6Q
KMn6rRoAzhCP4E8DXeQKset65DA7iU3TtF1Hwon6h0Cjxj77lHwUOWe/9C5HdjtNi9CwJ6Jviozf
ls3ybqxsRDoMSObhhwDIx+DINFBIFBTJWaMTEkrCxB1VNTxdk4ctZK7zFydPNFytqrlqnH1srgNG
U0QDfqJ3sTtO2Bli3sMX/bg5mSMPfH+RkcGOOBf2JBk7y99hLBJhtlG53vRexoElp3Mp9Lp+gMC/
vAViqHZbT9MeRHGe2iWmxqpgqZ7rAnT4vAEvkNXpNKyDbFcvXb3loJqrLPSwjZoY1CX4Xv+kmTHj
sXAuVwlVVhkM+4fzV8tA3nA+2G298XDtu0NssHm0n6gKl70tUbupwJCrSMUdmtxEdSd2lXJ5KyJM
JxwOB2O7wHGFrr+z5OgMt5CspObiVdhik+/aT6jSu+QUxrupdxxu8p0IhaQ2xvAJ58GQFr7FeD+i
w3hzBPw6Jh075PiD8TjcenNJsQwQgaIszPlc07BwoNGElHgQ8J/M77QaXEc8cjWp+KsINKAjzaEC
bQVxBHNNQBKmFeTOZjZjTh+b3jK4Q0mdKAtMOwhCBrbew5FxyYtb8ppaNsdK3UI3zbax0mg1POng
btVRVBq5J7zTisLcxdG9WmR/PPDetjzvRoWMkRweL19JF6V/bwjaIpdVevn0Mhukwcx5V5uXAemh
E1AplksYbyva9BHKykr0vi0tppqfI1P6Tm1MylrMuX+tfkGsuiJa2H3sG52LSxbboazQTp7c71yg
j3nzorFVeF2tNKhMj7F8T5sNd3ZEIZvZclwqaLi/2hf8w0SbZYwWorYiDmrps3jGvjOOqetrIQEd
Rw64ZBgL5prkgS46aRpkHTEPNhQThAYqsE0DXsOZHxsiXOlodegtiE4Kc77/0uhGicdPTHCyURYj
oW8zmflSzujxPGIgBEhMN/dygOfVCPzT+pIfbqXHI2qpR+/QmjeFCwV+2t8rcEzkmFUEl0qPuJU0
oEpo185oEKrzyAhTTSoeLto+AT4w5lnl/n/+WGe0nuen4weaamgXBl13jxjLWL57KhA8oNo8dkPi
BiBkKCTFkjrl+uysNUWLBU2AZRCilYGHXvRh33Z2JZgBdK4AboGohffwtxzU2ZiwdYW+JOGUKDRo
JCG2M2Dtft8SywObPC7VGdjZGlQ9az502okwgky9bj2e8WhVmDhdHMYe6KnjzAB5flCpx+sHpWQE
mjHUSzOgCgQJdfHEKStAC0GWoPtZUDSjbCFJRJIMwE6SewnzBqHw/GMDYDMuwMT9HM79yXuzAxz2
NZME0wHY9XfR1bOSoK6A1dOUsfUGq4uzT2ZK36yXAS2gRnNSXUW3Jg90DmMK0mmKibvYnge5CRia
wqilQCUuxnPRaozKpXaBiqdkCgcj0Zhfimxk4mfVLrMCkxgk4xAqAIMmoW7K4e2GDZKfKzSOqoFy
VOZKOvW0yWbzFYNzvpOmQjmI/+yr9uHKd4ZNpWSj1SoL/7hbmZFZHTmlWUzxbh884Y6bBMZCk52O
kkNGJV4ZS+AYTcvDu+nks8gTfQEGOEVVaefcJWN+zNxXuuqAbtwBjFhN98zNZPRefU4dxB0iwx2f
qhdnhi6I+q8guCSxe+ExSe6QbDwfSP1InMdO7YQ7FU1cK/3ZekVi/bwFt05mcag9wtSTnZfnpUGQ
4VJbZrh9y42bO+4OR6k8EYKdR9ebKIa9vsqJxPRoHaTOEHc5Qas6UuRB6x/u4uVLjS56coD3sCF7
49elQgoQ+calS8SWOrxdEYwGJ/6nts3aOKDIUXR1H9qp1KENM1e00tqhBFky/tLIZAHhptyTlg0p
oR8fXZbWOjnQ43/jTvpipimxg8Q1fHBn0f0YCc1exlkZ5YCwxgW9F2WTbQgWhJHhuYzkGwQrNjsv
nIff0W4q/0BSqi/0VRQ9yA17Pm2VeiU5woTKuOyCPJfjfbVFPEfSkmSXgOB7ft1y5I6YVLvJJ6BM
A8JCTJw5g5dO0yRLaPBtDbg67yu/X/iMhjGAv55L8NUuYJLqLmaGuNj9K4pvMZ6+dYmFfKGL9I5J
RHbOpfxGGScyU7gat4gGAYdvOsIuYLL8Z5loZcSe5PI/b7XBFLQzLkC10tDcVh1lqY/YIizW30sN
2rzpJ2QZl1p4B21Wf61lrTZ6HuCkHRhIWCs5dt2NYOt2b3elqlgdUqJVMhOzRgq4uoEcax5ZNyst
VEsgz1T8nADgV1TI5WnGXTD45V26jJSXCXuFg2rYg5Ui/sWzO8zlvy7W90fb35tGI4+xZVUIPkHF
LPlmfl+kJBYTBr2duNzTV+n4CyRFUXSGdGnTZtrTQXDxZRdtTzZN7D/AN+O282lO1z+TKJK+3e+j
UeDp4X4WivLTIFcZliGbjhAJRcVggrkuBwy960ZOjFok8wSSHfNKEYS9UopXWcl2RhRJ8b8rcllE
mbf5WeoSaJS1FFHoA73rtSAxToaJ7xSoTG+80DazQd3f/zotChzULMqnra6xFYwPBzfGI6gBj3h9
MB/aBZkvUiYihP0NWIf/AStmpSz7jVkJylKe0f+TBPVEa0/6n0lwaHpvttuQxSgzrRzRI/nejmdh
aNarJt3yptvXoJO6e1lPgdf8EUnU5wRJW925MFasHA+ghaCQjGqvFAEPznHJMLDgjJsq4UpufBuO
QL56KIVRf9xVDnS9NXBqPuTEvhEfnh3oN9+7jN9uSU9g7hpUm6CIu8lXoj/NAerPW9L1idj9GE6z
oqtzUkfEcY7XQKkh0xtjYeymQ5lCxvv50Y4l2elY/Ib8YjZivOVTGhA51GtDsghE1fCHqHRNVfjB
POOFCgFnZPddNLc3xhHll4Sy01DnD/cT+jP6p9edygdW/A16lba3md56XFGBPNZ+t3bhvwZmEctJ
qFvJLFZAlGUOKIoVDO9c3o6MMzZH4njzLKvqwkSBKaU+Xe/gEE8W7QESVHtCMNZx04deZYdzZ+vy
+3syp6dQCOkzBDK/zrG30W0e+wgR245yKMspTUWjjCtL0P2qFZgZewttD+Ro3oP1OY0yx/l4UHB9
oniIwCv3gmt31ix6LvtC1RUAYzWYEWwiOM9Io+8TjXbiVXYCvGpnNTmuletM29SJicQ6w7tMt4TK
g76IrqEzKNDGYYPzKBj/80OuqZ6rf67COOtaZKRFyMWDc7tuAW3gZbsY3Zg6hmYw/cspA57RdAvZ
mT5Rw5l1qtlx3CHkL+L8/U0vWu7NmbzDeSKBRAYtYmhF4PqzzrW1eRjIxehIU3dyQj/RrXI5P96A
WfpdHC+vJhfYfI+jQQw2y9FQyP2VwNJ5rurYdun0Z96nqwpfqjW3Ch3zmCSyl3eZ2fzVLGZJbZHu
92v5YuFj6012h5SUO3BrVCrFix0ATB2ZsoZHAMsUnRoqs27vEUzzus5e5/M/3nuzEHLBEvWcIAHr
jvfGfpgmPVl1PpVZ8BgIaMSx1HI8fIf46OoPmhHeqMngreYdTRagomLxrbwg/irc0Sh+T9FQ3mCS
2bFL85oVgCBQEGdmnZRg2Xu/5DVSzZzFnhJrf346njfewIbd1tZdzR9bHD7DhZEWPP0nERMPS46u
+s28wpibaAtK2q3CB+mAzOBBxamNY+Xl5ms8fBpNBSCa2LcngqIgmatPqxoWB8+1XwfYzVi2Vpa9
yGFm9gtDwUh8uWsjaXDX0L+HfY3WAwGEraMjdOTqgDV6/vpKbq4TYhifAOkWqnXZwli0rmfP7UAj
b6R6BXBl/5casptj/xer8Wo9doUjyOPGiF5bJ/AaSDDk1yd66xyU3Vi1qQtRGUb0qZ0a0g0Fi4uF
9tgx2xFTi+Aj6npmm6cGXS3jMWf5SuagNjHMWN/tZamQZG+dQ2l5htakCZrBhgCMnUFGKOdjdnxf
DXo4x+0GLhq4xNpGazTHWvY1p6Ews2eKW3SwwuknFnZeRwa/V13F4jNHYh3qLSU9eKwnVta3XDXy
6LunxXcTlKxVv9ouB8jAr6Krot1kSkbkir4xf9fPSOE6fu8a7nGHYQI6gNP4CsvApVqMHgES+Fv+
6qPza5o4bZsP9zm5oZCAagEztqXV54CuA/XEZdUhFP6LDgdnyvAceR00HIymOO2LMqlv+70jNH5k
3D5oMfIZvHNL1zaM6qIGiJJR1UV6fT5OpTEpuPSOGlHgOFUucde5IkP0bNacAR5mBiVIiOcvaUX8
wjVjX+ZpitHB1V4LQf5mKXW8THLxDDJ2T9ct7OGOvMN+6/hXwya0op128SIjRk5VXPuwMrW1j4Mk
I5i3mPUwj7jxrMgjpTomm+auECfX3b1kp8ui4sQ9oKvS729BfnKtx7pWvnNYZDyk+ZPGbMhc3C0U
pCeGM97ZvvweLWJ5gdtOnlo3LiGcMPopAXC67mC9TIOEXM0c94lXzQO5P4nNafJ7b6Yxkqv8YaK9
APBr8aGnKSlwm0ptP7D9KgUl9jxCufRN0i2K8UT0G+mq8Od4FlBD3ZzReG+CCjRrVQcOFo9Z17+Y
cX/y1GCsLslGDK7SA9awsPlc1OI2xJmXofBErsKvpD4vpO/YKPQuSlf23CH1dhkJsRZdAgqf6Hh1
CT+gAEWrwIF+/nvG/bYAdNhoTiQxa4NN0/JIQaV5CTdiR7HgHnSrRW0zcNJgmPkit8TU6A1y9I4D
Vlq9OM0HNjKBfWVizQtWrO5UImi4rYkADCAPY53MeEMYU3nP36nUtuxVH8ktRO/SKOkFOjIhff7H
N+NesTNUoi2SwEcz3ha7HTL+y8Xw3kHxVPXxdeuWnBlc/VlTQkmq9/OFhIMYC3xQZFreiWj+JTYT
I8fR66S/JJmCTlxayoaN6gClYdXqCB5KIAZmg0sQlnQjtZYjObuQW6iVcHgOqmGOaQHHR+DnDEGI
qy++EQ3XuiHlOKT4iShRhbpmwQr/p4Wkxf4Ra4aSZpcDA5QKE37hAl0QB9lWrAC/bff3jdsbGgUl
G0KW6r8Yfhctz2niheJRGqFtPAJ/ZY4fkhQLrm36CM0s+0OeAzdqYm/ZyDOXehyuyJ9xCeP7fb/6
n64CWZNAaqPCwXPqDIMHSI9qwq60+zXFvlPLMQCDX9lVqplvD7jAwxD9Hsp+a1pi8KdraKAxoss9
dPlx7ppkXsi1qEd5oTOHLrBjkBOlUQfcK06kMRHQOh4f02/eBWFFO5x2iLDLUpGN1TvY2L1jArfx
3uylhVufGZ1d69/fDwFGCBKtdgeXVblQLU/5wqsGWD4NKuUIDRnOFPMK9C/+DtG9e+9cA+A0WBAc
YlQrF94Wl44nGSn4JIppSAyAd/Mu5n7w+Zkso8dihNjPLeUJ90kzHBBsnfsUoiZJv8ZrDITjfidA
PCutNnlFJlDb/iOvwQ4dnEOCIgSWqU48Dn8GR01ukbc+q8KaKrOisExKyDfj8n52YUxH+wYdd17d
I1EgKoZ+NCaH4MaKKd613w4skm5Cp44J4Tpul15pW6p9rU1GwAoQLe4ni2hFZLFXCGPxjZNrYq+S
0/K2+4uQvOc9tUKR+yGDq3vFQQdDcV4sD0o73bAQIWdaDvZBnNMXOBWPnGKM6TLMLHdEI1KkB/jh
6Z34gBcsXz4+IAWfxEqYdG39YnENAAXqpjZUCBZTOSvURZRryEjBv2NQBrdETv1i7T3iKZByaR3k
BEtwQFh25SOpG1pYcHJx+s+23QUG73hVtJmZ8F/fZ+i3l1tmpKtLrYc/SNrKgqwh+BzDZ7ZXGjcQ
63dalWjhcOOv/woAAbEefShe6TuovYBEm9yzitDs6u547UIPOpXFQpiymsH1r1IMHtIovG3u0m9o
G4jFokNtvu4jD67gRGyZMUIxeweoe4m2HTrdyMCLrifmejRoGTjAyxZZ1GXF7YY9Z7Ub3waWLG+J
WZ4Q2inPO7lEJAo70sDAq0ngmZ6Ffeo7UBgxJIOkJ8H3Vt56+oxOsH3OhJfcLy9+yqJyyjwNUAdf
G5KW+IhLgznmN+cSXAaTN8se1LvxAnht7mvBidpk4CS4gX+CTopN+7DSicQeorQ4y5Fkx0WHni2E
SuTowDIo0hI9p7cGLxKhrFTcyzqwsHwgmSXNoD3d4sugVVyPZ4b5CyitpgcUcx+cMSY9gaFcGzfL
JP4UarD9qZX0CdFyyxL9q/nN64blcalrdIPugJDrtm3Mxb0fh08bmOiKi4k5IY4TtCv4Sa/smNB4
Oh+PjwFjkz1zaRepv4vE6t93xhwj4jA/LSM9P4vcQJL8Ewbrt9fZWUKG2pgX2cd0opkqmbyqJ6lA
CckpCbKsZjab5YGWFMpmMaGRRZs/bDbBoivTuj1swIodWS5xNT/SyVVvIpefhkliGQQPoD+SUZNz
rLYR1qS7hNsfLu8u8cjnsSHHjjlVUt5sMTrzBSH1RitDDfxykiZ1j/ugrYi6j425ejpurKLzSFvx
QimJnFWP+UgoTJxqQsbcv/7lYz4OX4jJfHccSzSsh9YOrbYS1Jw7vAV0vVFYfZDrtcTg9xi1KUfZ
oxiZ5BkxQ//DmyB4QbIROHy72DErh/LWwyeOMlZIlHZbam9fli3wR3mEDSaXAYuKNdAIVV/HM83T
2MxSM8V2dx9HNYIN16Sk4kwWS29EHiBW8bqax0oaJs/IXXdXss9FEiyht08tYOgPLmDVmI01JFb1
wrmIy8nzcBxLHWtyx/C7O8/bezmYjzNpF5Mr2Hk7dLDs6ojZ6I/VClLlZmr3Gk+C2b/gUv2dTahI
lGhPXGoBNpD3YiBoZPOtnJGTtQrteDtlXkHSD0WmnuYIS3spaq2b6ki2Yt2ZmCDDFNc8Vqm8N8xq
quVKTwXITrJfEp66Ko4QTDC/EOA4xBFQ71MsvQFwKSh5HVeOaV+ReaZQWZHn+8r5+AtjmcFwHZRY
u0+fZShB61nJTr2lOkODPM7NhEcbpPC1b/31KMBf2jDQOUXCBi6z9D5Cof3yVnmGHc64aNY2THnp
ECbZ8rECbn8GU+a+dSElmMHy6V0/UzXVUF/CK0mFhuPlIV5MR99lB9CfWLP8HO7sunvlMb5xuCgj
usncn/USkuK1R0rHwoJD9nKmy8RZK2lJ6C2F2kH/cZsJVefv1TnGyTCPgqUizdEWtxte8AevBWXl
FyDRyveDaS88pITQFSKB7CcfDlvNOxkWlsOQJRBtrfMceBgpMTpnvtRAvce5cY/hj6SimtrC8GcT
lB5QYtOjdwCJ4+VEhn8cawo3IItIIpZTIwZSbMsZQN+2O/6mjkbanns5B/TGDbAM1rGxJJiAI6mo
X02oqf/tZJgyob4hloGcJ9vAJ93okdjF4lRFfQAihI3AaA2L0GjnlBTgIabv+RWfDsQD71n0xQP4
juZwzQRzdZ4vTBhKEP+mJH88s9PvG5XRki1ry313rZz3qNwaugFrc+99JrXSmxK47+jtkPRRdpoh
jHB9asstTXxE5ZTr+4chejZJP2ukYi/YR5OWc4D2ifodXKmPy2m8O2Zf+/dfNK6rM+G4AzTuA2dC
x1THLLjY3howdB91CHxF7PpRsPNKLm5H50hTvIxryOKAOihNLh+dy0OuZbtQ91IRXEo137LDoRJx
vulDfp/bgFwDfR8xS/Wv5Zd9w43/nguewchE8glg0AVLYDa8C0ZPIBPxNVh92gmuKJSRBaaE0wYI
MQ0Gwvp83PDiLZ+zGSj4J46J0+/AmD/VgnUB5KUxhkVT9y8ZGk7479ZDJPVffCeVg20Ypr9bhV1W
Ap97IC4ZS3J+jPzsd+QaMU791i/B6I8IeYoFdTL/cVUnyHPctDlpDbP/J80MulokuZQYIHsu8C3x
gw8Wyq2Gpo1+jFjlCvQ8BErDqFP5XqO3fiO3qUXvU+5yAgnTczKyGktN0+Wnh6QfU3RJnxs/4sbi
YZsLub2WsmaAalT824u0Eg+oABdkFzzphilhaWw90WR8fY0YaYJnubSImy9CAMOANPFpgUwdwShY
OGRou7tT+vBlI5Jz5HhvKN6XyMA8NNo2fmf5rRVm/dZIhYo25ggpOLXps/mKwxLQiC5sDIpBJ4Jl
d2ckcFtQtd1aGtyR68sylmj0zEQ4NkF3q8PLZNaK8tGMLqZQt2qdscd61kPzzE1QSE3rCvqAno50
uLngl/y2aEQ0SdAoIdWcXfYqDYRF8oyxXcX05ndXcaLwTRjEODG1zyxJA8nWHqZwSAn6Tbp5aTfH
1wIgw4c5drXb98JYxS1myDoqu20nWH4RMx9WJFpHRjdww9lbeP2+9Xh0hZM9riqVowpA1uCwRaud
E6M3F4hQ3BvY5fCx9GF5AU5oCCkaCdxuN9IQglNqHCyY+cnsAMYCDE/A6N3UGy/C3OSMo9GVYvy8
whcqs/7OujMyB6uP5IT+8DdO9OTZvw/bOlfj3CMFUHPnyKfNMTzb2S/SMdaTxOWu8bOKcmKWnL8k
uARHR7vh6yBMloHnseO2igkt9vhk0nNjEXR3bGy7mUIIOZoHMzc0pR4s8pMp4JV+sH9s/BDlqDt+
z+p+xiDNDRLIc39bVA6KPQKR8F3jfNTwthLAbrobh4mxKTC+JqwbIZEerlrToCU2tNrCu5e21iGG
5nwQVKZHg5WdDYIZXCIrFR2aHro4RPQEh4EczvQLmXuLDTZFoV4UyfkWNJObEVjEZ6ReFmh2k/WN
ijPIwcX/xQD3ZZpDyW4Rhur65YFSgkEc1nmLCbeBDo8XeQvBj8sk2/rb6as7yoJHU26bhUL5Uqej
j82yw54U50xrw8ohzSVq4uWgFYngBGCsvyOIwToWhFPoaHPy8ssCZEulV4qsi39Hbk/v9h7hnWG6
y4uMZDq0I4bzKT+JutdluzxzL+aGDUwDsDUX09gMZlqvFmpdkbZ0tcr2VKcwXUkKSR7eZ4MwHuGV
BaDoJ7UqZNwZg8Ds6wDSitwt4zte4Ch/IEX4C6TQ+X0esfM8cUW4UUZEqLx5mfwKhaqHTz0ZoNDG
jBw2rW7l7srSSGo0P3b+XPSaqQzh2eYIuudqDF60XNperNj0ZLf4vsHOmyt9wlxmTysT0eAGvl4p
fBWX4i8TvbzSYi0B0znSXx4k7Mp3XgY06s6Sa47twpm9B/UVMqjvjwnIasB2Um3MxL35b4Ojkdaw
Yq1pSAwEcNeOxw+SS0Q8ommHeXbPlp5jYzuMYo5FNGvxgi9ok8oj/o9EHzkV37NRu9CBKDXy2XP5
bfOlXzUBUdP5uiuan4zY2AehjdDlrmgizDxiIT5+/WcL5dFhbXgHKe0cL0kKVDaEqFmdzW/8mdNI
6IUXQ56MYLPeNlQJrFPBb1k7HSZaAIqoZqfXsa5vIYCI1I0WITjvDPX0oH4VFXBEyoLg7dWodR0f
/gz/W5YjDLuZKO7kEkbM8ve6olfDpaon278YuQu60Kt+maRrYpCnp4NrlREzFWZ9jM2umYkG6DES
Y4aBbUxjYSxeOg2DQ861X84VWiuq6Jx9r7th0agoMWFKy6abZbUZVYESJvb7wHM2Pq9qVZ8JA3yJ
sUMbHpDnjfo+A5kiwUbIBXxzEqnkDrkIk58elX654pnI7/dZ63paMnK5ydcZbsKtsQ24K/91LMoe
ktT40ExyAEyJE6d9o//RqZAoTek6cBzJmc6XLD9/nXvD2nOfi39PlBrPjQn5x1F8z+u1PXrWYyTN
iLqes7cE1+yGx99eJMheVcRyu/Odrltr8TvS89Ara/w0FJhUL6KNNHYDhMX1EDwY9pT+tWnS0z/z
nBnGZHKeOrocTY/eGlYmty2Uzg6O0zmFa64eGPcFJWlDEk3PMyG4Fc14aWJOWRa7h/lOln1ZrtpD
3lVDbS8FPJxkFRtR/L7lSlxKLS97alkP4AeJRr1qRh7VwmMTFIEy5VdYbcpNnY4QPE6kN8ZHkC8X
iq/EAKgF7BBd++ZQj81KNc5PV1ZsYB5ev7L7K1FzmAa//Mo6bZoS44MwlpM6DvHi9JmL2iy7ee2U
hvSRIxogYX4w6BhUChS3nIwXFU8a3K6RmO0oLtjjQYlbApq6TJVZ+GX8cAdSXYA+0fn9ENueNAB8
2NBY1/tnsrDegbeC1REVESLK3Um3JWKjus1/tU2KxCZTlLlLOoUh6i16JSiZ6RZDlEL7w3ZrH5ES
Z7X5LJK8txY8G7MI9RPPAI3oY2n9TOBYeLeHKIK6SKpORrX+pMfmgGofAcfCqXvEO9Tj6B/8gMBH
SdxHfQaSE9dsyib+tyFKKkdrUOU6zteRlwtne/CqUPGqltDVvy4ccuOPdlst5n01IDGKdilPx5zq
D5Or8UHRdGQ6yxEtQLo+/RowCka+wNk3tIKXAr1MJqPZClbubc5BP+ASNUFXUL/t3r741loyoJkr
LLEFZzWATsgdkawPh9kXkTkon8caJrVgMPX+wAyfYCzbYAjZJm3dKIdO8FYetACR4cDnyh5X5U7w
iWWZVSy1/cJ5iP2wsPyq41PSQd6AjYQw9SIoLw9T1dNVBn6cS2gtxMda3tKtMQws6EVtshos1Qgm
4z5ovWlwwWs+Y6F9j/rQDji8Tmq6RXYr8gLAL54PNEtH8K/ecD9ojM7Q6OJD8+hS82D2RcRGZtAF
Lw67SvFaVZZIt2sasm/RBjTq+wt8QBb3ZVZX3UgmsWXzV8jJeftrUO/RMWwg2PLg8tC17gwx5KO2
mQYOuJF5jmSIoquTp09DV9FK6kV67+eY+zONMgsPQ+lg6Gjhy99wRvDEweJc+snAARaOxOdnES7f
1WAyL1SvJnJgcodl3r9Lbf9FvyAokVfqSAUYS5y2yBqJgK6mmwgsI/6bsGYVIKv9puul5VNR9wUI
UOOGjlIt7aXSPkK0jCi9wSGWOSjwpH1rkfvIxSQ4Aqx3HfhKAA2ygla+Nshs6hSlh/GktDWEoDYc
cjHpRZgVGUZnXc1NSTpXxDUU3TsMttJKkNH9QJYzGWxk9mCkworEMnC+3x2qvsuN4zD6LFFftWbm
Ex7UwgoLP2MixgDHM6+7WpRRYu1eF8GKmUX5/aXWbqjD1BQm9DE4JBVfVEmeDpJwl2yJeLUpffWB
sox1cLazDkD2moiHBK5kNjZ8Ng/G4CEVUtT3yPBJD7fa44I/6vd6IUDN/4ACPSkM28+RALKVohv1
//Kthilfs++ouha/EIBTCJAO4P+PXLdk6+i08RqHv8ZlyarSI1Cvh7cR4FdXZcKEBqvBiEpoYM5K
XhF/F0kExajnoh3x6u9RmCCJq1JKY6pkOHVE9zPkJ/g6PC/Tnv/5/ZsTSITp2CL7OLpzMTkZ+PHU
9G+Vs0jRSTtmhrrmEwJm4pa2KtcXP8MCOCV1JD8jH1AN9OJRy3lPM0DEdiWtG1sYesaHf0lHlmJ0
4okqzMZ0j+loFCxKv+tBxwCXVLPcOLSKNR0UeHLWF4FY+I7gxr4ip7WUDiC6gNjYKAGQWiTXHCHf
xfrmaD7TAVS/vkxE4v7k1wzNYJHPAF71gPdjmRAiGOcRpDG5lNJqgSqBlYw0QSj3hbY0+uRFafqZ
FQJfTbhs2mxxYiaSLvrNIC3a3CMsEnchSL5Y1/NuLHPsqZ+hTfBsI/z/BCDJhGDZQBsNDlnjXO3S
7TBK9fR0bPqKEDhHQ0+aZFigu/b/HYdUOv1GxozMcx+KPzbAxcFXhMS/q1BR08Ir5QNUVNZLCibZ
LePDNRkachROWKazjolCQu4gw7wst3hYN5dOz5LsjFYbXCOeHlbCx80y8BSypqMdRvAah1IBw21k
H4/qoxsiwjEwur3zl0XVjDosG/UNfVLagl/0fKOEcgBt8x8XlrmhLlm1v7F1Ps0dxiCLfUZSsar7
+7j+++5l3Dj43Nto5g6ALocM1a53DYuW0UgAXaQQmTvDFjZ3LcGajzHPxtxjVoJjI/9Ndgq8G/RJ
VLT2WMqqzVRIpa2mDD7m/eWvJXxF1E36DuLgCusCJcwDpaI7BLcTaiP8fL0FjJmbSCu9OAKpFG8b
m+nO2HF9n+NPMspZnO+/9Gg2kQfhrGh/1yfsMR8WHrc24s61+FaN+jn9hgfGslu5kxbndyAf2HUS
72Wi+WrhSr6IkaYFectS/c7PvukUJ4dqFmsipXPTccpeuUwhPhiwk39V0bKnqY7PGcpeAK2leOuM
dV0kABnKURUx6Tzbho+DN2pZxNZIaXhAkUT2YGfaEdQJqhurZh5cgm6InLvPhoQg3EjDeut6lYYf
2qcwMKFyPuEiK/Z9RzG6ofrGT8OiglBpQfZ3sNanfjYda7Zcp9JcYA1Z+4VT3e/MNDFAjT+nokZi
YkEysR79Da1bcqgYPL4QvMVlOuWnILYqN2z4o2SUOqzJd++UNeYU50MxZtnq4cUQEp2G8Z6T+bt8
Pt5cjcQ7K1j0AAL+IOwV9nUzoltuTFkV6Dv6+AmSewgMNHqn8xwGHtS/twscPLlPdAbRQCsAC1NK
HwDJ5zJ95PJodTnHBLsKylRVs8OfAJAfolwjSJE33s2sGwgmbGFQAPTC21PeBvZgbQsTd6WlQjBg
gVXzSEZ42AlZlguADsYeib8zBmhm/bv63/n66k8Buz1rOD9wPKkzDl342ia9JZ0+KRcr6SGD9Y10
b445Z9LT/5B/koPQ6Q3CI4MTUdRK0WWAkHG6DSHD/2TjYvDTofoJJq4g/FP3TgdiUgjkapsNG7of
ex4VBUKSAkKmKuGi4QvzF2h3PP6kM/X32fezs/2D6NX7jWsEFAITE60s/G6WI7udlH1AaoDmtVIu
lDFnzHeE/UDye4AIXtIpMeR75REmZ2YrOde0/vLyAd9kWbFMl8O/y0gOo7LmCwjy8aPQUNfE4jpn
EivaRqM1PckW6ZT5XH3yFWW00KT39czuV8gE64YQZcSoyeAyfpWuJisSGgdkXW+v/nh7dhiKIBJ1
RLBUNvBTKtcc97s4KPoP0n0NSoXbn3P7M6Bw+P13VlljvAitZpJ58KKQLMwIlUhcmu+7/wrk+tBl
wJRZtMbo+bnc5DRqO7I3Q8IiGoPm+JW+bSfaNeIk4LB2OPoinoryYNYxhCjLsu2TWBu6l4+Wb0X3
vEG9cJ2nzozG8jE8QHc37KNqsUqzEAISuE0vFcSvjVut2PP3F4vTxEjPdXWVLRGqe+Mx97O/39+k
wyBw8C617/uZdE7g+RdwCmWqUjyy/si8pz0zrun7iBA7YAfau9Gx1R9MtU2Wx9Xi55vUzyCt3HSc
x0mnQ27P9ydUvdrrrTvvXP26qWjS51M8Pn4hI8Qfo6O0EWklthh4tkM2NWQBayZ/36hDFqaZPuV4
4qDr6duOIUENOuaTClvQ5rJDaojDsz+GbbkGf0I4E2PZKDBGNdGDI7gmoIv0T2TPfcIXtEB+2b3l
po+HuDFH+xqPJ1Ioob1D/ZGDDEkiohE9UBfi4rMxHzp7skSvTSYeWSTEbtZtQXmg9cAOGuL4UASf
jysgmFg6PcUGKLHKHk6D3wbd4NfthTsgG4cJf1UxlxUnpN33h5yTRWrS87SLJEoDZa3Guc++x1nJ
PwHN7ig0y/yv3ar99cpHAToOWS7LzZXwC4T0Pqf1CnlZWRGc3GOmrxtxfKbJTf7NqKF8B2NJEQE0
TR09pTSHnILZMrx0V4NkJZWomqjDgnDGnDSBGRyY16thQ7uU3A5xeerOIjbLvwSjHUidRnIaVQN3
eDzCe3YuRaiFqqNr4zsTFRVt71sDhPACVgbOtmt/Sky+2GmA0qHVcxNFrRzDBxq4aUagEy5D2ds8
Zi3mKGKBlfpEpPikuqDsQbIQArEcM09+7ZBkBGG3ya0KPTh204OoaLaqkRGfvbQsehzbTfIt4dcg
rzgMg38XthDXhabVSsGr6tA+Ytji56uiDx55WsMsRGiPoi5qKnEEoxuR4LwC+5ksA9ThVFpMjxbF
0ULhPUSPADgsH5jODlV3YJnkvewJw3xSkqKOVIdV7RK0sAttkoTSeTJrRx1ORDEVh1WTaVdpm+Da
Z8ve3h0bqjvN4ZmsML2B+Mmw2eaGINaze2pBflH8eApa2vegXHfNRF64uQ14RYDnIjRzpsolecHr
rNmNjLoeISXVLqGwMOJr8PIpIp6rhBND446qtdIiC18Kh4FQvj95fC5mSCWN6dw/XeSlgwTeHmJT
fa1xI8AHF+iUJE0rpoOSEMAnXq9MwJA4pPg6twRdIpllSKN4cMZObiTl7Mu3yKu/lOnHHMNhLhMk
lQerWAxFskS3cFQKJsR/xpkwW2nz2UKf4YobxFG5MPhGfinkAx7l2il1NRRYMP8s9KBVzXwEQspD
Bv60uVjMj1ip5a2yZntTPsOypLSSA8oqUxcREVQVgjAbU7hWV9/b13rFh32zy1yhe0E3FciQv6eJ
qr+/EFnpDZ9+arx/NP1ayucqWQZ1/qhwFnGBYwW77NNo3Y7BugeoepoYffJJQwP3/bgTA8uugJVM
t4/5z4RTrsgHxkJgPymPWecIBFbanu1z4eq68KNsfWmmC40Pz04tztOKhDEwl9b6/TNtStSltcu/
Lh2CKgWdU7IwobcKGQtr5kItwBsh/7GjSrp8QX7wIpLQMK2KJO61YhoxOpasBn+soEO9NPdH542l
wT8hY7JS4e7gMJ4JVEC+Y40kqjHgXshFEL2dfZCPOoYyrk6UKqlJYN1gRAWaqJ3O8RQOefgjLoKG
vMpPpgsVEn8lg5U5nOGnh/kyfjPy+mVPIG0AbTVTAZv98mT2SZFMuXSOKzNEkxh52vbEYdqo+8R8
rGpcySimgf2PJwa3YjlzDDHPFExXuL8/maH8QIt+GRMvSHAE5J5TvngCpssh/m6R9IIiMsql5/xL
swoF+GFZMoj0Y+DrdYMeyFA+kERpIqnx1pSxN6e2tfLNXdt5r1xQQM1mrSLej062y3pI620o1kVI
QnVQ1H/wP/UVutShPXgUYgMQaaM7OABUiJEGsSQg66sORYfa1vQ2tnO1ti+2zUresJOcX2q/4i+y
KeWkg94s4UNyFmE1l7Y6cO/mT5ZN46hVbjc8DNVWlHs0ai9yVUdQRHFne/5ewdUZwkITAUYQWNdA
vRjVt5szVCd9GWSsFmMwKokYQCfO56qyPEJMLjCnlzgv+xA3omYf/8/KEtUgnbSaknSHga+PJSjO
LgKOHTxv4ZFFhBxJVnFs/gMXlHbJMvLllQtGQ6k6SVeYWU8W7l1zzjxRRNklg1ruODw/9vjBpFxF
wonJ1SO9ZfVV18TzLmCN1JNfvPnq2Ofqf5GCqRTzmEsSEfVnYsiKAIhySw9HmXeM6pPZQIkUa/gE
oTAS4+YT7BLF/yHP/w2hxbpmNRic2dbonAf/JujED/+vx8tdGeGeclcyUmGH+MOAIc1FTEYmIQQv
GcUjzNbCl6a3ThfrcKUmeKEeJRZMtVlXq6pWRdLuEqWpXlCpOFnHgRygwa3S1Mkxrnw7mR8AAAsj
O/yzfwyl8b6uHvEkJCQuqlTKy8KmGCyCWiuwtZLgTXDGxa3BcZSsitPFwuLeKpK3SRkzbyhZ6OEo
1KLMDUF5GbcQ6ofbc0TL1egSXmZeRTSMJmGcGnkzbT44Hp5gVvIUXQ7e4jh8SYJkJZ+Gj7Q44lol
rH1nGXv/4S6XLgkbuMrwTHp7iTNP9VTarL6oEknrpHPeXru0z+2hKu04OZu2mN+9a/ILkMGtMVUP
7O5P94WSv80WLm4fgl8FZq3DQ5LR7o4xujhgV4YeLT0sJBoFD2r0QvFR2xSqDRwViiVEn3s2KhTj
YoPOj3L0NbIp4t0ImQVUkj7lBdLJk+XJXdgCzbHVvNdd7nav4TdOMvSUs/JZTMcUPDHIvP4bNEmA
gz4z4g8O19AmFOCuIRtOrmvr9DupDEFKy2jTAv/xPdmaSBYIdqHwepHU0/qlYNOBSDRB8k6bGVOF
dcAZ027a+UPwJN8otISDW7GYoghiPJsgOQL+rYIWTxtSjqtJ0RHrr0o3yQ5s6IjXKIzR5q9czzTN
znweDiMbFGbKB/a5Rcb5hnPQbHZGkHefCaHC5HPTZEt3mUeoypBLi9oQJHvf6ybSmubdfj1+KXlQ
9M+n4Ac3nBNVtx6VNowJnaYLODdty+7RAOtVzmKhq4KdOCgJG651V8w2NWqubJd1MotAOSs5uKHl
VZz5KhVz9Go6PB7sBalK51UVKxZHY4u+c88GEWGnPrKVTN1XgxXNo+Yf2kcJi+2XBaJpY+xrIrq5
eSNV/vOQJQcqA3ctlv2g5ze21yK67H72hCFLSsBpGN2ZvPb/naU2HZbJVggageB2SMWtY3hih9q6
ZZc+cJOxW3gvysYsuskEgiiV5ETMdX+ytaVyCdv6aXvyJXNxkUtf/XweZBqsWMw8aEKZTB7l+sG+
462IKuVNJT+w7/Z53ELpRcCDpOvHdm0e+c+nEEmaz9lafOhC4iLHfOg/j2m+lHfCzghaZ+FQCPle
Ot5eIbtQ03Q+p6an7LwrNWEUJHqbRMQSt7qtCr4rU+uUm8cHNCKxnB5B72uoM+B6x2XLobJOBPrH
wEqkPkP4TMsB+1l9d2bT3gBKb3BTmZOGFiQ9UbfcETpl7izckIWG/HsjvvYGFNX0gU4EH5owl1Js
3TwL3jVTah9NYSQgE45RoDq8X8zeECJhhiXhb2lAyvRncKnhex4dvMnD0jqYrW/bpHGHO9pijGOi
tpVjXcUBgEe9c5Hok6fmr1WlEv0uQdB+FaRQXUmAaysMZTb9jVkDMmLJbNiHdkw6YyIaJCwPEqcY
ouFe28NswwXXuEwSecyzQnLdKev/6v64oi9ptQH5ru3DcsbBNY8ZGXWrnQwjpebneOPate6W1AT/
UgIrNPMgSSEFjS1P4tux+UDpJu3WVQW4VVp4/zCH+T0vr0ksVEXUak9sflUgyjLOaiETR0bvUe0f
HZRNYO+gJyqq8KMgBfvC3/yvr83y+TU0kddIr4WSHfqrMRPIm9+1AdFzk5AoC7JGiEJg5XhtdVT2
JrOuSJZ4SeWWbSlrpzGbqEg5UVgvYxh4WLm52l6dakDikLGiXcPyMlDonW2Bt+GQdyflgsfs6iD4
1xQcCWLPKxO16By/5FF9I9mYFvq5Q6uiahzxmHo4JRUbAotpKdHdOoMXkIwHkjWCLFuxWRlOL+oL
JfV5bBpOlZe4ahZI19jsja6ati5PhyBjjZydBzmB95e84pWnso8utD3Qf+Ynomvxnv0obLRDycdW
Clf2wjhrREb4KqQPOBkz3JCHDJAXyh4O/uCznYTNXjKppv4INAWy0imMiEIdMac16EWm8asjaxva
dew5RHhkcY/h9rj+7OCqgBtPR44u7WoNcqayXWODtYOB7AcAkziEbZtfmgKDFja31w7+IbJNOYVf
VEKtNiZszHSyvSiljdorQLzaGng5+sufYhLjjQViIfKDq61HTOU8feIKDK/6eJUTzXzhhlC18aYs
8St95xkH3r67nVk1/VhO033/5Af/OJDKuplb0RqUIcxBz6xUOAVH1Y3XS87NSLzrpHQAelBsV8jx
u/EcdaB76r0oMwT84cyXrvVAap8Tjefwk+1lwtK+SDPzI5wgw1bBBmWm9jekEGqwpjljfwmX/O6e
rnnKLZ6DiVTrplIuemv6kfB4anw7D1YadYX1S6Tzd09m/25N+9XF35FLHiO+cii0zsGE+qwh/wcr
zNaCfUVwtEP7Fq7uqPjqB58r835d+gZhCcyHchCpzJf2wjVMc/GCbAFMO3BvjRAAwO2/y2is90at
hRvGiSK5IBhTL+1Lw8aVsiCQpDnkdv28lZNN9kf7ac1NLyqGEoRw2p44rQqcsFZ1jW1oF4SX3qXf
Hxd33lr/T2Pg8Pwdy1BmnOThMqhB2mlimbPrqsEFLp6k0eX4TlXmV56TD6RB0SBc9m2DTGwoZcvD
ukZUoNQObu2S/OBiiwFDlPbm/c5Mzv5hOpuLyV5tfNqq+uAtyDNnENm2JVKMKTfcPFrXc5jGKvLO
MrJPMunYiIlRl4TWNq126AO3jGAihPoq9DyFXSlHLZiOg7tsGoTEB8D7wgmqFWotplM/15b9eIcH
LeaCr6k20SRopIgkYsaAIIuz4dw2MBGHN8LWDI8xnPVV/BGtVufuTgnC/RzajJn7jAR2rECoCbFU
I6HQwbPwhuyIt4JAJ19SedY+KHwiYADM/Yfkfl3uvdhv+WKREb4cBRqVGAujHAeICal0avlBandj
6psf0uWSh6tcrW1sgEU4GLrp6UttaVyQix8+VvYUEOPFjJtx7N8ivWGKYf3x1xo5jzx0hS1ALY8T
qMEa1icA2xIFE2rpAInGDwGGk5ISVTt0FzfOsKFNn2WWNCcJJ5wvv60kP5fDXBSKF01Nd3p1vWMD
Dz3zgFgS3jLhb5IRSY1K4QWF9rqtA030a8D0oUtZoMFz27TQxmhbpgV0bg1UnV8CsRWBfjWmZ+j5
b+34Yjgf73Vy9MNk08uD6sbSsHfBCTihXZ1PFc9Cnci/SlYuffeBSfvb1hucNh/BOBYQf7xnJasw
yoeya5P4HRm3Y6IMaGHez/go9+lNLftwESnj/LpFovNeKv9Clb8Gfpg7ub/1jFlQDVDVWVDhGlNN
0nI/7IDWqzir37fnx8iFFDDQ3SKByAkBnYuVtrVFU1CaOuDMTwBv8pCykQaJyRhyK3uqomv/SMYT
k+pw0bS60X3HtuGJY7lcts071qx9JwatCUBXrA3AH2wtWIPOWLPxkBBDe4eSOFJZe1xXYrYmxgUD
KBoSE/lAcTNz+qIH3Ntb9fQAFb2NnYT/mn2APQIThzASDzlM7zRefM29yVdP06kLkoLO1OtSeUi3
GpcuUIYtwe/AhNlBVPNAp+zG/on2qL2unPzWyl7EOEJ/nRZRAgrdWCIP9HAdj2OGyusrauwbs9Wc
wh1crtLpy0wsXiCSJQ4PoUXMGl+QvJsfzM0o9X+NEgtS++cToQGsblMcQunNPpUcJsCvqUm3y4Eh
XbCQlxkvJvWevYvQ/a+RVTQJWHeCzdNOsMcgRgk61lOn8CSPtZVwJk3+JN0e9QoEnxpcQMUYpuxb
Ne4tLXaexJ7NSJi1gxSw6lYXE8Xr90EaV1pNLLmuQv5TTfxGldB9Vq79W/jS3WjMOpUMmVKKYXmJ
3MfmS6FJ4njhOZ7qDEnyy6Jm/XccMGv+j911ZRukaA3SWZlCEoTUIYMERmx1/hPgg5FGbyUiYt5t
f+yhynxAcBSnRedfyro4CfHhPC7j4T7YGnBUV5YBDkjXQfT2i+mR+pzhYkeMBBD1ubeLfgCBr21d
egLI1A6IJ50vlM2RpaBUKq+WtplN/z7y9Nju6pSfNZYd1PwVjYO2wufDz4Ac9mchWr4pJqukJZvQ
nycsolSlQOTyj0kzT3MD0z+sH7XEhAE32cmH42wQVQbG0FwR999QpL9AAqhZAAJog+/PvQJAXZvv
d5yKZxiujxiTJKv71tTpP+E0oIrb8noqYnXuxLVVFkdCrkoZ28JfnsakgAaOZGMorA6ta3G4zO+Z
Y15EPNMf3BHgUzrVScstHgsajTLte6JPZvtwXKubdh/M+TPEBkNvOFu8T7AxUqJzW9kt6ps3stfM
vS5IwvBy5FBIJgpHFsvT0tzO/0eOAeBIODq35sySVrUBKA+i8N4DhZEh5guv/M26ySxS9yAVGCgU
sZweo/+zpcji3zqrsEh+14MnHqCrkyEfLrztYRrjCUfzyOYrMFxnk5W20G5gbkECljhXnyHw058f
M2iE1Q+v6tAApcSL8ngev+0EO7YmLrnAl4/cJ2OwlE+3FJcvTBfFrT8eXpBm9l96tRFzPXSKMtvE
6Vj3LolI7vJ9+UXj9AvOksxqWu0umOkzxViEid2izYnqsmAPal8zO7w/K30LU0otZLQ9TK3lKu6i
mjR+6NCwerabzTaDJ5dI0pFp8cxQIX3Z1CQ2ZvfRokod8lkOvwPWRivuBC6ohUMgA69XdILbahlw
uBrLrSJgr1vMI+qdF3d1c4c3SnmdDs4o73RiwB57do3yuyrhMejfgnpgvzfD/eUhOJgBkpjdmISe
E2ywgTJx+xx7IUGY6ZryRMzryX6r5KvwhZBg8w448s+zb0V2fZfv3j62zxaVt3HWX4DzNody8SLu
nMUr9gfnK+a26zLII8LQCG8pegjRv90+QhfRncCmTELnqfDxAGJ7moBUoH7h4hpxzXCvU4MLAoJ2
dNSlOoC674GreRk3Fls0zpu1pOAJdqOMWhPDLaXGk9VGk6W/Hvo6WAY5eME0r7t0NqQELRrRgKrK
w3fLciA4plpqg925EAk8s3b0fLK2UBZuZbwY0QLhji4+1ph72E1uagCmaCKFfqLXdRgCmg80oEdl
L1NZBdu7JGIieJDxiKHgi9/yQJ8pZ5z9hqvEiHo+Ey80SX/SENLk/paUeFJ3afDJ1DBTXU72dChq
FjHrpv8QNAuiXdzdwYEHC19n22aEa7Eg44diUVHCOu3q7i7OBQewCxyDjbcLcsVa+NMITgxaEyHp
1WzMzMQpv2UPdHv2QH49jOU/KYnghE548YzOSEP83+peYPXclb6wVD7a1f9A0QuVYXlTNZRszhYt
EpOvD/CP0MGm/O49KHl3AD5ik/IK6liJ7n+4Kb/A0Kc5Ca3eGAdHBTXMDA3OyjITdQIjIEAbuh9X
Mkx6RAHro9pUiyVrChnvY6fAx4ap6ZnkDX+qjPj1xsNGChp6lcExm0fkGXu4kwdQ1YgI8gvE7rs+
fZ0ikcVuQKnp0fdC3NWeRiXKe/DH38ggeMzaRCLvS7ahZbm5H8xbSiCdaaGs2c5nxV+2fPyMbETY
JzDRsGgYulOcxPypSyV5LO+obtesXNCiRcgUd6PgUay+QdtV2v8moFv0/tlyR3gYVtYUkH5d021D
jg1zT/zU11JsQsu9Qwo5zNIFtO2DyMfeiUrGs+FAgQXq2UxjL6euBRWqhUEt5qxx8eiHMO+8cTjN
hcf0niZn+CqVIM0tHuG0LoIgqB+lbt52vsktNQS/4ZhoXIoAaC1H+RYtDn6gn8zNN9y3ngoyDSKW
AkwFG7/zNKyH+zASic5nw/3qgSL+NhH0PU+Y+gnsnYl89GrqnOWeeN3Tf0nqplFrGkGQo2xabuiX
KTgC5CD/RNmVYBjVhuRcfOzlYVTu5o4bVB2jalioj1v5N/qZs1FrmhIz9rKPWe0t/KZWLfN4VHmV
USVCxbaJllhMd4puz3PT2/lteztBubtgl3XrPFqBU53YBgNjHRU/sBV9VcqwxyrV9JDBFUhx7cYf
PqfstOoIp9C7SCePl7/EY2eUJvKUpxda+Tixqr+3ep0Lt4iMlHPS+b48MMzZG2TwCQU4VndJuvuU
iTTZ1Cx8aPK7pD+dm1OPAFcHxCM+oWVxe/tkKu+nn8eYDg5Zdo99DLPVZ2UKFkGtrzgXymN/8TU6
euOTtcLFVdWnqGMKk0F6x5rZT9qmUdSCcl+ASFmzKID5jYJzurRfcxQ52S5vbwEdMigFF11Jrn2v
+LBavzKChKo2ZuX818loC5sfzmNqx+IvuH2ZNfv3E/fr7uI4UAo73Ui6WCzfYwIdnsrglwwI4gHo
56ttwFp1TBednxkjq1Y06EDNsXtpGld7lHvoVD6pKoKxZbhMQMb3ErgPCGewwaXg8m73Uctqfm05
w1HbN+YRwG39gE+N/hYX+NwwnpSeADOGnlWyA2mTPR1wP/BlpRZx0B2RdzpCzKkGJN6npaFMgA06
KNs4XNIqvbPEkCJK07VizE4ZYGy9jqW1+yXJk+nNr3QaXw3lBXLP0hAHuljbi5P5kZ83U+IlPXgU
uDfdFrwhDJc6iwzZ7TpGOtcc8L1ndmIB79lygdrv0NLGnKBu2rv3zndWenJtuspEFXl5LUCqYrpI
ehb5voiMYv1hVT++0h8T8ZkWSYnUk1I6kv7W1UZeRsi+EBDSZubj5eaEdzm+EY1t8W1crn4Sj9Zh
KKbSLhZ/oxR5YtdMfzfMt+sDnITCuen1NdAseWcx5vNCLJ0ptBwMwOAnuGuKmAtn4A4WZvnG5L7T
9ErpF6JAaY4QBDPVWwcXTnCoP49JfL8CWiQd9azu1oFDi+jPeYqeku/zc2cDOfPHaOhVPU32giRC
10YSxMl7S+5xD9vkR6p4fbJmfNQQ7RyfRpi9tKkIqj8pIbSkDZJnTbj1Vd/bcG/tbFUGmCNXfjj1
+2Pdd9h0ztN+U3rAqm2aVYIgIeLEJ9baSRBj5a+NSltUsKw02ZRi0LCJVGaBhy7aDgb9LUUf9tcp
Xj61HvAoZYur1EjD4d6ta58ygleBDtKbN70wx+24zSDFcxyBbdy8kLjaNlkgj7qeEUlxNNO8OLkT
k3P4dPJJ2vnT7nU9Xw+O1lTlyVQ1msjXtFe34hMyqlnugd2xJFZR5XfGSxXMYksH1ZRxxnHfkzcW
jJSm65sgNyRh1BgDtqanZOCpG1JJggDBs7JGrvyaxUbfVsfxDhANplpynJpQPdaweOORcjwdA0Vq
AM1sCDEWKdp2BJArK1XSDdL35ntKPvX9Cqo4aA4O6onaP/stGVx9+gJtN62R+rHrxFUombKSTxOa
0T/DstQyL4QzyODr2N+quOmKfjWn8oVBKhpIK0wQIGP/incCFBPXw4Hm2WLJP5YuNiY0Lzz7smWE
GVwhyAb0ZP4kp1X/OYKYDlQ6pEDMN7HjKrU5ML2kKDJt0HOfyoUSEucfFSeSPuQkIVghypBi9if+
BVE9VxgbUi2Ukz32XrZmHTCHoRigowPx+1hWP3RCPbN5kVw5hfHx+9xt39yWUHQBrtBoCQNeKhWS
2QRZRvCKLx0JEJV+036ogyrvEP1vmsB+dlAI9TsT4tQz0SAyKWS0OPHDGLzatuFEHJZqbawMQ6Ob
sofyHxU7ikwChFDmH5VFnH1d8K1vCXTmtBG9LTtY52DNzVCeqLmUfUgz0ePKNk+YSn32B421/sHF
mDCFyVUnTmJr3w4wy2JEQzkYo3rjZkewSXITPdFpUhsBmVVIB3F0G0qDmxwm5Uz5nXl/5vZUY3iw
wqB3RXFPIdybWAP3fXJfBTMZ68oM+tDxDy4Iid/apu7Mdo7YXno8rdpuziWL/xe3uUB5gdFiPg3n
J6voZZn+JxWs0UrIco397TZ/1KLfGsjqZvtaY/sdvU4Ctvwud4lfn60jl4lb5WMOWStxOfxZCgXd
lDSGEEt53Pp/OOZAXANWUekPpVxWLBdPVcPRzcbWGvhF3b26haTb6JzX6YaqdJ/nvHp/+xw+eTuF
46MUPUfqBMOKEUCa1hDHTexhMMO5IplqptiqlkMfRmVXZ0IdIjHAPhl8z0dizsKXlOTyZvHGXHvO
UWhHSXWbQBrrrRyoZWW5vgFtY/y1/03eJSW/BpgEs0GuYZpwqZivn7NJXh5P/Y+QJCVgFdWO7Cct
Nf+gfoLCbX/p8GwuCSOEgTlrB4gocT4zFhpwu1AgL9FLU2ulROwopWCWYSZ2m3QzIhTwd5ziOQcL
t4CD/FZ0P11kDQ/u3CAwa3uFlcK16gaBJiQYpbVg/x7Y1jmlg2Xf59MP32udizxUgRu6s2ztputI
6stBIcR6OURRYg7Q+Uqr76PXo9Mk5jQTLtHIJEtssE0SYIjwVkniNQMBtSaVgtHn25/tzVm8lIa6
PVSmhSiu8hMtVMz3YU6ZboISaNkoMGVGQuGXNCaqmBu1Ft8CP8kwB2uPN+faTCAy5dlhS+JJFkCe
E7Hs6SzbSVFrp+Ns5jca/BZJWietknJhO8z/FmRXJcD/roieIFiEiQHpGLnTcWucXl0RwbZW8CB1
Hhi9dFu8nXYfjDtwJLn781HfhRbXmpwr9rjPyhRxCk4ceu/cu73qw6ecinZbCyoR8g6TdfewgGLb
DPr1mKmptd6Q9cNYYpKbNnng3KniMh0/jZvq875kenL6YlF4zmv1BtJj4O/9p49/XS6lasgeNABU
46htdUnAVH1RnoVYOyD0gsSIy2wZkWiGkHq+KkhVUgp2aXev10sGV6ms9Mn3DxgCeaaGhs3Ir3tV
gqiE69yfVirm9+mVm2DJxNSdLPZHNlzAJ6/9VVJdvv0xB5c6JIcVZZV35bUUY8C4lQsk4kmj6zN+
Ff3ym9STgnJuB/O1lQtKaa4v2IH71KiaCMbNEPaJfJ2cZUuUKHa1ZbiooV3JzxRh5LJv7LvQfB5C
nxa1bSR7PMBJuWXObRCDP1q7jJD9i0zJbn8t6loEiNSzYYhhYFaOWTw7gs+NltOQxK5mJW0ZgDpN
vAUYnqdnpj2CWfKKCqtuzsGbyyg1LYQkh8pgMBZUQjL/UGb8UaqHMr2fkh54VNweOJccekSfw97Q
tZKXKxm0JeiBqaCi/IfAJRol8jwq7DGErn6HE+BB93wcTxme0XWyUoj6wKdAi4IAzLfdwDa6TMUB
JgfEKCKyHd1BttNwkBUdEwuYYLXyGJYvD61aLxPtSZRyh5/CZV8mmCq6TlHqFoPe0SCwNROWmyW4
UAAaRwEn46UAy06RHCNMsXF8O/aIjV6WakLLaRfVUPcMA+6Yu++CoQVPh2hz/nY6kFT5FPol/Q1l
YcmCR7W6m1gN+ys/+kpy/YzkVH3R1d9u4wVvJjLCM4JF3PvZbmvU8Q0XFVbMOJ9Sjc0P0q5GK4Ro
/ktkmyRdEnx56Q1iRNj2zY/wTQN/1rAMDeeD1G5D2odshUKFrZSFNAbdDuIrQYz3ggx40zaZwJD7
0NhEillwxRWWisdskwkUpIsWt/VViHQMB9KFz8iwc4N5RXpr4h5hiKtliN41V5+MGGLysP7tpcPP
pyOlBBoMhWVswCccV/5AppRl4wgDG9GVdXGkkNhshoSkPSMECS+X2e/obWxgTk+qGqjPGXS4/gI6
rlazRtSLgmJvC1Vqqun1K64ocMba328QA6OgvYDlhdf5rzD6TFODHUvoHpglREBr1jv8WqifKQGP
BBr7slWLshJU794AtXtSAxW9Smsb/kCcMMk42vctE5WoKNCxORLLZP1DJg9TC4BLj3ILYD3APAGv
WvgRbta4229GUgBtK8MDIMRt/cLT3RicLt5V3e6+VYDoI/R4+ACkxt6lD/EujSZktR6NbkqfQF3L
e9LcuqPw1kxp5+FrK13ohoA57AUzl7UHFvTM+Fqtq1r++ixl7GjdjRU0tfrD1qerEh1yTDNy3KSi
iTIMeMV22Nfg6ltVd4v4d9k5wht5QOhrrM1FUO5z3m8VGBKVvld1sCc7Jnk8rNth94TZSYEHVJTg
WL+8Bi26+VbmNnC4PFFv9fhyggP+XPMcH8pvn4bP8JZ9adp7N1iw88w0KgspTvA2xcMKipeOASWF
gZwQ1QAhMDZENaDRitUwooMLcD8jLE/q3PFQYVPWPsUViOSCJDOuHTmw8VaFavm+0x4/zJDKJeQt
el8MxCZStXsxUfEQcCy0PlLuI8QqsUOOS1Cd4CMghjp7VY84KYgKsP6jq2/OcmMmVGWFx1V5DVjp
xyabma9TZq10dcDx7IYzq/qV3F9AUNnXQtFV02pRdj3HVLzhUGltgow14GRtYFqKVXNfxG9kCo5a
GPOoGxUfsU0IR3+JJomQERiyFVJY/k11Ads86osV+iw1AlLjXk5I56nLH+gtHTGAUWdYuFFnLzRz
+JXdigNHY6eMkc+hr1VdRf32VhgfcFjE8BHgn1ue0GBLp7B5mKSlup7TZBZBKV20sjq+xZIw/a0s
sXv8dEM54AvyLzMlP/6HgdhucxaJmpK0o5/+icb5Q7rHRRVpfrOvjBTxngVT7jqv4WvIQVcw7nYb
UQVMHBP52TiQPe69+APWh5Zx6u+4Uv0l/hkWP2rcoglRQ902hL/RAJbK5jKrpHQ/BiAp5d+CbXQZ
hVSwjeaMIj/W/3FkOt2vBVy9gQ8XFgNunfpNNap91UfDmoAyw3VL4ikUac3dNdOh54e+JlsvC0aR
PO7VN1+lOQ+hKk6JlygEMSxW5hBbVUO9mmv2awQ0IQB+wCp+cxBrnPX6X1HI7SlaBmWHG7Zh693f
oR1+jtSExu42y3nCGF8DkVu0LbpeapDZEBDVyv5INq2tuFaltmannMtFs7OTufFfRAOE+pKMJGtm
+JWmQtSzVMlqD6I3mDkY6X5tpIK5lgBFXg52JiaC+4v9ktCeIlvid2yaq/YpJKNuh7IAq7Mv3LKs
VGgB6yP9Z2xU4+T1cwdSGeiLC7XLKz1E3RrzMVUV6csMDSLfAFRzelz+SxLMxd26Jg5NS9VvQS+O
rchMkIwSgMfzZZ+nyOapzNjeXYQS9L25kcayUs5cNRaOBNBpD5m9PP+jipPVQjPm7VK71NhYW5fG
skDFyGCxQqVxCpzFX5fLxwGjQNTR+1oHCnt7k0PJonWToTpxjy8IJiSYioymiYW0FeiDlOt/l9m7
Z0KFCiScGozmpQv/+SRQY4V7Jprd1OFePTxnDJSQNOmFfuWJ2tELhacDBfEXtsNqY/Bn2scR4p73
Dt78ICKHXYHKh+ZFPHgf6KoQrLD7EW5Bf0Kw+4O8jmCJXshGTf4eZo0vBgHncLxEN1eTiDis6wsA
KYZmwEg3+OGhmUwHsL+bGfh5xiO6KMJX11nehbr6M3RM1TPaYlWyUSUQ2pjlKGXO845lID6XrXMI
le2SIa3TCG0Gv7L1Hi48qbxQAOa+81AMpSML6S7CkKIlDw3mCXdUfhcq7nriZUpL6C1G/mxJiaSb
c0WRzc9pDUClFS9sOBepJdEMxlo+JiKRnSTHodX1SoQ8nVD73A5zlk7V33tfb/e4TziqYK+ZDnc1
Ol4NrtLSbNdSWB8rx9dxTdQ6ms4+wng0aG5ulmNPiVIjUJFfE+9A9UhyQ3usEDUtlQODA4qXImQs
pLkXAzrRKB2LhsiOySyFBpb5x4STfRaLAdX+CbscOZITY9JeDe2BTTxiPIwa5NQOQy8MpwPeJqEZ
UaWltVKuyNyrYZ3umKZRL5n9xEIEvSHxq5JyrgRe8VKlCkZYKmrYvdzmK0bxBk8cyOAHda3mzXTY
ek1JRsEAafdi3iorDRJMtgD9T9wcBccNItuUj8rk5WHsjFH1EzbZt6YxdGhjwXEE+Vbia0C1xfpG
RNdwpf+QiYG4LdKoYQbcxi3f0ekVfdWLfbIB9sz7/ukVW6qplwwkgJdWFwaSUfJ8alxS7+3Ddlch
9fUJYyI4BmqoKx80TQnhe6MfyiRmkJyXV6JUKRgPb5LBROHND28MKtDScelSnHH9UBcmVci/BZkn
JRxLmAaBagoa32YPZAeWHTsnsF4bUKWJH/dU04UVnllOd9ePr/kKzgCPlncPDUIl0YMmdCecxSiQ
krTYEwK7lYJlZmK/q1dJsTIdwtpyMsXE2uJCK8BVv+mn515c3cyPBNqkL4gKCzMTs0xA+JsBCnfR
yIgn7CBH83z1Vvj35b41qZb21CffUtRttht1T0+2ElK9uKRQLLEtTeFphqT/SKg3DkNysdEyw7yY
DKmbHHLUvdbLQHL+cVvYw+LAacsiOSZhQ1kS2IGJI9BGh2umKW4QeToBpCBXdeFtuposDGeSiF1j
EPJ4pMCfprr09Y+9TNN3ACo54sPwGCat0+zgO3CmxFZcQdzWd1uLsRauO/+hzqSmRbFvwPzXCpnH
gtApchZzDPT9DvpHTrSCFAUP1j4VIgIdgLEYaQA5/UrdbXfyW1jk8WcDZT598NfP268jqwaluPKP
nD64b/F0OpQxMmW/u3XpUle+DuPP/bhRQPKtGPC6n+0M45NGGDw0mV68hvd8vo0hLUwvEz6v/h0G
X3nDZg2fc+0Hrjq/qr/Nbon2DfRVqvy9FwLb1ibBS0Q7vPNmgVZFzNR0Azwl4uM+gh8NchfhJEW7
2QF4gilUefG+xZJwXrqJ90FTr+2pTbL65qniVPB+cytVx0A8vNnrJ6Ty0tGzhERONcBkWsVh9ITj
lyQ6XVDxITQDPPv87J1Krq6fU/xFZgqI+VbJGuLmrSsiikGKxQexbYSjTZESf86PQyOH/01NvRHO
LCuXBrb8n4yoafsUL4o1+fs2SRlE0FBoEPeZdk5U/fij8VxUToZ6ivw+IKo6ZwF9gza37jj2x41C
xP2KfDSId/G4DaORpykpiOZ8m8+H6pspa56ZfgLMpNHr88gcC6cP/bGDxn5rzQdX36Rcw9bjmKIx
YrTNPTAdHnq0Hb5Auqt+AZhDKl5Mrt06mzTx8msxmV/WHI65tMk85l7zTjaC98SSyXO7DhEMD9HH
bBfFyew/JSDosyBZJARpKnS989YEMQvOwx6MiLY7uQeunpYAVRkSel5SBnOhFKDH+MAHnVuamiDI
yptr7pUm/MtcAtm4HzzozXNT9oDUoivoTm3Ag+yNbkfRZWyYdLchgWUmzG3mB4oCT9pVGMQIEioa
b00Vm4V/2fST3laeSjXWRw7jMX9a3RoecmqtSUMjcusoD6Y6AWDJZ35z484Esxb0wk0U1/cjOuLp
Pe8U3QAoupcrPhg5h8kllHeEskirf+8giVf2z5pQUFZmfc2zX6Gl3xwN6esqXjbuSFDIRI2bVA+h
MGIb3T7iPNt2C8dFxp5gBjY7mPtISafrP6CdksaGxwNGCLgDPIBRkeU7oTyTHmnh7GXgITDbpgP6
Qf0aeWezgZilQ3WH7o3VmdhtH7hUAMPyXi3hRhrVpvnnmAFg+yJo7cGd+XWi1adbTYZFf2IpYWBB
O2NKmyiJhhtGZMNor4uP0dUcPeMINRiWB9PcD42KQfOjZ5+x0XfOPj825nJcDmS7kZh9PFcAZJoD
/Edj0n48qKMBYJcnSUtsaaLrO7tB4UEWyScltoUMpkGTt1d+TNZxNMqs7Avpi3I0jMehwK0DViee
l941+5AsHTu6BUctRC0M56w9pcah3As9VpTUk7RzU677yB5jtHZDaJLOiRMQegV7MX62I6EdKr1l
NppETjXREwmgYIB0zmLspuLNhY0mXk4w+fj9HjW5VEpAoyACKUtRG4XjuaCqdi+sS+j2s0HTU/UL
H6rit3i3AxK3H7rS4MrZd54c0B5ey0lum3UuPGNdl0DP8KKg8VNK1hk1ByxRqUZylS1G2vj94GLN
hjPPXOIRwb7J2ej65RSufrj0aZo3SQUZrlBKQKZWSLUfeEbOq9kuBzNYqNceo2IZyLzcwO7aSC07
R6AWTRXbDLVTZhu56YCIL3AOGIFOLo7ZCiTtBJ3FegVrzbzum8A4mye4sZ5uBarTapz4ZZbgj9ye
C80U9WbmT+7mL8QPPzhJ5ptjY5AMqeGrz7DWrlxtdS2oUP7HtDxhuxn2eCho4nnJSXGJD42BjlxP
JRKVwWSeEPQ7zwoMznQtuskDENxOhrkitudUeteu+RW4bjzFIqA7JVjF6W0AGunqjZpUY2h2ELKu
aEWbz15Cd5zrm6PF8BIvAYMeR3UPPLLaSoEs9GL8iMK7C3ip7VQXon4f9JFz6CqXUScmRYFv/6Iq
F3ul/GOfxNGUxP4E6TsJpqXy1hgFhHXBVZ/cjfTve/aKexTAe8DSdBtezbrWN7yyOqF7p7d5sLEm
VNYBOJtWA9DYYbcmspIhdDHkbfyZd9eNQmGRqk8Pz7A0kJkG2+TM6PI+p42lgNu4v/xtu1Frzocy
lsyJhUaJNAcP+mqP7OQ6ikA57I2muU+EQ4iLMO8gmWL3anx1pQ+s6POn3h3oYvzGeKT77g+BnAZz
vWYAuhHSgzVKTZ7P3gKNitvHnmv8GrOzmdwAHT2P8UrkjXMPuZQi3PapLf3A2WKvf/3CRpeH7y4r
plYG1i2uu4bHrAfwtP9dlRgmt1+h2cz6Dg5CYX9F+GBZb25LyH5k5zSAXzvqx0PwoCUowjUo2JtT
ylHtFdoWYy08ghO9trI9Nj4gfie0I+h9AmbMrGe3AuMRSF72KVEiYilw94DKc52KAGRwQmTi0aM8
RroWonercDi5AtqK8N9+CBfB+jSd/0fHjOihWbLREzbPgILa7/nYzhRNVmILxJPCONSsdqnVtjET
c5XjVWGlHhW8Xv6z9+BdRHdU0V+QhF5nhurgvceJ83dJJCQL1/76GpJ+Zej+UWVBH9L/tiLKo6vL
66HYipzR3DLcd2xq0wlyodCuQ23yZvIz0rwB89c2xN1Z8caWmnEnCeU2EiVuzXngxiaDFHveEoFe
aqXLaRTi6XrXqxtY/KTV+Ic1uozYP83HmYBOXBV0N/g2cxyuXfvMLJrME71WTfoudHINU6/QLle1
Nl+M1y9kKAELm08/+kPUXiOKxdm2fveq0/OoH3pr5h8VOmI+0BEcXFT4q+Wa5XSCthHQ+DxnZTvW
ZTKXfkxUYltC6kBzUN8BCexYHnStdT1btQyD+nnXIMgnJ3ihLiVlV1q5kuna4xXE3yVVhxCighk4
HZkITCVl/reCi1stW0WUot7NFRNK2CcPN7mVcI1d8LyErrawCgD9xrthaD30t1fHPQJSkbsrT3rb
MMTWF6QCZinft3/n9Jp1U0z/wgxU5I2gGpGQ40zUx0GRfzMUsMDHPveQcTJycy8vjWdZVGoTXsle
uolLMNmw21gIUTNTOcbDGNVQYMhZcU0Gp3RK2tdUnMRub7FKBwtHtFdrTPtGEdq0mvIdWsVKpl4V
Q7dl48yMOoxWJ58uzCGxbLVID+g+4i9l0Se4doNiL0dbYz2J4enL+3ZYuRKxFPUjeKLOJZAvbwcN
ebVOx1/y0xk7HACnRQ5mTF5OnFK4WwTJJeHZo7JMovYi3F9G/oVDGtGps7rtZAj+8QfZ9ggp4ub8
cEH4zMYkl1fJ6AYv79cLx0lOKjRVulJ7ZUhiqpqVReAB6lIDV3rN8KDFZ4KiQhugo1U4KBZpHwgs
+XKVnvW/LnCGdR19FjSY0T9f0iBLtEwyXfadIHkkhcQaCd4rrJJgu0ABsQdtJYlYa85hYzRqdQfI
dYe7OhEY8FGT/tePTomu3uxsU+pJStdh3kmPq/pavv1/gjgJmd1fwSh2UfaXfPp4mhGT7p99v7ar
WKW+NMBcerMeLRiUadpA1LqEpA9N+fOEbvfpR4h5B0nkWMNFXsduQUQDoPZrcKU0Bdlbqg403EdP
ZQvGj0h60iq02AVluk+qPSW3OQh7CmdYGcagw2K9ntg2ZMGAlaGR3wET8hMKHBe7EKB2XCO9D57B
BfXcYiMnekVhbMmnIQvUSEU4h5zeIt3GZC2WEGlWonm09y/KCP4sDCzHJOYZPTcjZL/l1NpyKpeP
CgFxLeF3E4HS+8KDGqBq45ZecGl01V3lAUUCrkBIXOFPmdCOZkoMzwPsNKplcLSQmZ1OjA2nL2ye
4HMfbFxynmk777Mr/SztAqhuG/PtdurnTNlLKne6QFc5UkLLSVo/CyVcCz/cEb9gDi2aVKHV3SxJ
uzupd2suILuMAo+TYa/U9idejoNXNi47BKChLekEYlwcuzBzetTaPGks9GWHuotQAsIaeUtB1rWi
5c2nBuuVOKw7lnGgcC9H6r9N0Uu7we+X/ysaLPUp0dskyOEXem8810XgAQd+O2hHjmIZyltPySZg
q0Y3pHWIilsR/fIIZCqwW/ZxhC+ebbpbSaONFo74dd00d+bv0fOjz85K2DoiAlWyWcsiCjTtExnx
C2b1xgiXLDOk4zbECuuaVl9T0tuoAA42sl4meGxssdwSF+xZms5bobswDA7+kR5vcFZleSIJamfj
yD9y7CmVDGNviZ9fLEtGBgrqLq89KzzJzGQYDzi68fhyc4TvYLfJT6MtzWj2493/itcUwSIAyrXh
0wgaOpvDKVIkvdfd7vrFBek4ZFYUcoU4Zr1w6pj+BRyA8TVQ5RHk2Kq4k+V5WF+ysTWDJhVEWYiK
uYNi2tRnXf89Ty0tlKUwhU0mLoyIFzD41j19GZOFOozYPOMZ3ppraRMxYYmiSMq/9xDnzrfowXz7
nbsYm3Zxfnj7rpTiEj/IVkQqxQL5IHjPV6gpfDXJF8y96MGgLF1jqks+P3bXCo8GKNJYE0yOZJDj
kiMk9LD22bFYti8IbYywtjCmId4uR/K84UhYZfSp9HBzPcoDwsRT8vRaw0qBwS9AWRhE1dP1aux1
2rfAuIQNdujYzf13a+NtfFpEUYzhF8Awo2rZ8rgx/qyenVmFXzy1RuquVcZmFRlje9bPDf0pNiyH
nXPnJYUXxsBxEF8dCjof6UQ+c9SEjD1SXikUnWVZrdRZR7ZJXZbjMVHebRTCh3ZT+ZwadDXwxXPx
3R8bYJabiK13yOvyMK114S2uU/e3+QkY1iutE8UgYR6fjt2VvGTRCnUsCvfsCFI7mSRcp53n74PF
3+sIxGF7AzonvwA1JPvmyMBxUi5rEzTlMLoWNNB4m88TQ033J0hm8o4h5rHMkflk6Y75/mIyNae8
Ezvnd5GsvzzovQBHCmmSwxawRtdo6rPaxd1V+2D8M2MR2Xj0MeNGVtxQHC1ChGyjeycZ3Q/gJknI
plG4kWcDL7/pKh6WvFad1I7SD7UhIe7gQWtPgqgse2a70CE2t5eiGWd4HGlhlG8L+PthYGo1lQt7
sqbj0gdAfb4PwBW2VgHlfMVcYd4qbIwlYrC261pt6ENX2ml0DDiyZo2XdbEykWYFDgCQCOSIyv10
elW4oGaF/uKwrbh2Y+LH3LSm7zZ5uC8GCbQXm3tJxQCCiT7eMg4RV+XhMeQuToZetFUZPzbOMoXw
oot4bH8fCztNM9gARsbbSMQtDLgBcytX0h0SjGDHyTyRnLZZbnYfCPQ8FU1g6/JxLH2mn0Oi39Jy
KSp9p/4+SDk1JVMw2ffJriS2DcbhCmG3uapR3OV3ELOYXE4iD+2RJXzvRNAcu34NOLGKM8JVH/Lw
9ZYr98KwO6eK5BHnXtsP5Rc1n9NlbMwk/BtN6jdLRsEmVQkhXz7sBglJwaAUUW64iYSejHgL855+
rGE+OYJMxm4J2atK91l/0B7zxiEgE3/tmWHWEFLJlaL/MlyKy0IH16ZwzI2Q7fETB9hSP0Ml+F/h
m8ewmhIbVjua9w65v4GMsJdX7rb1/nyHREh14sDR5OwWFPGSq80c1oPF3sRDYW8mB4YeOX9zhq5C
FPjWEjXzCetFmjbiNfH+46lzqimM+sT6RxVbDy7VhUE58sahBWArYKSvR85W4cg2vA74GbELe3ME
DTSoNYXNyRn9eknyGB00g1A+6jZ/5IEXa8ySGsHahcM/ey8Ol/h6UUu5QhD59Iw9f/2cdOqZ/aYN
2ON1Q0okGcr/LIWhyRnBpbfjD7a4NIqC/FGlWm9Ww8wd2mPa1lA+xg/u5fIIH36Ax9nqDBjmLLwC
wPLrCYrpZV9+b+K3DIp78NSoxUNkL5yWAxjwlI2N60C/ibPX9IWh4FD3MYQAmohpA8JkuN0zZa8V
7ZHUyWOAecHcxQxft/l/zf9/CpJRK8suFzyV7y4Zw6xJ74eXOJNIWE0+JsUZuOsAEIvsDBpXiC08
F9Euees1C1f+EoB1FVybkq4OUXQvO7xQ5tMiiIKDgvK7jOl+ItQ/4sVjwPwk9DUn58xGhlj+Wg+t
7m9QdljaHg5k28RPsCoLw2WIYUEgf2WXP2CtQvabMEgTjuOxyq5CqeX+OYwQdo2/X73184TsKfzV
3huj1WqkXHuKqxCn/IfzsBtcSHyxZs0wkihm0DCpHV0XNRTlfG8GlgaIQdIglES6YuMgS11n1CrW
6yEXh8QfmMkff0fsgvIi8u12bvQpNd0tTvxa5iGy89Os0HV9nDSIX8LdgqL+HEGpKM35eo0pP2A7
xhcbH2fE1bWCsN9U1VrCceyW8xukEdFujzV8NPQXLR77eG1bqUqrZGbShxDYmkWmZFGmn1iBiM6P
AbpqQPgNyEEvIv+32ZuZUWF8x7ySeaPCK6pNPp/wwNAU96rbrPsARaZ8klWBd0TGQnVUQBfOiY9Q
d2Ta6rWyyeJeXTYeidJcrRa9iO0Xi8UK47Z9Cl1Lb5kEtFH6lnp6lKOOEcnJovZ7VTS6TvjrmGYo
J7eO1fL0l+af5uD4gDeatYqodjVru75E1e0jZkUVsAsSDoeC3Cl7bAeYFOvrV57ac2P7gXf9bJMv
ae5l418Q63kfZMZL90hcyNAUGQuMg4Tn3SJ0qb6kfdbHeW7xR3FdwoBpWSMWIC69yObqADlG6crj
4u7Sho6YR79Bz2sQIvKly/caSoscY46QwMYk5sddMoh3RVO5gK9xwdkr1bzQLp6iCYkx1JJlWlnk
JYpJajGfDwrv+FlZ/+sJiR+xdPvrGMHTZ0llb2LaItSx6hrRphb8hpq7kfGlutMyw5nt9t6ler5Z
0+lD4Qh1Xyc4+5P5P6RINzF2uYB3EhmWejQ2MrBE6A4LcoSjQgd6saCrRrS96XZlP2Bhha+QY/uL
Tb3Y283T9yJzyFKobUCYwU2BKVhl/5hqa6mmYw7g1/HYGjrflv1v2x/LSV/iVPZ4TQ/Jchog5wL+
E1DvMOw7BENzPCENICm1iuhsdHo8XHvHTzTc95a34Kf6bm7LpmL3rrPzD7lTQJNQ0v8ZRr348n9n
Sd74rnMSm38dHZP4XgPpTfm0dWKPLi5F+1Pp3otmTEMYtpOF1scsAWXp89lXgpaMoj3kSIdSNfAQ
8VrezNGVfilqS0HkhYfnS3Bo1pCWkBJpUELFoVeWezseICJ2U1Bbh+lqVsZvdWTl2vlH4Oj1zRQa
26Pb5moHtuFLIa2Yj5/NszdtrAHIKoHckFVQhacc6Cmvgxxs0OA5i/f4FiLmGvsDa37NtpsRxR/g
ab1Ksy6OTYIKdutXM2hNr4yZ41lZu3zCp6j5BTgvyD8iBXXRCOwcBqOPNnPXnvpZx2A3vSzu+zpN
B3WvwmC4mwTulxcGUS+JovR6STbz58OxKcS0XDqk4G8c9lpCnDjFvEcKzcpkX2f+blOgDfGD4zeh
kN2dJ44/fMkyU7EPpHwalp0I1HtxPTroOCFkbJIU9Xa4OP03AO8imAVIbO743ib/ACjW3yYtw1JI
1/hRT0pz12t+9LMJ9d8I6kWGAS8hbERLEve3NfK/ss8+7Y/F7W/F3cELRD0jnLa3S5U5lQvTZ1nF
mZcVDla0NjZLnMh2pL6UQD+zZPGkeBPgirh3zUOOnLah3w+EIGKydy0wcOGsYZH8PYQ/NT3DEJV6
1T7qRRnPc/f12Q+PsnRPK3iY1A8BvJEUDFKw+/W8BKYHgEPa/bGfEPU6nC7usKdSEBmYhPnQ6+ZF
JCnRi5aWezhSgKj/T0ll0GzmYgF5RsrhpmE8HY7rt8Z9X+PWmbN3N1qwDr6URYfa5Gz/oKGcVA0g
MEEUyzNQMoEcq4KQQ4Pa+TOiX+PmEeeK1vL5Yu3dEAhoNikla1oxenlG5/I5Dh7tepazeVBuN7D4
FE1XmVxqoSOU5S7e06AK4UohBvKFga49+Z82WkOfFlUYwXW336V4emAGaswhcBAqVJcJyY5SXtF2
B4/i8EBoZILzu8+3WaB/Hb/GLjEmvVYJX3+dPNSEqMiM3hngQI1xGkObstiDSFnfhLbYEkY/+dmk
M2fgABGgm+GrDi3rDTaiXMX9MAsb5Td+Va0rGOdaMs6OaFqZYPdNx6TRTZJ3e2zeqfm3L209BbGR
GlFCDUFghCuGxCExCpMnWjzbWaAnGClQjhXhulxOxORKdnHkHZqA7nr/QE1hwKahh1rPsMK5xgXG
2Bi153Hc7vyhxGQ+P99XtgV27aoYbiOJSVvQ2rddwKJ0Eb6QzpFgERb3za13LryHZu6i1mtl/jya
qZiYwyoj95fbzQb4/402AdC4xqaB/CE8nLXihxZ14FhR2KLEGQfzy9u81gKD+s504j8l6oRJw5sa
h1baJlPupsw5M8Gr3mQtr2uEGE6GnbTIdwv6vtEUIu5KsSwiGsRgBUbZgOrJvwREXTivnZExiCg6
slnCA1XJvbS6oDLntjrKqgZ38qWDyrNUZTq/Ln8OAjaOXV0j8MOb/Q0Rq9VA8WoHD1YVIkDed7Ol
6y2bcf18ckgATmr3GWxozZfcNs3Qy3oF7s2LeLGqPmmntFeEBYoo8MUcPRPf1GjcoUg8NS9X5RUf
wGkwWAvDMCN8HF4PTOBSva5QzIMe+uG435DWZN7GwHvBxOle82RSNYm73nr3+yyzPMNAuX9R+yQw
gfu8qDG+uvpNli/SppNuE8GH2jqOrO3+5j9Qby/NAF24iSc45WYltqpEAvFj11jUTJgoygv0qUFQ
H3/PFrkInUmLTDxf4ScBPlIj6k+TlA8JX/pHVPFKsOnQ/g/CNjK4R2VZ2XWO4oODWZnC8gnKsike
7fnoNuOtw6aASKaWMB08PdjOu9hZZHoRTo6/wb84kiKlS/2LCVkoSHOCN+grYFXPsaICtJ8w6N7p
QxU0L2887KYBOhaE9ZRiceybz5dOQxvDiJJOqjp0/7ytysTvsTpSXuMaL5tts3UJJkcO8dDGCjTg
2blJXtYEJKOklIixa80gcnbCiokmr+wz1I+rsI0BepC4Yu31tOcwaWvO+jlRj4E1hOsH9sM+pVXf
zFbloOMCLh2GnOSdwQuKlySdlOsqrPFUM1kkODZ9CifHiBYFNCYX0pM180lNlPZStcakedJV+AlY
Io0vINFCKaX5tsT3F+6vc2GZuKLsGs2x6rj+oMsssijWICc0b8dTzQ8tMq14N765//MFJveKrsjP
bNELe/IETItSB6gIshP5Dnl9jTOg2TG+3xGwB6PX/9UKrafndJNm0XeTEjw4VxlKwB2LKH9dsQQH
ZfgOdlskk4OAW9xmaTdMtn0o5r9kLX5WZ0nk/skz5Lm1a+I1UdIv2bmmhcnU+FCJ9yOQyvpq2axn
QXZPXxFcZ0egcwdLHV6AvSJ9IJxsqkhLKiqK5tUNyCZlJJyw97nsUlbTeR5obzg9gQwjRBbV7m6Q
bM8F5AfPqncwai8notiE+KmmHf2mfrLEogfncThhhMrpsRflXMzEXzsCUtP10OO2tP2EfN5JpRj1
2fyIB6JA+JI09MP69gKHmPtAmyQYE7ypxp06YhbUZKlpMiNnFtCY9eYAt9/IMOUEyRRv1uWcFD2o
qLd80mCAVdk3dnNOocPzG1+eVklS6JA77ixITV1IVNQ3eaVAegmlv11FFRQDiCb5K3B/hznoVIE9
c6juLml8gtoxZHkMAcv26P5hfcaYSYjptOcex1OJBLIWcw8SurH0cUrMCgneeJV9NM1h/bTxJ8Rs
YpMkpF+9ExrsXrqyBUth/ZyX7omF2cIIRFBwUiSYkVRQBLxs6B1Hon2WBOjaQ1LuDG1jDRLBWQNl
PjPi22EwpYHhiDWp6E5jh6Fta52y5B8fojGUidnf7BfOfKKvSvocHVVq7EXDoRZ+eLx6D6D/Ar/m
vzAZObR7p2z+5Maws/bLCZ1u9aKD79UhSIcQFKk6Psq3n5OP9nSfoxu0BqPSt18Ekhsr3JtUXOBu
6SYk/RF2LnF4vozpc2j6G9NUiwmtGgex8tMJp5UlJ8o5TTa1Tj1ModhvLNbusLI1/7kDuuMqG43h
VJFBEFDI8Q9xnutBBICMv2dUotJvvQYvsXnqacTQ4DZkPSAFN/3Vf/UvSxfmyIEFTuA7K0Et8Hsr
JD2tuQeRfljNh2y+5DvdDvmaZbMMrX3YMP7pFrEKxlUWwG5Sv3xMjbraFlJ+qIk8eilXoTKy72he
YYuKNAQvt3sf2pzx8wfJ0Yaj+TBQJYO+N0aNzgmRuKLN7ppTRFdizMpdQNFCkxCiYhm8Aq5nLMGF
V2jcjxeMIah9a88h0SNcNK6lHztakuXPQCz+5msLh8nMIWtAEZkU/SWkOMTPATQDg3zzhpeu4BVV
c+Gi3qQvC7oQpsoU4PiL9xTPrkMZQ5n534jIEn9ZEL0V9oQofUh1UOmmLuyvL6MPNVcpZBhfaG4Y
lnNaxTS04+sLyc1FXVOy78EPkQJmHFsXDITCV1HYmKxCMRqBX2Ox07q1nBI4fzLJroSugZ9e98Yq
ntoTNmO8vYAdaYXNsShwG1PGLfLR87f7AXrQsN4tBLKAs9usyW4eSlvGTZXDsa2h8c06XDNQZS/F
Hfdkb+Izw9XC14b9+3YZa5mvCkSpSkKICPs0CGptHXEp41I5tTI3YpVar3MZkAjUSc2yCAR8Accm
I4nfiWHNlOXmjv4u1z+wHnxUIlQqMb+4Lh0fJkj2+DVu5IRuMq7L0AI82g+c4uwN6ydOMWL4ZvgB
xVj9bXWN+mCwlO3CnqJqKVmlconLE5bPCtQV6U9pUl6/R7gK0s0mE3eYYjhVZoYWUzYpGVEoHupw
Y/S4T+xcdBH3j7KGIv9ToL7y3ig8C3xGtPBEoVZPLIqQXddmPAJOCPwqUB5Fga3ynB/CKpoBs5RK
jahD/YDFVTis9dt5ezxpHQZqdFRgibWGtYueZvezDXIoQw8+PyzM2lIP7xmFiHgXZT1W+sod15s5
02pCg5gc6kXm4ETXR6D2A0Owvin6wGJmun56HPXcpzPNYZoUza0/VtlXGcDu3Cil3E/atsq/KNtm
MPaOVuFAW8d/LJsF0TKNjLf9xaU0RpK/97E58zEc0QjIa20Sh1NvsaphlWJ5+YIb4rD+aPW0PsOp
jDUoOomLU0mD1+qQHYaVJlpOnBxBt/tgLC7o429D7s0AQsz6ZWwNR+xnJvw1yDvc05S8yd/ScDfe
+WFn4aCYbKZIg95DtUcIfbee9H++Y+4u2FcCed+7tBqrhCEhA6Pl7eJFTilbP6oaVsuCTF15UhFZ
9gs6B4b0616Za53Y2r9ZcW+TiJ0lj8jvMshqfpmNJ5utB0K2plMTB/GI9V0AJuGeioVrzWQctBq1
UmCu+mp66bX14C2VPlJNgP9Q/APN3wX+1atysBJ2BhjKTlaNrNsKZn4zmmZEotIOXcniaw1denX3
CNs54aawozff0FwyHxc9wtXkWiFhN/UwxhHgRftDmb7fv50tXv0dUvwB4H5hTShsqNPqkeR+8l5D
P256PBkq5vcapS8DqShe3oSMgtqO5zyQYBA2JnQE1wVpYC7TtSN/rziAm2N7yqn4kOL5cWGwJS18
uFF4b2HbYJvPSfpIAgNX37dHYGSykDpVQ9yJ/kbra6T08mz9jHZ2c9S+QCu/6DNiMr2ctpV87bOm
tCT25SYbzlUde4ASlWwG9DhK+nLkrkKCbDNXbbWwASnOc1j0llWXjYdMRtDKJzwPVeJFUOcF4uf5
pEiQQdgVI4f+k04jyWd/WqdyHE86LuM+VOQtL8IzOoFlGVEWUS9S2dqK5SsyfbDiOdQOybSz9LZa
gF4aThb5nayjS7zrPE5Setn3HCmPvaSW1mU/Rzg8Xxtmkdkx+GMtg3gedXZECMGJYOWPqJ0rJ8g4
Kdv0uFscpsbdFFdj8Bkih+ZK3irOc09qZ/oM0ljSrcoFlmKdBVBA6C2gpddTEvTbU3yB4NFDYSlv
rqx79C5M6yBu8RXuzyk6bTVT4b28Kni9aOGtNfpsnEzt9zaj+VHGdHYt7me0zVGVD2Ngs6lJ2gqL
oNt5ozaIZPWOEJoiIz9jGirD8XHg0/g4VAGXLfX1jtDv3leuLB/ngIOI4q2lSBsp8TbF/OFYLMLs
qLX3BP2SXAcbOhycqQhUhy7Yj8B78JKZ91S5pfuh0YMpaCfyLpA8WLtQxyOSmo0Mn/6naoniBrX0
1yr+lOlyDsu41mgYYFwRbYjBWWjvCPwlVmIIppCR4rhE4j+n4O2o7/X98zWpZjwduH+L5NmYkEb4
kXKclNE8C6Z2tdDyJrePSdzv3CwNTQZHMqdENhOm8yOMeZcoQYIF6isZUOB5Pu3Eczrc9M2EiTo7
5x6KbUt4EndMgHmYRfFWmS4n1BaFqy5A08P80nA1/2lEOqtWk5bum4gPJIE2OzOu1jec+37uZVJr
vhEIvFxB4UJq1KMD8xcanf3iHlL/eioJ4lcnkOM+oipI7QcchL82v4/30bAOf1GxeYbqO3nkBjHA
OHj3FtKgYvhCBrYK13kcQXhViLQcBTWlmqwCTwX3BTzeod6rQ7IJ9V6q8L/zuvY598Q2tLj71J9j
es+4aXPTD7IOtOcJJ23tAY4nVu1BMBjK4o8bdsGqNGveqyuR9Jpf6BSgM8C+VFceiowA5wExlvFW
IWX6EiAsUkZiu59K+JRQ5O8jOXHl0PG4UulQe3m0sLsCf0rcWErKVwN8kaoa6cj2CLlI6Boo9riU
gwFIKNreirWreRXz+EbJFZ6WyMd6pIUUX1JaiAViazwAhBdE9jxiXM41uDaj8XdDNyrWxgDvpgun
VHwDZIIPSHSSlMmAl2t8jZILgPb6U+S/RWTYsDrdroJ4c3XxjqGqBHWW3XfoE+reIByGp17gc2ne
eAmN1Byw+OBw0wYVdTEZywRYOBkyV1CBYxVSsJ1fejbpejnfzYNjc1stRSEBFSSpR7fgwPjZ4Oie
5PRpyW6hlqRw2XnS6D4bIJTD84y8XZPdv4Upg9OvaRhY3pVgZ/9Bs8MLOunmxbW+9KVlSgS/VEWS
xsAXSmY+i5EL3kfOOVewjzEZH43SW4JtlOE9GpeSov6NS22MpJL1vpKlsGACtRCsFtNowhFoYFgX
27AN2YhipdYiiEHuEYH/uu1o6y2dsa0r237bVwaZ7nV9OyV7a1UhR8EU2AGSk1ARAU2NXdSRAmpX
ry9pnF0VeH8EfLgQr8f+yEO9KxQe5qGYUemHBp2jrsly4/QRej2L3Cfd2aZkN/3HoHBxcN8I1G0y
FVVLbgpI2nf/ZbTwlTocbiXrPYQPddrCgqzTZBCaW66mO07NmcNbDMyf+3wTyzytSXlH7YhRru2V
pCLfJKv1N1DyBQagPW0CLcyk9s3bDKWjLSwst0khcdc1mQhb8I5JlJR04os6lxA9DQayBdzohqKY
Z8DJsHiluvK/fXWo8w7tBkMG2mPorjMdyz3rnV4BiQMrnsLWNrOv9gJh9ErCnpOxp4qRsWZdtvd7
fE4fI8+/jVZXUZcAShB1B8rfzM3Il+4axg5cmd0Shfz/W1f14W5muAQqdvs/m+9dU/1UgArLvgqg
oCPRQ5/CwrsKu+CiiRsTzpKHE9m+Jp8yfRZEUYRp76VgDz7RKHgxXmYLCKJvKs9GkZbd1dG57U4w
GuQQXcnO5qiC50hHPRM8DgGw+DLwGQI1pMLhNRpEZ+V1yRrSrhzdIw/jOQEQHZOtS9fZ2bq3UaTr
Be3E91RJc/vEbpRRswb0BO0hK3gG8e2Hhttg98fUEutD2Lv5JArkrAut5z6SNgfB4ipaqxvDeZNc
aHuWa52iTAr4TfHcnBy6E2U0FthbOWluLxVNaeFrpw0Elg8gIwPa8sqfWGgkzl6YcafLRgS5OnCn
YJXns5Hdcj6pBuV7AdefZ3MN0EtRjOErDvBzOvC9amtLdhc95PmjSYt/z7d5xZKRv5Ch/yrli3VO
jWULYm9kwVJ/yqNHfN61LvK2hC7gK9DmFs2XNoqoMN+lAGK3+ZmjnzCtTeBZ/yR1Q8qYgSd+PfSO
5OGDSkcJteXfWd2ngfnl30eLiEHvfczl6GKif3AbAW0MrfMW0Kf7m0IyVuTFhdiU38ux+0XKuV8e
Gaj9cgvKUF8SRR1x5cjiKjtyYP7DoPHArGnl2F1tz+mlGB66q3j/hhErZQObQtKy/s5SXNe22M9r
YCRiaNhQJeXo9vbGB3BtTgind4C+t3mih/Ok9UB8sZxgk6aciWiIKttrPHN4fY5cNFyhmZA4gYV9
rGlp8mTK5MqaIBp6LhHR36rXTHdZxEC/F3BhWt/taqPuy1DkzGPjErtZHVvv6qjsijmNfNtTm9ng
hahJ98l3u4yGxxdW+DbESDaL5WE5l4l3uxgrXBJrFmGSJxwe7wHUn8hrmCPUSnVhZlNLSBfFzWA3
4axoxYWzpj1drIWSKQmCtHVfUYEMR98jWmBDEK+xG6SVj/prvc99EFi6tZQNrlRgmPPnSrANZHIO
c6NpG2GO/vsScpPhvkHRHRoY7pKglEMsEuqrCYy4DCz7ZaJXfZB8p0PI5GJ3re2R6tfTT0S/n85N
5bRFfRsrUnZHSnHjqOactkQ4h0NcuvotR26i7aCkYyBCoq/4NQeqdPO2sD06tX7YHJ1/Ouqb2nB8
DQMXSHVFXF9B4YDVInR0Y+XxWtoIENfnjVXr4lGQ0Idw5rCJgvTgS8YF+926lWs101LSlHZa2rJG
Wqq9b0c2HZ75uUurD7m7jZk7tZnQefSLMlryZPqiIBNeZDzKfc7xami0EwoWlSzXYzw8eZa4Mb0J
Fajrm/bXQsKjaoo48/O2EcsZj4OYD/HO9ufrSjtL1pIJhLfnEJZSqcqPDD1xOhOY+WJ2yphQQp82
Plk8hd0uqxJiDkfwdoqqfw4arwFkcDngkAmVjWTBKeFeH8smqSnGiTlOMNGi9xQeUNX45kSQ3gVn
0di5OV0PkO6eZ+HA1x2kYKvP0goK2gbRfdvhD/RH8BFmc//PqFevDnzfUpbMAeVo9U1v6NbZgK3D
Zke4xRhmaELuZCmLpgbNaAx1AgOH4EfEq4YKAj3aPSyfg5QTd+o9fwxj+BRqc/l1XDjC5xCFgMkI
Xplh93Wcr8fdG4HXvauQ18QBjO1BYaKf1UtRKiRLE4sU1cWA4niGkt/jW26MfztTtjVAM1b0a/+A
Of9IgRYTI161S6NEUMHImy8gDKV39QaY94kQXlMoONi7YuscSefvbAyT3MMEslRruBUTO1X0qTSx
kXYsOw0VVb+8dmafCIN9X1hcMyYuziYygSLWy0dF9v7lsDvIJjfADkTjOF60cz3oaQdRwc26W7f/
atQ1qWNDkpcJY5GZtpBug6V3G6B5jdT2FS0ILAvPuxDqBreOPtfufrXn2CchkTOLYPO5sHAHewej
Br6lkrUine7v1LzHOHXJKISi1aac2FZzBmBYo+U9Z5iIvyys5Dbh1jxHED+dM+036uiKDmoCFY2q
63tlnDsYQvYqQUDX6GUnqK3EVg2CRafHy98+/yOC+5yb+eaqcD9ZhfY+dnpiHJ74v8Y1X5dsaGjb
9BaKgC4TRjLdte81QKMXSUVeSK1A8hz9SX3EOf0JSdFuDbTcAipD+H/TbCMiUfRk3YU1yv6vzADI
yLJ6R8yZ3i6F4CppXoU4+6kAleakWz+CzImtSCAcAaFd/uLqkknUyCTr40tRrSbfOHBSI4btWfZ7
FSOsgZ3po8gGZ0HRC3gnwnZvNq7Csi40S4G/+naT62fIe+dTRQ/sDjj2+/b31sCsqY+Ax4H81GRU
8VoEnGsYN5/KsIFWnhrOvJuQGQyxC1t0PVAgGlKcmSo557dGBXaFxZBAyid1ObOUKJb+ac/ZxnK3
ezUlnqm7TuZzUPZRDyYiaNFvljWlURdP2IJwd40WX7JDqEqf8Q7QgKjNupBSYUQptiyJ/N4i3dyV
9/+Kjyph6bOfxwFELu/RTy562geyrMQ7Cp868arizFa8yLK5SuqFKCo57jI6io5D//fuwM0qXir3
3n6ePgo7UbaEtUk+mVaYfw8H68O9VMAd+yO6PKCZ5WlAywzMu3yNku9PzjVOkS+Xut3U5s6NOY86
eValWi6/QhAYM5GfsTc9v6cvdzF0d9H43R4SjZ6c3tHlWkX3xpRXN29RuxhWw4XI/9uDvmEfetci
kxFiWeLlW8ywVGvCS8OxmzAzmwc/DQOCvnXPMJLFAz3Uho1fJhP1GwQ4ySYEb7uxFACZKdv+i6bO
I//i9h81WRIiBlaIcUO5AuhUImC0uHSxkTUbOlK3hBeJM0V7Jr4cZ/qIdh4NAYwVogIj7RVGmvsW
FXeL6AEZzJSzZFhByTgKtFhKo6eV/6q5jQUpiGWp78Wr8rtMVqXVRFWMM4r+oqYa+/mJhmwwxDL8
of3TOx+UpGBNyurcjUFhJh6U5XSaynAI0LReU9pPAjW2u0/SuB6n0xGfJhRBERI7UEmyW9+w1UlF
Uxs4JS8AY1mZij0bPHFLKV3VCvmrIBTNhlotE6y4RBMNtJQhF2M2jJwq2dwWcEh2+jv0xhXS0c/2
v6TZvsYMqKAqYI+S0w+sIeNNwxTS2giHbjXJuUzXX813kq2i5l0Zb2GBkmhOFHhA+ZBfDA5kekQh
/okHpQgC8O/zZPcByQMS/OlFjUXWODP2bDZFM9bZnsxKAYDEcA034kxJ3qcn5HaZz9T0ZQCbIiz9
N2Bx0rvMtenq4yOmFnyqqxk1aNMkAkUdz+G+1cicmfc6YO84mZa4qdCtdZz5TgmbBtg1DJY2W0b8
bDVNPUwl2zAoRUwUPDHvFSwUfFjjHgS02PIovyVTf1Gq14stbLIgdY6MbELdNyiXtX9sEBemsdhU
rhl+q+c9qNwBXFZjRKK+qr0iFalOG54cFNBFYKLlv4y8wXWtJP9YziFXtQB0cr4G8JUabt5c6Gk3
AFPtcj77AuLU0oUnmRJ4AgQUghKSy0L2TIP5J9u8ntrEfxsbCajUjd2OQmKXS+5wlLzr641Z6B7R
7QQ2t+ooTZ9C/iX/xJAuiPuMDSNn4hDzBfKuBuTDb+Z+GPdrjib5aIrZFv0Q/kMDhZja04nRKlfz
yYfUmVKXPn99UePv62+/DvR0YbaBna7ll3jN7n8Z9zFAkJNvGq6kfTp/KWp7g1HbCXDqsYYjz3zU
cG3V8CiEcea24yXpwGx4TIkm6RJFpmbspyb7rwt6b011b9otCmoETlNb875YMt7bC1cWSX31GjmZ
R52lBzuRGfl5QNypSDl36cwmjLsAJk2S41EuADfMfTTp6a1FhZVl0UKxYw4yDOC8cOyrK/gREYF+
ZSuG36j6G6vpecA5woDDhSw7ATkey/hz7FFENSZZEPTBvNls5rNELwQbQeaCexCs8PPbq3vcoKe6
arBRR41X0qdi2Xe/pd/3ZHCTCXYCk08fbyAc4oU/EoWq7pTcPjpd5djdNnzHvh8k2gsY0KBr6L1K
yy9NYPQfh3M/xDTydK+SO3++l1wcRi2rjMgCjMsPps/X1lcLyX4djmjRY7TeWRF8tcfjLfLsGjV2
o5B04yW7Qro07R3CVa0rApXr8iqDJ0y/hinSKaNZgNDOXwFzltPznFCicr7Wa+Uso7Dyf3639bm3
86UN9fZ5bZ7OD7WbOdyzA3kZY7RejRFAzkFTPRao3yPgV0vGmTYZnsIGg6CDTtHp6WSeqAC8I5zi
1cp9LkpRIPi+g5JmTNe7DKO9OoMZr1LlbhPKdoG6uF+3F6/elVkNyEtibjRhJswNNzO/PoAZJssO
T+oTPtaoeR7OFP9SW9CdT1liaRT4aP932Qhafvi6NZrofyC8szG/KiJIk+qem6ttfZjNnfLs3sud
8yWPTtIDwtLn8zHnOTCa8f8rj24W77SuMgPpAX/TnTLpYRe4n2IrTZiu0wGyNF4GZu0v3ny7k4Pu
f90yIIJlrWaWR9kLpaXH0g6n4UAM8A52nSO/Gvq2ck/+wlic2HprcR685K6KktbC3aUagdHl/rje
dpB+0Rqct1EtrDpsF+M9DJFjLd25iY1yvdThXddeo2QGjtw3hzLMJsY983fn2Ih0W7VlO+zhe8wM
mMI1lFff2RqO7owuZicMoRJJGcHQRTNhKdS7k2bHcpXkeRLQO+b8lOp2jMiqTe8xC1R1xBybaz5G
8zdurF14y4rXOBhl/A23exRn83c6/eeSMliTMUWeGHu2NFt84H+eUbdbdGjI8NIP762vnVEH0MkS
mhkV//7/l2Yai3ZkZ2IXnaeqNsTy9wHGwPS0y21wV6qmbRJ/3c6JmQXQw8VIznfrFOJnslEk5b1M
0qDFaVah8C/g6hbLUi5cAzUs6TdumkxuUcuyG0/L8wbeqjBdLEciKDI64MRo8gPV1+znSJ6gAGrU
Gljnu6vYVc1ClKB+EMQiBnSVtkdl1vJdX9BTSq1k5JEP7nRvdNFKY3lZYmWI5myq3IDkubwnGSM6
W4677k5uobwC2UDMT+RN9XAEkjPUOaJGujFfYAReLMdwgIgXPep3deRuuWONHjJxqWQxtHCREq7S
4FvU08wgvSFfzrhMX/gK7TuZ6fOdFdWZr3+9JA4qPB0jTjViBYshXpgEGhh59O+W4b8pLDHzRu/G
sczFPQAmuQzNbGhS562Boozk4/FMCmddB4WxfIoZdZ8FO2ScjPTNIK36/gmjYnz6MeQxVw8R1NbD
lKev/fD8OihirzyZihw+ToQRd3Oita8D/xzWqXto9v+1QMKYWaMna6BEhDyZVNGokwHQlJ5siCPR
JYKjREXOI5199YCSNA3q6G6Ea7FwO0SbBrrl3/MJ/Cl8Pg0kaEnaCrMOY5jne6txabVolU3kcGld
QR1VdrusaYIGtbD0yKCBjZE27vjmpIIS0wazh0HZy2oivyXrLgnQ9kuf4QmSD06Ld/LXsaF489km
J4AS62w5iRdgHVvUE+bT1w9iCnvfBO5Pu7UtESSPklrR3dL6F/z6yXQS59MzqVEt0N9cCijsv7bd
in9Mz8JzaQgqJAfIlsHO3khJEn1wvLQfZQW553p173GMh0KLDLylP2J9tMhhepgWlN1WAYWSC+np
KM8r4ScHrCfuutI8hazXmOSjd80Kf27OTLyEmWwm1H2MA45eevmuEpAGVxw/LSsssXiornAP8GVI
n59ZesZrqaQ+KlgZc+u/rsob2Dsm9+iJkkUfM+fylNVUVVw2hOOiWTBAeTebO+sy30I3Buwvn8Q9
4bNUVFc4KLEfmowl9V0c3cMRSnnyPQQGv3AcWu2+JI4Q7YGP86X0RTPQVEthQ5NWd1TzGPauBeBw
gDmRfSMLVpfza/Xfd/TK1/LDERl3VWqhiHq6z6y4RK82AyaXlcycrbzH0maSAftg6grZbbfqjLsW
WRZyhi3Tk0YuVkQsHBtPWqBjVvJOVpYPJ4Sbf7IYlraJbxyatz1UBu+9FXOtoRuqUbOJ9EfmMrHz
ib11yjrrDkRcdYpvMEwBCfEZDvT8GSyeksgnAIa0iCXphb50HOB4mXuGrrSIZSzIfsBVokING9ej
zEKZ8e2JOx/59sTZ6XqFuBUCiFP1y0R92HT6DmSwd8L1EOjNPzzIs3kmP6pMisvQwTHcLeCsVoFf
xlFpvBqB57bF43NMyzf2WTdF3Q5BsFx+A+I6xMogDBCU9x6tKo1A7Pc0VB88GW6awe4NBQN09Hd8
ViYQF4uzHrc2YnyV0RQ6z3/2I+rDh5xkVc/O3WAdJzkYGCwvJd5F4kQcKQyT0Hrw8nBeFH/Fp5Yv
xAQtT8kX5pSMGMuEvnr1gKMSoehzfQpNNst0/i/r8Iw/VwNzBy+BN9GOxIJyXeVE387wZXa6Vfv6
7FPVpPKexeaUN//tgCrNl67EbI8u2eauUx0XkGpZT5szIq8mAG2WtxOA8GtyVnCRH+35MbFVHP0c
dxjyywlwCYkoDnpf+dGOon426vRIo1WPPlY9tpsZIaWeWLuL266HMnnuAEO+6yNt8jdi+Gr74I7E
pkUawtk6jxqtLhSRqzTEPCES/HHqJaaEPl2ZyN1KwUWNCeRTCgEVMG02lmyJwBx/SK+GW2jkCq7o
nJt8w9xAe1U+/kipcZlNRvWNHknw9IxuTUl26W7Qng0SrLITFQXGIWgvSUrxQ4Ql/vJfgfL7URkJ
bBRQS4hlSwOPlV4SlNaMluGNeG4f0QUpVR/FUhIZVrEyYiALGj8MPygEYKI3KX8o9os62r19HG65
+zlQqyMpk7erbIHfK13nJbm/KHzzjxL9qy0tERxmpcjcyeu5ztfND7awVby7nuoQYYNf5NxXlwqM
ZVl27nMxTZL71dgNSE1bCDMMz8ydkZIqsjIPBOniMZGiJdL7xkR9nS0tyRSLPSh5wMx5XzhuYOG9
ebxNYMLjPEheEmte8ziiWX6SeNWh2ysk0USTgfrm1jpyrrhWUTLqGHKgLWL1KQgGU6xkHFhbaNO/
/lPxz6mZhPncz4qETVaCWoRzY5kq8rJkCo8IzGQig+NVJCpE62WXIVAdHq9YN06OdAtX6UlvEuPJ
viqY3SwoZC/HjNHg1eqRn+xwwRs503zij7yFL9OGRXParzWQ8Q3+5ZwRTyWLQNwj+sgOCvQno5Ra
K0RzSfaNH/7Nh851ZS74Ixz6g6iBkO2hXqQB+gZ7pe56H776x7IG7Yfn3BmyB4qvh+SvJx7S4j/O
ZNbk92elYYQXv/SpIiXc0AlX+7sLIRM26DdN99rebxQuuCaJ4Z1Dy5MVHdjLxQSlceCImGCZKrlP
c06bbfN9CAX9QWWLBVH9AwRxUlYXgw7/YZLLivaS7a2FQlQqgo9cWRFTBBtPgyBl2uV104r5/U7b
/QIbMsVJFKO+fD2OE7EiCtmXdqmlY3Pxk791SGjVY3QiH+5rHNPIzGKPb8hVSeFQIcY0oBmYbCh6
mNSkPFv8mqor+Z0no+52PyzofUna1lC0SDaRs0b0QZcWWY/5AcoDGPFpnhpoO4YoD2TziNIP6/Fu
ADgy38UmQFjGkxgyIFFX5NZ1JKQVWlF2C0QbEI8+Eq6th+dWThDSMQbzQ22TcvKl5hAUlwMd7R40
8wtkOPZhM+LN2HR0sHxy9lReNXgJOFfaDFEpPcDTCIagCfWYWKg2yLsH0RolmI4jKY/IsMligdJG
euJURRc9GHV/f2inTKc78VhHePobKAtodINraOja7hqSU6loeDClHY0+/zSYlXkhJM9rI3Q0STY7
kCPVO30SbyGquFkchY0hqCwCkC/oJNfiuxmYORL3IUSfxpFygBBzOEyLTUJvPzhQEitKEZSHu6B/
rHbklPf88gM62emX2qIgBVI0slZM3TB9ZCGHMndtaMKhWXLc5AIriFkXC/qi/Z2YxfmLRhohYcFm
atm05DYGNvNPI88J0gBCF3jQN/AgPEoc5h0B43+BnLIDldfV69qkv1M13NZywx/MJu9a6H/+7PxR
t+DSUwwsYdtvlUIrfmF13d7zyp4uOXccX7HpRam5c2d3hHBfKGNkluu8BETxXu8gbsi/j6X5xiw2
OdpysO7UGcvFc507IJ7p87nrz+n5bNc2WChTKoYEY2WHAIhgvoSrEZ9rERmKv25dgdlyqaUkEITF
C35uZHanSe+oA/KgJTnbDmcwRKvEKymgUIOuMsmx3LEd+0lzlX/G7F9cpr6ovuJYNm04OiNOfxbJ
lfaHZa9rpqFFDS+tAXY91V4Tsacu8XFe3NgIw23Xr7CR1dFaxQpcHqMylIJz8pHdzbXQaG4VhyP6
M/tHPg7CPLvcZ7Fy4c5giU8sQbBBcFSLimj/jvAz4rNGbwF5l1S1pGJq6Yhx1rAjaLTA6hHjzbLx
uzS0zm8UaYNZZ4rd4N6lVeA14jHT5Pwo8ejePNYU4gfOF3las5wqHlKunR7/d30vkJTtZYSk6rOu
Bqs1eYzFxMaQq44wqQYdh72JELnW/Y1a4yqE2SEHdF66tLan3Kao95N9vHG/sRmHZ1ehuZWT96+p
xXrl4smFgv0YYQK5EZF7uns9pKGkerWx3de6q/iLghijEn2T5ZzANhmKpyoZX6ESk5HNyiJNVFgx
rAHLO128ubqeBWdP9z+7xZNCVJvC7dV4P6/olQWlSDzUWNE0eUZEvycPHlKlSj++ylRdPH7sAR0D
0QqyEQ/7r2YQMjLfEXg4Sbe8fnD+l0JVPuUjqHduseijWLLOaBMLGttio79HaMo44e1/78jDUPd1
uc0oizNjcO6WHImOJr0OKERomrR5X8npU8SiMmynqSTipW655NyLw7w5jx8bih9Vf3suaf2GlTWL
dLJqLT8K5bqXwMTsA0841OICWroSSJAk2lxVVAe757cwZpZxa3TYAH3vJ7/OOnhdJp1oYKjZ2ij9
Qi9D+A8AQ/TDisdEEijdjkvpH66G9fyi7e/58YfNtgIzSUSfHjZIJZiGTi34ASE/DFtRCNQ24q2H
BQULd+wnQrgnI0cpZvo1//AtY4VF9XljhBObCMc39hqQOdDkUxCI2XnqB+4LsQDh0GYYNd+OD2J6
n6fHaRgz2r10/C1o/kVT4LPb+kfV/FRHc/5tED5TkQq7fqQgpErm/OuRRSmZLyxDSZtMzQWVHvh2
jbqIFo+QpJmL09ct8AFPzcxnS+T+tebZQI3DXLiUC5BBq+b5x9hEKwIcLbMMK0XcV0OHTWwhJXhX
nehVi6rCvOTtN3Flgg5BLasImBhr+9yRMk4PPIrZpaKRhgIedaNbL0Sf/SGhLu3Tr+QJH2K3UNzB
UinzdcoOEnQ9bb2LQn4eWZpH2xSNndsG708mubcw1JVHOq2Qay3oYct4URgW3XKMKEIreA+jmANY
CsRLPR4hfK+n4FGsIoOCzjrHKDXIgrVek8+UPdTAOP2CSLFIw7cB+MvBVGz8IN/6xOwAffP55cUO
oYT83iaZNmAsTld30NwVu9XUEVnJerSMHHozJINui1iDQ46H8xYTpXHNl1UA2jwFWic05QjQI4hb
4thG1IZADgjquQaAbUG7/lw7ruiZrKko8Cy7RLNEoI7X5erma4TkS2fLvHvXBwLXUmbbhuVnaQGo
wW3bmPgrp8Xk7XyWARUsCyZFEdCyAfKpzxOaPSn7GgXBj6o/PEgU0VcAmuUAQqt8NHtfkYAdofae
3Mswxu2SP9QI5wVULtRry3FX+KMvLGLHO9J0b1ClZtnsTvOMKLXEPic8VoukkWWNDA46aZjbAkU8
nd9vFu+RmoH/F5ij6UukHVzNEF2xqp9u71iFp0rPdf8ArRwF3RaYfsGNcMyEDcAHQAxLzFHUbYPe
oWANmxkzWk9GWeWzU4aLCrO74qX5ju5ZKPZ81VEmJMwzBpD2Ts7ESweN8bdSXvLh+6+MnliDqMH2
Jh8qpRWuj6f2zg1Xb5aOJx2FQ6a9dWJQPfDKjvueS+oljoXUQxgyqrYczr8mR0qf4FXSEjSd6hQY
38Pi8wrp/rRqaQ54erHg437oZAgIyLZSBPDN5sNlJQTm7eZO/ntEL5w2E2MZNvLvt3nzHYRnCami
1jZzW8BqrYj1vbIexWp+i1MtB15WXR2ddj7A5E/l+iNUsZ9Vn7l3BY6m0EB2BMeTqaClC8iWRV74
uijD7IMPlxZ/qmo8ilybs3URMdxVU+sxN+810COr0ju5HqORafNUTMHyjjbO4YKwd40ORvubzwuv
zcR5/Ls5zhlUGrIdG4Y946+DB2+e5Q3gUyo8ZqZ4Up+QQ6HUndseGBwt3TDct1yrEDv4uDabVNTQ
Y0zRNph3KgLbnJGLAUQN2OXKCfKGsLE/S1Rr7TzpvIT71mjCG6VT8mDy4V3rQznEXhKbni0nAz5X
Ve0h4BYHuc0QNhc7TK68I9ren1Lng3UuppTcb9g/FRDcaf88crgOb7vJZ1goLUxs0EepB7UOik0e
ZWl4NNlooYfc/Pn78xvGTR5YonbGIPvDpPNNWD7q9PvJ+n2HKY1S7ucuVA4Nwn7rrO2KiMbZ5Z0p
regA/LpZkvCp4bbEB9h9rJurcEmk31QckG4KiTda+zHnSRO5GrBNFdbPhpaFcyrJnaHWuT0fKiB7
oH2F+l5x72Ez6rlMv9bfyfMpQqDgo8AGXbg4euKz/AG3tylrJioIQMKh1cyaeiXl5DyrN85XY74z
VacZCdTKfPP8oBa2GllJZVax31hFuuTLPOwSAyH5uvMTMjgCb3wD2lWuImp4dTl7tDvymLA7Pvni
5NPVhBiVMmCruGDnJyIAlXDlDaOaLI8Mgsbrb1xt/eSHrZuRxv/BTwuxRpxf4jaI/sayKKAFu0la
bpKqNRFtBRO0leqbD/MyYIwgLv04YwfhijNoz3Qeg7hsKHyU2dvqKhHwGhKLZhSC/xcNMvBUyQQ+
Rgsq0r4MtBlYGAHaASqG5ko7jGulAFWdXXo7xc+8lQx7tk/YgSl7ipNEWkOnAzah1Sm2CEXwlw+g
hUO7WiZ3SIzrkG9E9TF1E8r7HeHTR3gxs6BeurD9lD1QxdW1VdX/JxwhMY8Ls8lEoiVGPpB/9dAa
7Gek88vXXdwfAO03xWhBoFAlbvWlMrbzxM48M5VbDNqGfUUNB+RrueE47JShUPcNqb86TcIcIhCF
CZYgDA33qdgE+MfnBB+eKYj/E/i+M3bjAFm4u8TRUVmfqCAATaQE2iuHPEB5fV+912iZrAiDX79A
2JKtUd7ITCs10DW+8bMH+730DulcydaksWunsDMn7AFL70ZO1CvHf0yAPOxFaSC+eh24SQR6jzgz
+MJPa41FwVk6DT6wjzyCv79PEbnzUfwo8WskWg+BJCDK3dYtJUpP0vWl1llgZdmZNjs26TvoBXZe
MHGEpLWE2fzZMvbNGdNRF5zkKh03gViVbcms4AU+3+C0KToiop9j3eaf0TrvwjV4oVcb0y5BaJmV
Ein9w1CdUIhycqPOOwDwvSc/tQP0jm8vPcojJaBFDRosh55KpJNU4rRGdNY1rRc9DBhNOQGNVM7I
vHgOOY3yBzVynKKmJuEq+Qiiuc8kh0z8WvKg/a0+U/xPrmYwxvrWOpIj9XqsYu8XQ2uKEKU9zFmx
oFwcMmx7G3OffFusDVpt/MAWM7xguLR+KNSgk3eFYAIVXyNTxR8PjdBQU2SMy/ZJbKpFPL+U3PVH
Kxct2b5C11mzB/gSvpLUOVRAHtwz+jOoRv/8YBe1YXNWbLotNUzovyUnL5w97aKwQzhLLFjZyNEl
PAhXIvToxvr/rxHckG9uR+sD9NCN6BD3fy5kzF9A8Rl1NvUw+oPTu9Afu+S9Annk5G6hElK98WQo
Kz4EFsl56g+PghJYM2hhDaXxdWQ0uBQ8hiQ4xUS9BEPZoNyazQ5HCbt53/L6NPVXD4dVAtUV5tAy
0Av4nCcxQn7hrvcF+TgDrE0b1ylGpdzdCKBdCm33OhBDK5+HPdWsVhPUJ8PVsMNrFg6hnzIGuDWR
xlf5X1zyq500/dWJxJggrJbCWje0KzIal5kfcnGoIZiyNC0/iwzPdCe1cVi7Vy6fMDcqYWyLeWMg
pwmvASIanxIcno9NuRGK4Agg4ooQePElkp2lFrk+rsLitKkRkGZDwucarIH777P0SGcrbH/HTmdE
kC4GSJRns2c9ymwpT0f2+YcCBNyfThZXsVYPZwfqdos3nyhsZZYsp/tYKh6CoHYOVftCQGt2A/o8
i1U/lW7L6rL/J07hOGsx0XHzwd2/38PXKSMs9ucQ0GdQiZwQVDVd+1Qr53I6LYBmkrQFhegdM80F
4Gtal6jrJ3EPyYViZ2z5e5YAxd+FPraCuMqJNCmYSg9zaifu5XZ1NzDog3SZnklQsSOD6cMRaCee
CLZNTJ8bKEHp3DYXMYw69rnDzO5OqwV+9cLizu4OH8cx/LOnqrrM+Q4spNXBQStzAiPbWfVe7qbj
5TjIflqXg6Z6bgh0bHG9190kQFRJ/srXOnnbFjDhIAVja0k4iBwrKW8eEX3j6FBWFqy1TLp2Ivui
hJClXUTYFuLgcXnqS77OwW0f5AoIdwrolXDOiB2TUrhJ5+Ib0bz1B3mVIH6OvTl/4z5svzdFOz/Y
Ac9jgpqy+A1kvGmi8qyluWgisvyZehOV3FbUde4OijfHYoqK2Xt6xQ/eNFOVfdYx392pW4Rv8+XY
r6YSLSAcz4wtuuQc3kgFc573wTp/JgyY8uAqP/pWLhdQnZ5XZ+de2nCTazEAOzLCHEnM8+1l23Ie
RClv7eCRCamTWfFfK0j8o88/aZBJzk0pnxnzegGqY3Cf5IFXW2TqLvmDBJE1zuv241OyFqZDe5r1
G8Wg0Q8W2QQrStL9bBTkOSDNsP/BFpAvXCG/ZKKV8ReyE+iTDa9jUn8TDYRDbjPKfyrGt9uVPO90
QviI33Qp+8gepf6IsBGMsn3ub/M8czjdnP55AJIxfmt9PGfjvhXkROVuL6fiatytNQJUx/uNTU28
kVUiebQPkOEwkn2LSoRsRIXuO5Ik4KaG288YV54F5CG9OLFD8PKNeWyOpya7/slesoGLDXFoB4DK
OgHxYJartM4iR9op54MyhDNCQyTU7AKGjuuEsswNpy1XGZJowwx6YKuShFduj/ijqygh2YJ4Dsn7
RlpQSodpQfDPLoGjrURv8GIa3JIkGwczU8U60WLnifRlbGoSdVJO7uqLg2X/HwxXxCyvwvYukaMJ
InPdCsZDRyEB1f9XAEwtnEhe8dZGQuOYDek1HweBr9BEImyOK8+ceApRDR6gyE/UyQum/gDonhBI
d1aaodzZ8Zjoi7Y5IQ9xpkBs/7TIJh/uZvgEwtP234G+ldcE0cVMYtxNIDTVaEoza9TmuROiAEh2
H65j+4plLpAGVB7xrqRhibRX11dfRXFZ3prfgB8jayIAyU2MC46KBTygFo3hXa5AbQ9GDEUhJnKS
qdyTiLuzFbPfX3hYbaA90Nft4IhKJgf2XqkSL6ySDBkkCZMwC1h0YCpEDHesmRQ0EpIUniahozhH
mrj6OpVAiulKpEqB6aIArSH/TY+CtJongleNfkkbyVBucWVjKvV8vKqX+g/fvt2fnLggM9bcocZ/
UzhX0XNK0Byh6/+P/jJxYxeuuehDqh8rA6Vdi2wXLZ6z9YoOENAN6jCQkodFZLmRI+NMqg5hWfyl
vclOlILg8kOjTdlgS8IQg5U+hgEDpHjsFpP45NR/pdAH9DXA0/9nmmuhmPTqOdEL0iecJBvATP7s
w6EiHBaHP5Jr7vhlR8BCedbbuuKvb/Jq84tHAyhGly7P9uBQWhBoXW4sufoMjpv3EOu5hMN7d2hC
j4PhR0uowk1x5Sk2OFp23skX0+wDp+jmcExBzYuGZynRsfLGrqiSADOMTKYfcDKoK1AcRNF03LXJ
L1I2OyaRFNgbWkjrkYhEObAV6VyM2N+Oeq8jdHHPsnngrFdZCEF05XY+P/LeqDo3bNg8IW4bO3sc
EScoqgeNAYfMj9SS8ZhV4KnEkOO2xDIBiVF4RvQPZh4hjSteE/Mv+ypvnqpwcudzYqMkNqUCce80
ilfkEzUsgbyOcv5LCnV4mRisAQtERxeMGyO0OjY37lzsIW0yj8cHqGI86jczABouiqrx8SxHV71k
dWy4okb9zMj+dilgjGB+1sNZ6hoUz1i7sBO8uVLNdYCYiUECfRquuKk3xBqAWE0FCHAoAd7VcjQ6
zoHd2TyA3mH1SqLiVTR69LzB+GjJ9oCOIspnMzAjuyuEw1U6CSeXftuoL1d619kC3F4f9x6LZVo6
hbbo26TkgjZ3YMyHC76mVXLHTraNx5ube2GlbXLA4ws8LsGWqaYrPpzNUqM3Hqz5QUr8ucTa2AmW
1j9J8Zo0LZeMud28ggE4cJ4AjoBcbcP3HvOU0sO0h2D5xyrKtSF8PQpoCLOoStYzGgWnWm6cNoM2
ae4vtL4buP5OzF1UDDKRCwhsOWI4Mo44FQHf76Trne7guBeG44hsDLTTt7gQ03Tfw/41OH/ByCww
2nhomSO6teLrH6ax3pxNRol7BQ03FFuizy4I/b6HdXsursKQAAsIplrsvDCd3L0lgHejVY3tYILb
tAGEOvM3oYHGPNL1P1Oki4GKDQAp057IF2i1HMOKyUQqPCdkyDinhEFZ5FGcbd7/lC8Vo0SdiWLd
F3sQZoli0YjWNCguptsYVuhznXDGjmYUpfxPDej+WpxtpCGXQB38y70wacSuzDujaNB9m5621fOg
vfMJni7xQWB1n6xZGUPK/djZQXGFaZXv/V8ZmS+XlqcdMmGucsovfvOFPGOJ/5z2dBo0VN9h0xJK
OJxqPfm+W19f/BMMh1+quA24UdvuS8mPR6RPnU5VkCxq3mB7lQsM8iGKFO+UEcRD4owl+vJffELL
OntiXnFTZ79qrOXjauFZlJplcY7ntVDgsO2da7iePjG9hAXGwisUs+64Kg1LrQ47Q2dylGgaHQzy
PrGs6TP55KzhPsOrwax5GSHw7p/FEbGQE56xByt4+xnOxL/A+xYzwCjYwDAmHarZ3+/H+73TWITP
xxUcO1+ey9RlVoc0w9tJ7mKta5YAw83moI6CIvSdUahR+gF3FINw0SOZoV0BovHYKTwQ1/W2coQc
/QqIgUT5ZmqELKJHEBIvtmjpuP5x5BU9Ehu0dzEGOLsv2CoV52V+FEc7a0fRI84jA7S2THZW6CXH
wWTvi/DZ7zvANbmL3xnUywtMuSi2YCcQnD5haSfTv+x8XAyElrm1vP5Y4xsefs+d6E9HPVWPVMr3
55titbic+obAk8maz40e6KuZUQnEZPBo2z+vEYzc02YFGH9/gc0Yn4yhWcRyJQN1DsNVCV9K3a+b
lZqkQe/HQ2yprB5KOsReQ4iYq8a2GyALxAQ3lCYC0/Sk0lxso+wqHQnaBSEfD+3A5Csq4z6PY2sX
/FAoWaIoui+UVBOut5DZ2oZyhembVrhqwqB46p7U0ILE15uzv0l0ugrDNp7pv+DQ4F8Q2B0dHn+h
i4NN4ml0lJcwfXERd++12nuYQbYux2A0vuxEIQGaDA3D4tBJAkAzSNLLzRqZLSsp0vsaxoFZkRDJ
10kYwXeTmyjZwtoBgo08XBHBWYqBOSW/K3gYEwteG5Ul/aTymKFsvJ+CUITV9yntKS2/RBFomAnZ
4Ye6+np6SZKn+hlFJwXdRp9OpVis5LZbREBTpn/gFq3Lxjr2sEW29SghmiLTOByB491okDFFlQGQ
6x8vMKv7p90AUaaGr2s47yV1lqT8HpKAfMOYbR3kT4FmyEuBMO+SI2j0bb1Ofcz9Z4oxjNjpxq5u
g2E5DGJ7Jtf/l9Z9hVIvCj0y34+Uy9tHoTkRzCFToqv+fOm6Y0rAYubiVFnVbHI0t8VVYfLOycLn
DuVVL27Mk2xNtBiyVRoJRPI0iFN0laqJp9ByP7tm2E3lfRghbDGB6CstmxarOr9CY6VafUbA26Q9
Z/JYZnLWXzZEa0x31Nhbs1Vx0eIDfzZE+AE3BM2i9d3La3aTi+QN5nGLwlhePyE2vfcbMm8NmNeg
OUt/gndUvbIKsczgUKDyy1W9yDOV6nGoImHrzpO01Eb0WcN2ejB9KPJjZffKfG4iQibX1czRSLkA
vSTP7NhK9C29N16gaSgVhjld6gQwV7plhnnavmmqg0pX3dSZ+mwaRR4fwT5ld1R9FEcF0r1M1ICm
8a9ZppGlQ25QXS/G0IVwHDn04vtf3UmrYCM9bNT4inn6YRtML1/ajzW/wq58h3l5DCly6UuFXI0i
9R9970bPSECgPKtcDd1ybOEr09+/BUByie7ISzBl3kdt2xtGxaonQLx2DXkjVy2xlqwSC6hc8EgT
hubVPo0sQkL+v/JNk83XQ9Ic3ux3okI1fMGt3dTMdCbZKXPiibPbj6sc66mCR6W1AOzYUNmGFDlU
Gc/ff5nqZnOcSbKIXs573tbCI9G5n/0/zFC8ibDBUlXfnuwcdFK5Y+THXhXTeC+C3fQdJIgARbyr
JI3+yA/0RBJ+I7pBAcs4aySCQsh8rFoOtRbGv8QFj1p3HXapI0IRoATAREd0l+jR7eGSHFdRG6iZ
BqyWKQHMGgMLHeb5vUa8ORNkf+NYLFVWneaA4nKqlz8ZutsrS822jqOGXLGUUdy3uJLyAo30u5Gi
iQNTp8pr0iR6IUcD4Do8q1iC6gE1LeWey8UfJIOx1/kzqn6bTxgHqpJkN/BR4Y7cVUdUkSXn9ApX
iLv81qm2K9ED3OyJzDGUNO0Rh8RJzZ7gNwxbrVp9BMEfod7h0TfHTJszX0dK1y4LlkNBk7qoCP9h
4WszRALVvlVP+nrWEudQibllgvL5uhjPmhby56Q9/dOr3g0EHExHMxzkMvJJ441gHFriTmtquPnO
hhvgBFMw6L26+wc62qs9Z7hDfaJSllXEomGqccKBsAj3KSzL76d4ueGFXynxGwK2W7wdPcR6C9eC
vFbvxclmoQiKA4S+Z4GZq4AiWV+iKgIh/RnOJCJP0nPajCiE2/v6EfX8eAR4Lam9gMicdTMn+xpz
7x6TpIIE8ZN+W1Qcts+asWWg3BdrufbEz+B1RaUtAQW/zmnaR1Wx4DyK6vXx9piQNYd8lK5pdia6
B3celLpAgs196Gunk8wXEO4Tzbhp5AqHUHrPG9EUjnEr5dTExYqMCIRV527gFmaKhaSxW99cyGu5
GDElCDPD5U+6tRGiEvy8N8xDcrqq1XJfwXkBDuvBCy92fWuhRZ/LMHVfI0UMkhKEl7NEqGwzTV/9
TX3bb//EoUPhm8gDt4i6grrZBLND9cPnsaTGc10hLy+qVPtmIyqDaeXaeXeBfLch2IeP3Q9++vr+
rFTthcTOqG2BzOihMPLBmlRFk8jTH/d5BBR9d9+xbVCvm1syA1qQ5GDt8eWoYYV8QpmSRagosDaE
87y+F2GiBqggCFRlwWjS9HaKP79tjxjQjljQhEn87SCVrNupZfeSiBs71UkCkrN3B6n5zg4HPSne
DbRTGqoz7t3BTquyXadHMfLSi/GXayj/aJWNFDzuUN6cjhusH5o6Y/afRJ3cKbeuDgXPMlmZto/g
v+NrHLwzoFDakBUG0M61TH9pXvklItw0IXY6g4XADmnKyY//LTHRwbh1B+Y9k1Oj33BTAuHHK83Q
OXFLZZlmLyCdfodTFQkFpPAh9pGG8reFlhogt2sBEKQyLdI4ljMe9NSIgrah+QsHphvm/a/bQSaU
bnrvvsaSVQ8BVc5u1BPnoeyKTUiaQNNhevMVgeFbl9HFX6q4kHvqnwb1cVRbfBvJBm7I8vhpgb9A
+o51vg27yjLJ1ghySwZJl6xTHwAzrndexn4E3uIy30vDjT5qbcMTOleKeUhEq3Nc2XzxU+Cx7cPq
6RJ3wjsfPQx2mm1gaa11C4kgpRA3iqgwCkEqVQ/CQCEBHC47jV2UIPAMBUyO28vOpLT/Ss77dkjw
CfblMtp0OAfUV+NVZznczZMIBxxa+pkM2zJKQr6aDk+FDFnFBLkEvU2+PJwKsX1yfc482zYj8aQE
jEsL4et/IltFP8CrFSw5tgkLVGNPuSiB2/yhMmfq0ceqiePbzURRBDTha7+m/g16p7vWEr6bO+OM
eUxuJD9ZYOIoYfBrUvqzM5S66yw2kuAPdxlUyyn9NiR6G5CI78uoPCkpiJSFpBgefGGHZyjg8Bbz
aMeZnsQR2FHDIuM0aOixx88ZlOlU9NreDoIQfZVME2kKeIUeX+xQcLmeFSnQtktwrxZOolNx8REx
8M66uL8TjGz05+VbYJ8oCXRYRVYNNR+Yt5DZ0hC3yTDxsR9i50jWKNC2N/5xrHVBCbv502rJlqkG
BCxY3wbjRkBMfUBhmQ9tdVeJnwmC1H0aiR8X1B+GnvJYwv6h/N0oXdl/wIxIVtKpQLfBgoIUs+kq
WXvuBIwM1TX+t8/7YYPCOIUmBPn9zapmfFgUbxjjJjPAGsOqpJt32gp90W0HiDSlys9hV1Y1jRtO
7/VvRUgr+KLZccscnalwYKzV6cDS1GcZuLXuGutP9oEOl7Mu6D2y0kHuiCzkZABJeOlcVQbbOvlP
lVdkPpa8yvuPTR2zzKkAgmgploSB+YN6M1cgNP7L5ET4JAKQPYZ4FoKe6FyGfSWfHLIG3AFK3eXK
WG+o9j4scEy4lKSBFLko9bCWGOTbW6VfqiAoYCFn+kZYFiEX7V6SEHw3drrvylr4xy5Pvd2Zzaj8
EOSeCQ6FzKTAhWaT8JNKB128hNFIH+hfx7LKhYiQxvh/JwKT36pKbqhnS1KVVv8Y1fSbfgcLw1Xy
ZtnUQUcPlRDVeXZsqX3dDfH8TrGR7LAxAQN2+PmXCDGVk3CcI4FLCRbgwhqgnT1dW3BE1ucrbDEB
Qtpl3wbP+O16T0T7aXE7Na62eOBoKAo9GvwGXyTQuh5PP1H11YHwZL+nsLuFi1AMlXdPapkb+JL4
pAW2TVb0EFpsEHTjYrYhXrKMrH1ay7m4ceosLoGtMl5ieyw09wN2yCW21tviJcov8QMqMeh5vgsv
+jBM8Ffn2nF/AIslG1iu2tTd/EBlAEtjsHsFHqIpaUsp/M+eI6PC6MC8OE57w6M8PryRm9cKa3XC
ogkH5rQz8sDBq/oJrrFecm3iiVdHpKOIeHNp5sdmlgo5w6SdTDkCpfp+8Tf57MOIKEoJgUXEL26r
ZG7VcirZdrKB6ub30IWpTchc1D0gszCrPXZYHef5UWXyO2xO8jtR/NQSj2CNfQNbXQogcaGG+st1
DLK0/RGZxlem2iq+vBoSiJCX6UyZ+Q0XDU96rMyUTuKs9rYQ0xWMVME8pl0XQi71zYK+c9h6VOG8
1CR576ETm4WUyKlp27ftjqtS9pjlYRKeQKmLF3k6SQdn0Gee4SrvjkEnPRFFFB16ULjmbvhUCRq6
AqtiFygSsctxq+p8IHmpocwMLy06YEBIDpKilDuqsHmsxPQqkq4UNEbWPfC4DjEMtyZmdKtNDdjJ
QCYgSxvAuAVQgiViYQcgEB5ZIP+kL1G7+ZUhZhT3yfdcakCHlIo+kS9m5lL/BCFAGwCmQL4FJUbA
urd0uK103nmyLDlngu+Fv7atZE3smdOVjRiahsI/b/s2LlK3C5OhuHCWT7W7arf/ImuP8t6geyV5
FECr9dmv25tLtxhwZVX7OW29Hh9ycrbEDzai8SfMQLYyfh46heybTQYZo4m9PZdvj6FmV5Qu4G1z
Mf2PBzZZ4OIz4OpFsZin5mXxE0Gz8mNFXtzJLYtwOlP0Zk13O0dpUvJAhZX0/0jQ0/N37a4dD1JA
etdZbVpQypZMhNXYLolYOGUfTHr/g+T6qzfs4h4dHQ+C9O84V9g5d5C0VgE5IR2vq4NuP2RqWSqm
lbq/PFsVIdorkCUrAZNvnArL7c1hB8QUM6Nb1EBZocXoTLI9+L+IdFkiQf9P72PZhrsfXXPMfJbp
G1p4rGAeJzDR88++Rm8ZsDkoDncRFMwaiOwvOyPZ7rPzxPL6zmKC3LVe/a60GM5ERviLVJ2sIEJH
cGbM52X8meNfZ/j391psaxNeP7vDF3h9RD3UqyZp+7Z+i9CNdAlhTncj8RgOzZ9HHRRu6tzdWcY7
iQQVygHCqnpS+e1e0EIj8YPIwFq+ASrrHSTNAt5MeK53eBc9Rfgq5nGyJ3oCQeTF2OC64l+RGWzJ
tTOXM4lwOZgoQDduFGpp9NOKv3m9CLvzzuyrTrUKoaoONhElFGVZX3/qJqDLSTe5zNQkEpxfo88q
o92/z9fvCXmrwi1KOUy289QpHP+xI9eoju7ZLuy6kHM6+yMomYe81TDpFkJFEhH5IDeJ+o2XEQLU
SPGekEsEoNPsP9immb8dCKvpyqYPOSd+nRgHXYD2265s68eNwVqCiPllvxg1Tcs4jU16iQAIBHqG
ADpmoSGq7Kd/5wivdj9w6CTkzUrMfVDkRNFG8q/Plyg1Fd83Nbv6F+zLSsgYkbtF22H4M5PvlW5c
zdCJ7lkl+s54WNyQo1Mg0IIWdT6hnKWrKwjniR5f7TldKk23VLQE0tzH4lLld18hn53PKsjrHCUX
P/FLrBOXf2VD+z8IG7O+4U6fKy4aRNIA0jKIHPUTczLyRc4J/NUsMHWWwrYoPEIyhBEdHL5AFuXx
J0Gwp+6uiIEckrGCiUtgHxYcW5+6y2kmor7IWifMR7AJiHqJuzayrfy7SRBg1tN4HFWbO2BRcOXh
aIHZKjjntajLbJXZobluAjfZi9TNJinvzmLJ/m+1mGFo5gVJ5i3um1Yn8LnZBiFwBfmZRPBa6I87
RfbPifjwZ7s3IA6QMzjnItuHQlH1Wcf9cuCugdJ4+cryqyWqAk2vWzwN75Htb/1/q7WQxr4Mwyjw
iZpvv+V66M0z5VmlMz6sCO4ogz1DX03E4cwCmU+ELm5l6GDE4wHDebWvYM5K2cwhPU+5gY8QRn+H
3Ehm4piSETjj0oS2jIq3M9PpO7L9UCjy7o0X+V66CpWgpLI1/iq4wHrIOAO5DtgfXUb737qB3SGg
GXOH59JTkN9H68imaummFYlWCgfHhQFWAFdnZINPWJwliLejzBfzcGNgRYrNNz8NTImkSHba41i3
Jycd9sKihSbieYSrZrGqRgCzs4v1AntI0Ec4W5JRO996tdYet6fPaJPffmgQqjLVgGV2D1t82Hmg
9KDUU62wGV0zX46t5FtMvvgGFozvoipSce7giYbwTCP+pwTp35XhnbxbsDRP739kRHuQrqrLBXhO
v97QHxWeetlkoyEh4I+uGzF/pehdgiOPLhQpODEu9Q9+Mx2z4NDq8EAjAI2eEZjWEh1ZdfiHmRDY
bPGjUygk8xUdzBtTP8ZrGASH5P5ndqtHMBrq1nVfO00xy0JxKwPCxAOhTp7wjlbVSRfW/TTjFFDn
ZD+6HwCfjQ8lEIQ8xJuPpBAIduGIWGK4tjL1ZqVCDOPE3E0jpKyvZK2YrIUH0s04tc3c/SNc02i8
gqA8bpVU89+GwT6bIZR/Fh5p6wMJC7j0J+a2sHEIrk6aEyKqXK/Q03hualdNA5QVf61ALZrf9Wj9
0JMYVEdyjoiGCD5xCjC1R0DRtxtXbCzLGT20Z5mfbLzVXuOEyu7Y2UrJv2iW2hdcySzP8iNubUiM
ruIyNQANfKOhN4WlNsvC3madh0Ap7Yo8ZEQj3zcLb7ao1oiDgZjZMAZYNvzyHr4CC3/Y6tYNWlK+
Z+e94F/P4yXFfzM/waGQW+OZJiH3mSr1jM6sbHZS+axXkir72ulUNfrCcJVW8UxJmdbs1smCYujV
woVJ+X2fsK0GlqW9qitEvF6fp2eu6LRPq0dL0haBcltT5k7u6VdTq6aJ4wN1nr9F3IIcmaCr/mDJ
z7aGL9yyLLGpoxJ+vQV6D6fQ5bhD/EAz1KbJciIEcpym2QqVsB7wznVDHkpd0EqMvEaKM6WdDgZ6
Q1Eshpi1GZd06OnJ/KS+zozy+1HbOfalLxyQGiEDNjr3lw12v3Yie1XaKN05lIoWqCCMZmniHVqg
bv+KJ/VdGQQ6Z1Yk9SmqszDDWCEn2MAFm/qViXRvzMwFsffkIKJ3//0T1aAkIB8a1NUNx3dRl2i6
IYeAcvSGT+xeLwzMZM6XiDO+apo0H5JX4eyjvqiy2n3NWb6Wf44EBBTbcli4zXFgDH+DZldVs1jG
tuvQE7SdZGgydxbvcq5sh42MNid3hTpqaQD1dwDT/Tk1qOINzXtSK6gdxAUeoICaJNaNqzZxq/Bv
zGuxB+Nx/2/hxfLr5flMFVaSN381wwGh10x8gDlwfcRG6QipgWciNIpw+Of8cd0bjkjsRGYaeD5p
5aJoPL4fXuw9wRGVaPd4C1XqPzdRhHFbj2CXOlCDQ6Oa3RFmYGuT1h4bsRaZ0pdhHMQOTglONwC1
km/5w9nWlm7N+NEQ4aDRXhMWBj+Jj/0nQq8SUADxL0TtF6LfZxu9OmhVvlIVSe5y1ZGbmd9yEzuj
ZMYrrOt2XIaOMFVap+MjdNMQmk1caohRCvdqgXBfVMYX0+RS/Uu0ezDGIyTnKKHKAt3OHFJBaBar
xTJxifLMkmqbaSJapAIWLYOED+OL3W3xVXpnflzB9IeZ6Amqade5rpRzL+7dKextaC53Ylrp9VzL
rArBhq4QZL8I/AX6iWw9rptV3uMB0CI0UQhtzWiB5bYQDcyhuMR6ccmItgUJF5xy97DFa0A9ekLc
tjxuzoV1RX65w9DDlVaHzSOrDg/mPopJ1HDRDyFwK9hU3JSVm2SyLOMG6x+oGTQjZudCa3dLNwX5
b6Iauy11qskapuMOY2n3P4ixHB7bkxuWO3bdrssJnZI3m4KiMySUcx5ZsxTnhZaRgCP6Vg0UHG9r
ZDOnJ8g3AyyPrzetZ/5rvMym1aRvrvCKKSd4MxC7oXOE/4OOxzRCU3z4nYxj57qS93QMub1TCrbG
nxE0bQOyJxxVFEJkqdtCYiWAeCUus+79yCnxzfsyi33/4MoeKNRAPl6JD9EbZGqA4rbmz00rtMEU
Z33cB2/ETaE/ORyqCqMMQ1Yl+tBCi6YrDTUi2M0ByfBlloTbXpBne4OX8gPc/Wz7JOm9m1GGf4J+
vL/4kqp0yvBDbrPOm3oTwMkU2xi9tac/K8Ua/xLv0WQrBNtU4drwVkOqKjTEuFbeTLCV+OYSTNAT
41nuxPzSSSXwnVoZmQDPbrrtZUjH9GHiGDE0qu4r+h2CjTSxIbbhxoRsYYLZ/Gz5JuPJMTjU+rPj
4WeYHD0QHLzftRynGTZKDB/HZ7MXqw876iFSGwG+rvC4QudFiLod9fis7x5V83Chh56ZgG96ZLfp
9/6BiXRORdDuDkQZOISS4xuprZvW8BZ1319Nad2c8u7SHw+W2tJ3m3t5w4vORhYJeQz9d6pCuBVR
65/iEMtyf8nplxbn09FiIj/wMc7pW79YVYYHjfSw9G8k9vZZpJfWMiso1DIKBhaumEhLsVOGLAol
P5OOwL/LgfpC78Q3Eixi7Obcrh4tL52MHd6p/wrqXskNgUMliGpciUWJ6TACzRQ37zNn40FfVY7A
VmB8OAW1J2spLJgorYubqhSsDJk8aeWRPZymgFFi7eVyH8a155oWEsK8j5Z4eVPw+pj8FLJ3OQ+e
mZ/jRSdUhT6txkTr3DYQFMc6aSqi4eX7ihNt8pPG7E1a5cfaV3+nfBfUJn3RwDUIpihkE3Ifq8h1
yo0hOsH4KNEspSD/pQbPf3Xfmrcd/GcYvKlMcB3+9s2JYo3nA56hbgZW2Q/KxsGbeDuSqtMiOOuU
X8OoutLw96F/4HF2UfRIqstg2C7F+eZ7ONUhlmymO8m2oXae6vlvp7RnBHapOIOgDRhrzpObjp5r
EG+XNC8c2n4eV/r2769QOHNC8ts7km/tetTG6W2vZINvnXDCRXRxdyBD6OjnpLeXILDeotkTyLYS
lM34RRJZlO/EowMbApZhHLmL3nmnepgTEQWoM5vTyP6xRBBCB4vLS0tnUsjSduEzDgoqIxuqYMvf
gAuctAHiCpdnOSxa+vCkYv8WoNKT+PA4l/GniA+nXIp9h603RHuLIQr8K2Yk2RuEkvNPzuag/ch1
Ie9sURocDzykyg02N0weUwk2zVoSg7BGCdc7tz+2b/ZeKtOseYBRdWbnsjoIu3HtmuS5IscGfvU5
IhcmBBEEhvKiUTKdunzrlfzy9JiXchrt/hKphSX6MrN5PuEjLGMltPMuYNqo+bW8V0iTGyGITr7a
qXFAjIss5X/lorqxlB4xf2h83EWbevPnQYtB6YhHlr9SQKwCucuie7N5ItjWF8oSKYmRfT4S2K1x
vyznM51sT83UfFqsaa5ISysB9S3TqQ2ijUqznbedBGwKRJ/7IZ7oLg1+eDrcug9HDTQNY7gAWPdB
ixUiq51MLljBXRDeJIO/TzhGqy/oZpHFs04sfJe9meeOMocgaqgzh+gPxQy2LRjMpxLLq6M3Kt+U
L0tGxdbFt8N1dHQFvSw4CBq+KYeACyTHXiQYre9SdiS2b312Fn9wM9hRK3Cn7fg9OBl3/il2eE3E
KsdceECkNZjmtEohgLMTCRu6udnzOfgwJKkQ1CVdI46Nt3ZnICFPMlhfCZinRj0zmJWI2jMX77LU
N1xQ2RqyB+LUoML4FaD6ExpAINI8OeOwp84P6+D8xDMgUwUJjWxmAU4BNH9dB/HQgUMeQFp8t4/Z
7xRT4R5r+ls0v8Tvi6U/NQ3EIn0VSkQDKW0qfQH60dooCvYQc6LCGB7yYpBwGvVImRIUwon+0s1k
4Hig7Jj+sA03AHqAM3SLLwVEDhnnmEvTyZC4pvfBLKUeVde8zCTRpIeSgu6Yel4gCP5K6yXBMymw
5lNQVicf4enoNZKxVyFJEvMNzZuKIRLl5HyiaFGCTJAoR/svJELNYvxX64ZnDsLvAFgGfk/E0E+r
4QHPpUSQ7XfH72+31yAEfsDWVKc8mH6rFDjSxcgPakf/D3xL46MegkEvYqZMD0TNyDjC6LEHRry3
cSpyou18phCXvI4hj9cdvbFOkBmiA1qgSmOg7M1aj6BIDw+IyaC5EQchM4/fXPd1R+UkVSOssn/X
oRWQVBroXNHaofA8pXJ8A4A9gb/oQmV0ppPbECMnYZoYwDInHQ8gpcx/MYSS2vCi6t9qZgPaoTCi
qYIFb9E9v7Vtja4W6F2DfRu1/7bHNA5GeGDkhLZPIOjXTm0I9TLJHrUipbMQ2fHXlNMODyf1Zmcb
a4vU6SeXnAWhc7FUdQyBW2im69QI9xkfsQXkJrNWM85123MQJdMT1laavMgxd9IKEjCYRLvBjyfW
0Z3Ko9saz6XjAa+JULBSCmMJc1lfSt5jVYBhUf4WQLbIUY7c5GXBX9mtIH/1+wwNNutunoMMgcjl
7Saz8fiAHybKS9GumUKGLdApGkstjjC+K7nZarnnNxfmxcuS+mze/WV+GWtPvns8Pg5vt63HNW2o
izLm5TIUWRV427rSLCrKKzhLc6w+02v+mSCEm8QuxbZI3rh0Qgjw0AjFxdhdrcvS5QKYggEku4RD
XGbxrs9vXTjHK+2xBKxkjkP/pjNR4VX90Q72pwvKsPcRho2WKM6auZlQt3wH+KjxG54Lc4UazVlr
ZW8+2+Ms7Iu6TAt9CYRxTH1AMyUeO7JVXhO5WovWRl16rREe3cEFeEnMffZF9rYDGdwpisOM6cX+
bQLAjOJdJl5PnstPczSzDF4sAcEsToVmXZPh1rYyeddDPo4KMipDWTnn6dYP6bSn01PdyF8Tmipr
KX9/iIKy9vcPGmfABn+fo6Q0FWYVp4bBMYB1hu/TGSQLKEeOwZ1avxkArGg4YEH+1gy/ObM3w6fF
xhevmFcvbesr1r72ExY1UvB3BGvsimHqC6E/8XN4n4+TEYbwWcuQzqzBGYQG1fmlSYyQONs3qyWf
vV7Qe88U6pgvtncddhIvTavjH9yICdZsBu5SDrdgAJEf0aAWk59X98+WlTcERcdkHjOvfQRP4KPk
fxjb9pPZ3fTO0m4Y4w5yCBWosd/ifrAvd1d2/EfCU/+6CBWqWHrNTtpJWnnFQKFapTiwILpZ2MlJ
x6q1NEa+ufJ/C8CBRJvjwXy9Ras68lwlyUw6nHgS3PTY/DL/WnEn2zfaUm0J2N+xODZ96BveZvvW
hZiZRSpYukrb5CmHGETbIvyKXJljGsovRN0X+qJy8ZGWEtmkghuWPThF64BOM/e97Jp2HvRTmZOr
NSWLyo3O47EnnwedI/AL+P9Z5F3HxRciyEZL+1ZSFXpdNvtDgavNRLPLLJwM3TOtPa4baCGogDzT
Pe8uHAUpminsSPpczNPF+9jXxWs9Xir3SeMuij883WUFWGuxx+vhF1YhSzsCFBq5/sSE4l4LM2ls
uAD8oosjCAD7q7RQmokthzz/jUga8CxFKF5TLrfdw4pXdDE/JTCaQwAI3vZJC7fkFmDTGVzdvvW2
NS/LEcDd0ajpWGdkkgU27pDQFjRgoKmKAivT7MK9/jKbvQ8RZI+OmH9iS1H2kcOX5I5YgldpIIMv
RXuBOKlyeA2/uUESYqRcBzGbm6JZoggM4mg+6UuVNN10qnwLNw1DttBbqGvQo6WwQznNnpbwEElc
L+GT5CQL1vKiTlSW0kI7IdVAYhWCigKLkWT/c/uP+473o193tShPO6zIu7sUunAbRi9spM8Iilct
ot8Gxh+4U8u5BOKBNTQF56n7B9r/ILdJGU7IZJfU8qYbRwNLKWhlUN9YIx+bHQ6i7okODK6Ktt4t
8m+8GwFvkZIgopTtpB5NdMw734u0FhbJxZNDxJ5/Ysp4YCHnf6sxJZkG1GU7u3z+FdltDY623tuF
APonkcXwjDE4eb9AyTsPnWsGNXXNmqVxi1dB0GoUnGqawo3wtOrYq2CoDqDiXnnJj1aZAfdagKgE
JBKzrfhJ6Z6BFGNK+8B7J3YBqbhXk2wdjFYvjbthRv4njGYPVa/ornjtmXw2LpVUMq2xOSylcMV3
O86XZ+gV4mE5XlsBKcid2OSmSqGpVou5bP3NQKmC6SSRvqUA8q01HSYDf7VI7dcrf1gUljEDO2hC
UJtE3mPe2+nIR+6PrPpaLS2aQ6OaZ/5Fd1tOXEmZ9dPW0WvnxLZBld1SB2OgVwLHT0MtY9R+gGHq
DWS8pux8wji1R+dx1XcxTX3yJxLnm1ogwDHDXypFXV5x+ETyDjzA0Hqbuhh5YB4gpwXaBBkMEZIE
GXAe19Jgg0hLfBhxYjPzaQZjAdKqUcLWoRXUrzZOwBMlEksEJ8fz4kc+P8qnf8/XO6663Y6xtgZs
FAon1OzeOXbIYo0KSWTAPphg0gH1fGqZiwmZ1iQ5OrrnmrxoPk/h5f/97HWdnW83nn7nbNf3m57X
PfOwMFKD7z6qdGGZGYm4SRITxmPZwVaZwuZPob6cfsndq5fBRIu/YyPU3in7jhirgU0AhOmNnmPh
Bb0dJNhUxtXgUWs9eaQ914Z2kLdRdpcXRkqY1l8igyb5g3+J4pEnmyuuq0538k6mjXuF6dyU8XqK
BK+/CKSqcHEa3W06J1sm5zLNDytIR2Ta9yyyqN7KOMFjIOJt59zqtn8lj+2Tubm3jzXlxBDRgol7
/tQb34BU81dtPwDmm6xpc1k38ZjOCNKO/cu+iIGkGfgYG6KdAv5oiX1xkffbMDhgO6A9gapAMQTE
a4JgTlFl60ULD3rc33MsxHSIsDKvZLVFa/JKtTxWGv5D1vjru5BkDhYqJMu2O9iUoki8rw7CCCy5
wKNRAWOKdfJeLffNFA0Yjwt0xFnUTLz1A6rl7Gw2c+Y7YIwt4Tomm5OX52p+nGQfxd8p9SM5dofD
H3BB62Qb48ZixqZA5SBOJYKERhzn+YRSTwt7ItRKPrHeCW7v4iai7+cE4letV2o7LDruY2r000Yw
rEjadccOTsQZ+dm2eDYj6dcLOW+yyK7vyOhnQibK4d0Rr5744+pplo9IVmX9P85mxecGYJKg1f/L
3f875M4lTYf285CMN3j4MmPv4kqYf60tCqhKr40r/jWipj0mriw++Y4vEdQXMKYt+PXh7YA0luuR
baQGKIa/5Yry+PQIPOEm8qXDEOIBktQ/xnO8PObyGh0ngCGy3PjVHPSQKiJl8awP0HVvqtt9qVwu
HVVcbSy9xKyiyShQ6WdmSxn0zdNm7+afwf1XOkiamk2szQD/3BQz3zwbwJUEg6LRa73wYie1Xz6y
Izq+b9IX0e4sgthGEE/XpHXfJkq1a931Gj/J0JFrFfNWYHin0xQmj2Ld+5/Qws5KmwXy7ucsuQHE
NBKWCpfvkv8RZVx4XlhnlK4x0fAfYdtP6hCDRRO5/ycVe7pPvOeoiM+QI49UI40ZH3BDGmaNTSNs
QExSyEHA3hgOpPisbRNBK6oYmZx4XpEDN3jaZqMVdbqJ5bq5f2xoS0eMRpm+IiW39/dDj3VxB6MD
IoNf3zwBIwoIerhp0pFMl7LuKUOfmW+RN+F5ORDyUhHNqSkRN/n77VA7/GGREQEbG4aeCYoEpAKM
qA57srydLkOBAMn4mz84wPa+trBvYAZnwaKtMPZT3uP9XHyiEw1XQ13+KMzrkw2RZCouEBOA1DtH
zVPNuVsAJwedC3Nz+5a6zAAZlMFVFVLmT+B8xpis5caLFheInobxgK+VpdQTCWZy0OF2jHf0elA7
x27hxgYYE7F/v3NCdG5Osecav/KuaSjR/S972H1gndHw2lF8c99lAHrA/MCOeewIzukfI17TOLqN
j/wAaXm34khG6IqIP4L2nnH4VRmp+9xmDRB39+s3Lu3fvUhzGklUfLXfN0obokXiWC1vbgH8/9Ke
1HDe5t1VEvEWeDSdTq+yOmFXgb7BDLQg0MGdVMYpPS8z1hViaswiUoTdO56XNw7Ivea6dbchKMi6
uePEIE3JAXGNuuC4vut6Xls5KhuDFRqJBDLO/lVvZtRPFGN8ANPa2YsA3FM6sys7QsdLwFXx3deF
oiZ2PSkf/V0VjDLDVvz3oX1yoeGqiGGDJG6Guu80TmTYP+HvxILhGAK78Jarc5eKSDhawrRtZqwS
TPISrgUcpOyynyTT8T7v84J4eAazr83iFwlt1E0Up+Nxr5MOxTVZJG1cN7frrd9wh5fc3LffQhIg
P7yr2QSlygq9H2qV3dKX7RDe3Zv/DInwXx9SnKmru1Avolnrlu1nmDuNLHe8TSIEQyfrhPC9ckPC
FPoMI3wkUcuybe8+wrpkhFgAdc5vrwmuYXZDTw0dsMM46YUjS2U1C9jXxx4+4JKO1KiX3kM7FRBX
r0ZjKTDSVBV0B1mtXjWXNhlzLEHibuJq3MW7Cqohqc2G/4DvnFBPUR9BvAPGIG9MIjf/TO8vgdKs
1d99VU3R2C/6uu5+KQF9ZZ5BaFdLjS+Z+fCDTrQl4yoxXQFv5pVvtw8q+yCHNr/FCBOuGdGaDeHo
AxHRZw/xDDOJyPJaKFeXYvcHz3a/cksZMk69lS+8qZQFL0tVRIaADHC4zSZQESX7It6g+oGFXVgH
/xzz0gqEPT461dZ6hwiG6CRHkw4eqwig61LV6u7YaLca44mXYpKejG1i+VVkl+xi/NJrmNJehd7J
kUHtQsGi27vYNzLU1JbHfDDpP6UawKR2v2a5Nj3r98LgJT5Gb8UI62FiVVQt5zRrBk5P4FJvrVVt
asQfSBmTOhIlu5JNPonlb5Gl70YN4ft3igrxjjhM0sOsVGP18HtoqadL1Ko8aGquwkds6EDZUnOw
dmxmmE9iZbp5bsc3Cbv8uGTNaYFRT71Yo//aemc4IQD+ywZ6n+XxaUagivDAj8K8Y485TzAdStEA
jVtNf4BFqjFAooKHLaCVSgvZkGUFVx4XBouD1TF7adoWjV29ly8wuGTkYM8QXGi/5WxeYmC00iJd
KyAY6ful9iADE6BCpKblqQOcKDTkrs9ox+LkM/Va+Pz/BgAWJnUxG/KpC3aKS0dA6jEJtvKacOxk
2MgU3TWGh2bLFVBiubjB0/TjuPfuhzIIzdZkGJRYLmibMFnQK0wcFcPYaL6FKl+sTcElql2BrZ5E
EXu4FMmALx6ODtcASlxmWlUAzdWhLB/XR1guUv7dhuKV5nhICsDyplr/xj3eL8V5ZzKSQSxS8Xgi
RwIEs8PwVYCU7+L60KC0fEN1VfNEjazJXQLM9Um/U4XL8Kb2Wqc2BFVzVIZqewo/he+oXPShJPey
yjJNJjrxlGZEl9EVz0wzgFmczMYU8PZCm6KEFg8nA3g0aLkhkUYGT5NhpBO8F6uBDVMxpETYXnwv
5Wq+moXxicUHa2fZZaQa/pJr1nKr449t/NO1hoT9HvtcPwHfx48o2NkGKqHYn9nq3kIK7oGDiPXz
ZBf4D/6DCWiH28sLNSOpxcw6VJZTJPxYEUwj7CP/U6d2HoyYY8K38fVXCWGJ/32itvWkeiow9/zL
boyHjO1PhS0oG4Xi+MPZYnZrqQ9XT5qvHFLzvHQjJ9WvMmgZzKf6zCaURywovRaKpPIwjdDZ4U1j
4ABmwqmX+3HQxT63okzvSJc7pEO0Ksaa8Eoy7EcMDa875Oy1vfs6FsYcmBukJaTUV71JDk1W8OCP
GO2B5yktW8qDLX+0S8MyMYbk8qnZd674Zvl20Mj+/+NVJ1iVNUMLfaUnyNEhxNUEPN6YYu4v/+p1
642187BRmrB5tvGRcJ7cG4iYjliw/RVYtTdF2XFxa+mutMeFqswaXkRLOOhBB/hOkWuGVXisiRS/
E5mCuusx4v3pkNIV3hh9EX/CF+qaTgCV+5flaWv35KsBj39qhmTPx0XxVuw3pikrSNG4AyWf+yAJ
pfLxh5986Q4X5e/4yELFHSLllWlWfhdU7GkUMw+TKIch+bho29mEnippy2TGQIRk7DjpUOyQxL/P
ILU45e5fz5t7WP3v6FP9GQpqgBrblv6aYQ+hqs5lpEaNdFkP5imMYUXTi8Gnt4NMGoLAfF7q2Amu
yhZlIm3yeuZutCd/5tMqscv3LTgkRjt0E3aJMuA9koHS9/mGCCoY/ETJL0Qwqwx0DdZiGhWfqrMW
5+YZY9SdVMPGz0bZ4c2N9Xx0GpYDsgdenDNES0WpyP/8HCkkFExm0/A9JBat9vZjJsEjpPZ03wpC
auOZEWd2dwnkaXAyPYEwmoFazVzkx6T/ubqR6BkorUmxxxdF0MeI6ImJ/PddejBaqpNoSkolXseI
TcXeZ8UFagcsyq8QQFGJsCUhF2PzO+miGZ7t3mM2NDNwvFgrhgywuutk/NkItQMaLU55oIGXefx+
7u3wcG31sKJ5HhNQ0dZtVleRASmmKkMqktiok65oNKTOEWFMVP1FKYoWNuMkBxmK60R86wyfVXtK
h7EANi3tqL0gPTOG0ekxLzbSDC32FN9fzVrKZrpJvQAFBKSvJHiKHSG+E+0QBxhmSS8Rsy9Nq2aM
EGz+fSh4Ppil2XQrTz7ohTkLl/YzWMYd59d3Q4Z7FokQ7V673K4SvIF61PSFVtGP/dGlt2pSdyvs
gHBLyrk3Yy7FBjLTJZUghLpDX/wEAyl7Gp/yql13R8IgmmF3CawT68Wxp0y3VUXf8ylS6gCDQ1FE
w5IBzbrhNsol932w87eIEhFW+jzZvFKFYXFzjg5EI1Xlosi+sM9Nt+3KiwtJC/FhnYkcC4WtGUyi
4/IqUCQxdVq5kmyXqACbmHkMlDA68UcObpy7WzX9rsRkqGy6sFXhbWG3S1DsYoiiFRD+2cdIDJTr
l+ustQAe3oJgKTYvLrPrwurFs5zDF+6WgTlcsJaJ35qnpuF+hSLlqD+oELnTwlGLyETVujWCxCny
S8svF87MlFOMMsPCbY6Mp6ozsfJ+0RBZJuMoZwA27XoYEH2vq16IZtS6Goja55VfrCdpCc4g9Oyd
b+JZ/ROFUsKloGs2iaCjtbWOD7AWT3MOqtBn+wViKyzFK38vvyWCmB4wxdeNMCoaggL76iX+qVul
wMfdMJz0jxGOoUbTlvTm4QOA/bMu1NI38cUDvoxh5ZPJjuftMMUB+DumbydTH+j7LOrgl0t0FVMf
KhkeUY8zlXAu21Q6Zzo+1hn3uB2jaNijVRvHwevqA/KCYv61QDVMdr/28cJa6TlFDles0KMcP6Fj
NsqC8PaWxHPC4MYd4RrJDbgpRySBF+wlmpcPRhcNpPe0FH56MYZJpy0Ry46mfCslRsq2+7zR2Ida
lOxK0etb2p3BZLcwGgS6dme0kkRYls3cU9Kmg7tP8dFb8E1ntpM8U7tEAGJWvrLLIepwu/kAWheC
SAyIYvW+3ehtTHCp8BMk82H5nzNmgTbKBXQ5Pr5n4ttzI3B4ABJrG1GG1O04yeKYlZUzHF9Edw7U
aNuYt2vEWL8895NDqw6mgqVNa1CjD9+DSY4QviD2kX0aN0OEoi0+Lqw14CRAJdgx9gIv0I3jObtM
e01caUOMPi9UwDAa2l4QHOrlbTM14bU6Fne6TzqozxYmStYDMJMK5MHjU2pU1cPHtSem51vtNX9M
19ZPArtBM/to3YuwPDvKPbgip7ypEtW3IaiGI0q8A8B1HhpWXb4VufDP4Cq1PTPfHHkJCK+MPP9S
DsVHICdTFt7Nx0r3s8naF/JiVWNQ9dZR1fvzWMESY1k+GNSnaOVwU4jzcYZP9N13iDi5xtsF2bBb
Mgo9WX+pau6KyiLrGNxyQqR5Oz0V06EsdJbc/S8P4+N7hWICGXYoBQfW5mHodbFqvn6jesmDi3Yy
1EprCVWlYvsEhPHN/4Hx1vY7Twv3mehncx6ZKIGCv9Kab8bziGeJpbM/u/Py3ETAvDOONGOqGD43
zwUQFX+osPwh6OX526cPSziaxUqSIDjm0YJkS1SoKrNfGS8yZBgkSCOMxeb4AGo6AT53YAqkQUWk
7vT0rDmJBEUn5kMS1WMfJpbWbgwXmPcFKawsFOJ/pLLlIO2DhZffTXf6iUalpE4ZvVnBOPniux6I
VeVhpC2Urr28JbnCH4Q7W7RFqkRkCRZwXJTZv8QSMS3yEgjpaDf8C8DxqMHhulFaocreeMXZwQvJ
pgGC+vZFlolcSm4ZTbazmnqADu6/8lXc/EiicNXlFYL9Y832ednDsCIyWn1dg3DAPXdhXufd2nIK
QUyCc/pBjgWR5eFiKhpLubdWgIEBAhzCFbmxjr1MwmX0LJK0+cuR0VPVoDYeNDXrRry5IZqWYxIs
BXobN5vlF5zbm/cvkpr15uMzREhDqQGhIjIQdq/bRkXd+K3iRmUwZv16ul4MquTbw5oaHoKMwSX+
N/7G0XBCH2RSrHbUuagFoK34AgXoYOT7y2nIjjkuVg6GSjuSMcrEQUS/4gkITEqvv47AtehCWYYt
zueqDQzZB/I/PiyLP5iZeJTUZJKNGaQzVteUz9qNsxC+kMsuURA61x0h2ufwQOHn/oc+GoBmidUV
IU5R7KrwRMOWZbzOkYBoIlEWoymKiKZMkWRUbSoE3CkpZIYTpcYnFBhuP99qhirhd6nhE1PRqbkT
0RPf/6RA6yglen2coUFqJRrMCOXC1RWN3vpmtSnzZbEPpKfXSXOz+cbEQF8+orB+As1URZxFb39U
J3DhI7N3sCvTFgs4hE0NZjuPrCG2ih8G1kklOTxrY45C2nArMkaUY++Wnu3dSty8Rze4PcyCtNv/
LgwfWyjeq6WwbyC1HFSQwVc+2aqk9TGfeMHeZX68bcQVou+0O9SVosUwx8K4gGzQAZRTy43Vp/Yb
W+HYX2qj0qQgItBzIv1UolSuOELz9+YFT59p5QT18W3LxsYdyzIfTOz6UnuBJW9Y+lFVnOK46HJb
Q34hGqe52XSPNidXXRjXMBqjk8D4STeteXCpnEa2tWztvI8l9JcAhSs6NdtHksQPfPoQdv0mHR+g
lSyaktJevRxFgnBZFblrRtpemST6gNgSTTzduO/0P4W+qEPCLwyOepc+7+LmH3e2eDcszRc95EcM
Ekn13jHqEJwckEBmtmOdQQjjvCZMQVj8xELobyZRj90GIdJylba3bTf+2R+odNqSMlKiyWXQDdr2
BDoRtUDY8c5bffb/OAfrmV2xL7GN+zlOeV94roRS/HuUTgPVfbfibH2SUi52xz0KGvoVQ1qLH+K0
CTQ1uD8Bwdu7GzrMe1TykGbYnigTTOrcbfyAO2vdPfkETRAq9vaLSSmKtXqyfEn6vlUIADaxqjp1
/vs0blV/jjhou5zwbuZ2XxO62em3up0pC9M2/ssA/r93btTmjcy5nPonN4KeQGXTPgqrC34lMfxz
+zkQyXK8JHw9MdImTNw+8uvdN8Zzfz4mYEyNVWhqrbWJOe4FZ5G2Jp9UgHUGZukKYHfIvPCZaZq5
no9y4gb8UZ+Z2ZUosRUj9+E+A/x54q4rjVz/upQ0N4Hcn2zxAe9BWl0t6tTITJ95IfWebGSC+ZdA
ly44IDmBzcGe2Bs9rZju3zRRtuIb4YJTRBCa3sBkKyM0VPFQMFf/4CaiyfPAS9Qd6pKETGKAnJBt
A6cKAC/L5CiWKgOOF97VMhd6jeCDphSFBXeVdZRyCHp84uJS6ttXuq6n8uEcIofzggsaMxF5wsg7
9WihOPvyJ4rQ6EGSCi1WZLAOfm+qakK234j9bA3fWZBeEOQeKkZN76XD0ekZS3KKsszXr6Y4NDMW
eEbljboVNdbxQbK9dcCjCsstBSh6Th1xdSAWQ/kjk1sPsuXLdR74KNzilSqARA+tK0NOFyIm12/8
02Wk+t/63adSNMJb8oC6K3EuRdehjl0nRSXBoL3h3/Gu/03D2vrjghMELW0wPGQ2zuD821+79k0q
E3xqFG01NuxujYLXA3GBGpAAt1JPq4wtdPlNTWKPfK4Db+PMgFgf74GCLTwa/cZetn58kN/dcrgu
eDm4auiqeItiMyXfOyoJg+GlQA7ASTkrebmLSHhaQEXPJC8aSPV9l7TBAPZevmZpNiHM03ar35R5
yW10HsAWGhxmLISxb5a/SNnNd8lkbk82KssUCKLNXdbqjO1gFE5Ol0T0Cbp4r+qHlRUk8eAklm7B
A6YPmy3SSktSyg7KevlHyqrQ0j+e32wPTFnLiM5nFOygaoh0Q5sbg/k4k4aNvm+PmHhrRENgcAqU
AheGIU6nWjzvwnbDTHwj0LcbUJKFM3xLSyCFuln69rnli5XYut3+zbZNElt4rZydgBvKef5iPSsK
WnMQODRNb9labWXmA5gntS9BlEB1y01vJh789+RYpR4RRh7UWoNnwwgxeRE16UWP+c71glUlCFfy
zbFFWg4xjWw5kreYtPCmb/wBuB2Ic+6OwrA0GddAmencUyLv26Yuc5tUVy8WiMiCfPnXtseIX+wB
3sPGRcWeaOUurXbpuu/KQ/DhC0gsnfo463r7+OVdSGpBY9kJ+QTQ35NIy1M/js/5g1dHVIfpXaZC
xHjvEcnk/MoxJWtMKTsegOJgBNejhX+YnD5lCGYjlGYxefdV+tp4uWXx0M7aZw2A6bewCQCmclpt
C8DRc+IUlqElTM+JtBF4mJJbFHyPkwQh4lbjfNrzGW1XODtcVAt9j6pfvwrVy+RuTXh93cJGHhnM
iyGMqXuhXOGmzMdYFB5TG3KmzCHtp3ToNu5Y8zjjPfgQjMN1j4bWYGwmDvug6ADpZ31qM6/5hEOP
VO2s4yXMOYd7uz1RDJ9vVNU+hvatUmsiavQDmCSc19kOol+bwhSLRks7JjZ6yeyDQFr1AqBBVcIw
2dJ/LrFlEjnJMJDKUrYDa3uXp68+otvwnrR5IaLymGCfUalouanSeoV1ZHFiQbCQTVDsK+XJ75Lg
4w2GD/nxUMHigiDLWiZndhjxtnzL7RYT3/mGtx0zkqztPXGQs8HyCf9KxVsK8QTFghhHhNGKcLCY
5eoiMBWhMX3vqF7SqBQaPac4N8/3uhFh6YN3jOKNSYXh8l4z6at0+ck3FJpQh7VjMBzKTaSdiY7p
tH9pd/WtuJikULg3voqM056WIGsP/WpxbkgZK+ho399ccZRZom88Bdy924igxdCI5i9TYCY7NZfc
pEUsfPM8ztbVEjtzYxfe2lM/TDGEhhJmqDNpjBRrPPiURFdMlwnBiS08j9a0YoH0zOLAdTf0+HGq
/+mOfL0E41GSdA6n0TdZcxYpZoeSb5A3nFMY4BU5PgONNU2LPyV5Fc2emvW+30lWRrcKCVQRfWli
oWPQDaaqJ8c80xi0KPjPBgAjIX0RcKJxoCSeteSHdOUIn8yYt232kWT76URC7n8n0jnH7fwl7Dzd
O+dXVJ1JQBlsRgi23if1D8Sx1kYzd9b6u0Ll/Rs58n5+VSy8V3r/Ky7zcvKvfpqfoCXaXnCVDOhL
kbecZEqAOF0nRAbyDYJTRhFavb1PnqpkpzJNd+FPbxBE8TzbzeGi4aXj0ub0sd3qi7z75ddAxp8T
Pi6RxmqW5I8T0imPbRIIh0Qw4Knnmc1wYfeq5Oz1xi7vm8ZIpsGKlumO/PF5RnMVB61dtAzpOgX9
gBFKubC0yG+RmdP0YrWKoMc2+0nFSCyLtPkTDNgqerqifI98r1KVWnkn4W1IIHw0sb8ZWyLBaIIy
M3dGonQYxj5azqmk9J4oFIkTao8mCc3A/IXPYPP2hywVbapUY6CNKt2ABEf84b2AiAT20Nxtv04d
QSsQ7MiwH9Ucq195vV7KmH1eO006sdzlX+J3D+BARmM1593rgPeITetf9IqWhU53pxck613LyyUZ
uYS/3Y4/fA4NofHySS4Y0A2v7sNoILDxPx0GbvftsliusCajG5kGJQjgUuxNwpE3JIV/fWlVhijm
XOrVXW1NQNym8YeD/Yvy0OyfrqB3paD+slbI/kUUZWXjV0V/olYMWGOBDKXEvSViUgrjr53Nt8m1
5idSpvPGFHhi6/5EgONKvZFnQOhOMTOEYKe9TsI990663qmGJJSsMYzEyG3D1mk0iJTx3WO2kw46
dHzhO4O5l3EQJqzWiJCZGS/ZzsVfZDOzc20odfMPaZpDiDi8yrP1Z82PUe2uWtUJu3XfpF6wYdrx
7X9lzSgXaFMQZCXc5htpUOv53Vy3a/pDuC+bbxm8Oug/6BhqiXSBXoGmC5VxaBNPB/q5mvY5OJZC
qYEOwgo1y9keZRQIRiW7oUaa8qXmA83p8xSuxm7cxps3IDZEr93xZUTmUB1y5sHtTeUqNlt00t9w
XxPDAVgmPV6zU5aMN0j1Kd8Yey7HDVQuhh+CfPzEFjlWkaCeKa7IOaTgKBzyL9NhKB5gHw+x7XVa
lG3XM4ic1h5BYgYf7E+cl6yS2hVLoRxqU7dNWh5grLCiGt+uRcXh1lqbf7iEym5DNZ/xPo5TPzDA
G6xP9xfEH+hs9nwOE+HWYtdEfzVo9P9G+2eZ6DjCDVUIzIO8QlJfyEqCeqWxW0668TVnFuKdwzhq
Aud+ESz9YJV4gZaKbAKpUfzLAlQXpuIW+bJNLWUqk2ex2QWAsRbMDyqGwyrZGI9BFw7KWC2nAxV8
O+DdPBhV6aMpSWVaWb7BmLD4iIDucfQPao/WiWzTNfZDddaQTjhTOgz0vpblcsowycg0VPiFrrqE
AzAT+nOoJPnLA1bpG4FXn8/+cGuDwKGNfXkJLQomE/ZxJdCzuH3mIZPLcK5LFlJTgRmx+OcbeOXx
3UHESUiS1m6gLJ12+3Jrs2fY8fjfb9qzEaDeh2UgwrLIzFuj5pGOHdmF1ll37dQ9etmwXIduJcW+
dS1LkJa7LgZp4eHFw7I5H92Nyp+7+nbPXfeLU3lPa9BxmT5iuDHRq/MGyX79OL3KJ71N4LrjFvAB
LfHnjrkgA4K1Vu5MwFJF7g37iBVBZW8QUG/7ZK0Orb4w6DnxzbbOkMb+rDM9apjSuu1OJYwyvTeC
qpVpNjw2wDuO8AIkFuxTUR+82c0oiz2Rp8w6he6CcGWVWIkCbca7G/hszv+G6bcGVAkuAlb44mdg
UGJcaeAbB5JZXiP+YseHM7us9voDmd9AtjO2sZyS8CakuPpcPbZcL+ZQwmm+SIt7/GA+icnlEKZV
tTo2+tFQdeieC4CHC85xgMA7JCa+ZW8SlIntrX46KYAj9PP0e5BLTMjyYcRdVAxoVtXo+rEywGkv
LuVndVbQNbvuWCnuwPMBWXxFlJ8nb3qdTlcqnUBmB9kH8+ZN4l42p1iabbNmuh6zYF9NA4EB3+/X
IL+tvItUJ/sAvVOqIHdEHidxH9+WwDLvU9LL1Qahy0T+M/wSmTpKbs5o/e8bia4q60ioLhSow+a2
59Z5YX7q7VDwodqUiiL0l/gAXMdmTBlmxXCcIl79Vec3YeaGXeGkoWWTfbwTrR3pOFC9Rulctm8F
j9pMaxorCrJN2f0KQMScb3L9lcsbNImXsKeBADTroGZKdSO2TsUjqZCqYW2D02jZcmlYs/iUWHmv
FJREsdxV8/QgyhIdNrxl0pqfIuSBtb57wyc0s1BQcGJl/yPpy1xg9q532lwF/rLcH70d3vl/EI7R
AyJ2l/V9idhT/8xf6uix7FCWupQ2zzqGXasnsP0JWfXwFP8ikY/SKDq9AmGWHkOu2iD0Ja5jf2ZN
ENnjfBHsQfKN/hlOkH2R7BYAmpq+Bv4MzFCuRY9MmK61sCGxkPRC6G0KwAScyUyQr7ANw3UHBiW4
1rWsJLRf2m/INX+d0KlJYT46iR6M+NzBOzU3j9bk8z7HZMiLN7nJe3kzqp+AAj0pVHJaxAgPHwOF
7SDf9OihFiAIPqunO3cHZhqp1/zdGVFpFn9/kKUEmz2R0641zbohIACaJ4mWTwd2fwsRmubveP/i
hcuj/C4YBAr9mCyc1/DuFM/q5uF1yAkO5l/cT9L5GCyBd1/ayVJVBzrA5bfww/M7HqW2GqlvKuVS
G+Wax2VZjHMf01FMQUUscBVZX9Sv/F6Ld8Z6WBsRLg8XdvaPTl3DcEXn2Wg26JN/No7pDDNg8akO
yAXJlyWgDDGSs76G1SSCmx9FVi4d05QM9Z3InYyCbC5pYV5f5rOhmZaB43H0wOjRsZljE/iZVaii
5tfetFzXk/lN9RpGTBkSjhJTCRIO96LzbsjqhwQUYXx26AIdQzflfSNNr2bE9EyGsbPVNIVKVxbm
BwTxM+QDvVIE4ZLzSGXjjhq1v9l1jPSeQYHOe1rIcuDrOIG2NmXpFyAGn+1Oaz+CJxEDlNDFJ/7H
KzXSpMx2NRC2UWiOyq7BjZoOH7NX9h9/uF8P0WL97hWgMFtwZyCryChO7d0Oo0+rJK3vilyoxDbW
oAAwW5AsbJL/+p/bhuZORtaR1d380dk3av++w3+Jk5XOX4OTLpJNZe0lQTbSk6ahzje3d2vxx7YV
OK5dcyFqtmlqoR+KaI7g4JLvFZ9TYJyGvEXRE+0rOas88HZ0mA7f3B691kWyZpmjmPrxUYubbzvY
091Mwv7OIrMbahhioKTeBKGh850cZmJXwe+heg5r9gzcu1QoS9xrvoPszXrJFhbu1Ooy9MUQs4Kk
goAxY11L+ZhgflWZvJJynLVrEDPmtoGle1s0VxOsE1QbA8yxjlbyn2qWpv6GxT/fGW/V/h8P5njH
G2M6uKvGd6qyNV3UE7QviZn6IMhkydhoywCi/yYtI1i0nudtJOJs6GoZnSOTEtEyRRy6Dpfh3anK
zsoeJgi1iGhj7GF/StPEnl1dr7Y4mY76YEwQZWWh2yoscwrXu70vDbTpec4oR+wQCTiXisna5PKf
p5orayT+KYfacJnGgqg/ozheKXOnSwplcvVzJsj1k/wVYdnkTJYrtFoCBniJEz5LX/vBjH/teH4G
mxwz4tCM6atbTwzpXmpABig/Kpo3HwCWaT/SLiRMGk9mDfS0b8GmvtaAfOxQdPb76xdevoweZbuF
OCCs0bwOGjbbMvUTinwETfNMrt7iEaxktef68tVTV0tcn67SwBT7O2WPg/oWtfIs2as01JsjU6cc
TgS0mTVoQjPiWHdyTjh8u3EPprAzPzgm1MPu/WXL3sW5yhucKKCalEe4wA5u1J8zWFuApPd9oJOJ
STJupItp5fONixzo6vhdmYk/gQWF9rj5grQlJ7LGqOHWkExecZgNdlEMxriqdmuEYxkofg2Y77Ly
bNQEB7o2Cdt6fHgWdy7OzfiiDHjY5xnYjBW/bpCiYI1VBoA9kB9A6ghILlh0ZBnI4t7PAgFjwt9q
M0n+JvHFoE3UG3fsFKVu6GgZSyDMuxPLZMaBLBxy213LdthDNzlkJ/oSc6Pn5NPXCTjunWMyjKDo
aI7Ie1t9JH+cSLYBAEE7B8Kw/scxT9rVi0Nncecm36zYF3eHjajIggosTvEpuB5YRRG73UsDNmm5
hSdimOUSIImOJUIvHQsifB1C/E2oSepPz7K+NgTBIabhM9We9G5bxZSuo6ubfBv7x5qHo9Nvso5a
Ci13cxW+FMCXWLAgFm2NerkWq/MSibdt8SdG/SmkTD6ihy3hAQQdHx4bkeN4Y2wsE8+dV+bFbdBQ
OIEbZcuygzW16AwZ6QF6s7+MMqq/aYqE6xcW7xGLiFIm2AX5R2aEa+Oz3cIJc9UlpKI+FWWmaSx/
QwNbM7CpprMXVQ9CfGn89ICRGIVQ1/oCVSYU4n0h34ssZsFsRy+JtHd6taO/ihT8VqJQl78fEUmX
sq3cfiKYnEfu14zuvSgx+zXfbFNYWh2lPxqo82M7hopxtFRnqOZAzSGYCwkEYssPyvS2pJVVs97W
5A5rOn6CdKILlefuL+qf42n5xN3lYPjlZ4Dc/0pk3DO+MNQSO5dor6CBiiZckCaez7kZF3vVpCIr
qaPkSt+wW6EeX4uQ/3WbQNdPFKPaeecngkkLFjyk15NzKmGjtzdG9nNlT9Q5lxkvBHkFXdFqS7Zc
40fyLRhq7ZABNKhee/fsfTPhhTkQ9ECQJMPZE+mc5VorfpP+wlOrNrMIdUnRjppPimnJsPxXvUKz
uOXrUFqWM1Xu0VcPYiWL+wJsYJnYyMG0rriF7cjP0AyKYpUAMdvhCMX46UjurBpVPLmQMCWQDPuQ
q85PsHtxV0F+8HqxTQK15gNai9Rmnc9DrW+p4v/CLdnK/hkQhJ7L1MnXwNCsa9rauY+RPUOLCBCg
Y4HRdATC3bpgs561pns90C65c+nnE7Li6ADulsSUMD+05RTuGRJ/V/l93Xqibs7M3V6HjQRIrnNH
a94hEGX3or58hkVr1VC6oJEp6b5w3AnYazvmr2xT7ld1Qqb08LaX50hETQzh0A4rc4YTQj/W4f9t
xKke208tZRFJHZek+s+GmCHLU2YepsAsPzNLq55i1BfKSlKZFz8mcUpNIHZqbdxtaxylU1k8NUZH
iUMRxG+YDynQa2KPTnudoqA/TmVIa7pLXqdBC0VqaOlG1KkmvCEGutKnlqshdaVrYG3fmh9xa/a4
5hAMP0WDgy3Np7Yg2RUCcaouf11pFc7XHrIkFXjvQ2dpM5C4BS3FiWHmLxWN6eXb6a2JrNQIEOnI
aZsrVKBenA+C/ToSoiBwhuKDg8o9vD96dww0Kp6ufCmS/cU7tgGu2NwoUkSw5Vg0L7+SMAJDFbUY
nFUwKss+AneazA8Q3yyBCUMMM/uCFjJgHQTEmh8PrEpS8XH5x91eg8sjAloIPubmeSXVcZKpHxYI
s+OBfutvvXHMkYCrPhr2aUR4uTox6/GIUg1LagISjoSg4Qn72gnwFCMgzV7qhORPA2sHXLakmvoJ
37V092o3klmsE7JkWO00ie9l4jRFKTy1l3Onwk9LUUHsNSwBD+7qvzuHyc1OhyjZ8JArwHnplPwp
vrwVa7NjNnWt4A4Xj0eMrkR0JgK0HoLAufq0axgW56OaRZ13k+v+Rtz0xjCSats3H26wKFhQCuCz
7lU6qgLNt5HxvNf3H+FooGlb23utgBPuT32J4R7YK/HR2/EzBWc9YGVZyjFr6wRk9tgNni+2Ac8e
/2ORP5PSr9PmRsCRdEmkrjyrdjVQwiyUmRck3oaUUDBOq2O6MDbHsdQ4YrV7OByNpNrCm+k4IBgZ
3y1YoVu5bRJdanDju0u9XKtCTsEGYM+P5HNlM9dZG0dAXgsRxhzVgVWkydSW0PKiRsT9Xmf8cpqI
d/Go0ewo7r0t8um8KcmcG2Z9VBVWQ7UAuhk8w3nsVfJIdWfolfG53RGSS2WODSM1d6qRHC0+JY7o
zy5XDHmmnUczCiVQ7ZARkRh5OLoS2Xjhmvi603vijuAuN0cRQINM0krn3lv/Gj4BKD1xYGEj/Ftv
PJT1B2RuiFh/aHLY2C8Qly87D9zGxKQ5gWam8SsKcCF0865npIP2uHMd0k7HPGOwmn4UjV05sv59
xKxUJxBq9Oko6RgVhynHhLXTNH8t2lwXoTT7dn+1APd4Nvo5Yhd0BIX5a+Fts9iixjF8Sbb3NqjT
aJJsLt1y7gCyVx5/DTkO/9iI6Y09+XcZr2xwiDp4jorOYsCQxj0QkwyZmar+k3WmqZBAIoivBxn8
AsLFxAKCgxZpjklxDXK5zg3DIQCmCU++fPj7Sq+TC918yf/k8jWdV4wV/a7MYEuk8ddM8RR5Pe5R
7xviPdsZyoZJX8AHcYN99oEOZTIrc1cc64tAWKwsbZrOuXsYT5ANaP8AYz1IZFtcf4KAONmtE1dR
bA74udYwUjseWJVWtoAGaheo7q9ggoqnOGw6aqDFFtCki5JC84GjFEl7iv9JHMLSyYvMsXRODnq8
OZVZQSrMDUIquXURzv3lJfX9bWHilap9s21PCbdyA9ffYr/p6o6k3i9pz8SitN7y7qrUcYcSLIRr
79tYkZraj5Pu2+78JQdKr7GtuHBz0paTiH6ghom9piqMvXmkXzyPdPsN8NchP5dhrzOpGyF65M91
E2WuHNQb+jVwUZCs/EZnZ1TQglUOLmXtiA1YCr47R6EShMwb8tha+INj849BOnlkpnYupF+7O8wY
50pasL7PzEXTGbfyOqH3nLzRg/pgmmW25pzf5rnFV9qYZp9ko81OPBXWLozmyI5HHFoa2qzUbO5n
Yf/NVzds5N4Bo6L4Vdie5xT0PJZcsTrYIxUsp8OvYa5Pmkn7rF7xTSwK/6sB5557GnDwa6ZoyDti
EG5fYaee8vbarUP5jUn+5vf9oDXJpyn5GG4VAYI8464PJSXDBxPx+Mw5bE45QVXxnN1U7UqrkEAW
eok54jHxYsje5v4KKO8au2+4vreoaQwM0D/igogOOqPHEMFn0f7Lf9HtguDlfKiv0Ut4ozXsh7wc
wxToC7Zonjm/Xe4CJHxZiazemCEKCAjfjvx6gKbDQbD+ObAjMSux7E+7i7XxfWdpxP6rdP2dtEZO
+bJeqy/r0BvRvPcfoxjmFkhmaOSlJKNkyXWUezGebL7jvxcNX+6LDIy5ixog/5jQxok8ovChP4Xy
Hfp5Y93BML+X/KQVsFK9+rcB0eHZiskR17lxJrc57YH+DBTCsgtgpg7KsSoigbpL2r4/2j9LZFnu
WZ16kwmxMIywdjGubYFtWhZyvdI7uix9H6lNynYp2o7gAI5TaAmLbY6jB3kfeM5umJhZYBTtlajv
hp1plpyFGq67z364ozaJvFLfiJTTKgyVaCRjVl8QXbATA8YrOi1R6+rf1NjCKZrFcsU+ExJOl0LV
NH8H/rQbhOWCrhTkPT0vpCo8SXNWhT1L5Gzhsday4lczrKKmVUNjywKB9og2vkQXdJrI2jmxFT95
g/QyqWspQzVSy2dw5DOPzwWJcAoupRufkkdUFvJwTYOFGNrhAaBh9f2wQUrZVVddkYy2YVXFSWlJ
uspJKL1sdtPZcLw52KJkwQXzrk+ztIdpu75HlSBcpmpKLn3VytVbKi/lv4qggUIbwluYZyPPFM/h
IyAawW5gK9gsYDa/dNjFWp7dpAG8KsuLez0SNWIBa2lw//M8PXWTuxuqMiRTQ4u7RzcGzIMNWUj0
FW2cbZcBpTj1FRfJ+x55wtrJtPDyEZ+jzLxw5TXtCnjrTVxVOFU0AJT/To8GYIuAxDx2Cw+HNQqB
hDDKOpmz0e7LuFEttlY0HNGtdkFl6f1Ia2lHlT9Q/fa3u9k++ZFmEb+M0/DxCZnrSc3oMlSiutVX
2xQf6QqnRRXp3aqUZCKLJJK9ma7zeeXx7ju4Oj8tsm/Weeig/4QrsumbWfWJfeycmXrMy7mnfu0n
LvZYtBUks4wBVeJfDcStGMmtnz3l8hkCrbcfYRsrSqdbwmA4BYW56hVR3KzL80DQ9sspk9BenNdx
/2bDQBIxqra0DFn/cgXFZ3//bwmdM/wWPzfGXyf5WTUBhcpn1/XlTmMWGGya2HI3rQBw7tjiB80T
KP8dwB9o7SNXbxqsVS2PWM1IocqbtWh73wEONNzIazU6DRGyG+Gxdv7FIE6k0XU7bIc6fw/u4KRO
gD7V+tAIA6Su2v3mJ5C6y7mv9C/mL5WTHHVJD1jw6Lw1NOm2441eAHQACr/ZbsLlhAinlpI4yP2w
dcOb7Rcmugw/SXxYdheLkjp+M50HoJbLUA78hZaUc6Spf06TOXSHG7JYImID+BiUVrWrrnmh2AB5
vFaKkFr2im06JPTABFj8tSv/GBBBsZuZyrJXP3jEo5F/w/Ap/V2jEwIt2fgzQ580tF7SoUNxmqTY
jZQuLkWKcmTDekAe9wzJX401cktZzruEdJMxhOW8+U46f20LpazAFzGArs6hDfGdE6apEKz4P6lW
E/3NM/OzrMeeEwfkh68kH5jb3mKMPxPwrN/slUkMLSR1RH9TZF8cz1Hm21NrKYNcavR8+pmM4pBx
givhC0jle1rGfHcYaLohFTF5cLN4kXf3WBjO3PP4gQWpUGunzx7F5muWa4vDm5FVDwnIu0oqsV0g
Ftg7IGsKR2b0Kim4ZSrWN3TU+Tjp1/qSNaXLw+b2IBZBKI+WnsaLgvfGIumcZX6/NM/QKtqMWzcB
8/zBaLQ5pAMU20hTBgbduXDwpilsfwpSxjt3xTmtkWrhgsOe2UHPEKe2ia60aDRVudNTjTe64VXf
utuioJDfKi31+3fwlJdl/OPJWIv4Kmgrc7vkytAiybl4RzS3YqYX+l/sBjpwYlT+E5OmH6e86kYB
/qZ75XDDBi2sfZVMKq8WjamZdkFYzzgTWh2CHUwiaUHLXIXW+r69Pkw5R11J0vf9og6awCl5zdII
ZroWWFCCukjsdT9xiWWfHm0FhIvK4DhEHb1qOrEMg6+FpPN8EJNVB8os2eGtZbLYSPCA1NxHsNQH
WbL8UFwpsPp/W0DNdBXRQ4+Bdl18rmeaDbsqOCkx05tmEN80aEMD7+LdR2dNlTLja2EeGfiXB6Ag
xcKT6OSHLeCEPRjuy7CVfdi/LnXibZlZx9WYuXKy5+vGUE03eq0QtF5mlShsMoUVg8euW6cZ9BoX
fcH9A4ayzAMi+5R4ucud2HmIhUvVbJ8N+5cUy81PrVL9IH/dV9D7bOcibeg60PSP9i0g6N1DQ1mU
aTqty1UJKkXXmOCdvzEceSCSz9GE3GfEXMdlRwPmhX6XbLlJcgS19KJgjCri5ugojl2Uh/bvmMwp
cjscpUe8WltTF9ymx2NQMt0UZtuse6JL7M/sAjJLuLoNkIgyB8sf7ZCg14V15tWzUOhC3PBEKJAC
dx3axoaBolf3UikMTaAZOK2Inm8a/9gyohrTh6Wo1IYdUCbA5LswZr3VQt2Z8oQm4BaUe4RbTity
TNrt2HA4C6Hun5Q93ZbZtTF9/6q3xVD159qYaG0qqCWb9rdvi8vIdjUn5M6wtj0Jbwm9PQf8yzlB
MvwxcKfPkWTP7CNQCCGEfZTmoDZ5Gqy+zJo1h1b82QjCsa9hVcVrBJpMXZ0IOPAH3gpaB/qziwuJ
g1SBUtmntN6loWWUEkZ6z1oQ8oOpWs6FjnCF1ZCJZzqBXlD+CY/jhrspWfQWHPVS0QZBYXXUEv07
Uu+J+e27f6tIPyFt6ywsU0qTPZoozli5V0p3qQMYfQYnIGDNn+0bTsKDUnGY8YUTa+8WnB6QbVaz
AoGkQQLbdzG70z9vQ5TWTNaMWewSPO8uHFGU7Eg5CVSUYXQaCAkQm3idVNJ0rcAR1TZ4Mrih5vvQ
6h+4OYMuq2DWRJ8RTBbfFPEPCfWh60dBpUAf4xD22Bo0Rycop2oadXAQm/n1gxhQ1zW3Gee6rd3A
oYfkRu+P8zdm8XoTo08TCi5ROsoq7f77nwHdl8W20iuO1okXlk58/hUZGNXn3c8bD5HkF8lKx2vP
3gccBK5HOITFrRSMU9pM/qIr+cNmS2nQZUWXaZ5S5xtALrOy7GqE18iED4exntuUk0/W5TGvqpAn
R0fBpq/zqkEV4ffJpCh2VzfbPQf6ac2tnP4XdjXtyzsx7bAARcltvgzn1gFxscKQK7yqGarV8blt
7QTk5S3gps1zt87gavXKP0Z0VDV1vy0JgD17EhxbQw1deYcFnipyDRJJiKju0MHWQltSxrXaVtcf
HygkzGIjv6A2eWxrklHHmMJTdULg8x3MYiTKh4kcS/36NbVEaJJCSvkoWSAyYzSfzRqnwhFWYaT8
JPXsz3ozDB9jRn3tPtazw4DceTaihZXt5sIStvW0awqe5MY9cZ+FmG+ps+1IBgkQ4eU/xMwLEp/2
hYAxv2ESZmTAxINV4y4pC/jDvKtR2nivOIo2i0t7JqP6B283a4cid4Z1Gbu++oxFWsoLMrKyPFbh
KFff6QHBgeL4bRpSlFENv/e2ssTHh5+HGPJk4UEp9Vf16ZSAk5uLvwoGncuvbX7BWyI9w/k5hwYW
JOE9NrjMTwX6xQEnsRiNdsLdbugr4vDf6hs6tjrBn142jmRmuwFXXDSRD9krxWyzkdU+sIhnOaEa
B0TC8gFQ8AZW6bnOVMQCTBEwaUq6bKz9kyphkQytNSnPxTUzyn23mqV76/dmEJ5yO1pByKhjmI26
VGwYBz2OkZD+IRNgJGmNsNiiZ5z8bwkJWGFfPfxssfzyGiV75sIP0o5WIp9W2WhR9JWO3lrb/P+a
b931fXL3q8odJ3uV4laLXKtHlx/w5Vlynnq137fb8xt8x8pixOSfjUuRwbIfb/0DNuLcIclN6xrN
+tTnqWywETXtMwfZxQrGUVIhN0/0ThyZNhNcZEMvFy7OGU7J0Q014SkVpCgZzrG70LjjzmunN7Ou
StaOO+HAkweIPT9ll0VeAeP+HQV4tXwt8tgZz/v1AFcT9zxWPx8PPP0nf7g7gE9e2XLOgyNvAFC7
a0OZOV3kfnw4bRToBWSwP2VT/h0bF/VYvcMabiIuemf8LqPS3q/DbHnCYJamLz5gzTqftFUr87ES
2GZM0sR02n6A4w5eJ0HtckRHUy+c3mFuyjsphtGtTCsTPA67tIEExmyLhS5R4M2YevkinQYFpTHL
4zVgIdqtfDGdzc4EbfJ9cIedWPPnlqCuf4bFwq/FGBU0nOORU+SeQzJCO0mwZILSaXz5ctlE9fqj
QCGejbO5d8/qJ7xbrbePISxqcKv5GbubDfPfKFh82NGrnLwrlyRpoOJKwhuZX70n4KtVRxppKtts
uq3Vz1xAuk8JEqYnRVD8K1Sa1eoyjgnGCSPpQCySK2zy+BLEVWuKLVwzoqsU7quyCIlmpAS8mn3j
Csw89Vd88Rvmc2RaNCMFWogkBPBtCcHcBDiVXPK7Q+R9v//aSukqRLlECjb3sug3Jvx9XznKqMdt
J9AmsavaQ6dSr02O7XW7FAzEdqZ0pBpxbcAEuT1+pYe3jdl8IshZcQwiVd4PDX8Q+jRgkwbJhHzB
AC/ukUppL7S64OPBCu37VgkJ+K28lE7hvsZjm1D3Bl6H/UcuLzi7C7bR2pMv6TXs9pt9j0fj5uRc
6OMRXKsTNSvsoBI0Z2XRvppIQOzJc8z69yx7JCDWFhpnC49ejOyh8IjnZ8lvRjvdhFDl65/Ucw+v
NBjyAX69k4XlQ2cfhfZZtdkBEVkf1sD8IOBJE1HyVRLYJAi3YiekMIYNdg6ld+HOWOa/tbB7sHbe
3xJi4ec2/TnXaKmU2w2gA2IVTwx15EtFUZ7jTiC11bse+UztJQkzIrWpNKi49nX77Gggf25ruJPd
5RP5CZa3xpTr+m7YwF3Y3nn963IPMNScwJxx0K5uUe09cGxBELq/mImAshnjcDDqPx2A/MK4O/b2
hgvs0UM0DIR0+NHR9r5LA++lnds0AdU1oOSEl8gFGXzhCZ1AjXgBGWpISUx49a0D9taGcdOUbUt0
xv5HpQmRGSZORLHP/q4Uv0dlRx9V+ShhmhUap040CaQjtzznir41CuN2+/nDxydFYZvJcull1syM
4i7HtuuPdgc/hTrtZfoH9njNZdChhx3BVvX5wuyb6Cn7WLFyftX2lIYNqD+aOKQeUpM3qAT5TKjk
G4TYdP6IdFsPeDEL5rWRWuautPc+33tFA1eMW/3buN95fBDLGeoiVNbZYBIbGkh2SHbCCUpz2xlp
tnDvrPpm3ZO6oLMGP0CTQUh/bYQu9v+cP0mvrO872vmHG87yd4c5DM2fKyJbw18hPf/K3z3Y51W7
ciBLPkFKOxQB5CPFIHj5DnhbXZBJEzofhM2gvA3JTvEAE3OGPtkpkH7gRrrb7dO6Oj6fTgxsT6gV
hhCRCwPxf9g9ZytQHA/vOX4BkNk9DytSsQKE0cwdC9lqz1mMTlLCB4jcaJc9hEKnaiUmK/9/yzR7
rGLdOYuXdmGMYPhJm1Titq1Jtn0X5ZkndNvkSs6WJth4XceAqoUXdhJKlFI9tn1R2I2uUiv6pgpg
7IR7AtOQlDMcFUgQl364DHpM0V0rHwO7VpQLSmiLW2znL1blCYB5csHAIotbccKy1Q40LqRXPkld
oqlgP6jpWC3hWSaTyGHagdGkLx3FBphcRUhby7IzTj+A3ncghAzN7F3EjulnCtKHBE8aioNikDQn
3duI+/iAuhTO4OhOjWAeBOXdZhzAtrVl4qhUm/3gtIe/fAmL6ICHfM8Dzl2TXZtqavP0y/TcJcuw
SmxLmfDlQyxbJmKXle6yKToe2H9lmObUF6174BOldJjfXFgIIccD7qBChXb7c+2/4+gvtc2fzRyN
tsS4eR9Nk/AnBe5TiheJiyE7QW66YuWiWoZsHGF36UrAENDmObLip0iJydF/Wk69C1fT61YCyAok
BdOtVZq3bbuZC1g3jwKjoSBBnNoFhbouLUZptFsqq+BUon0MSAr6tJBzUC3qtXhHriNe5egNqzjZ
wqRyp9xlg7xIuslCMcCBOD6QOQyzuIj9hT0v8YSifbhfx0MhLPHrTRTvZpAcFRWHxQRBmu+AXyAc
87F5D3Ppbmifz7gl03He+kWsof01G1hm9Py0YhWNQAXOX0EPE7qPrLNqfp8hDzy7dbAPf7CW3fWw
rOcrzpKn//rAaU84F2S5b365T0pwJ31citSP9KrxQxEpVVSqY4u/kWBfyy6ACDDEO4sXV6fzz7EV
s8emmtiz87UtroUvNXVJX4IaSJNTAgSvnTRYkOFxlb10EBeTgVb4OB1lS7o6dhXZejU4IPy9lJ40
omuwd2Zt5RkZC+cf+Rj5Qyl98tTC6mn+nutV+9MjRmRif0f7X7SVDuhVikB14ALpGhDpCIk1EHjs
NOEQORu7cwripG++5NuVyKu2AYR/UxszFAESLjn2jsVlpT932zuV1u6aTpqkQb0AKZyPzjg6j2Rb
TvOgEp9tMq0dTWnFVNy1bREUy2iDCaw52PL3bXcMO6WiXR9h+M8bn6X1tSQ5bA83TIiqNaCrvEw1
dj1404P76IeoxdcDcTVTmKQ/cwqNDQn/XZYRTyz1jSvrfwWOyBdI9tu+plOZdzwy2IDmMFbPycZ4
ETJPgA+bTi9hDN+AmT+69v6IQUwCY9SIoI4YAuLF99P0/Fx1/koRtaZ/B7DWokQfHsMxVNbpjQ5d
SCS21lDS/gKtRtCggBMkUtuW5zdsnwP3nu4ejdRaYhzFCW/gKqEqIWYFbCCGpZ4rxRBMdKExH3Ca
vo0wBG7gBgpjZ8ewyscLVNJoSlbujrFiXSkV3AWpxZTgAt9sWFhaZ8qodPWj6PNsefhbk5xcKN1j
zjIKUKgBx43CFGjTp827FWaSuErOC2XEAD/xDvs0mXFp5Qz1Rhmm02wVhtf6e4oH0DH9Xu4SDRzJ
jCZ7uHy4mh+8896sXp1wR1uqt1vMnMfFde2ReS1okNX8/wBeYTDZI+2UVxfBKy33DnuaDXtEfeIr
+4LkJIplA159bh3agIwKjSXmNkspwtiSBd/F6vj5HIQrc7iwS5flV3Hw4YsMEN1izuCWIQ8eVPtP
RmWxWpFt1cCzcH1afKWg2hx9IbIy9XyTl86gIcnbItSPMWNa1aTR74gAYqxgauqKeyzRzi6zU+Dr
VwsyX+euxkcf+D803zc8pr3nig/PztsFsoZlSE+kO/jK49WXc5KP2yEFfpv55Ss9JvDs1KwZ7SYV
wmwaNgEmMgV4i8+gP7z2WXpQiB7GYFNr16p/+6bI5gGEnZcpzI8qLtkt76j+Rb6mmnDaosjMzYDv
ss0mH2BEh47IJOAfwmhRM/ZdblZQfEKHCACTh00M1qBgBEqmjrkKz0EJyC/PWMN8DJW2pRyZNI5M
qHX5DgP9/y0YaJjPOuk24mePuzxzLIwd5EGH4Kt393uyP13G/a4nvNXh1BTyxxRSCwCiqhzUkcl5
Eh5res7gnzeeCan1WRqrpiTd15usGYnASXkhyaednd3+YvG2dWZS6GHM4X7UlAQrUEhvF2zqSNml
RNBUTTYhuJ9iRkdbcybZd3tyloX50G31akaqL2UFPjM4mWgK4koisEzsNeqYaUPTZWemHzW7a5ZP
KtZjdSevLG3mLC/87LUkyJjuMhcMJSyOlw/IJxYhpvbfiJIHM+OwjGwI+Y549PweWmKBQhCWmeZF
lh5od2JgWYsOD/AHVPnZVrBPj2XKuw+5mK43PHegMOj3TySr6qgBmInP7rFUffUAYZILSgK+i7Rs
dxCDUQcRIIRB8TvWsy32W8ZFnJ+MYTPB7JvojayKhh0qcuhlRgyz2QqiBUfmY6MfdeUGL7+IZTgG
gCh6OH5RFFO5MkUI5uR2v7jOz4oOHKKap202LDKfhL0/fO4rGFIwOK2pA8Rsv28m5dqmNiKtnvLR
ZaL7j+PeGmle7K3Mjx48iaQWr4Dq7DTBlK7ltqQCSG1ogGUGWDih6y7Cz3iKxx+DH7ct55kuz60M
u6mDEGBfFWF7MgZAvjkhVCoh5ls2VpPJNybwSebM5AJLwCPCMC5n5y7be5rzWq1thewgGL8tfVz2
HcIqWHdKjJbRky1htJG8uOYp8mXtLI1OHV326VdDNLLGPc9pqIEeDBqZz+EitBgIZ692WE51ouv5
g7txJEsEyo5AdRg13A9u+HYBH7rawwyEeNRhKG2mqnUQlID7mcXSZGZ2MSQ7MFD1VP2IMmuw40uU
q9guldEjSgjTx0bVMWjQRH0p+CFe99xyt9Q5D+4RKCMfATzAQ6u3cr2hvsMR4S0XEJXUtFtObAzg
nQ47weN92c3zQwk2B0Cik9WHuQ81ujBY7vpu0t8aVTbQw6KtxyqT5wLEUhBEU6PH782O6V1TdhkW
OytpE9v1k2IoCSzqWTIfk+QAhEPhnta/dvNt7378qwi8Ch5Q8RIty09I/Bm4AJHQQ5XtsGLxN74F
giPkdtrTxZvfdaDTN/Bd16YMsVaRCSRa6BtU1bqGOPUI+4qR5oKTVwCQORMYk7Oh65QqEXdrzZjd
u/EBVK6L0w8GfVz8GhVffKrUzTqyh144PV+KLyuxdniGm1ZJ2+j/ibEidmbsCWK23ROgZx6ixazB
nRMfmQNuM9/DDILlMikgWyRgxnxFq8KptR/XzL63G/iJEH9aMhAQxvHCYER6DewB7h9pG+yG5HiC
8svszLBgJBOQNGxmv3Ygw7K/lmW+7Kwf3iWrx4EjT6p9C8P533UNVNbKWIm27Jxv5czWMLXf00wS
gRrtEVyAEPDFE1BReHZsarHlcBhuJCb6NgyfeUPkMFjya4Gs0n01z4xxUpPWMG6kRAuLHXS0/TXM
/ZJX0yFkvzpXbSv4mHhNIgAftCtEi3troGzHMuaGD0udkGtyZ6nRfWy/V/OZrOJs084EBgdKwaHQ
C97OEgDuSZinuP9mWR3wEy+37Fsvxe5+6OZkTCkbthpKOj+w7pqVz9F1coKJZyQWmYsDce4dvID8
S1YcDLZ7qbBDicoCyMhuTxi6tpni5WfirFBtXKfDm53HKjvFt5cLwhzWxBty7yI5EVnwWkA9BO6V
T77dgXUT4mDTZDZ4bknnzDwEXeYQ3M4MEKlIwGOi671AsdUsHxEsZriyzhJSQ9xg2PgYlNbVgZIp
/zze+XTcoTKrmbMPMl/Q20Y4vb3wYXzD91EvRe8FO419bErBBCwrJKyztHSYzZ9N23Gzai8IAFUA
9rEvllpm4bGfQcBKaWe5SRwgzPKewwGBiuek99ROt27puBGr+ej3V7/abf30ybGo8gdJYx9UG0O2
pXz69ECJpBPfCzhJTuBQqQHEc0aW4Jrwk6HEsfDNJuFKOj/UWYKDhrOsjSooI+Zi/4DM+2M5VLlA
z4SofZZIMWn6NUVUMKOx0zZK9Y9A+4SGk1pu1MI47TdUTcy1Ui1NSeq9eagLKeh6mMHMVdBuKCkB
EV1S5Sa84/fBLs3cJ32NNBZ0PNJy+oofn2UarWpTxV+XoGalUyut7TTRcnwKu2xk3634QglqLLS0
pD+uxdbY3RIDpZ2BrfEgnhnyYal8iqH2YB9//x/UQ1IXMToVItzRCf4tREgQsI2lH5CjuV7SAhtx
wignwDWIUCKiKKO8XUPRq2hDwdiJPXu9epEOAf+9Kvta1pk22Vr8RwQjMb5euhkk/jsAoTC1mY4+
Svu9I0EaIdunE35fbE5YAQ+NGSi2GA0H2OHlbu3Jy1AZ6mc9saWZWwkovvvr3vZ3ntsdYcdGYjV4
PEvrc5DxyrYkuDlrFhgYAfubxPRi1Ry4o82oU5EwW35ywuY77Fsbhk4L2CGP3Mo+kOF1CXU8kVDI
RltE/4kSpvslvg7QAx46STUE1O6vQReXxeUkLpCKLPFV4K6hywcWiuQNc2qNBQ+4iEsZXNHzr+7l
rfDXpzZ3NmYC6w9JXcHrHoVcbb3Hzm9P60367Aj7OpK0UHihIeVmUdtZNrR7xlrzYWnctp7o1erW
yTgSQp29Q/qGSkBsZEXacUdFs8VrqENvhOwsyFBIo5MWAmbNHLKkVGEl5yTjD6q7DSIC3Rt6WVs/
wGXdKaUxUyJO+t6Os9aa72TOdQ+tvwcq87VG6ROU24qsoctBp6ysKpcASk4wWRnNclzA/7/t6GTI
aWH9d6F8w5z1P8se2bUXx0TU34G+OtSO/mPXkcD6GW+oWS3cMkuAGOb+9nCQrfvOeit7HtNK9k0N
MnZ8eHu67oGgbWCko24xnCkzZNYQsLfEDqzM+g/x8rWcjzx9IKvR/zXaXb8ieI83O8H/HimTDw/W
1pJNrfNnEG2lKaQwQXQ5PAhebmORPq5+Qw98kUxbcEFoUJJS8eQEGJPOeYJWuslDZ6eRkC2vBqgI
BSU8YirWqq5oYmhCSaw6RFBQwb556Ltj/AMhRmraMF/l56zN1Mzt37zoL63V3dl4MlLXGSzL5iPD
+hV8JX6a6g17EgHv3nscOQBsaYZ1c7IOWgapsSVsA3jywjRI+s7TP7XOSxhC+cN8vM0qDtZa5wuR
Q7UGlH9h4/755nkeclP4ZIMThFOb3dOXEsjaEsbnBKuOwrGPhCA4hfXsAkJReugvETJGD5tcOahI
OANrVfXR1xh5BKXNTq1vToSqjny20oYuPqVsJrQSzX0DAxmMhA+zm1fw50kjL0R7qSYiWWJjJBkE
gTv44vNH7F/JSIflcPlMaMGy3f1ZmTNZfyK+HR0QdykuD3n3dor9po/hPyGTvQXyfTkPXjgVl/v6
i6OmvHoOeZkEl+ktqlQSP8iZghJtUF9+6dxsgynNtyo/vu7A8t+yQZNpaNF8yfbPpvOFeh8N+kz5
h1cF5kZZ61xXTggmylbl/tpYFk7mvKaO+D4R74DTgfanM+Y4bKT4e98EfFCCE1U5x483dSL9g1/d
n8KCWBe9ERzes9EiFACth3XeB3B1O7f783lzTx0wYiYyHkhTCX4hKFjdMHghpTm3lvUXrg7eS6Hf
r9EbY1Ie5AjyXqVYl781FlYTfyMBuZn1r5oJwTgg+f7WG2qg5JdOeya6DjHeSp+gi3CAZ+w867xq
JEnI/SoS96ToZMGEhsz4n6YfMxWUqfhnJUL0eUnK8jeTQ2VdZJebH+AG3DUcMHLF41oOULeUbtnO
AXd1dNrEj9/IzLYmL3bI5grKM6FhT2bLLIrASCi0epGqX4wF04oQiom7dzanxVy4NwOBk122H0cY
MIVKQb5W5AXm8BTS5pLDhyjBIR33vWjXsDheDdkNem5+QBzlgoejKxYD5W2lBiDWfGwBvo5gNqcv
rNeay7hFMunVOpDAi/WKrYrqjgh6uklL+Iqy3FP0PZ3jxZ+KD7NdcH1BeA0/KWgBM2M13RZtKBAA
0eZF9lIqqxheuZGFKpSmmsMbj9zgX/P9AOkyp0u1fd2uA4wsRioC3AF+ZNKQ8mktbsoCOtmHObWv
q2ss8K9B0tZmz6sRtNGdOlBLFPoV+KhT3BG2yXOsllH/B7iufJGUySMFHvrP3zGCRQrmI6yix4Ly
wgSZZNriunyQvpD2DRynRaxTZyGULS0UBzTqLqrk1wtdZgrp9NR05gi1aOXmOJbhFyzdO4Stfa7Q
NiaQJYuJvCf4abuccL/yWA5R3arBird6yjaintz+/AEJ7gdcw1jbPyLO3B6eDLhY6u8w2DOIfgUq
N+wDo74grlTiCKyWokXwOK2jJXV9AZ8Pyt64Ly18aN5IwY5yAwe0fkvtGmz39ac34DTUv3CJkxW4
CYYqqP2PahR0sb46HmRGaue2OZkuchst+oIpunzDzLNBRCOL+QMloP054OnbUraKxskRCqiJtDUL
IGYIQHVF+XHtX1GYPdN056y87qPlWKW+62EyYwLoY6IYu/y7biDlQPqv76GAvMty4iz8HpYdyyg8
StsK2INtDyX/pCJEs8+Jh3pVBxQNnvasK4FUjWaRffxyo3Zzuw3VQ2t5imJsbMYp81wmFAidgwjD
mQGTJtc0YJpsTy5X9J9p1GCXn8YBdbEgB5zF9mShTMuvgFlMY9rMqflnCSW1twHdwi81dGA2cEf4
YV5cO5CsAhOGwhu3GQVFBjKk3Uh7wLpOEUjUWFio8gzPjmipPwUKsPHymwm6X4+MGD8gBSRFvvPW
9iW9tFfTNfYnY5BhPLZQdhDhRuARxrwyyi0jCQB8q/Iw400VYm1p9Puiq+i3Yb/ptb81MnYQJ+OX
2FHXCkpa2bJr+UnzUyb7BSJwc+xV9APF2Lh2grp8LVCtq1zUXSkpxM9RJ497pvVWdtBAd0mPeXoH
Vz0+WPsfITf0GLjZAWgcUurdGDkHdoNMjcPpwWKrZGlMA02QOHmnoDzBlHOXyhZlmZs8Wx1ZAjaw
9JnX1OWM2QigIXwSAogVctVb8YarnRy5ZBRmeJDsKxkawwAUU2AD/CvTSOXBshPPfbin4BnY1P/D
DXEmEOGj1bTK9OgdICZgJ+FTq79PrZLWU5Ks1ZkKSx+I7EZ9eBgNWpSydKXM9HN6haPwu8mMf6vc
1dqn+XBa/Ip7CY4r0ZABYRSHtGGhjouFrDwJG+KRa40GMXEqyg4FrZx8RsTFtrbb/ucweyBPyPvd
Z+g0zJcx8dNJoGtrugmuJqcEwkC8w93fElBJd7vumdyQ+UFli2YQq5m18VFrpgRXENMgP9vEw4Cy
J/QfpblMSJYwUALxQmzRaqDgmhXbvgApKIR3RrYYqMt5iXdUwoM/MrRCRgw6ZXRTbBT4EeSk9Tqb
GIvfSx128EsVx1jv+TjXL5okmxV3zZ/mH4twYpM7V4uyAkRedXfdDorC38Rnfw9QszPiaC4o/ffS
wUsMdkhocuPJRT6A4Z57k/5KqJQhrbGjcJn7/UptHOJhRVOKDUPEhByme2U2jSlXnkSjGXc5uXJJ
HkXsrOBdYinEGfGPLk75Houe4CX3JPNjV19mxzHDYl6ZBxkQt/kz4Rx9/QvnZ1MSw3R2JKc/9Z8d
h6+gmcoSbnzRaxaUTgRa+Y/aL6W+maqqa+bcWuyvyvWXxnBA55nqKp2XYZxhfwWBOcpVewlTI/m6
KaDqqb6Z9etc5Xu7LF+pG/jWnZvtnRADjOqnPsMr4PMfD/ZtbVxEpJSYQcmuemkobwaeFdDEOaSM
eOqxCY5I87gsLvpZ9ocwZ3o+VfHIusQxQvvLInJLJ4z4RbNa0X9bwg4Wqu87MFajt+33yMdpOX54
Gf4IpxcdCPm0KDVeh4DDnR2f3dsenr+EF9j1/AUXhl4HJmBbCPoVSaiKrAH7Hjv8XFvNDw+uNgtz
lm9ldF4HC5JHGcI/gWUcsctciahftZaQMpSOKI7gsqLyLVm5o1rGZieRE0QPgQyfYutdAwB7YLWq
e0oxiT6lIhbO/2juXKPVtdaLD4Zn71FN+aOV+SB4AW9igeDhd7NFezdDw31gLDSc+6N6hl7uQfmT
5G7GIplUqXa1Ry8yqsaomrJeLDpSxLC5vLZvcjjVEOrF6VgzRwulgcZAUbvIaE5bg4uWqs7zv9TB
Csa2Btg0O1CwwvNGYPgDRYs5Y4ZNQhYmXugjuG4sKXT5B6snYKuy31uW3ZA5Vux15dO+be2SWDN5
PJPnG18ZpZHXozcxEatWbAHYQVreqBPP7TvC1TgIHy4Lq9MmGDvOw+L3Ol1gYFhcMZnFsa8JT5SO
Y75QMyRr64f+TlQ3w3CEZof8B9Oe3viBPlc4YeA9LnpK0MYRCJHN2KdQcRk8P/TNdtN2YdItqyXj
caZQ8OVVli+v5Cn0KKTSb/kbqS9dRh0xkuHiQ8RVFIKKpwWA512sSrI4oIXsk8G32/h2hhPHjr37
UDeSnSamf04WflQKfzifcdZ6PWtdUnDh09dpPkTdPxfQFCsTAyX1Ha0fqpKZY+gr/+u3Aj+PRtAt
PHowVvQtJn5qImZYe31AxhV68Z87ATItruU/5LSUieZ1sjGmypySIgEH/EpG89YDQzHX3Ir6kcM9
LF0GCBV5dHZtctvKBsT1oYvIiYGaad4pZEO7dXRh+Q5Vz8ngSHA/YUdgRQmHHUB5GJ4WDeD35jDx
MRMYU04R8NADnz/zh3GF5Bv6UlLc2otZ5R+nS5FCZh3ZwIzuOx78CakmguqaSYNlabMuDtxuHdFY
/2gckRk3g13N/LR43fWkR7fEbW4ds5J4V1fGkOjZ2IsB5+btHa+5j5anbuJiKmkUbyW8242uL0bL
TGccALqLrJkG0MG8dDDcoFB5Cxp0ef1pyetNis2I9aPfLmVRtdtvU3HVaA9eW3U/stVl5J79kxHC
rtpEPj9T+rCG9+KKEULQRY6zwES2Y6qWab6jx7GRz3UC36z0uyTxCU4BV9g0nDmaipFoDf6qKHXU
Z2rANkocBc23U3UklxWJovBHzNwIywsqO6+pbLSYvzDhg+UU3WVW9Qs+cJOEv6VG1QGMKjzBmV5t
qXlEqon/5a0wHeTEz1NTMzid06Gjt/2rhWedUMM0ruuqGmEp6u3mrKozfM2yvtnJ4o5oP3uRtUTR
jMwhiaBF/c9lXWzKRfirTAMlQr8vQZodwHJE4++U0XxeE7jnySWmiaggf5OkOJVkb8hxn1ta5ltw
L3hVEz2QoHpXQKoSDQlnmtxgkQo4Gc0NQ8oWalCMG4jd7Wh2N1NWA9d9/2nTLn7QQ9HLPEXjSaHu
yOzmxXGmMreuAfvK8xOzgltFbV1OuB07opTtWCy+nXU5Zf/HZYiPVO5me9iTofKAGHnCs+BGgQ9w
eXp2EA5IWWxIK2tOHR2th38X4U6g058Kohqj68JRV/y56voD3xQeQsUdO7Zi6i8vPneYWEek1Zoj
cylM5mkunfv7KLaRouCGJrMgM2gqh1H6jKG9IbwKx3JY7afdzE0AMRxq3fZvo6qHMcYfux20rm1n
y7fD4VU/cTCAY6RUdZbaJORRTFyN5+aCfMHOlZG5yP/me2iu9cZmSZPfg7XQbPlaTEWqdOEq1tt5
CdWgBWnos5QWh89XDmBGQCKo/u+p5bPHyYUAbN99kjMerpIwjoI38Tgcbfw/IipAfp86QNTu1FHC
QbqYn7RMVXIKP8tRYbJoGoiW5kwAa4moImAp1tgA5oSTFhQ+uNpi2Nq+fjIRN7zKUlakZRGl6+RA
I90xZQcYvQ9gB8a+IMmyKAyZCTAe2ldskaXE+GqrM2EefdINXpjghVWzKpJUcbg8nf0NdJs590i5
KhW47q6DGo1xBwYDkp+gUZT7lTsKif1M6SB0m0a430kBkUSxyaoIKg1VvWGdtZ+uqHrNIB5MELfO
zTyRnWLcnWfmkL4ZyuGIYcpWWDylwanVZKIp529DF07eEDXX7VDG1jyyeug2Sq60o98UBgVCsoYH
VMjR1WA8EbbSKHhjbfk60vJDdKeDfPM8vO+Do7hHQLUMx+/2NGqBpZUyIPrph4otPlg4yHAHFvyv
xTPkc3OrY+z4aszTvIIuABslBtuLstN23s3JZSwPjOLoveVmq9eNqSBBQXsVMl8J4GcP2OEz6Z3o
KaK+NjtdD8/oOZU5MzNdlcJcOCT3t/yyxs4yhH7JV9lDyaT0uDVmqLNAT4PAeVPS96ITPuHz/UBR
ptwDkP8CsPbBNeLoSUXPSgIgJdoewzFqWqO2uS0eV/ChB9PkXbjowV1R/cG2vkRY2Cvpg1YyKxKE
2qUdZoTx1Wz0648YrZjWnSsep0XNiTFQqqnFirBAx9rXZ42nII3a0lXXjrbqrQSpHklmF7Q0pp9v
8mULG0rMm6D/cYDSl6BBWc2HLd1gqkK1E5055ujfq+5f5AgNhNbcKH5//e4e7+nzTa2SShUXZ+1r
0IQ4xYXL15Fxo7JIKa31wc4r5PqUsgSoD1mERVMQpTxv3DPtvNsRL8n4n3ox9Cru/l0xz5I3WSTN
MMgk1qhwV9e1NzoGic5oQKhKnU6q+LAoVE9TYSVd6Dt7et53HFM5RnhuSm45K2OwFBzE53g0c207
9ub3v8ownZfZsEE56KKpsbIQq3BjrRxstNicaybiyLeiY9jCnYyejHdcwksTIzFfJNTVLMCOCTeA
TIQDoprgGT6GGMBvtbz9fzXyRhDJeD7iVbsjZE+DAYfVZiCX0YKWERnhPi0RulfyHx/G9IgdVQAZ
5j7GEqSvPJbxS943gKgLhcL5Q75c3R1vKiXqVTYMPAL2Oy8WyvjpKNo3xfqN8CY2qRVveWFxaWDp
pYwB6XDQT66wmii1GQvPWQqPKXa7EE+VVUGwhgrkUnRxK6xDCp3EGMH+YqJe2jdP5hmO8F8vPOo5
PGZSae8A8NMkTW0JENBW7OHYXZIZYGV4HRaVbVrL4XlfxYDgGCjQE7QIikpE7ShLMN28BxBb1BKm
5WnWfp0Fh5zqKmk23AfMusNYcm8qLLilgw3prZ92kaTTD7sjhx7r+Yjp9Wz2Ap1/FFx/djcJjdJg
dpUksDj8VUgh2HBXB0INnd1oKLepUpPM1mkbG2z8arfJj6HklIA6v+A0ngI5B7l4QHbjMH0a3cpm
7n9Bi8NXwXr7hR3tqG7yRGaxCeOTTicoKG8uZ7tnRif17Y13tnvWaV/ScjNXQP/xwcxkng4MGwaM
VYeMEpMbsBMqeJi1Ewom2XDVOy10syBfla8knI/YrCPhGSC3H6tSDXh+RZImypf9+hvKIP6/l03M
0LkZ5sTuDUft9FWCQnoaD+MOjD3QnCdqW0/ZIfB5PeWTWMxRd3l1SlZjFy8m++5gBKma3EPmxs/X
vls+Kt0VstK8WWq4RokW1mfgeYs3Deet4B9fXDvbpnThnCl13M3RpOtJkLxVSnYPGreiDVlueIF1
FyZ1cB3JTAtofumEO56uL9i3jRK+UMXlWqtvT5daJomgC5V5ld0OmeZi3ZJFsrWp9mgnlWCvW6JZ
rTI+qubduXFX0+AKxadvDarkcCSB+HsYo5y3YM5tqZ2TOqNJbwnLfjeiwx13Dy0zOjC1kz7cU4fK
Yu+iLCL6H8SiqpZ4YnWnx2TatIoUs8LKOtkBb0ftVXLm4++gFb5jPOq3mDiWjplo/VFTy0l7jI2r
AenkZfp/zSBktloic75gXmH3FfTxfm82U1fs/tTIlvOIXoAsA+rV+ZEtFcXN+JhWoojudw4lrlSA
y8JV6jsCwBJrAa/5JvZTtzLq2Sjjcy10wWkkm/XBEHXjjRkbKU6XEbJHBjm4M4H0BRL5N7mHACZY
QyDsnqwTfxNvE5YcUWDkAB0YtutBw9UI8XRercgTaqJPWlCjI6qz8ZK/3TmCoAPwpaqJ7o2p0gJ2
0bXb2ohvVihe3P8+ycs313PLrvPJFQrg1T4xPnlBNeTJBYFTD78PoAdm7iHGHmWhly+Jam2VZcsq
WH/Xzih/h/rCY/eeaD6lKnPPEkLrowUykwz6TeZM1V3BmoZEAuUGiY+hNqUja+63jOsUMBELq5tV
GNXfGVniCZfeviD+83GCfwMd648IenIZKRjZp8rXO/cf+D1W23M6blv8uk4E8iIZtkESwUZHhYyL
DyKCNSnq5d7mwsP4VlHhJ5AqEn04gosUq2VvNGPblo4kxav+GmmWd3upnJNxn7/Qze39ogEK2HMI
MEuvci2eXbmrwIiMWxqazwJCGtO+yUBPsfglXD+04nd7LfUejsufKFoYhoqFcz2r8azHGL0aGzbw
vmHMhfiDvq+tL5VL7Hu1zaqYN/jSzRJfQltn+eoJes1n20pgypBs5fnaq5HCLqFohT2+gWAeMktU
vBOl85pg0vjyZTbvJpaYUm/WsRLpGUHFghD+4o8HxMUN1SoRwTBIsxAr4QVHs28c+1ddYWINpm5I
7amKeL4GcXTe8omoKoEaTIqgx5bYExkMCfpmMSaueBgcLq4H55q1t2P4gULky0iXyeJzgyw0EpyI
lT+e01Wq3oqm3pXlLE5KpIkPfxX/Oj7XUE4Gf5IdaBi5zQhO5FHsU36nQNrEsi72a1wQkwAxUY14
pp7y1xhNuv8Q+BPcMErb7wlDXGvOtjhviGBlXOgdhD3wbFeFWFHwtvOUtnr1aYIIh6T7wEyL1Ij9
2jHzGNzec9OcW1v6SMsnno5l9VljgF0DLxV6jaLsqCpvMbwMcULjpLxG5WvamUnvmSDAv7qY/y5z
ixy/t1E5TSTrAZ6uP2Vy0CgO+LYPucE1m1ilHt5RjaJFiYJnfTa2injP9RRiU5AlexiHJxaERA/z
xer5Cb42c3SNTKIThpAamZ80rDnxIAltO9MPur3Dgib42v9KwQc3cC7wDOozaAowQIFSR5b7W+ID
TfYiJa0yRaLqw7351rvt7B/z6BM5KaTLEjVSbYCPVQvgcYP03ZIdYV2Y9EXHoL5OCn5oLs++oNAp
pMSuXQxtVBAVz13kzqNLQYjpYlSHROUbTgIfAMdUzSTr0UoupKt55JSuwA1G5vTKmYJA4OhzUqnr
RN1YVXbj9V5T4lO0hbBmQUrHMvr8cPAouG8ljgbCkd6GazI4m2vgl5vT7Koa2C5rxP/WwaLyl01F
RYcMxrajmsMwOIcGrkiNUvZcAQzgSTYmuQFLX326OqtjPaZ+rfofDdoJhh2V5AS+RiI4dj366/72
yYispCwUps9+YE5ypV4mH3H5bwH9ZMgmRdOyuT6L7+DQdu978hgopNz0H/LaA1taX+9D+oB7Ub1O
bOFvKPUv1TtrY/L0HxKU/RlC09UWkiE/1/Qyz3HWGV6RBeRPJwte5prw682NOQuhuDjiB2ZN73p7
q/h0I66iUElMkZigGNjI7nuxA3RFmexnSA9o2MgoUkPTcvq+MXj6acszqEsB8LJt2Kk0TT8sxmaT
UvlpV8p9QqCEmYfn8qjyDAxRZlJMAM4VMELltuJf601jIBu8cxiJod5zEVLllW8OprWZXdEFWs6t
KYAe43pYjVjVHQgia27xDQaJUe8syN263UWu9K7cn0YL0xqUudYRS2No47Kw5TUUJYDlhEnlmzvP
ervd1GPVr8hKN5byGM3cp+HqHLMo6WjKiCHUslgv78TCZpf5c53fg5M4z3gt42mZ1cfRLTykMfIK
Qni5xlyKJLDBtDb8U4NvbrC++cAN014dYkU8Zi/l9vP6mXl+X72Mc8PL9wumS+UmoEyGfq4JKZzd
xmbLyo2EcFT8d/g3kEKVxe8qbgIvtJNPY6qnlOU4FEi7wR9bfUVS2HWJ8gZADYtFrR2LDGsdvMn3
2DxKURMW7tF9SZ3lInPHYl5EWvY671gxlxyZuczumLuH7fCVE91hFtrJBS6ZgqAUTnhBSpkf4dgx
bW/Rh9h0YFaBGOUEt+K5JI2/5kZ8NQQpqXVfXmVwchxEcojYsZzNaNewFIheQHs1ECNpF0KfJsIc
VRtLGLK6pbHK+pVWH4Z8k1pbKDoMZaSgLthQLgUimTiMvDWkn4VVwtAElAHz4EcJnSrxuXvc0hIl
DcVf/Ig5Wufwd9lHVY6a+RT/W0ZNNClE04DT7sLd2E7X8AgS2P5G4BO6/YHT4rKEdaSAiz8SKb6C
VdzPgmOKdfxW+9lPVFwnfnpWSzJ2aLseamaz+xc7wOIizzHDKZZCerxp72o+Dvh9jd5Gtmu3wCEp
svT6DalZfindsxPs+yXtYTvSDX/iB9VfKUZYblpNG+3fV85y1YqliMAUh8gv3yV6r0DKX7yfUIVx
Zc9Q36bPim7aLuweWnEectocg8icLGWRfseU8g6AaZI30vxj5bcILRuLgx3MnhvPmx1XcTNGZYXN
FcAGfJ3+4/VT7qWY0aAmH/p2vpS86fEIDAw1Ko1Z9KudvbSIo86/h+dtejzKjUtS6j0oFg/yakSa
mJ8aO8BoN92cBlysGOgHHSJCEcboR1afa7FLHLu8M2wKpAYaFpxNmbidw0G1ydtDV+hXmQQ++9a8
zIugw8of+k8iGPrIE+jwwKAuZnqJN8UV8yzx3F2OOKklOnzFqGfzpr+eSjwEJxnI5CNWE4xkn04s
hPcWVD67awQth3hRP/wjESqDhqX52sgkSOojN1G99qQWh78D3YNOKT68aRgOciWrBl8j7EhWjbWY
MZwriDEoDeXNzUJ5EMTmCIaD5CTT03CUj+Lzx60PPdHH6VG7jZPA6o5trJuz3Od4tiL1KjB6enGc
m3A+SpbuoL8JWWiqnOPiVktdRZLcDb4dZJgBT2CYNWM2D8K6aiN+aUHj5PZzaG+HIEh63jWCJO/+
W1+1tZOfErGpAuCkGlSW+7DaGqDT924jvBb1o/qStwTgMcwj/J4QS7dkg97cmptmFSvx1V6Z7ehu
eR+C/D5jdxPEVwHzFWnfKwDnTHJz2f4KUFBu7hCEkDhEFs+EwgpQyx7AvqlfhMY5PYpyp02URMm+
/DMbPQ6bKY1WKxfwK7Jc16QI+q2iPEyTLnq2M0XSfkyY0774Q3y8mlqRhMLEe46awebNjOsjZ/oc
/hnn410W/sqP+O0G6tkza7hgX6Hdok57gw4VxCkR+pWlLs1fCAZU0CHajEsuLOHnfgxKRmJwgbm5
ZPkWT7/4ettUGPSceGDEE02Uvz0KHqYOT8ok1Ii6cNIJISo6QQIVFhXy9idqi76NfLzV2Cinl38D
W0lzlX6hadZ3tBiwT/X80MTIIbNjf+dvD3LW1jzgEEEi1xjksmyzHohz8GetjZpCj4UVkbuwbzWs
qAhfijpPQFuL9LRj2igbOsKEnBM1Vo9uZQ0g+tWViefzjIfE4OvurcrbVKCEVPQPCnJgpitfEhjP
J40iFnRCUXY89ri4VZ+1htDnYq9ww7TufaknEuKOXL5lUh1HIVWqAqi0UElmi0ZCajxxb/dvdfd+
22PWPt5hFqRAg92c/jNjg4R+5FA44G+6GcyzhzADEA89bq5sFgo+1O6C/fzUmddorVYMiCsJpGwN
rrI5dplxbfEi50E4ENTTEUL6ajgsrhXTCLMBO2XEPkmF6aMb30DyPf9yy8MZZcpaub25pbwMaxdH
Y0jeXNGlAzIgYF8xNSAM+BBws31G2i/pVNoMeMA9okPluDEnR4FAizAvvy4MPP3NQyiU6W1kGft/
kXDnWTjtGH+eVZiAVG7YXK1cfNA+TfzdbuyJaU4PZ2I5dvTungUBLCgvwdYnlv42cIW2FWr9B1mG
r/x53ad0Egz17QlLshpRw/rM8CkKOcwyy5MhZzJzAJ3eoq9BYpMK+FaP42VS1CzgpvxDuWMHbOg5
fpu99vLJYchVAFbDDJXkDb8/Xlq9wlko+km79EZ/NxdWimPjXT56dWJnlZkyP1oqGyUZRbeDv3OB
cV2CNxK7+tjLzHJVA0jLJ75DavRfmVHUORgdIQqsMF8cw2OYBuuvUbiVlb5ohkFoZdLlVOMPTf+i
5TjT1ESsDNlyH6X4V6lahI5N671QP+SLvZsIfK6Pvss56dIbUbUKg2sAiNOiOeH4dgAGVPy+nkUw
f1Eg63DklUiOhcFlAf+ZldNt1I24KIPNcj2S+oCqfcc88RbjQcLTtAfh+4Wl8/2o5TxVYpPncOU8
hcpSwTymJ53CtzbpuNdT2GgtpVxHHIoFiYpDqc1jIvQnbxu+RZVrU2eT4f8bTDGkE/RZq2SKJzmf
JKJd1YUp9ipzREm2SgI9XS2WQ9l1izYqK5by3Ye9lnG3Kn1aUGq3MiJpt9bK/lI2c2iw4Ums8CVm
NdnXfKK3OosmhvMxCwuz2eiAXNF71SQzB7XbEnafkL05o78b7fwXhKQkgI+3RM3Qlwy4WeCDO6in
g72m8cL+F0HU+XZbXS59cT/RriErCMEgHlzwJ/wjTXURkg7W0WESY/vUK8IVot6DVhvX3L3d4YRn
51piMvdzRAv1XmppY+K75HJhcKlOl6AT65hFOAG6YmRIe6EHgv58UbRh8qjlKr+haHNi9YqiufBf
vO4Ga/5OxO/TYFOIOPPqt0UkEl5GlgJ8RcNgI7pXXpwYIublV6iv02weAo9twNBYMt5rA0oc/kbe
qTfibydFfLe6mUiDDLdttAPMRfLP4j1bllC35tIJvOVHX0HT+0uIQZU78VElrEsOaCE+pgnQ8oUU
WiaQiys3xkD+6AD27/ISbDu2AWtRnUSz3iPXXZjKtfQN0jU6ocM9MXkLiALPLtzOzx4fsOQADYjE
dfzk4KweP7dTtb/9yoAJVnmhWmeYsqeoymNBNmBcncLTLqjZw4jDmI225n/xXhz+Z/l2ZD7tgoms
9XZioqlUxoW3Fmg15Ad/QGQUOr26KKm9824QXTqErusOKPZi9uunZabNjDbLx5NUpOe0wXu3TyZF
F6SFJ3xZiU/4xGad1XFoVVczHbaXciBNS1JZEl19EP7U117fJiV3aVTVZ7RGNB6H97JzAhjUOk4T
2A/s86esEQN0zeKO9uuC4mzqSHhqQC/BGy7Nk/a1yaaEtRPuawXLZEIqRoiv1jQPRtwfKTU1Euev
K7qIeAynxwGAkqCkILx8GFQ2gTaM27HbxZa5vuNtznMfqg7QTTcitTdD6HbjW/Wzk32wqmK9nHUi
zp0ITqcsyYIkBsfuxt5VQlNdgBh65n4PbHtRsf3/gFFH4WITmRNidhoKddNLoer7gQ6KWZIts+vn
hAssMXwMRYwi8Za/qMwW9YH0OPkpxHjwxQQYU5mvWIir8fi17CHaPCjRcfcg1lneTiZmQiIl232M
AkFywjSIkrlnjIeFUiJRe/QzvXfwAwS89DU/hp/1+J3W2FblbugdBGV1KHir8GrKXdFavl+l/s5a
GhvOMp7IuBXcTVTJtBMxtgGKnMRWzIgJ2CpOM5EtpB9yw+/ecpgVZJWrBhCCfkR37ueZLZdzDAtv
Kc59ydegGXyNjuQGO/LGFyVW7vcLuUzoOOhaMORz1v0GlrnUGuZ6Nvo+OQORSYbf+x1NkGsZqLho
7ceTVYrwzux+C6BtCuowfAWtaZPQ1OF2EmgS7lx3Q+ospfnLu18/H/BNXv8Xnv85aWjeCxHqJLhj
qao0tyT5zlTf29Woifvx2Zfy0TJfUkdsjPvkVMvNjJtEjFV3YJbMA3DqXaPA98yFVbCPZKYGfL5o
j4vt9Q2HlG4bCLfvTrnmzG5s8uWLGGgaZt2lR4uq0zOKTe1giRgYphUzh2QFb1RGcQVP5m+nmJob
f4hN1b7QvAQibDv9DkIbt+jla2ENp9xLGiQ3nvPkt2VY4lmLPA42EH3xsN4CRwrzxl5Co8nUlXoA
+gVpjxtR5JJ2JeP58JdhSrEG2VGOPzfX7d8yHZZtQEX8ykLZuFIh+jQx3LqWQrlKKhcRNvacnYhe
umopv/2pUx1J+nfQ+IYoKsRwSXyZ29Lqk4ziXhwb/VSgybqcKP5GXttw/kLNRdN52ECkGqEaMPik
0nf5EjQPfbVV1bfDMZolQYloEC1VzblB10CFjUTKa6UStbizAEGZ5ZAXk2qL9uIt18aELdHUNvQL
3ynLcVEkOc2+js6tnTO/AEE/XMRnFCSwp/b51xyw5lugRhPCF2VNey8LcdPX0ndo/N3R4HQ0U5YU
4iNsWj2Pv48k+3FarSftkk7yOYWcdeO2cJ0zive78NpnTYPuJUJbBxu/Te6mlJm51NxyVRcx+lV0
i2N9nlUlynE+MfutPmEZTDibQWAH5CLNkceVQtHABHpziL6BLfMRpO5koA9+Uy+irCmvdQ/p0CGA
BCGjZCqRpoMqvZOeV5Y/teclYdFuMEvS/+LBtkcMRSAliNfDwVWe/oG183nTqApELqyG7nTJwePQ
SpVo6ZywG4NGgyzI9Ito7tTm30olHIJgTktERG+ywrAnTB8d+GNCg01es1CTvWhmRJ3AbRWhCgmJ
b64WXJE6e9e8x6nszf0izSu1mcD6TrFVwn8fia92a89uY/zPhvvf3d+ursBPRiLRdeEu6E6rrxNN
xtLyJkN4r8YCbfmx/X2sxkxcH3Kv/5HW5ElV969oLhBV0VhXWMkaMaFT6JVkRpZzRg7KkZ6gxtc1
Ej4fUAo5EeDVgllUpKgZjSL/qrzczj4OkkIrkkBrxyHfEWueZsCJW4dnQlXf3YbfCFWMe9LoY0y5
v0xtS2v0L9bOBNtuRF2arQkeqc/EHUuWKY6aG4kS8tNotRWDyQ86g+zdOkxSYZf93kjd5IDkg5qe
iA70zLiuEKJc6dlC1E7LTE5lR0uJEhEuIJtWZZqFr+JwReV9CIkHGUf9lssImyL/9P+Iw/kguzOM
KT5EARno1kRTf5P2xIfYUwc12QhcM9xZojUWpM9EzlNaxvc69fjiUyNVK8vpY5bkaFUmeG5PU49l
l7MkauV//C0vjILAzH8Br0qpADX+9LRLbFdqu9/T5AhA2D3JHmSSciVlpeKkDOm+7jWkYbq4eh4U
xuMwJXMxCNxAPcoDR3VoNUP4kfAKL3XSZlSuIFdDUO+vfliOjeYvySJMCteH1yZVF/P/MEPORfor
ofrf5lNFqTpjAXqjN0FDxniCeh+5jAcR8wgEcWeRe04boxrzkJlfEb3H6v7u4nVBCoc/t51uPvPG
omup0yLd06He+4ZGDmmkVnjh2XzJ7HtzmtzXk21tuvHkH82aZE7fI50iTIeeSk1euKoWm+ZORuKW
UjLZQdnPh/WmNc7Yb9zeD4FKWczh+gEMWY36jKttEmAHzQWE9CslNzHCQz6Lb5bGkYv30Iqa4YzL
8SEFVOFa+iG413pX7Ra1Zbo/vHommD4r75EXjVs0tP12RdQ4kIthE0llx+nOgjZQJMnpOqv++fWv
hBnyxREl63i5I5/cjgVgWpP/C5jc0JbqANGiikaEThyRg5RkgHMCl2m34JjRnXToQqzlxp7Uw4EA
5et7n7lUFKL0coRNnhJdUBj22kzgh1Rf/9JGgQSAdWnbOE1i9eviVDWEmbxrB1PSszXjukQOPxio
LAS4DZ9Q4owr14vAnFywmDAw/cwylSFIWoHWRJVtmbNl+oErADmSXhlpDy0g/CsQQzV/OVitegCO
LkQxGe5RgdCyRLwmqVEy4gtIvYZZn43GYzCuw+clWdH2CV/QI7O6Nyn0T0imqc+V2sQdGyYy088Q
I8T7f6eufWGhW3La3Y2tTTFPp6SOTDgq32fV1quI17p6w536fT0qRc6xuy0iK0VX9DaxpslaIRoK
l3TKynnpi1Pc4gkKY4VMTgzl4yuZa0qsXpLAimPcwXZGdk6s3yx1sk5sHkWgC8+a36Nod86PrA06
K9sJ28aFIdpRX2fKMW+hXBMjYbFL4KkMVZp0tIrxlsdFvwmZL8KgmeshjCOgQm3m/NhaQ2IVlunC
wyebxhAjCMKPufOlI2sBxiypWY620dJbVHZLcPC+GhyfOVKgF4v7aEVxNVsBe+xaNLJaquS33RhZ
ikfumPAx7FrBWByHqBLABrp8AcnaYVir4qSGNaodYcdQ2q7sugZIym0HrI8A/XhXv6Oc3fM3M/YD
nf7/VIfi/du5SZNNvMkJRcxPo7d5sA8yV9fZMylbvuOI0CrUsCXOatFYRdQPzH044wH6ZZbw4U6/
kUQpIF3iOZvX/e3CYtQre8rltn6AoT3sB3+5AiKV5SltdQsfT9NqDQbjzJqQ58/nrp6RpaUp2kJk
5cGNQYj+nsvNivGRo1KWZWdFk1Eu3WRh2RZRNGPRSol5/vCUzMuKgi0OR0c5oBQwdwxdNjM6PByv
P2b6te+HL5OPaFarv08wMVD9oo12NkkxjFwvLpNRMuXyD6rJQVGcNj0ccm/RwPf42GBnLhGafimv
cfIENX+Oih0K9UUI99D1HUEr0SY+Qif0nPTniKQNwKXYubHjPsXCD1Iz6a/DdOy/REL8zxtlGbat
InOfQnPo/NkGVLNWVdflg/agacRZkGX57qrCGm9f5vqUN4f/llPBgrTGGcroXKTAJ3Un/IV//2oy
7hMCOQzKFpTNqX4/QcQ1Nc4lQXi8V9RlBut4E3SOaURhWEVznR7cRvZ5czh404Itlx8JC1SPR9v3
RFPLajFygLuBrdH01Sig+ViLdGftxpClcRJABp3UpG1SaakW56KCNf20VSvFndawbmXB3sRrBz0H
hbH5a6xMd/db5ct6CXcpPCw55/Mr1r9nkWOX0hlZ+MzR1lYhGTQVqhygwGUhSJ8z6v1OEF78UNaY
GE3hISiMZtJeBGsO5FNcHs88/1h+6+2eW1nj2tVhCSyt4wk6KET4DkRgVl6+bsrw8/S5PAi9cSfM
Qa8I7T97X5ZkaHjqAsBSa1pG1hM4LkXgC4s5QLRrNaxu/6JdWMA3EMT6TYbc17cYJQIC5OEOrlhe
91HpGMhtuGowbbLV00dQeawyDuey24oPaxOY3nEM49cpqKLbMNa5qhPlUBUA4R0NevdQ4p9HuciA
0u+aiITUh1kxiJaAjWLrftKsiHBAOEpTz3ogQNPDWS5fN1EyPfp9rv2RIQSB7+WM3khXbeWiEi/1
CwpzgePzGMlSyFLOBjBmGZEMk2QR9LsExTDJyMLEsyGMwArHw3DgjeJSQ+x1vFhSABBpzXuhkxf1
5fHjDVKyyoLJnGMpLJcEPxJv6WBKb16rZ3SkwYBZQqYeT2SujxOZj3NowIUgrmky4oxBs5Cy9c05
j+ja9AGke2YCdg4qhRPRrYToAFsU6NifU/F7lXlcj5K6//Ah8VfZAHbAELKFT2ijJ/KkMROcjV6w
eIPgs2UD0ZKMoc/j9/j0h22rFF3JxdCpAu/Zc4JL8KhF2czuv2OkfgPSK6JpkqL4MECShJbL20gz
UeKjlRchXMXOfcySjeUB2HOiy71blYB6r8uVz+yO6uvP7WVdI6tvpV8yqHa4xuSXFuAe/kW+YY78
XSBr5OdhOHN/mPJZpHH01u6YGnTYHhEM2mBb74zSLydiBpR83LwjgqZ7RjeU2bSRBHpw+BdBZ4AY
nyGvpkcSKHNAhz4CXtUjmG/QTaQR18mZKZhuD2qzb7PAJnS17WkZwKc/CcIvMohkTpTtCXAZssHZ
vwoP8zRkKoH5AN1y+xGwseq3U1HbFHFPcwu/R8iT2nNkkrOyjWMBrA+0P2aq4LaCPzvFr5tox3eW
6bg4ciYzAUqsFbueUX4TlkS+Lpuz0vT6Dr5ouMAn/FdQdEhA8D8SA4av13GYvQETnpJQU4Z0nuhq
tUK1diFu4q1JjWwXkbYzQGi8eouPm++NDsKF3Sdy7nabfHX1IMGlcGS/5O7T7OxZIDTHAMhiFrKE
ooXv1qTSWr+fG1/pLaLKo060LrG6vc5GxD+JMpPcc8KFpeMw2CB2xuGoigbVbG16cuHvb4Tz3j6N
ipnOQHvRf133DXH8NIIK6KI44nX9I7bwL0xgDABm6M5z0vheQ7+OCCXsz5QCAwTcuqOQTvhxXwRS
iAyKSdA34FEVOoVOzM/9/YI7Eu9tLig1W1kxvGgqFD3yNh4S8oAnjiFmxi1o8rd3QRxG12u7P4OL
e9NLN7z9q4dN62njZZAJg1QwWNVtO8+WHzZVis7tFhggmeDsPQ21miEL/zQ0CA6zhEC82Ja/uidN
xh+YPyJpD15eYNF+QMVwcYApnT0YbUjaW7x9pYq7BvlUGrvyg+deHVkHE7KNmt5+v7azU/wWLLUf
Uukh+vXMePmrSeFKF25v6y2MVORzgQUtW0wsY5fOtSAIH6o8jbcGFUUdWSQG/01JI4F0pcu5ri7k
Vv6QwE8GVTWcahg+F/uBciANxKHRSXbuYyD6bqaMtPE9y+0KduIRBHo5HTYhbe4R8dKURYsI2dCu
bcTxNNNqMWimARqbtszatJXKPHIyPpWUVtSIkhhZZvilIDuzZZd0cbTO3sZXkiZXLtFTBo+vnlv1
oeUedbzMvAYd5xewhH0rcxB1UKBRD09Xj+Ze+FoNVvQG6re3+0WMsGp/FIkhhax2eTNc2c1H7vX4
n/hnczgPEMyQSpWhy/rRaCjs5nF9Sk5tHK91SJQMv/qbB0pBLDDvIc+4KTm/Ks8D5ZGH9Qvwa5pU
hZdTZVE+GudlmOK+oP8y0OsSIaNAzLKaX4jWsRH64H+klpIPb6pz9nDIPH0QpBg2DKNIsdZetX8e
mZpblCXJ8zIVwObdjZbJ1E3Qwi7q/DiZmTBZ1zLe0e9Iw97SbigN66jmkpRPv5lECTaw7TzFAKkB
LKmUheG94fJcsTMg+bwhQ6tuIvp5YMdTsFrpNLi4REMI4QgBbVIkXjBUvVUvMVMvlaQxWovhCmy1
POaHKq4tafyLkGAHzndlZGRNFVnnEipARil5Stx+CY1qumwBoz0ozSCeyqdEQxyoVIlw1eHBzyrY
n81VwbbzAaj7C3DMnGDzigExjp66ywNhmllhkr7U1e1d8OaIQ0fPWPvI4IPWVZhM0AyScZDwFqq8
IUZGGJ7OSrf85eaR/VTwmTNkAZRNB9THjPqc+jvVJ4tpJQaePV9FLVHbY8T/KcAFt84TRXYa/IJI
xPOivUIvw5LZ/Sj04L4SzCarYCEBGnYhV1XZaEBMSsV0zOEhLkW4wK76RBMOIR4YmSQLAsvJpf7e
w8F5mm1XeJRtuygn3gWxmq0KrP8FjWeMDj+NZraKR/Mz7x7bWP7k3d7KmTahDH/gVLZBPpIuWqsq
+j0FXtQEyIWlsdkZEYYxp3DdF4vpi6Hdn+H0mH5GRk5YwXl+Tvgxu/83CoyDqYPk4se2l0Zy8ll+
9tu/w3SLjuTBM+X0hyHqI9qy2vJMsV8KrXS6QlKpTwqungSBPcshgMaasKUcOQP0ecCKFzITiYG3
tuZuxKZawfVa8d/iITw434T+OagF2TEij0C6sGvTspqzEWZX1RUbD9yVL607IWKxpbeJmgSax61y
Hd/3DWsJKz5OVmes92SbtYanmh+9uWAdQctQx6uPxLPF9Vrk3Lgk+iWKru2QMWhIIEje43aN5b3D
/EbQiCf9Gq4j6xrz6a8ChZf6brUF6y/VhJlXCMwvAA09QnX8zBRgJxd/3qXfIY3L1H12TkqMoESy
7tVpWOlmWP212SVY70rRTCO2DMcn79ZbM+Z4ov2gKX9z+SNXT+FvobFIut0J9zD4YVc9669FR7C3
zXiDpJA80Hnndh0+b0Z4M3I5K722i49gGjjc0WlFKQmsdUn6NZ1e/+vXKAZ8st1SsFWLm2NkTRwe
ya2cyMNUwrvB1QnzYFIfJm433rZYZmOous1hsWDyCXPDkYpdVFdY+rph5EBmNEHCJ/nZ1jowU/LU
F/+Ztao//2e3NSTQ3DMJ6jIPwAsllfE8O0PMMjlTpvBQ4HrMf5Xnoo5iNqqTFrIQju25svHpirME
46j/BXGueqnKZ5KmDGH/wuN00ssx9pX9FvsH3hX8h56U8hhpF3FmtTrbkw8OI2XmNPavMSw8S6dS
O7zcqdvcmn+kyWDnn3LkEiAfNP9xMJg+UhiDT4E0WoSuGeIk3QyKjpKC7xMZuDOr5+1uFf1G40WA
BcAXfZ8hV6CRzogBZXmmeWALvHOGAZwcVtRMjCehyIEEd0AQN7ElvokrHOt+qovc9pQMVm2KP7Pc
cfNsbQcTAxoWL09DNXFX6CPz+vke3CLEZbwoJT1jISMcf3JfMdecRTXEqqTSzkCJ3YPOLWm0SVS2
Jm2r2nIE6wUCqJQygFVjKWomR6BQdI17bWBitNlyWHVVZjCwsf4dx1HhH8I/ECc4JkhEelxgDGa2
wi62hAc3AwF/x6W45h1BI1qOsS3L1MDEKTWakmfK5GTMWzfOvXbjDdq++WKkQOCfFjnPyaHOIG2y
oED6bosS7gLSSdAB/lViqFHafvliu/XfNdGeD09dwbcBLtEacyvpni9XfTBSLvG+oLL+xkWnq966
r3U2D7aO0xD4EdemKyTLni+b2XMuknPnOt89hwfPdpda3UGHeIcXinKM9bVKcoslirwp7kCzSbT1
6XxUO05CYFjVVEC1Wt0hVu094IewvfHgIAUfMFtG8TRlKV0HG3K+ZvwFso+Cwllju48HltXZfVAG
l63F8LXef+6XatsLIbzHgZFSOKoz3H9ZUWmDoxO0c9vOIWtZsVikN0vYeFbiuFprU1yIIXCmgtBM
ghuMD5HxgsKJL4qVZ4pBKZljWxtALufvvvdstPmSriFn7zMdYqn0/SorP3Ah+a5GoqRsokIGGvJd
obbtYxFcH5BQVlINHsjkdy2K+woMHpMP8CP+gb/89sxdTDF98pBnh5jt7XkA1er17+5KYxNH++uA
ZOXGNjzmFGQsCjFgkDcipUuAAAQKfNDmgy7G+lT/xxLjvE4mCpIh/Vgawx4KdMPSWpdMYaKntMYT
rolpcxcSMIQv7yLZkL7hrbz/S0WmDG7EfIhtjEF8JZiwsX3KA2LHcnzFDvGaddFF35A+YD6t5AKC
3RqAt4avAIc6+IzY08z5quZRFJTbSdQ2hUqly2JiTRDoQ+Ag49K3ZCInrVLuW4SWre0Nz4FFULxn
mbdehunos2YSA5ZOkwRCR9ux1jyZqP3G601pDrbQMqClhyPp6dTHqgOK+BfMcsSNrKwLP9eWmvxd
hC74mctc5p2b+anJiibky7rQv59hiKKAZ6SO66aiOnYMY8sn9BgKrL5ZSztzHQ9oFVfGHvlpRA8g
BsXGIMaIKcW/JThGDe2aCeVOuYsbZfFcfdZ7yYFVbcwgmjzwmOTibC0OifaulNVRQ914vHV7byge
igNKVGBIOLngYgSJHljpQafr/zYJFpE+KsbC93JM1ll0DGa0t2UmTl8JKEGN5bK0ucfUBZvrdcqb
jIg6r7vQUimu5nqLF20JH8L7hxnNOMqXqCdgDsKnW8rjtCBOTDSCjmy/E9NzZqjUJ7u1JDs8wFbD
IJQ1nWyVWlgJAE5ZnA8kHvPRbgzPCWxRg8JEzecCzbGbU7fqwQ7IXPq4yCvZHWnv02A9OsZDylPP
D4bD8w+ft8QZQk+QyVbfg0NhsVxzqS4aKOPo+SC6BbRI9CdjIfbXi1MynLYXP41HB1TSMVlymnJM
Dl8buHIC/IqtqG+mq72C+koj2oXf28dfYGuDiLEKiES8/Fcfcw5JZyOGZ49e63WuTbv4vdNjREKG
77y64qXovbHCJEMP6EguEqlADfWpblQ0nQQl/f+9n+kRbvOh9uaYL878avr+2Nl/K0gcvJHefSy6
TEQBmjUlv4itsK4AcbaSe2apWJtbAgVxZQRsffcL8HeJT9IHljupMU7oNf2C5Y3Lzng9V8T1clbM
o6fozV5J4OS+pXtdKTvlzBUnsf4G9RM4GkDSjoQ2q/uZ21JZgg82N2ZlVYIwHKc/IxWS+QfbBPO2
zw0IG7ATRLH3FPjrk4yORWO+if/dmIREYGa1QW15srAfPogvrHFZxAD0fLPhZjZKQMV4jQmwWnHM
ylPsXnmpPh3H92axTfPkJhPRQCggeDue5RcESvHoL+6JNazUJhXcKehmxmXhbe4AhOU+I3Z5eKMJ
O6mt80oWrHrweImWR5KaJGhUv8n3M2ViAkNZX+2PGUyyzhi80b9nqVECUIRa6Y4x9cAFRb6gp/Q/
VJxMp2Djuup/soJyokF19pgLsqPs6KMclWJksdFtTEWKeiXZDuo2+J7v+60h0m70j9/HkyED8u74
D9n8+SOsrMc6kKAIU7eTBrr9LCLpf2ZQGQQCqsVT+ENuttodyhx1cXPGfWHrBH6sv4h0dNfddJRl
hYJrF2TvwyoQonDkfiz4MaEIPfPrrqJFAlPwtfvgi7BjU1g42YgIc/hgzk3rR+LIgaqJyX63VrGx
Mk3jw68g7CFQH7XZYzOw9wKJujThs7lLeBePjBW6H43au4FUw/Tus/0kgQ43qabTvJkxgt/9EPBg
rovOC4LisIyaN5X501jgGdXHekqiv9Nt9LkbA8hUvCDyHNSIrt30sM9guTwTmdo5IOMUbEjerwkC
fg8IHTSUg7CoYHjskWSPI5CspeOiiiK6PIFAJnOMRI3VJ2gQAV8BNlNPnwyNfZzWkfKj8i2e7P/G
mnXTjF19u22FAg5JDjMRAzKdmBSHRsJUCioLx3MoymLor6cP3hvWc8AQp9byOfNh3rRMvlBCIbV8
o/AytY5vV9jtH9bG918qRPK92u7GU0Xf8V2lupWdXYSszCo6Z+uNFhC1nBrpa4sz3d5f7PJl2r/O
beSvpSxL1st+Tgj4u6hU0ZZLqOocfFXnLJQO4XK3GmEUBXuDgkvLZmWfvRHdYGrLretbVr0IjdPB
pSVPx1VTwpGaE2g8nD42PmGEcTlwnpwq5WHwaC0Vww7riAkvIw+eUbNXCRxINCauXT4WSpTZve1q
6KEC01ly8ziugS09KoK7JdDit2LTCFjIWVkGUItcCChkikWQGKxzMDEdkI3LYAqJ0FUYl+2RVK4k
o9Ulam/g4HgbD2ycMkYOsungig1+S52UMsXhk4wEm59zu4mNxobMRvIEqaOcOgWYVLPsbhtMKvku
sqo9xJiKgp0L7lLnxtLFXDHoxoHWkFkHuoqslRVRGqWtslHtN5l+XBjcAv3vPhyF/vt80iwn4zKx
k9xTCWong4pDSH0scQtP8D3qTfk33zkr9Kwulo5rsO9yZTE4GCh8HpMqnOQst28yaHrH53Srgoum
zqrf3Xtp6kQp+bdjp7i1AkO/Vqtr2ViiArB9Uwl+42Z7MkC7E+E8KcLOHR4MdAPnETxUNEFqSyUs
JCm0tpr9h4PXfF8uxNeI9hbaJeuLmQvumu+/bV/S6whg/E/uE1e7aksbKbIiuHKJj4TEMIIiauQM
M+uvPTRq4HlKDurfJo6BfEPUFv83kVYnJMzzGGBLjilAZJtQDgACy2kxWvO+YAvq7fojWC3nLVJv
XrmYZJPXMkMVBApTp4QO+56BqjiPuyI6kyluep07C6Jpv0qEOHKVuY+Q5dUE1n57HDUU5TfKJknm
qB9OtSYcwjLZkyejayNXI0Hej59ZPS5ixzOv6ygwqbYGuL/Nd2ImvYHnygoV4dhCGGNPuCY1pXKt
xlGXfPOfzAFAPyZgJ1tjyBWfpR6lF/bGR2QdEwiVySnNsAWeqzmjma4jvwttxdwT2VYm8Y06O3as
Q4+cDNzH19/1CmB/RNwpnBQs9DxEavOk2bcJVCInkulShbjj9exKUPuwTR6kjjrt4eRWD79pkSX8
PPNrr0J4KP2uRn5t+X5ZHRkFP11VZ4svfpGOYVY22af4id2pIYWCCsrCEDzONPQbQ5tFMbdhApDr
TGoZRQmNsO5uMZkdYKsG7uQtBts2vi/Jh5pZo5dU50bLDDoXgsbGTZSh7b+ao+KwWbk17ip5GXF3
HmX653i6YtNmHGyHMjvfCucccTp1JBj68WbhgV551bmSf/vJa1+Zvgbl3xNWxgdbJJVD+ZYOs4W+
weyNZYDseNlsyd2/e5WGMm6DdEPKau85d7cKyYZIhaSPBw9PDJlvnoHa4nmNSL6LDktaobVo6odW
89ZtDLavVwzEV73xXxdRuuknLmYgZupCHzg5xP8IBVJuKzHTC6gAhOUOLexfWFHz1FRQuz75+vrb
aEn3BKj4ZrWmFRlSW7UV7o9Xm/MAnjcbHK/QB2+Rq/TZ3JJGIVMnmf3W0wk70zkZMmkWNwrC9L1j
Z+i7uQAWkJgRUQuNFiCq8DM9e6aI52+vVsiNgtsHcK3sPnJbEwdBLNrY+Qg3FyswiB9/8+1hMv2Q
i8Hcb0P7JeMUliKe3/h1VgXVwyQfZ+xjld3ucYC/vCzECwX1TSqOTTWGZEczX+287r7cTvKdARGn
Gq4egx+CmjxBBkzBZVth7J72ffq4Ii4t59Ff4G7NICYrQUlMwNiSczwKLDuQvdFpR1pWLSNEfKPt
KH24QvgIRc7y4JEf3B6ff/fIoxRW4T1KNGE/k/o8z0Cwp49gRh4E+A7GKIb+hr/D7++NqhTZutEr
Xg2MLhqSpIKZ1Y/OSiGVW/y2Syr0jUJLOO2w0OpHMJQOqv0YIfER9vKt3Bip/jfvrtofUl/31tGb
Exp45CYGtJ04LMP8OK2gbyQnMY9qey93OVAMTmzvqIMOhTCQlmzdlHZAQeWLKEsytjMbagDoyG/H
+UnJbyLAQzAWZjjiRn4saEfWV7R+m6yi/1mK/8tpXmUW8gNMbvUdZ/qt24t2zlxYyr1+8A8lkw3r
VmU5IkDyGxgs5Myk9BQamKSAT7HeWSSWrygx+DjIE7AyJL+Dst5PqBUxXsQpYRrihoKKMEfs7CrV
l4ijZpPLLD6I/r1oB5suMd7yATRfumnDR1wSx7uZnNRLb/gLQNhcfgW3aaLsuIgGGzalHnR9nc0X
KdvkW53hGmEMUkpT8yceosASX1oMxinKpXoGXbMI9O+reRmq3if/WfNYw9kddWQDEb4oCFQyNV2j
Xalu4vkFwX4JGctfk/hWz79XI108hkoy+in7HvBxhNa1lW3aK7EAXnDodQKMmu0nqvoxz82zCW7a
tysVbUMTuoAdyszO8hPzZRhvtcYufV6wbZQhvXYxKMiHo1V0Y8hsWJqiezB2iTxpZ039OCWVybOn
E4X+tvDwfwfe/kxAVlNcxp6tY5/lp1HDHAyrY0kTeWFE+079vK1fLEZcrJPSmREHsR96ki+2ArN4
kB9twQmLSHEKNEbdUeKOjJ7k/Gz+vDl0FcT39RIqZSxoNSTmfPFf+wpU/IyGEM9ZEmlQdqEdtTkQ
2zgQuAov66A8A4Sx601X80mrfJoomhToitSXRP83JlXkUCuQN6Pxck3YRzAW10WKgnvdRlJhDMef
Woayw+AejJWsmqhgSsRnkRU+fvFJ+Tmx/FSMwTgl2v2xcc/a5f0X86hSzN23JRDeVFdPRprWBS+z
JnKyLvVU/fYu9WKB9hvBwj/pXc972GgzqToYrkX7i63C2Scd1mUS+jLUE0HYD7rsd7jVnW2dafBs
U2HWt2pRQDVvPIvViz0vI1nntw8ywHKZLeOTDRZYfTVCVEJ9AUdSuIbWCog4qEO5CwZqLljtFXNP
RSU8GeE2jIav9VHQJ7ttXZtdx9SuQaBvuH23NgwF8LtUqj5hju/N7MWoV+9fYA1NwwtnTjQPeKyF
xwJv/kB+1x4ZJGG/oItKN82sWGymr3yMJe0nsUPwiL6vBUEwEi25L59BkxXfaezkVBQGFTjW0+Px
AP0KuJKC4EizhV67UGHZppvv0gdx4rGprnYpBZSEPWHjoERouKtIR4IIoKe/v0TSdQRIpLYmpoEO
LfbFuIdSUYEUiInbxL6w3rh/8FIFmhe2nNw7SHKLhSLqLLJUaXGhjVVFpXMLHRQ47YQDKaBbb5GA
M5o3pVo9p8sdiELHkBI5WxNcuiScxuTaW/tlG+J5bWsPR981PWYmMquiePXSlSaN3y9bl00T1NaA
FfKIyTUTHnnOelR75QiSctVvQec6/xI1COcRmlPnmB7KbJ7gRdnDsu4x2jiwRayO8Z/irny5eC20
ZG3UvgBQ6/ZPuQhhlV2IX+t4BOJuutb+7ZyDW2rvx/fzZ1UAJH5wmwOf89UDSQb+KhQ7XnC7tCcG
YuP80VjrXsiZAFtU3amWvdat6a4hVJt+PmfIEeNrtoAal0Wyh7t3TlWIdHaqW7SocO8ulU5yvDfL
QYgQpngV6rDm58hXwCMHMdwPhpFtS9jw9BHTCtSVrN6rzPOxzzjlX7VD/bV5DR3ppdMqJYkyz0Lv
V3DlbRxqsFR7he+unSCryF49VyYsQWqaI349LW8pKzDN77sH6JC5imOFfBiNaMNIETuFrZkT9COs
MXCrWJ3zmxMjFw8h95WIO+ZWTucYGc2I6CtKZIQIvlh1eB4xEYuXckeIoGhYSEy78h9nFucCsh3D
2RS1SPwNksjcfy+YXAcF8+jSOVRsdT1g1Kir59LPvfwMbSriEOoaxn4fOkODe8J/8w7gr6N0xpRS
vdbhy+FECzwSiAqCF72F2RVOltVKyiRtJhip1M0GEtc//4Ou0F+NusOPYFo5b+0FCfeMU6jKog1R
Z6X3mdyAhMcJzQN7h6sKyKWHIiwJuYGWmCqJ8uZQOhd2es2VlhBvJa1ek/TUdDup+sCD8ja/sLcb
mCvePw3YOeuCQjT8fygPRJ99vEiRUwkNT8TP5yT1qe0TXMxyONE10atHjN6LEJ8zRMH+Pj4PxhCo
cHfoqCLoe/2gNo2j+7t4e0Qdjzy1Pxl5YC0zZGVXG9IploApS8rzvQYTc9i2ayWPCLtUle1tqDWZ
zKaVU3qI5esu7rIpgxP4ZqUFmNU2ypGlyLVNRhvf7O5HWjyPuDd9YlifCN64yETRepO+K6yXaEqR
NfHD/IpNTaALByKTR+V8pDwp7eZi+UA0LfuwD6eFa1nv+AcPmzBOV7XYXkusmZhXBj2y+D1GQHFQ
Zchh6bhZARzP/9GxRfOQ1cetlElJkwoJI/Hs+FTXSyYNfwmdTAYxPpy+bvUEDFfPiFIKX/thdnSe
z34Mgy9bpsBFqNFPlGeRYT4UMQnuHtoZ3L9YQ4W80XDCYexobupnQjBh9yT4wn1HW2TRuch6rTgs
5zGG11jvFKb+xNf6PUJKG7oz6iamB8kVdnZE3IFY6CwMeqsPtjQsXAvQSnXqYqOFcXcc7+tuIo4s
ragESFqiKPiARMx0x2lI5Y/3eCQ6GR9zPVjcUgflLJgAk3ujzwjsOZEhxxl8sDQeWhSdmtnrklxJ
6SFaXRcc1sqTGakTQZ1E78xBHPRLFP1T2cmeu+juwbtkBur7+sQ5v+MPhsBBPIBsxKsws3u/Av+f
jiMi5mj/Wk5GhKgahiODP6rVg6Oo+YBvob9pDC5hNGOvHCJqrIsG6kDpQOS+peQoFoQR+2nG0Ws+
UloPxhj5Zo1eOg319zr214b8r3c/RmWODmKNGvxRZOC7NDREIhOglHz0mzwbyevt/Fv1irxRQVZE
uQoMDzZhEo4wMbNFoFaGY38igZSgAq0qeX2q1F5al8r/PXzWMIk8vaBqSwmw4mZALMBXPSYkKrF3
H9Aj0N1g4wnhMMqrwotAGmYI4vqeXUeABZhFPhNdODuk3Dag9ruBp8dQroGiA90ItbmfQXkuizAe
y3WlbJzzE/7IokdtpITPE7s6ZJB3N5ehDNpE92fn1kret98mzT7y8E6cB117oxPj7NuyNTlDYXqT
OgW1TxOX6s6lmozTN/l105vfWbTL8rKXs0HwXzO9nvxInrA59wfRafrm9St/bG7sxpun1L20itOC
d5Sdj/ASIlj2q+HxhupISlUPtkdKqWJY+odD7D+aDaetPATpqn1JFy5KdAxZXsmmJOsWUxCkv8oV
CaQAUzLyC0ur/PPwteqTzGCBC6yfJc1csS+zuCzeYhaUYwqm2lJm1o4WtHD/fWt06WGJ3bURsvwg
1rouqSX1WV6fBv5krRQXv77xcrSqzWPwey9QDr6rM+U0VCUbAd6LGXeeeosRhKEwxaTvsVtYBANo
ozIWoC6IO5OKXfONNmDLCXq2ibt0ZhDhYkS7nJkvNbQa05uIeCf15DCRF7PDKfFs2PrJ0Z5HEusj
YrwEkChTLQI43cgKpG5kaPlap/CaeGhKFqrqFfI09n5lNmFgOE6V5jAjILhjQLfEnS5IRlT/+Td4
J5BMCIrTOLzWCMiQ4l/6a2ahAIU7uLOONGLH+YSTuD1kGAFxYH8VfYTTugt6uxzgk4xd9vH+ERh/
o+cObkQSTwcve+3I6wlQx8O3ZRc/7zGvByphSWQOnE+KopyEIGKSBq1bwIWBuiXgt8qovEoPqyZg
1b/qOXy4g2ePhoF1t+mC0dsHmMXXNAG0RVlRwMVdhBI3Iy0UORAVC+k6zRDzjNULwkNmTLMwGTLr
5NT0Bf+Lg3UsmD3pSoChHd6rzp4LhZWkfJ7vNYNic32gBS0isxtjs1ttAOzMLozyETiBeRaW0gqp
Lpw6EOdjCIpnedU5NcVW/1rFZvViqg70Hw+uIDEGCShjJ9MfkiRz2vBOdRt9RbtSYPBLYO4WN59c
gOz2Xp1Rqg2CuaVrMYtj1GN/tp55VvTOLMi96Hm3RomiQ7/uwshe310hiEUFt0U6nOx3aqlpD9K+
BRAhtOpucaXNHyzEv+8pzCdol4N1MKoSC2wd/w18Ysl6J7Rl4OW9YPKANWZGuUIhQ6yZenENo+Z/
JTNNzCp5K6XabltOPOOXfjrvGUFw8ClPscZ+Cfv2qrsr7oraJ67is3vpGzdvvjJcNCqhBYPNhHRy
hXVEdwVc0+DsXjWDpZauRPlOXcWJ9Z6PLEAIWjIXAZv9ztAqf+SgytkI1syl/STrGZKEtH89lN0C
kjCJCcW8lcBw8GSQ4ze3G3CG2y+dOpzcxpJ+jGYsqtREZM19/Fif7iCrpavLbaR51hu8rEeplyzU
UG+SdqHLrSo1d5vlnJEC3Oiv7GL2BcOaEYrMc9XopBBrNO/qBeBiejzU0txSX7sZydaO2n+gJ8eW
hkyOfwGmm+RgXliIGUC0dJTzo1fMT8xt2oqWsizPY/eEePpUlZA17HIiFJnlMKDlyBqGj2M/3Wtk
EYWtXP6R6o+xHHUZyQyfkDr9cqf6MrI+tCwXP2Puu8qqKWtO6oBj2OAMvYHJ8j/5dTtasaTg+tzI
wI89/w922HJxvHkO0ygynbZhuLBhF75A4U6qWo95YVWslDoO+4C2aAvM/VKkyLhaadmdFJ1S/qm/
7r9UHFbCu3yG5mQ+BLQpws4Omxdi/OEWvPPe4iS1vwm8p4GrFssGXp4X1ulAYJ0ZZJ8hhmsjx2Om
nof48oULlMUTmI1Fgv7cm742oUsfTCAY22dwpTdgQD8eD6QzdQFTQvMunpZ6mhoUL/GEVxwTnr/m
KAyhHC4Rrbf0Om/7FvB3c+BpAHS7DaNm8G8oumBnfW3QapHkuRz1N4TVytO7/DI95cBK7Bh2niT0
hi15+KSSFm1TF2A0yTAap40TFA+3ChmBF0oRT5TINs74swYONIi4omSgsHVHSCBtQkZH6sXRIPhj
XJqcsEVPXkN8pgwv1b77hIdf39wFT8oQgCcGvJeGPjuDsH87yW3ZyHW/lL1VTwi+Zf4np0YHXxc1
tEac//FQ3eEL0vo1cI6zERzXBSNkDNJAwhJ3FSdu7OE95hd/uyxwnyGmVho9Y0asQBsNNv+99h1e
XT3RoRJrDut03x7+WxzyLuTJSv/F+e1LFdav2okOpwnvmj0kOgbiNw6P673iUHslV5sPYgHzIinJ
3Xw5YaimBAaa1UMuN25dI0jZWqJx17KD8MHgtk2XZo8Dkf/3WtZfrPKUruR6PVk2yfLBZyinyD07
GjTTeZCdZxrvcUn3lqm1gJ6q5vdx/WeBRAbf2yctKklBfJd5kQAV65u958SlU7RkKPlnJcLv5fTN
Axx6XYCMwg3E7WXG/jh9vnyuy43wLOFz3Vd30l5mbwKn8Sb3ftGGg7OuS3x6XYUSTP0gHYOOMCiN
IRtdgjZTXHVgOoNN7kvJKXU8o8T6NdfoayueTTnBOYj1+HOPf2qalTVOtb7wTLaBGxmnMsh1+bJA
AbNHz3SZ3CKYmIDApTtwMJlmKnzcHrHKeHwUoUGlQLDNFtAYyrgTI6/AS++oBHCqlpmnZnWn7ULF
f+18SqeuYWH855aJ3oLl0zalZjv8NA12RG+fIIXF7MQ/wfCpM21OZU59n1Khle8q2e8fPdXHpsxa
1X8SXDqhhxwMIOoe8jGuo/x4cn6jx4EMpvFH8bw6pnmxYk48kNqEY5f+t/lgLwAXOuzLmAUHp9qP
Z0rh/FBSPBoaFyB+XEQLJ1QNh7+SOshgda+m+RhF3Q2ZPLvvqJWTCSE6uFs1rNjCMNywepHQ6I2k
0OoNwbKU+pM5ihH0BVUWx5O5QZzVJMfYzn0ja8JvDJALdFarFY9hAdK2U8WqTkOqTwnZ8fXjWsTP
vue11tnu0LLCavIHJP9t45xaWRoxIJhifeMTfBEnWGHSXjMJ3339bVJ4Jpxjfdk65zoB/3NwBcWA
eCXIXCv92NMrdDPnvYTcjhNn3K6kauEpuI+yl7E+V10kSqawMtrC7S5aejozljkot+ytiGZCQ+Yc
1YBb8wREz71fFJwIXdwAqeeyMYv3kPtuiHppSwkeNELFdMWQIkAR+LEy1pvqCqeIR0+VaQ1DX5Vr
Cd0roq9yQPQC8B6hfvunpRAXh83Tz75FTj9TMFwnC8W8OmiKvvwEeAPxTw4inXZFyQ6AhJ4nhJEd
baIXfqvU0x7+aTyXxj98uPmYLjClrGKhkDSGZG5qX0j6+nRob7Y4IWPibfbhhVAl8KDxKdx2Was1
A8yK9nXEJ3vqozkIQAOR4t6FiVsGqsYZaEe0i5T3QRYUuJP2oKz3rfzJX8CKuTU7ELdSIf1iSAdy
paEvrNh8zoHXPMes/e9eDtvn74fYoBOmEVQWELNnkkWU8fGVu6KcZce2Otc5L6/koVpn215AcEks
7ZfsTd0dqT30/FtXvwO8F2TXYzsbGuFkjYT2JyzQDCkwfgDJMjLPFC6hHvfihLiXIK42PXD9MaMW
ypaGd7qWejK445EufE7JXKlpRN4hRixoL8Xmbkvd+Yg4MVNHoUyaOgchPDrt1hfvFJkgdspgKdDE
ieLoTEqO4fuwM8Oow4RJ8UECgiv64QRWD7c2o5XlDhuhg0y3lYqKGcz9lImCYljtAZGWUk7q3boS
5bXGaMAU6RFEo6FLnhRl/wJrBJPRowZMuWaeXhtkvu1plXq0ijfvbty2ypnL1km0XfRjRSOdSzg1
R1mhqare2BRhAPNIaezhNfe0E+zyZCbcymf9gwJg0SMWJFwHVwQ4XGDdb2ryIPg3EINg6sGHn3Lv
BPM7EbNB+eTnU6gjRgnGeffX6rEKwET0pVj2kzw3lD99tttYGbufeBGntnsEf/ulNQ9qRRoZYo8w
BNUHKJTVIjxIH3ork1JRZSxkOSgMzwrYHIorkWk4/DzMjxdIs3oZZl8+50RjzxRpCoNPo2A9Vu4k
W5qEb9wdk5IcD/L5+/gN7tS2Z1d6ouPG58tQq1+Uk3VAhPT/VhdQsDMvsmpm4RpbSIgrvCYeZ5Yk
0+yobi/4mtc5pdJoRfmyVuq0GJvLzRaXg9vY/krFrdnObot5IEIi819WwgwuVvA67ubdrEGq0H/Q
UNxn6MeoCyLm4IpI9Ygl4l1Nr2CjZYkyNaY7UDgq5cw/Z1eoBjaFi1v6rh8T2bslG5lcnUQhqhqi
GgRwvxYmImJNT0QKS0Cq1zmrFnPLsDHONjM2dMAy/CC4Ej3/D/BrSlphqJhv72pK84WDTm6DGrCd
/NBFQspxyqQPv+9GHahDzPweSw6xWwHEpQJDPNwZEUuK6k0yEyoWJG75ftzvRh30QMNvi6zZWKZn
3ciIi5ssykEpPZCo9wluuC/u140w3bgFFz0wU5qPb7gJp5PG9Yv6b+RMnwGjLSQCctGDhKZfr+ml
A1ChnIV/q+ciEidoKW8+FsljV6JMt8YPJnYOje09CVqYWLtkQZKMFm6g7dWHRZl7SmNfxr0xe619
pSx9lSAbkBxoXP34iFO+2B6jgD7BYBuoBHJoJWpUWsWtvy0shoEJ7S4BrUyrvy8ciyL8i48FnKh5
eXCIGumttOthmEKgofzLwVncKIMPhtcN13KCGt7leWwgD3v+bwIJDrkTQ8dS5DU68xQqTRW7KTK2
smCO0FB+kNIf7KHc+2x2LJvXciZNbfPSaGVr0Z7s0EV515NcCCE808ri0kOP0OwydH7hfO0+QUM1
vZwMk9oZVA8KuiN4g7DE1Rg07BSJ5fIH5igodn/K5aDya1LY3D4xNQho02kJklPt8B/i3vaVebFe
LbF9iw1mKgD9330YAyX/PHYvuLWHN8z/KJlyKanMPjcZVhs7OShqMYHvqKGLS0o/Z3iZ6yZSrz4J
4hsBUBdpMj4FrBkbjh+PmhLfi4RJQLjofk7+3iMu0rJSs8eil3DMB7Dk6V/on2yHWmM0DVq9t54p
YMpblV6laO7eY0iAAvRCYKT3vcBndzaDTIralTGOkRFTB8Yd1ZiKAO5G7SVDo5hPdHHYQ2urLRoQ
xwVTcWdcsYdpNN2JkO47bZYS9TcIYo15eKeyK9u8nelM4loQwgOCD5kqzcW6dkMMWwK1uwYDvk/6
p1NqLLgEWk6iUZyaiGhmFD6HhUD7b52mhsv3V1bsNXRbNoByfDXlIwHhnwDO+3P06loBNprMf2DA
dFAkjFS9Fjl3SWs1aBDbip6h+j63yCgQYRGHlIlrIm3Z3GoxLZ9t4nylt4GUAg8MEBkwjkdQHdgs
NX3MPTQYYbcOMiUSb0xBpiojxym/EOJGIxBoh37wBkM/COx2Hv1hKQTXQz3J1FbJGT3jeeU5Nd1J
IPJhx9iIgtcXhXgsZqKh/QGtsWSHxKDS+U2Q6t6WLuTfbv6xzncuuLCQ5ctJobdvrm9ggY3gpzuq
wv8FnIovEpp5c2YrNfx/IDZ5yF2uoJy630lEZjICpar5zP0ysqrYHiOuYFPMAj3QYFVXH6nmNqdJ
iw8PPtsjjcG0NlzEO2A3XBZ+AjaVNJowYfrx4WoSsa4/yenbc0EZqYbPDoxQlISTo+ybB0g841Yw
TTGBd1/Er1/Vu5sgPqrww8/bYZ+oeImlczTG9z/JgVQKajalGj0/a+4bMi2qTDDt6ZOBF3ESL5FU
XreQKUbJBdTFpbz8k5wkmbgoD/7lPjbzA4Vc0IkQFmuZi/MRLMo4F9qQVlYyL6m4vUJ7l2xxjhei
5N7rsFYQqqGXawaSS9MdDNRGAQO14rcPWn33ER9AljQre1L5JtyTsSDAeWSA6MxWNnZ8XLCPzyoN
+hV+x4d3MHLxKsoobSuM/FfyRRef3WlUgLn8ZOdeBAK1F3m/LaAolKWqqee4SEcZndP0YoZ7FRCD
6L1m4+3nQ/I+rGO8S0DlKLewoNMjtKDXtIUfr9zLOPCUYCXzXY25wFXH0fwr4xe1veudlUyPxg42
mcQVXTNqeBCZqRIEY1ZN9VsbOBGv4y7U1aV4AuGcMiqmDG083dbp2Ua0t9Vvqe3JOu+oaAc77DS3
Sd0/tktiT2X7WMi9hEscb+CYWO6vQaPKr8mHJfNRkRj1erSVEZrCknoFF6Njq/oWM/5MoNaGpusn
5XUG2i1zocu6ChIQAlTA4poER2ocwCPMx+Oo1XZgXMPQHYeF6j4SUi9F/DvDIggGha7s5154tGMu
F7Ruc0r12O4sD++I6j4deH/QfUaDduWLon89gVPXF20Kx7rBWooqM4RAezRHQQpSE7e9PyrA9el2
OMtRjFafWysI4fQ34Zu4IwGsWS8InqB7VRVRA8fxofuvgQA4ZwWN3cjUWwhVZPVmqK6EW2av4DAr
VC8zYggv0Zmn9ETILy3PePa5dCJoRb9TJX+ZaTzzv2ddYJhP6my9mf1hY+vbLJrcy8wyyIsS+Gl6
4/7nkXM1gJPTZnIDYhBrkdOoGUQtORzzriqia+LkjNWLjXr6nM2FVO7KFmqg3ekTHsF3d8EkbaH7
rfF03wzi49ZMUbcE5YwzJgX+vnL7tsq9dJB4Im6G/ir2PJFHK3XScPycTii58s1J7BaaVLgfjr6p
3CtFPf9Z2hGE1N4ciT4g/Q3GzwjNvYU88ETC9sLgIiA2XWePYNAlevyTGC/BQyCcAY8gG1f20KCY
baSlT4I6WS8qKlsZKR54YFbgxDVMP1SQpIMm+qkWMK9sR4yJjf1a874Qmiy9ck5NvVFpVNjydvC2
tWyzHsh0Ks7T2eOVb2diplpjzrk9aIIZgBbP7+2t4UKe7r66m5+Jc7Yur8KQdTCuCg0YAOiwjR/X
bsjnug+ya0MJFLbVzpWDLlfs0TsNidUPiwpVkAE7QHHrtBl/mY2f47f1Cybhzd5kntEIAVOshOdr
+QOpBSVQQLGzPJvubPy9DUnQU789f9zqdMnC31Mxh9kGUGNek0agv/Hj8knIz1JmdyXyu09lHkqQ
5HQcTG3aGNRqmp9EdOk27NakwgA3JxJTvyrgQUX4mMB09jJrUhZSxvVpMdS1G1rQScq0mG/tmPwb
r34xsLJxyHC1aPJq+519UtKU3oT7ADnkO4l1qcurbQW/6hz/unKbSip8d6F9VkdrxPcqPg5ds+1k
bU6QkTIYor+vUtAifnVekY+FnE+MRsKkGeJFh1d6hKjKIKU4RLXVMuYoHhAxfvvMiy5V0J2dTPRb
aDIf2dA0kFFhscXkdqyFIneCvGYEQyBnnYbL5Ol2RhyPJthcBxqnltABmbtmeWBftuYZe9FERm2Q
+3uo+hsvJDnZiTgrFUFnPIPMVjoLNaQLmG4k3eDwXjhzmP8ATGoHvGXydLLG4mZMiII8vgWZ0qRK
moP2h2Yw/jhzKEgaeigyM7hVdFHfIWaDJLQgFzmdK238413jpV/ik5Mzm9U9eNkDOWjG8AQJrLaC
z489qlRU1jn+WjLZpxyIwGz/rocV7/NCPVRc7JkH+rc7IfewvlbxH1P/uFLzP76IOa3RGHqD0Pn4
IdNKPMl3pOCVDpziBTKRuDf/ROv+OPjvkzl3RX2J7SdvB7+C6p2Ad4etekXQJnuboneijZNsKqwx
LgdmgCHQAsfQOQRYwW+2UVptLFuAKJi/3xeHzyyEhD4zX4MLBJQGFdV8WYZ0GsO5oirisCMYebr9
MneF6PkOpBi6bOEcHWXtF+ySFBR4uPmm4b1Kp9GMWc1YaElZXmLn+Kdgfk68C2miv73ZeHsmvSNQ
hLIHtnODhF/bxpUPXhplnbq2Qb7lKSOt84jn4kU+7uDnPGcVVOgqe1LF0LuO8H57/d/3VTISTm7N
CaGpMXeAFH6YS6eBp5ScWl9mBAZuSEGLdVc+7u7+cMe/LALZYym/F7xQc90s+mOqZjaE6L6enplJ
vpjt4M26m4na/dYA/wLtKo158fAw9wKGlGnvbn/ZGU92D3U8fixQPltsOw0p+IYJEWBe85RcVyXm
W2FhFscL1k/iKzfHTAegqk0upjMc031BRiJrcM59dqSUEk1bTedb3GPsrEOPcMNkvlydDc9TrTln
e17tK+Gj54+KvT7nNjVXqab0I2HouY41uKZ1OXWRKR7iWguB6kMRwMMWLeZ4Q24xpDUc5L4ix5c1
kBqIXkAbI+KimflUljk9I/JxApRfObGPIZ3iSiUk7qei8ignsOESdcFdoXM2WcS0ZsmCCJPwJ1YP
6FVMbsKhbU76eFKbnrSlnjp3I0BmMWqSVswlCLNusOYoNWju0lFUjOGyulSms8nwVU3q/WAeW1Ko
2Z45JaZaocTiQlp8Llbf026CUeV6Pj0vSOgkHR+RKPCSkpWZJkdz+D6kNW/ndDS9tknQXX9hQHN9
C7Nlte24qX+shMX2Y66vTTJr3pwwfUcomGmY2FEgm59lQgzLld9/a6rYuH5rEdKkdNR+ZBuw9MOq
D1y62oqZ7ceQ5x9Li9MYOE/xsQ4RmYqyIHOPICiOymJTFiKvh5Yp+lHV9C++eeq/0SAqIWV78Wug
rMLd0zp9yp0vD/bCoCAfaR/hGWW4nzBy6hWEbAsCtm8WBYKvs+PvijSel1EyvdXP4kVUOla1YAKS
6VXK8PeqdSTpVYzm+rupLZqCc2MFJvKJ/X3l1L3JsbiS8UY7IdJNZQRfTSpsq1AmlInSLmIz4paL
iYyhiOPLEr6/DWnFX56g3A9thcLekbF4s6yNgB38MdYaKOpBewYwP2BZF12D7VrUIE3UeIWkgUv9
+gto5MiVTAlSjR/aVzpcJCp/s98oWlAsPZE9HSLUm+xnSaXdrHUZWQJ1ICT3xkaXM6Uh7F7TI9lE
sxsoiKv30YRNaO3SbNrS+KjK33yCgE4PbCzfZpD4c/gLM8TLQriDerdWS+jKFB5zALu6sLe+hF8g
HF4ieCqVKNgrfz6FnGcPG2sumyz0L4iRsSAVVNYAApprR4DAKEPelhJmLe1ZHmaV/z69tzRdy8pB
mbTzmg5YObZ5mf3IJ2Zp1WlWEfOACX0wK5Gd1bpTfaXfAEbP5aO6+GwhwK1GXrlbRDHvT4JyZgj3
ApD9FqLrcIkL1fKEEMhr3/zt6FOO7AoBMnZmNu1f5h8cTpuCfFkOBcIhawFdpWUUXBROEBYswsNB
KDwH4zoDExRX1SCXvZ2MUfVLl8SvcQ0pKIYk4OMxtShjE2v44MNy48Dq/hCVS8nlkUv2AzTpa4Gy
rL6G9j3EV87y1zATvmgz4Hmhq3fVD3jIJEAAls5eQSXLWS6hGNWJJpwiewCUhZkk4zjEgwXiDsJI
JYUusWcbOqz6gRoUjpVzPIUAtOFq97cUuyP5YpwzuskakzYY+ONoBFZ+JsQXkcJ4Vdzhf32Vg0Li
GXaha2YqHIWRfC5ROirD632Y6SH0SuqXQk7nvoRR9UP+SyqOhWiHBv0da3jrSSkWaoDdCTlMkur3
Qf2rpHjpn95FdpiNzWyDzfsin/LCMZVB4zCKgpHBdoCYHlkrUpVImTaj5ntvBMMuV6gvMiIuVlqT
oBxe/Z8Ravu2UYGZCSgcDIHzRXg25LS6VEt3XRcaXENfZZWAx7t+crwRcmhDKYWgaoZkNIxRpuIq
3yYpBwxFNiUGrWu9iWN2rRJaI+zfl/nRSZnORi3RHcDrKnZAcyKgAoKuwepRXhD1HWOHqlHu34kj
muNzMJOURZJcEdttW8uTi43r9iV87KEDpgri5oarwJ47Jv0E7ZaAOlKkZGjaifaMBfdcuiV2nRQj
YNclAiGNQ//0MayomxQ9K+0Q4w9LmgKOtEUBZeTz0KgtuZk8cnGZEwSWQOjRy6e+uVdKHAG1PnRU
LoMHrFsC3IsdY9QAK5f5WkjbIVL0qFDuXXWrZ/sXCyX3XF3HhMkoZFYRI1T8sHVP/V+uttSrAU8t
PJj62/r+PzGC8zXUHR0uVKKE7fCmqMwz4o4iUOCeKE/Y4UD9x6POHpH+afsrRaF9ZPZtE8PnrbHO
+ST1mOBFpFQ/YwdLGkMP9YdBd38nW/5A628ut9SB2qx+gTC2Kg8T8/6LThbcuBcN2rxcR/H2Uvor
dZtfHfcjpJtO/F/nzeQAx0ZAgu2cz9h6JZv5S8V1qUQitqLB3Pgn7+NoY0Vl183rM4nh+/b6lhyr
u+3cvIIjtXwwYvtUZjvmqHW/+I+N34pLrskEdmOPy9SMg+iqGcGDUmDZEehT8+R4eWbdIWTDpwGF
68j55Hgp+t00RELw+LDc3DJ9ZufhFOMO2bjTD0fE0VgsEfZiWEhFkc4ubdsq/K143FpL1EE7tJNx
jMeG9U35ch/b/U9jlnOiXC/FhmPUR7NMuqtVfjh90/pM4trTFgM3L+vsMNaBNaEAU9R+Wz2EU2Qk
2UoE/P/bdXaypOCmOrVWQ49eXILXEkDlGX50OaoLWRhVZLTX3K2GCXuoqSP8NkEHnciWObpdIz7X
g+KbXY7iOkJ3NkjNbOxhLUm8Ilg0nSIKfNYFtmQ2c0T02T/hLn8oVb4wtWmPzRmQilIDeos43Bpl
ljrkTmWj8vxxqDuMGDe0GMxcK8IcbSRTCHAK70B0/vKwTMY/fIfyfJBycpBtcjxsS/Xlk2HjsG/7
l9szkn8cRl/cN5cTWKG7YwR0s5fw0zxD+q7oJ6V4Tm0msCfxUgDgE1TvjggnnFLdLgf7gG8tQmxa
BTvhG+IJE6BqejETxKV6U+nbtt3JxjZP6NZ/k0BHYY3gV6yYvLTYsWDKZkoKI1RBInPaZooANgc8
MrcVyQ38Ue4aorqn3US+0jPmCr7ioqYgMVj6HkhHMISsjXjRW0FcKbQ5nDFxQA7viAhx2CRmRjSj
KU8ICIqva/yM/5pQhXoaYXcZomonoxyOGdv+P+qsqjimab6VZEwOOkyVFY2BDlhtD2Qkud1FV4Jv
4HnvZMd5ig+tW7+QNtYEkIjG+deLfd+f4Kb3dCgu+hKAD7L/Li+mx5Igkda58OUAcBUl4FgwPepd
IvzkQSrtmifK32mJCWZjWHKbuVxIO/p7sBdFto5aStmQXawxMtKZoMsRY6GViC8KkKjBXQrRPpzz
2FGGxcJKPu9P1IBmZW2W5fHqBsJtaIDssQ6gAn806gR3w4bx9Jv12oM4ht/p0Pew/xvDtrYwWxhY
/EJ5Zynhe3wVvpX5rtjcH+k6wsCT6MlqDjls5cPBEw0W9aDx7yTqjC3RKfTS/x9F/LInIBM4n+4F
ChI+pzkpkfVnRIRBUzOyb5Qt7ajLB6r4sMo7GpzggWbBrw/PETYvd00ihDiw5Ve5I25/RxSNxr7a
v0APejd9W+taB9lMkbullfW2vStv/mYhLtgUUYSBfAua/dTMWZO4DWtzCTf/6LzxO2IYpgMRNkAR
fqrYs9qYleN/g/zJK0znHALLOcBoXp76MFm9iYrJ12qGFaaS4GNM0smrrKsbg9SemHmdP+S69LpB
U5alOEm9cR+GdBzaKgxsy0WlJ/DssivZqmY0A4AyHqhy8+OBbjhS1aOEKTC0/h4F0OTYsxJ3b9gu
I1K1nXfG+YlDsu0PVrhzpLJ8q8CF86BqJH3oKZDrc3CmG5b8xOMahKVSauUPNdyH3Ztvb7Sx7yB6
24aVwk3gHvYtbhJCC3qcK5MPzjLXp4a56c0iXEF/x/BlDi/N/yGazrFGDCdPG97ONOTwdDlwPCx+
pOMcXgePvrD476ohi9XMgnnPtzrgDiOWI7pKNVw1L/VkASuN1M3ZTQbBIc4llK7eF7n60PGD4YVJ
eaLjBnJ2kdDZl7Cege1upiat2VuWw+xTk3YFMTNaANZmBA7HXV4Ho+SpZrjF4f46Ojqtr0wbvlYM
DWGGs4s8Nk56UZBzl3A5eWlHjGC+N0n7BY/HrUdDw1c/reA+s3aYs43zwgRiAVd5g27+2RaHSwPu
qE9qaXZwcx9R/3mFctMbDdGFiP8qIbDMfjxTkULcGR2EUQ8012evwfvXpMaP0ZlflgG1AM64N4xy
RqACqqZhTmM5xLzSJxbIV77WFVlj6l5JJAX2WKrR3B3zjNjYJ2EtExs0AP8eqXAKSjxY9MLfzGHA
Va8FWseft9uhT5hsYwdSX+VFupghmgHfIYzK1DDi98dfSH4HRdHgW7k0uVSYb9pGhAezy3VlyGLE
B4cORn1HLJNSz4v0wJTUAqvbUcJ5AdwDUioT2lBTrwGorK1aS6OOB8zZdA4KjgBBGs+ceQ1D1dqr
s94lqwM+vJ4i3j0i2hvOFhN1GLn8LiqARXZTjskPpa+hAsftQI5qovV+inDFjLkvPOK+iDs/QKaK
eXuCUFYvYOW+S2aKQtS8p0B88e0nmKn1gSal1+oFvDjyJpKJlNLlulhKdLNChNMyEqC9ZTFBkaCS
SijOtJF6mL/0bgl3h5DtFCSPHm2MWk68+ukHMOIlZIUD1kDBe2XOgJoK+30PWDEC2a3EtbmPtOmd
Ke1p52nhrr0+Q4VxMTeXSZOTw0Ymk64OebB38AImi+Cdr7/uKuBbuOPQRSvANnmceR8QBiRfNRR7
PXAZe08WlrZrUj9ffR30jIonmtxHWOiMzpgPI+EASRTdyc8NLZHGDEcBVAbTLG2QiXF98CLFE29K
pfumgTlHcMwL9r54X5tICOgQNSvTNS5bpzT8oKsyjL7jE0D/3orySeQQTRBukfi9H3j5eRqut/lj
vkdsBnxzAI7N4xkHC1DwyUZxM9+V5WNK6xCsfn/d8rurYIsF4EhGWcBKySzOOZwPVRPqzgtrOQTA
XX5kxO2Vv3EgKD2TLRFGBOeveKTCGA5HomPxIAmUZ1P1HVRxZY83CnuF+bPOiIkoS4OlAYvYrY+E
dzZCZw7QTxjN8c2j4vRTJEcaxWaF+faM2pR6f1jOPOmw/prLV5w6QCe4mupH9qvYliWjsf3MqRee
kuJyd/ar9Qrq7nBPrOYVJceP/pkRKx+xV006CnlOXMeD2qhyv+t0GuIJX0FDPT+aEZqlN+w07MtS
aO2f5PeifozyTgSDXcMOA6YxoKP0fgdr5Jsj9qEVK9Fy1mHK1jP9QVI+QV21/UGvIVS8/AjoRLn2
mfvsInnnMqaJ3s85w/XpunoIPclrlBh7dRhr3K4isBz8ffv96n673Q8XNGmpHIDbty2GrwEML/QA
kJFj3NwhkTw0J8aqYBB5pQDLBopQQidK44jQOvWwHZBgO7raL938VfhtR7+Wcktg+udpcARBLVXy
spRyX2xsYx1ddGJMpZtGBnPp1MdYry/4XdQUIEIO0LGW7tAtAORtqSyErp5+zUt2aSm5Yyj4khGi
4vJVfAUNm9jzznxK4iVAmp+6XGx5WXgnW+UqLLAviCD1Ask2AP4Ra6EQK2/FzgdqZpPjObxn7tAs
Lca2vFut7hwpf0W71ua39+lR0JUIEe5mE3O5HlAzhjiTcdFm4yPY6qeGL4R+t9praIdaVyVUnFIL
9dHUjXJjHXRh/GY0z5qwJb2d6cgjfAeipebPm9sXCRkLoEjL3M4G0Umuyl2igSC7PEtvXObrPHcB
9+q1p7t9nwx03QOISrDeL9NMVyxh/yxYXNaTmAo2t0DPuB9FuhCZoNtUqnyFWqfEnPtGATakTJb+
mNGS3ky4+FV/S9EydaX2kWuwmskgZqOM9jO72LNdW7DDheg0XIbT/IiBqcx9j9aR83xd6/thfb1j
5RjMEjPVcHJ8IloK35G4oSo5Ujx+usfepuyVlHmAW/0ZFX4kGvBh2dJCd10jkLVRWhj2PGTolRzL
hEYHD+DtF+EM4vzER63JWfQLSLvhepIcY1vbog6f7NLkO1nUzRMB4IogzCL26AFnoX2CIx9ld5Tr
v7HHhN9069lykMQtdjvs1RqQ3LtPwLr0wij6IZhzjxRvQSbBjCFb4yi7gP6Zynf+4AQeQMurj541
XkHuXVQjkdVRlBomqhXhQ6kfrDUjCiETWzknQIGHZlUXhJ8jb3wVmI93yQ4XDFHNg/HaQzzKaFkS
470fCr8rIUCaGWEeiCgUleBWnN9mnFpp5qf7Lm8qHSuLU0WBaqx2AMWBf/1Cu1CRXh3n58aUFRFx
Uy47laQziWrvynVRVAA4lzzOpQOQjlo5Js0j2vNdzX35x6RxdRzkdTibcQV3et91jJ+7MV9a6B1D
o37sOcg2RSMwE+dRYU3HshvAfAvCxEEgiXWghnXYq+DUbAfh3q+/n+x8KbJyOF7pS9AVaMaGhlUo
JtT/oXeCB4+CxF9tvKY3fwE5+a5+ZO4zrmeDGexivDS479b8ASK1Q+U/mjVlcDaZXsFQt7oaT+hs
AcC8CiAeN4RA+bqMQ4gr2zno7w3zqUx8sqIdGoGrs8cnlNG8yYBBJ6UxP/rT3WQSIrqy/lneTK4Y
bR3T0kvGxFVaYIU9FLEYtEmf2ug1VWAUZr+qwcFJiLgsvVj0pDEN3ScNpI/22xPGZj8WDE8FBPGn
dXbWD7uK9CJkQMUqN+hk2szl1s72nX+uq7l4bKaGQ5A9zL7peBwFYnV8grKjkS+1wOTJEIy6uczK
1uwmBuEODXjY2J7iQkCtCDWg3XqaKUJXHI145HSB4CqivJNEHAvj39lWp9gCO3siVRbK//eCdi+H
5E2LYzI+R6q7BurcUJk87SvN7yhibsE5ubOAkLA4nDEvyWMhjYkFmkdNo1XWfRz8LPlYguAnTSg+
iXTrYhRyyK0mrPcbS+XIc25OKMa0QDcMlia571/r7wT2KZ/KwhtqwcJ30xU6Kr0hbdUI39xGLjCU
z5GYdiaysRyLA/I16pBbTN4p4v0W9ckKg47v8Z5WGHnYYmy9T5vAAD4THGv/LuZl9gKpvO8dO01z
RHvL5PvFc5ANFm7FyZoLfWBqv4lsVTR+oIQ3mbvkcmeDop4STew5LJyrRpK/Y+yVWjNKggP2QXWe
xfCyqNp6c4uIfxwuCJy82LLCIt3r1svVuwXCB867ci3JtD1RDO/qRQ4cEHViaZrA0eUxePvUILY5
9kPoOaWYLKxI/fvtx0BrFZcaCcMiLU5NbMNHHRCeeHisEFzB+aPiVT+8gHAWD4z4cK2Lp1b8xmDA
QsicsFXBxPS54wzuA9dEEpvpKLYWHJmwBrwqsoa0rFIq7c4SEIPdSzD2kSG9YXk0cZFVeoiRTkVD
iqVHqUnJGXPwPOjvd8MkdTK6lYGg3B6HngoKqf6xoygy9+sm+HuSdFaXS/Vc42Y9+oScGdCuBYKr
c12fLzb9c2954lZD0B3O6N+ML6ABCz0uHK2Ejqpb3YKvJRU51tIJrZSiHn7kyt3ZSsMHdHUJoUdr
VasUwvLEncCX88fGnALMLwYYxgIkW/Fdo2LyIhrCqyiprnUFjto2i6bAgGxkmwQavynvJvo/jmMF
AqozX1wYw+PHSNBUZGjcdrE4uVNtHwprbjKw44FnTCy7CmdoiEV+ADweGzz/6fcFZjopIwzaPu1w
Wel8M/VaWOHWhtSdJQ8x04gWAZYzFQ4D1sr8yjzjn6kruGX6wibNnVMcgm2noTZvP3kcE+nNzUjZ
1QMS2V7hFU09FYvBsOesAXyj7cvXhU+ACZyVhkStRPLmVN8VU6cHLtwpzRYhnn7U/HlMuSBrj6Bp
Vpho2lSC2tCLAJLIlE5mjUN4HBXLtllas3n7s4XmbpzF72jdBnWbozsaYCDjmvJvppaPviIJjrCO
7x/5KWosM5UgWg9hY1voXklVD2lPA+21QxFUqWIqg3LI3vP5u+sp+O6V2rCnXdiXC5yjq1PFf+R6
6HWNuMjuDMZotPJPiezvHxoF2UcW0cTaUjBPnIfKOzmeu6jG9MI3RbyzKIce19/vQ/FivfMqn8RL
V2q1O29cOLmuT8vMvUQEGd8eGcDI3w+njR4F22inhuGjPGkDPeEFgl2im4iK4CRTxHOwgqlfmGTM
WdB4YNfkXKJGzadQUWysk2RAKV3XKdXSuS9YKbNC4fw5qjDKFf2PoD0DEOivrLT9+pFShbivoCOy
92ml2pjA5bsWsGveP9CkH+qDknCeJ+unhlno9gMPIX8mU6SeGXOhl9eZ+bzk84Ia3Id51ewoA0id
MYM8sZLh+7w53iMfm45pzRI7VdRuf9WA7YOOPr42txRgotgGQoSooWIdjwVSciiJvUO/VrulJEsC
Kqp99fNs+D3r62vEANNEY42jakC1lCgtTe3LtcpqAxy+Eg0YcuQW7UWaYD+ZGnVptTR8i0lG3LNE
HDXHif80rLjeiBvd+MluDe0CEmI/vdxA/0xfykFRKpmwX/HXqKxk+yqnFpdtNYNPIyifzluODAuw
FMJC0jaw/c9h2km13tz9lVqWp0ZIGjxoPfT/rcs1a4snOA4JVerx2aj2guIb32qWFwnrU8aTwAlc
a5y1T8QhsZFn1OXkiMrZKTLZ7dTxnT4HC7vm46W/YEFyeOTprsko8TQ8IbuVihPhnKNXTPjOx4fn
lDDNYb98V7XbcFeD7MOAZvtZKpdOsciyPXOtQiCuvMx80IYIhc8IOs4FJ7OrV/Bz2qsSOzXjzvgX
EVMqDM4rH6QnIPOPqX9WMv0riJscNbV665qsRQ1IdgKr2geQSUEXeaCwusOkPvJcFME5ZCcWCxPA
Lna27wYbcMVSUY91TI/cK4Yn8dCyP8HCIqp38Mc2j8Ax2Jfqy+mKti098VEu6olA0z5GkSS9GtWE
JXtcGqgGYV22Y7tbaVB+4sY5FUcvOBs/CCcpIZJsoHnwGqgJ2xz8+ROzodu1OoM53l7H4/1LJAew
zd5b/NTovH4hKXSzaBm7wRWwLVzG3C296ZYRUnYOk6BY3Ir/uB7XmH32e6c/VXTpVVIUHrd0hdiH
/j0HjLup7xp1ynhQNpcx1ARS3hZ23Kxmo0YwV93LJwgoRCjGT9xcDc9X48uT1nlgM8WL7z4ubpZX
q0c+HFpEdQS7jQ97Jukpm28T/1AHzVNZ2bOOba92Ca99OeSIBK1WT1bvCd7aB+Ny3iIgyWXxEKtW
2wW6wgxEQzdmj1u/aqRPKtHmGUG0nvrQ2DsBxTB4q5j2rv4QthkEuNjdDHoWMHSo73eyrpYaFKJB
i42ESRiWa52PpQp/A9zXB036rF/7gLy4OJzDxia78kU/yJv8HnWGc+lQJNvIzlW1dHwMsRPtoBle
oxFoRpokvr1ywNlJRXR038UU1bIhmhxgqXWb0gn5AFTvaecwKClczqgQkx8UsN0ghhbP+ywN2kNG
glTE5+4naIl3HAV3clh6bi0b9KY80Kc73DW9tF1632cAndFWN+skEtX1RA1UolJcpuLCJjSr2aXp
IRHIz0bBLFxsZ+7cGbKZXW0JHa5NhE9k5ImS/6Q3GNnlZ6Tlb+GAFihSx412BCLTJAGFIEF8blCc
GLrteuPBDIfskoa5Y8cdYLCGWHWLCHTgEllb75LuMNlerl6b6KoYacjiUrVbqXJY718uvg1sfPOD
m/rV6BKEdxRiuazi5iWLyATggK4itPWzTCElcqIRvOC4GZw0BuA0/ShuCLnNv1Gel4P0Q93zsfNS
xh2PVSxGCSpSaQfySRbr3U52sSWfYyjE98oVyZDn76+2ya5mUdB8t32dcSPWYX8UzgPli5pKCA55
pTvVeZOZdLi2sMO9+oogS+5WF3ieK5/5ZeomUuM76FaGDbSlMoLu002AO32u7OhgnHPabaE09+Xq
xXkszHCYBh+hspilqp8GVwf3cGkYX7flhGO53kiEg7vin5WUOnDeSsPJ+WVTUW4iKVxQP2Blrc1X
Dq9SVT9HeQCI6M95YiHmpzMh83l51LyvctIHMj67CIOX8eyVhCAk5p3IVYjNmOv+FfiCbeGpaXIn
CSB3Y8w9fIZj/jo/FszUyGghzE8E0mNHzbAXYSeO/jozrINXEq0+TLPDeutyD/dGK1GgtfLsauq4
5yEtVFvx+R7qvneIQklAJFlMK8k0+YcOgEuCJE0Jack+C5302J/Ide7lS04/5tTQ0Fx8z76a0BHQ
eOQIy6dLk0kwCOVrLiOtGFV5ScJRgcNnKhqbl55nW2OmirJRQ4F0c9Dr7QSirFSPFfhtX7H/XFoS
VLdNK9K2DE9GucdO+brZ7yyZuDNOa8743Fh2PSgac682rnaEZe93cuQVV7QcRRBxkWzNB6k+yyHN
gtIIWvGT/8OR1ybPFAK4SWQXFZkV4BHVLlUYHKZbjvhE24Ag9UUr0UVFYiITbI9GePJkf+D/YZMH
HdhK13SVEmKSzBR/cW053LMwE8/E0/0RdmaJy7TYrIA1o4OtHx8s/zTV900FZEyHyEJAF9ZenPzH
ITiX435x7UKuikb5sB6SkVl2iNr5oA2Tv6y37vQkvMCwhwm3uGFYd3F7U1KnRIy7F03gA1W2do0R
ipvYXS7+e3Hbwc3IDa6NPl54OEryplCIAagplWsU3Cl39zefwGPDARSfKoXlygzMdKNYeHZM5g0S
8dWd39GbS09Dn4lDCMBqMsSLQYRXDO4aYGALwqvqJMkY/q8k+EwNiqlnT68DXM5bzlugnkEkpVAY
s2B2BXm9eTcUEfF5FL9cqCooCm3/s112ys4piblIuJpenM51ORCAxeciHZPO3sD2b20C74XFujuH
GsjroHjRFYTCnNeg7vJFl0DLRQNzlQQvxUFsle49swIwhcjRoKgsjWl0098jNbcgR3y8elFWVVLT
bsASceFikxneQ4cA8IFDD64MRK5LF1HLP1CoFxKOV8xkjH+Vcdc9m4/19K82INfCEOQxZNjCKM/J
KIexTrifv/iFpEV90LwloBLBljcNimmwVoOQ5gM4xswJxSHocbrdpIFiaC4LVRrg84kmehi7/KMV
jRvwWAk2dpnWJidTwU6VYaV5nwLN9dUXWvehV2p527ujZxoctij17PV6GkazNDqkLk/gqoCU4vTN
Tu2RAss3BC+OigyZJvjESXV6hKrORzZmFovAOzS7hRsUW/f1rppzkMdS2o3SfCOPo9t1hEjcvJ18
P14m07rf+gDdVRsxfAGajBjbMls24xHuZJQapz+yL+lSTcCGdrPTf9rzvBtPRXE04zYLtnjAmfgr
ki2n4FTZabWW3bhZkPbwk0NWakY9RTltLVEqZHjy9RJlJSznGa3Lp6bJzCoUfpZcUX6fjWis5iMa
LXCZPcYFWMEKZSpKjDre0qm+gHps5v+vSt16uxu3iw5sTRjxkPWLySaZt/+O8aJrYAd4fTXcUhWA
TXFS8LaxvFK65BLJMb1pjKGammWsTXf/v7udJn2+ngnteOh/Z+4Vj28ifCyV0TAG8v5HrxuL0+pw
b4Bn+z8N0CJkiWCcZROte8yXBvArD1ZtVrGpZgbcLmgI7FM/dZINdX4RUVf0YT1qU/r4zAt6uIxP
k4czOkZIdn/8kH3g55wLqsXpseyaEhqIFe9mkLbzzQv4A0Kv5/3Xtwn3OfIQt2QPWMEpUUBWbpg/
F1NO0WgMZJ0bbUjjNJM/K9fFNsnb0FEH6aJ1650M2XZ1HaH5UC4+26pipbg9FDzoDhb4D2TJOU2f
lL15zTtp9VQ/6pDOHIu7+lEtKh2Q/KpukbtzBwngE3bvGwHs80JiogDWlIDgv3JHUCNtsZWexCNU
mj2jzcXkJf8sR3aBSzKNW6FM9wyEfbc+pkQ2uXfNLqPXaQlr5HKG01TIBAOdZQHSpG4Fr3v4hZSi
wQluTskoxLwrdKjbjM9rLHguSY1sR34f692LmYp2CEzjsYj5DVPNuoUprJw1yG7JJjasQYhY8Alk
maIkD86toYymUZgj5eJzjy1wSiWDvTOev5Z19YSy2bXXOly/8qnIJJp/DQpgQH4hnLAWatTSJrvU
TO/55I7nDIesm/j5Y50X4AoUPtnL+DEJvJFhgBuR4jK2SvhYJMFhVlu/Z8gy5wHHEHKsGeIXIZ3P
KHHdo+3J57bGHNHXEaZYKBug8/l0crT2w3y9WDlB3xHK5HwJf5fdDp9FGsgyQiXH+5b0JyH9LSB3
QVoeXQA2ssPGtXa+UK72C0k8gmhjwwawE7gN7PLVR0/62W0ECa/BhmQC2qoQl3EEzNevhfiMk/DI
jLTaAX/SSIE23idEx7lDpV2v+T492stPHlYyVwx5WqZQf/G43WVByv3+iTpM0meThfeeUZbsrMnT
p1KyVf10nCzs32ugnb4joaVQDHFcXjIwKtSsxva0SmPd/yK+2UlthLS/7slfl1T1w2y1ycAI+VIs
5X3ubVQtieYE8Zp0ggyV4J221cQKC6L8XhRuf1HoxwKhR0jOf7ZQNELQKFycLPucz1m26t1l8zjB
ewtagUo5f4yL0vCbd4XP1yiae9ncf5mrRIfspg3B8NdPiX61riymraHvFtbM6y6dhM+d2noKx7Je
MXZhadHjxaLkDDtWB3w6Lomgy7Hv1p8hBVYb/fLAQaB1wTDjKRJDecdDEpXtynoP7OYnhH3Ys2w6
ToGSNPxYwsGwY6wclvyeh5AmkBmFc8k3BtiXDkeetci6nMCNyjkMZYd55/CWd23C8R7Vl/D+Px5n
+oaj6gXHzyAXQG2o+5GKRDDal9jwVolCkg3Xqh2qF3AZMggGgSbEB9BT6qt8obwoZIpi+HxfbSXs
a0Zm9hqre42dbyNFKiqcPHm5BpdRZ74qJJdHJg0g/1Gn6HWGFzq2N6usPRmmnZfNWQbBLpifgxjP
1dciN16vOcOEJ6IqRdxAkSmD5AncmU8z6xXSrbSZtV93lrxoEPvv8bjk/uDT24ZK1XYyWBVfwxgy
oZzRrTQ4vZjzCSB5wxrqOXjVjs31PWFeAQ0vp7bFCsXqO6HOQWy49ylWtcoNssMp74USILcBLPQO
2i08YJwCA4mn6+6y1PTBWYbQNKCflmdLr1fRtV8sCc3JvQgZ8MGsJafDRtSi5T43Cm+Z35Z224KI
hhfkHb0QsjkmVm50eupIjo6R9P4x0Yo0Mzi/8ICcKdWtxDSGq0DntaIr2ckXP/NF293Nx82BL3yM
bJTK0lk5Fq2bj2jpv79Gt3zIFkLvEg23fELZ8q304PBBLEsX9IyGbJlhof2Vd6i9N+rqrPQ2TLCn
lnYiz9367z94l5piHya2FBbvTvFwR7cMXyk1EYHPEhWMqbqHLqinkg3hZ4hRNx0inzApa12orY14
3xLDt6OqVu8g7gQ2ZDOvgbf3rocmaiFlxdG5pJ6xTApmPogYc1xksFSjUKzhwLja3jXUDmFa6R0P
2oSJyrVJGvA617oDVp/qTGAaQ5HGdcrZNKcXICmzCub3Yajibq+6Uyz4zfxTacIDlaVh4UnM0BTx
MQSmuQlaBpHuOHAznOj1tp111LUTGHdiPBwkSDFZC0JgMC1cZuzwsUX0neIyjDRGFMXbwxAz55XQ
TYVp/i3xW6n8FCnM5n0Qg6LQBeDDvLWLlZDC6yCrEJf1pike0zwz3o7tm5PpwXYXIKwyGSS0cbx6
uDqaF2Q6D7+v9qm4G/a6O2DWaejMckQPOXXp6QUN/DAtzSBjeI3akkVzgSwtGkkVyGF3UbZZlYBZ
+L862hXOAixIPZxofKdE429tmElybV0THhTBaJK3Vgy9vWR1F70CZEvqiSADw5wqqgzHPM39MFYg
uQXA4T0g1uPqS+b7pwivAd/n75JjBDCD/57/sF6k88dDBRtCmb+0MifPGv/M3A9W1dSFlCaOIxva
tfHViKPVSEFuUBRUw7yCQ0vEHai8G1Kwa6/Ym5eMDxW8MLVGjn2lRLYqD6WAbPpnh/YgD9GyFx8k
DDvU7KinPznBUHhQ8c+HfCSuReM5H2kmBQBCwVbK4FBjUbKl+1PcLdkpqIktwNLnGJxZ36dajnqu
LTm8wv7o77EoxrALGVHYGklVpaYINQ8qf0aud0hh6KUTKDE+vccv+d0ZAuzzMvppPaunjSFMK50k
Nix/+KF4p4Eg35tl98Q4ZcX+LClmlE3dWr/SezLcQGznK0VkWktZ6MmydzeQkJLHgW37r4Jovp2j
Bb3/mFS8UA0IY90rpHYggDuoT+PyXepiUabk5fHmmfjvSy06RbKvrityPkQfUYEn9CPC5smzy/UQ
1q591mbFA4nyMv1KWfCwY+Mm6mv4/SJpRPLCocqxiIhHFFj00oxLxhhDECgl7Ifn0Lo7yi6HcJdw
kedduLnmdEj+5mHORM0wFB6pC6lSg6sxcs4VLHaKwocpnSsgq0iM4sHaM3kc4SMe16IwZQHTuADb
//DL37bjFbX6+cyfLCf4rGMPV29QpCbsfS6Kk4WiA4VQCUwfYCjUkx/azutW8gpKpr5uFUxjAQ0d
wGtV5nyZ/Ub+oeqi7GSaIEH8r3ZbZFH9zum6BzIJx0A0gqZ/zVvKSUMlmur4O7ApAVJrcoV2u1xI
ZhLeKDrPLF4UjhOwV8HN6aEaI++E2kSlibtlFM66a4z+S023Bnh429uD4jM7MJ0LrN53frGozxkm
0FnML8FDxHMjvYG8rsa7d14zjw4HezgP9BqyqrNtAlS0T0buXftefqjkbvIqx8dZm+Tj5DXKrBKR
Ta7AUsMY596hRPtSTbUGzziTs25wp3h5AWC8PlqA+S9UfvxLhh9iLvY40XOwHBXpnEkja8eUEUCe
uP9XBU6qpL0/+3z8Wum3F97qX8t7mfGIRp3WVbVoX+0HQmq+cChzS+zqNZt4d/G64/9R+Fp5cs57
p803HeL6e9shsX3zkP+QBLKN6+lJ1NwEJk77HRKppBSqBb5xgCV3cqdg+I7aRfMiuMVcGqAWRM+7
t9iYAgR4ItYW/SbhFV76X+HEcDQF660ebeCH2WXoujrqzpajZZWz39iMVKHO4GOuXs6brSyFYK+x
EDsBz7+UNzH3UNl81Di9hoymsMQmAgXmdCh98cpAQJyx0/P66fUpWH4kowwllT1Wd46CAWuIavzq
sqpZZjvtoYYEkkyu5ttUcxVKntV6XD5zVVuFCwC1u4T4sW+oK4jktmqSWdV7UfR+oMH59x6m4Bos
LLQAw6WE0Avd1ntqQCNTxCpUuOHOqVGYoBrku9eZKapm0Ya7qYsvAKndXH1zQ+CiTnXX1/ZEzlBM
ZqLJ13/KZgmpl0lP+qSDvrloGusTdkXadezMDl/UAZHjrRP2OgEcS0fzY9JUAfXrYw3EWL4ESLlB
QJXlPbJjTnP9LunJmwUr+12Hcw/7UgLU39mLM5KF00ymqtoEzEihZ5rS6I9R3/dnydTtISrVibkA
MB6xpYCU92TdbDWK9kG8cv5wy/SWcCOd4eKkba9vSCGzhbzVn3HvHxj3fwZe2lxfp54P9ttUwPos
GCyC0P9FwZmZFYTWaOwmhGUo1IwJkWdDnlG3MAWvGA42BXmFCAj+bcmsqBA29o2HQBPRxitqlCDI
Wjg1cuKcbI3jyZnW6qMUeiSEwxL4hPLSIPxgJEApnG2xxlTJ7tcUf8Wq0vGc0PA9k7LQrjToKF2B
KuXlCmVqpzEBnINhD+98D0cBJDeONMsHGcaVk9grdh6mA8EPuI9pPyy1bTrY4qz6G2iS4wtT4A+a
xWt5V2VA3kC5M9HFKkHFdE8yhbdUlhe8BTRFC8gVAxpFfoP0Zb+ZcFHQK3djz8gFJLvpoCTz0mX3
KQiM3Qi8VkawBMeJduz4EL03QloaM4dJYYJd4I9Xu3OVy2VlnCYqNrFjfRqYKpghAq/EXmwurSct
iR6J5TZs0KtWA37lq86QW50ZZGJgrX2UuFZXDSdx5zfUU2uaWH+gbU8jle2RziIvJy8j13KZ5oec
nobSu+Vcn6lGV0uVwEY2t9ZhEwDY8VRt/Prixn5W2PPIbPikMgv/mYwhcfOVAihvGTTPwhsz+8Jz
vb9Dr30Cx/Hm/OXp0zmNmzzF3miplSAlggdmLLvu2uS3Nh2cQb66Gv0031eqpvgo6E2dO7z49Gax
GRGM8c+/77l72yYSj8yNHsfEHlHZUUo8DAjctnoEXxKYjZWOo0oHafBCRUiD2Pb5CmfYKbgr9Qh+
GAd/YWzhuUyPpXx+4ieQUrqUO1OcgxyXYGpcSfUx34x1O1TyYCCjLdl1WHV0V6VhwIQHFf8P5X3e
QiPDUc72RI5kMtvOcKUQNIsvkJ2t22mrgTZAPPnFIncSczDVQ1MeCjhmolr+zCRh8s+gYrZyckWY
ACMguGpyYzAtimbmAJK244TO/q01GXSih4aorf7sQ0uviTJXeVFftK+ELvZcYCKp0Tz1RGvyITDD
2KJxDxCvWpp0zmqQyG//ws2uEqR8U/bxqf8NyLEwppvW3nM9NdgvVPf773aU0zCJpV7Lut2jw0po
aw+q9JFRa4qZdR+6PWaKjlc2aPB+jVnVx1urgSxDQ4in5Jd5bJlsZ60pTZgpY7LY+StNhFCDTd4H
e+5a6GkzP3yLcGtPG/zZjwSfwVPrFh630TCPgoRy5XWeq7A6B65fPnS1cNTEuVP9QNVqtLs54Q22
680fxZ/Fr8nGfEjQmxc3PW7cAVhZAj+falS5SLnUoSebZLcBZ1wQmNtXRHLEJeH4GMwse/i6obpM
aLJEQTBEmto40wYPsr8hWD3YPOxZEive8Ma1BUcDxkX5GrYME779Ki21o+a4xjd97j8ICy8goTXp
5aunl1d6vRbT3c4cj6h6CU8kkGPie9LOTzbHiO2Q+FP0zaumLLXOEjplUt6cKj1WXVkNKGfwL3g+
Jb2bekVbwCV/0ZFa7FSKXWXESxKUB2z8t56SuHzsxhTJ9O9+9fN1IQzJfd27kYlt4D7qPn2m1Wel
BEhR6tx7eh53Rngh9brHEmFNhayp3dxA1rqPQ6/K/J6ytxOzrfenSIWJ/XD6s+5K4I5catsmirqB
JVmPaNixrtErjZAb0MqWXyvzNZwfQwA8PLC5BczYbgXVVaop2qi+o/y44n0hMN287RQHKZ2xUKzU
hJ4I7ZqW6yO71XpM/Szq9U1i8+nr5ZwKKM1TNknKPKAEST/M5M17xLFAVpZySDCRhwzHvWEI3gyv
2W6wpEU4WrfwX70852H1TYG2WxQ8VvF2YYOGFt0rWuwnLB1y9zs/BNuKh5V+w5NG6LODp7f3m2iP
viHgw+P7DBGwHReMCVSSFe7RyHguEsinE4Ld2bmGW8LiRM9TbyC5JQe/pXtwL0yrN1Z7lhKVaCKB
QQRnTgvuZXUFhXyxXjj+MIZSUTADVFvjyLUojppf416tKna+2hEracOkf+hqALEfbPB9jM1/OjVj
XD/GutgmYH+bg7ysp+N8FMIOvbbVqw0qsiWtcWoHjytyImuz8e6Gk7VqMXenZnhjK0DFhIB3GQE7
f9qN5ipCvCbn+5IrCuB6w/W33fFeuMKLWR7wXY+qbNm2ctHWWOYUqUqa+vml9ctiFSHy6YEKN4/f
aeUPsoQsN1jXXl/uRqFiJKbyh5Fu24cQUTI6ZsUc/z8BF7pVJc2i+J6itN6+U08wFZq/Oraxa2Wm
ZIzNTo0K/frKIoNZaRdykEQc9NEtvT/+aDE/eUQ6v9+GdmyrJ8g3YJCn0/71SMOgPKlCrlXHPF/0
UjobPyGmUrzMIC8J2NXirf6Ec7TzylTKxgmEfv/ab9Y8S15BWz28eGys/OQhi5QEgKZMXKMtO6Wv
ryMOI3iPCw98aV4WMf+Y9D7/+hZzvZN5B5A2Mlhv2BCL9LW5RyzHjnZPaUWWyBMwHVCU0cJG4fYr
7i5gHKdmoDRR6XRqdAHWniJXQV04+qGSntFFdU9ChAcKa0ScGraRKPX4TUxORQXyJDg5on2Oi83B
xhFApebyBqKxEUTWzxHVw4pC18T/tBxaJ4VoIq60WH2gNMMqif5HQ0bKDjO+1s2hKeoTdtjQwibU
BI9i+UHZk1DJszczn8h8wwGJEScxoy4jlvbPj4ZakTpom51DSHvcU2u2hk5mjt6N+v8hQsBcCkqI
M8a+xO8UXIx/uuef2NKYqARsrKo+Ing4Fdm1Z5eGd7AZo0HSjQtxfAfzC7stuItsUv+I0b4LEqxa
t9cf3BX0Bq3m+ikwGqkpFJTDXPap4Pai0i8x2tZji0I13F9XckhVXp93ebBoUseioqpsTw6RZEqI
jZoayrjD7hB1Sf7//S95e5uNLE/V1/aF8S+J9hTt2ewaqPuzygttD99h7pubMaqgMdTevUtcFH2X
+R/Ka3HzW9fNb4oBNFo3G/mvWbE0yiGSVUXw9UI0a+ulRCJaW76EPSTlE+s5iR50bI8VLF9o5jgS
k8xadTo4T5I+aRWTBv4L2Wo8OB1WiuH5oEp9OFp+ko55Mxr1omUc9bJIr+0zkReqRj+Xf8iVdmNe
CpjGQ2R4a7pFxNirhApy3M5ETfnvBhAnjpXZoV1IAxw0wgSwlAmMS5a3hT7U0/5DDGAh1QAnoZgf
X1+UScQpnzou77YndD9sHJp06ZGLigZCuZJnZa4cE4zTapjzYBJjJxpDb4bcM+xHDQJ4mR+YKKVs
WgOZfVJ4gE2P613WpJsf5kC1lmcIZDuE2Y3ZAaRO6UMshWAr+OeOEtzqVx1WQbXMzmJAtVBW9812
EzWZwpPkh6N92tGdoZkVgzaYt7RrK/k+kH7NqVPuW8k1b4CSRm8QO3C1br4UNVMccN5yU+gt4jJj
+zMlCjIuKTF1riWo6ELgYGr+RUg1fNR2jt2+9BIMyb1hN9GYy285NWzNXkiZLshRQPWMySrD3mmL
IZJ56PzxVP5Gv3BCIolhnsPNakxu1ryQmkyQaOmBqS8zx6omkOLB65tYkxFl2FHuEIfnpGwW5zJL
q6SeyOy0NrKX8Wmx3kEq3Dbk+Y6Hnim/omGKbCyHA8p5Jzdq+JpoDcx8lKnFHJEPkRlorvBb9LKd
AY5lx2twdOYT34awIYSqAWCQqqyylea2O4nxSKXlOvnfmO1ophh8jbSssqbfS7+v5ZH27LWpDHfl
TKPIzvl4cX1De2+rqzJDonIzn81QszZVujABvKu0q33GnPkgptoKVmxpBobsln19/ZsHK1oZnVrL
fuZ7YWXTkeqEvoZYvN0dZBzdezG+WQhylLBKflHf9KBhrzpkMm4Wxnzx5c/QPXVcPJEKTVDuY84m
xMMWaFT33IPTUXVke8z127vsvj/SZaewpZiDKKyupV7dkcEvb5+8qBay4cKh2dqcVWLBC6gdrvCg
bJImYgGSUwV6iVhd4fRkjWx7OnV8G/A50/yAUU/6XtRfRr+BY5FKKTZKZrsdQzGW0fC3g6iinDBw
EsqdZmHvDoXBqHw8rn7oBne5WRunnYsCUMxLvf/YYwVdD/LQo6psxVCoHBlcZWCOlV/plmiekuRw
doQkOaLJK77IqF+ei1HF6sdU5oPNbuO1Ey1AXlKwnG8OVKNCQpHGOMibw94v69QzL1agwFZ+/sI5
NwZUJB7qJiXVV0Rm50a6mSyGmtzgbFKtT+xq1+1lRikDKmcWA7fk6ZTnsEtcnZUvz8uFlDQyEqis
bfyZj/abqBXR6oKWdEJMdn3p89YrFxtP3Lz0CyP5Tnn2yB4NRXsfiaPKWgW2bdThi+9wZuEANx0/
47CneezTY2Ewmdsvzl6nJ/GvUAnHvzANg/7l54HGWb00T3+dQ0ovuZ8+iHoD79xbaEbbgXQZi9Et
yB/Y5dv1F4prswYrxnMaBKV8z4hA7dIP2cR0PM+xY85i9ZPAbvV4+8jreYLYB74HD7EF1fzWu1Gg
ErBU0mb4cICJGMAHh2wCFQRaZ6x2cBgwBKypJiG2ehaDsVCexAMrwmKqPvNJE8o0g28KnX6enWqq
Qvqc4Eyv6XLSFSGZV9T4GMfrefrMqKlyPuV90x3OS2s3VUzFK0vatJdb3vCJ9W50nSwHTClUKZB8
EZh2hiZTpjCfpIx6A+CKWnikKJXepuh1nGuCcJ/bD/Fniy73iJTLaL3cqneC9qnhIqiA56F/QId2
MLaFVj4Hg52VVwx6vTNUf8xTsNs2y+lLJOzIR4jmGP5ZLxvH9uKwrTB4bhZMfDEPYGxCYOojLNGK
S7XsX73PpiZUkLrwEJWZDj02/9QrSmmbYD6du2noTzBZbY6ch4DERyRJIeKewdZeMP4AR50lQUIz
Nrm2PVv25bXHhv9wzVnli/ggIkXxNe4hgjL6KzGRulACR+kR/4EdZVJF9wJ5iw0Z8xyXU8x5egUF
b3UQqCrY78Tm/fJ0pWW2dmuJoD9c5eSwFnj/Epd6ULbyG4O868O+IAhkQLbIDulykXLKSpKmtUgD
Cg5OmLZu3Ovo9peUa8ZZdqEGlWFiIGIQzDJhNLW+EJgcY7aIOAgGPmxtX0snWLCs8VyvwcMRsrP1
+3ena61/4kjzkP/5EJj5OB7OoGFTxdEoK+suU8hVrQEJOM4nQkMLhjac4kbUF6g6XlzrQJGSmsHM
lg7xa8izAzRI9fUhSccLBhdMiyvn26TjbVntQfMpLE7nSaSxXBIqmh6lwjzwrLaSDWwlWlX5KS9r
YIrd0qIWdi2fwaWngFzYELRvzzq0HdhbP6HFLriY2OxLeZMiEd8Mpp+QF+eu5AnNOiyhXPzcycRx
0ADzS7HhcCZKYG5jIhmhioVMxbC7AvrrRB4bKIYB0AKCRnAulMOBNh7FEFOqdtjJxRLpfQ2cAdDq
esD610Kzk9xi2wuGBJj0fPHh0QNjppIWK0N3iTqQn9iNortEbxZxw6Lm/bmTJQ2/JTWI2ECl6ELj
5U0vvnyxZWOpTCbKrsqx0PMHvhA+1LKUjwQ6AGLDN55n1c0yGZOywR8RUbMcbH1szx7u6pnXNxul
LgrqDYCb0TzvCIPj8BCgPh+jE9qHWiCuphzsNbraNl2ew86RiCnWU5ayxmwd304hVH0kJGMssaRP
drZ9VH4jbwq1+eT5BnniM3R6Gyh81NrhGD/gQXM84izLbslU7XGwKBLlFR4Zqpd+buDvnWaNBJcY
ypu/igUQovw0A2UDid9f2gPBMxC9PNN4aczIAIWmbHMzHQtpIP4lyEMyvccpMQ0zNh5x9ceNT1N/
uOoakvAi/3yEZfjeaH4Tqm5YbHpat9i0iE/2qEN093PIX9/MSk8BfdRi3kQjhE85QhLgTgM1nnug
ZwRPs+RNn18iQ2CwYpX4QetR4taDgiQeIml2a1GnNEXr9lhLZWVmaojdNK59jQRElZbtZhRcQhmE
YUmqbHQ2ZcESNI3CFSfiqRSbSeTHlXlFSeMHj1R405m4RSq+3nIKw/rDRDA1bGZJE4TUSKTXnouW
j2YHKCLCw3O+YAcWS6s6TzQm7cacMn+k6sGmhmA+QOmql1+ZpqEk5iaiKtabrowC6LCaxLz/Myek
OBE22akmEB4j+2CWRDKlPn33k7xeTWBmJHC8Kj999I9FF/5c0rqZun8wNRxuUlHe4O1y8ffZgZUb
g6asMSkWKr6+hx6zBtXV5OCLPQANOXyvbwFQuzQL5a45rUNBg6ledzvxbgzFwUaAxOTBhnF+rc/9
0rclC1tV1QnHkeHawXswLtH/XyISnRNUk5ux8T2wCaIAUIWfVDQOw6TKuAPJ9Gwt54gLvNHDqNkv
aHnfy9/y45dVxuN7LC0hZ9YtEP0sO309MEs3JKpAXOY/bZpTCtxDxbZkH449ksgrxi0zqreO3x1u
090Lu8X132Z9hBvOPHTldisaRp8RNyfdsw9vvzk5RNd2bnpqLpqYlY2uJtn7Pn+G3ZxxuuK5f+vq
cR/LRtxQiznlt80Ji7a5ZRdA0Xl1ZLN9GH1qMbQcH7AmThc7rzIF0KOvB1uIoDvnw8MgGroF2D8s
To8WY098VChb1kALgQ/EnIVx/4P6SQrBO1VZxy0GyRF1q42IVrRTV5hymifauw5VzdX3TED5cf02
rpTEEozL0VdxuI8+s0HldU+16AVPihLSCRjcBaKCz/r90wK24khBSruikr1U51WJeC5HC/fAkLQ2
NrGr8/RtNNikv/DrqpfqFwM0z9mtJgmtrpEsA6YCJiup7QXYRoQCvJwDKv9J0tj9jDV1DZL1dakp
tOT47BMteY8XuGY+SQXquzb6HkMJppHH7PVWEdCQmIXvtfktYoOaPWo4lpMuWvdiUc7cOxO15stx
HqpNEfeZXzqXVH/TAe3y89UPwxIIKrAhAQAgZAz1f3Dt6N5BON8Af4X3Q1rzX0VnJC9W2aZJkO+P
d+rxhmrsjkWCPmbZotQEDNxM0hQzfEzlFVleHvIDZPqDy+q57U8wPlmZqwD6kvL/VcMOeVLXK4D9
dEl1dX5VFdsYHNTfNL8T7NIMRTpjEQSWeXtPn5xQzva6wrsOOkUWweksZAc2Tj+lBm0TbZOTY4BF
yEdENRncB7XCUPNsOa1tUlnRI725ymL8zt3uK8RFxvKFetZ4UVEIjScVhOGWycfqRjDCEeOpouJ0
dcjHdk3Z5APlmVpzsbg/4CkSOOIKIHvQ73BW7uMTetxz998GSLkCUDnkATnV9fCMXhy1I5fXULUg
t+UC3Jb8w45WlTZFMs8wI9HfuxLlNKU3dvO8Hp4U8WM3YFRg831EhB5ebEyGQxpvBnxLv193e3tS
0Ol9/wVvd3NwAVJLeqVmuDQLgVm1xJhVPhI1h7NkfKf88tiUDkwBwA1LhOlSDc2AunJR4w7Vc4Xn
uG1/NDiBBVJUg/y6Gl5ti4OlGmdxcaompegVmBmk6Vk2ZRVEe3+LFnARJb8WPd0hn2CPv7LqknQf
1nPFCO7dbm+Dz7/Jf4BNxOOIoLYcUcNKXuO/SZvWhWRAsHZY9YhlaykhpJvmHkOTk8RXUyI7af2h
+3qTeoD7Lih/VYUwjatH/EVKJeTZFnfLlVtGkounhyspBbWkSafUlseNBUdyT5lcd7gOCIYdhMMS
u54xCmYhPOjG6c2ppQVN+6kMApV6cY4Efx3g9zVhaYAm2GeBsKr0pn92bxtYwfsQ+xx8ffYWBvSf
tSQl4MFcz8s7qfS+EWi42rwqGNsoLhvlD0NpfCT9LYsqSrapbEsd/MzoeVUtkTJA/0sisJECRFnb
bRZzr/P5m7qgdj1mSoRCO9LaLizoOTqlkKrVpAFOfb8t/tjf4Bc8ehMb+8H9wzmkxZtrrMdq4x8K
2XeqYUIdHJiO9HVlVOc9yKnalEqWiDsZx4TzE16X+5yBWsi1cUanNNBmsezEL4GOJfbuTLTTwDKY
tiSh7sQypotvUWjWIJNKCB16AdIBEpJW4j0qE1jz/N8ChgflhHdnlcD9baJ44hwwmcqtHV5yrGdz
xkp9eNOPK7a+9x70Y73EnEKTrWuh7g1t09izz6qENN60BsFWjOElVQxGXS0QPyQN6LXCC2T0BDeI
s21NDchh+tSWDX/B546tlauTK3dq+UNjBgyMdbyDiyXMeR368RZViB085NkZq/Boqx3Cn3DBPO5F
IzFspZ8T+fPxfS4GGdY5IFEEf7HDF7IRD5Wj7TOmR74pbr0jMQaXlwx5B2iqxdKsEyWokENvVubD
jgu6Ga+QGVRFXO4vzF/f0RSmIIA2/CTiW5OVYF5fPjyU+d3KLzD7gluhSSMl2nHA4j3dD1pys5bd
CBrtpvyJGDJdxaZmRmgKyVldC8Whr+VNJOpP5KNFO9uRMAPuGk1KW8E2bDn/kSbpXNARXBPj3y2Z
u8Fb891HNlKdS15Y3LCItajFR11aCHbk2Cvn8DTIrkT19NpPAPoKyo+a+I1UqZMswjHiDVDi0P5F
4vkB6xBV6md2v76dvGKlOkJPNaVLitc9cO+Vz8hb8lq7cy67MoAaHrhwpFqKg4pCFCZtW5Kkczdg
4+4cvH29vswh1vgo//8bFLmMlMGItI8XWtR326ifmKBiKPVKIGbRBYW03xtCxqQ50VVB7dWR+ogH
yPrz9qnNIOvSJqcWVoUfU+b6m64Pa/KcSuB6bCwQ0QVw6K4wd6TId6SOZ07hPTe/lEtr6qAKSzMQ
VIbXvHIoFya8KzgnnXkL2uKu/+B2kZYvqTikaJv1qSWFd8SlXbUq1M8dKb58XCTp27HBQGrHl6wp
VH1VT+12Fvepj18fNk94mqA7dIBeETtXEUN2LwMg9dPDRS3tOBp6lYv4TyBg7aoVENkey6hx3hfT
CHVJUN79SKXJJDZMJ8cJHCSyjwc//x5VFb3Puu8nV3pVy03r7Vpa/2e0mK1pICtgQmnxeMoB2ysp
mHdANX2++Syi2bew9s5faMrKBDIQgrC8bsFcZV4djxnn8tXvizT9D9WoaWq4Et8/zA+keXlKeojL
zo8JF0mOMSguVmwVnG3UzHbsz4ECgtW6E6JPx6mPtGDfx68ufOdpEfONTGcuOySgk4O9P/gbcwLC
BAlFX7X2UUh94M70dRTGdqpTBEH33j7tSzzM5OX8IgXMNOjWdMH3LTEJuxQVchndU2InlRTLGHMw
NFRq+NoPRYEYBIUjKElPatqmFS/G3MH8bCkURbdUsN2A9v3H/1lU6ZVM8Nst1uCmo1F6B41oo25E
czouHUD9psDQ5ZWTCzB1VRifL5WGpVSp05RUPOuAyYIpzq/3t/1ZT3oDVFuqF4c8VyVC9A751bEe
uYautbcAJMM0ZFG9swJzvfmhMsmKHHZOjFE7Sm0gQiocqRC2Oc1hGNRlBHwE1rhJJ8PcZBP2ByXF
uw7dvRHrqB9pukTGOoGQIBer/p+VNpM82GNhu3esWLY+38jUWguYJ5S1UpTgBjfxInjiqz1uu5+8
MzdJ1+H9WxbcwliafUbm4eLvEXdQp3KM0zwO9hUXFPQOTzW/CpYZBF7q8Akd7zkFdQY9ynDpEIJ3
eK7DvcF8WP6o83PaEW2qigD96i9zOxjWP5MXlEouxoH8kSiFcOI7H2Aa8lsOOfxybah2TA+KBo3n
V/y0lq7o0gUqrWNs0GfBbA97e1nj5nnlISYFVaA2P2Gy7+/xvcl9CEaoymxCDFqB5rGLd1kP+YVF
NUV5ru4mkc6FH5NZTWCfZpQgamAT/9XyQUv764XlQRjHNE+d3fUlXFOl5EA2jn37KkI2x+z1d/aC
n6WJOLmADjVUBrW9btdFjW5b5+ca023svqzthc3yAwcnHds5iSIvNjnxMOb1OCqdAydNgTtCLI71
TWinpYJ9JxPih9LMfhVkzByVEVDB794AwZKkpJKu0KgIYjBd10AD90OcJgiQviZsr/9n1LIZ6KVM
NC7sMTVS9ZCSjll1r/K54qF7tX9YQWw9q8ZnVet7LLEjlDLteM5ugcC80xPP979uX3CSgGdafC8b
y6cPxY9e4rywPNKdcHq0B0nJd1pdNbFHJTcoD38wZknaV82gs/1FqRWZUKvDFQRUWxIpPRk6NOpn
V31j6UD7qOpdb957i/EVRgJdnwXMRjh5RaJl3NUUO28ZSUAsek5ZtPEs8N4URBfyf3i1BK8rsH2b
kBk0uFSDVdWzqhgpHlB0NRTWgwG4UZEW9LLabg7B90eKrvpYr6NnuaAK1nkajfprHo00boC65fQM
5DJ0kbgTLf1sjWMiHrhUbgHikEK9ouW7bt8YfmG6leW7+x9FDrDJ31JyIeaPa7dkP1RfeOBN34Kr
saW9OFIXyvHVpxkguiTrh5QnCsOqMfMNMRAh/4OzLgFMIXUfVdO+jK5gO1KEehajY99dPCRbJCsi
GSP+qJ4DWyxbvnePPnAGURWwDGAldOR5rWojh1URyE6N3yzrZk9L1uNqLR+gWfWz1/OqKlH4Zvop
GZIB3HzDAav/zQrhNX51TXnhb0I2SgQVsQ5YYOnVr/BO853A3dSgYHUWO+JO28lHRa10hKGS2h7I
twfDiM9qZwdDCoor3Qu1yJvkOT5T+5TFUO8d//YvMNAT23wR8a1XjJ1TMDrJMUi69ZjbJ9ofxkbF
GLJUQeA0yxrBi0EejjxON+90p3ST2KhUhzn3uR3BGVP1qhdBYqyDmEVE+KdjGlqPcdGscYaaDZgt
D6gnRzTWtGoGhUQd6lwKl9YdiUnZEwd3DcC9tXg2xlpm7col+sL//X2hxz8tNvdDw/DQoGv9+CgS
kS7qyIX+MEs/uKBVFxVJ6T1gOcKwl9UPuFNHb+MADtJZPe0x0fdGklTJx4DUYogCZWNa8vyJAxel
K0aoriEnNnKiAn1LQOnigsiXbcMDqO4KaFoTtVAER9/+yukdAiKZyYlOkrnijf2FSpq+dgrLI9zb
wadrl2tOqMUhwGnNhbF/aQs/BTqRrai9GhwrQ/1u7A7tkHVGgRHwBI1CWRFzWZLiMsmi5Uk9u28L
1v8J3o2Jr/rlV/J+mjAUQNxR1DyPGH8vcjWfF8fHkXTmHQ66gcVZzW4fmSDHNYqiD+HaY5kYoeDR
DEWQu076ODEeXRGr30j8zmkewNUXJ+s7rtirUO/BRMd4fD5heUfZ8eOOHyHwuz9Mc9wNxM930dUs
4NqalN2Y2oBIjFRScWKwDYjOj5vM0s//BL3qO0eGiwKjMzAcms2AZ0WCwlkkV7/jccsY71kCsgHB
/IOLXdsm/f+JPnAZyXy4RSJjAPvlMwhMwMsarqDwJdDCuFt5xNAS5bMfB0mJbcid2RXz64ffFCC0
aLGx8yaH91cnWxGzmNilwsYE982AiqTFGyERyzSzVjVrVKAJl/JpXLLo4+cEhonzzHfTqxG99mE4
iTtHfYWvjJ9Bzw/EJUWMUnvLRtG+F+ELernTjsuDf6Mkn9bY/m7vQ2orguKd0nvpOwG0Hi8rCoXk
/Theb4s31+shlHgNAaIq4rtGQqH8GZngJshclmTa91GDJAXLZL1oeN77iMZTDK+bcOiLY1B1Vjct
dhnjlzEnfkdxh8bRFSOlkusmE+H6WTXCOA8eF0uHSBLSrsTaoXPAEgSBxydz4yyqX1oLa7O2TMTp
82n3/JGcWtoV68ekQ5qpQezF/n7RGk63SJMfNyRb6dX4F2ZD4DQ1/LuIwcS8QqQgennjmsM1Sik3
hluy7nXu7jtIlMq0u9LCjm2tTUBr8dV4wQB3xM9nHOW9tiQ4HUekH6Vm4NReGLo2JWDd0VoAh66u
R7UTZfmDB53rrWZatFqiK9e2utFW2ghIpenpLn1ldZ/zWBQssdGwEONb+fK3YwusC2F/bSBuGpGz
pSQVEVhf1lU3b1uy/p8TECLVMydbEJtHskzGgxSlDgaOWq8koJQg2edSk0ZuB3RP5IV3D4sFukhy
D2oX6iBLjV2bCQXJzmd8Dj9zoKxl6OVr5mRmhLGkka9fX5HqMeiiX1Gm41gchqy8aAI8REROyU+y
5XvcsPTko/Q2qZ9gteCuibxkfAs4dYBMbmCopboHDpXI7vBc0HP30/OFmj3+c5PxHMRbZ+F+OB7J
+FghjJ8vs2oNVBOMVz+ZjWx5RBlgrpnOK4960xH9Lh/0anEWdAFukjTkGsbIHJxg/mK72XCe3M19
cR5yFWQmI4lPZQUtvRP/nyntuncizT4TJ9hakkPjc1laskr1+fOL/sSGTpVS4NWTs5DHys3vW9nn
BBrlfKFTHzTK+oXbFHpg00FJJgxqXWFmBXZ0x+USgIqA6p+REmIn6sZ1XJ6/0o1GJin8b63lMuJp
sUlselzLiRD/D+B2A4RxhZi0VlB3doCJ0YmtuUeS2fvFNmLHHggXDzIrUY6YAYVkh2qy0AmCwtHx
muN4iy4dfvI8nlwzRMC1aSJ3Wts1fKo4xb+CgL9+CTE/tcefBnKNx1KI5JndQcHYNtzIaEDldb25
duMbWPK2vnkbaY/N2KPnXJzmIoyCMnRVdlzbISvoX/zXiLBmffc76vlrTilzosm7lpUdYjuYCEpP
yuu4U1CyGQ42pSvNu6eBgaC5EyV7b2lkz0XblTmduTri2ubN7/8t+is+WPZIiJCi9+stPSOX+KsH
9HG2N2DtbRzrnSnwwvqBs6c16zwWvBF2jPzF3ToBTg6hpnX8oix2ZIKVurikXqRUlCl2mnTRlXWg
94ZaMXFVsqmwCOYmbxj2SaMBimu2ewWIc5bFZNwngxeTHB4G89sv0vsMk1T/OROnNEbaA/MJLjVi
RJtLkNKs9uR3Vr5cQi8AVYDzUXT07v4i5xX0aeUjty753oFduw20Iyu/mIt6l+gKE8zSUrdEpB40
lDaTceXoKL0Ne7vnB63ikgwIzIssuw99l9/Cg4KEZ3rdAURSniLiy9CNqqnC/TS10QrUUiS4DUzr
VP7aiIcQgurDzyqCbsLsxSaI35ohN7LaQQ7jRNbRxq+7eaRVqGrjW7cJ/QV0ogId3QXnOJwS+9ty
UkRHWxduWVXHEJ0eKFEDk+75gQuYqB2Bwhoclj8yHjCb8e5Pvh44KeIllurV9hnA4k4pFVm0Z4jI
tPBk4bxGIzE9IMJdBkWfeJiCi3x/JJ7dyO3N6LdqJS64HJSMIz9ROz3A2aFM4BTTjykjwTSqnG6F
+xE9lTsMvTh0RFkuOra3+08ZqewEVWmn44VVboVRQSlTl8whCM3UuhUVFtUaN+m6mJRAoGnkk8Yl
ailXTbgkrM8IUIKuppdMKm3jri+YMF4bU4oNbGa4BBNDjyp46fjl7SThbtC1OXycfgxoFHFybt2P
434FjQdh/RIdLKfw7cDZjFsSYJxxjoR2SpDQ3v5+px7ZN9shCSurP3jV2mXAErTZ5lUJ8hEvZDyN
3m/wP9IyaP8YCQrhX0mT8xKpT67ISx8XIWnFt9FsUwnX2BCxWvPbXwCHA2DxV4nVrCN/nK33hFbG
puhKgYwQoiEGiEvNV+u1eT593nUzt34fcKIAKSIySCRkwQQ6aDoCvBmmB0fOH5Ykfi7OeovhmUUE
hdigP11pxpBiAIIz89NKchuMzHRPCjMd2+jSr/H9Nrs4zmjdxG2hZYKrp7owB1rU3ybkWK92rBz1
q5HnBw7MpdI6tXdaskpFk4Qe8VpLjeaavt06jhZCiazdF0QJ35rHnylKtPhZ8ArNRQwBF03fI7Bc
UZ0w5Smo0cAAgSPG7rioLsDEYpy5ofp2KgTDU2Fae/zYjDnctvJJhYWHOV0jYTeaxCQ25AO0KZnG
QNfeZY10wDMnVDyqMXmeFYcXT+mWaL09Ts6zaDHd0zrADYVTiIcx8QZGkT9IGNy8b4XA8/MYhzSV
+vUng1/Rsju7nS20IwRX3N5xUwtwLkwsBN8/vg4Ydk806CsZXIXDi1h8Ca8d8Bq7oi/DGOHvYRLC
2hiJULhicmFt645AI4Kyuji39PMl7z4curQn4W/GPGPl+jN5/CVrlv0FGugqeKl/sDVnMWvUhvsg
UIL9OaXRJTy6a04oRa1RtaeN7LQiv3vMDoYxKNx/nM9n1vfLXXl1Ys+V8mA3RAnWl4kIpkSV7Vd8
fikGfU2e2mYiiFQdbJ2iM9rMO7u20LJ5dcxRIFbTstl7/XqqJyopSwm7fIDJqdo4uwEPkW8CfiZ7
CIhQDRpytnt5UmJtghwYtESatYgFPZn/Bb58l1iywbNxuKW8MAC8hgU50BGCip9EOpl5i+mHOrV5
30yfYBVXatym7pKzapo6ZOI1MXQHwcfO+W3p0+JKJgiO2vj3+HEy/F6FJr8vd3t5jEK8H+royM3h
hvASPqfzqLcGU1EodqZA6Ig/qVl/64i4qQEGzhMz4eY5baMR2HoRgYLLbmmnDyblOCSo2kR7dYo9
7WPMzx4X2MMN2Wz665x6IgVAsvrJP+FOQ+KoZU9SfnVkqUpqb8EVbaKyu8tDOAlZS0lKPrvJry2V
uaC4HM6/3pVTmU8GfVFU1dy7zG91XcSsxFdfpxKYIuUDJ8YkzX2UqliM4iz/OThPfUmdz1kMVNGi
8x9o/zXRr1lNjc2wA6kM1OZ2CEbg3n0PP67nTyLoI4xCEpet8xRrUZ5yygHI6fWhnJQehUNbCZJh
gr/904Hy1oz1UjViDsybVdKMD/ogXujH93l59Qzr/Xi6OvUMccXVRHBycnqh/K0J6bP++q2xROU2
+3tt+0Rdt47bht8aLy9QFYO7E7posOd5F+GFeeauMh3zuMJC1jI8Duk9wGK6J/ExR62EkPfKoQs3
kADJBcgqwwvYzwTTSPdhdY2QMMLUV73fpb3ICwe7Ai50v+ZdfmWZ0Q0Gix5cDMjwTCzsdn0q7KL2
TvPyMzKGdirliE48BhTyl2C0N7IxCiRp1p32IHx93xFtLhTrbpA+M1zE+Om1DDD1TUnfbF09OEPk
M3G8rZJwf/7tzHpz10B440mz+pf15DT8I+79lvaeQrDpUO6vKZvkPJ+5pCuQc4a1H/Pm2yq37H/2
MSwX5rGr8r9qHL+sw+07gCJ9mfMw4NzC3k62Kpk8+Z//4ewziGqmiSY0U+SFqPHq3NZxishBFlSM
LYgdJ42ptgQz00DitU7src50tEog6kqTOSXC+4HIUBzNpp/by/JHIsAnJfszXeVRBrfhTl9YJvH2
GYGu6m4ImYVZQ1X/fWheE3HVoiaOKYAVms3kZjcIi5t9imAi9CedHTJPPuhARA5yQ7WenzxIDkjX
kO6BzY7dEMmtit1xUO1RdPk6F4W6CEZLikzV1fHW5F/nSSOiCHD9M8Jx1063KUzz+Je/78tlpada
Ctb8dCoFiGxPB38uWOIoo6bAAYhkVgODHRnModbnUNcXKKK75ej05/td0tTOOwNvLApUHpQQXA+l
slxeML16bl4DQW1LR1YzBATn9mpevP0K1gRxmDjeN2Zd7IW2WFmMBW8hEHolmi/40H060PT70o9X
FVIu8UychtpxB+JK4vQrD7OO6HPfE3b+H1oSffd9e+Q0VzaAfU+HVsMiHRTfYzKfjvYCU+TOu7Gn
F0iVIYy/fSPL2lDXMEh/5IbjyvTqBtgZjr1YUkganMOrkkI+llHgAaeobI42687DocrCphT3tkYH
tbtE4727E8w5zOzkLApUf/0cbOdKqWrPQorkBDAlfosE32Fma6ox7n97YQxkhozfbAUqJ5EanNjn
z1F0KVqEaFtbaa0eGk7dokzVfcDYd97gPpCNW1pDhPhL0jx5H9gUafN/RmBlsjP0K5MpE0wlJ02k
nIzgoUUid1mib2QSna7AcDJlHJdkoBO4VufhVvLJc3aZpgYrwr7A8IcGmLCoquNk5sCLMBtxSw97
24mfqKAl5Md1Kn/YJmDvmJ5OYeDrl+LurZWic138DuSwLgzGBq63beUjE2WOj9CT7Uxkce7IQwPd
ZerHArsXlMIY81Lw+kLnPdjsdIRSsk2tOTvjQ0aSAb7uLJxBkQKpTHRmtuEWmcje1KVKF0Xz3S9r
GyAKobgIRWVKy+bF3lp/dU0I1JcNARMhRkGsMbTsetf8i11NIyfFroYUulD1/1ASKCa8UEwA4hSf
6sdbqhhs2zPbDEg9Zfn6+Z3J7mCtvTOef31CPUsj9ozbIEtafNgCUkIMcWKsg+oVtizzkDoUcBmi
NSpOBhRnkp+UuiSYo6Q9vL4gheF82Mka/d16GiQUqXzEIjxxl48Un+u6AD+dSsNMncxSa+wdL0Yp
mDODT5b4fnCkcH54lfH3IeoNQ2Q5lR8WjCKlnUVbIRDFNyLNx2e9sOpuiPX/+2Eg2y+bUt7+DIlf
WBVpBuVjt4WJaEcMFy3/ARBhBawW9Nv1CmFKglxhwVCUNO8F0mzzUqOu5KzSuR3ZSI0pkXmRZ2LQ
JRCh2cNCgGdICe0WWBIgarHg2pIKFa2qSNHU5HK9CB8140nPV9p1w2f32idUt5fHm4QmjQuRk+x6
vzTXWvSBEE6SZta9WHekz7IRxGvH1YhBMZcwwknUPJbwq7TOGxHnoQACQzKJzHead7mOQ0qET1fk
F0dg64G5iPKj4J68czoVCj4C0TcKSOUY6V9UmLiqaJ4pKr/JkSxdrOUq7Jph38TvnhktZkREGV4V
xxFajeZdju60rCzszNmAWbJJJMyDCUvUKfDlpX+Q/2Ua89r0vtYkGo4KHrhdZa5PaJnuhGusBx5q
EeSTzkzTB0xKsflCtq0Xy+jgKJOeWoP7wFbjtIUAgReuYQN1mJXszWEL0I76eCS1Qia7c+Zg2pEF
w3C82K7xk0+j+lQJ5JlQbcHm1l6GRcDHor7oF7DCev5FVQJwDf7jlfKhE845fBSgUMdEujvvFKdl
YK5lX6jXX4v73vVItVxkagKQXDUiskdedHdWVuCpyTUfazaNgtBTUrF3DK9GBR8RKqhUElI0Xjm9
ftiwD8V+Lym3/ZW+m8dK7f2DgbNCmg2SU3nvjhEOYdCPpd3gG/6qSkbETv5g4BzQcSRU7664DpRe
xnyZjVRF1GoJas7TjXps++Gmfnosp0nBjuwus/ZhNzOPQlqihRIRshaXJ9U5Iz2VEcrn6NzqCegv
gkKF0o8GJRqAEILN9ze/a1O+H+pepQWty1Lu+1ihYURKFAORfkh4TeF/NAVNJg5ShAluDPllIIkK
4NVu9tySlW1tJ6KyA4QxMB3Y67aIiqKjW9neTi6i82e0keweFgpx5b8u4N9XI2HCErmx1dUhaXHv
k9pAdQsSlePI26E8DjHEHw0QJx1OjXIEwYj2WtR2kL7Phrh+UzhQG3v6hwx9Du337fQ/6uEY8RMs
VVYAORD+Gn3gUpb/CcEbE4Su0XR2g4Yao2ybX2v2D7G8h0NCGGauPpOuqZKMqlBFB+bAJ7gKTjDR
GshCTP1ALMzYLbdofgiR6VBr4mzpcf21UCknQYnrhzWi2a53T8dOrpaYDK5+1Wv4Ej3SkuQtBqOF
6W7Ibq6gsXyd+oXWo1Y4cxcy37U35/dc4VxXThoSAHxt/zCH0nQEROeL5gETqzaXaCXGLOA3N+ii
807GfEB1ZUpIo65WaHe+AZk/HL2JYCP3kp6O1eyxWiGT00ytv3ywhrAXCk2bKkH6DWiugNvejtrO
p+m6zPPEAgnHSvDX2W8eJ0+/whhG5bdsH3Uieb+KDGnA26rqg7QXwBHEI+u+ju43CaGPKoxQyq/L
i3Vm+LkpDEjLo15MRzkm3T+3QRoUoUMHOB52H6kv7N/7llU3wcrKtUB248o9wkMHirm2/Fldw0NX
QkNFMJjbTsQRZinpXieTZbvQUICGGtoJcqIR9eniWiSB6zuo867McQZrV1Ccso5s4dnnuvBqS9mg
67HvEANp6yusIBrAwSSjsnhmPO3YyGf9jkTHNYurNgmZ/7ilYhMe3N7MljjKqa+QTXB4jKgPvKgO
4slI8L60MwN9yV2sOkFcfQkEqDR1vNZzb4Op0lwJRa2DFwYZSwglqMgiHHQMXDp+7Es3PdjujcYR
R1CVMDvUTR862v5Y0c8kTmk3S3yFzsxsxBtQfLhQZk3UN+r/1GL1wrWK7hwSFhHJJItTa1X086/h
t4xULnBogouQf6+p/pOUwz8ltO1Pv3Kpa+NoncPj/N6hnh5nytNMMWsjO4xhvNVEwbwiIwG5+vg4
NeRccmmHXDdbtdMshF696vy+oznufEPQm1p41ubEgw2/7KEavbuEucaQnySXMAXW+HVoPdF8eF+1
bmBcPZsABvxTqSAJvIKzFQJKxd2HOmKvVKeXh+ThvK30KQZ/NjcuIQP2zEqkaDw9XzinhLpobKz/
uFSGaxdlTE2CMepRQ+uabeHExaRgCMQnuSqx+5zNjHdhhLHeChesYBMmNzCAppLULR+YzxeAXSbp
6NRkxL9UpCHbi7RUhama9i0+vAm0qWmzThRrSQzxyI1VGHZ+Kn9TtEKjI3kcskHzr/nCLhm++hkf
2A8hQUThYKACoCOKjjEZ5mxKU0GmtzjZ8II+LxLShBQury0gyoony+mkdZKnyPdybSynf9EPvnp9
DI9llcPrhmpZEyVP6UQ3CZgoUxli/mjtL542fHfr1RmwkI/EmUoDSx7wPb96kZ8pGAio/zT5vLB+
u3kwb4u3AUs0JJH9Gtkn0UnzxzT5tQVbui+jWHSdmJUjYLHJGbqlRj6dVVeTxmQCII6vQQNOZkPU
2/RzIUE0Fde7AQM1mVb8HDR2zga7qru6BILNEqvIrgbep4tEcjV/f+dMCJIx4D/hmn1GJDx2XhZ0
cIjpJSEtLSOnt7R1m9CYL0lrNDi53KAatoa0kORQzsebeM/EbAOpoMpE0geCC9o0jBd+dRs2ah/r
on0+qM3oGGMbvQ4AXqjZ2adHQDVqD4Y24hE93jk2z529yXJKK21cQK7n+fEL4DbdZKHk7vfxe9nB
L4gzI2I1YUA+LnmNwfiNpTWNfkS5VrpE8XwbPxI9l3PWGqJZ4666Amtc31eMP2o+/Pvu1+MgYfjE
bwSfkjfVn3plMLjzJlGyFH/jPfZUoUXib4RnvMV3zxs2l/MlclMlTRB+pBgbTbJCobjxZ941cZrY
u1G7/G+D/x9PaG2qh0ZPd459s92g++V+8gef67gFjnmGNyjeYMDX3bwS3aMbu28NV9OOUbMWHMWn
8EJrNWH0n0+Hg0CbGSuyukez3WmJvteQ+/dsNv46wAspIm7NfZM5rgHKSgPaw1OO27IyeIUw9Kpt
fLSV9q4pyqUC13CB/NQ9uVswb1HRRpx+wIUYEHgXz7EF8Fx1BaDkH+Ls5DSoRfCMnA/pjNd5ZHTX
qUEKpxqAOccGhQNn41+kSQ58h9SCqfXixLAjarfh3KW+mQmfJvTvKzF/6dhu8ICLYCSgWOAe2C2C
PTiKMTpZytyg0uDLoZMK+8zMyYTJAqzJqxsv+hT4VSAJbsP+KxZTnL33IXIO+j231XmYS6tqRgJs
8cAIdOhP8IXtwEwvo3IMfl2UjaPk87e8MCvXiIsznQwGBXwLuC0s2XJfdyzLBEcfULahd3tv6npj
Si92Af5p8opSzv0cej8BBGpWuYZEZWojrB85/tUDYk8TnBGXIXwT3RakJdRPPtDI2ZMghpI4B3U3
N2IUVlfaGuegaZP3+Gw2NnBNfGE47f+6HvfzTpxgELXc6yWDrEL1L8q7xLGAGBWhuq94mX0Bzco0
esnvn/869v7NgercLTW73DrizFrdNWvK9TpcEu/GELZK2P7pPnlklbDjHsd0tnTIba3HPFREIb7a
RFakNPrccoP2yPDIMPi1x/lZZ/F5/PqkPu6JJRhismyesm7QNU9g+ZFgOYMzCaxaXsNG1hB17HeD
JAm6QC/DDteB7TS5bxwocytJr8LXCOTB2aKawxN8JkaPHxc9y6v/qLoFYJFMmtbYGhf3gqLbLU6J
iGec5qGw+uVg3tLCiguB2Noxw4aiIfsqo8riUbWWmXjTesxwM16l08SrkfBuNJYF5Nw09Qa4wlIQ
vY2oviZQ/Qb81I174DcfcT+A1dFekWwVKfjtIpv5UKM6wC2M0f7zF+ZTkGtHd5/ItjR2Id1ZQKmM
bWXCffHnJzkeZ2D7UeSsDhI6ZfLlcg9iaN7OjtIPdI40RwHRhvSehRq0Q0NcB+RKEONBSLuh71lz
3EXtsOClxYyu0hoPEylFoIgJ2JDQaEVF12CqywneKQlit0RwvP/OBM9D9ItCGBGX1UNIVjW2dK2g
NVU5tFJ6oZOaVS4ToazrVirnnJEgxIfYcY7TwElj/RdXz3PuJFSSWK7lUO474AIx2gtcJ4Q/ZxxX
cL/nlAkX0A7hR1HhwmH14oHRFoBtBffbxVNGhAyW7bEzlNNH6XIoj1V2cR8UVDXabBD5V5SEBG44
W7h0kLBEUxlt87V0Q//LnyyW/K46HabmyzecENcEVEf2VLv8ugsK90scfc/HRqOchrDYvASbUIB1
xO5fG7LYU57KxjuDmKd3KiM7+MnLW9bHD+pdgGV6bO235HapZ56yhEn9htobYA+Z4INaZ+jddjEY
zWq5sjAQ9vx1N+3pFhOiE0m//fnHLVR2pvUIH4Hwkh/vy1tSfnTHdMEa3VbWjsO/5pFhRyKTnpbB
qnROzUvOQXHl6k3I7/dPNo/jG7YyaRcxre5VsqaTjPmsPzln1of7RPjbfKXB6QCbIt2jy4JLxlSo
rMnjN7iHeUMJzgEj7qw3UwaBKy8JcFuzQ+yG8Je/yBxs/Bxo/FgmHA0zXLvTelkiV5xs0pLxCYAB
IsWPDJgTGc+W9u7zqOdU2RIPl8T+IwMZnel+sMg6zc6XuA3hHI8hkC4QCwak3lOiyT5uOlB7O/Y+
fhV1Y3rNQwE6RTAsgai0PbhHjDbm7jPBEbE/lZ6lW7M8m8mHwb1zW/g14/ESDQGwwIJjHE6XDPhW
mduG2Uu7g+Qr4x6QDgDDQ6gitITA15vHem0QDvkFu+3ribblj3N/scD4IlskouoNuS/bzqw9I7NF
Mm8T0D9P0Y1KdLcOqYg2lkZ0jAjYj8d3CMjyBBRn3NPXkwyIf2sGaHRbghPSbUjZo/QwtZ28mAY6
lyKufMipgxTV8qy6BUmfXlg51A+vblLXqEYxPkIzl+xPIhBI73f9ZGXaF6WAnfMxFOs6x8WA/VuP
oSnAFiCvsSPsgItBPUlXuK5F6T+P2DVr9x70Wxvr+M/461nGFX45C4ZX3K5VIWhKTVQOEnYDgfFf
rsy0GfJAI/sBQ6tmjvvIAPhkT+FQl8mNqySONUfOZBkNHZG75174HaXyQLa2adq+s6dSPbkKcFbf
vXxux7z/PtfrurVnBI37ZSYtq5Ujfrwk/L8hKQPt2ynwZKuG0ilaOq50yukH3rchhll66ScPkBQY
q8JbnkIGeOf+62aswN6TN4do7av5v+NJyUi0+8xHQ/o03M/T9TZwP92uQo/UhenAKev8EGshx1IJ
mboETkfZqjQGGg2gmZcudzbNaEnBLiTk1VXhDDRIJuVL4ZMUnFqzLLVaBjDX/CfuCBhRfbz5v9jX
eZfx9BHhZTz76v9CmM9DjkzpY36luqhBTXlRyXdlo/ZWGo3L0f3n46oK8gaG6gkiHPkO3K1SM3y3
z3H36kuBcBOqeN+w1wSAqSSVUDsrbI37UyrFcuA/X1klw374t7gi8D0mU9zOoqBk+wi3LeA8LvPq
jN7YgGu/rn5LqcSHzEM+8uCP6AAxrvQm9WhF3pYOD/nPpPY3FgM+5XvSSHzLDgkxDuudiKDCje4i
UOykV5tbkYQ5WoKAvsFpFb8Ik8DA6bWkzFYXgZaP6eQwgot0gV2ZBqHR0FlFfuJmaWRJBL/kogGK
eq3EthUSv/HUrR2KF62X3B5pmqfXpLGq4y4y8EO++DOqiooXA5SXCWQITvQaSP6nmEVMW9Nou0IS
6kxBNKwN1tJLPOXzGvVo9jlFpgl8c+I3RzFzLCHjC6CGz9MXicbpEApudQqIaZoJIQMx85LKapUW
CkryjNp7Gr2fFq9NE88JLB0UiPYtpre4m3ss1vi/Z2ZBdUUmISga+hypiGx8kICtPfk8QTDrH1ew
sYb5ehOIR0uQ59p8kYsZhsMk5LzMa+udr6iTU5aCnECMihgIBZhGueA1f/YLrdMI/vLoVtBgZsjg
Ce9a4atjlXWQIaNk/CpWatv6k5r6x6nobfeoZn/FTHZXNvohgau18Vf4gpFLnxYJxjG4i88smyYx
9UoxkbiYvAndHUAEdoESNCr2r6Yqq8wcV/7hfH3s/VsPHewz2hWGupPrUYKD8VpDALw9ttRUy6+t
TKJspY0vsolmN0KTqP4dollE4BBXbs1B2CS75BtEDMJbckKlP7tho8e8PD6RtS+fvp0ggEzerfBk
7Jvagu+bALomtf3jCD1dBMY52/NCvvuvs/uzYIlrj2DqUXAU1qyIQ9wFq24POaOzasseQYWOh0dQ
dTZYvsV3kfsjebUbKv7HF3t7x6q89D7A/XeIAROzBWPN6JwqMiHdXCbatTMz3+1Av3szjLvm3Goi
FJwywUXb25yLbmrZmObq8CNvva1dDZK4f2WaX/GQNoaTYq1B3mDC3lfRa7fKZt/xWpaeT6W1CH/2
WRc3NVg14GKyNUWSI2Z4eh27rXXUSobepWBuyss+gTUeDUIFBU05Nct6V3easWOy4KIn79EBvS2d
a+1UqOyOeIDCN7Boap+KLMBZ0MYU0DMUbY7/H5+r+DYoWDWadvQLGcr339TX5VnA/VebjFQ8ty6A
Br3ubjEwnwER/j0ZPhoq7sd2puwKZeZbJhR/dD0q2767ulF8u0mYY/NLrB45REsq9O8ww7p7wf8d
xQhwZ79LutQpSvEq3qrTfBfP7919ND06Vynp5lFTEjaqAoMbg2gxJPWWkWmBHf3I4T7P8CVZV5bN
HOW8u8O88kb6rww1JpnDevxhNjU4CAC67Nc/XxbbPbZOjDAVtkBpGGf1iqa4k67hAYkuiINjaERW
Z8RN0hXNWBvuQi3ZrI45BshVsqz0BGd+Psz8v7RC4PJ2cj7fHL261PCk6RwZpgMTyJK83ZuD3bbF
Jc5o9I795nUCII3Mp235woNVR00/ZTecaqln17uhZCORnqtDjUaZVUhiDV/6WqsuLqMq9NzhPyOs
TLeTTMuApNHnUhjOmle8syqKA436IEklJTET9WuvGEicnNJuXlkWrRpxjtCej4k8hdkfdb9kTwaa
zt3+YxYGWT+eNrdWaax/7m3ZWVM9pEK/wFcBHfTSbNB0aUVNEbxVA4K+6LTW7qT3FSI9yhT6SrXH
zNbdkKHn6on7mVmP5BPGtw9iuk4C7UuF+e4TBmsPZ/S/LUFJOTv0SxthJEnNeqxfP3/6pHyW1t0d
n2DPWTf43wjp+gbKLbkAUOESDVlssBITJ5tnflofJTg7zWwrR3Mn2ioRdTLASDoTfFI37eqppXz6
2vbd0jYb919ne0hjTvwsr/On1TCC8xP/XZ8AAFZfbojUeqaiIMahw0XspqrdMRb4PY9ThnWllxdK
QMF1FyRAu9hUgimAEYJC1gLD5SnqiiUtPmIje1sT+owKnupmJ3bLoxpt6Uc6ahR3Zx5mZnR7iFLr
Rq+IZnOMiN0T6arSnCqf4ZKs50KeUbY/ixnCi//KiwOm/PRIl+FPjMe3vUC2NQvmAm+LZ7GLdL+0
kEBqvtZH9tUlPiSFB2E47A3SC5T3PaeEw3UoO78oSRGpWxyrQTWLMWzTMfbWHiRKSjlVUVgmeTTP
RE9vIcZje0ldaHAY2/06k+FS17tS3z6am6pnc5v9O6QaOYol2MuP9zCxROpJs7pSJmtb3EbYO2bV
qX1meHHuGNYRnnz/Upus4gpcTrMcKGc7tQfTDhb///VVfkpmlRTrMbklL/wvUT8Deukz/EI4v6ki
628P4xB54D7pTC34dcyFFijkgeEACrfCoWFk2x3WYcBfF66UF9lQKbWI+Vp3dZr43fZNUV1QBOtg
JmVzfkX9gv4qtT7hRK4bkdbpl3s2aFmG3jEARCvxZYVEeZM0fIJr+F1AF1vUp23jIcqzqoEeSrEK
GmapYUp2PAf2cGpsT9OG6KixpyvaMijQlkIpwnP4VxVZOI5p1i7UW+RNwJ/WVPrPhBkBYz7aleU7
S4lgSMmGPFdDdnu0B3yVF3AYhEBecZ88qV0bFKVfW5WBIPh0i2VqZb8mlvVK4adJnTd+ZopFBfJ3
FrNNuQmtsCLl0sgzRKDNKYmxthFVxGDQlF8PJcS7fsBtCd5Hzge1iQGPZR9JH/4mV7j+Wb2jr3bm
ymxYacI33hs3OJeIhMI0DifbG3wIZKm3/O4qg2TvUPtjEGijOtxyeHiKMSac1xURoE6I5hwAUadJ
3JovcsGzwZUQ2znwWxn4XzInpglZRPVfnFVRY2yt816WLZjk4X6dcgfBm06a/V62VimzJkjO3nLt
Vdoq1VOTXI9rbHIcYGZgZSa5HD53c+I6lSWb5IMH/9FPuJTO93GjLWUsdA31JsQz5NK8nwx/EFNW
E30GPzAYpDSKhg5mguyoflVehckaIcf2GNQVbc3pVlyEbD6OO/mkhJGzPiEXgG/qMQR7/Cw5D+Hd
Sddh76hSAyWY3sfEqHfrkqNi6Rlo5jjPye1sDvjAuZ9RGHRdfJAAxyL2P02fj52l/qutGLrrmL50
G2TmdOqBc8wrCWF7BbyaPqVc1RKVFo+YIji61Fg7dJ23QIgucRbxeE2Dn6+ALvK9I7Ag8KdbIRuy
eRW+UCMGSwCHM0hWvjf2ARScrM6olhuui35fGfY1NbILcJYTlwXGiEIgCsFgYnBDddMX6dB2ya1X
LwEGa3f33ezqAJ4jPACYwTlC65c9X5JeCgnBuIg8yjb3blVwxjpQhRTO6m3b0a/N4ix3+ToVo7wM
ER0O0HnN5mNHF+cjZ5Ivbzvdq0CNVejuTVZRXFV/+a9ER2UChYqzdpIBYRlzAx8Pf1Xe8SR2XEsd
8Vc1TEyQRKjixNyQww6bXRSbjFHcWPlPM7rO58bkKo31PnEdUJZkg1xYnG2bOdymNFEJ/1zYDvhv
pBkNv/vlDxDsl8D8W8EIuz8s/moqDPbkeM76U3/m4Ty6DqIqb9kHqBEe/OQb1IDcsSXsGd0Dwz8W
IEe6hvjb/HRN4PRHEAxOZuid8yp5wG/SGpSUuW91GPQnEyY0KSKSKtNdxkI1ySGr6Fhr8r3ikskd
dMR3C54xoDqDMn5iV9H6neUr1hsOu0pDdOLfVr51IxCRDcxSFIB4c3aBfTYXmfOK/ImqC6GEPP1O
6DmDQkNm/V/MtqBhtFNZVpCGFGozLPRTvzYxTwUCrHGWU+OMoFMpDkMjtmBRH0ZIrFXj32K7VFW6
2hMRfVZZU7WDcXAyeqv8DSNJ46zXlCf8O6QIA8Rw2yWV9FC5aKGucrYk1zggwm9n+znx0zFmOt0f
5coT27qWRUZLouESpbH4zUR2HHAshmA1nA2xOP3TW/PCN4RGBqDLy9Y25/HkMgqpU/HMGZ1do8QL
1I0DQs81pkcfi+rTQlwymqfQPHdN+hhuPxrdOsL0OP713nGj0fAtBqUhloB2N+isi3lsC2Rk1E1H
36B7V/liIe7KjP22nPBERPwXNyXcBt7wQIP0EcwEFUn9ErJO8W/YYBrBydgxxGZy8c/e+xP9fFuZ
/mR4+4EEt02F3NWI18tl93sWPpMoIr5f8dOR4bKiGvS/dmkxWfbqGgtSueFlyHXm+b8oGP4kqh9G
7hf7lRhg2Kh2b8fK+qdWQtkZHgRKIIQmN/zAtdRpCOx8vnMCkIyc0tJFOV2cDbeW9wpzNkoNWLhn
ZH6yabQCJNz3s+jIFc/h3bG8fYsI9yyJPYWHjtB2adZTfQXAtRjTM6ZxOcAewwaQYMbnDEDuggJ5
7/zJdgwWMgZNsbo9e1tkkUi04lV+5UIw7wCyrVguOTxJY9xeqz8vEDf1OTsXJRPPq+0irsLdkaId
2w+N//FmORZwuc6tepVqHJEQG9yi9irfvoIp2c/11yloho0pI7FNEKWOOF1bq77KgC4rxhibJuvP
MF5OSnTMDtwzF+CWLR8gTcX19Ou9r8mRKdhS+NdvsrC+lPjRUAswdg9X3PBdUhJUmRxJYCHguwej
qx2S0dQZo6K/7/Irrkye0Qea4jq2MxTrh0+S/W8ZV1McKEtGk8zsKCllu7/KTIRiBjecOojC1pLY
ry6jPvH0Vvj+Vyd7digrElKvI90X9N3QDNeVdR4P67ByVIlIPkze3OAUlrV5b6wbr4dkFX7vXZQ1
8FDQHijqpbTH2kMYAagbNfgA/97iRWSUS89D/NIkeRAAE9JOlt4AHmHgB9pHQKkbOsdWHs+pYf45
fpmjoCn654oAMrCqryZnmcizV8eLR3QYQ3Kzb1F1FvwsM3Plobn/o7Rq5nlWEf8UlqMHXwjFyYjx
s0hWCvJWEWDVr2mgZ3yCS5QElW5Inb3BqQcOxw3S+Hc8qYIGHRvgSgQgZZDzLeFXoTOcHIdeKVyk
2fuJGsjJwe8KsonyetIsKdOX0OC1ttTIBsoAOSLvNbDbkVjFN7AZlkdpOuYz1YGJy53eZU6/ZkvA
P0utvWVv1amBHgLLbLAEQfIAnifb1634+sLCYfY+LP7AYqtp3nfZ/ONetkW8/BOVOA4GpcKRZ5un
XSwuS9jK8z08wwF+Xgli4IgdAhBEo/ihc1kupDq1rpbvBjBVgxMJ8VVoHl5aRMd09utH3z7upbMn
OYrF0J56PhBJ1ry+fZob2M1GzYLwNl+aqvR9bO7F3Vyhk4zSpyZmH3eG/A13go7FgYGEN/lGpXH7
LaqE9x3mqo77Jn2BjYyf3VZEb0hrQl6idjivyESnHbgdSFStYtHIxjWNdsfQIEwTR/zTkW9zqhf6
VQ9QX9B/6IfwPV/pODKabuVEN9CL8zY+bcbUI79enrW/irUMUOQtl9mbhEtch4YZxZjPtZlCnioL
6n3aFE8Gd6M92TgrTe5D2aX7gNhoXxRrLX59PBvviokWaVJYO0SNsPPI9gYIXbX2hyUvYFDKotdk
VMMGaA1uZkdTGrlHHE2b/etrLiJ+9mmJ0ezR8rEjXtVyI9+xn19YTGnoHbMYYQJNu9PJ/0xzhOZe
lq2owSBegHBFBX/uLmy97Y1ua6tNkbkQ1oT3J3klx7N+EqoOoO9wjMTnyr1ylkTlkoZK84oClasW
WEqhO8me+MDgATfFmsBmBUzNGdHJECqDRp+0lO5+Ht/Esl+42vw46Zto6psLjBDBP+GfPJqp6GEu
FhjLAn9r7cgeOLFwzDTpz0bo8f4Hd8xFs+BEs88jB+YRF4d5Sw42+PXkIvumFcyfcoQR9c+FdK0m
NUVY6Vlu9MQasxoPnY67oUX1t2EHbvHkMcfjiHgj8VGYgSVQygLqhUkrPQkgtGLYrQfRiEiw/oDE
hpI2RZSIN/4Bsxe9y2KKaGLRFTdhBLKIt1kwZoPGPD9eEkgx7c0DmPMkwBVRHr0NESFfkmacFp9h
f4KGLFtavG3TtR7HegpEMH20Ir7abvI/VMDdF+y5xEPReTvp4jT1EzgO7G6APf83B9VH5UPqKer1
M0s/dvW8a4aqqHdd0we7gmVKBHtYJ/6Epji8dsCFlbXJ/pYHMZ5XxOfIdcqIB8v0f/Ul7kaW/zz2
aW3/VPkVTxewgl/+MzUOZs5745gT+Cax3IlzE16hOZkRvVO3IevBBzBDrWxD7/eMWXGAeasUYvgL
nM5HDMHI87lh6MeB0RB1dWrXzSfCcqJ/9yPBVoYCd0OLwA+5PNvkvyl0S/De7UZTRNYegto7xnGe
aIJRok42/KeTxsbMNP5nlmlNTmKpCnp3icFeBDxvO8DXDJ6NZtJC4t3WuN8u1MLyXlGPtq+RPP/B
aPVdjse+y+F7P5sSrrRhdEQ1iBqqgkblTAXBIRQwvAy84DR/TZdmJQ0hsH4gHYB49KbQPrqw8iTi
q6VJcyjPtFFXK+u1B7rUdCnkTthu1r3KxBvG4esq6lKW0CQqKsyP606i2LlyUNMkm6wpzxd3Ecob
AZbSuxjo8rcxbRgk83oOGpXN+Hq40woXxUAMCm5bwTeDHlkGR/fZjDrt0N65y5P+BQXv7kZ1C9id
mX7DIvrfYFazfEqwS1Tjg8nHALkJXBBj+IfcDRtQ3HqyBtP7Y4iP6xp34W276ZJDZBRg4GOxCjKh
bAd+uSHtg19Djyc4ru7JpbO90T3Iu0F/OgagTn1d1D8uPuWmXcKOAHmSBxYCN5c4fj2+XldgdGDV
Hk2anKEXtf0xzoeimqeOF+Di+D+/U0YO6atiGQWq1wnQoDQKebQxCHXrBTPSl7pmJeC10/2BFeR2
YvTUL6Xq+PrL/9WM+2ce3bOUsdGGEuq5BkVujP9lAIJB3Y4ZMPAgGCerajUj3SsB1fufAUO9aXaP
LUqX4ZuzjB4PScp7TQlDG2R3GkvChbW1MGbnotEV99+7Gi5F7tmhkI4jeTJ7BcjMSAmUv4GMj1a2
phhawZXDX/0nlyICkGaZ7F8YUZ4f4SqIEorq941WLnmGAOJikRCdbWpuP+iuSXBuPA+4L5/TjJLd
VhymeOU0UbWvH8k9VBuwxeCO4qJD6yThy2OO7t+If0RbjyWCBpkP/ZxKWyLphQJuMLcGkVdlUt57
oenqcTIWjO8N+nDTwWjpi1Zj9mkyFhS9mFQLZA9hO/0IjhsodOkLLbv1h+sQya8r61KkZ177L38Z
x8SIX2cewRF+anUVSnHKWeMuJbPJaUKC4L/sIuj0ZDNV2SYnLM3EiKDh0NotREn5aGdUtyt1GLQJ
FlJWJRR5EYcARoz0qxHv/9BNighHq+gi2Nhsh1HkwDNOa4w5pmZdKvmS1YWpA9tUkwgbPL2G+BmB
XBeUFGNKdUhewJo4sHcuQA3VHGcZTw7OWK++A70rdC7v4o7Z63WaTRdIwsWhb16NYaF+UoD9YJbN
4c9gdlE3LSN47i7eEc8ednPS8qkeyK528LxXWbSgZVpZnsn7fa8fcr3xUfOwUPiA89tqHB2Yl3kt
k0I1cKi4WAAaqf9CEkoXCCOZ/okNlBL9f34+5cQSLU5GekeUK7xpi7TOpMZxkpgSDEHvJ/3hVztH
YX6LS3lBrOtZYpDmrj9cSCtLs8cL7y34LGiGCOmyi+KYU180ll3In+S6FoYtxq2e4fhJpkD0mHfW
yAIFzlPUZEKmJYlBwsQsmAn66WzNhfJQ6TqxpfbQCr0c299Fsk9HS5zu/lxVGBj0U0K9VdqmEUUs
Q3ceWoq0oKQjzbuwmmCL7+zeCiL3FTAlBM7lijwVKbQuryjeJylLmMVBKLHMCJ/QBQzzR1n5Lxuw
XA76BQnlptfI1cV+mqG0c1WONvMoYDYtXWy/Rk0295g8rBaS4FVNreoooHOLGxHgI8iLJbFpDEjm
1A2CU+PO4OuNrptWS7tNS8qanssJi36lDRciHU6wHIxkKcT72bVP9sTytYvH86jc6TXFmk/ih5EU
BmVJz/NmwY7Cl0qs3+Teh/J36Ld9WY3d2PVrqyrRyf6KqN2wC+7aHDmPL5BeKOhsuD19TQBwCvye
Teo32raXv0u0ChbMIXSVbvC+N2TIzor7PI5BD5g4quzJO3QcKflUww5FTPl83APTWUSSOTnbJfVE
ggIRisMjnLx5apKK1hQI9fsu6i6MRdERiIl1cHhA8qzDYXZoqP2KTuMKcrYrKfXs9G7i0C9rDKzc
OOqFkmcd5N2dj2C5v+rYb1QBsYiW3K2oS6fZeOcsnT6y6TewiAVq0tHa65zjyf47CBDFoTwClZvR
ZdfZ43GhakZ6zGOFB8kEA1lcB+v9OZJJh2+98RjHpC8XKTqz0UvZuvhAV5mfSC6I/w/uU1x9NP+w
/nKSxB9PlfhWcTaRFu004Dr/xVcZqOO8h/XfHa7wzNcU3YjF1HSPHGjXJHErGZVxqLC8B82Vj/pW
yWeyNGZ2o+PxWFJniesulH4xitgewOrHaq6AM+D2FvKhtxvRzsX41x5AJMAnJhe/HBD67EFl2m4R
MuaiVoIJ9sZKemMiBCngQkjuB4Ew1tmAOoVzUYD4ixZqwopgpzXafKMvu6uIknM7KZWfPMcaN29F
0H84xFinOb/r4JFTsj6DfjAU3GewElv+8reR0UbiTPxkQX4ZDQFa0QLKiYZyRvOMnDkmNgcfNOzF
OpQi4CBQWV1Zts2OCmEd91Doi/p8kTQn9xotQcUdt0d16cn0Pn9HXKDd9tYLXrdtITCiRTjzDyFQ
jDkACQ7LXROPcW5eZc9W1wG4Vy5L9DjJSL2kbMRDEjtc/ABNk577s68dBHLNdX1k/2QFeMKnw08O
aSpXTfKshivtJcYgIpPA0jIgbVsfHkTpv+lciUP6DH7xdn53PDVBH9BcF5jEgs61VhrEHiQ6y2X5
AAy9OQNsD/OVYxfEdCcOEFhHMqnxLygCqOCinnEoX1yp30iiulm2RoyFQ10rZxB2W/khK/7OR+Lr
UDYoM1A3vo1mbQO7yJXmdZRh6NHOPtdIA3AwWcjJqScJwQiW7fZSgXUcDUCAxfDqFjPEdetMK/AY
VJzg9IniNQcxBP1ZHkAGAH9W/5gZ92xK3q6JnoRZTnVS3JkNVb/7eQUmf0JDypbYWjwToJj0kxuv
F913r+d3aZ+VmfMgRiMFXX9nKkMVmqYrbMZYPOI7xyRPHCOX1tTUhR1gWMWltDZqUPVIF+2MjezI
kLEtN1yirAb4MZNt8Ul8Rm52fXBHF+Ab5Qz/+RsOu+EEoNCude/8q/gwLFSACJeRFJcYll81AwpQ
KygDA7jSss+bpOUnNSpbaQ/w3MolUFK2fBMd1C+sGGV6h5T3JfngiJLhSUir/apUhpjkWsbyPhf2
Tn/6Jupr/iodc/QvAzAaHGpT3ioOn/d7hCLwkYVs6sM10A3yIAgvWwC60ksJwXNq4iEun1in1i71
ramFhLjfkLBBcWmpMztpHNAo1DCM9YDTM74ZcEwYZ2PFZqQ5+/nr+AAOggyzsTLIxnfAg0Ma6Xx2
/3dsDDnYXxd8MHXlSVPVcnSNEDqDd6WHGOX1tBhJkQmz2Ly+fzfF42S2b0lUnsO+xkWMlLoRlXr6
YEITrz68LwEJebtGLNfCg3MtToCrqUm+ONlyPes2f4gJEfurAYAND+TzY2Y9Emt8Kw5uOaxWSCt7
F5JtctpHPF9nQ8PK8UEhjy8Z0Tur/s7ltflz0rf3NYClfhbyv/Fl6L4rBSjT6LcWEmzTsw1Xi/ud
RFdDSvk24WjM9c1K0ZrJbCSjhWQHnsAdG2xC5kFv/5wY0qTjzMu8mMOaI831tWJ6kEtGsclVGW9K
2nnEbi69lvWjXzo37gvh6OM/Ms3ED5gIFKsHOo+cHRDXzhVsP6lXhhNouSOtygWQbzpsESEH68US
fwg5VXDaof2oBmb78Pdse9E9rAnOTf9svZLwi/2TBhK6zFE/pAVWIiAujZ2TKIgrbGGzq4ERtI75
SvlAfRe4QVzLhjVRkchsYHeyiMgORXOBn4owdGXEbZsDv5VpXD2akAJQEb81/zi32dIzvmwf+XqZ
Z29vxHrblQwaPk5EujYNjq9jx7UalIdZyZVLb+dHBpIZG3uvQpGS+ZqlX1B9HRVK1cDOlIxWDvze
l+T4f6OPKaYuEEUeeSpngjfrFfWJzYWi9R++nMBOFKFAA+8N7vnvHDOap193/IX763GY1FfW2F6e
rZ53romn+XhMKdHKOSUjudqEWC0io1KtCIRTqMlEip5D7sz4cnBnujD2W2+DsgUtgJKWmqnu/wm3
N3AZWTJ00LsMIpWIlFS4hkLQcnuuJRLja44bIwBqcCt2dmrY7QiY8fEaVI41s8oekwBM0Y90bYRq
KCSRzc4DBeHjWG+6uHiP7h+jLAj4o+hvxPGqR7a3tB/NHdzIFIYHWRbkuZS8NGN5Dm6wcbUaais4
WzADparzS3r2dnMdD376CtKZpBlQoIIEz3l7z++dkdKLT5lgbWDIhQUypTRrZewR99It/8H0OCiI
qF30egYcRidoqk12x2fMBO7sYZPuPIoO5P9YOevay9PpucTe1fYR0XHMfWcWV0vE1Lfx2sptEMWv
C2q/PrnKpPN6CziS42q8LocSxwuASe6k7EU05DTpyZM/HmV3djQ9tDFnVSGEUjtPDkl92ws9dRoE
Lr9BeIU11K8FZ/p78OFD13SbxROMGk7BjRNXdWHL8wYrkkpgAaSsE6khtSQDcjL0kJfnMokv9NMu
TDJxWmyXnK8eX254ec0eGEwX1L37rGFXKNI6HhOgEslsgQsCpW0CNkyNpCxPaLjovcY1Ij/44zV2
mVvQ/xejy03eM95Ro/o0YgRVMg+iUtiujOTxnHqLoe+bujrRBp57rWNm/IgVtfcpyoPuswP2jdK/
UtDLenPaONGjzE6RzqoReEFKYfYLUudWpBDdsH0J0g7os9foERPVx1QUb3sAnwERqk/T3DOIh0Ri
1HtWLQ8nioIjO4efBjwTKXgvPGqMUneQEQ7UE6ShJuNuLDhxw2JigosjQiJ/cDBlONCZhmBuE41G
PyrLNnFT6h3mWUgzteUcN4NiVgQSQVr0rcqsKZESkCWV0m/qIznx5c/Kha4eYduMBaYAPlQ6N5wT
Jht9XndFVCuDo3t7R+wbg9flLQnPcrTCB9qggDiXI4cAQD+51ROMEKcPa/e3jmDqZbm5OKzM/cvV
dkjznidCWRoA6/ZjDN6MOj70i0Wo85HWA19iWgpU5bmF4PN03ePcfbyZsZS0Vlz9dde6rk6DE2ri
8g3Ld+2ldElTD68wosKTBnWWAn2YGdV2VYROQpUrgMguKXhvtNKnq1QPPwAmigfFchN0g2P7gief
GxjGkIX10juttGhnMPP9vZ6VUdcTWEO06RO2xH52w1eL66bjy2cLWI41FnvYcdkmabtn6oJeFAIG
pT5DKq13qjvBMFv9u8mpI9HcO0uzccDtuxd52eAq7rnnPx88DaIq+ftJw3NJo4LNnlD5ajvEw4sV
argqsvmWy+C08Vbzg357SZF24KcnwuHJ+eLp5TSYpg92+zuNB6Pzl09SAIjA3XfbY9CCVUZnWwTP
aGaZxodXhGyGkLkGHhc71cGhTCY+Q2zs/MiL3Lrnpd/wBMW77DB21aTOGW9Mm/ZBI+q9GBbHpKW4
s/0uU0VjraEeo+gA3MzjndPz8cl9jAqnGQhthY2ozaYo68o45ekTyHs51mzDJUOf3RjAXCPN9EBI
FW9+ickWAnl3DukUvy0ChP852l0awufAa6Uwr8gOdt2xSiZ/3CrmNOZa7asrw64AbIYsoVtg6Waa
d4mylnAq3xwHUhFHxHGtuT7kyfUOi3/vBXGNsISMsjkW4r8dBQltTeUV0ruIapGTmX3fUrkOe+h6
YHEu6gFxC8cS6JBxfPbdNv9jpF98xQAi/S00AVMQ3uH0ahvyjhr14xDQE/R72cnWJNSFYtISMrqZ
bs6lcvR6eRO9T4H2W5TOpHudfGoopfj2RprUqCbwmmNy+YztV1nXVvZgrRYmWZ/kN/muN0L2KjPV
StrbRnBK6q7Vc3TQO4kvmQjU3uQHjO5cYtUEaPWd3Rr4vwoEDcAiIMzKj7voX0ECxbYS61cQC3FB
FVYk2f73ZU4LLJ8cZN6KlJuMO+3db5UDiFEyLUvMVGOFe5hDTnj+lrqv0aV8OHz7J7VZgp5AzN3W
GgE0ZCtOGEkPl4IkYUBJ0ShXYSYVmgL+P6rpOMEye0IExaz9oZkme1vHPOcD2SQxi3/UFpnVIB1c
YVG+g5PHvvSo6nJtnQiRiXj96FTOM4DU7/wyrRnf8gUSEiKvip6/32AStMXkDZaKWiDdCilkUNuP
EdPJ7QK2E9G8QyMGk2GH4mwBXipVpVT2bTd7mG8lwnSTdYvVVYv97FdsCWjGoZVGbjMEvWMwG+P3
yYsF3Dds/FE1Ln5jXlbhd8PCTTsYmW7mU8PzvuUjaDJjpoNdlzrfKJ7zjbNb0bKkMSZ9BhNfYxeI
VuIHB9cOXSAfixNX3yw0WwuxdETe3Crjx1YHq/f458ScxNWj01RvsTO9OLvKazBXw4/5Pjl0oK1B
pk23OdtvPOhUf495GbsdMOTSBda24OddVCDBO1ish3OeEFhh9LkVY8FyM49MNEJL3B3Xmtw+kX1d
twQFjSNApzUs32P6VnOCF8py91R9qNqKfAX4g6O5TxRqwXH0FdGo9ks5gr5ydoEsOeBWcGm7Shp2
Msit+m3lK17lb6VPamc8LXIwvP5XIxaL0Go2ERrhBsDVW/HtdVGsU/FRC2OdRxDxB2VcSBP3M52t
d6iYdpuXYOCSFcLmh2MwqlbVj3NToeOr/NFg6xLtvA1umdgn/lCUMZZgDK4EHTtLfMuE6z7lwm7j
wQOWgLFsv+Ttr1rwS40blhzHJKk6L6ZO2ueOeQ8zZ8uA6pvw9wcPX7m/9bfn3h+LbbkXL5kTovNT
MKaTZ7F2VKyhitD7YHcc204nX1amyP+FnmbQ9f8FN5CP4YsmXnIBrafc/kheyHXEb8vvDcuJ/FE9
mjk29u9B0T9JeFBEGh6ZPjYSsxNnlsXy7ltQ9bssqHzLTVIPQCyPZWprTbUjESq8g1Hzxy6GF7Ja
K13ogRnqu/83TDNMiYiHzKpPYJXErs1CzFJWH9L2e70+OjppVrX9ynbbn5VjDXLIUys5cAanKgH0
qN3sobRnjtNcVzNLOaMvfduVzdLNNIxUOUk0qWHa7WtqTeqKgAq7YIQueulFewUG5ftEpeD+lS5g
SVpdkVXWbc1kwLDggDeeahVFX/F2IjpyhjolhzRLMKzd4uJyMPFu+AdGwgti/tnRfenEfPwPQzNR
lV3ogIAXgqbKNyckNNSYvyWq6gr7Gm9hsLv1eU8mlfcYH3a8x2+ykBkTOrCRLTCCiFwgj7bpctdT
YqZpNEQP/PVjbFKuQq+MNVlf9K5DPt8YHYAsIIVly3NZCiX8OC1dLjp7CcKxwJ+2rCQ5obVAqa6+
FUH/XXZnvod3gZlE0EtdIJpltIAIHGNQPgZGcCYUVk2UVKDX1RDjrUeWAzhIxREf1RLUEy2047Pz
ITl+D08ghLqFP5EUJrTzTdHy47INt4J+CK2vpXBQ5PcBENJ4RdCO4HSXsi90LEk7jeVhE/tKg35B
peSiAU2QIivkGUqUbvuYqJepN9RFKEpBrFcaKHafE5Zfr84imgw+XpHgZdC0IACsVhSRxAZWrNoa
lpgOhBo1KFJOpRRRDP95D0hIgFDanSqoRya7FyVJkWf48iJG1l2aOjyX7VCV7PVq+q02KpSlAAA+
ed2Ci1RsihfxLDdTP/cAaRwyQ9J0gnIm4vd+PuY7dYr9fHldoRHrYRfjpxWYzbBwwX0C0HPnG0Jy
kuEovHUPfBiFG7q/QSvcT9Hd55HOAa01N7WD66l5s8Ei9CEfkfKmRH72UND2aDcUNqdIgZaw5BuB
TjKRe0cuSkyjRgSeMCAw9nhnB9I5HnHULlde6N8R215g0KHI1T96N0Sq5bGs8BoYodovyADZWAkG
Hb87EnbDTZnkM75uVgTva79xWOCoknonuQWNd4A6Jq5Th1xsyEuM3OjxeTrNjTa1hgPurvFmd4qI
zR2+V7+/w/3pzJ4AXN81XWgPuSrx6N4g3UlDPFnf+uSxCAWic4AxH5eDosUHK6Mv/z+JUAYCR5vb
dorRlGztZoDlaJGkrHr3PCjoXV+mDAQ0x6JjM0COVCQ3jHy6K2+gGwu3pc+y6lpi3zw1W3JJTX6M
qK6Mh4QGd9j6o2Bd3xZGGWe30e9+zyHn9eoL3o1rQJ8ICXHL3KqqFmc9qaciL8ODGHKmxD9bkpsA
D4FzThVAx1DsDfa/l2vHDoo1xM9nuKx+Dnm/48k+m1DhRQ4TAYrOEwcnvWovQC2eHTTds4n0v8pS
87sE4dFDmgIP7SbEDVCEZY77zMORf1u0To5iN2hMsESyp8Y7k5zpqyllc7fGByE1VwtrZiCTfLqB
cpvzdLp5fKH2p2Xt4q//lSPrt3eYWdsylynqTnhzKFW/YVOGpxmwADm7Ffiu3i1jnTz3h74zIwJG
6LkE0n/0URKMzIfkloATNIjjU4oc0OiWDnLm9tkQJGuwJ6BlSGGvX8yx3fjKEz8+ogn+UpSljwaj
iwoZSU986rKnVnwT9AUih3y27PjdA0546aqf6kcIwFmxhN3tIwPL7Wp9Md78ZNJZ2tN5VvoxZEwk
IBaNRyo8pq3KaW650WRV7imIuSGt+yto/wpxCFScEJJzCW2Br+QNVBrnYefaXVmThcwIih6O1XtA
O98VM8PnK4DlHyD7AIXqz7crFCtUGfbJhDjuW3B3smE8kZyxKc7FKFnwXCqhyikoWR6JL9KZyGHS
argnX4WxKk30TJCc7pW7Gg8Pb8v7MTtbx5ehTzKCPENzrZUF1x10TICpPpf4wWWKhscUaQaSG3h6
UbQ9chSImOUmv7Vc2MbxmzWS++ByGGIkVL6IDI+Sm8K2+ENCmgQbc4v9k6vpfGF2Yh5qce+1jv8l
yPHmwmwRmRE3dlRwFLZdMutLzYsM86urQGo3uVYKYvre4PLhFmZhU9jtpv5XZ5to8cbN/hBqDdDW
v9i+wzGITAwvu6bhA/2hCHkSMoEwMj+FcgrtutJd0AdsOAKY54J2o1JmhdZlA6r1CsiMIstFTHjZ
5Aq1w/Tc2NJ11IRnteyLx+B0iElCYR5uqVLy7gWytU3P70sHO/E5LFdnxVFVfVhjiMzhtOlbfceK
3z8/iFmZbn8pAuLwQ7YNhY3vbSOMhcbPl+oBQUnammynVhoA+dcgyy9llTSyi9xZEhzc9NfWjnpN
FZpWM+AOd5HGF3cTMNS5UyA7xpnkzF+narHqfb6sd8x1g9J30+XfKxtZBJoPLNNwX86/y54gKeY8
9kdD4lS/CYT+L0It4PQtTS+yGjSi4KcKvPG9iyrnMrl/s19ODk2dCg350dKHTxE+Ga1gqQqm589r
pkwyp034cxhSl9i1tRUh4uzKv9XKrg8TVcJfINtf6Key6L8PNQo58sk1bpl+Th/77TtWbwLz2rbI
QiDTVvHPnQoOWttYzVq25SrfPVgDG5tAdO8BwtH230585SiQaoJmo/mm9aNh+msx8l37ljRzZ4Ut
93CHGvxqf9i0+U2txjo+bzElPmAKeehhj0lg0H7w9xfy2DV0FjSxafsewPr+QTifMG1tet7637d0
VLUs2Sbc1LfqoCfnQP7G1lI07DpcNQ+mBhuEL27aPIai4EElg8HjvHksI/uomsd4JSU7uQjIiPy+
iJG09fgXjmEVo/NhPsB3AutX025PmgVHyA6D1u7ozUtUHAlcxMRl/Qhuwe+OBV6RLysWX7/flwhu
PAAGZ80V5+2RieVz6w0JpWU51knejrVyuNVtJATkNH+tGTXw0aHiRZbk9B1IkYzABiOalwPWhbcr
mXDIbuXvpZFW2HWurCecNs1sRBTkNPHhP7mOCk8fzxJ9pzE+2MJpUgPROhYA2xRL8xJEzLJlbl/d
aFuNFo2T3dBjx1K7DzudFo+UUsCguwX0JhrER3HNbETM+JAug88MXlhJGrRpt1Bkzo0Pke03x4/V
asZxdtDpE0yvyi+DSU2fO0HgH+asy7yubxAPAI0szrY77ueNu7E9EONjmwqgibK1iwB7/ccbsCvw
+PNyxL0wCMVVlOP8mYUsbWfz2DJ6OeRlibwMg2XWPCsjzMCbxdsO6MJc0JtKxitYww/2mT73K1Dj
MvaMMMA4STeOnDsTe4mFjazG6ZdKq+5hcf8crsiqgt16fSg0vg/pWimb6RfSukrcY6P1XSDA6vSy
eOS1/ybHejE+xOOifHtLVe3Ko4F9wQqW4TezmdK7J1B9C9RQQ/xRSCWIc7+Po2Y0wp/ln69I1WrD
wcOksEcw14jUt1LiXiEiB8oHvioCqLaZXLbctF/LeRqul3C5cNDVLzMNd9Ymvn/Tqe+2e2EG1wEF
vf/CatP2iAf3ivzSxil4o3KR30zxMbKbgwYUD14D7ByG68gCtyhqlSEm5x70aO5SUM9S1N5jJiMG
b+49YHqD+u7KjoiJeoFd539GqHF4Dzzw6F4yia15pQKNQlfXVh7MDWZCJ1TZaRSVoIZzdakLGOXm
QFfkdfHn8MvJ6xafimMKOeUG0Rm+C3YNBW1M8Og5jJ05fQi7ECzpskQkM5m2eW4UNwE3tBjVKKBp
qnL9ckz60iN70hYyG0vfeMxH/IaQCNrmm3NFxSEPAV47lRloSgiFrhrhY1RPZRYPqvTyPnzBLXLy
VeDy1Q2TP7xPt1KDZ8Al70RWEske8bTm4t2gVlBaSUqEC1EDe0xZkaD0+4Khgf33YBgfNebhdndp
rxuxxZqBDnW3c1i1quRkeyR+pIru6WZhIWzoktvJKKhTSWUA0W/kxxcLQJGn5LfsmJ6CrLNdIXTP
Q3DQ2Gm+pe6GIR0i6z4i34COS/pvkAWc0eIgBuc1WqWKKiwlllbX4Wa9YM1QfTNVUuzxxEEEjOSm
Wn/A0onDT5YLwmcFRGQiIg0TN2RbNWJ7EbOJ15r/cKRAAmFAoMjhg6qpVPJedDeIIC3NAW5B3nl+
Rb2Z0T30KQRfGVV4d+hTVwlk/TEi2W7TRDFROXjlJQljUhUt3iDwg4vgpp+QA8MLzHU2Bu2EKQ3x
kf1knaJZ81vKcPum6E/miyESP4ub84YySXOqisVgBGt22qcYiEmKqMA77dAypSetZTrLRJIsWvDM
TAGEqpEkJqVKBnpDJT/OjNngfWlEUy8+4WIPlc4YB9O/FJbbIQnjXPL/G8lgfUhpqE28dbECFtSK
U4ckIEdSK0i2C7CNBx5WFwjJ3vNFLrTF1onLHQH3y7tvFEWpGZK/7Omlv8Z0ufl5mxUtQ7c3CHDo
peu+9jqafcplIPNzUaRZ0vF3dXcBeAhwkQ7vZApzY/1mxXaq2ur57RftYZeOoZrfR2qCWkGElSlv
ckWxxRV0riq53aInab0MwkmqyTpXHh+C4dXdpkqmOsozCGPeqIGPWovw7zKU7D69KQ56Nl/U8lod
Nndz11srxNe4prCqO7327ehtTvHaSrdsQoUkOyl+UsEVI0LMQ2sHmwG81xFJ3Kp7dPIQYfSAOpmO
IHxk7YJM18WDjLciGYhE7uwgtS/6uDgr1o9LF/wB3J+XXCA1s1AkBtZlCYZJHu3oABjPXmYkxGtk
C182RfbCnltulK2aF3LUrPPqYktQhFUmjI+0znAcNCIjkjxxJs/XfEBGV8v78evugkMHzTPbNeUQ
XqfmTSc0cfyYsleh0CnhqAjz8YX1qFTk5xw4kL8E4NwLWp2HtcyC+pwL6VZcn9i6sMrL09SJapyh
pJE2dka2WxTtJ8Un+4rV4yF4m5+l1MnuK8YHKQkgnnIM3udHsZFfk+//IFr2XJDnjOsExj/0S2dr
5imrT2k8xW5BQ5ForQcKTsIzxq4KMnczRzdaE/8xVKiN8raOIaCCIRC8XcU9/m5JqortHMZhiN90
IsNirkEwmYqnJVtUmEAhUNUkWK6UjfOXXDbmurluKS9tTGmSx0dlxitvG//Zab1ZrpZhLC03cxtQ
KuqTrv+xREtPhpg+GFVws0YQsZOq1b5xZYZUkCe9oEq3+MHwaXqUiO2QnxftD1uvbODNmNZSuEb6
bUoMG6Jg80lgtgRVoMBTzGrcHjSCPrGSJDa2ty0QNsQspL56jm/g14zu79yTT2u+XUhCMg00t0r6
hV/ywyxhV9gF6ccxH1tKM5lNASTH2Ni0nc9K+1QIovBoC8PojZrSGR/SbanaJlYLZV++yEygcPvk
9EkYvKqJ9Eyngj9L9UctyMsxvamvok/Syhd9uXYQ33R38mWHiA5ZHbDqQ3pMFk4LNkzrj+50nnvg
97LGpyz9yYqQNi9qB+2628Dvh0/D1XZgdRfdIVclI6/bEdvQofQl/y9wxjTQqPAEzEpbH8YKwo7/
nMBKjbBSD2JAoNa6ZdORTneMHgVIMsjgg4nPkSp+e/4KLD2tWwDoWLR9jhar3dhl8cX4tQW/e9Ou
7+WZqVlao6z2YhVXVCcIua71LmL9603ozdNFz/JEI9bWeLNJUL5WTo3mRGqAlQPBXzuzTe37zrpA
HPbSHWIy0WP9lHGDsevLsBMwEXboSAsNH/KUB5b25L34xVFrmD+Nga3gODCBkc4hmG/ceX0nm7WG
zhQuX4AT3KULSGGUmNnh4O1+4iJsVXXhbVfQwbjpJPSiwYOTMyX59/wkD15JtIX3g5bE4oTEyC5Y
OX0HSO0wGc7ShG3MOD5ZuAy5X+6y73O1bzgYK5iMS9M1Wunipp21tQeyTOUJD3vZ5fbINBzhlwKW
N2bACi8dzCpNuSRD9Lz9eSQIDmB+DdSkPZhuyCnmOmoOD55PJZlfOG+H4j3QHCy/0m9kotADrkk9
ThPsCPqTLKxrYcaZcsoE/EEzSVjCGryTbArLhTqLdGenZnltl5X0tv/f/W5FLsg6JGoHx5ftahSP
nbK8picSS3zQMZEaEEyeUYuTxAhtaTa0P685423XcGDWRyq86/S7K6pn01eDEWVDSWuI1s2fIEoJ
H82Ej/t5jNGe0wCrK/XwgBkQ+Lgvt9iuXzwPrWoAkp08cOVR38l8tTaSSbX2SYRAKIvw+KTxJ9vF
RNrBX+KQ+SZqmFPseEGXTbjxqu+UeE/YGr5xjv922CAbB6vaBg3NDNU/DIO8pcfLcAwiC07WcdUz
dQPLttTjmKbMsTwVD2/wY5c7xalnfT9DhP1LPMrppU58T6rNgmGJjw+YGKPO6oifKHP8urW444HY
3rjzfWS4c4ffdwNZSmkYwOXrnSyYpJOJ09+TGr/bY1+1allFzdyqMalALJZfp72eSjJdr2sQWPSw
kuX+11iMhhWHoAr9tJunUDBU6Qp12Zo5UfmiDtyLr6tW10dAGCtvum1cxjj7gS+JSSaiB9LltDyC
Dtkn7hNApsBf5Z8omeDn0Fezwnj+PqOqPatrecQkNNM5l/ZjtuqwpZd2ohm0xKOSf9T4RxN3wSLU
eYzWOmdzbbYALiZuDRCsOgJuWLOZts42AbSwJrjoFOd7YDu6epi6VgsEM5xRAcKtJFlXIQNfhnYV
t3s78GO36EBGe4UFeWy5qtIO6DDr5LGLHQG21PD6YG75kFhNXWSH8F46uQ/nEOdW0ayQK1/IwRG3
YIEE0SvDG72Z3T+9e82XStbaTDGJlgg13KLTongl6bXrUFyN6lZNiqmmJcipZ30nw/YWWA76ZRtN
UEFf1yAHWFnY5SQasqpyIjbCY3U2VBbnfqHiSP0r1n7mzSxG1WsaF30KE8Mgow08M0bAubbZfcgW
cBMhJQDh3c1oDpgP+gHABlpo6tX1CZDsj3om8m0lubRWdB5DxUHlmEQ8u3wCy9+QQFGR9zh5JSFJ
gdy0Bg1nnp4YOWShyNLvV/v0PCLgLOO2+uUW9evX0wIvuDbU+WCzWUUU1IiJ+9mMPcyoPbBQBhgX
vi5yE9PLSsCU2GQwcUcfw6jFIWnDHrePQSR9qQFzBEEO3r8Q4BSf9Z2S2QRf/aI8N9krBrOWm5aZ
o8Ox2naUGMiIgdHHbOxpCFk0KUHlcD2ehAWEFLDQp0dCuuDVzqkPSYS+2gJiBJGb8T6SZIhZ36zK
z6J6G8mBGMkgoCHokHYTTwlJLtYCBtCgyAFd6ccYyAmGq/+5HX6A1hfiDd9q+5ZGNatiEt71ZGRT
z3e3CFLVfz4S0pgOQEXaCUKOj877NA0g3zhjsG2ibY9HgG5H/pNfn1m8cbnSace6DiQE+DNpca/c
Xjg4vSUIi09Ks5LU+pR9flGzlRQD2+HjVduEYvNxZwzW5qAK9Z4DvPNHFmrDSykBCJPlc+7aADA1
2lPa+VKtPID40dWyW/noJ38LUD9M+d7S6F41eoFS2h7tPofbiPl9jUfr48lmFxoviCtwp6vGAfRY
iIBnqNuPcpdCk/V8cyAgH/tEROT/ppRkgarMDR+rim47wH3uiQR31q8lHuHimhyGCWGoFWIYSGKy
u/WuD6moq6kRREUt35iwUHVHCoF+TffbCL3FiRKbj+kvH/gT1CvSMgp0jcoG1xALo+i0jaALVsEp
Z3AL5LjkWZtAIZuat5u0zqMcn1iTcBPE9SUMYu5NOu0GbVV4MuSe28qvfdoTUFqOny9ziqhtP9s1
jAKKik8gOTd4APhA+jPjLFzfC1cCBtph3i3wLpu1SgP6PMnb0aKeIXK41coTi6Sfw0UysHtm+hAq
VKROuhOmkpgW71tk6ldML+k9F1FpeXGdlcBl1cLbally7dGTslPdMqj0b181hZw2UqcLGrOpxMPm
H9/DT62nCwKL/tVeuCZ0rN3GWt+25zlCYq1Na808fdbSj2y/54cF6rV/G1zD3qHoJe5lBG5b3K1s
kwU6e9JrePspWgjDdROO9TgpDK+DaaIQC3pBgS6E+7XvKfgeAxrbQoUFkgyTAksCMR3xxj0+N0yk
cjVtfewDw7gMeaK5jEZFR/vGlMKGa4GdKgiCsxrD1t85pmoYFVKZ9tny1LuarZslPIluU1dRBzdL
TsApIvcoZBZxco7tLxgc1N1m6YoSPiKthk0DSakWZN02ZhjHUwyswFnGodMZ29on+I9r459bWXly
UyFUMrN02EomK+HwYt9kmc0MTSyTD2qYJSMXh50xoo8xw51Ym0WdVOrT7TKcJpoydvZgq9iO118K
oS3OEg+/y+A35O3Rt5vwFX2JPWIWCIbEbKSS4nbz99CYf6Z8GRv8ROnZ4KRIvDar4ml8q9LVDJAK
3z1QOfKPZomqNF5J0cRCQsJjKLqmdvnGL2cyqR2PP4JJqdFuLBipKBAui4MIdm1LzAfWU8KsY1y3
ImBPKKwEE8eh+o0F46GQtMN8GbtztjhSd1zlH9+/0a4q5bFPLJvMJT/EAgEO2Bfz5hcDcOFVO1FB
mvpBQiSl30Am+bQi2DeiavsnrCTi66Opdy5jOmpKN6zLiPziNITWTqHZBUNPHBb7atnNAA09x4nx
KmajlUDT47UDNg1KFe6i2tyaiBju3gj5TwpEFP3B9tfw4aibyY5C7apJCzmkLBTmcKyMqpQoAQAQ
GEpJGQeF8mGM+lQI74ChD+6jfcdJsSQKnIvQg/XQiWOdyp65pNEZwblYyP5rL2Y+1FOAXmfh5dqH
wygHQMgOsBaYTIInZ1wAn39fWVFd1W/urwjAK9qTyz81eaHZmoeg32eVFuoQz9JZuaFVjs7kXGLQ
TxekhLfIePZSxADn5UamxUXG+jux+DtjXl1HhOYRR7bIt+YUBwJoR8GyajkHEkJPIQc9Y8PRUcmP
jnQpCIA+iHgpvryh0behOZ3FftZHvrjl+Oaf65WbgJXXFxZNUBk5vCILA5I+aVaMruEvpyLcfcGL
J2Ha87iIIaOr5ZmK3H6Fl/NxjttdoVq1kS2XILkBHkRr9+xYkS5yPx3U4zXrLhslwCk71MMBrZFv
fJ+vQnnn3zY/wlNKicDc5Zwqu2W71shQQ68qRfZu6bGaTr5RdUGW6ig9PmLThO/8SUj0SmPWlapg
8/3Je8W5PKELHVBDwscaGMfg++FkHIJBi+C99k+Ua/xCUBInkbsCHiW+gfK+1lsVtBd/uIhgFzw4
cJZHDdwlhA0o1xtFAySOuVchJZDL5NdH/hb5599YfBd9D8QRAqLoFriipCnjgDhWZDrJ2TTvMsnT
1JbZQZ+OjqdiP2gq9RI/mvGXnPm6R/MN/HtDRZQBJqc+YR3NOrpr4krWEHMwDKH+tmNaXJYX/xvL
beyx+Vjjb8/CLkNDDM9kblY+mp45vHxtVJ0HzcNJZc9MVnoufhtHl9yt99/2foE7Ee/hoFBEXXkC
w7rXJEJh6TSZpzAboOAGlDS0g7QxZWqed3kNEFirtwb6NaVVRCKv0moAhtGu/PBLkO2qGSIk+QKV
mO6Lt2UlUcvXqtHonzvkFGtkq+SLH6bbjKZrPyUG/rSBAmH9Dt3XiAujLtQ5SDRYukE7YMRLOoE8
gLL1/wvort/4UoYMfyuELWUS6IyqpNPM3wV36xO6uzL0wLStx4g3x9wmYUDtuPn3Cbp3zHgSxpuA
THWvXEMOS5IVk5jV8TbvINsoyuAjGmypIb/l0N6kgP1zgCbq70CFbG/oRWDuc71WGaxtjyvhMelO
FRFm4iiQtLn2gkqmMLMotl5vE3xrM42uasEa/ds/dA4cWdD8wkqyYsgrs7BUPAxKcXJa5DCO20XU
x4iu9EKzgDI2WqWLv018uAHjHeew7LzT/CbnPr2G4Dov98ZoAo12/1TpoKMcyqGMo9zu65QN8UkP
VILG0BHLqvxudUOBYP813D8fym8mbMnQe9Mwp9RbMzwnnYhFoAyHuj2h7y3VuKkmh+rK6xfSVdDz
GKjKT/7kMi9nX32I+K90PbkFiVzk7LI3EII637ip7rvKPcXxp8PbBWkcpStgpKeuRSy9ILlwShO/
1WdLKuytF5nTc8bNAbQNaUrvXN35eajWkBAe0ZWzV2Fx1gRa0OBo3GGtfAefkgYoD6LSZsf4kzqN
P0UIsaa/7Q4oe/tm1H9eAvca6myUzX8+ugMnGhCqSvU4FfaYUkuhx0W+JRuoqYiv9OFny+8RMwv6
myA2PhgODPc+HbGjLrA1MsxxhGQLmIeVVYZUwYc20J4FvzNpK0+xeGXJiWjh1oSRf84yyhJhOULG
KCMwiTtZQNk/3CHUgFt1yU7xf+jvQ54NlQNoNI3OVHrL7AlJhIn97kMIyuIGxr6BiO03Jv7shHjU
rUfSeiBhnCnw8zgXnEd5Zx3JGBVpLbd7ifTR0Z9bdXuXviCYoSawHqfsdA/WiTH2hjoLUsRMau7r
diR0ZaU2PAzogzaGnwibUZdW/Xm+i0lxW8gLmcOyQ5S2VAXxaHuDsTFhZYPvwNVFcoHpys44vMcd
gi5lZYlAEoSPpmiywDjivmhF9elxMbn9zj1ZTmQ3GVRnz3Bb155iedCUNAfXB+HXgT+Zw7TqNwQJ
qZiQyYVBMJC8vYBeUEOGWndG1uS0IIbj6+omKtRielZ0Yhoy6yhwsndOiK6wbCxaolk9MbUrn8u+
3YDIuzEnSmZM7cNEbiNTR1bofhavuR8TfksVoquZBUHUdDaRGnsuojhM+4vTCmhFqbFxBIeG0fw9
SanNiPVNVOlCDeCIp98IW4JJVPeyI48mcYq2o5aFoDS3N2rgmSOWzS+mS878lUONdxmwqRh52CWV
gc50CCD2TkAsC0nlNwWL6j+m11wwSXV8IL2lMEcCjTlSVIXvvER5LYHp/FEjD3l9YSr1dtgE5hj6
181nhHTBJXXawHoGXucJDhXM59KgF3wCjzyZp8dLtqFFmgfXLhIyShnGUt4q4XMDdTxP9Li67KZg
cwk58ixClCAIaBnMm6UDADb8+ibFwRm33pNGOqUnR+egwETUQIkOLnSFhml+f8NcjG5wDYV8+T/+
YvOpqNbAly7t+7eIpcEDYGSftzSDZytf9pXF/JbXeuLjc4q7bOVoEoIR4fQn8UKt3bP8xWMMn8jd
uNWvYZvKlRhzAc1Gza1sHhKnnoBwoaZRSBI1yRL/5oLYPSM6gxXe/Ibr6iWx67TNlz4qJ7ATI5cA
QNrBro3wSMUNKYNoDs93n9+uyfjHBnQJnK2cDLINHBfG8hl5hYGB0XmynM987msif7qksgIoC5sz
nn3fw50gVDBkTK+6lcMR4v5u3LAdT044GvFNPzQfwREjyOpsiol0Ric3VaXqULvHKNFKCoUCaa3B
uH1G0T3wWABVWxIu2nMQsgO23fyx9FaYgNsdAESDpKHT5FkeTggppsskh8oIvNAELKO3a4L4Yw2p
HPr0YL+j9rlXLw/RkCd2dD5YPkgsaY5h0LbZfQRHwIOCPwM1nll+VWaCYtsfrFuJ5pq61ZVcvIwb
OaagvwhKJwfz9AORDTuI6G19seFYVeBbprSd+HIW9QzDVsxTCp7FpwyKPxMUIwWuckcWMlVxmB3n
zQFhz10JVPUhPn1KVE1NP71V+y7/HHc8wW4pBJwn7oYHcj+UVsJESix6NFPfez6l5b7SVZGStdau
w43CobfV3U07dFwbd1qmz4aeXEPlg9gUmc0eScHc5WjwooT2uogrBIrxttJbEPZ596g2dmTVuRG1
Qft7J3gNYbMQFWp7WeCC3uaKALLac7ZLPi3mDZE5HmK64Ops04pCNmJTTU4gMmK1Bh2kXfzQzdIe
2miB9L7MtX+t63vQ3+iMZ2w0xWcqVfU7qxrXJiSuIw1dqV7uphZP5XFgiUDFqOwx20UXNdTGeqJ3
TTcBNhkBDEQVVYwzZASPFgkoJRNzcpO4lUWKEFl5vkTkssL8k5w2OTKfQREu9hP3+Qbh17jJgKDN
jtXAL6tGIRMQcEJnEBSfOagBlFQIVzpF3wrNW0mZe8DVoGCe/f75sJmzYsdDLbaiXUUzYtR5kCHn
/NgMS16LjCpPWwsFEAPsc1aBx15QiGWCu0J187csH5n46avmySQflL3vFlQXLUfUx2UGzg82+AnP
iU6AqAmC92j0PqnP75IzmtfAngU6wyDmW/k3y/SBrsX0twsF+LXMe8OXwPQCF66wkAKvw28Ubbe8
ImNbFkyXLIiCp026RwHgxTMwM/0zpJIiv2h8DMzbQQT4skzlWAGXEudWfw9wZJpWyNLGfUc/NIvy
q8D3Pmdge3hG0vOwWyyZ1Slk8xJjo36JvbkYuYyVWn2K3W50yjpnCdoac0UWdZjPstMTrJxfsdKr
CYPXyRiTIW21j1V/OyVgYPpqynbZfBhT/mioUxQBdp2ponlwDNfIbrKZ3gAM5k0Aljh3tWI+H0lq
Jq2LWbm48MiUAUhNvF0zF6AdltkRMvKLOJXxaOxyqEzaMXK/7rFB2cH088Hispia+Q8GGff5SEMI
WcDfZUImLalVfDoaghiDEYNDIJ4DIDyNEPhJZipboLRyw7vn/+Bh9IEjeQk1tFKF2ytfwGBHr2f7
2eDMWcPEpQs2wICPbXy6tpYCvQj7z+rClyHTKgXG3CqkOINnsmDdJ0iLeBhrn/RHRpO8iKnAjla4
uRXGOsIvQno7C0oStiLYsdqBYKCSeFA8Wx3FKYybsuc0jfiwhF2W8mBrA9W34tIyKuceFLpOLieu
HuL7Epdywx5oEY88ILytWU2BAdvK2Vu69c7dy3YloqOh7cxHhcXi9RDeRGqK/Sg0yqxcI3cP2dlM
PDB+vAQJbBOjIc5jS0kZDj3yYKlSG+uj8DqEqQWkPZDIIJaM229J6+TLr/qefQppf69ib0bCT46p
++2D+hbCY25jUsIgwABU6KJ74kq6QVcjWvklMnFQqKufovAKc14qeVTOdJJN67PHJ21xB/k9qtVJ
eXS24zIpRC/nIJG5Mcg8/WZwjzvRMC5vy+reJMSrokvVdG08pkhgokcsu1uN3paf6JcM2Rb4mo9f
1QIEKrBX2OUzUM0noH7kLlKxDUE+O3DYpB79vpKqycZ1CTTTQIasD2bIQMcBMlsmePM0/a+wzjC5
x5Ss6dQ60A0OXbBEPPiS53Ywj1LNjz0LArv14eH+3ICFbQJUEEK3YmFlg6bGtPyhOkbCxKjeLejj
KUmvr6unct2solKZQ15esQpcXQ6141qyfM6PGC0Ia+/FVoDuafmYjt7yIGTMAI4GGG1nxExo0tsR
X5+ici98cm2qVq24cGKgE2mdi3jD/nIqW/g7p2nr/IzB3pArRHjY5P1o+I7oOkReOSTvDgI4csve
DX8K5ofwKucp59WQeimVCGXfk25/J9HMs9HD6dFKfO9sZSjB2oV6BxECanJha4M/d/fGf8QhhAAf
aqBRuib2lRp0eqC1Hx+N1Ub54bCJ36t7sE04R+xdqt+rXd0PRJvAhJaq2LSE0i9PmMQ8Oinxl5FB
9xMTB+j2VJFnMVbBR+US9JPr4u1q01LF8mi2uPSEcstkUfN/3LWhwBTGSHgW2Shr00NOc5OkkYgO
fUsWoOqmDwAyqwcEFDLmBsB9FAeudq5WrsvRI9OgoK/MFUkVVmnttOrC8Ykg+3kJM0e6FsTlFd4V
r0NkVx1KDaH19KO5aAbKILU6BKFuyMTIqMwGZnAC3svtqGoIu8UWke5sdn8K9AFXvKaubjKW8y6w
t1GBpy3xBf2TfdSB1QlaMRZjAqOjw+ypN2VZXbq9AYBJm/eckoGmNno9s2olPt57rBTCaM7V4rns
IXq35OKlCNYrCsLJcrZGbxTbDNL+eXYHO4IoHukmqs0xS4O5gW7cw0qhS1pYl8FOhAl/0GEqId/R
wPkhZf3DuHGaDTNS9MVGbCNjK+8Bcgd8W/j4Bi/qyDhsUkGyy9G4fj4IKFkhfIc98+T6IN3fkSOn
LJJIgOgnPa/04+2zOFRsipe55TqXAHh6WiaNmlJoZEhxo8BJQPcm0IVxwrH3xFRznyQpGHRuN8vq
2aEE0XqOEosMMbo4f6wVefsBx+Xpe62Ue1d7GNO0eSIvG/43k+ZIQGsPrnXKvkmUnppfeNz9TCmJ
Fudd7C8dYXzFTe4nxtyirdBmnQhKae8nayikCoMEiixF7nbrOqb2aasF7ZSCU50nNHrHiGGiDwU4
cAXDaJB/vOggOV/t+RAuFSyFXmzdHCbZ4iE+bWZr5BDqbHHrOl4UKzNXq4V1Wbv7Z8vA1hDct0Wo
afGreXdJr84GkNQXOBqOC4mDjSZsw8ZmRb948AgsA9ajYUC2t58t5Yk2cU+NEN+QuMn2CVsCn+zN
N1KvsxqLofLtPgwT0Dzp6xXpFDzq4ZDW8pNPLNABsrZUWo1Qj95m9Z4+pGcr+hDAf1TyFpsiKBps
n7jwk5Z7fjd9WZaDYMdextzSFDhZ7bi/NSPl21gZPe9/Mk6mvl1DLydYbTwc4R3RWyHeeylWKOKH
DI/uYsgN8QBOWRhKqPVsa9sAkqVaLoQ2bbxTc+TMWkx74F/p0xXyNjTuFFroB9AH7tGtiegDcxBd
KhG8ch85uW3OvDm3zFv1RNKglCr/XYPtEUsY+gi4uKKJCUu2NUWYWVClXQrQBlE3ntVYjlRIXAYD
sZTGKk8SbADXckCmQHaDpSfyzNmwTu3JvJDCBxN8zkiC8NQaTUzwv/3/fyKyIDKOdOQ07LB130Gg
eMlQZNF1YOntecWR3KC5YKnB5MY5UqJjkODut9HhA/3Jt+nGajK0xbJjsydU1nMQTOaZLqDiFJZ8
0FYE8bS1YqHoXB0RTWGe78Hwgxh2bKF021/k63N2QfU5uaqizZ09pcOuxSQN4G9aHbYPMbylJxb7
tUuapscZ+JImHJyAWINIqATlpJDz7tx76O016MMTK5h+DQf17WGhK5nbb66bSFkzf0c8m4yI+ODb
WU4n9ds22h2ImR8y/JaE2beOAT1mM9uErTriRqaFOPckNH+M3r5mngL0wCMya9OXPWi+QnuGq1OQ
XP8/W5p9+ly8rPKRSWWWuwiXL2idwNIE2yjw3uIfFXIapw9dp9xWbwT6vzft+22L98EnlKnU5tjY
HYW9QpHeIQJVo+Od5OS5LdV1sBdMdTgGfuVFx3G6oKqoVBWpSSI0C/qa5pY3jdVE99B/VaH0ddkx
rwua1s6hfbZLzMKDLvkZZMBUTOgUNH3+Arhm9skXdwhZlaJHEJFrEfXpxdHWgE/d0tcPO9Q08NX+
lLfG7L4Zgs0j/Cl28dtBCPzNMKBaAjvyBbg0uZZurCGnANKjD+QUk4T+3LU+Vo7yLpNZLbUXZCiM
DOmvVmfdDCDRBSI54miyXidDybxASlPYDzeY7Gsz0gV1c+dxVzSyTEV72zay9pigek+KTe3eORWX
D8R5v/pcp9IZCaydKiut7S49avz9uCRNDWliz6S9tZwP45zhcYaNismiefVOdDdypUX8IQAFzOYA
PjviuUFxEm6whVzlV5dKitrXoft6wxSsmJZYv+vpKZdSBfuOrx6lrlF1/xOAKVdxF9pjQbIv8z9/
YxFymW5/ZuE91FagBov3X3Rn+tnstGjKuGeluA+Hi9ZtkqRR1SxvJ/b3kntuzWYRCXFehKnGQZaL
fKFoVk4sF8WnSqEegAQ9Gwqq1Ky5YsPSUtMDSK4HW2T0L968U1OEJ7jwMcsd/PmCLKivDbWVUV3L
RYwabtk3muF6rCG7LcIUqCcmNK56EI80TjB8uWHLyr4myOm42PNt6+8q+DYTJf39cv4zlN4Uiu1x
KSOhFVWxfQC3+2bhzEsn1VB5TOdFU8mKz1qEutSZ9T/ptjmQbI2W8uMR8Xp9dRpRldikm1D/CIqR
T+/zmTr3QDBR+FqcULTOuKUQ6QEoZ2azCff+bqIEr9JC04MRjjEazfDdJGTTO2v1ncp3JWBfOTxi
feC5ZABTn0wD9M1imZNb+F+gZVQSVn+G7KU8xTE+5sgWD5/CYXKXvV9WunJEPDXkICXVudVWpIJS
vhC9ifa/L6rH0yCUOUMOuYaPx+W/PbgnMfnqqCeFLTMjvstJGnnocMzBrI4vF1Au+73no2UiXmxN
W25mcuZbzUeM4l7E08apLectj8PbK89dgOlR9p3Uw60GbKIDZ6Jrb29C7Cls7RaTC+Msvtm+hPDX
8famq9cYHej25FW7aR983dnnZSGH7pJDdL67gx7e1+c+AJiCY6rGKYsMQRz4li+nCquh8ROMmaUy
aeq/ei2cmBOa11VjzywoJKA1UTg0oE5wYeZl4ecaQOA00sCdgtIuWuMvM2mWQZUwTv9zcsQTykdb
5nPs7KRl2bFt631+B/CN7IsDLiUoki7utGIjftN5Qm2H+s0GSzArGO8HBzD3EeTYD1F/9PR498Qu
uwEeYRA7rWtpMUoW8PuEU6uh3u7UI9w+hl37uzjdxOLLA8btAjKu06YbTXZS6uySAeFlL5TgvvEu
3XVqtx9/ttok0KEs5fTz+6AeuiN6eTPg29jJUxsCpemJ2KdQp7YNp6sStl/EQtig/EHlsxTqgbss
icMTKUDZpxtRtn+D/XKQBtz9Oo5A7nszrtvcp64D18jfDPaFTgRtyODfcbr+5bXmqfzu2gagHqAt
gF0rq7cfw9BxCnznX8c/f5z8Sr4v6B+xTMxJ6Rdw+iy9+1Itc1C3P1ojgxOV98pR9WwfvovhJaTg
SN368vW3lC5jpmJBOYKkxKxnUMAsiXaXLln5fgXBftQEV+1wsOSc3TgKrNuY4QQ2yQPVUQev8dkD
sLi1aqskLLhFb+s1Zgi9kFx5lkP0J9sIvzivcWMuj9o7m5373hYwhIchFq5olSimxsXf2N1nLgvy
SXrrfT1B4V3pv4VkLevCcjMYa6ORl6QxpaKutOceRhoffxWD/kNqVmEYhlyLnVnNuh4o6+ioS7j+
SrChSVyMIUjjE8LrfOu+FKqawPIoR1fv9qiF/AFQzmZVvj5AiO2Z1tv3fWjY1Lf5XCfA30IzQ+AM
wf20aJEf2+1Ggx8wOWAQFGpN8GAHelvJivKlwhcWbE7rp3BVs/tBE5DB9KbsJvr0Zt82LHPGsq/Y
Y/N7Hwv45/Rj5NF26OLNXZxJGhL1LSBYEWYbHYKo8ARJd/n6pypCMsa/KhbUi8G0PXipn5gnH+9l
waVr3+E977jKTTLrrtfLr2K6rBeTp1g4Cm5E0FoiCBgwIo0vN++61DpCw1Jmr4rs+aWHjs8eN0me
CEHLBmTsoJ8cL4/3TZnw8SMxBE3GFr6Wl6OibOP6gfWVvXmX1qKyyoQPJR3jN/3A0rroEJVmWBJQ
OeZSvOsq7JL/2AIpXUIzL0OOQHBDVUoy4Mq8hnN9bKuaCrgfbX+aP2i3Obn0kk8EdQuqWahmirKI
mmujV7W/nraXs7dggOh5xigQrNnAxsXXWCUPhcWktTTSA5l3c+/oL7Fo4wc28tQVOM/3pI7yLux5
fHBFGUJYzIFYZZYwwfwQxVHpbXzI3C5FgmS1wM0PSlVedraASqUmCmUpox8r4JT+0hv7wpAt5U5k
cgqAb+rz9P0ltu6wGhl1ekz5spuYoCR0i4EPhBJqpCdn1Cn4yyeal/4xYSX1jtkr12Y6tECmKqYC
nx4zMfvFMa6Q8XeU2RBG7FtydedOgaHt34hlvDy+VkDnkleCC2mNx7jr4NCB30BivKXF9QxAWl1x
R/arsmjMlh/0qen+b7Pk0lRKOr0Lm1WPrBrE3NdYDAe1u75i/Lxzm8/prPC+e2/8BWzWf1dr7eVl
ZB73UaTCqLEa30ix4RMjgb93PWJJh5PUrgeporRt/GSUbQqBpOrAhrZ9Ji6YS2+J51TSc0e6Gcs+
GOWCeZOoaCDsdtjyuBFWlp549KQCPrdIUAsIiva3W1vCT+gIGgoU9Mbz5hBAsZYxg1RJJUQcdMb7
0qIJTjHZK8MtekgeOXFlDCNelDoZ767MQWjSpifyJBCFjdIYznKfUlQY/UeGyq5inQM9CP3MHoTH
Dd+pcUDU0vCfa7VfxVJ8hmFWgqY7f2fDZwblO59/8/iYjzsSvrBeUmsCBn7NEU1Be4IzFfZDdc7f
lIXskSCLYcXuKlTJK14i6iQ3IGcn4/+OcKrlY23ARmy3i7dymzaI2Htj5rRack4q8TImdVfpvJWE
deMFDs7hsXopu912Wdp6nZ4jtxpB0F4go5RsnjGZ6b5jEF1wGZsXyLxhdxtIf5vqXN6e01UgXDw3
N1Ayelh3MsJSYWFwVNmHoSXx3TAGXFVKqcPrbv+KznAmPugdUWHGFFGEHUXoTCU13A72hE2JkKPn
d4ilDEXfuKUNwFAqKb9SZVo7yiQqVpuKZM+3hgHX5baL2ofOkSbMqjQL/NnqwMNv8KD7YB5hkqny
TkhWl9jmWG5HQZ1jpaWcx1VvIgLi85VgG6LNUhinIF9DQLbM8Dejh1lJN4xyRwrjdUfyo+3Knskv
/BGXQvEBa9rXuX5GYCePB1gyl5ggZ0xAFM19LW9/elJvagxAhrVh5BT00Iul2Gx9UAJk6cuzw4T/
9sWV7VCg+4bM65kv1Eh5Gn3yB4EKBRmZaUogsvjflS/eUGZq03J+kjP25HPxYDRG4jAkxKJYKn0K
fUVzG20q1I7aPhogs8IzHU2PNwIySoo9qT+TjUFolKa0zj1v27JmO5Yi+4fcCIXqxjZaTA444vYa
ANyOuvxdDcdY4nDPEbsmbyGKP5IYoBaVHf3D400KRHjdkeae+vgVURQeQawJZjSB61VdZVsy16al
hnq9+MwMMEsljGPSv7igmr89X1khwJuKF4Lmb4p6cxgFHcpHDDJ6hyvXizjd9BuUe9uj3s0T+2Id
xdd0ARujIFUoqNIfgHjQG9mmSZVo6tufaDjnZ64mDhr79voPm1w3Qh0GCPHEKieSbp+ev8SPZ0fb
D2VDJk6tOhgM4J3lGiE73xLyEwvVd2h7RUQ+5tZLqe1fMPWbVvMLnHw1N673mOMYg9HJH9be64gF
1AJwyIEB9b3wGV8xHH2+EORGi9h8NzhsdLhjayDWOkfwK1OpnwqSpme+ye+SMjeg2mdgjfGkp0Uk
c13v0R1Z6+nK+u3ZPn660SzXmmkJx3r5g/haVtnlZbm4N4zHFP9at624kPWNKGNUTx+ckWnudMUs
eHyNR0QNa1pT3aJ4lPucx9drEmkXPlhTAhyPhD2KKmCibnS/gGYdcVpVW7VjTzavfxdrwA9jdGj5
oZpU3DhsVonDUbqUNRZhwL/9WgkYth7DNEAT1W/YAY+/w4FZnRIVbctCRwH1oapUsbJlETYQMxgS
050SR5sB2zhxur21BOqtPuSxbHL95Sp5QqlDBCuxEfcoYR/bGpmnudlYI4C681pIXtMyYO8dBpgI
wwShoD6LznhbzlFla+MFZEmV8nbaDEMZaNrh6zpEGT42Di4oFWc6V3yWNbjUsVLWyiFpyZKJ8THL
aOQe6B8+7EH6A+5D4fh8GmbCYLBj9qIBECMgaInsdQst2MVLBxqE1rjebEN05v/YBomB9eyr6gb5
FGOq/M5i/1sjTCW7HuAyMjuJ6wr3B/36dz1XMFvjxkm5uJCCWrOuWA+b/xqm6xmN6x/5RkqjPbeE
KX0eSknQy9l1AAPFuce6s0r4VEy5Tof+jyGyE0BRv1Fa2MfNTQOM8V33X1jfwFPXiLTIutrylnCI
zljNAFyzw5Hfu4WpqzT/h7p3HyT5cROK9Yl+oUHCVOz3NburYT8Qk8bK8DeXMVgz1LaMY9BBk54H
XhsZVjsGrdTtX+lNawGGouHVoKENoE4HqSc3lh5z59Ky7aF7vdvJ25IQPJuUsw0jH3ev2CnKXEOb
Deehvi8vnLLjc1mzJrZS1LDF5JZBEaIRAY3cJclbYgbyriPNkpho0QoNc91Y6gn2DVujWf+hocyM
KUFxOZyENY+Ob9Ejk+wZQSjlkzL36qqVWzextlhQ4A+GpoQpe3wVLVauZ4UpaRbXKA3NWC9l59Fr
LKBQSRlkpYwc2VrIVaT67TobbJtnzpFPV4Si3jTr/XxkZfSFXfZOerPVAHuTscO2+A7vwvYBKFYm
FELZkyyS2e2g0t8GRSCB05KGBNi4m+lOOkInxpoUM7yAhwG7tR59cJzTCHXUDFvSBFmMyrYthJeE
asqETtWdIOqtPGYY1JC05mr0L35BuxWHFd3o0rUOndN2DwcAG8/aAgko8yQ0VGN1GzYvbAxvLeb3
bIJoy1TMgQGDXaOGNJ5SSn0KTliB88S8VVMOvw/FJaoRnz9pC2zYaEzEmloLiIClFN/wwESUunYG
zSa+GHewupV4bjC+H7vwBNH0KHT2BfoplpTelGDZqkCBrfjgv0LzUZbw7CqifGXJHavpPzh3i43y
tESOAxExQqpDrYkNphJB71lIVnecdkqCPFnFtorRXOBQvFVAH1yuHYligzmNa96b2Do0GT1uvj6p
5DhlrubuRecQBYWNzoIFmhTl60W7++pSZSpklleSR4ZGvDhjHzgeak8GeeX2/JeCLigBdyLpY8fH
hX9Xbtcxv3sAeDeFwOmceZSQNZVePoIXdqdgRS1AjBx2nL87UKXpsdiE8TKKhnnm4FOt7iTowFfz
f7w1rkIlhSTXde/AjCO7xSpAGhKqC5du/CK+t0zG5Ww8I+qImZB9xNdjSXT67mVSfktgRk1KYZxi
3rT9xadl5vYb+uV8BPqzioop4/IhmqwsOjIu/5zE/9UKWB+ecs4LPxuH8ODkz4dUncn/vRFX6UXK
YQH2319VYk7jrl0YhY4d/1x2qahLy22yRzZm0YTCC5cvK2S1wnCZPMHqgiPgGRQmyDDM79LVcTx8
KLwAau/upHHu62+emkVkf8a5h+2vOSiFnvQrdwlaPjEzs6c3a8jqGoDz8IGd7U5Kg+7iWuQs8AG/
qy4EMBURR54rZvT58o4Pytam3OXLvOSq3H+cDTnKFaWaT2xTaRyIJgxs8f4fGhAAfKtyhZEuqz7C
ecya849p2mYa3rOs1EvUWjGesIW65NSnDuGy0EeESj/oYf7LVRwib6uhrpoSoCD4wRbMrUWaB4Yp
6e9u4Tw6Jy6DCi6ui5Tk0tKQN0d6r/8M8gxSVp2CJzmrFW53L26Ah76fhKqVj6Io4WL/gFbwBIpe
LExaiLy4hKWSCyQnnpdGvPaDAyhw7RgYqUxQZ43YrexePlyVpTaVDm2OM4lU3amOkMyYOQ796+8M
Mp7zabRnlZwfPoIwX7L28pY1S6nZaVidUPpYIMfd+RaQ7uxJr5bF+Qq6UxPra06uKdACHOEbfEbH
7T5PT7Tv38iiqEHeKGhobRz0VTlQJOz/ngDuNL5WFf3AGVvrDBeQD2igEj/KIIeRi2Xc7q8mE+1k
JGRXXv+GUzaH9rh9ExaiESy0nwK6KMCR9Fc9/j5sErSwSjRne4gIAfoYr1v9Q6OU7yIgv9fgrlN0
MrnQu8XyB+F/E8gtR9Z6OjRJak7qWMNOOn8QhA2sikO8WVsOOzjKzhrg6rwtMiVYYV+3jmTYPq9K
l0ghcg/BS7y38JKGqi+qoURuZFQrAgWJM919M4q8iq6hLcWAiY/z722zH8xcU78D11MIP5bngHQ8
VIsF5FILyF3+WnRw7Jj5eivDnQ4B3EGWaRdgJlH4csv99wPpRXKnJlV1WqOVLKfWs7aFdyJuGBKK
WR6kmWJFK8bjZAS0jXc0tDej0CeZUYQC+8pV2bgfsj9WNDXWlz4e/AA6/ggizSUwEz9OLKTlygYQ
yj4CoJxgNd5bNnmNzb/YGcsxjHrbZ0DxoqyFM0YJt6bh8StMkNinzjBSoaxAmV5xvGipkYTr0I9m
Vnn2tl9V9WCSRM3uc4oYNJxySuQL2Edz3CTuCiUToyz+co6M3YKVnmkBflppZH1gfDKSg6tN2nPV
BUTfCUDVycwcl/VRvC8wEnmSj1jWzVI2aomARx/WEvCvY9VOgBRUAybpLCNLUqGF6pqGM8j6zt05
S9lqzTva4L+ZuInZfsNrv7AbzO6y6u5gdm+bY174xfnXQ5Ho/CaB+UVAvXeP6PaWkG5sEoLG7rwY
hAebH/HAPmlI45WHQOTfdRgRtM6NQO320F7Xdd7DeqOm5FrmZHrYzpMtw9DwNOszkWBmc0MRzmqQ
sPx/Zc+SbZa84EpBu19JYhgGxcOgmBSYD7hOtl5MuBJzfH/7DuyCj9zBPMMl2ZVEfcXOAArngygK
c6OKDuhLJsJrOiML2WQ2njnWbIbwt8EUREkrJBh43Qe93OHJSjuuX2DTs64v6cPefxW9blm8n9sP
Hbalw900DsUOobxboF+6T4whCJp7X4idlAsKjzg7jBblc1KZXHsIekSHpV/5jpcLeJ0umyDmE0Lp
/5j1LrURaFZvUEEpKDO3cqNVk7pdh5amNNnMMupi+0+vt+HMou73VWes+vlD36flSrrCf8FYH9Lh
SyYppkIs/iJ1ys4CyR51qg2wpyb/hmS0jw3tSVf+idJIUQx09mfSjNGPM14lwrYIpkJ0eiPFbjab
HMeA/h+4kvsApWr53DdXSoD/RL/uCT5AYYSV09WtbDnAI5ZsP1jXaGwKYzWLW2Iy9TL976+GEqZS
Ug8wa6gWCwjUhMfCgtNq4O4f/rfMefPM6EPbVluZ1llwEpI42lDBDHJ13zktvwoG9762UfTq5WJH
o4kmyCG85ziS3V7dOf3cClXZ9As9H4YmjMQZNbtYhA5qL9av/3QUME7LdFzw0V4ngp03xK6fJAHL
Q/kF2uo2h6iF0euotdizDjWF1Q70GellVo+jUM7bXNDZtgbhspQ0mII9E+rLp/A1lhAQRDSTjo9i
PSyvSRHnviN1UGrDc864nNH1YYVdjyO7J4yUHxAL+I8rwqIUHLfTI45NypiX0pLZyDCgXdpnYkCX
z1g9y8vojU0jo1QcAQ1e3wsjzeLjTSkgz0kcfo+D/ADzBYM94K44/ZAr5f677u7g2RvMHlbn2+St
8Hs3eKlXEOOgVQvndRkkBJCLszM5aoEGZm61fYI9uScxsS18iQZBdY5Byq9CsK/BXT7xnSr1u6YJ
DmKVIpNs+uVTPGYDPI3Zy3M3WV2s+b35MLThzU8VRmXgbHP3IU5BIifxPloKUwGpMoP+sc2g9uEo
2eKl6bCB0weafZ3mj0i05lilhW/8WXWMtK1y/TZm6Z0zlqb9oXBW4A8k3N21zZRSK0qVJEMlm+DD
dsHadIZNVB2tNoBAdql8+O8O1RHA5uPJsKIiWq2mwYFDq4MtDF+z1rz+kRT8BZjzbh5ffEaTSt6u
rTu2a+q6nDnXUCo6fs/VMcxOqspZH3F3wSYqdo6vsYThQ/x20bPBv8V3j5oo0WzzH/h3rJTLUup8
oQDdtAp4Xbi8lG4l8UmvaOdK1A331QasBQFDhKPpwow7NzHHHDW5hnf77bPYgEcOdxGYZ5gXmGjA
quQw3WflfickXURZiV5ANhgr+wNhsmlZGvBGGILbjYe8/1ilYysd2B+vYpHI/RFLoF5190S1fCnX
tG5lW2uVVuTLLVOwGjqSTMgHypTTM/QmI2VibprzEsyalpLcHfWyJxcOT/Lc0H+GiN/gdfseFORo
0Gu0R5hqfUH1lFx3Zu7+cw+4C5ygVUhKxCPReJWPcLEtD0NJcVh4l/S1EqVRIkGMqM3+JRcJxHPT
3mv0lujiwEnQRGYj3adMcTLrUbzOGQuU3rmPRf7X8TIU9TJPo1diECQVHMK7lTpbsaQ98xgDc/pJ
qfaGsFUKKhrS06fcRDbABd91l+E6lnJ+H8LZF5Z6EXVvvMC0oUokkbwBo2e3XQCffCa9w6taWCjQ
9m/vFxN+osuTmBLC/wtTPTvOXjT4tiQ0vdzoYObjTq2kVvLhjQVvHiGDRt+EKGafuXq04ctL/4cf
BDvfqwodwCl8CAHE5NQh0Y3F5OZS5P5uDZneDp1qQxs0Ai9o1kGvmp9jet3rzaJF0O+YuGnLdHxx
5gc/9xbCrujPS5m+v520iT2LTN+YAxTt7Dv2q1dtBRBFw1fobPk/aD5tlulUTAePVUbNlV+r3t4n
k4XXLBfFZdcN7soZ1MC9CWsSjzjK+f39eCNzceqr8TRfreT4G1RaKZBHI82X+kNX134PHwNpnnU4
4ZhUHkaD/MueZeueKzOXf686kJGGurlRwA0toDKGiuiVxmPUjsbms2epoMaczEBIuvw5QtnOjIpO
VZzyesJLBBNgl/1Hd7d000eYj6Tj8qOCJqIa4Z9PkGGSdGminYAyK5+r17Y+E4ElHa2pDJg8vqLj
fqIP9+vR/+RWa7P+zcymC87YnkraZI3vPld61Y6MdOPnQN/Q1JJRV5e9chG1fPD2/bnEw9/4O4OI
HApV7XOtDYm/dmV+MPKF9H6cdC5XleZIWISCKsfEhAoyc3E5fbpQBMsPYuc1Du3y2uheW8VseNR/
2+LVQNTQtloGYDfCsgGZmMQvGQX8j5Kr/9jhuhF4HSYx5pwx3o1kDqh9X8xfgEpHte07Ms1lAEO9
8mHZozUmaVRzX5sPuLc7nv9rOkR+nXjOz2OVqRs9Abz5Ekw1MK1PNvS+MYg1ZOZoZ8sKweqFQ6RL
0LS2G1V39ZsdRbyhWmdpn3vuV4TlZ3JBSN3ITOaY77lMrmRJf/byVRJJUHu1o5HKRO4mJ7CLbnwt
eqMB3DWBtxMeENePGJxTXNZfBpzAZeNUkVYMnhSIxdNgAVOMENa4C+wbDv400Ypy9scQhHBH78+/
YSkIF/MmIXnl2DHA6qbC7OJjTiT2PSoi81zdS/PcrklQVP0V/5hRSOqp+i1KxRQZuR6Oyvcf8LR9
bGI7QrDgCmS00U5kknBdqnTWQzry0/P8wilSMWadyZNm8B14A6RLByzwZgX3FjQH9d3jXxYN95Y0
MCes2ufD2GZec+mOdLhONjaQATpGkApFTwle8QGC2xQLjS8lMmR8rNosuNh7dsSj+4UdgB/xAkpj
ut0bE0IBCA4yCHbLlyCSDknLyVTbKxgKuICmpkIWySjxu70GI2nKpTTG4erp6qv8mcLkWr92cLc2
TUYlMHZFj0gSDPQPCMxpLFPiD0E9kPWh/0bbJlyICzsC0BVhg7SLuzfslsoIhhcTrKUzu/j19Lzk
UKlpbX37tD/ZGU/E/S2qiKLlyfeHdsPyI9xVPZzgbvXCQjAaFEdZ7DnQyacLuIXESHfOVswjUyvj
rjUBot6JrbWTz+oA5j779WafSWUufvsBQkmbCtTITQ0cru77+QF9wG+U3K3AgWg4jKFdI4zKIeRI
Oko6PDlEtyeokHF1s4lS9jXl6j7KdgHjsGr90pgOJQKEBG8iDfNupC5KzulF6aYX9/5xN2aE2B1Q
gRNWGzxh73DiK8ejXtDwj3i2pF2k1c1WWfA/UwJhqsDkWHyCzJnT9lPJmXN6qOVL9fBW9xx+kIub
0V1DYDZO7Q9emMdQDvWvAIFF6LBozjhNYnn9d//bsHXPAibwtd/Tw6uWqFYwZNHxMCBQet1fADzu
Pg1Td7ujYomaJn3BuqIE/0udB41G/YoVV+K94/3gmw+to1c4OnGGWDW9MXf1+DIZ3IijodUHApEM
7z1B0aXpgeQQ1PbncckDz0t6c7DWhTtJh/3euokFy4D9iQnpfAc2XeA6+12Bth3ed1ZJGokAeT04
5ljnNC+RPC8nQaAwfr5dXqdh1AnvwW5RmfmMlwz+yxeyO7m12TvVQhFpWNcGXsud3JzgVMiFlyTd
o5bobYBYnwQLlBduCU7UlG+x/juu+Pz4qLqFoJC89nSZtlSuI3g0sBM5d40xx+FC4rTdcNFti5M5
zaPrpvTrwpdAK0QxAmFGZJX6o4cjFgMemr7801OlubpwIKRwcnGuK1+DyaiLWp9EXjbKRSaQgvfL
EJ3eRRJSZGGiqU9SRIpffUxQoVcGceuI5ul2WuuVa+73JEKLFqPvytkGmQE3bjBWzBqGKQTR4+3z
k817ismklxwXQP95bYb1MMG2jb3qO740xI6F1yqMfXSY0A9pg+vFp//kZTurNfmvJ4HafkVpU4Io
YKhDnZzRIr7KLqXZ691FN0ynHgE/cjJHmsDmlvwiJlYsn+KEFJOp2gRB0kcryHAdzKfMmoyBthtO
yD5h4kJ0AbxPEEcyl5XrtTF/+Qeo8XDug12b8sT2NGeP7B+yp2lWcxLPeJIvN02jc+vp/bz/eXB/
OyBZoF8L5PCK/j7bPja+5QBMZtP3pcGKxw4Memblc1SiGzTlVXJgYsX3gWItqS61Y3GyW8sK9SWY
RuTc9DYEJyrSYxENrusGqty8HXKbVlqchn5JaFzKJsT7JCMNE283UxZ8THKc307nXJKYQ17Z7KUQ
o7WBsoQOVTOaAaCNupEejiGkyNfrJmtssuPeCgkji/jOv8q4MOe/GR3SbFqyhn/Lwlv4Wwqoz0h3
LRzsd5OdTkoDMeNGdhRPq6N6wY4MAufBkbxwVMzO1dVs6NHuh24NH8BAGjQ0TP0ED+8asQFg0+rj
kiDRA/TK4m+hnpFwi4EUAPPUlNRq4+ahmXEVQqqFYofDaQ3SJIXUv5Tji628zDPrja7inWdikakc
u5pLM6J8BwfZ0ps4D6Tzl3jbqgfQEzti7z3Cajr7iaFFCrDgGe1MTri9dt/sHGBezIr9iY4aZ57D
+n1xIuW+nk6tlo7w1azvG7wVDwn997zSScdT7xavpnYr8Q7pjEUEX34y9sz9cD/nGAUVzUo9yH9A
6uNpzlxvf5heVXmXFTzzR0JAbqSAFcEGcj6dn/FrnikgTaSnQHQxrBxQ7/tdLTVCyg+quHeIAUHV
diXAu340ScRKc8P/GZE7E/qUkjKvJcJ5rKBjJgVGaF/BqLhSkqeCJobq8cl2j7rXpBpXGiKw7DyM
1a+fPKk8uqKCI+C3hjTxMcIAP2Jl1N9ZVRSSbD2v6A7wLdZLdmHC3RUgerE0djOSPV/JEP5cuGzB
Mp9azX5ra+xO3Z3CfReW1PZhvEZz4cvqiHgS2brHgMykzItbko+oN5MLmZPtZkjvi7BA4yYWnPKs
lL0JYeWY6uO+WOkkWEHl+ko/7J1MsdILryGAg57KaoHVT26/ipsdLNz4S/uej88qmnyn6Lk3affX
erPtGW6PcOH6JQZIXYWFR8SULaMngo/Hplx3iRx/02dvNykf5xR846xzcsPFtFLYQoibv7chmsuF
MduwyvqFS22CX7Y7btVZrEeE/8+kJ+B0rbQhA//WCNzabVQxmxdNk5Vex2uGFc8DgXgZjDfQa9gg
49wbDJuqFzyYU4EDS+tHKZunE4kfwWs3sUASwXundFXaE6Ekfx27DimW8ttDZdWAN2s29LQ8X4jJ
UJJxO4//E0yEuuo3dwGGlHZCSC81Cybt3MJDrILNDBppAJV8aEioaKon5kJ46Cw/OA68jIGZ1Wfe
VNE0nEW1kwrp4YC1ufdgQ7HYhIKz98qwl1qjrWuSU0PvPmCPz29UcmhsfPcNjrMX/Fg1t94zs38q
akd3xkuP3O1Dd+MRtILvo174NDU77R628UqN3jCiZdzcbZI4LnZsR+bzC036Xu1v0dYChyvyQefV
Z3gjlbM6659dX5Xd5ooS2aEZL61pyQsyWi7tzZnRsngjriPezzuFK3OTfMN3HuUi5Zc4oLqncahc
zs2eMw5xBOoK3f+B8ADCZzkLukWdgdK3F2iNu3vAiIMvCz+QhG4PCFSyy0T3CJTnVwADwalEmqvw
E92YzDyldjwiSErT6Qy6JpBXeAQNnrqnLHTSEh+CqkwNsJgbvFMPXlttSRQM20JzZBANuIfPNOr4
OL8cjDu49a1ZylCsMkmyNbvPt0wPfEOsWwN7qcMzjk5J3wl/eei+NZx0ZqsyTdEzPgm4hU3PDulD
KfJ/J5HO8V6QogVn8Fx2N/LKctf7nh+pBC8sncIKiGv8NGhtjgw+wS1g1DeAIP5eqMK79HOVsSwS
7f3EjlwtYtB9mn0Fv8P0OQobqElyAiIOz4X5rob/mAZ0QI9Ad7Vuj/yi/k3LHjz9tz7CoiNdTR14
xgKhM4ecv6sVD3Q1hOLklgQQSfljHyIvZGAfOJOOWH+lg+CqFC530nbeCFr/MMMEUgO6ZlUz2PEt
rnlP0jl/DsgoudGImXmYFob71aif7QVJ1tfSNTeIL8/B/MsStWq9dHVwRqIlEg3F3+nCgZR1iJ58
JiLtsABxx710+E4ZDXBd+OX1HJQZl7nB+OD25VkRESnkZMQ0phx561NtVPZLtV2KYDkKPxKVR6zj
Hs1wb804IrytqdDGogqkqWEN35FPuVhEQfKdzxwlSnBqsMCXF21CTvI+QhQugU55zBgwpuf8bqSF
cms2nC3NCMiXOi9twQ7R4U7qNXVcomkXLhuB4S9OBWgN3n23kf7Qu2nC7FYBE40WewCQRwjdE4Pf
OxAFN0bj2Y+eRiclBXG2ZstdKGEQnHxOlxkc088latg9IulYynYy12JHI6K6zhirr+9rbGIQh9Uc
bSgN3FDM/FHzyIYht4M6E1UrwcvZ61hIn7NYRd0IBhj94SnlJFCPB0u5wdBcAmBtnANEEf5VUbHp
g7/ogk2uRI/np+Ysp/zXlDAqVwQD02xlijQwaq+sx5l29sX8IRl+S9Nz3fRx8a8avCZaovTQfgtZ
Nu/E4wnzC6+RzpHiysrgnf4ZmCcw3U51ChQk+/Dgw2XjC6aBjsUz282PMb+18MpE8Hm3Uz+vvg5Q
WGENMcMLjuzFMZXvMO62P2Xkn02DzAyJStxpxr2bC5nAvd9mjuHe59CgDDFy4gb0/EQ5inGm1yds
RtrodC9nYNNbHHGrW9tAj7BPBuzF4rkInUvO0LfQXFmcCDlTXeZUw5Pieu+9npf+Ui394h++AGUY
USaPaI0nDcSL8LtGYR6IO28vO0Yt4sOsPdz7EkEoJzOEzSbjtgnv84ynTV6ko6DTd75dra3dpHb1
+l6H3ne7hUvij+cpnRNvHz+f9gHyMn7xJHveApihK9p8Cwi3AApx0CR8GawNM1RtiFl3X728PPJH
G3weHoRu8E5srJx4fF5oZyGQS8UVUSI4AC0DuxTqcAXbCgBblXcQTIhTknCg+vFSBELEEg2FJJsk
1o37CsX/bxBcUQexyXVcN7zMUlRnJ4UaVUQFB2ZstOgAjAa6/InZ7s6f4RL1VX5nnyV86zbJMqg8
YD3s6drE84OdTHHdvzeIxow/9kU8JNujKzEJh19P0hUJA3HiOAPRgzVDRpOFerbcm23XOAq3zn7P
h8P4Il+pHEgcCFM4c7CDaWyp69dChlepIjgEhp7Kmvd3kKQoaXkKFgAAcwyoQKChLkAKWj4hHErO
nYxyuUrIdurGP9SCugq8XUk9Dadcyj8I3EjiDYAaKZph43tEzHi5YXoSSDAUabFhc/yoBQZHFSDX
7EGQawR3vaXNDw1k6nwYdkTTqpgedcLg9Yn9UtTmUMkwIX7OzN/26gRbLtgkLYrhzVE6KZBd6O/c
qCVJjihox2c2Iy2bNwpI1LybBy89PxcCrgWgX1W1WlX5qeM0kumQGoVBh8H3lhLg5coJN3yd/91r
WCJtO8fCwZN+8VR+0OqF/2e6M7IBRtBXG6zu+AXYYa566OvyW6iAYSzFnSRT5aAgbDRdbUMn6iGL
xrC/NgKhFasIFMhfQtI7e0GixNVKW0lYMv2qlq7hiIXNsL4yxRS8ql4iKoG0EJt0Y+Nw9sGyDrsI
Ko70zGouMOXEdUoVsV1zxd+OO9qW4z2A3h60Voib4cgc6ZoMY7gDC22mH4MVHWpu0HwB64V5Wszw
5Cm0u5zBo3qQY+WnArmqBGXvDale7mdJDFKozL6yzCobu8gEE79kmiXIzzZT0YkbzvSs2aTQqV2R
S9gNXIycUNTvXiAkjs0bR5Og0juGZcbdoUvkiZbmJ6NGPMdiQh9QZ++0rRtoLa6f3yajqDFsbQMs
xoOqbAgFIkg657/K5/+V9/SRnuElfwGwF0VTLNor9gL4qqA0oYPXC1ELsFEn3jqlz0r6PNdYhlWn
Vzs1/zR6iLXqa6/qTyguuFy/AXWC+u2ITKojt46XSv9HJiA5KzTwFP3cHAfZajyN9QO2L/ThY4Pv
et31YvblXKhndedelJ9Fm4LIBJ/dEOXDtqsduk8eAzOgqADxikoIo0CqqIg5/E/hwFHwRBCwISFt
7BEA9GiK5Qowua2zqYX5PfkY8FaKhhVo1WCqvWkw54SDIbyoBNoqcl2r9vyPKRQ7Xtj62Q9VG+6l
2hYTFB3//xjEnZpItSzRGlVoXKrBIAChEkuaaQkQBo2yNxM6iyncQ36gnrv4YL8TORO7zSJ6fT4U
I8UL18sooYrgZXdoWV1abNZ/OBt2FR/rUsQd5/EH2MKYZ6LFzQL5zE2NTTCqduyvHZVosDErLVUw
Jur2GhZ/hMb1WwsGlmhKr+0zw+bRq/LMks0Xkik+/HIWnRZIDVfPUTOzjK4QARzWw4UroLO/niFS
FgZcKDv29myUN3ppLwRqyGsaxILY7IJazu8fF3NAi2keLTSzWbFBU2iriakiwPxfo3nveuigTpPf
tGDZCqEW+YKi7ZZACdPIsMkcDXmpqca3uAFh/noY/e6JMeHZU7fo0QKhfUVHlXzoSI6Bie5sIn6i
ZVZHVjX9Ax+mGG3Bf0I8uiEbQLqeBH0cZiWloZ2srJ361mkV4gqgLAGDZ8RhxrkDeDgVwlqP4Zn9
JzS087gCgF5f/frPeIMJ6pfxqWgE7QDHM/+h+PzvdCVI2f/24qQcBof+Ln2kDJyCAXBSa98gSuHw
Eq+IHhAle14DVjMMUQXVZtRmi197nh79gphEdd1N0GQKfIKxl/dN0DDNGfeL7DdMjbjYyneKDyDv
LnXQq3sJEZDln3Y5ANW9RrUncjUQlDujutu/jRkQxn3KqN/pqhv1t8UqhKTFSXUSWJBvXiLIeaZw
tbTdmTBqlmvirG6kk3UVwdvuUhPCaP4pf7M4BPIR92zPC9zqgq4cOItWsSxEac4cOu+ChlH42p0/
J5HcdJ+SaoxpTS3yx6moinGxGQHTIed5sd8aI7Laht8iU+QyGkxyiAGW4yyzDXJHZsNLETonMfIH
t5jHdJnZkZXaC167tMOoY5cbht2wrSgkkodnjw3alBIF0O6Idz2NeNn9CKJ4tOLQrkmYESLSRpJ5
6q4fL1MKX1Q8y98W0yvylgzqoaewZgV2uv55nWdUUgUUNv2sWNxC73ZiQh1Y6LulFmpUe+q+OXuP
Gks+zUz9Aq5dXAskZv98j3GM9YUzy+4Ohl9HL8BzvWCNuHdLdO95X3Xd3iDEn7Z9KzZNISlK8RaM
TAzrcadJGiB2SCXQ4DQEivBgaDUycDiU4ldXkJQJkhs/3XQe2W4FJgHG1l/EYMEcr+J8vtX9j1bQ
1bKW6k9Dmipv5TWUnCZ9H3ZMRS5O4ZJ39uQePC7i4Npph4vPjrJ1m0NUAcGfH7ZhJIuoFnBQOdNF
S+9B+nk15UWoaHmhBAPEr2w9e0phtC5onRTd1C626cM8FRDL79H1QjUsZDDR2GpWqfxUrlsHE2O3
GyKEfWvxZIXMdaPUq8Orwp/rkjl8fZIzqqkwykJ6tOE0DpLVNfjTFrmduw6eE9tyuAM0M/B8o48I
Ppl3Rt3OwhbCBze7XVF+UVEl77WWmYo+oZtqAe2NF8OM5+U+vDcv+rbPr3pQYwTjl87lNR78eoEy
9djjQxZFrlDWl5NHnvgz7jssPhZxkXVCT+54cWJbBde3JdfSmIOMw98RF+glAZtpDxm8xv/Pkm8V
NePQglSTa9UrPEokEut5LoyQlGRp41rz11hXf8UA9l7Weh3XYf+OtyqemWEX1NMlwhVlx2haGsSM
iLztOuTZYkaP66UZKn2u6JC+fNmZ7hSdkaqI7H7vN7bj2dkEpNH6VzCYMJ14DB/jdvpyd8VVqtbY
2fEfn/nOIkJBXg/JpczdRBwostppXFLJxyndPRYCZedHykZ35/5b8ALnsRibpDE/HkSnQT69lWi9
6j0qRZc8PGYirR7QdUzZsnB5DfcWfleLT49oA34RMNnEmbLgIUpr0H3cVxjw5MfxfJfQvUV2q8WR
LG+ZERdSyPaqWahjnO8CqmvqN2BiLLDktmoMemCmxbtbFckv6pYRR0ziNfaQ9KyiuCZsLPnNiC+J
3fIXZY9lUwhCi2P3IzmXq4WfFwFCuTfVB9h8akwOOCKhghy5QYBkrKJYiVrEfaW84DKRqIEafFf5
lGti3vHLPM0aSXpHRK/polDuom/ci6ruaF4llOOgK+WVo84738Iz7aVjqaUQoS/V9amGUKtOaTdp
ZIlUF5yq4LIsqjq14EkTkTPTMCfgB0dfe3WgVEmdoKDa/nv/jCHxG6uKhxpDd2Ba4KGX47Sw3gm5
Guq8MhJhCCpzqSmn0sR5wMfU8pjKEHUgtq/OBI9SYyL9Ggc7p3H4EXMXUK48p1N/Wxd1kU1yVDU4
1xMpQyBuIlKklYNYCjXFUP1CFLb67Kze1jBgcUea1eNOriYitHKEhMujrqyBW4YTojL6xuvIM2jr
3b38OX4PHxQyDQZtdO4je6P2U6r/gf9myHs0/6hW3/Tf62ys0YeLlKF97gL2dtH5dvY9b1dwhzZQ
Fs2tFepjO8pjgRMYQhD0BV/GvFJkNJQPki4a/S0U4s6Io6svFIxlpu6Kpj70RT2MWfLX3ovk0/Rc
QvTnGbOsBLviKJ+KF4GXU3usFOVF3+w6nVk46QFfTrtVMGU0JdQAOrjMBvCD8qgsdZnHfFjaYzXW
L9rTP4aUhaC545i4wHugJre+2Ycof7bPJ6/32pJcdEQJl6J62/xHTg2Un5yGulyRkgIK8cuFOzyR
UFrbxAdRzkcEyndFyW/ZVOCn4sgL8k9wL8cTmugYrOW5GFmyMJT/FVzp4WhgD4KzQ4kG4ueKYape
jKbOZ7I/ybKtro3RLa6TGMtnB46S+R4X3tRPq/fgltbS54P4ehDiqxs6vCh4yiRLYuxCOVXkg/aA
bn6+kZoK6UBoqW6mMEKn+REkGv77oDDYoaTB9c5Qm5at4xiFNh3KMelNH8We6tMYkzQOEMs9lR+N
ry2ergXnoxWT74MI7tqHndk8l2y8t5FrL6KbLoHEdNIrSy/fyjbhXJrfcknXHw78OkUqooWC7Ed4
N4nL0vti9QmUBuJ+wyBcNFNJh6G36fbZqcIMobTw+YvWkAKKNXWRIvZxlc3syO62OOm5vdSV0w/e
y4XvSzNX57U539OEoaBr4XWYTEWF4L7W8wWanFyd/tuHObnDcLuPBVBBGVDw8vai3pYaY7IfCczR
XseOFRPQo0IbUN+hJdh1zcHvtVGK9BGP0u+Cth40hQZSiJaVdJwG5vgoIBZ2DT2A96gWBSTusIuL
Qmp1pRp2etF+H5K+PNatcM3Z94NEEhLfxJaDRHJbxfV6XJTo3yndBxmGhMcpg9bytSKzN18HPYuQ
vNOCpBpD4o4pbbaHLVzVdX1WCjIWh6kQg0W242stcbU/xgpPRJDtUS5nVZRUHIF1VbkKzWXnzcQd
tAb/eTB3K92JtM85u32AjCzhsPGR5fmbOAuVFyzgKOe3Rif45h0Hn3C94+grG8/u/OhB/ZWsHqdR
haKYTCfI5te2gbnKP8Ky6Ddk8iAOx0PCayRa3laFkxxMdmFtF4wTJt+OcHVRtOi6JnLETMr6ThAw
aTH7Tvip0CtflMp1GyWXTUqn7s695nCTexsSSvgivfeLj88NeE7Rpr19HIbGFPTp5HbXu0Qed95p
K6NB8d/vD9Y8BRl/1jRtoeAWzviHayAkv/BvU5SpFNiRK1k+wMiGthmzYFxHVqqM/7dfPQkyxBuH
V/1CI+QKkpYDO5OmUn13B8ELwKAW16xdEv2BWJuJnqLhdwA9Qo3mVHdwgvwnCIhjtUCPZJAfsr/H
zsMP9VlgTrmU2kdgkRy/VOY/ifmhFSv9v3ok6mJ8hzhQyoRWlq9NI3OtqmbvKIqPWFycJOOLG/mA
ybCXXBabePU1m6aEgFbk1QNEGaZ1+wpgojh0v5OSm0+V6VNm3ovHymlEvDD1v2sahyX0TT1pvAxH
RTlym7TETFhdbQCcJ2OK4dCImU7/lJcLcwVYojnUk9Kpr15iki506PDQf89C4ES4iMeo0T+YypOM
Ql1GzsqoJ5nzX1pj7CCSrRplzX3s9kZhTb6ZZwla/UREWluqri+HAzllPqV/8a+GXZ2dY8NRoiGi
ro1FdO9a7Fb14xjdraa+YxRrOGMQ9mGBQqohT41pdKLkBd8lOvPbtOsPwzJcfoEHoXwjhhVR6K/G
Ww1ShhsDH2epMWQg2Q3v11j1uLmlhQtDNnMt1fRvvqRnV10grp237KEGrNSa6yNWWsKh+FYlfHVd
7EgCgPWQGsdjARi9vYEN11xwU1Lxgo/DPbY34CSRSmSdv/YQ3oBr/km8W+RoK2Conk+oVLg/OmHS
0bvSm223naQEus9Ms7zX5GUd53LEjrNl+xzdRC3JXymjaSV/k6WrpfuWxRum+n+CJi03JrIbZa9S
ydWsdXxNuYj5Np7qJwuep120HVXWqgmkBhOFlZ73rNZ/eL4TQUhfDZ1KyrBip86eUUgZI0+fuiOg
Xw8n95ZEPZaJVUt+Q1HO9hgBpEkUDYi2/RQZQs/0qbAXSi3dGcv6omMkS7IBkAeh76doj2mkFrim
nFuhkIjj/orYKl2ISJHvKiS7Gh+ua0qXEYfdrbGLeS8LWUNGwIVPe9hUL47IOTxIsKIIJeHhE57x
VGS5YDX3gaDgYhUFRuBIDTgd3gVibXBW636TyOsisI6qx1n5VHUtAxk69A68pyKm0P26fUWCMmIH
g3ovqu8FwBIx6aGp70mhyxRiEtoTVuv0pCcqeLjATWkxt+fQfRdS+0tTkKRfgb0v7ab11kPohSyb
JY8A9LvG+gH2/CdakxQpsqd/r584xSuuIbzPBgmp9VBysr/oM60xVGifJwG+LnK+86hpedSzSCPL
vljHkKsfVHSQ1xrx8bdWuQl1Rj/N5k1WAm89Qi4J5s3TiP2PbdBKGNqjqNPp2luBF8uV5Osni40g
Ezirwgrhbc1HsNTRpMw9Exw77sBO2p+t4SjrK7Zyuy7srxg18fu6MpTQbcOMMbJyv5+Ai8j2DEtB
C6CVhBJRB/XD2ZEKJiwTavH1RXR7Kpb5P7aTXRzcaSXBBtRjxJ5dSIWpqIF7rr9GMlfPHXvpxT+n
DmIVG71AOZ9PC7ZkFVZ+vxfvpHHI7sLzfKURJFVpK0kUWbz+XMOmLGl1wcHzzOfBPYDEHYlCfgiF
8UnsMaY/gbctSwxtNc7LHtTpAFi9hdNtQ2KoG6jRVKF2eMECggX68vyDO/wezmPZijEMldADIUl5
/EGbgxZ77rr4IMY7qi4F1d0bVJivIHl/MhbcxoSFt9EovMAWewbQkbDu2rNdSVr5ojW+GkiuXhu+
Gf3eTnuqTbekox4Zf3TJVp1tYHBjvTxodCk83TOvrYxMPHT4L5mUjm42VjGuvc/2j7CBIIQjM9/U
oNYOexIyJZK57nUpOVw7W7ZMFLD7kHq2WPQhuRig3V2pT7L5Gb6uGkLPqrmquwyymoxMYmrq0Xyf
lyVfqnvgkh9zyjROzcc0zr0iArVN3w38Z6HZWw5lR4Lj5vkv3y07Y8uFeFsIMOkruvQwjKyh8VY7
SV3ItfTcOspq+9EcRWG24lagtjtNXL18I1atE83QjivJzJSzz2pUp3ePeKGp3VdhRr98a/gMOnym
mBxMyVkKVNJHRugFviMsRcqFkSX4uCSKdeKcQZ0l8Obma47l5qKAHnAkKQ2OugNHc/jwrMXKSHiY
Vx3zJfJZpT6oWYfmKJQM66YKsVZvC0LrHgXYMpn8QlQecVrEULKSqmy8+/fJd5EQlgi5fsVT2zXB
zWoga5FvaRqh5rxZ1deIhuzqcL0tARs3XTKUj4PRqj4a2Fy6ih7efHDQLBJxLK9Y+iFyjs6pU0DN
mhVqssHEJFClFDryRR993F+vACOeTBj++7yVKyupnP60cFm/TzqX++6MrxAkY+A6fBw2ONkLvei0
L73NVDOlmoQ3yaRSH1I3awCkiMQKEATYE1oeNCObkLIH8y24I3psl571Y9VuPgnZ6yb9+EweTiBu
7CyJJdnVVHmW3kOpKsbDOO8lBHsVc6y1+9AGosBPsiB3K5ptpZz4bd3FafaTrvovWBsBWLCNb5Ad
Dm967lt2XSZwmsIxtKLf38ZIvQwLA91APUGVddzX9LPNdSD9QGnLoK7F77UabBGmD6bb7JVa3bT+
BiRMPrgbsgvBN0QHhSP9uRpN7E9QnZ1nYTOzrjv1sTtq7L63swCtA8BveAe+LTdNd+zxYCxeSiG4
jTej9z25BCc/lNMzvgJ1uGtWsOFkxyzRR1uqyjP9xSg6NjTnIgntppepRudY3DXAIILB0J2qLmdH
ANdp7iKzlJpNDmAt9Adrd13sRgsLMYOgnu5L8Fpw8R6h1LQo8YN1pc4n8GH8iK63MMISF/T03bJK
B7umBnYxW9XcZBFSjjWeBx5sv06PHNpyNgWNyjv8wD6iztfrn06btDgmSibAXTDP9DsdQYOFkSxQ
T6bHRcjvtnhHZ5DSBFtl8to0YRA/+9lyqtgEUEL1FLP3IV8tWGz6toGlUaE++pu5amep/K20TZ+v
TmkjSAKY6GHRHgdQuSbf0kMn1kYaXxT7lNehjH+lTS6gMYXAq70X3rn6/g9+qlUPEsVNzyAtz+Zt
nyooVeYVoyhnLIZ1aAFJ/Xyk393D05yUeP38PYn9tmqWDrWTMddKgebvxfc43phBex5my7GHObEQ
egr/XoTWrTKOM5q0kGg//kFI52az0PmkdKe6460HtY3v4+CByWknYQrWHMnowyrubfXiDaPgit3e
LhBbvLfjlA/IZ+xT47ThDk/ZdN3HG2isPntugwRWT5tNc5UED4ZLN9wsB8t5fJf6Dzx5SELGPE1/
1kga5msVGfiqDWYwJ6AGe7XQ7xozAseSCOEjYT37SSrPXxpzA+9FJJ5eEz4KO9OEVBFB4AOTEcYH
Jy5KBRe9Pjbwoszewkf3XK5wtiju3Kh2x0qjdjFtOY/khig8Dujnz3+3C2hwy4jHWRIDcE4/FSPI
B8M93HnHnLJlMWMPWRyZpzIhUKqsnVVw8K4buNqlstXPpNv4Cic1YKN7T0esWO3VdyIDermm5KzG
9dTdKcML1mgnDrdokpYR2qbDxpbNSvStlr8DqDgv5YlLk5ULfeJF5ld7PY3rDgzkCzvAoa9Vf5lV
m2SowUWOxlMkvfZskCwuigKUcvfi+/EXCJwtjY+uSoaAF8jrtTJ7by0Ym3FBJKXxcOCiIU/TSnr7
KhClx2Eac0j54Q9YRWqSslRyWa89zAahhUUaSAgXX8ryV93mTucdbdttUeEUzPK12spdszQRc688
91GMFybtFizoZsTLdR7w4/OgfmV4aeihXe2S2B8mJf1oXT6lWQHMcjQGzB7oefukuNZdAS3CaZuH
pm6dmptmSo6GZ3P3pZQRXGpKgUlUUs2sKpPR6efKL+CreSmncP4FnSTEy9tQ/bGZbyGphIk67Cgr
pHspjymqEFOCkj64vA1kncwRNXd6iDk5MeTIbme5dXjFzO+xYo4SMhBFJMulPoUBTIoe2A/8sxbk
um7wZ1IO+CVVkK9TcQRSgR/n52Id/EHl+boRVN3VgrDKvnWv1ik/imASrcXhZqznpoio1SaDKcZn
IwwDhlRbetqv+n/jh7dg4aP+VgaKWSecWOcG97zKV40CqlzM8opOV1yJ7qEIrEXl8NgBg64ripF1
KyulTXXw3CSE/PgdMIANH42kniaDEEUcs+DwOlzT0dpqmBFNKIJHI5lwZletX/lIfQcp2fJjtxFb
F1GyyHcQraUMUAJEts7Tk+Gp1AshuoLgWFRTeZ+p5GZPeCDjHz98cyaaIYzHQ7djVevVeFEVtcAm
mu2h8V5bSXtkX5TrfInCMaI2RPLz+DXc3sUJ6lNEuhsDToLwK5TmQgQ5x+M3fQ1Fax4k27ty8aUb
/aEOd94I/tpuvY+JVijtnWbBOzkIbfaPsaLa7O0+s5Gq9YlU8E68TJA6ZBCwDuwmnSm61orb1Lzr
nwSeODWQZzpbqVpI36209fHZLaF/nr3shWroTnKp3MNNXNlRXnGfkmc1YV1kCl4eFz4F7J2EB1fE
d/tGKxC1RpnuVckPYWSxm39HhnbHlu2qp6IpTA8o3DAzl4C6n5wYFPWiW2CIPK6duziQEWLZX2sc
r//n1DZ0rlXgmMZNGcJN0TOpvSQptc9yd6YCJdAleqbSnxIcfcfV77QLA619VDyGnkPgTyZ9lnLp
vuszGDluoi8iMy6mK0Cy8RYk9SD9eZb7Sj9NGnGZpbtI1ifCujuXmgpfsCme9knF+m8/q5qIGKNY
ex6691ES08Bg1H7pcv++BusG5L8nHaSgSPhw9ZT9E2KM6tvMuwBuRcM1sfw0Z9AU2+D9Rgr4g3us
oByOuW8kdTkH7AccJhLEpgyQBQf0PNMjW+TaKeEQEGM95XDfSHVQvx9pdgCzUu+nftvs25Gw+Twj
G+BHufTJ74Rhn32YYoCEvMAVGe0gnUYtazeqiYKj/xbBDdray43Qj9OrAue1kdI85lCaYQJ6s14W
9o/YLRznVzjRjXH9HlUkMhdCjxmJewDchhHCmKczlP1nh9vQkEWZofXZKCuJGXYj0iZ/U2UAT+qo
LSJ1o+48U5rGlkCRt4+jpu/yWK04axnKuwtlHYaCCIrDj6sBAOmt8svC5bonfCV6JTpZdUuPRC+j
+rIVSXXAbDwJlqwzagFyJQqu8f/Pw/UZoF9Pyal36b0sV8izrivnwe1lWnwRF7epKIIwLv/0/iRJ
E7IGGdhyxIxVSThA/jA1skrCVJwk1fUWC4EIuifaxZGAJlUoWj7NQRm1kgdTnbO9ppv0VCX4IWRU
sserpVyGVNcmgzM7Qd281AsSO/ds3BMMW1AjVl0Khw11WUJ8xintN7cIcS4+t4K9iXYNKUdvbpja
DzcOzn0HZ6DnKwDQPqiJN4I4f1dsMw3xPLeRI2X6g1WrOkeo2jTOn+OhqHNobtHO3wWYpn4vfrch
ij3M0f5/PIc3A3ZCEfuqULszhawpN2kygNp0lJKLpTmvQQcAx1Mr8AzPYbBi76dSYqrfu6lA8U/n
zRuaoHW31lB6yxJNCnlcaAmLm2QE3Cpbjsp8/r2QyRIb6FhS4WzQAri+ry9Muk962TNW5p2v+ZEG
QlgLX4F+hwlEFyFXE26Zsl7hbAkTwAe5BDt/7RSsXP38zYFGqGx7qJJtT6ISd+Edo2eLZ9AmDyrR
bu7GxKVY2W9qtlD1uBsZ15FeZ83fdYMH+xeld6U0Ytrag6xgAYsLHuAuixqK0gfOPOwOuK5Oh2+U
AX8EXoQD6JEFahiJKmdPk+VwL01ZGs+WSecYAHhEhJY6qty1c1FZ2T27l9Agi0ag5GlqvTNmPXRD
mGWi054bJH2CKMCbnIknMGrQ85px0a70PTMPeOWje2JZ6ktBbaWzIzgVODl0azts3wbfVmLyd1eO
n0ANMfK8ppHx747wXUQDGCMq3adIQOWtUIF5tLQOkxJtjvF/9ekhdcxhSDi/uHvGmos83hwkuVI5
ug/gn0MXjPKR97ohPg8gMBc3TN05H8KFeaaFJWq98rRpAoiBXiR29CyEBwpN9LwSSUtVOaLkZtO0
daW5oP90VYRrs8Pt27I+qHerFk1NXqLckB2GAhG4uDm4soSh2nxEbtKfans4fjL0voCqK+pNKWiy
gVMHXS9jO7rphsQ0mZ7aTKe9p095nFst7Bqik1cswLBVWyN5K08/DkZQ2Nt3HLL7AkCmVE5UR0h5
+MR9qGh78yy2YXtiBANO3JCBPyiP0BPnzThc1WZJORhs0whEkKRpXidXMvZDlPwVRm0sC8TwiEcq
WQlT2WK5sdhol0fhlctb9kwojILd9KNH0MP2vQEbm+fryiQ3hO472csD74JLrGqlwVA/MnHqn/OC
ivDe7pvgbYo/KdWyAmuKhDNMD7U7CzStEwBdRaoWYtWwhHTcDoK50QRzpDyrKhpmFgZAhSkwz86+
lBqR01MEEKfiNUhfzx8mlL7zJUmurEOtLII7+E9eztRuswDye0Pa0/rOkKSgDK/tAZy0xAywoCFK
EqAOYDZTM8319zT6M+Ti+4WnH7KpRHemQtxTbvyFodgGPlO9sKmcOIS4k+H5zjlBUHbFHWeDnrL6
VN0cB5yUgU2KzuYWoZHOWwOJRYI4iCCkXDMIenfmd3uqq7iEEnX0JrIDNQrFAsT+0+yBG0WzQEPz
Fw1u9r8oGSTzcHOcA3qWsgUZpHTU/jiJywZXriMxPBDe3C8+YCWS6LxpuwO6ZmvjFDyZR6fP2xPw
ESUw7Km/UclfQvhpeP76m44tyleM+xmX2nyx7YATVCjBycsYD5dq5l+xrdAmnMlHMQieYj6A5uX+
8aazmxzlR5tJeN+VK2zS4Sp+wyCKsAsojnCsl6plE7HvbwxbZwoahNqD/OFXAO4VCMsuEJ3xIFZe
sC5Ww0ZkNdxzCebZdLy1Nxyhf8gVe94475PD/qcNet0tSw7ja6m+ZLJ+9UCQ91YQI5dQzq5IHqCV
W2AQF4+kHI66eEzBW/qiig/tXo1p0VOsnyUD1uaD5C4B3J1kcf/C3E5YoHSWLEJqsclyMNB1dW2R
kgCTH4Oj1c3/DjL0Q07KGYMZYaf+ohGy4FNzlyfGZ5pMH3UNH37Rtlk3LjZQq0WLAYiPiEmmi4mX
KMbco6yv+MT539beYbPKNZmP03iaukhQYAy7XTYVAzp4U29ypgl7v88Y9nRpWwHxCcSNBfuo5dea
BLwp7jo8iOyzEPQLxUr9yTfoTMAFIbqn/DDUharZCuYUnrkGcBdAXjFF6XI1sX3HTjgRKHgPkyQZ
yTzlZYOv63e6HllIKg3kvVaZ+SBtmdguT1gTdvLeKFH1TRriGhMBDRNTknxgTnnvzqonNXVoqeli
bYv0a1PM8L8aUDMGmzBW1s56KlT74SZe/9JjKbN2xG72/rTA8UmWMJ3li6X+su9vLNYJZxVFnA2Z
xmxjAZB1BMv8YGZx5JGyG3PPUG/KUc3r7qyf62IgGvlrPHJI01NJR3gvr3uyMR+AA4S+539Ly54K
syYAk2KEPNjYGbyTCNhetKP2gs1AnmA0j32ybIAZ5q3VxLLn8UhAgrY18WMzN93Djpb1/8sO5cIF
bbuZ5iwan0DvoT8IQ4K476cBh7VuqpyAAWt7NOlgEjgFTPDLGUDisXRavDiHGnmCQk33YhYEP69+
oH63fiQxaDe54EXIiMP1e7J0MOKenRNIce1Uaj/vU/ESQpX5cWJiohRyCF502fp1S3zqPVLEvthH
NwpcaOTqb2HnfgMAaTatM+rbLSAd04kM7I4a0CfQAI9HmDoSxVTXMOKFC9b/wbDv9TX1z6ngZnUM
FNIEXlt8wrQIiUDBTZqPC7rsyoyBiR1awqwMZnucOZphLHGXIq5dsEQ2McHWSYnEgtSWAABuET5+
CbUp0KnG561kRwgkAP/sZeU01CFlPs0YhEsOiQokSNi+ExA6Nm5Y5hgOT6dZcrSAulUqDHivJf99
rmoSWNGGaHXbqqL/blzUSxOVS06ti0iyx0sY8OVUBDbaZSaDhvulFWINuD4Iqc0CbGKUgpW9sea3
xoRDth5hudD2OAOVBwrrURZhpHAbmsiL7I2bvmnEsdBwjJzS3opALnTX9CdWGrLRUQpY6amQ5W+i
k2fes5w/ZtqygALnaV4ZHMTdHwrM071HKNFY34U4lolUELy+Hb726o5Spy5/tg1FYQhuYo4Qyl4u
EQNp2Tulbb7kr9mqMPwhLnRJnkIrpktJWZuvec+08eSLTsLcu8yCe/aaYEaCucPEgoisctZGosdF
VXboTBLrCY0bNIFBh6NoSWQGbGXd65LRia32XeUdzk/KKHe02kFUShnjxw84BhtBbcGCpQbI2Mo+
DkoPsAL5cxXuhfZDG6Mbt/SP1mD9YilMs3VmbinwRs9lBQtYvj7d8BRA/B2K5cPX7Q7jLbfTMhEz
j368aYiZbJIggILfZAnyFajVttRnwgOwrwk7Rqku2VSzBAsxEX1K/lTvJXUbCySTaeyR50I6Bfvg
FLpSFYuTHwAh7hW9cVx60NOcp3wK6P6qAMCGnbhK+3UtctZd8ViQtuwC3GFHfQ3ZxYkNBtDIrWyj
obCVLgc4uZvTE60peL8v3R7KBnEa3LzzKqTW/Ley9cVP9+S7uSXYQV3tkXlWds3SYWbomdzlnLM7
HFI6f+zWOjlyofp7GhxttVWBt3Q5hIP76UECMItCJdjbaq2zfzBXg0w+3RResuf8lysgUSkVJTPs
OrKU4Q48rNNrtETWEz8NvKxAklghKyP4/GZ7NHdQjhzmifVK6Wsy16h7Vtan7G2riqtjZmkrsIyM
gWJxd3YgdwwokkXZVArXDZbwQbCnL6jYDyDrDE+xFri/sPoBzWoNkLJULpwSzweMyVIka5ssXX4x
FvZNiDAfMl2K4VWL4A9GNI9qPq+jKxuS0j4dymoatSUgE/OvvXMIv4O3tpIM9Zp1McZp+w7ZzPuQ
LzJSuzMxdsX7gyns7LfGZ5g2puVHS9BMhDpvSJAmQ9LM+UDJvG2yrYAbnfoRs2shyRTXyG3Gt9B5
m3jj6kwdp2BKNT31zUOSsUqxIRWPyZIPsbJ5TcpCHGlgIEoeztIXIQ8WPYcQ1G3JCD5SVVwYlFYR
p+uPrKm44euJWoe1aayL435jWZ+I8olIvAzqxBvonCkyijwiJCRM8+3doD9c5dGlptRmBRQPOagx
EkdEKAEWKIV3HgTLx+sdTKga1LCVRI+y9yj52zzyqxu/wumFjF57oiORGIGsYEP1QwFtM2lVjWxH
JwWE/Dc3XXx84cSR8zGyt1WIauNntC/17Kxh0KYOg0e+OCtO6FeW+HeYe4BJTS1N2doDkqB8Fzeo
y/+OXq/1R8/PPL9HGG11HsiJYsg5HzV6KgqkARG9iQ8z6DH2mgzIqUP2yuhWMhtEI+ikxFt2zkD9
z8NkwlssgcQwzb818CbCF0a1FfPeosFwWgcgi27A44kd48SweXdlmta6vyED6lpMvqbuHxj+YdO4
ZZOG72zAT1kkZiPsHESG1QxFs37lqDzjR6zzEyftOAMMCuYcoOZO7+fbpEJp30pt8qEiz0Hh2Rk7
oNOutWtXey23ydOXkgWbPaz5VzgxV9ljm9O7GVvN9Eds9LQKGs9FWj6wXo6X1PEDYztSLEcinskV
RSmEL7CCUkGDFsOrjYxoS5QkvPdYUj3wDpY+cJeyvv0VCPjGt02ds9K2LwxleZVU4YmF2Ibb/e7h
H1RbSLgesIMbZ02axuMhEyuE3xUrN5r1zo2KLnA81YboCw1MnIOnQO/6YPS882P+43YThqAnjUSp
nWnY4xK4Bb9lffPKRZp18A9fuI9gWBrBTPy75gR74hUWYaB8ErFrkbzQnk3laz4EhkYGwrH7Z5Yj
s5HCWI9QlLBrHZkwE34A7hGIw92LR/9rIrQvkcsU8P1rlT1PEVUu85cZCl9dWIuYiQUMahaaybQ5
MlLvm1QmVrIVvo4S9G4wIjHr9MELBEH9qQPBsCgiVvjcZ0WWopkjeqrz8LpaSm5Bk7FHXKeXzlgD
NzNUuaMlifKDXJCY+n0G2YPaNJ9JHo1KQQ2BY1GrVVGfgzSSlhnB/GbaAqw5cqvhj0u7ldZAD8lO
5KnpL/dc9ZsrtvFvgrWT6jPHREDLKuW0DdW80Os9v63wm/2B0uBWokOH9CwXkf+Z6ei9e3CIh2iz
F51ehgOFdTEprnat65hp/D5EfT0uAn5pYgqF5jNIXtavEpvDV+Kw+yJHmOSOFIHvkgkQoLpmrN4N
K15XCGcgpBLSK+nbX76f9sBdGmhcIHcMSF1vuBP+ITotZlgYTGQ+kjMxIFWGM9t8h3e86zYHAnOT
6hyti5bPq80hUUUpt0VXBm23NJo7bt6XFai5IJiIsj9ITH3FVcaDxRjoAHGxBrpLQlvTaDYTiaG+
gX6JV0NX0jT8pzXwnszYK5osGDsMPrY5GrfkUpmX1LcRVHWkh4JG8ZLDnVMoXHM2T4hqjvSW/5Kg
nH91WbI98BcOKnXLMhP/SbhPvzldwGaLmytU/4NTlp8FIkENTzsn6wmKPvh0u+ibySyf2rxyFlmG
dTH0fdm20sYrpPkBCt86IW3zDr6w4lqa6/IJ9ftVPWE1xw35p76/wEfAbk08FQwNOkxICbZ5kKtm
WP+aabxyhTjVZueZ4wVcI5HJrmNtRWUkHT/jf4Upcofjk+T0vaUxkvR5TxgPGVtahMSq75J3XsGo
iYIS085m8RAThmcgH8/hbnsPF6VSNlbEFQ02LRZRZo8X5Fq9R21kth2GStoDIGchAyLsrm9ZRFNJ
LDLpK2I74JuWxxD870RMA+almwuLYTC8dLjrRZ38mfNdVTwf15BDBOZIx++qL6fJtoQozgM2q/dM
lEoJvH9oYF5WIPG23WX0RRok8Hw1Nj9je0Fz3kt+zsxITFOdlCo6bBj5mGjwS35EeW0FGx9RJBxT
r1BBKFJclIwvfDz3/z3F9eBu46knUVPMbSrJe32YaAdsubtcRWlpGSWC3tuc1xY/MmURdFON5cH8
URFp5Pk6hwgI5A9iEFa0cJpi/6EW4eUubujzecs2KYcxFwd+wQ/jBQualTbEP/BIqT3963ifhYBA
vUWsb2LBIVvDDCv/oRBcp4tdztiIsqRbkhxjAJRsgpPSHysalxMLI2CAq7vpUV9yK1EPC+3VJUCV
dGBbBhagdAbMQqveT2CwrRIe7KSRjsc3RdPvrNtOw8n2P8w89RZQjT5cD1EKdePkw+jgz4xpWq16
mF4eLvFdq7apvUx36SUz91SMv2+oAnh0rWkniUsgEna+Oc56QNytGbgKBIjp5dRPqwQQtPfeFWu7
NebyCN0SfnU2aN9DfsyTEZ9WPTq0Fh8vy3HLAOlehCGNG8Xh4CE+j3YzpQpZ08NOriA8esNwusmJ
Ti+Ihhw/pPucNISijpOTS7f0U0KxGeaUH88S8KcrnmwCnoED3USTkHc+C3elFjcf5bzMDJ1pAef4
zZZr8cY1epooZkg8LPveaTn8NBEaLlGYH/dhmhNY3R3kkBC2k4LxBunUxzRCk2jd5Gp045diQGt5
BmeCGBj7l1B6Hzmm45WITA3IG4+O4xj8Lv0ZuiE2keyk0yCOPT+CC4TXgKVbgqVVlW3y6/dhUJO1
sx71UEbP7HeMp5M4ui2QlFQj4ON3ME5IDXkKgGM20m5Jj7r7FnPvxe3te1LQ6XQnLry2npxovqR3
EYk3k2/kViZCqxrVsIZYFdbONZLyB1j5FwWJ69YapYe08ctEtSBSoDLZ7St3wvUZOyXKDL8WsAVq
6tG1VlwAza1OMhweZpHsUTkspLGf2OHaiLd5aNAJnOAGWhtDpV/tsIOP+Jjq743lQ3O82gHAXi7J
+Rdnlw6q/kpXKSTAO8YbxUnFGwI2zQ3of6jicStc0MHB9kcthsHBzrK6VJcMzoBEBrah1JGvz3dH
FEPEAQT/wAVf5gm2fCweAsvjmzqNOshRpJ50NPTCW5sq7GlLFvYwFVO8Q87mPDV9ZDJ/yhMRm/Zv
psOI+KDt0fguMVMLkC1xtTRgpC809yuPMVvH7fnsCA1WgTHZlJisFBQZdjBHRIJSKxO4YP3EdXYW
xE0QqeKLwca5KwI+NDJIa6AhrssLacFDFrDN0dThbGcUK/kQqSc0XtU7NXmj+j1HL7qTinsQkUFk
vt/CmStd5yPySEHSltzC2h/T8zsj95JuEzRNyQFReJeEJeMmsWHhy2XzRK2TXivP3AF9dWKsfTnC
Vxdf27lhpaCh03L969haPQERx/fqepK9KN/edbq9KEzPNmeuhYDMKn5/o2riatf7nMZWs6CnT8/j
WauYsQdtmZn/bAhsf+KuR0N0kOstwxLkdcYCrdNflJaAT8mQ4e0MAoHhOvDzMT6Yk7K1bRy5loxD
RAjN4XidQJ5WolwPbl+XNsAHuXM4DSwCY6UfqIjHmwRz8w9kEAfRLNXVK2vWY61zjwtVy+ENlqyg
Q4z83it3sojF8N8m01NjAdJakjIXGiJ8PD+IuPm7gmIyGEg0i1w0QSL03i2ive/AjFtJXNLmFcT+
9J4rfUVhuKSkviCeEt5KCrEAayHxnr0GljEnOtFHSTWGJssQEDX1r4aif8ur0kS8HzcdO2SdAKIg
n5zcBOMjf9IRZiRKgwNfD0X0ISCMH5Lsw+ATpJhMqesJiKe4eJkFCm/97Ln3ve6oVJocKR85JOcD
gN5ysKa5SmLb2/Z4O0Mhb+5+mm8yK7WpgB+C6KDeUgm9n8aV71jQSuQXLzZkIOXgz+slfJ269KZD
4LEF00lR7YGl49Dd5JqIxQMjawNoJfTX1NmTaIoe5Cy6IVXgkvZ1/dnvRovXpjmW+7szBqiPHaHh
E7mubI6Er7Q81wtkfo6reJjtTUZhn1ycubIq2rmafdjyl3+4/WOMe7Pt96cb2hJNgesGX2jaAkYS
jRwuDae37x1eUPrhphDVt+tRIGzm3xkFymobF00NQ8uyo29fAWMGhLajgu4iDj74zqawvjnzVQOl
vWo2tDFXqUbnGgXHKgKt9LXNGGxpcPVZC0/5K+NrUcFsv4InjguQqbduajHUNofLP0U5krAaVbNv
4rhAjDvWkGkkg6fKp4vvUkKLbgNeQ1reGOcHv3ejsuvk8FNPNL4E/dDStG7n+NEkDK0aS+9rghq3
jMfG1FnVOcnIBH90w6EE1sudA97m/cx+UIP8yFf0FZE6y6On9jekT0NLIqPFc3RiXuo7jG2BtzDR
URn4njfjW/bPmAQsrVZ2M/D9cNzm3DTUygpF/a2wwu69UDlu9oPEtTJKfcFMB1q3kCZAM7aDiL0U
eCNetyz75FUT1hOGuX+lcS6ij3s0sGmVjta7qiIyN/P4UVIrCUhE8xnsfzEDPRv+fF1LPctKNKMp
QsmfvxWct7xnfcskokwpj9bGAMZZi86chpxwiKz97mkjd4U+LHlVGoxMpiGl7vroqCq+U2Uzs7cf
j/9VMEVtqe+MaWYEuw9bUKRbPK6Fmx+TR8SjZ9K3piin4YEcDgb+J1DyyQC8LNLrZqkcMGnQG1Vb
sQnn48p9Cn7uPvHPWgIEebnFg8WpIvmovPfScqmQjBtoD1bFr0UNVmb8+kvB5447e/zcIc9KP0va
whoqmUgRu3nVJcvTAPuPqodL4EZzoO00OdGeEp6RyBfSaf7TprUJDTR8VxCmu9V8JhBolsksTNe5
eKUEcLeI0aPxkuWKL40VXBkrsrHvxOBDdj1XNbGRoJcaBTdI14f75J21K9vg3cc/Sc9yOS+WKd/+
sidAR/9ZR7ccnmUyC1txRdILyLAEqzHk2XSd4b5DToATNhoNRRz7zGx6lnOszGOe5qS9TmvkwzuB
mkHgPHazpPtNdEhJSHDvBQy3EyaSuWbQQ7chE/bOk5Ed2TK7bxuZcZL5CY30FVEYJdOvuQsAR+GO
0DEUGjz2SptO2emQzMncA6nmWc95HggCe+DmW4RqZDZZf6+jmMN7Gh8pnWx+6OPDQI5MsVjf+T7I
3EWRmCQWJsFoRaTjWRKxnS82K6rY2uSkbTCsn5NnV3L6+CVw/dDnFQ6C+fVjelO0GmG/4of8qU9N
vx3FVux12P+qa6oJjD+iGCSsHuqvxc/GOJpFcCIPguNAwp4eJZHcVYmbZD8IXM53FMizDnwxdZw2
X6gupa4Qut78XS37bimdm4Vg/8Ib5h+BrLTksVb7gzSbrBX5p5EwBdcd3WMT7t3z9uiLTuH55vPt
oSsK79kagz0qxz01drxlh3f/4t9jcY88UA0i9uAbg3ZDcfdpYIZhJzGcHvuXo/WX9uoD5EZAjMmu
SU5I2zahcVMxPpBCNQM/1OvCVUIu1klFn8JSdLAJ88muswfj874EeCyzP+uuF1LVgM43nu8yugrj
g/RBEYrSHZyrtQC0279vx9Mbr+URRi0KVFo6hjoPT8u99xLfaFUipz1acSYydEuCONUDwLNsqfqq
pnRrmDBLu7qjBL9dVhrkr0ywx20laN+3S72z5Eyy03ipv1WSkvsQ8VCyU38QskKABmuh7q/WxVE7
KvBklCUSVzLyWtXXapAZ++7l9P8g8SCoH3XGpRu96ETA7MErYL3kE5NOgDM6vGekLoAQezlOwkIH
4nbIB/TaDkvavnGoI1U73AxAodDJ3oepwiE2BRFs72JUWLKtUdWGYvA1gYECCOjLoT6e+om+tzTZ
Tkg9u7WKAH6A4rH56U0+2s1rpOOgk6NQE7wwOU+BrHGQe9nBy8KeEafkLHXGCcmIQ/1sLSNykQHT
dqv59onPNO8HCRZLb29eAYBcG7rMl7uENuXECR6GhuXaiSqDk1la+dXlWg0/mTQuNOp6pprFN5TU
8xCMc/NA7nQoFGZbteQ6ZQlWzaZtWBclnsQKTD3hQC6vyOMfivqOOsROLD5ZpDAwuZtfIv7787UX
qEOzNJN3oAJBPdzGVHHPwyAnss+kdIttFSzWcbETcgqFhkLnHLlv0RpO2bqwTfX3ERq7PfeWneqv
GXE8/3l+1ATBRVV1jsHyMkK104f+lHdmIQzyHMsbfzsiOuVbncZp81wKn4/zNX6Q+o0u/LDw3ntB
6l3Oe4y7S1BMPM/JLyxI2ZZQ4rzuLk8nCKCtZAvrZZQa4YH53vrTHu1FXvNKlik9c6f2CjF1JFwA
gVt/gUm3V9JY9ShPgQRhRDCo9WoIflFOzK004Ry8U7Sc5+GonEMEPT+KN3fkB6sDL2uw9msnyBES
s48dWrQQZsr3NAWtTbBhK7p4yKrTqQu2Tiq17kQUmNW8OpVTyGUgnbQS9lRW3GRDZ6kMJvw5KgaI
T3biGwKhIiFuyR3wDDcJbB4gKO8fR1ni8fD8QoCBjf4Hsv0ao+AWvz28mPNV7PnwMzSlTVxkN/Lt
T5k3WD8qw45sDe51mMk+YeVoC8WISdxlmQ769RjKfJAQWN85VitSqHMznIMiKjmgc9Wcbi2as7j/
Yfg1DYeoWwOFFLDr2LXMP7MxxJizY2Bu8dNi4VqCRpOimEBAv3xQ+5Z7d5awgODUM35XSVGoP1C9
yw9VZ7aOwHZbrqAsDjZrIy8P37TyJdZrt3k7/27Ad8iThhaHPYcLKL8gWBTtUUW+1mRiWiyIgjnF
1gdl1Iifa4QhnoEYok4hTDHAije2SNc/OuPGX8soBO9P1L5ZsB+ZKfjThE05rk04cP5mjYJnL5GU
01OOIaqKt8NJ430KcYvqoPeBk94WhW6O28YoZ+5iIPHTtztdRiUfteL8Hj6GBgT8JIZ8rmycyM8C
HXVQK+unGGLTI4XyCnoigYQcf0DAejfZYEgDPHVftFJzifboe/EeYkdenQVVEODf2+JxSV+maxMJ
qDpFX9p47caBC6ONLT0JgRdwbFD7mkX1mHPFMmsEZxXYcHFdE+nE32iypWGzrGPF8/wnI4WhakIB
vZ0TOFOXijrlax5TpWaL46JU7Rnxryl2ACXappaMd8ZzIi50VIxh7++yu7iGU/BNh39TkGMQjtcE
vVDI6JWP/EMgZra6yf1IRgHFqHJD+FoS+MQ4b7sp8L2/xrz/iJ9FW3ydmxKIgDEZQJVq8FExDTXa
ZcoVGd7DmSNGpqaW/8vmWrFHffCKC6B52hhzdToOf4bMy/co+NtDCCmSXH/SWOOhwhkU3p0AQ7+L
0Cb3VgFrx5BjmfIRqYsxUgx9MYWwgUiJ0cTWk7glXUM374676Xl33bY7cLZmifsnLZxOmkIUfr4O
yktpII2VS5aHujMHZ9sYDenpxZHETlei7WpX++8yP8XPZ3f3zAyjgVAVoXDmfvUhfFkaf7Bd31ww
Ht77uzNnVU7Kqqaqp9dp3XVONex2rmDyVHNsG4DhGTRinXq25/5huk6by31Mf4LBPeZ0m3OOj8bI
rA1ic60FpqjTMmQi1iuFBG0ngBWwzo+zd9SeHO72NNNJ5Pub/sMOUaOyO2AQb9pUgAgNlO6QjjER
dbCwcReSsYrWt+KWaROX9bCwtdY/SaCVjvZAS/GjWJb80Xt+4G1QtAmtt2oLZ2x2ckqB+GQw/SbM
wadCXgMvfHUMpA64rNleRPy/5FTozTI4OB2j8Ntjlk5XAWxwpOgIOrRD/uAP9XcCRxGIumWaj+F5
1Kob9QC8AwhIJ1v9bbfZix3+LgCHOS5wBcUYbpX9jMFmtAvw2vk+hmOqqI4hJr5Z0rzokyfKVZX9
Kwx3Fl0fsGhQY13xWzP33AeoGyaD3gBBzShHCnuw/MmHVAJT22nIl4URP2JlgeQ4/Ek7q1Tsnek+
yfjXlT9U0yd768TpSDwzTSUmE3L9za7QXEVN7ctCT2wTTOkPx3rU/hmktVc/9/QfmyBzz5vNtDpC
rWEjtc+H+Aysnl/vVnkYKlXGl42eM7B7M6l6hdnHrCWlLjPuKGchc+SiPJ5oNWCVFbZC8EAM6Q+d
oXB37K4Pzb6ToSqApYy3EzZHFVUAJAnm7h5efQS5Mi9yuZEufkBF4uHfgGQvrAN5LV5jERTZQLBX
xWzaONJ9MY9xkY0sf98B/FhjBktK4qxNjTXt/hBv+FWHQTL1fdNWew8mlOeCsfY4FOGtr2gD40tD
VKmkHe9oIbVoJV+MbNzVyXXnS1NxbNUvvProCQLcoL8fKaY7boT3uZD1RHRFKME+K3homJJfIzHu
TrCGZYhWRZqLpp8oVIC6gKQwVH0hbQtC2NdbA6TyBLXqdaqhDqWVJdvs9hZ57zp3mUojdsDv7s6O
Qo0a57nZNeiP7/ZVXD3aq0dKPvVST7CHgG2OrABpR5166NIO482ooT0I1CCG4jGPUNTWPlvwEXFc
DTrTPapA+b5zykYDIs4dfK+ZCSaLJoLagdslbsm5SPhJ8c7M0iaGVA+zJFCxdGrFhH8gB3Yaa3wB
QdOhsYjDDMO6WHFEbjoNhhVrj/TWIsHa3vKmp+uRYykMJ0nBaeaV64JZfKivUMIJ5J63G+QzImKO
YDxWg5xpKTO7+ajNeTcjU4v92Eg1ZAqCcYzfgL1QY9Ukn72haiNm1aFovbXoPaeYfDuYw4xcUEpB
V6E72hs+XKCI8Eh1Df97lhhpn/JXwHeOBWjP1F8FiP8/irQr9KHNe2UAZWOwsjV6TTfiIEKuLdaW
W8UmAHwO5B8QaCt1F+2MKZGDAwehIoOjCV8Ubu280mLWI5Tg0XZ97yw4EcFILdauwNKFvwmK+Rki
FnehSBBThD6e/5WCH40E3d1Dk32viRbCz7jStmlXCpX2xHrCwMXeyK5Gjh0x++vrgKR0NfJElbPF
npir+zzoYrJifig+ixzS+tLddMGn/MS9PxJNyQxbZIh5+kffkdbbDO9dcBZrSsjn4oJtsTrvGLDn
wpfpuVY2u/BIHA63JStmvDLwxNYALTakS5ApLq4zJRrdXAmfMPiijZzzNVCIL2NEcDv5kS/nOqmJ
3RHhKwltFFPwQiXq7iy7OygnAzT8op4XUPV+xruXLXpcNzw1W/YVMX6mknsgdJlU9nmZom4H+DEk
HDMYC/ZHXv50/NRwDMA5qfMmoP9hNarCG9G266x4zrBqbucEMIlwJaUfN6BE6dB8mi2yl0TnlAzZ
VMwngn/f7hrQGrT4kH8CTmceuBR5//jS5z3GkDnyifDaz8UUF1DQWvhHUodbpubd3iWhjXQQBntM
8C6rWE1s9AD7NG0TaDBKZl20wVn214iKSs0EsAuVoqEAN12HNkk5rQrUfQe+sTqFgrRFMwfw7FOp
j+xzx/SXXhCGsGq7O6P6w+gUyRDGyd1o+XXzHNikHztFWHshyWMZsNEvB0OuWasy/O00qaxaUNPb
wSafl+mUfCqPrwYj1328NErp/PZLesPyDbFyLowqw8d2JTv2njNe2qFe1Ql+nsVZkciMMWL+Wa+o
LIDn21vy1TgCYdQRY9YP9pPdbUu0gELKLoifrwIn5SGRDzcOoreE87N2FuzPDvQWu0VEldiYfNZi
s0hWolYEtruXxRf59M3rr7FDAVsjxnnrN5lqgpgHDVOFso+OquzHVtiyPJIeD4nM5VlOm+kh1YL1
qvv7QrwJPZK3uKJ7zgMhi1hYfJVsmteWHepdT1/g3Un2zTzET0dq/QSxDcCcQI5ZTtBkV5GUNqqr
8MybPHDxcQda5hphxlgHKOmn9uH8hcJhAYHxmpIZtClpMslwGeym2qty7s9QZ/AFaYVpK+jY0W3r
6gElSrbVZMd4u1iug4mewr/90J9aj/YTah9EE8Il4FlCPrbDfZpNqDZG+TQ75F1GDD5HmeRsuJG/
tsRG5OhWRzmGiftVY8kTCv5sBe8ncRY6BLQ7Ph9HFBDkqgLNKP8xWwyySl0all0kI7LzFpFGcSkh
81hcI7kHvANK3N73fdMe2bN0OE7uX7+EQg/HgWd8Gv1KSo9pm0/KWywfEpwD2FrrQO+kd54V/nYO
/jzwZlk6435JipYAgATsyxFMJzB9+czWaBrL/W6ie0nINhSfHd4/XYiToNC5E1FKJrMwq7tOwZgM
Dbii9/5OILabEkK4qDSpO4/9oVuWv7hbAH79Qx7Freip17ddmS/rMcEcbBdQeGyEQOjp7/V1dmaB
4sipqxWS3e0fcUNg5Zub1w/5JS/gudTS+Ornr6xYYk4Pw7TBno0MQfVJeZWsEshch9Xyvt9DL/E5
dsOgtZvS7MdzVcbG5BK0gvrED9fCR3g99YOXuCrFq8E13kGn1yAYPwMGAJ/6XNNnaA6l/cMM3Ah1
n57EqEzPOqhKU/k0anu0nPFmqe4W5UDR1A/3cnRS8OfBglOLKwcj7QSP3rycl4+4fGEXVLGnSC2G
Tk9DhBbyYAnCjvGc9XmB5LQyhYNaG43gRx+kJV53DvXxJe6g1nRVq9iEIM8r54CIaEfmsOIponsj
43zrObjJCIn8Q+Fnp0S40OOdHc13kXo8esZmPuF9SsFH8aVy4VDHzWpkDByprLwobHjRdJMv5MK0
ibLn8Ib/ljGhIThLEs6vtasWAbwEk5kNyM0OKIqxMEG3wUUGez97TC9QQJZ/rPhdXYx+StvzBh5s
AbF57MrGFAcF+BLHkYFMo/DuTW6N7PkeGgI1bLig9acsqbmDoe1cG5tW/pEx0n/OgnEfs8xgeY69
XK83qd8lykHfAsekaxp4Hmtkl730q0djvQfgHMsn020uwweatLPVqjA/7flilWyRRMgiBwpjaZ4m
sAQbGKMabbKRSQ8wX/Yxrsrqtl1A6/JkVqBfwFbqfAc5K8hGLZzq1bqpbdokSPU5Y8hOgiGdz994
qYZt2U+gECPl4lLlvyGWY/vcxX/cV5KYvv2fIZZT4o1Rh3Yvlgim0rAnOVSb79JG+hFU8hYctNka
4qvO4qpZ8/ampyx1VcOhm7DZzyt/6eYribqFqIFOZjteGtL0kAHEBPgODPUPpp7shHkD6eTrOZ6e
foTQqENWycvrDFC24BDl8ad/2B01H0QHNVonqbnxUDmTdqCg4mOywe0pZGdzcMSawW2MmCyKcra5
uywMYTWhK5PO1iA07MlEumhavTlbAqJEJAX6TE3/tX/3lMuh7d8TOSz/oBMq4IoI8mCnFcpBq0qw
mPo2ES6f11AUkg9SxQjhl/Iduu5Rb2m9rKPmq65NXovoym6od/fH/mbrc4T/qoXQS+oO/X9UiX5R
Nu6+cv8LLNR2JeAuo9cCBXWJmY5zjgp23HG8+u+KYjkk0nkcXYEVIsqbGkmh5z8aFAGatKos5Tes
DvMeL44yrB/aQR/U8ToRa2XQX7zP/y+bp/QJdxH8ZsgCn/cwJ7tse/WiWRfxkKP//BXjrHMbMqGC
SvhnrsNFaN9SNGz5r5ifP72YP6riieeOzVvKg38r1joAlB2vuViMz235ENJPJ0e56kX4p4zQO/dz
RO78/1YtAM7AzbHQd2QE/J0IDIKqOLk76nA6Uc+HVWFkN15j6bBhPrVuvKIYm5nezmAzUu2a3ETU
1cie3n3T+TucFc3AVJNwIbRNW+fQqq8q0WrUmMbR1fL6iPSI4VKb9RRrKW7Qu6uvldayh/EhFWTv
5iyvCED1TZ4VbCK1lCMYTmPyjscut+PGBxAd22oEvJSTUZ/kzTRg/0flpDKMo640a4Sla93LJCA7
4mQFhbO9AqqSf4xuBm5/j8XCMH0jcNgSs2sKSxVQtO3cwjmTtWKioowhBWBR5OFGINcetGnyFI2P
cf+wcmm+hozZpLlK5E7K0txbMutE1qKalZPM/MYY8DOdWfSUURQbpbyaRlQcp+FsobZfWpnBR2f5
ujntjk7+gzAR0N20KlkSqRkY7E71r/d9JtWAAjipvRc5KjzYGNjHReCpmI52rL2hQPzWHSsnubMn
DoicBdTQH1zPSDqVFj1MY/TztS0bZnwO5yCefnWy4olVGz+TY8yBf0VIHXcsmtgXrbM5JDQQONJP
NucjTRTB96IcKoYyb0u7EKHmSz9XbR3ggD04YRAJxsD19OnE5gJBrcYFThPdTDg8ZrWpAqV6J3eR
g2ywhaVtvkHzLOPxUhY7o6a9u3igzs+emX4XvRUx6CwSQTriudeo/DVGCCWHLAi5NdEMu2dAd3JH
alDH1c96unrNnq7s5YRXLVx6Y6XVlxF3T5RSGpxq7SaNf9ygk2wDOOfSoqlWkNhumXtIjqBrLf1c
2NVvSv8VG3NTNzoIEIg9XQqvbzpwRNKGjomO7e6R2/eYGbSulcSMvVFWd69f+4XpxVpv6j39HgLB
T+4gFJzZtKDDv/Jb+zNIlAdvv72YdAyD9Ec2giP2QKZI4qTnYvjBFdA/f8pI7jJ3PKoQ2Qp94UCV
Ldon5i7jlUtE4wgBrJMLCcHi3HzLQIEIQYvVTz7fYpGcBrhrCy79USM1V7WCKD36esWsUwB72pR6
988VX5x0gz0NOCDRJ+S2Y7ueGZHedVvC8AmpnlrW8u0hyuwzw2dEMzNKQ3esPHsfhh+jjgIKfbS1
/Ei8vA4zfKLeichDYxChEZ8/GRzlmpOI25Oft3iI4YD8OYOREWFyf2/MGXZBPVg+8TGC8Pl6Ccem
2BfAk9HFhS4vutzSeHfVJu95amD2eCpowc46vizAxNANZkccGm5l4Mh1mnXolrMZhOQBVZhLhaM3
NeJSD6mgM9AOAxB/CflcKWb2x5vakrZ3rgXcK4RW/YUuHxwwH1ivYIVxahn1B2f751DY7DLfQaMO
ZVWVn/O8n59/yeoCnTatsDF/2+v2cy8RZAS9AZA1DL7DiE/xtDqBX4Ej2LWMA4h7/6fmLT0RBx93
gOS8j1vawZuWXpt7+KodCdkT3eOZP8piYUU0SoVHIJYSRa3SwTkSKU5RB3ez2jlE8+ICNRTIE1r9
mA5kWVL210E/zVlCUThTZPuEvYVVE/gz1Ib7Tr7b9F9t8StaUY3onaVQQG1jvaogeTaUfHgtPtfu
tifiJWbnF9QH1xPlZeJjpieSK93KCR9f7M3oGupTMLydfh6t6XGZovTO5mZlRaGsgOe+KyD3MnQS
LtjI+iHnCW0R4APzrzQ+SECTQGD+aj3OzAwXkqkQl9zpjVXTrhdSQZlnXrIn2aZjgEgsEjlpw8AV
nrRR0Ua3VSJbw1dnb4/96sSu/3hR5vA9rmtzMcQV1AgEnGVlq1tovIySBZqRNNy0JkvpqpucYz0e
GN1R8A8X4rIGTAr/7/DwAOqVRAfDRqoxk3056bh72tOrEMGCG6lHbt145dCMm/5TzEq9dxDNuvf+
291ZqD7OvYLUi3Ih1OcOLBi91afhS5suvoSdmHn9rkPmS/2xxxAfr0ynp+9Cvzv6rjcql36T2v2M
Dp3s2l2DD4jA7dfg3oNmNGsBnzGcA7E5lSKUNCefS9FqkmpTF+KB2pYqy/XU1l/M1FcH/fhdLhBl
qrScqJiZm5xEQWD6BdxNgJO2SEYFCmiweRada44Wi6nckW23iWzodd2rAHcPmsdEVLvXHnuKVoNj
68pTgjwnyUp7zT3sb+MhfePEo9a11ouo5ylJWs9E9nSMevF8ceUj+918X1B65ee4L8DxDc0kOyFn
rvS4Gi3AbuIMk8yBlhiNSPk2fyaHrNjDcyqIjqfNjNAg07r01NQc0hMCYUNNT8M2oI6+yNM68oiI
uIh+tX8FDVklkgE7lSmtmoPTBgYxYyCeVTzUb36j+5NbftNgfDJUXHXxi5owKP2X+naHYOd1ol2O
WwEKqyUDylxsTGaZFXnSaPHppv0R+KqhIr6hQk17xE8TBNxl28OcvP8hyURcldR1gApjdol3odXc
MgxT3L4MERca14AYODJgXfxDgJUpisIMmJuCWLddqzuT/brzZ4Dp02KYEHjRZQoEpl6yPwi63c1L
TbrGZaRjksYY1+ZG/ZXLx/zdHWjwZfJXVYjCLGKD81JlwmUErSDK+xziHJ6Z1o6DuNqMETsRY4UL
9UHR/i5IpIAh5igf/bR1CNyWmgfnvKJBN5KGguU2Gb6L9zHDsghX2lrnsH7qp6y9vj9rxiXLYZfx
Hs7pF2m6ztHaVWwfeBaM45QOJ9x7iGJkiW+l7SshFkM+5J36bF6y2L382oM8aBa2umAVcwP3PyII
Df0tbqRIgfQuWTcw85W8+E3sgXcSK/X34/DcslDLT5hwaIFsdMYA7X+kYPRx+GdO5CMKC2CRwD/u
+f/aAcD4Zkgn2hfPTRoIc3x6+y/+VmcJUjddBSbxTJ86WXmjcrqDq0/ARvcsWNc5mpZpT+4bT94L
cpzNM5xtP4S/+OLWUNy58G0h40PxWoMee0C6ThrVeDCPd11pfMoD9Jd0c1yL/UC+Q4VyDpPphl4e
s1lhEUf5Uy6aE5b8bDUNPipmMuOPefpeTRd5y/53mcD6uWkY67OR99FOeGX+NcQ8j7aW1h8XcaX0
fNeQggJI9dzVPpI+rZcQyEsZPIzbC8GKMOqfv69pzm2dIIbh45xkqZki+vIBYMUGsU8uynQKicrJ
qTUpItEpOZ9BRYIweYrSoTh8M1dgdmKINgcVLkIwG4rGINTZh93eWCv/Q4VRiHzW4tAfoahDpRaC
fMU/65N48kq516hHuq4Zkid70QF75RHeeH0DPdsjK0K3PrvATtVAtNbWQwsAh2nMuWeGD9uv1mcK
WFCFlPQguUxzPWf6XbiWPi9lpmxjwZFsz0Yd3heNFeVAY4n+TfYVarj/gsCRoZYKoKnTv4KqUIVU
++gRea+BUXeaAJyOQ2uZL2Abtvzo3t/HOsP9HKH1ACpKCB8RqCtwHxZTXiq1X4zaobG0SdPyC8kN
jBo2UQ5V8zv3SADMf11SdYITQHnsw5VaHUwtMNg6NyjArsSDUW1Q3M9HP30LOhQUSQNRnBcgo+wq
GKuz/pETy8NxXq1iE+kucAFpWgbZ9ZP6AAz7TyfyDRJtLmNfjZk2TXxneu8iKt18yKm/On84WI9m
MVDtJPN93v9ZzzP4aMi2izRCZXchN6KT7rHFdJD57ldiAzNnUmgp756jNRnOobNt/nhY2IRgrIr+
l+cKtmg3H+d/V8iRF+YabHBUwhH0arwottZHj2HXh3pQQ4Z05D3VDzj2NMgwI7aq6dIl+9agYyAV
E2POTD8kwGW/sJvkkc6zHOgGjcEPCY1J8ds1vdPC/7TeFqpySRqDjvDVLR96GZxAKOisrb9FX+Wy
B868MYBaps+jUdSY9mO1XwKScmL020wC6+0WWtA3gJc5pXWcSRGrQaQqPNAZ46K1p5ZiNjJzDhG7
UGOzTqBU+KHkq4UmUPIubDBiPnPnVawJvfdxOzrpYpfVVrDc+2ReYKr9wODi1eWkmLTP8A+/2B25
3c4ONKdRlnPHvfSNHzyjVVz0QxK0JgQFtLTe1OABHdjdcm7mNrctfYNqQk4q/P0Ybvgu/DQZRjG6
rIEROM1dkC23npAgxv1LtjxvZs4VMK2Kt64nsSY6iVG5uVQ4Pps09cETPruz+Myx68u3bRal+YsL
7RcQZi5SYuXabXsLQEe9qbj9Wnjz5RcC6AFkaLr5nGbcz0dXjEkYZOexOkb4n+uQaIXOVGSiTVm1
uXDkwTysuKcCfK9Tkk3R94KObLPQyVcE/wx5Xfho/mxycTj0kiYy/1UKyjmrfAmZNX1fA4kDwLif
PJbFZbNsmIlWfnYa/cXJRNcP3pX4sqeHMnU5HQZzLB3IUP47vexbkVzDmhw9Uji3ekGHYzUkLumC
0xgerwloTsfQFwwl6/K76EIAV5O1NC6gdh3JgU9mZ4M4nmaV3IQdEJVaguOY2/gkBuN8HznXkIna
Ku7UuCnIEc8Y0fsHIfGZGfnecXJrMlaGy1Re2c+4fs3+f+wz6HxplAJVWyOlCwkx+5nz/2Kt5j6r
ndGbiRvTb7p/4ROuGP/x3kzcjNv0Cme+zhkUKjbYMvzfzW/p2PMwFEBr0ON1YWUKBMhEJytpbg49
mF9mqcY/xROTRPxK0qYn/edmM7T6iChJL0K24y+Z3C/4kemHbvCitQsXeeY40ke4ILgRQtdoxBqI
S0W9NUvFMTcZCki8hmK/eciFqZl7c7oXnQNPNa2RS2G1xQ5jGLsOG00kbiU25sZVOGtXpJCO8flO
FGHKArXzJ7/soIwGD0j7+BaDyQDepUDrAheS3baTJOqwTj+Szq8tiyszm4JVY7PxQyGJy4J2wEQP
A+Ime2lln0pcQCeSlRUyw0U7uY3yxwLUPNdSOWvq+e7T6cdoDnWKLach78ddmwJT67kvDVImbWKC
5PKx0rDvcZ/gzIwuDrJEsr+22gIrBVVDXD5bL/WjZgnSJrcKXo20QIARE3xYeMF8i3xzrzEtr7Yi
yeGqg529JWAkUzPA+wlTdVReMai2mvn38+y3J5gFyA/FujiMGqGqlzna3NFSlIORVFxZZCPZymYQ
pNYuxpmOo0/DZJvCOrX8Ir8OJZwca0Kg4CVjS91GZHUj6gu3EPHyiYK+iKyI/ieyYntwTKm10dO9
rFII5x9lD4BOae1Midh7mTSq1Cpb8sLQk5WS3dY7IviiNDNVEeEN8+7tIyuW5a3dQ6ZkgH+M0JhZ
LCfOc4Q+2ig0TXKcrLMwMFX11gMv9ZcVqbDdpCWj1HDCp9ohBg/wa6tTqe7sEr87sNmgCIQ9Jyeu
PZuJDbpCcUNK9fB9AJ1+DG1ZIQZCIehajsraz6aY1slwWRSiMX/d8DeleDZUDJpLOR0P6Lx9Aauf
i+uj4ruM8g4sE8SG9Ym6AKc71EtOCCHryLt7v6PSZ0aQhNYlSJhHECsfgj/h87BKOKGw/3u4MArU
LeHe+Tw6B97PAS4nji8sbqvB5K7Rjds9davRhzfTvcB9X+JDzPrA6zUObcaCz/icwscqv4DNP1nE
WOXf71ZbnY+QQBY1xeVMsnERPuNooj1tGJJsWX03lCoq2V123CbqDfvqIy3pl2wPyA+m5JK4xUOm
fmXlp2Kd7eNdFNk2lmhF5gHoD/BUmJeot55e1oeZe0U1EbcASuzSEqcHViuDzNk4YfOyzfx49zNA
hTn0o4dq7Hump3Yy1GuVyUfskJSxRxS4OyKwbW0opc7js8WnKOQ1hrVAGvuwC6dQ4/WjnXjb2v8w
eRqLCKAChAqrg4cc4xWU2pfCLpK8vpsADLbY5TLm+1co0CDRfw+4zErhEqiN+i1cjnxbuUFaSTI2
iGC+ndGAs4APx9++0FjBm1lRuRPgI/5VPkx62dSTQwVocnXoZa5UlOTfFTFEBN5k2Ddn35K3cPVk
5Vd0vXUTJnRnQetRmqUjMFaM1Gx5TXElOZhNxAAWP6U9kzqbEzPC0ePOFxzI3MdqE6OhdPYA7AvV
VwCYmNAlqflWIyWMszTD2Fi/bt9eEzmzKX9k0VV0bfUgb0ahdXiRIOrO6MkiB/uYaZ0mGJf4OU8F
lOcwwGU/1QMU5kWA2h7PmvyODkolYWDBvd99gz0HA1yLBF5HBbDyfDjO4l23VI/IqoQ7Ey4xjbRf
bM4IQL1c/AIrA/fSU3+fjdYwHFDGxNoNDOYWgQdkEOwAzF5FT9nrx0trdMXUWnYnGvjWS83uZ4VH
x0g+NNYe4zq9Y2TEhs7Zw3dL/OWz6vzEhpo366E7qyZja9zDGrywcbpsp3z4F2eLDUCzoOvTJ9r5
ZYxFYU1WTBZOQRRWx5jcnARXaB/X1D2lnoh3LjwflZalXrW22dqYM9wWFpgTMCWtfClbLtBWscv5
+pvGstLgJ6ZeRC9CO8X0+Pa9j9Y7xjl4Te9JGynXRFfOKyJ09WMEOBO4FgB419oKNXe4h4MfdXyo
8PP0xU2vBbG5BB6efwdaNTCW1UvKk4kv1QhBrRk6rxr8U7xB3tK3dCUtEtKLze3ud82cgI4piaNi
btY3rxVNf621so+SlT4zYsj05UAifoFZnPEauuzGAGWlzXxAmTHEe/Xny7ygbPmz0LwRdRQAT1R5
wyH1uTkRHXq8lF5LvpNH1RtTknY9sDyS+iawSb3GqbW+MFYeN/K2UjqOnYx9T9VlEVaDMLuFxohQ
FZeVi7T1pD9X1vfVqtOHTQXDwxoCZcXxHHHzpqniJ7lbrCm+p1YgjaxkaVrpNFAt8cIPWsooL0C4
qOEFLdmVtlVWaoRmX0S0pmxkqXleACbP+q8GxZbjrYU1QconfRnOFKpFuNQ/HuI7INSkNgEZgW86
V+newObmntkW2BPtUyfp19Klr3F9jOg1oJqpTdpbken2sUDkQ5/YtSEheuJAQ2gd/XK/rrN7BCHA
+f7PJtbQ4ELdwI/udObnoNw3CtdDu97RV0Y0KaFM2mESaSP2N41DIshjMfTPb0bGEWX5+BB3xP7S
QmGMw+UzbeJrHqIZCA7g9wqkHEPOXjKt4OLNrgLQe1bTadh0grEL8Y3qrfA3/XNrPtBeQOrKmcUI
12D5GFjv3DiRSCgYhb2Fu0tk0Xj20l8IvBT9eBnLS8Tgmdm1r9hAdIOhYMYM9dIsYraXfCnnarlm
Rb2bZ/oFAavRSypHbYXOaqStDCA0A26CtLpJoGPgtJDsaqYBkfGdaICZe/PngxK18CHJDxFp7slC
+mdhR8VZYgNVr4KvV+NC/n0oPMlXyzCmgknJiyHNyWmcv2O74Vw+vm77sWYXqiTDa8v/SupqMt1V
/i64jYRKwx4oFiwRtV7nC8sMER8de+A039TbNu5IkjjTsMvRe5VpJMpXyUhTjT0vz3zl5jzg62pt
7vdk5kIRRR2Ssf3d8g1x3Y21GvPnFtVnwB/AU1tq+79wk+pKdE6vvYt01iHtJpZJN1vEsAWRNqC/
qsP231W1PbOyhTUJNlvaNPafxAgtBYF03eFjFv/cLIE/WM7NNyhDS80iwtOrIRoXMNrds4N+ulCr
IM4pGeGyFez0K/YUMEj0uiCNs/jF9ZB0Wl+dgpTOf9DENghzk4hEdWQkEiPFr79hJhURX0+gZ/xn
rphhk2MVGXbq3eNCMyN5K46yWa1C/CRugMRSLkLng+DWCpPLBL2h0GCZdSJkxQlrSuSFn3NlGGk3
kn/2SAr4PUMjjV+qxmOJrnVbtr/p/gSzSD7Tzqs4XunZ54xKzrc6PWPZsTA2ppwxDytOrOwo8CNE
R0XmbuIXAPYo98a5oABAGYcyJI8+1PZUDplXP4esKOPel5uUahNccVFWp+zkaZyEXGWeiY9z7W0a
GJAmdQDBOBZXN8azP4vggi3fWTbcacDnUmb6MKi6TeYctk28chXqJ9dF3lVe6mtXXyyBWZq+9e7L
Tt5o/KwLnWlHaY9dtU1tNo+rqflPps9biwuBgEc3sop3mlcJ2pnoSmG9gwx/O23iBVdOJXXh5u1z
d8xRY/oIkBTGeoN7dOB8ttF67meGt2kSR1AIH4KQRqozfeyGbsOFNe+eDb9DAtZ+4IVWqxGICXAS
+6zF0X92aDl44btcPJrrMaccKLzhWXL+iC/8Dy/L/etLxcIEj5aYgvsdF31G1SY5/4sGsxEsWmKB
L0CJuZEDUiqDa0wemH1AVrFEmc2Llr+vplyw0LzjUxKs5HSfZTds7g+grEh/zGbwDsc1rW/c/+LR
KS8mwDHraCQx1d2oy91l0OfbHoBxmPCnuENgHxA19vEUNRdWYVjGLEB3L44V3kWYtjMLMd0WJJmA
j+MLeRN2DPp4d5VvPxKKj+qUSkZbLONNtpuZ5Mj/HBwV+R1WOC0AX/m4qEwQQd0zzgN7cJoy7Rk7
dljOwGGTjL3M2kVBPN2/xUXURvLX9qSqTT8eodFbK8gr5Sdby9QT3lnUsgeNL+IqTSv5sPS6xaP/
KMv9h6gyHwscEbXLzn2cJFMeRQGoZnFcVc2+iTBPiJ8DJNwEH1OyHCETe8koMUbNJHV3giN+K3uN
JfjqDvGDen64wsvhKlWzz033BuDiphwmlCf8DXb38OWEQDjBPEShqOpfjHZ/cs21yGMNujt/UnFk
tzEPjX0weeXoxuLBV00ng6i5HvQG/0Pxf2HNhQi4Mdz+fTcaWaJj93clDNBU0P1k3VoB4ou0PG1H
S6kQZu/3Lwdlxqi+9NyWQm9wwIbXJLBEq/FrYGs8hLFYgSQgJdXXzGyb/kARZ/Z97+M9l8OXlwvi
2lZ7UmAc2oJkp9llbxD0Od69ht413i9Tt9m7zXr3YvOXUZjaGb4EDh11IFET1bGjp7M0l3CaUYfF
ny3ZipsZNEShoq5obVkaa6TPdeTYDhDI9laABE5nhNajrdes1KENAhZ9d54b2ODcLlFOj4cLYGNa
odmDdCNmBfL9KeawC1lVmTa6VqFLy90TWZn0zUzA3txch59HLN31rEQF2CmMa0QlhpwSbx/1hP37
EyodIBdeD3MTfGjj6rvDropyjpxhQDXaxdSeOnVFFWySVFw/YcLOi7HA5rdL3Wzqyh6h9bakk1Py
dWyYilfX9KciBStXXKKnWpE+Sezrx6+YJ3p9hopu6laeYRtJGcsnqL/h9pXoF7Q+16az2xd5ljRN
+lBllsGxino0SOD7j07r5HxK+VAgLZFlxKTsbR5W4WsijVVulbybdBL7CSAewxEzlyXgfmN+G+Ve
ydbIqWQH92Yzv2KJyZyhib8BB4Peo+Ki3Xk0VWaFHVRzt6bsqDoHF78FVvrXOb5TC6uBEQvt+k82
62BdJJ5Rn6a4ZFQ4REW2qo2BombIBr4DkcND8dCX/Xn0BG3FMaey0jV4VVfDg/KIZ33T7hj6O3oN
cdDx/BQL6XcfJGbJu0Qr8mNISIN/myqj+RZCi8h0kUOLcnhbZzdT/ZlAWHKB+6vuIdjzAD9UWw8E
V6sB+IZosXPljJEL43X9nuzpoU3oAYyVMp4vp+cxC6A3mzBm4QB7v8k979KGKOyvSvUcFExNx2tR
Cl+1WmOcY+kh2f+M+VLVYhkDqzV2hPIxqokdd0EGJJ4mFoSHhtDwx5u6mkWRKF/3XvD8SCmYB3b6
6szdnPIEhwKalmd5JNksv28kwg9VtLz+33nEQ5iyGi1KPv6zk5GrDA6KM+K68gPIeSeQm8imapvy
+fGerrJPwwdcj0+yPs5mQoH56QzHIXbwDN+VVinRJ7chA9aOqyBiB+WoO/EaKLLVVKBBUAnDFYSo
sv9nGXPvUvYoc7zeQiD+OD9Ua/q67SMFghvQf5TGRGuTHcopJB2NNMQIREM9dLjPr5NiBXULaDsV
D4bbQqpxLM4oVv/SIi3t7a7ihznqr2lclOUjrh0F1jlgzh+xQ4R6lFPbsVlbVJvnvkzZPgU4aFvd
g4rFd0OwrejjQAsOC5KXDFsawWfQeuBKJflSCONvkM+4C8W/NnHqc4Oa1ClIxYIlmKKb+egAN71c
b7frojDBv+OAI3alX7b1wLPhD67fH6IIsDpbyCEK0DBlUNrwlZnkkyQVvNiERrKx1qZkgBAQr8RG
LAUy6D5k/gLOJCZPzbK16mK4dVQw0/JUFj+vvUdb96ONWNhNELMguGsFDnA+BWTMbjGZRTJ9SCQB
5STghUmXrCgxpxoplAuYOjLV61XAXkIeb098ECIMzwmwoL0os2B8NdGZ9muhmDE1B8BA/UcBhH2t
sudI8gUMVj1BoIKwvLGoNWMjxnl+Ouj5ofH+9zJ220ic+Xt4nbvaCjhvzNXCmhPHjZ0ryTe3NZFw
iJ5/cFE97lHdVBiOUJBfsKHeYubAYOHmX2mNDZ8PXPd1uofPVPWJ5V7/FU/wTW2WbCDsW/Ofq8dl
aCqa472WW+G567Y9jUUGwyJ5IeWzZmR3GZUK64usk1VDyFcVxqXrG4TlVPesDylKRI7v4tnItKBV
H55yO2AI3un4qd7xIMUP7/YS/2BA5B+o5R/D+R/Hz4uuZKOWX3OCcU1NtvgBh61ylXJNARbsKF0r
croLmNc1oAmorAihZLLeFh7KRj+pn5ZYZPfuczJSIblm3iCDwnvV1UBNrCYhaJ2dNSFAjd4emQx1
tXcid20UoQyCmtDB66LRjfUY4gxdSa4QHH9onBgkLLOQE6kQ4gOZ/uxVmQQHr9vlalfyZPnTxprh
Non/EvOu7QC0TqUjYtR5tgLwOK0svEfvXWJfIbuDHN1AAj+NR1LtnJrTZRb10U4wB0Alvm//xGcI
nRuC2hwPFZRbcBPkO6h5uu0wSrIkLFxUSaufkmbGbPWsed3w4CmxuW46B+K61LbaGIsKYYoZHGPg
hvhJuiGQozjIzyjDGCENm/oR0d5rU3W0MdvMan2hLktjc0qs6vSCZkjpsYbRllL5P+churLqXkOt
Cmg+pAgN98fr2BnUDQXtc/ZuUfNJ0Yf7jb4FNVTiuutQgUSFd7AenalYFZPHIvBqrWuaoAIZo7Gl
7IcAVEwi4Epdww2CEOarV514pD6vlcUNalBqE5K7+G7zpT2tX4SY6PdAJkXM4+FmJw6+meXyloSf
LqSYxd3TrFvDmkzTZn5Q+zCcAr8NxK7ngXiw9kApZgE8XtdPx95puRY7AovRD1VWkUewo9Fe+olb
GqpiOXjVihhQhBvVghGk8pb1SMM7HaiCJDAaHWAFetclsMfATCG5tuGDm4AhyoANG/T0ZzYAjxjF
kyRuPaXSDfHC0fBFYtRR6CU5/7/xd+JP8m0mZz6dTnWYdJG7786qecQI7GLjgCFC20Li57PY7Cci
bKaj/3uXtvn9Pz8eBinauDw8q3YiaA+vuAb1eyRybN/1J3uZAl4ZnGpWf4ywWa7gmqS1zacVpxyq
Zzq8JplQIv0SKM0AA6XBkb3ihYDbZuMys2quz7tcuW6sivNUhVeTvzkBPmI084P9+dfQKTUT5AZi
IhjWdGVePSK9rPsRvTRywcjb1dVw1tSK2JorHMUk59P30z/bh5BAuqbC3P516SNtcrpxcp/Hct6x
snuH3FnXKHd5Ft6kxvifRdcNAKFTP+lrTTYRd8c5oLtzdL1SfmV1kkVi/5i0wOEmgZ9p223Kww76
SvQREgIWa4i2A9A8ObiwzUZPIlbqmqH9+gUY//0C7+oIVBt9FjczIGGDAbUzh5NSl3uMUW1ljek9
fyuzWamhSLINVlTXjxXq+mthAcn3Vn+k6tWbSXTbIHzuRMyJCdzpLj5gu1pj5by3QWYxx4prbDPD
tm3oS/1vLpkz6n4WIXIkbGRnTdv7E0HoKApAcy61mIqB4sL7BFvXsOSKlzn/ywpM1muo9DOjrLA5
oOpRwy8K1GElUeS0v8MrJguxC3vuxLhzs8FLBMKevtpXnEvf6Neejr8Iza8MxLECWmh7r/NY1xWW
ZKROhIKVOi0Hi7fttViRJUTYRqGKeDOJichKn5vn3P/LxEdixRA/qhTCYSL2tb/IKSsJIofmV9UR
tjbMBlCReLUWpu0Knh27y9UaxzTPGtJzt6FqvwvBX5ua4+neeOybxnQCzvxTI8Z/1SAL/o4ZycM5
ZTzDJpcr0CYCYmPYgurPIAIkK3Xa3rfm4gmj8gRiUxaMR07XZROCBlJraOibV0A9lJrBLw7HskC5
6MlpY/h2O4JlanwPx3llBVBJYOhrD4+VVjZcdlha8by7RYSvCHWji+BID5bL/oopv3hnsAg02wBM
J/ybF8ApUGmOaE8IaCE3P/27X36JBdFEPY16M2ox7h1UZfKRQD20JfKGcX2//7wnjIKYH+mt843a
Cb7jL1n1Zj7IuKGe6Db4D/V2gvv5O/wsNdDc9VVJQB5qgCFNDC+YRuH3Lwc1StdWXoRUtm6QcUsc
GdmxYHFLjpC3oUaRSkCLngOWMeOcw5V2acDCh75vtKXdkUiLwbqkI22QpjNujBxzcnSG9NTkBzQC
epT/ADezXfVet0xwsl4sSQncT1r3GWSy0EFnw9+xYsW0kujzbbCBC0eWL73Ada0pwXjxxTznWpmN
wDsUzb8/WLMW9QxsNMs2kxma6M7Yd+LxMWupDdxrLOMUN64CPmu44NB7PlZ+wYgVrTlHdBHIfG1a
gPrdFKgeRilUNpkD0sv5FRHif/AhY8j7rwcAlD8kXEyklIvOPL2+WKnjegBmk0vLK6Cw/aF7shk1
IrQPMRIbR+5SzGl+fptHCYW96oST2bOGAprL5xSFhOFCe5CLygiLWq5IgkbDEEZJO4qhLyp4O25/
tvNOtBcsxRbLSZ4aZM5q7bfM7moLGgJ2DbFMaX6Tz9mvEnF6sUyPwmKc9OTItqjoSS5nK4V4E0gs
cVn0Z3mvMzw1THuxSxgcdNTOqvzXo1c0boOBHVT0j9jNm3DhgFZIQtJ5yXpYikCSok3NkJkfyJ1p
g4tv2MbQZReIfpQGyUlsz9N86/lrPWRUaKJJ8cIXeATDgZvhwioYoialRd3yBP3mtJfy56U9tHHq
HF4T0IqFfmGuXddznQmg1snSDMnupIFaCeo8gI/sqYnsey59U+R59qcUrJYODhUlbJ0E8XQ5bBX6
PrWOtMctnVLAeuh+zo61ouYwLBholmL+mhie2F/7wAQz5H/bNFy9sMK8ocJHkMvO/GoRpnZxOXLi
kNJvdzu50JlKr+RNqKTbbu+eLGt1FD3bIVoQ8Kvt9biwjczwUPX+wz/rF2k/6cgXXGkAA8cPDd70
u4ZuNQwzYmCZdhfr08ezK62XX2XqyN3a5WCKDu0nd3RR5KmD8FHPSmbPdaOeoAPxzQvUGhqzyNfY
0Yf2TIt1xJ5fkXnzoQZ9p8IQtatJGhry/p6b4/wXG3Wil5j9XjcIm6rgp/bavoXb7OjTn2TMGf2C
9tsZtFkeQv3YEjfhcaN9TumDHnd1HYk2pAcd34m6DtBhRu5f0P6SBHtOzErPuboYp1/ZU1W9jYtu
8RAuLtKghDSY0Y8Q9MMojbJ4qRVjGPhtScATYrgrLWUSpO4LL+gdm4uDlBhBPVW7TQa05WR8a8wB
VvqQeFMRALRRazIviNdX1k6OstFVBlGYN4ioaM9IDJYhPeTPCwZEnNgIkLrCsK/IRWc/jFvkQ/7R
MlLD45e1UTTxrQlJNFimJ+dzQzr9r7S/897k5mbK4uxRvKkbWXtFqiIVut6UI6mHzVZivI3gaCkF
3cQmKAUl+Az33JIXBTHgflGzdN7fFdxgEFsIsa+qk4RtI7iaaMppOelLttfnJym3zS+3fezxLTSF
fVoqUAnWDUGwvrmzsZHsjVz9Ov8+IuM4vBRAQpClYUFZR+13HRfKKpWzhs1XvjWwYmItFDCvie9P
nWt93KsEDLL6nVZsHyU631FtDL4H/FNuVGOxpY9NZJKRmHQoJHr+RsXacwvPxp5oVBZb1kaAnNxX
jHD3Bh51l8bdLvPR+mgNAQUN06kwHmlTXiXjDO7UxepFpjs/sLDnE+Tsmr6QjX+CMZqoGBqazr8a
8dms11gGfx2GojCPTeb35DrMouvXiQwF2NqjCxLVoWYVrcTkPF5tDcDcVQHiX2jPH2yuRk41rp/5
7+9jaRQBU71bXPXEU+z68lZlpj731NPho6r+DFu85FUDfj6HPF9n7Rcad3wDcnMhn4dKO2I8MvrJ
Ymm7JUgwwYKx1wzs69A6pr9n1lByMGQoYj9K4ZVIVo605zUn3968NeijvIoPLnlKeMaz+9LxgfJn
u0d9fYwQ6fyg5mHTLBU0+kC/s2vG6fxEOo//95BMvMAZ8EZkhYwSqXWlF490ithrmxhKIM0X53/z
f/3T01AOQQtIntK0dTaB2NHsf4hh/ftZHqYmxPMWlVBnELsUEcdsYHs/kkotu1XEBejvF3O0329a
c+OoICXxPDZGAxp2D7gwUp1pR7+oGk/pBjfkLwrdszL+XrdAehqvw7/Zk9GKESBBQk3trIUI4awX
8iFG5W9oQyAkFMRMOoWU1qy46pw/OcqsEGcdNcek4D/Ayxy0aWp/G90aL7SZc7ySaW+To9BUuSKk
IknbcKINMofUkkIEvxNI6jkn+A6ab7BOo3l5FUsB9J4b2R660T7ZNOvdCP0jnFlmDTDqZSfaSm+W
TlnMIjAnWzTXD8PIFXbOGVb+EmzKLUH9fqqFUVOLZFaQU8jNvDiq2VC3I4OwDVl6xtjn2gXRTDXh
8yBcURJRpc4FrBy3CcIBSOSb1OOf13nvr+NJM/CfixWdM+kWp3SpTzs6YILvVOTn+dwlToMkC24z
nn2reOwSNxkKfytPCwW4bt32Rq2eeOubQh7hv8M+G/FClmuGb4ifeuwplbjqtSZheV18SJNFFrwm
iWvCPuj8QP8Qoc67FEmMo3sP/1vc9yJUouP4mViv8Z9Ba8nlURK5Y/vjtjzZwXpsOFheLcc6ZMH+
Teux0XH18Zra96sHLudIME8WhdPJEWY9/NZ0lLX7kfMR6E8BJ/7e0ZUDyP7Qs0oQHKExLcqoSVCH
6FElNruiAF1oVbqF1ILiw0ier8k2efzcUdIwlnBNKN08jLjPMCSGm0o0kP67gvdkUETFNnpqxMVq
MjlR04ch8MLAksK4aAtagFyfv6tPGft5ET8L+j1yL9dRk3N5eyXWlClQn0EjtpqYFscfrrYLhxHB
sbnIrjF2QrMVzYwh3WVqKYvJ4cJf1myEB2mT2kcjUyzrF8lvZy7wyQ+2++KpFpQ/ceAVwlsHISFH
ea4QVusj8UjQo5BV5dE20hzTUm4Q87CyW7623T0EGvtDtcH041sjo5VjtkZ9pS0sgD86n6S5XD7t
0YMB+574JOexlBNDnjUPPvu/eNhca9lVgK9ZVJLyjFOJOxcZyqxmHrjhSfW85+QIJBx1URKEyJar
ojwo2xt8X7y4keL6s+W3V5qOXSdMU8UPgfiLD292ZCLAqvlN4qloVOFs+oRXuji2F+W3odPYq46P
njMulDvc4dmXba6ms7zaBl5iqP/J/xDa7RXzo0sOWmnW7jX2WVbtQBRRGjoO3zJ4T+eBbca6eRNu
8632rSzDwVWA/soHR0Xg08vBFkCtrV5inlTvnynRk4018LdAw100cQ0nBmwqBhPMxYn4+JWw3uzb
zfbuxKBp3lcOpec4/3R7aWM8bhKlfGQvN9t2HC+qan0wyAdnDDd0LnInFiUhySWj5br6VdjVAzq4
wTE3l/6qSzm6QCEnmyQM7nrVWC98K5oPgPaY4PG3vsKozYOqqxVigU1iT1a5/Qn3dN1sXY8t3V/Z
447MhaZY4xgMEzo6nkOSwPsZPbq9QmrCEWvqvZjrW4wST9EEk7yrQBHijb3vXn3mcaB3/HG5SewO
Fxmuq7UU3kbosoX6ZhAq8ACmyZX2F0yj+Qu1Rk7TUXr5ZcnuPbRwRICVq+k4d0oKAwhAT8kS5pq6
dbHQd4wgs/Bk/I2pVXRIGsycwfJ4ZeATeWT+GgjNaPBQ7IVlfR1BgyDDI7VaEgGlZUSmnR+eKqns
neJSEKRiy30fJAc6M+kwM2/v/unjBMO8AWsLQEy3BCLFOoof+CXZr5FnladfHX1+pZzga7jJaOeg
0b+eyU7mH80xBf/GqdgQBQhICA8rrB2dU7Pcab2FaS85H1yIdf+t+wlCcDaYO4w7/LZQ1jy3y4lQ
hYTDvpRCsVC0MUGv8zJlfit0kctZkWb0xYD+rqLkX2T6UnW2GufQJs4crBZqDx93HPiZNRv9cjMK
665mIB/CxipHgrMw40lE+9dKG2ha4YZY97G3tuu7iu5MzeI7VG72zKHl2Ig9hQl9NkzJZYO/rnAR
Hp1h4MfrUzIrzy7ECDrFgl3owqhJSd+uDIFkxjNzCL3npgfCpw7+p1EQe0bUqMC79pHpQ+qZGA/L
X5W5asBci7uwuGRXwQxYAdH0AMlm9fB24/781EtvMxiJasEu7biboKKTjfK5UTh3/rnVjkZUL7zM
oMr3O4OIXmx4eUMmNalfUo5rOfNMOXhbW4RjNGn7qb3ywYPx6Cn3t18sATPQPezQNUh4BfJ6VOVp
Ae+nDL/aP60s0rOvOGRRWOoWKhtYPUmLkosj8IG6IgUz4u7ihG1xyRrOHXcJ/P7d5xMhPlJB0eKj
nfq1p6qro3WANe20a4ctW8YTiGneb4CC6VqCXnJLmP498DBuotzoMV413twTFOlfdqXi5ayJd/Wi
kXAzZ1tnXNEe1wJsbqRwxF4rudV7IlNVjw96xp26Si2RHyCa5CAJ4lDWO7CTDa7HnI66fC0FdSJf
WR55TDUtiSp9qju6mhNzQ+pVarlzrHeOGu2SihvKpcDykWTjiMK9egouil+QYgZpSPBQeedYyegi
/Ekc94PCEinfnaFHV4I1wqOlHW8QYjVbtnyLt/fomqVThPe6IAGNGJzL81qm3hrjSBRxcFX3IWhp
WVYcgc/Y8iBYpfGoSpmG6eLnmjYZl2gwRZzbL/WXL4wvvW5Yp3/u11JEZyEHYZgm8zXTRH3yhuNY
4ifw6ACnbE+cjlZFKvp7HUmap1Y15zIu0o66AoG3/NVWR1CRQhKv+lkf9OmLWBhdb6qwhLevV20q
ZKs4P5ig9kzkNaXHl1s42EoNEUnZfTY9CjKj+4IhhZlQzPizdl7fsVN4XjWJCQxlJHw4K9Znp3u5
OsrJ/E6YgdapoOpmLABl4NWv+enPUBm3kOVXfwc/2Ly0kbIDyENCsEcDP4qWnIlVkqgKLQLlogK2
Nc/OWCow3e4pCsGd5oKC3itF2AbI8S+7xoQHFDCLR16HJPBg7pxPhLDfN/F+pYhrIFL/W5kpu7dO
jbvKyROL4D3ceenAAIwwUQgLVQ9kCKjd6CoXW0tODzs7epzsqUGnxl3I8VW4w7EM+99T4uQRPj6Q
klYxyImWs8IqXr6lUn1TMJnbHL/T3lIjpu1ySktuhgyWpY399afSFjjtvsEiMliTVZiQFU+D7ucX
IqstJgdV4WR+wF5gCwKngqqW98zf6/tP84B57R0Bn1iWeypMydT0i4Crz4VNz26jLhTh4/KHLDbt
gsR9iYZqSfU12bRu0tQ1pMBsxB4rpCoVpA037QkUeAvhSytLKz38+qt/4SqA0pC8iB5VEWmTB0BZ
6+AKOEhrliKHYoZkTBH//vysxleHLvNqJy3xQoK4KFesbIXlz2voIB6UIkxueIQjsILHf6caYb/8
oaMSd3bR3TrTq4sGHfBlT5ReEa6o3d+tzFKSVAonXb5I7IQ3483+FMu79Yc7kX/KJaFQLrUGwZci
vuoo3Ap9/dPUpA146XsNYTaWe+ti+v9JpDlO+M9ZXUaoo9JCnoR+l4cFAFfbiZQoWt4AFsWd3wlz
Zsxc+Ulg+1Lkkqcas4Qq/gO7cC4wK/LQ+HQisnJgrwxhRV6HctomYs525o+8Q5+mUM2/qJESNeCH
EUHgryp2RYi+qNi3/jN/ukRbufCtAfag26HZsKZDvvaQj5oitT/lPySbpONNwlLEDFWzYXFKeRpf
hf8kK/bEyNb/d2ajj/S1qsyGCghEKpzG015DOEyvm1/eBGtTkHaDX7hdWoiSRQGOyxmDUX7Qwlfv
dP0ou4NunCiotzlg22pAIGSo60+cWtaGZcDjzClGA5wvKbnZDP045Eycj4mgZDYC5hqwqHqPU+zN
pMUy4QLmlC6lb/kvvt0ZRq2MZqwK4/Aw8914XiXUs1fUqXGhmgaGJhKIrLXsuvPy5tXv1Az9V3mN
S0QH9i/nij1oaCvOEVn52sV9bUrvsq5W9IMYUrPe1eI1fr7xyTX2Kd5LyA4bhOAWal6u5sz3FUb9
YLdu8Ewk9IQuP0Uqwxhw/YYLOSxDti/byrY7FWCXD4+Bmi8EXqL+N+By5xorICIUzHFPs3sOCPbe
U2WFPj2CK5e8EGFWfyTW9DgF+EA0WpEF2CjlpeECsDlaP1hyNXfOW4dSZWsNK169dWG3ZQepCzlN
LRYjhXwQhNy5cSATnh2eCFcBkwOCqLJro2gNjfnrSefppH9uMrBTJBhPPp65FAXPpyOUjAIFY4Ml
nqGRuefnwXEuZ4UYcTQALcUpKmqWjo8B3GbY4oqUM+SvUpob3vfCPOtEvif8KW2GE1XfGHboF3ty
BBzW9ETvAp8p12EMtHmFj8IkqSbaV6p695KOTOigqggIRqbgnlAtw+TLGeFf8YBLgLp7ORaiNWc0
Ji975UuaPDcYZ4OQO4Hua+KXAyugKwPnuOFP5tEsWK27CKtQ3hL/kgmgDxCEYJQ4xNDztv9Y1ISs
hnwhpotgaWM4FZl6xwmF5zS7EMb8Xxfgregtkd4yyVV8ktdJQyt41bLU7PHC72f5XDnidlVr9wft
Rv5R8oerhmoYnVJLAKc2jlhfZEbZYs2zTqHNJ6sUEI4XpZAlD99yvFNjuHHOM/3Zynof4sn0j2Rg
DgYz3Ce5F5s6x1Vjc9B2wY96d1M3Ev+6FnNtsD1EilbUjrISQITreZE3McuNN9LOAWQ1UojLXYTq
VWhIDcsg51jlylYSpvz+W0l0Nfl6yKBOq4odeftfNlnTJffY3z/cA+24iYouj/fL5BL6vtRQlTfd
sm6tEJUpTxg8rvk2Bfc/tv6C20mimLbiEnwqNKB9Nt6ZdaVml1BdJTmlBiaSgsqWf52j2PRqC3Dz
eSsmo5EtP/7K/LttSLDxhWmuLkeklpTQE1EifQS8m/zecXcPoPIBjVDggiQbbZprZL2yFIqMohvv
fVF3h2+ADoo/aJj5NQD31lQGV0cyN5kB9chmjuzZZM4JtJ55btItgrJcC7D/tzQW8uRPfMULtaPN
kjbxOzPSViED8D5Zqn6Z35IHKHoZLmNYlJw0MYSXeixHNJLRtc8jxG5tlbhiIG1t9psf6k57sJqd
opOV3P5xFqkF0Vu3PC1qxxUowm5ICmcdlsWWl3r5H7j60im4FwwQO8nIMkP7LkNxnYzHMh+1PHBl
F20R5GBW3rgBVBsi//dT3MyJPnIRhAL0QmunajRXImN4aExT4EyhwBmRs511rE0j6sd97uFi2HML
KWwsX6oy1rlTLXfO/X/1/NKL3BTiPbmFkoWEmnqyBjsPo+8Y1cFrxwfUfClRUj6wo6XJu4fMM3Qf
l7iaMGgYHU/127TgGHvWLvXtH9nEmH1gepwAGRBrYgd7IuLl7RYIIN1gVhdAv3uODyQI14T2kkIa
HBiad4jm8maYrGaiofGx6bvr9sJbfbsv2KaMwldmAIyqvevzIvkWy30hTpFDcZjVgzAWCtlBBAbp
MQGxRG5B4q0kvqvTOQzuFRJ2gnVH5wX7Ubp/cCJjHBT/1m+7iEpFnAYwiDQqJSDxdYRmx0UQRjsD
yGHkIXgvvQmyCzQ5prGbGLa1sC+z7JOBHx1HjRK3VpV5M2iG81LrKRZ8NwNVYF9raFoK3axwDs3o
WfOu489yt4UnnQ5pe0xCFBm9DaNDfTA2Tk5yCvnRS1qTNH1gaaDGImEcOra8oYDVWRc1A1mXf5mA
fzYHX8V86M327eN4ZGibESKUDELMpwlPTExmwrgZQ+WCj6CdJje9Ao3fnwk5WY7KvhpwcOuQAIM6
W5hz2Xpc1PBkv0zYkVRyWIwrrj7skLih4UyecI6u0UtqSWFz455kR+tzu68mVyUJCXcxPmF9Ikme
Ld2I9nQMwGOqCRND/y8xTyCv8wV5olG7m6glApDH7k6E579yUSgapukdLHD0A09L9okIRaAdlVsf
mgHd6Wa0+5Ge9F2xeHB8DDaLbN5HroWPOz/Jq9eMNRr0nCcElvxIzEiZUVlRrt0vS99VbA9pLYIL
f4OZgGJhnh7P+rii1vM1pw7mv/Pj29cP4L6CBxrU+JgLODYrfXWBD2qCtjUqQ00dvWPUVk7KXAx9
b4AwFPVZYFEDQ3uoOcUQnu79atMF1/T7vs0JEFNJ9Sv2yFzjDOK1cmTMCWcSNeYj6hNVlI/AMOG4
E5qLPVevJMnAwafQxS4Ktql1/J7CCoA16Lw/UriXA4H2HemlEsOxfnoY3cwuhgRR9FLVEd+yrLNG
vt4PcYw4AFCsl8xLTtPfukKGIx+WN7irq8M8kc7xVQfe0RXCqwZaTcCz6419WTwollfeONpcCDGm
NnNivxR5H/g2gS0X25zh1SaI+MkZxO6ZM8c9okD//zGszQa0XOOYTwIwFvHJXqm+W9uaEn42xpxH
hTVomdJJRIcjspiX9IokWtGZatjZnbGldSXc0Bz0H/Sfr32GWlbzjrQVvuxItnnN7QMqJgdWbeLO
IX8sx5Fl2R7ncuPFtB88X8Z/HiaGNXVd0FXmYEjPhwHiED8oWSyARlHnbKp+5X8YUtWSY9gpbd1S
qeVdLAagL6HwcoAIBq6OAf73nRUP11MfTIIw8CPA3UoCUpKo8AepNCrJo9XWy3HsHLk8l5IE0m/S
7wglEVphWKwEhhzwbYI8AteAujJcobSU02xgUExMdR4uQQSHEY/a96YKy/vGB4UrvTF0JcfUJ+DS
cvJPDNOZ8jkC1vZimGAmtO5eX6cS/uW4ihdUdZhgIwDlDhiN5u71DZI9plVk5QFGc83+mltrDotM
ZOAViB4ZjH+booDrpE2yYmjXucf5YgKy3jsIhdEZUOpRB6SSRwC8iCBOJzrZDTNtAbK4YrjnqP2h
keYQOFx/+NL2eu6ANr8eJptfSEpK/m3XpmqZBWbYJtvEqZVPZY/h0uYj3wiqrdF+sJivUtUy6RUx
kXUHQt1yYFa3JhZuMTnVXqpAF1dYsmqobmIfgYR6w7ukm+6v+wdJfXm0zIihP5ylME+7UBPq9FAR
Td4FBjEd43FYmVcgyc1HiM8844tUP4NyKAguduEBEWEkUZS4kDqrY96MGwsgs0/+Mo5OozMHJOJj
OS1E2VDDwVwb1r1VJw4gos0Pw1hYBEJIhs9MmbGMHCW8VCAimrShbC0V5x81nGx88bdudTNB4iE3
FkAMwN0OW7KQiUXcj7B81DjqAM1ysChT67Urw0TUZdn7/zCEiPrthjwXXd4277lJOcTNsKRoRNcC
YHiEXZ0aH/h/t+3SwSXvjphXiOkoqjchbZZ0owfXP3FpzzLD4QUEOWsS7pQN/9OlHk1vwAEVS5hO
JclnihHtie4GbOPw5onfYIOv6BKwPu8WOM0QuO2WEkqUAsNTGdhQHsLRRK34HTp9E8HLfFIf0ccz
NkxTUSjIA8wrSdaFc1inhQ2IPhLTwRnnN7dmfoACIa0fzVB81F0UtM8YPSHllULWVlY/Hq21KIDv
MxPd2LxHcGt5oKv/CeBCGFc8z5bVQ7SDcvYXsOKqHXy+xHoJxmq2dYufaGyuf24sFNHBB2TTLVUt
7gEdwkZ52SvyMrr/9rsWIbSRv1q/q2wAcA11c5OLG95PUSnIGfASjkiyzKuIgRfoVz+iNUpNM+1K
5BQppSkNnyS76KuHlokBLWQeNVfDCN2y+ChCPwWQQqH3RXHlkla+OJ7zhF7tCgUM36OGVL6v8yEH
cCDx/NjM1QrEPtJCYjiBh+hCZDDdQdzfxb57vkttaIY004BcjUrzKtmkjYutEVFdkXOEwT5jpFS3
tvKE44vSf9KJ7cXm90Wt7L+BuzzztFuCIWje/CN2gsONBGYxOE0wifCze0U848hgkKjbSbhCyMC6
DOa0uWxlKuuq8NTZBhyb8Sr05URMF2UvkFWLUpXizuya2ZxMyW8/vQGJawapAAb9wg2UbXIXOwgN
kBbVhPM6WXZE/YcPUrHRykI1o/MOrfJiygFl8bAMJz8bhegiyKW8gH8850yUrf+M8Z9Yootng5l6
UQ1+4GtYfTqcnwGprJpOsmLK9Q72uM7Oxhf2JF/2C8yPApm6NL3kt/NL1eAyrVCgwk8/wcYPEBSg
0NGB2PYoITZ9mdLaOKYM6zsV784xcrXgKsqzQocLpqKMHsZCINnZU1WUuWsmNyDrpYgQOXAYw73v
h2jRRpzNU+cRRVciqtGqDXhG8uWds16t8S9YF/c2+OScRKRUiBTHl7QSXJr1tW7E6GDBEwwCZBVY
XsPwQMaaYDA6KGkKBzGvKRkzTIvuMcrpPLS15Ps1zhBxkNq5ajK3vwJOrJykdY0oVzbeuYjRolBa
ci1aMIqxHwbqqv89mfxufzyc/0VJvf/X6U1JkouWeU5GBxNmEWKicH0P8sCwn2gHb6TwXe+m/hWL
+GiE+KIV/iNboIINzp9b4AxS7lsEwf31Ta8XzowhjD7kKx2JYU9tHJiXMWc/SE08qanG9CnFDCTt
o6C0eVSFsyMOElMYBTBrb67Umv0W3vI7cxFXbylonAqg3vvQsLLioyEl+cttvDbHI9UEhJthvWwA
I7fwlb5QAvrubDu+szUqknAw513BWvoz3Iigpeoad+5TV3GXlTa6D4QAczGVmo6IvmLGvCq6shGQ
mfDzkPXa8IrWmp/J+GIP57X7SM+vDUgtBsdPHnROvM3fZDnICbCLazuG1W2X13e2P3EMeGzHWP5g
3U5ugCRws+cq0eJ0VWax+5tR+elwUyNKc8HoqwQGFsSq+mau0NUmTJwMnJA9T80g2iKEdL2jr8gp
2CBhwwwzZCU89c3l7P0zU81GJHOciNYn0kzIorhQjS72r1x8o1+vnbcQE6Y30NTF7M8esCaA9YTZ
XdT6Y2mJvBvtrPxAHrlkE+zZ2Ym2oGlWLWB/sjvcAYPDzxoOF+M5V5NW4xWccmdREUqmERUajbhq
l9oYYUJ8FwFg82t65um850OabXi/CnKa8v9vF8Y889z6uF3KUI0mL1pyy5R/mwYrdfSrzjH9pZ9Y
Gv6pAzZwSsrUFol527cVOUaTpCXk54GJet3oQ5flOjHtrKcq3bAzkuSaL2NnCx1uUcHWqR98XtwQ
owriHi/5+Rb9dP73EkWtBa18F7kC0V/8o/RaCcEjPEe3XdaEHmop5CDqfXMCI+TiFrlq0HsVG42/
1sdk3uJtewMIQz+eQVcStlh+DpaG7gCUYFoHQ1SyCxCJtnuHjSOqR2DlN/mJ3dG0VL+0wC1mzYVQ
s4cfxiltXjlAZsguRNqOoiAV2gwFZaDEXtUsXKLlhrkYHWsm86sYdrvQunswC++jGlbHvffmY81J
Y2XLtVJmGEBBt/hW7u1GxrdI0/4JeOYrmI6rpqJCwCB0bJI6OW5BJQNPsc6zwyXMfiGXtuS9kZoy
PTwwVhsi3TIBeUKe6RUV3C3AewvlYaV2bnCKemgTGjkOANmhrZsv0Stp24Yl5eFXtwf1a1n+4aiu
qwQo6L3jQzuzZAR/V7B5aGnfoNal4GVfwSsmGo5y7+pnSb6GY2/2aSiJ/dGVaBLpTFap9+d+h21i
nHHjS3u+Bxc2oRGtmvbU9x5zwy5iP4tsLJ1JJT9L6Ku7eZkoqZ4DTlnFI+YlD3NS9ti/xR8TLoec
LMXdS4IHmWwQSzey/Hk+Z3R7ojorZnngmBCaBR4Fv2scTEXpA2XOOwSBOO+5zC2A+Ndb2gQJw5O6
dEdnMyZCM67HMoz3W0mU7MLxEvYvLD14L4GWg0lM4rqwbPdKUPpczmgHqrepTW6+EdH1GeRkaZRd
z/8uiCSaagCafstWglnwWXfsBiv7BGiQcYzqPQ0aVpYNuVje4IUCygwTkdc2WvxTGL2zCRcL0o0i
ig++pI1ZMs+3JNxQL94EIK2bnNjzU3EB/tn2M3NaR46TGx5xhRWImFGsBRPLpXnARXkkIDQKUoxi
Fg9eQrgHIfecklKKjbAfF+pq/rWbWuum0f8eyGaJwm7VGy/hbXBT0bPEsAiO3LfB8yGb51SkjIQN
m/vsb1imOEH/3GTQQ0m3qCXz3EOyvBHnKfcxq37N2n2HP0H2ApPGl9FkfY1FB81fEm4NevpDR97r
8BUsN9ZULWO46rLcVSOnJhAdqn3NNHbQ6T12hJJyUXlqfgG3Q9XnNSVTvcBypaKe0Zp4sVh+gswX
C+hnZziJCPvAKskXwGe+5bY/xJSpfjsC5US6I+yNwuZDrlOvT4lJx3rseTd/yoqDBuomjU/HHdOH
TZAdqzSuhVGOwJhyHibm5gVMf7iOGCn4KtbOo31fcpgF/8bI8WQiVt0zzyj3ne9JGNEG2DqGxPPU
wEmboNxxN2ZdGxTLESYd1r4CfupEAB10Vxvikav7KsKVVPYNGyRrco7KlJFUyhnkaXaZFHJSem7o
Qa/+tX0LN/uwss9PTwe5CYJgfmcF5FLOAzovJezXWL/QHFS5yQpvQe0YKLOPRR1+0COLID9vhGI7
PrNjCPJlVthKdalPB+5iT4SzhTzUyxRn7l3t4SWKFz9FO1yjxjAiE/vukJ1vYQxXRhHfWYiyyU/3
/0ZJha6B9JH4VMuTGtMT/9Q6OCKYRk0NeA16tx3O4lV5yt4mhB1elwjF9IONM8IGlWlJO4Mr+LCj
epMuBqkR/ULNRn3L1SDEFD2sPZv/WkEOiLymZpvf2gW2Tt/sj3LY0vBdNxOzSaydukhM53Yv/6p1
+1EYs1XoEYoiuw16w0kG9Xj8NZzJMk3zufJGmUVWO3TqLeimkGIXI+MVfTLmMXaGarHzBMm/FZQC
fQHDZFti3cVjsdnUoqjMndJ+Gj1vNevrbDA8Myczc+TswFH6ACm1Nj3NNmv7hztKRlMmwO0hfHVW
AyuMxP841SbS4Rj3BAUxe8GXvCP6iACZAlOZ/WyFVDNbsppHjtrTyCSFXwkARgOOD3ST4XOBQWNB
tqa6ATRYC/XU6Fiw93Cw3aIJQSZAm6GoltmREzMA5A2fjzMiu68KyMinjzTZX/2qN0NHUznGkXMg
L5hSVbDKAVTh53Q4TXKG6uLHB4s37+mPBlfijAJf/Lv57O4tcpvalYPg9mFyhOjkYfV8K4KFqR3H
TpwacuddnbT1IL+TF9oaRxtti5tOQ5t1Tvc/7T0VC9FgqEbbZK8YhhRLlO71dkkhQf0hsuPZuklX
IoFwFNRwp1y17sjpGfXK0cX2/GUqVe7de/sVP8vqyWgapGmlXNirNTXNG7ERPsRPHWwQR2fJRDV7
+j3MhSpZT+cu6l/IkHJVqK+flYYFoWZTL/R/VmanKhovj560Ki9wxC7i+gaUWb7CEMvgNdKYnQhu
QJeRV/ksdlskKZiOA+1K5Nxb0LqA1cutlaDjtaAZqwpJLFrRecd5fDvvAUQVoKhM8G6ROyUWzM56
NHAUFpVkupOnnPJq69tcSa+6tRqQudt2z0SaHzYOvTaJb7Jx7l8W3QEMLHHpnYtDf6Cdx5nbWlqK
N46/jzNj6Eil6SfLHvOCMfsJyKiewhmf4N7Q2nCAD9xcCuIPEM3J7ttFhBjqFEyAPoUahhtRxmM7
J9VOQV+Mxwtbaf/Eee+UONS8aJm23f59WTyzOboVK4QZCa/kPHBmea/XEikR7PBsA8Uneo+fr1ez
RCXPIXBtbMuPYuUlIq7NRMT7olPt0TosUcP1Aob4R0HgEJvR6c8yVAoMO9BDmJjm8u7LcwDMhJx9
iEl08239RgeJx0NZ4mWpPR2fm/pcCkvFM7LD29Fz6VnzJDME3nyJAIZGtfsw1x06A26LAdgO4h/5
nG6P70l3Nod3eW9I/sZkEHrFifeeK5nG2TdBZEmiyUxrEJN7+Oy04YpmO+QPCzriOt27M2vXPgPV
XEzoq9dScv5AAr4As9GQtf7iucCvQS9Olyf/k/sYNtkxCPJjTM08aDZCECGnVJXdCrh/IgUn2s1A
znQd4DxqdBpfnHLhy/z/yw+NzdUSHcHfxG5DoU1vFFR3x0Zc27UDAoPvMMTGY1K0Bq5+8ZVm2fei
+mhchn/vdlrmtao90UXs2b10Shkl7i7YIbLrcUq0DSbBIYEL6Y5LDuXDvFFv+Kb4hE26bI4fvNXc
z6C0POy+AE50XqpgKMS9FSuJkX7M9b3wpRl/0dIFBhJC6rIL99X3xUVrSld0QGAR08lb/m50lCKZ
UlcVtn3rBShMSz2oY8baZxtpREDxJEDjr/NNrAJ4LxEKLd0eIDCwmzHuRTuQPeUXv4uIOhKjnOAF
XRHGHuVUteWJyYgO9o5W+reL7Pkxk7xbqU6f/6W/ExGNWVoXtgsRge4/5OQNeknFDOti+apfN7nK
8GsuZ9+XNWg3Ar188Ur+kcN87q7pXl4HQFJvSulM1Wf+BPMxEA5pR9fnbF5xwNqI4JBmfn5nQM26
VhLwcqPFaihPi6U4dAuBosr4RynAkxfYoG7g/V346ZGPsLr1CkW8v4FZeYJmdQmLaLc0LtS4ODyf
AI3dVxYwjseFgp4kPJ8AqykEX1QHOdjmEBcadVHr0uweh8yO5mkrh6JzV22Xo+sZx7nVMkNSLMtA
sAWvs9ZZiif2rzZyYv1x3US0CDzJXwYV95/fv0P69RXZL3y9u6dhFHpRF1u1fTcKJJLwoYCZr3+P
HuYQZ+lulK4bBIClzy/h6OKrrW1mkI6uzRddmhZ+qGRkthbxyJI0VUWmUJsjW8GBddQuLZRkM7lK
5iSAcgwpBhK/1i1hKw8Q/PF+3CtazYX+2SFEDvK/rqq5KjQTjT8YJj1Yr9UbgQQXh+hB06A+hX1Z
tmyHaUVfFuVgBWIl/oqmb7DOjJbXEVLvvP/WvkCmkAD+7w1axI4a4L866fZZ6p4PT001ATUAb2xL
+F6ejdqJdMCF4aDUuAcxS1Dc8wYu1TiXguopxQZ76ZvyoyIUeSqheM6Bt3xFspvwN1R2WRwf5jCu
g5znr3gAwumOxYznqQX0qKAYzoJeLD+qc2lrFAUyfBKIvFez70KHAC91oJUTsbIBNn60lk3AEV+X
j/ksFMg6tn014clL1Eo4CYFLb3UTFnKNcH+CIbWP0wxCCWMMdYRb6ll+qvdlsyfMPNpde4TZP/7I
fpScTE5rgJaMSoK+IyPuQwKL48Zs86Va1clIo6NGG0z7k5MF/kHth+LdjRePfsL/s6WkVO0Y759F
zUy0gYSaZ2o3B9XOJ+42ap5ewRyXsUu1UqbDxmL4tWRIOza8ikOUTZsQSMkjBI9OYwZrGM4V69j7
jcKsfjgTRA80KZqHMY1rZ495g3MfTandaLSvKIPxLWTFFLIuhpHG954c0HItBUhNB3EMddOjilaD
M8B5IKjnjXgAPnZLp7gOi8uhmV/V3mZBqQC3a4S20+LxrSr2/PEFk1TqPINZhv0NI/nyeOESAERH
bD9oIvQMdU8BguC+JKU3R8rgfly7rZ/ysR8eO4E5AQshC5AQP6pbnBRgkpONCy1oNh/sKO8U5dYP
2UOf1EjnKt1yNfxsqGXVnqi5uSEUqlgHnDa0mabzfACwnUYCRKEoJOqfuwoXnrqYST485bt/E7xN
xrIrjgKp0sBopx0N0CphGehdeXA13lWPXlBjVtPUGPg4T1tlHTl0qp55feYoKwQ7m9ry1xxTMtfj
Z2alcea61sX8TIXRcgmZgVDawdtBzwMvCplE7RMJujAxp2vBQiEkFVsdvprmgwNCQMC1j3gpsZmO
jku/WYLSA27njA7c8OdZClnlCEbz/i5PkZNC7sAO8XqBzVxfAO+boU1/VxfgrxVNaS743b97OnbV
D2uX77vOOciNsQur6wtATVw1spJgAs6uY2PKlCY3xXIZUtOfXSLrD38C448HuOo0J+2WGaZYCZH5
NVxP8Aw63a8O2Z7YEam9JhO6ew/CS50keJ2oN7mc1EYRhjl/AX9ZDZ7wcLBUFQp3h1iDv5wE5+ge
JHsxI/nhDYEtADykNnWhBfKQlVeBSGWgvpcdz3yRXN5gChMTO393XrhicUnVLE+23JhlY2VCkuYW
PDIj6xN0qXYUj5fs8Ff8+Q0EnEP+cR7WonNYg2zJt80c8F8HV7TV89k0ncjQl6Xn/EAeGGr887q/
FODKlyeI0OpHz3O0YSLm+6pUJwvxQ/xJT5jfTlowkznGoQ6qQdhYr4n3zwFJH+IwlmINKqaDqQoo
7cd96KJDN8ericEaqhXslxq3wsZTLR1fqjGkdDEaOhIbh+Db9MChy9BuK75Jm60SUwMQ6DsFYOuj
PInfVhzeO3aFEJHYsUU6Db1R3IkIW9dezraVMR71EjiOk4fy7eYy8FziDZyP7oMm7V+k/ZB43Yfc
OXmWx0rfrGro2VEJStbCbD0uhabewLuX1jEUSaJkhateBVkRcPuTa8JQgRUZ04whFope091SIjvh
BjNqvfTfl1XMQEIymVtE2zKCS6SHM3k0qqRp5eFKRrT645RFltthx8Io0JRzcXgFzolCM2xSIpFV
1/c6PdyEpdi6Ogw9vUvrenIwe0PpSJ2XvDuD1I8tJfsqDNHxuK8qUANfLimonX+HceJ0nxm4iuKx
T5D6GNLccUMtKP30MEmmPoVKMVXbZMjm5HXk4z+1tQBywnmvRZ5RYNIucMcHszqhubGWnEllJP+m
FegLO7a7rolveC5C/oYdY0w4SJsAyDdKYQQYqIl3Uz3HSKKZDov4K9bzqm2cg0pLwx54RgUMuUP5
11B810szVTKLsyml/2XdtpOeXR5cB4zRV83Enyw5RVXHevNbc/KW6XUrxhpf2anGiabxXvxiBANF
ViW26xyzUaDzBaZ+RTPaFVnZz5r4XnIYkG/GGeSmVQX1yQlUHelogXDbh58ic51tw3e+iV+Rv3QN
tpTmOHau5Ac5CavYVJ24S+nkBNhECOqvfXvaU0bUpOf3o79sCRUSXzDota0n0dc1qVTNi/p+wz7s
Vm9T0DQWjCKMFoMrOpu42BczFZv4ecYf76NMDFJyljcFHcy0o/hvHkr++flMG/om6Iaw4N9UW69S
M3MUgoR3D43FEZI8ijPaXo3mgb/4YBtyCi15pp6rkWERj3q2bNByQS7SMASSTghfUgtCA95r0xDm
UMkS9EpeRoAt6YcKfaGJYbmS/JYyv6yKkaLz7kND2yqvODleYMYrXDbk4KaNseYg5ojRoxbfUj+q
PkyHXNjarsAI+VJQlW3Szge9EWyhrBmLDGRb0J4ETZo4c18yvSbn+q6WLv75ShK6WRHdO9R3oUiI
dq6BbW6OZKhXDr+O572if/oSHJN0TJTSkzXJwamfySe29fafY1YrFMWFpoKzS3B9jJUPTx4hPQVR
GqKtek5ETHxjU40SH0pQwAliMgfwk+6y9LaBScxhEVw3KKrPZKWrbAQFe0s+t9h6dCZwjq6SbOcK
BxFS5lwWfiC+z++o8PGB2grCGVpEjqeKfosbn/VokiQZo6bcEzHQoxSQryizbYmk7AhRYfFDCD+C
kkUG5vMAaUzBYfi43pGsW8s9Mv6H2DyiH9rUKUFsrutYCE3gt7V/t2JdhWR4H92/HsaQFBgQDhEc
1ORfXFwXIGvbUL0uuv1GJX4tQZ2zz8e72eFljrFNwF0Hd9OAxSzeQs0oHvqm5MmwwSKxLbgxuP2I
+lqALb0gwnY6HJVQO26Cq6aLLQ6KTCLEBUcVZYKpU33Ps/qbwwkKyzwLyT2JuagUhbuTT9BfPYbr
gQdu8/JMwF09Qb7OaMUfCdeNSnT073i+v2LFJFhwKNxuDna3Tob2kb1od6wwCkHd5s4WWt7O+f8f
i2JHJPTtOhmnt88Gs/28t7bagsdY9Eg+R5Pn0hu0l2k4giAgGwCyZd2HWWIQe43uY2nu1DWVIr4Q
4MOCSUK7Mv8iv0tMkWbD/y4LshvLv4wd1RpijXrfhFonV5daK133lNQXRNV/snYJfpZtKhghZpgF
m8UC3zuE8CdZoyTycpRppSWKMoE2PWCCzKSENFe0Qn26ZUF7BTdLEcly1WbcmwWKGBxqNpdTsrdR
retTm4v6g21ldJkAivL0kUiTuB5lhKJqD+CKkcFl4Nm5DPRbecJNpt/sHlOgk4Tv+xnJkREKX7Pz
IxFsoTTfmAzlB05vWJDLtE/EFNQ9iPtKtgMNQWEnx12WDClylNGF1jJpi67djei8G47nfzymuooX
VIyONGzSBNVHEbBbI54SWu3JKwB9TOP1rQI4fnInuL8PX3FL7sZfLz5YZnKhLL5nvwydf9enYYGZ
r3c5ZXRZ3ZyrdEL/F8KWHgUEtfG854lQjDj16nJpidiK/gr5R9TJhT5ud4Tdm0Im3hPBB9EdyT2L
AXS8u6fMQaitlELIhZwd6Kbe9zI0lNpkqhlARiHYxTY3FevRL5x5AHacVmih4/tPO5HgIQ829il8
FuUTP5HMoG+JF0/nJRu3rzfAmrok+qixBUnft7oeL5y4bY89DVjh0u8j0MKTVi8NjCMEbUr3aNYh
hYUeURLTbCTv20+jANBK766tJWQhx2nPpjmcl5ytWseEpnIhC0END+MqVsLWrYllGAZuwhPyw1E8
eVcXwCOyg5jfQSfHchyE4dxohLDel4jpEJiQ+kmZXo/p1jOOWh+vlsC4Y1toHSYAffCm2Zc8qKP0
Au6mQGFeCfIz2TAHE23kZZvwmgVcdVCWxQoRmGufe3CMRdtTVxI3iWOxlAR9HeX4S7KJj1OTD0XX
ZF/JwayB8DZxZT1PndLGTtgo6cXDRC6rFyq+yg4Wg3+uGTc3HFygXXB+xB38oMa0yyQ3t5gpC6qj
HohVH4a30b8kuNHAWBBgz/q9yc5mokNF4XzkwPFlYdy14xOvS7oxbqmJfRmndmQghOvzlLi0jHns
UQDasveaF2e+WpNcShkNM94rfZHxA3/+DNtB1ZtrLg7Cl4qY/VJgT8PO7prAs9vzOY3+TGN2U6qg
8Ey95me039ufkZ335fCdPlWC7IBLSRqZJNesjtm2/uMqLlpHDrhRYCAauEcqdlRCwOlQ4T8kLY4C
oL55qcxnWdPIS61qZ3RTyMQuaK+zCAir+mFEId+6IVU2meR4BR6xw34wLz82fNAi7MsnAFTQf7Lu
BDM9AMZoNFyhXoI4NvmbfjI+hRvhrAWf+HFmNL0B6PkKijjuUT5Fs6qbfbXUYcuSm4WefIDBgZyp
W86TGBlutBlpnx+sbnRRZJNJxTTkAptM7eyryZvUnnu+QToWm4ZU6AtNUacqcg9RMrYFH2utKnJ4
/fqoBAXkW2t06oYi3SCHAUwtQZby5i795QBHkGTSq92BNU1FQ8IiI6G9xVIxRNvt9W02/2heacoC
eV5Fgz5WKeGh5OpMDI+X7TzJbcgomGzTeXIM59JMd0VsB62P2SKyImzfdZp+9dtEjx6IfWzAoUAt
fCl5dzIjk1lHueoN6n7B8o5OCrY14EMmC6aRmUFucGEEVYzJFiBB4X08QHNUsLhiInfnkZlKDM4K
BeqCB0ymnM5zXo4yFpkJOiQnqIdNnbul5AwAx6kgHhDTswpnO74+3H+MHGI7qAup+k+WKKahPY+B
E+MNNoiCwCMrtIx9I8DN8Wpe2JYcc3cD8SibsOneEib/42uTe1NZMvu668ZSxTemgQiWS0l2Qqx3
93VWuC9QnW3KilIznBsFH0Yknk/L+9zjLBmOl+14CNkQ8u8ILpcC8FDjCik0KrlO/nhO8Gwh8H51
hTGSq8kLhHYN1SxpvZ7Q3Adi7fv1/70e9NITwgvskflhQyc8bAf8K3n7X6/tcH7QvLd3+bU3Czg+
lYPC+4ipM/rmwJ9DPBV4QzW9MKpB4vEAFC8N7/aR1PBZG9eyt12E+PvxxB0psfDdEX0WKBpFYMWX
6a3c5rlwlR86R7wP1zh3jf2dTctzRsV7TxUgzrCTNGly9IqYTbmiJMQnLKltmakklH9H3Z/v7E1T
Jn/gsWVG746oDgEZdDN8Xu04yWKXDZYpUwqGYQQoYfHK7BR2OL9Hork4tS/aGq3Q4SJgB3fu9bjF
xazYsdy1nH8+T50M0X15o3DN02qoKcmDOzOzt4B/VWtjwdw0abdGdpl/m6cp1XLwnjKXnvJGZ6KM
8Tcv7yc51BD2sWC56IXXEdc03cSdrVFZkDY2mWvhxLMPjKTSPDAzsPbMDftWer8A370i0RuGf+xq
XPQ809LF18MCql+u7wfz3EzFX3U3IbXYbQNqsTJnl3gXb9kAmoYn2eTg6Q11zno4EWP8Nb6Y2jO3
aQWzP3s2mnbB1YJdZBTtQDvvX/xmEsUK9X7s0VaK+MqOlPQsTw1QFnFBbO2+JXMYdA2Z6P6u/NJw
2l0hukioi1bxxwJUjVEz4zM4SycwPP3Nx6HOuJ9y91Kv5FcsM30SJ14/q71WcJjEdr2cOj7jE03+
fg5HvyRbdZNT9FeeWbkS3iE2y5bPOzR22VYMNwZ9QuXhf4jv6mmQDdccc+GFnFT3AgTKYToOXYEp
Je05ofKHzEh9YvW7GiTDKQJpggoa0Fi49ldMCiWtDzRNM9hfhXJszWvkBlYaywctjU4/3EUfSJeY
ugh7ix2k9B4c+inUXwlqulgKq6kI3ZwKeXFREZ5X/lddba4f7dMpn2jKgyijYIOHrdk72/qin3f6
t/PRr9besL3oo9pt8ADoV6JhRtIB9eyiscSldJGRjYweVihShPB5PbGOCSjcqstoMpUMZRIbrHPh
i5h7ZMu60hnnsEZ4e2qhv8ApnSHPpp1uU6bhpIHpVfMVVLOdg/Rg5PEOKy8LIZKqFiR30DZVptJF
vg52/MYPWp+j7WD6jFiZtIcHDzawWsl7UwoR5GpjKBbmaKVjB/it+3gokQmx80Cxgt1WICWXZ6hM
ymccrLygQLrSWmmkU9tK5/BuIGcsbjmWAKU+L7fLjGEhsfdW42hc9tGDPT3UXuwlefrmFlgg3qTm
K9jwP25ezFKWLfa/03XlKrrKj9e5yyaigBb0ivEZLSIZjgEWs9X5YR/knt9A5qcxC45aQPRjMg5A
GzsTe5l/rtMyL36xBhejMllxeISeQhwfnO8g/j5l9qQuUXjtyCwhgT8Tud2jsDqsVjNMZFtvbHed
yeUNMiUVj/fbRVmV995I1Pyah4ixtp3LKWCf9LkFxZII24veMrzYjtYZ+Ap1Ulq5RE94H5qKuAqt
7FSMfBT7WeUfD67/cPKyN11Z9LEqv5KcAA/gmRXStNNTnhxv3/4qVyR2YXALIBquK4Jvn3HYQwey
5d8CEp2oGfMIZ9maPfksRZi1XdQcRi7wqsBYJEFLNjPmZ/UpnOJA6QPx6qVh/XduEWWDkE/0n/yc
fsFA40HYChqqsyCANfYysV6QJjoIgXWoDhO+KU91wQ6I0eQMoFoZeWfwzEtI0LZhsMkZWAO4Mpuz
ZCY+YQGqw8heyEtJ7cKbwCvKhaNdUlRL+IlX8mc7RqliVM0t7TnkAjPGzlQ/XghdPQHpMQ2bsnpy
fHZYJUaI2SfLKYuszraPESQon2/XiBZsmR3dmmI1XHO6YNBF7aTi+yzabkK6Xjj7UlZqxVgJFyO6
tK4nRql8J2Si0NMpNbIWBE7L22AI3Rr9kdCmcoH/v/7JCfRAIi0mHI01wTwldDrV88CZ9f+v+nKj
3VFhucEuyBI/I6Pa/n+2T3rzqf5nLIvoz6jwn75VQS8OGQd8BVYx9yEd06cRnsRxdBTl/88qqJ2b
OnWaOmuL36o//IVGsymsEkgl6K0MVM1uuxSCaou7MLhB5qWZE9Vcly6jtd8BCSoSPuuFAWzbtEzO
+FXwCqADY2a7z1wP2r5FjWXeT3VWazJFi4PGdkkJIfbxiSnjgAD8ffL9pybkvXpuO1s6nlCQPpsL
YLSUggJrV9BjtFVRcEpFPMuuPjkpx9xB2vJ5aJwu41cjQu3TtUzzA9Udih5q4Hr2mAgyRg2+bDib
6mIxrxeuq4bSX7izkpEco9rosfSQvAUrboPJSrHakI1kgG5hOwqF4YJPFC44yLUwV/6eYqlOM097
duRNQO5rowj6mwNAgBboRv8CtCGmDCckMFa+m1ujgMHoUZL4wlMGph0IFMD3HvZ8hk/CHuToEAzT
i+oAk6Xnc7qNuzyrqVhvjJcndImF4jpT+HGhj+NFHia6fY7J74ebhnLyvak1WmvUbVvNdFOGmcPH
2ZrxrCxd1tdMUoW8+TKIoFV5/k/Xdjc5gYgIjPS5lEG9V4yKjXfA1XqkJ+KEOAeJItM8zl9ns+ew
beNyp9Fa1E3WY+pE4pg2DMEhWVW3M9lo58jOXzWDTL+enIiKt5oE/qtX23qAalCh1kRPrkmzppA0
XZ63tG1nfBr75vzsiZT7T+/GAdYFj4/GhhnekWONCtUEbU1XI+TKvegnT6OeDFiBMZsec3xZ0Drz
lKfgZhaw3CXDscDyKiMlJ7Pz/YUEgPTu8XWw5/UTvOunUpEsON3nR5QHYtwIXcRD5LBnUeu78XE4
ofW491QdChT1U8npogDgAUsz60v9nWEA8Iz7YmYK3mcI2QYTa4u1JuUaTAE5a9jxFqXcRyjJ6VzZ
CXhKc5IvpBVhXWAED5pu3pjpewZeZjeHFQQHBWTe05uq39uZb0YO5kLpCkW2duumiFX5UQRNuMyE
yi+88ZdqUMkHZLhHao+GZZOu7/hbMAOLP2SXNCWiHvsg4RLrUaWbhXDjLHhqYknle0qyr6ixlg0g
//eF7Sl8MGt1j80NkQc+ym1Vorgn7VgV7JfNjQClXnd/st1GhCRZqScoyM0x/Lb+cdJkyUNcuhi3
ljjH5tc/JUBqpCqLyEZNTBwV+izCQRus0aomUlM3ehfC2agqq3CD1CMUfA9rEhMz1sMdD+Y8YuMu
Q/fAOx9WNHZgrhAugjS35bRRjPUovimV7P6YSyAsmmHgLxpTnavbEl2k0ieVVvQwZ3O6l9v860rH
TBnZVDNMRYPg63Quv3sL0SyHJ8FHXeWxPDLweBrOmRm7pI8qJ3Lz6sNjx1/RUTmGZA4iVmKzrsOM
5onwTIMrM33zgGmJVeybHJI3BtBHSjq40cQYwy0gYAZD/xbVc+Flxq0Yxek/1/Xnw/AmhlsroPIG
qyc6ZJQeD9V3/blYhQOkgjH70ynqXKgMQRNtMq4XE1Ey4CaHguoFAabGEy4HQ67XPA01WjWq3cDz
9RslS4myl/HtvDobZ7Pp2dyNtAWjrB6suZCSitE22Q3Slu/+DAS2PFDqbkbWm4YvkpsffDC4hSmR
l9Qf482xHSS4hycfWxqugCSLzTq37t8SH4Xg9mGsd+ABCYfRel2P11h9PDzXkqgK+POR/geATkYc
BQBysPOdBpGLx1PeaqD8L3qMjDAn7Nuv6VRR4AWS4ck7wXo2F6u1W2OUn/nMVhRqOnSqPq2UX0te
I9PRI/MZ3xVdZNe2Lo5DwrVUGnDgYIjVIhxSaUxvmVSrwG4bp1Dd9R2s4oYL+UE8JHJKUdE66/GG
rpyijO/EHSFlnaDrQ8eQN3HhAr+3HH/RuQ/YilvpC4b14Qm/C7KfhtNtKKtRCapSgLDdmMVGkQm+
/Ure45rB6RbrxIFVrc/OaAJQwFuGz8TM5zaMaITdswEdDAz2OO2X+mxXfh7vZQRBK2Xv53SkhLMW
I2VEussbjBRJu2FXlJKH+LV+saVSzDcxx2nx70K9Eo83vBLHGKbwZ4De+puGVTaWcXgH40/WKwDE
B19fTSj3uwwnYlg3P4R00FxP6xpWAXKKJOZfr0ASj0N0pWqHcWf8NsQofOAyedAaqOjl/64rGPd8
e36Xb5dFfg/RK7BjeH0KuiDhMK+Da69zkY/vfINYi3Y289BJb0NX5B0oqlpu/NHutN28Fuo4JvLi
j4eaXPnO55WmhKpDYTZsIy7sjSucQG0elL7AcEE9k3PdsYLaNIGl3t7DYsfdEobVQR08LQdwSe57
KUCmqoOqTYpq3KVIUYgcwPiXDCxC+PPKkpxeshaSXAT+LjpHbcudxQ1CqT+mj3wEiSdWLyHF+b7l
VStHCuOtVRjLKL954rUtBdPyxaadd5VIMH/VDBE94qKAm1xTaifZSJ2uF5X5pwc6r7IL6A5qd9uB
dzrfnBL2tRHVOj5eqWbu5JwinsKdusVw08yYepeWB9IBVvXbPdwIlC4k38E9MfT1b8vTd6/s+Uhi
jI51ZjcizuqfeJi9smIRKn3iZs+kQQkohPp7ec2eJ0K3/ziDHUOq1n5Q+m+4/MBWITjn8+8h8msd
z/+jYlWs5QcUSFTOY8ObzUkcCdN8761b/8vcdU9u1lOcSYlEB49eFmizperzOOXx97KAd1t3kigS
MlMQBScetspy1gIDBfn1pcnP3+pq3AjqalEb/gLDXPxsAmesMMvnBlPXeJBekbYdaqCoPYxFQ6uQ
PD7dFhQ6x+P3TEpr+MuUv9C5O0WU5jPXHqTEJyStyX2bnVar6B5zH5/+Ua0WeI+O+8r8OAqmAePo
B2CBTz4/wrS1vcNaqj+AaSl34b6xQ70ND0gpD9sU7q/OTzVwj1n8SJLzCuqTRr/UL6l0jbeIQICV
My+nJ8ezdmE5aakpY5cyWJRjgGdX2LZmvpfbP0q2vsoFN0s+Ji6WgUBmX+6DtP1onhL1Z39PwvCt
A6ThhoA7/7cc7bxOnrtC/kNLm1J32UWJy+7Lw7V+uN1RFOZNI0FFZGDW+4ci04d4x24ChMnclNy6
K4Zj8G9PTs508sqINGaYdYQH7VpBfpIEU0VvHSUAvzkVYBkRGp4x/bS3Z+KtlEsXM7AcSLbeWkhj
T6aeStLwMsTv1KgbNrjiyWhKD7GWkYca7hiAh3XgYMjdP0SPbtdtVubje09dUR+A+wTFJDowe9uV
Equ14XTj6XocOkNXVUUmB1d8dtyPpIYSQcXGBSwW0WZqV98ruvEL8+u9vBGorhzZoCtAxPWR9s7C
OIr+7Uvk70tQ5bQ/mqQ3uCxb2D52/Msw0AnO1eS07nJX1i1ulGLduYwYbKC4ilXCgajCR2Po8PQj
gJK13Sj65ymJE+lo9b/B/UDCqLsqi57WX5hgYlQK5+C+WrAv1MDvtZmOyo/NHWsoxsxC/dSHLPLp
ZHkiK7d4+7Ds6Axo1bWc+QIS1/Kf9k8CamnDj3eJqL5V/ma8fgv0TtNT6Zc+3buFk9zKGW5aHDI5
L7mJ7zN72qQY3ngp5WvjCcCm2/M36c9iXca8fYzel0sRYGvWSZ1mEKpyGcziyiSo6+qLiX6UGVHk
qon5FL9ejWWRm8qdLUvfHcSuTa+Uf8AdTdpzn1qcSkBpKN7YRNkaSJDPth955pHQATZ49hLf9bn9
RVVMKNLjtTHD7OjFCMQuowACVsK9TCc3xtWfwdd3fikLOrFx8MUN9gzcGDAem8pdk0ouHmqhn9bl
22yWATizjfp+08kg5ju9d6BWgLVgMxrGn05TcLclDO3IQyqNUrReu7Qya/U0P1k4WZZk60Tvjn3r
Q/DWYyaPfjLvbO5XqggNzzNcVlk/3HwyKppY+2HUZrXfkzR/ryBZUT4heuU7luusEtkYfgVo+HLj
1vtCke9cUJRzAvUvA9r1sqJm3piI9cK3gzrdUcfJogUfKUP6Do+O0HMft2TGkGjWFlhvOyowJSUk
KdsF7uP0Oh3AazXeHgv2TTJi8O5TOlvNrM1DMG8QtmhGTxqap2djB9kJmCROztkJ6dRZ4H684kAw
5cwyP89tqCYHTjlStCtGaQ9pgped49wp23bONyec5hZVdH52CoMwuhycPcAyI4FxnMSNYVWqsBbY
8rA65ODMRR5at2q0FgY4+KY+FEVnEPRfOYq7gRt/C78O+3jnwEr/FG6ZnNhEoDH3sqAHCDX/TVZ7
L/dWE7TeZEGAIdyWiSujRDSeV+fOPJdKMAievqoA3XVrPgnqEsxFbBQzfEAiTlFxcvOUAuX6fGjt
rUvYCYPGOrrZ+DZPTMnLk7tXWKBCXkC7cBY/hnRoDhfVxgTSl1x9jsKHeb/dVGZN6jBCVv4ieTCR
7XWha1O7UFdATVomKaKj2+sJPHfvaH1ca9sGCUSKRIa03XEyPX1VydWMzcVJ9SmRg1RxDABp04Vp
cNiazx1h2jbIvdnpevd8CTuryN/s6/SfiURyugavtIx37eXVhtdAL+onCql9OI/3oHLcfeRmGvVh
tkDR5wQRFtTRK7IKei7WPfvdb5PZuGSbNVB4V6CBLXwEx3d02ZItW49InkV/kfKr7f/lsrirpL8F
qbAqz2NUZEF7tF7rX8K7A08LbZHwO5PIXnAnwZdmoq7SP58RbZMfFthWP1AZ8dyLFNfivZqNT3mH
h/XX9aL+bo/BcboHZ5/SIudKL1xmELEzgCc3VlQgywE/enEjuKWimnPTaRCTOgP0q8024FB0jHTK
Pq4TWeiJ1jZ9Kt18HYf6dPE3AgnbxtRKalIdiD18+rUdhV4HHzKVUS4cKCrguak1R3h/ZY0tZxZg
vavleoTMPF9uwJmCiwpJV+lMPwN0WXNEfss0kBn0zkYz6H27xCMMV0+OqYSWBhcbr9ajBRgxYzm9
p7N4zzRzvZRlc9uydFcoDj/GMYiRnuArl4SG5GMlEGWDmeeQZOItPVx281oVHKpfpbqib5zYSkbn
0YWhpITCwgZni5Gm61xnKSMh+ZOXzqlJFoe62G3CPyfuBK17jJojK/z4Rtbq9QjIMwpED14WIKjo
zah4LVz6Wa2MripHPG88v1k6l6b2zRTOWjpVJt/U3v/AB4za1leNvdUCD6VnVZEo39sf2SH6zmBG
JkJ6rAc2hIIqTEMd0wW6lxj3s4NNLaADQyAxNJJFWqVU+4+LtG36E+vbS/qCfHLV2hwErooCsplD
fx6PNwEkLf04t/C+0ujx0OFY2AWC51DiLS6hycPtsj6yFs3IK6Ih39nMVvxISca9SPJGtGzoMT3i
idAsbXLnmZVm4WX0zb84PAqt002oh6QIwI6/DXjIb9pUef3hT2QnoRe+7x+QyJ0co6aN59awY72A
OrFJHlyBirHpgoyPhMQ1P8RQ6vQPQY4WLaoh/CSXPKqtA697NNJuPNLTzRgtsaOWruN0ntt/WmS7
0pR/aLFegXzKIxOyKf4IEczDLRW/t1msQI8MpYbr+/IvK2L+9J7EHhtpfz8gTxZngOL6TxIQocX1
7zMN6iTmkU+l1Xx3KLqQnBu7HB9fIPPB0wKys8weX4jBAn4/lWRCnkyK+jzbBTNZj1W61BVN6ECr
Cwfugoe2OIIDiK8h6Qvxb+yaGtVIZyXpNiqjNdewL2uW68oKywoGHN9pSg8b62lhDjHbmASP0Qrn
V1XbD+vNzmweWsc274D8mLl0xJmLiS7A6kimHgPVncqO4YjFhkakMd62BhasrwZia9aWsa6irEFK
vyBwzt6O9t/vZncEpa5htL0Se9yck9ZxvuYs8twHGUlDyg8SlUk5CnlKqS3tKMVA9ve/NbIccuAn
miE3yyllqzPIoq5K5x+HME2hQUUqUzzSHF+uDEUzYOZFa1KfcDCpWLSz03xuyH+VYF+HjGwCxkE9
OnLSyDbxl7Cp9/qngngQb3tCj5+2XKur0QFWGTfEKvYkGd2jKHkgGWsyS9K42+yZaV+oFVEz0PsY
4r/qLIbQ7hrog5mja9zQXSW+L8vMh6vNjQguIdqJ3aqTp3jKp5Z7cL1V0Mnqu5EvIXQB81pgW1SK
HNn3Qh1l56AViQ1wD9//jUvhtsTvYpu3u66K/asARJbup680V43zGw9J7e04gQA8mxEgix4x+aZL
WE1cbfaNmu2LAghhqsBUZKv5B/kXGHpCe/In6YcCrDu6IWPE5iGMwbC2KtwATiMHGLIMoDUL1LEC
jKUKuupygzQRutJ1eamLie4E+/F2oPtYsaHtyKC38wh0+xYoj/lASM2QkJcCAFHKyJVtyjW92jS9
8MQxX2OwfT5J95nTaYUbzuiMHamuWluPIs3tFy3NjvDUwonK49b84TVJFHBkraz4xZBrB6ShJYGV
TooB7BHpc3Gw5gGtBpfRO4n+53L8ght8cdQaDZagxvdkNhCzI9d87A349Lvr01mjSoUJdDMDwj46
zRLrSAu6tDjwFlWzy5v9nnFunZQGU3Pun2OZIM8vpYcc/RsBZXWPk5otWcV+JNL7MtHLmaoH4cHL
AhFOYfD+ksldP2XtCKMGKAq8/+RTn6pf+jClgTpiXW6T6j+6P63FBbxcYoAkRxVWL6oLCIAT0hdx
EI3AOoS27/wPQ7o38dzfXkc5Le9/MXLaxCqmW+34nr7vBf7EpPPNhqU7hB+QnpHULn2wxnojZqdT
u70OFNzztCwDPZYNu/UCqqiL90KG1f5ZbtesPo0SoGhOAO21t2E29UvIkzc+OlVbt5w+eTl8b8Zf
bTCHlYAE1JsjLqtUf0eRyb3ROnFToMFeo8x1SOOdUrMKPHguaFX0UVUxEhFZsY3QPMRZsZfS6iEP
4v9V1T4KmbCTF72iNZbBrq/LwIfstlKwUnKdeEbsE729IIKlkFX+bI5FrT/mvbSu/E+2H/u1gfgD
dfmbqKMZW9Dd76lKOjV1tS+HoXbM2r38ki4f8FpDgOrxj3NTyf9F/NIMpIMaStRQ1vEE7mjjuGmh
euZv7FInDa+CdxE/mJYK8AkfOueymW4Okc0C6wUQz8PV4lmUY7DmNY/saTMnC/y5zme/uqApC4N/
jqstPQLOQN8LhGEy7pOqwk7Sk+bh6CEsv4rReN8v8ahKEM7aBOFSGI1FKQf2CVfb5WpmAUQzFFPD
4RnXeeua+Hy2Q9POusbhLdV7D+b3RJmRtkLOQ62KYLNUDiQSNHZXaWxoWcDgaKzgLR9PTfiau2zl
+My+FUFXbp4+HSwO0FVEiQdfi2w1e3d23OD8gCwOV7tVD/0hayTXhPDIvQwgFygwbJA/tQSMo6m+
lkeFf6VyQjXo3KYXvHosmNTOACKAOUbL7TJVRaWxKAto8YU/VwkyobVHd4TEW4rNvrTDO3Ao9H7C
Zd1XL14CLAlkI7PnQamNQdbD7srwRPo9F7DtXUah7Kew7pKG1PzeQWGTUjsZwx9IipAGXpFVTQ9v
1NZ3lvyFW89nJd9Rvy7ETEEotwusYiSiCLeerEt+I0G1+gcOfoGVgCxb7WtHu+tbHfZ0E5G2Itrs
pH9w1aosS3KSybQeHDsweb3/JWRHgkfeaQDKKzZrLnEpc4Ct2GjR5zpU0QqGaNjXjqeyIMvIb6p3
Ad3P4VTQCcJcZ21xkqBSsYcm7/5yjkFZgkyRS6xHe7Q4eROU+nCODfBG1voLzISs5LMvQ5RV+0xW
BuWde921bixExQsLr/eKGhFMofqFCQhuNX65NvI86LTdrKCFZ5JA1x2pS75b/X87J5AF3MIDQf2x
Fy0oJmXGpACdag1idcKJ2EmoPcARA5ivrME43S+xkbU1zyTFHYqIQv3ona05lnV/0iQkBgcFE6B2
q0WgCfdmGWF90NNLbGTlyBP0YoNEs86m/W5ZP269KsmQQ2LxS8li3gjEVPPWTGokrA1ueQ6AibtW
ATwDXZVQoGtpAuNk+juaOG7wdU3SBhzfa57PxkilSNzvx53SLWakuN5HduiM0+IgnEcEXDvb5ZQt
RZ4kMKBEQJZBRCH+Z2KekKdRwyOFpzfuU3RXSrtuaRuwBPIxPe7CkqpTQT1M3xdOyZguWPGiligg
xQi1+VoW4ANwf0L9ZTba/RJzVCQeGkqhM3SkdBwXkoYlPEB96nKHE2iW/BahHxaiRj2t6tkALVqg
btl1A8G/hevklzGmBpJViM15O2FHg3uhPS/LFLiOGCYVQGEscYU7RK4K/dmglhpSwLSF0AtyPeD1
9ldKrVLo6nz8U/4uSWItq5Bowtz3hZqz03OZ72oX+/xUom2n3n609IsOPhoG0wXbDUW+UYS8R6Eh
Nu4sldFYipcvgbHOUv/XAr/d0KAIW7Gga6LlTA3IOCIGAf9PlZbJfl4kz0G51zGZ2Ri6YBoeDbdB
OKz/hqAm1g+kEI9H0ZZyYEcF5UC3EeLG6Cy2q1Xs9PNqTQtXLsNeqt7hsNcQtZDyMDFSkCF2+xMT
qyl/OTqkXVxF7sjzz7kHokdl/oeYTK/D5r0H9v/quJIo0bR4v8SBqGg3V4Fp37LqAEUZxz9VTjqq
hK1xukarjFPRh6Q0JHQJi9KzadVHjr2Wi8yLNZAtVbfX/6COdV/LoT4D7IDelTDlyWCIsOUPezjx
WxFftAznUk2OiAQpqdIxms/5jhwsCCMAz6jQqoKoOYAynemxDcDkecJQpqWEhpfuFLBry1Zt0dov
NTXxm1dYx/XyktrxUP3SqQXMCShDSxAyhZLASZuQA+AHWRuI8mqAhmzzmzyFEE/Ip6PtjOUjUjso
NaoP82AQKz3Yj7o5dIwpBiGOs110vrNm+kfYwZh4506IHgOONpXznEGy51Tb77b0dOf7dIGGKW+N
CEPSAGv1J0qg7vEpTBC2yzZyc/UAiNSDiuwFO/bS34Edxf81SFgxLTTnOhkdS6EaWb/lh8v4avIL
MDCRXyUYSa9ATwjANFyKDeYl4FG2OBlLkKuS51zfs+kCaNE7xV3jHXclrkv4dSCY5D4/GWN9PvAn
vjyIQheMhNlhyOZv1cTnewlwiMk4USMepIIDUhtdCMJu2m0eAYhF+p3sbCOpOFEFv/VG6vqHgJXZ
Ehwb7537NHlPGMAhOKsjEZVdhzKfgAhEJAvrXEGoujG/Ykq2HqhSZcsRcZcaZsXsuL8C+5qcQTw0
HEHb0cVntNq5QWVIpPb4szvYQzXLzSeAAF8hE4eF1OXL8PTkS19V9sdNZ+9u2RmPidvz1h8GucvI
0rz0LEL3RNqKooGiJ5MpGwSVMcMEBXY+Eb+TocbnfkbJhBhMLBZS/TF4tzbW1J+wvhclYbisbhUQ
Rr59HMvei3X+jwdstrZxx6apL30vHmCUObMRsIsyg9qDn+p2KtTOU9j2tW6IF7MsXwWOMGXPR7dX
FJzRAJKwOBbUk3X9mTzStL+KnwIhB4jxUPXJfEY2ReWtza95a7TQ2BIw8XrNQOhELqAu8SMKdL+N
4VtkI3AKxWL2mctSOyrm8CUXaCUUgeeC/ZGDSX8d3Lh6nuefFXN/+xlJLwxD+TJuCQ+l3AmSVU0e
J4lWlxDi3JnZU/9i9+F3uf0rziM34zZYw5ciJ+qGNHUhTHUImL5E/r+ei7PP5Oxm9GmJom6uaxEv
AE5xu91oL2EXVqLi7U5z305er0mIz/AWrUaLZ4hFlG2Ik23OYN3Fc1yVuG7tQ8bsCHJHr0BvYeWi
Td4+JMEG+LduyXBx39z7Qc2CF1vP6fKUUEVthVFhtx4/whayWgT7i/8nZdsuCMCVugjP7dndXGcF
S9Nc3ka89orOyqZTxsYAqmIPH40+Ve9PJ+JoTzPWMjlWIKo0PjicdbNGscnfKbNHJ6mfb82vESD5
hlHHBTYq6wMLeE7e4BcstZRlg3ZhVi3TH1uOsBPLw93PdIcaFYiUBzbsRLO34ANh4B3nKGqS9JbU
ribZeHk0VlkxVgCc54leVMjivR0L9hnd14UnX7IN8kXhXYU5hIG9uv/cnTP9SSt0jXSZwoPVJkK3
S69qJYKb7dlJKKXBagIWnbeCgvKREbcxMs55civc9HjHAGFUX7/Wphlfmsdlfx3E1adbFZDuwEDC
wk3IsuZlXUPQq8c3kr5cIQdBulQHlTAmrhmFqtcPK/cqif/nUQwUdFyIhcVCP1v0kycLrwAk11wk
hwScSZmHTfP6hqH/wRvG2MB3aCfy4ddFKFc2zDb0z++JWJZdDB+T/FFD9f1A/mRoN0ISEfmiUM90
FtKuwVfh41Hv0lamFb2GlGY3DefPMwRsxBbUcnGgCJDzFcwg9XUkvv75vXZvlqoe9cKbFpZc+BmA
4zOr7kVLv9s+AOkNz2gi1jLhsVJ+KGVzrcR7NYU2jSPSl2ary3uchGCwSWnY4AqiWYSLt3CiIDKa
MvCbjamTNL379SLm5XQKon1saualTM/JuqRo90kuipRbOGwC051qTu0OJrTpurKDVpfK2G51BIY3
WN88rAV94BVb8J0sB9W7rpcOOMuesN+NPs1WMprjbVu3IhV0bNkMf5nB4DcYj259AZnlmtWv8wvC
xSoTc1ILNDrF4r4md4zA/tnnbsTJw8Dvo4dbQbqX0qc/aYqQpoJmt5udxgpsnHimcVN5oGRQvvAZ
8b6tOeIhE9JETmeAWCqX79sUdwuVY96W/Yubhi1dvXRkV3v4G1i17wEMes38M/+ZFujRsLHQvBI6
oT8jJrJNiJT1pnAnMvjkvauaEIJbi2UKBZCVJuxsE0/XHGZdxCQL1NtH6sSi5JACFxt5hhLnYehi
w7lKoDYXG5eRObrRrJCksAVaLINtQMOuR0w+NrkBtEyYBRaVcGSPHx8KzszJFD8e+sK6unRFHvBD
ZbLWEUdQ23O7NqRImxurYEyYSzCJ/O2J21dhV1OqZ8rXAk11h2ypl/XcwmGzv2XRx7nPLkuKKg/k
JLqCPPUca1GJ4PzxFgUnkqvi4Cm4tuFnnnYaQ9SoYG8taz/nqY4TwDCf9mwNBraadJ0aUSJkok1p
80ViLW4ZcuO/G7gXNJMV7jbqoFYqLjaoDY2DYDQuTI5B8jrsx2zxUFx2LjS9RLatPiH7xlBn5MWE
2WyVbRxHkjjsbrZvaYF8qFfFLipC35n7olvxMsX5YYH1wPQQCrPoS2HRpbKgiybtRj9UZBbnKlcf
yMu/+gbS8x3RrCoo7rMxvUGyYopoddfMGXL5X1Y6nFyHQ/EPqaxGtuC9q74HlzRZa7be+7TMwTC9
dyZCEFVSmFcfjTa12L6+k+oUwbptxfcYSY1TAkIlG6fafyvzUzPT2IgJnglevJksWGXOiS0p8C/+
yhg4/UZSeKy2PsGDcNalbX9XVn5kGvo4jZ/XdnVB2Fov6qSZGW/9k0Du61+f8wXJr/o5lKsCSd+o
s/I737tOewFKJV50suq8ys+5Rn+APPphmLssIiICRnuuU+dKni4uNfp5kifjvR4WIKR5FFcZupwG
X1fxW4xFVXkuYKhgw2azQK/uFS7xJPY+MH2Zx1MaR0cjQK/nlHpQ4tWL6AseVvO5VvGVAf7kbS8S
YquEP8H46jw3YHm4W299iSRMm92RvPb7bd7aHlXxAjXCOqWBfKOFelJKX+zCXJg66qsleGPqMK/U
bXc8z0RyP4jxYOBRACEie2eav0sAYCz6tPwN6O+bT/VGJs2wUzJjeKLi8h0mA83WInZszx65oH8j
aYl7uR7l7GEMQziWchR3yjhkr7dr0Ex4QlG9p/6jAQ0uRKb3tsr4VRey0THUzziRDoJwlsfmsOLG
1tFWMoGjiToYUA9OXmPY4JkhRFdwE471fkpa04oYQL5ENKf3Ct7gBvJYLWkHr6MGIHZoOrMFYLKm
fh5E2bEvXVjhn06u5wJBdz+hsGkszN6gvi7gKO18JOEpwQf+EaJkAcFhXZ9PIewwAwPacAlZs8PC
niC15Ym0ldrL5DB1sJkorDoLEOkVkNfn80KPG6uFBPvB4mlxr14Yc1EfhGzmP7L+tLBsUsRFZmeX
5M6smDxCv1XtDIXuQQ75cjO6QeBiH1HRDmXjAo8kvfzx4E4GKtDCEEMUjWYINFJsT5ANc/S9byK8
lHC4053rIxdA6pnYVW2BS9PG+3hUJA+BVTlIb1eQfdS3QCpxn9W4efPaAVG6rTNl/NoftVhW5qcD
oiVP+1WwY/rdbVg5TWsNNjiCzdB7d1NDx4UeQUxrVwhsFXSm3yPZhASCbbqLjyAU8FWLWAwSl4Xr
18LMn/gVxB01LcMHjtK1bd1zYPamPCdm1NowT+jF/yzQif26LvvdZ8G4rMmy5VYheoaG5YAPUxed
Ta3z/RYD5QK8QbLLYs1a0s9dy/gf8/GTX2BGcra6RPJuVylYO3vrV9T72TtuxxMsqxkGBOxS2m6u
1C+uLlEz7VfIHNI84x+kLtpqtx9VT8SQ8hxMnjtLi8KflJ77NXYcJdfHTy8K4QNkwY3lR2JXvlWr
ASVgsEsSAEVeeqai2GLrSNvpWccM5Vb+pBahkWJrZyoUR4+wlNHjO8Ln7p6KgF7nCraBPkAziKlL
XEdOKWiio6KzrNCOWB1L4cz/LFhcnRyLaXgNmp1k4wmNDtk9iF7OhH9SknlJOAOm0AG20UboKmD4
FEvkPFwHuGnQrqbJ/p+Rkq+F5MtsS4GsUy6luKmCcvWvws+s5qQsY0Or0qwmSSQkwQCfBHKc8NLW
ts5S/qTVRw9NRyahBsqVuVsMTW5Ch+DORWb8ZBafiJl/e+W41qfTOM5B8n6NYp5d3QjWnz8+wQxd
9vlbbg9FJydS+WyYs1his74WTMtNxLGV6Z7IuGp0UEbXrGy7lPr68dK04+PfxV198ZrMtVzPwhbN
kJAYgOR7MDj9SOSDYLUxbWf/J4erawyUlxxa7A/bj4ApbrvEKTEomG3upM49uzFMgS+FEthsQ+EX
VdO4SO0IkPAqJOjsCGdGsU5TSqlJY1ZTMSMgjxQSkUtIxjX+YkoWluuc1z6RMM0Tk8dFyUDwEQTk
9DZkvRNyKUz6O7aiiyR3r3AN8ax2pdCXLccfbxl2THXDsse+SURekYloRyVxLZObELFWRN1o3rbY
FwPNfL0PWph/+IKRwMes7Bki7XfFBnJ3hXeMfGGRUNX3aJj6lrwZ1ls2dFccfbioGuhKnu+o1/DC
gFmj8LBtbpUf/5oYjy3w5zSF4FC+MJgYAQptCS/Tk5uzA2wD/GFuFAiU8/8SkLrhgYHF8CuMdR4y
5OgE9bnJLAyXGEQj2iEg3XxIX7UadgdFVecMn0l0U/ZxiOcmtUBzAFXRRtKJSri9cow6092MP9FG
NXwpK8in+CxBY69qKmaYjcfGMK0a/9M3IeHcPLqAbPeHlD2Y65zaKcYcf/nDmf6/breM01ZYvfub
1mSs2ukWivSONnWH6hyPNZFvpPFBVHZZsVyIsADHw9BsM2A3/lugszCCmPwi06urfDMPzj28WnHZ
Lz2qVYtNE7ADz/ivZvtqsXk/i4AZiBUY213cZKIbxAfU9Hv4+uZFbvfMjWPVLvbLrQWt9PMGfVUy
zXGChRic7NttgEx7fKbb1RIXpLYMxrtR4+L+iEIFawNRdkrXscdYhJhYTn8OzOgJecgLA0OOBW45
fuzzTGgOfQkzm03cQcb1hHJ55XG3dLEW9GvVhK54YT3I7Y81IagCYj3NBSachQo+caiIUDLtjHn0
46Vv4gs9wNYvY+hUtvmM9LsoRruJnc4mNTuZhmZZBzjFMpmwJcRmDbP4F6PNohldrKnkYrnDUOOV
SMsIdOpNmgm1ZBM/5MiqKGDt0o9XlWbMhdnDNUl6ZVT80vSwhFGH6pqaNq3169QkikZbavPYPXPW
GDatEVwzZ+3hMFeyp6hibxy/kMao0dqGGIbdjSfJ8Prl7WkqpchfXJMiWdO7FGcxxf7Xgs74HbiK
VfWhrVMq6utjmnC/wnpLBZ7JH/aJzoT/Xq3yVXtO+z1UTZE5FPg5vhfr8HQrev5vnoPhbe6vJMU9
tv4bGK84BE/ozCJbMWcXpzuBqliwEisc9/RsecgTNSDMN77ytu34ZUl8cIdzFztcQ8Hnw1o+TD3W
XEZ5ffze1YRz5qx2u/AMsq13WBgE9bURKshGmxzIYAb8SQkyy0Wuh0iMlq0or4yISoSJRKsNGqW7
ufzXzsqkxIdmmwghDCOsqgZPZE8qYmZil+vRD1RMEze8wvD4wNED9DEB6J5poRaShsvgAkWoUsVT
oLJow/X+2MhMmD8YZVRqgZKU205aA0r8T4ayjGs0LXILMkYt96YrlMcswPS6Ns2PFYbkpfyL58s+
jOMFKzWppNW6WfeFAlG1OLvVjvXOdEsKjeXE63CglM3DkhjbD6GInwgd6XPZ4rVcrAns5ULCc7W6
klPbt7tcLy+c8RHeTkIjBM6mOZgS0ei/3g7x6niZklOgLQWq/4nKNtNozSesJnbtiHCi8UJ7Ann3
bNzHPhaoc1xsLFv6pL4MbD6wjIpv8HVvb0CdWlt3gp/r38IZ8xp/y7LPpMcRvQLhwWRVc+SmDWFl
VsP953LPyUtMoeqccsbTx8/VGi5jEsgZmxd+dySyXNoGVmSrSja/A7mJtvKTLBKekalNBIX1z/VX
CXLuUyfgcSD558u/2trB8+BM7nlEh2lrhM3U6sXGeVcpBT/QA4Ubtsr4H73Yo+RxwTeusWHbGRS4
SRiqwjIEfG+SOcg0uKSepFT9Fa3MOhqCnZoCxOOcac60pDdMlQ/KAPzUS7tf2YSadXAOg2PNeC/7
gUvP1Fv03JeodAIwhBi4mnzzziGw5errYqcq+7KUEckEWsjZNrcSRHz+SM32C0Cihvk8liZcpACY
o1RzEUlQieuaBquPsbISigSfMZVlQGPbKVyFpFrZF29/oeV4rc/kp60QWuOUFFHBchugVP/EZprs
55d5L1dFtpANz+pEsaJ3DmrOb9cd+YVP3xJGSuG/LFPVUCl6zQ3CwBLzkjMTreG+gFWlPZv3hPOM
D92B9GZD2lsIqPMpMtRWHHHWUuLXJUj2OrDr/hJtm7+L+xN5bjI5P6nzr5aYmlzSw9O/Kwz7CqhL
bKxTF66X7f+YjREh3TruPVI6uvjNGUGF3MiiYTnDijSSPKR4evZACa7qqdnm01sMes7SQOMsXg/x
hYBYS9OYvFYmVxdo0e5Hz0vJ7aofMioeGyWzUuzV5kcfJZgLzFg3tgog0fkA/RCaspg5hLVpCyKj
bhramnby8aYzJe4XPnVzPW2CFzJmA6Zgsm5AU1VwbUvUlXOMLyxsWYFGYAfW5BLRnFMpxKPJyDa4
VuemCDNJ+tknxGMJp8cHcDrt2l50wG95tn+A4POmgU3r1Ffqedya4XsFfyTuhzPGy7XHS0DiWO35
cRRxFrYH7PfgHmSdAIKKfVRNdGxHrkQgz41Kdr+2YpR2Y1V1fjWMBSOQLCOq0onKaNqVHRzIyuhm
WPMSi0xeckuHR9XXSg7+E56DTvEM3pjF2O1IYplGLNsgWUgEeVxQD1lLECtOMWVMTV1C4ahhABmE
J2O7zm8rDYKZHW/1Y62YcD01NRhQIzG27oDQ7e9cTxsQdfXE1StUT4jMnzB3OKesQNvPP6j22WUb
WQvfZMG/pekiLYMoWynZvc8oHqNJh8A4xckRdTvRN63gkf4zYbp2y1iu8YxP/RS2lCMIKVKfTQGL
pZd3yHX/2WQ1CaoTnLmQOjyg2XPPzD9QVXedU1RMWhLWpWezndLf+kWjpzhS04cADyjjkkbX1vwv
cxvzXGwhzkXi1YtaHohnyCIbG35y1u0M1EfsUEJKwNwAlmG0QccFkGVFopsrhqMmwHTioASgGnKg
T7EaYDM3PjQFtO5TuabamRr1kiQDy8C6PL/VP35VzB2uEkawgocklpesKOYJmor0IxNogmDFG/1W
xDksY1ILBgXzKfuJse1AtwsXKhgG4ig+d3053fL5dsnskSTZoW7hWrK4CAasdkf08ydJIBnt7oIL
V7yvB3eAM0qd6UtnfLLRTETNlylyONM2zmztHG+Tk95L0n/cStOA9ASe3p/Pv1OlTGf7N6WY+qYy
lizgU7QDSKTbUsEtvKxstV4ENk/XE8z8ZZR4Us7HhX5ItE0dqhg9OpYKH32kfyrY3Q/87swS1gB6
/rWLd3xxwF9ZsjJWokyc93N7eWwF/nSlHXRh0hVOfRbYsr/iy7ow6eNUw3SiqK94UXFqRPxqn9g4
z/eFoAXSPsmCoygJo4h6+HtmwxM2UTqCDY5O2TcV7e8rk3JhgL0SqOIKjRlMQaoGBsWQRYoVlMDD
sR/mew7+vie9K5wtjHZp7+QPzqGxKnkUjGMz3f650qhj89jsCFHuUtciuTT0WqJ66wzCU8uVci3m
ozGbriMcx0no72SRveM33aq62BFIrUFj9mQQ6zfsBqEENivU7BrTUVJQkZimYQf+AnVT56rNPe9O
9t4OQJDyIONUOe8Nwvmhh6hlzRP9bjZuBufHWkVoPN63xWECivo9UB9QBU2b2bv8nOdJm/uBNmX/
Mw253NBRGbwzTc/ssTOVW5i4rldt2ODeQXs2M8WpR/ssYlKKSXdXh/A7q67Kb4I6w4B68pKMjI5e
u7/lZM7eQoF3zC3CtA0qWZhwqb7GlZVhMBF79zXgtp00GoCajMS76d3Fglo3fi2vWn4MQKZdZKaD
lIpfZjb64nMJhFwVR+0SggD/Yn/a4o8wv1dxnIvjn19HcCADLvmREewez0FhXu92fm+am2DuZ0VA
hOwmPVqrIObykOWcT0dmXoxnIiRPYV/ERaWRFf30C/hQbSrhTMYlBWp8wef2OiaaB1z0JkCtNLP4
llWf1VyV2RjXDYEAm1n3pn3rkuojPp5/koT1x7YDqPeGOibJfQEKJEgdoZvHd0rwbtI8oWYehL3C
I9OlEVex5hhZrt3WAR+c/8rvRFRswZoBrX7NYxAouNXlp+EuY0QIegGaFQ9Q2eFt6gpDBZ/+5wQr
Rg0oSAUwS5DNCTYctrCjpqGFvyLkHQNIsZs4CBk41RoSlGQ5zuKZFo6ighxG6jL2Is1cXHKm16Yc
0jTEOn6C1B+HUBrKRl4dLX4NmsxWiMMKrzrWmxifF1ccIdnZj2TsAIjSylocIoEI4gvsoWf3NGab
j319WLMINgdahH+aWDikeLCRGa78eaLAktv2FYNdEp7GNfKHUoJc4TyEk27a6SXXnvZp8IfAHrpG
yYcSvRfoZjWCsriRvdYTB6LfI7YMC6Ib1uiefZ5ox6M2Bt6+/otgXn9kQwluaFG/vRP0brXFaZen
EXQxkPStIXfNAHLclnlDACqobWsZlWpsy2VzXsdWyOQMzCTXJnDSOn30/5CYPiVqsngueamV4zyi
zfvsugUSkLJ8ajdh4pH7ZW3HrUlQBIU6BL8fIZ8QqdWib6eiiBo1WkClGT3M9qwivPoqEEPbfT+s
4G8jthSRGTJGFASlBFqQaxU9FYC9SDJD3AC5TfxdxB7bgQ4pgiavR83yHJeHYN2D+cp/Hnsm/6Sd
6ZTDga+i8KXUAYCkb3qT2YgseN+rthCHzl9ZiU7V+JcSWm6M+Ao6BTfw9QcVfQsyyKhwHdyzPi1b
aCX+3H6oEHhVU2vy76j2XkbW4NJqk2Q75DFyn3SKKDrwWRWOZ/3LPcQ1wonKzR8NspHGdmRfuyHc
6Niqf82mkrnXNStzkCUr0olB5HumWPyxY/EGdXq13TWhl0vOkky+bSUlsCnihC0cvTSTt+dVLPK+
FbY+ZRvJb8YoJXsR6XgnjWWhTMqpoLK4nGetPPBVzaiciWyMG5AMifYlWUbpGj3e74HONSYqSjE0
CtNCOHTT/xbUbA7hY/KzZHXMyfTC3CSOrHgyKMO63csV19BQjoUgMNtOEeRtXd7a7opE+NIzvUav
eYQljzvfS/hHkulPk5bYI1Jswazhunv+EmtzCCCm3q9Wk+Gqp4d0QSTDvvDbTsim6Luq5yLH6ayH
6rVXIwAYg8VGjHAu5mCucfVq+w40YvZQ64Um6Fde2In36SG/80NXD5yHOSBuj2ACdOakGmx12dC0
Y/qVy4sY1y/ksPezGZ437JTRaJN+Rs0xySrwjvbtmtYc5PRdWbJD/sJmhioHURgkaScrno758XDk
5TWE/l9y4jm8KWKazTTi7l/DpLNMWSa/4McBUxnCHZ+mpwCDOD6RBVRPCAXGgsZrPzqKVHiBAvGz
6trws+TzlldxPof0C+3rcvnBm5swq9daM0/pVTsWrYJUiknzX7hOsZJ3tSv4fRXDA1QazyA+jyiT
W3jh5e1+pAqkFDme3v5lYdntukP1pgf5Szm1y37Xf1Zvd7wKqQB+LW+Cr1TsS/Q0wuR6v/kioF5J
BdCdas5gfD/40DrbRS/N3rsWQrw5BV4ukPR/mPu3h5jqmu0Jf3H2yBGhveVXuxU0qUlIpBN2U5lo
+vUA3IEoUhWx2if87vpv+oZH5XevPbvKEKk6RomJPhKjZHzmqkEDf978dN3s24h+gW7nf8s+Egst
T7jNVDR92G6OaM3GQtzKNO/UIi/DKM1YE3cFAb3sgDxlM+HsSfdRvylqy9UkGcMaeG8QsGCTVUFq
fSXpXHWfV8XKEQ0hUV5JXjXNzOSp5Rmeh+Hu6Phb8Uv/TuS2paFSS1Dfu+RC31fEy5lrZpAP3iaU
pra2i1VcEJJTEpci4yp5+W6ANPi/DfNoPeECdDME2LYGJg12WmJq4RoV0xkGMm5RoVec+VO9gcXM
n0jO7a/aD3WPP9C9X2Z/Sp5Bbgbt9HXLkml9BUfJCwh2Z+89k6NFtteIcbjsoJFjuZqgrpsIIbAC
0wR3FbRZTjNf49OGRGWr+vr3b9UpRac8W0FteOaaziEMq/NworE4HBsQ59FbHvtUUd3FjtAWTW0f
F3JTzowJK6liAxj8lvUStl05YoOLDddv1QKGsTurJN1DAnYS4+GkUEcZVihUo+5l4O9smMwJCJBQ
DnJvctZjkEX7Yrj/MaPBAXOOnXpWZ4V1Nlj6Lfcikabor0FyXAwcQH3BqjFg3XXpzcBl3lGdW5OK
zRsqLhkXHrpI+1jOIlv6lGvQnzlPhhFXFsTBpeC1URrd378dscCdq1yeA4UiijYFRNdOrDMFoZdb
qUp8F0bZgwb6Hfhm15rMrbkhdj4sYW2mvidMlv/I6g5DLTFm8bCEY7HGn/qdbn/OkuI3p+xe01kd
xEer6buVtIdDC6zXghR5TvnG4AqPxoLkI1K47cPE7TJeGAhOLYR/wZ8SiQBXz/+Vrhm9dz9yElLr
n2Y8bgSZeB0MNoEVJklJKQUa6gCIqOAOE0X22cdPuH1hYhThVaAfgo3AXm+BR6/DJ1Ijbp6iBjO3
Hcw1mqlE1TGJM0Lvmarwnwn+z/i9F6TKLAgY1o5tJfUKOJJLy3L6OCF94KqYmPFbHjla5bNgLWmU
UF+mhgifXiVhO6Gy4iHcDypjUiXNnFha2QSSaCYef2t3VWRnh0/2L9Hz9ErQIECwRj6O8B9zk2Cq
RlwjAtNQDsoNrT0FkaIMuFy/HrYQTsbFwxo9pxy+MESa2Sgq2pn/ooaRSUWHQE6Y3CTF3LOGDXZY
k8FprF8ToXGrcEo5yZ7OkYu3ayW4Xr9mjFAmLxJdUe4Jr5n4h3nEaRcyLKc7mmOLIGqfa7GcvxOZ
4AYFeKb0/WSk83PWVcZzKl4yMeWPnJJaYhuyr3Xh58oitfUuZg3iejKULdpm9JfO7SP4WQk77WK7
IqkUwh3mazXOXJxFTKn3xYwl8J8waHPIPv1TSnEbuE1WUMc2VpDs36mYIcZgWzNMZ+ytxMXm/owQ
VZLEcGYI5bVpQpHsQ1lnhEryo4BYnySGO0X3FLAoFUxPLIxFKldxlfvO1rfpgb10JEgaERlk0SeN
7sGu+eeUten9CmS8/E9RZ7T+3e0LNayOVYwTGQgFuysCF5A8kC3IDYr0ARmEt49kUzCXIDSwye+W
QUG9ZjGVtCpmTikmef5GUC8zhX3ik5VzKHjJoDdAc3i9UOlBa2NIfLVmeaV+hHqOaQ/OAIXPzX5q
bGHLV1o5f1U6ObMBd7lqekB5Usejuby58QaHtF9Ua4pz4gQvUbLpbdrgIvDUSofw/zlQ+/uZmhu7
sCOCN5CR9e58c89kiSkKd3PJWAETvVYWaxYOQSwV/DXCADYTv5opDg+szc0mry2KauYzI+jT2/2B
j9jOAtH60qbkvbpUS4Z5SHVJNxmGfGmRDG6mnaG3UWcnWETVnYWNbBoO/zrt1Micq/YvD3iXRsFo
0ZeYXq4bb8hwZGHd4hMxHrr457Hhv9WYYJxKkFcP1aeXGf3hhN6vSH6EAQdG8NGDd7V0Xm6wCTfw
1CLhz0EfuHHtdhKezcK5CDmfnSqMajCaY0NSL9qbIQF1sxhj9PTba6tTG/lS60xt0VonPuO0ThPh
w7Vg4RlaUnP1gMndrsj+zNgT6yqN8vEs/iSdKpOsOrSspvCM3rQPmd8ZOtiwnD+T+wOctLREhLeC
JuIVRbwvNQwyJlFVCLkYInP02GltC3z5DQ0W9G6WQSF0pJ3VlvJZc7qMlZFk38KHMowax9mxD2nU
SBbqVIXsO07/ImC7k7xtnOdUaFTl8a4g7gNiWQIJgDYY3C1eWLurfTTY3T1KWXfIw1o/vYJyzNGL
lAQkqtwRS28UqnxbHKc/AoCM5220WZkNM1e8Jf/9g+N+LZkPsLS1vwp9HQ99MWEky0M8zYQGhwpm
p6tnrBFR3FM1UT3SCL6d21FcLw/dov3yPGq1NrmpLlMDUoGKYbRBpokHKe3OGmVUvH+ADmhw0zYK
VY9X7/gnJ2/Iyu82YEp/B8zLe1mmaHffyJOayQufzBx4zjUgx7SkmOBJrcgbefn0sU3795AHcXPV
qT4tp80z13VWjVq+IVN1jbXluqoTvyPLoHAtwGMuFWJaCNES0PCakzZvLPcXGbmPXxzwtezHaZHp
Dl/u2H4/OBQR0Yyih5GuzMWqruEwql0QTDdSKcmtHeTIr1YS3hxNN6gdViFhF9X4IDg4zLPmwz7S
lsdTuR8g6I26100xs4UhegnEkXc0vuvkq+3woWjRAS8UXBWvWkHGfwIclX0koCuga76UYzK8+Wds
MBKx2FXpLUHH4gLJaom1RJ3SoK/mpki/TIlLo6mFveZ3klJcVvmmUF3u0wxHxYxmTnJTAcyx7Xoj
3c7uztevH8nr0Pg8ATknF4IM8KUA7Zd7u9oRmXQD2UBocVtwjLTjLYZePliAjfwMXjIFbluOH2zm
Qe4l+7scuavpW3xBWiAtFuNwGqySVMh5CIt+JeDmWGnbzfkfLvj+WxzqM7H99cp50UjLPBlIaDXQ
Hs3fRXzT5+blwry9lqwq+29GGuzWkPY+iKimdcKFVmdtw1Jlv1whqCK3Zm1EUE82aMZCbOBHXIqR
+sex8jeHDG+ZeISXy6uupSD4C8i1qx08iE1b91pongPxZv5jHKHS9BHzeUEK2roXEuic13GApXPS
OafOeixjQPwX8k8UXBqNqlA5yMbe51+RpqMxlWlsq4tbiIupAQ9yKFqYZZvX1uOx+PSNMS4tpV2O
ackVz9KKJPJwCab/qTnkjlXXlB7GmtSZOB+BoYt4LEQ6qGY/l13L3zljV2RaVYgseAI26R3Gc1SG
Ddja+D3AD7YpX697JYRjPhv7CZrhgHN/peADrhMen8Rbiyjma0yyCMckj9kROtSb6RSWLPetL3Ey
Yw7IhVGvJE7lRvcvQ7GYd3vfuKvmv6Rk44Oa6CMn9yvKp/vvfYygxQO3eEQdduM6GljzOA93CMxK
O3nyJGnw/7R2JqcNEN53Mz8qsaQEwo365NEEcxmDsL4BcmQSBrpAbrT3tYU/1M2apAYwre9ytc+G
4yMmEzKkkpyBc6o/Q9FbzohrMLVT/b3jz3K5pU/efHIbN8iFlPjmP4T/1Zrn0A/p+7Zc3UJ4BlGe
aY98A7hGwQ4jJl19kXe/PTwKepCeqVy0XCfmL+1bEW0Lq0D/VSKAuFmRNo28uWAI9upfJINDsBFl
wqsyhJvR4K29yNckLzxPbOofbz3Er5JDahNt/sazatiNPGFmqmnEZ7jIZTZEiaFzrJWQ07YoZjnr
FS/+PkcIuNwSMPQXn4QiaM8N4pDS0yF6bD3tCqDIPmDt9sPNzJJRnsiv+shVZQ/59HzJXNCDWDRL
xYoghUhm7bbiho4KXurt6gW9isJ5KQjfkqQDrh9uGxw+hoVBgqXMTubXNS8UozKys2GSYw2gar/C
yChCZzAow37oXhZOe71VIDDM2coLwStX6ozDUjBmXW5qYxbtnqxc7jgX1iwsvA+E7trPzmEvRIhE
f6GDicbfO8Zt56+xgLGMSOakjm/yRIgIQWNmO6uIs+CMY6/bJJrV2jBnds3Bo4WRRLKif8Nn4XZy
nixBt63th3SVyCbBB0Q6jYYpbExy26PbPu0QNxXXDZPYBT7x9VrbHMCaHWh6Z9zOM31J1xPIM3Fb
NMnj7oWz/2FiK3jdkPGWvniQETVbBWKpmyHNuKgKmCuxOlgdOV0ye1XIvStkXqJ40eN6b9YWS0wC
mcYG8HCQKJTByZTUFbJV7+GbOeqBhf32RH5nm7UaMNbRJIKdk+Nkt/aJ3ec5pqHcc2QbvFstXr5m
37ILjKve1kzpIKgoqF0WHd69APyXouvFHRKCM4h0ObfYMKd5kmMpXPY0wkzyLVgZ4MOXuxk6jOXV
aUZgJJIoIfxI8qxc5sdg7FYL8UMC8lxXpPFpIgOP5Xz4YO8TQOxfEiMXosWmt3YTEPhfGdgH6ipI
4y1LGkXP87SC8E+8xDeCdt0dq9R9ACORIaiDI7H25FEOtHbnMzSjfXRFRrLcNoCSOjrOCLh+yaNi
dvWZoLFmY/wTcwu9vavOcIcWZOGY3A4nsfh+azrAKb3rahb4SM5Cc484E0OY6AKPoUe94TihKwGU
XdCOwmZx/Bc1l3Hq5KPGk7kLX95xv6HKVAppcdNcWHNXdD5OXv5ncASi0PTksYPmPcreqg82trN0
ahMOHOhYyeUWAKVGISZrxbtsyeb14xtNEb/WWn5kwT1xCSDDWRvtk9DPmwRYN40FcmC2WO6gaUz5
3nbkleuQlDzhrq1D+/aLnoU+AESCLrcG/EFqS0SuEOB1I+HSDOkqohwXL0SAPh1wA/obHOwBEnqs
yW7dzYMDuZYCL7q0jCdM7yCW1tXOenDDZG+VoTPVP37NK5BRQclBIVht1pA5xs8+dScyCNGTp7hg
9xQCLBEBVNeXgXZRHzpwv45QQ8Z1MvuuibVCGgHd9q2A+IpQjk6ZPcdD9SziBGovN7+491zPn5RM
TsbN7Z/4oecrdQEF7mwAZXRCS1C1LUzR5FsQaN4aEaI16Xf0wTLWhveB+d6ewAXI7TjJ0gfF8kx1
vz6lngNYQXhVj9Y6weCxSKr3iLzIvlas+UWrp8ifQj9xFQ6vsxJYmmdyHUddE0yOs7RmLD3DbYWp
u3dRYW2TEVztAbVn57y/hryh8TFWKWXZ+hH+ub1WM7gyXcbkNaZRzlMikDKdKyd4aIuY6glzA44p
knZ77ZLen71b51u2s0OEiYZyQZCTz02Q8fsPk8y3TVcqSzKGUsk3NGCVgCffVSRyeaZ2WErOik+y
JQY1yIU9SeDpbnEFAZUT8GHAO6MOA6nY0jjtxbL8p8kPqxE2kZJOPFt8HG3bMekHIUW+ILzdTfiJ
AhETq4p4IZ2FtnUHRWp+eXb8JwjbTHUU9URAVBxUT/GEVBlt28/qIjmx3iXDCH/k0y0LMq8CDhWZ
xbUXyRAJdVIhDrdE/sDrZbA2dMUUhbEkVsTzANtzJO8hGtPkXYShqv4KKC0W+Eq7AvVZitKmFmmp
YIfBB2qkxCRQnbXknSaY3hH0cD6N5OZlsDKm6GBLixECHENCVml1qt5DWoxHbEotqlMGzZXoQd6J
1x9eF80nfwCVDH/6kpq6yFd16eRJuc6qxoNkafMzFek/eiPaZ2QhQiwADFJp+w31Ca7YuUx+6zk7
DaXIEMaoOTBWQrlrRDuQ/1YgpBHTAQf92cr9KRR25mgsg8V0+uQK19NoUB48Q9s+o4j2A29V7ymE
EjrZMW0y6ijR/Ng1zMuEotF3v8gaAYDTABVLbdPla1Q9TUNcKXvv8A2NjeZANDsmkUkgl7s9uzTJ
KZe/GObmK0Xc6ZMcvc10BeRrS4qoe3yM22G4l1jF5WUnoYOTuew1kbnBuHR1fdrB6bwuKiTl3ob0
39u69jw81lPU90L1Ehupqv5+UZrInK4T0RZKVTyxsq/D56awMUcsrzAEoOLeMXM04lUNPp8Pavga
G52SXW4xrQQGXJbgjdcTTlnkKKcJLla+Jsa4QKotBTcNaggV8nCkS9LURGgZduE0YXtaEMzAEJor
48ZDNoiDbsCEniSvvst9e9fzH98J64abvPiaO9bl7UH7QZSRgXON8gC7q9iT8WayzxCLJWr+VC6r
X84Wq2PoYTZSI3f9zmOdMFa5vFfPxO0GYUlLCHqeASkYIZpv2zrMjIxzQWC/DdVW6CCN4le/lRmN
9RoZgF8oqYWDgG2FuiNUA9sDdjHSHCVi93pQQF6QZ86EfLyaEybbjeyi7j/uwAtrd+tpJQHS6641
Ql7+EtR642xhmMFfvUj4RgUoFML/vwbSjrekTbnmhlXeYNqtxQiv6UI+KoKoFojTC3Uwu0tYSMrT
GyRfgHaQ7hfxUgZV6RQuWY+5oKdEXXazx/SrDPlmTg0G922V0NwIlJUagIx/A0xAoL7Rx347ojNJ
dODsOhbEBfia9yF21v0Kd1UlnpQZHJo5T/o4iX5Tk77G4N90jPhjCd9Nw/vwrRgV6PukhszqUEfM
ygX1APkQrJH3GfZF6XLhgQaPiqdEYR8pKXqoAGGD5pISs39tT2KQplDhmXPwSVxm6cjIRunoMaHW
j7fC9ZWVJ725244YsRpEFBo3fugGaBhIY+FYnuYmouLR1xq6B9yxSRO3BeApG8xfHt5H/2VLgIrM
XuwM+bZwuqDHlVmxXobEVfUKDUMbQ89yCN0F48MSRTyR3HiZvF9dqwsaVGnRKDgpZOhrnAhkO5vM
EpmXr3yc3z+ITkkIh5SSltPXtSXXMFy0KY4ig06QZGDRswF6SKYcYV64sSQ9wtga6jYIUIAv8rk5
fBzDM7d9zfkR2xXJIqci810jNzjZeuQYQigHz3Rui/JoLlUPr3YsZdfSvmLYefW5gaeOjgT4pKca
c6u3y5+iZAflX01OsoiuoydaKYjCYiV8IZ3grpelsPTsdLlgsZym3grNtfx+BPn5+iGeMW/+Kv1p
RkdmUH5KdV5m19Lazognacusy166F71yWnbt+ioEYe50sQymBpzv7n1sxMAHKpqfjyy6cD2+vVf7
eaubwus/m/mQW6a9BS26JTsK0kEGkr7Y92agdoTN5f0oly3ieMlKi+I4LZDLZScAVicEDNVdAo2+
oMIRcBsykS9jJc7+tobkmpehkcvYbrl645Sw5l8BUxIvOw3OHPM+4T5K7YvWp88hBd44XYLiEAgF
UTb5rjDZNQUNmr7weaHPALvbl/zydRETU/8XPU3b9MlPVL0AzyA9fMYSDyteVn8VWdBdUH/3W308
pmfiBXZt5HmuGvMdhqqQvsTwyBuHAuY8sNCGIcp3munOMFRVeYc2m4Vvxtmlne7qjddjjEGDhCf2
xU9gAju/ogTRY38BSv35onPx8fPXy52qUeqafgqRpwXJwoJ1EW4bm7A5cj4ObG05AvGb1BjmUt2S
8W1WUurcmTpNtb/iLrgh0b2hHYhZ2aygdUXlHnBXym8bty+yN/WKaMAtcQmup9MjZvJIdjHj3YmT
CiQHmd3Gj05kXIxgRU/+QY3kHPBJU+un6+XLT3n1a95t2C6jk41Omfkxq0c+/ZV6ECSkNh5OT0Mp
uH+OnK5K6d+RKGlT7yKz8zWUg3mNQhJ7Eal8NM6GVVhHtygjh7YSrIOX021m4g7XVRnThyWdWc6K
VKRgK811+H0TPZBxNExIQqwwx9LeDBOvID/uYdr0JYchle0qnsG21Lsx1B/dsNhNXG9uakEKowX8
XMoMmjYMQVvFFM9QlrSHsWBdf5wJu+phljj4Ry5OnpwKH2uqr1LoCw/Vkby2ubTsbluuJIAvUi+T
ctjdzQuWgAHGOeNSHbajAgvZx/ARl9DWoWgOoaYjcqSr86e+GcE/WCKwgO3UGo6ZKWyFSkK+xsDK
B+8+pp8ezDr2Z4mFWVYY/LnBahAlP22arLyrEYNe00ilG7GPYpeAp58VhmaVeyCWweFlzfPfI9Se
EoL+I5//eHTHELH16zOShF7gvha7k5/0q1Iidmx4jIIKOUgTKe87U9avc+aZO/EPyLJQ3Y6BhhcG
98a84EO08z8PraVXYyAsNMdOTRzm83KAf+yxmMmndo91697VYTtveKakcqbAMTpI+u/xBwB8+bTv
eDtvJCRc/5gx3RM3SslCtS5jfWU7fUf27HaGFuUeKZhrj0aYskGZj8gX8As0XJHWmjpw8ilQ0KvR
+Ji+sK6yzPyJvl7+d8YfTcFZ/CB62kIs+1bNth9T8jThwv6gVrQ8HwOhYMTwAvCeq119oEKkS16n
6/sKlrwXpno4+7jzEjLU3KpU9TUz/eP0scoScAzmT9vrnFuSbugWx08kaBlzKECv+7Dgz0/Hqqm+
MoK2kfwlr+X5jmDHxVyAxLCQbd3VjHjCMObPX/gcoJYFj4Os7j9EW102lRpmR/ycaR3YvXL/1PDK
Fw4qm7Q9GRm/WG2iXABlcZA5WiRUSrNy0L3jS/wv0Q1I6HNp5hBFdJoa6z1Lgq6EhrtuZjQG5dFj
tk9LgXUf2PvIQs5mNM4hPqayh+NGpmtrarZ3xpADvaa2CQest3oLmANqm4i/3ndG2fJu3+AS4OKy
Zpm2mN+1SnBOpSq+VLaTARmt4+4hEHdLYd8cGa4+33SfryY6D46IUo/OuxlocjDIT0YYE2CLpUuQ
+hpBawg8OU3vpdwuz/wBnHGymdEhLL4DuyYQcv0yFIPHL1m6wV3ep2FsiT8br9zu7W4t+ItY2Klx
qLBHM7x2N7TByOlWsQa3HJSEh9CKKLQ4UPmjn+81bkl1h1dqrywPJuEP/sZOS9VPNakWkGVeG/3S
PyV4NPQFyuxOh+HJR7oSih54cPc9yGJGSk/jHPAhylZldiMsaogNkLUKsSLlKRIZByA4oXH/aCzT
8Viv8h2UbfL8VLgTcPZ4mxs9GBUag0y6fryyKRqDIokaJHt3Kn15JKNyzdTo/+fuuMg22i/yV973
VchTUmOHy98bNc5vDkJ4H2FmirIOBfffL1mNQxp+OjGKNIFk+0xb8Uj9WiPc4fOazx/TCRSwZVjT
kdRnNHRVuEjXHyJ2ZuEprcWe5nOIQeG//3+d65VhXcz7v4caEYNhyctv9BzlME49jbQ/s6u69C0V
FHaQPuogeUW2Sn12P/3yPxvdpVEBOD5EQrCEOJkaF80SFMTtejmACtgziO8ke9QYZHCKsuEVu2Vk
Xqw2msN2Ya5sBHVPiHad+woIkJ5T2PV6sXWGJv8JIMVooaanM5gEHkZtXtsKHzKRRQSmbqPoZagL
m4XkqBlss6IH4FJV2YjFFLwO83hAhL5u09D6uO8+SqLXauxnNhdkaQjiydIjswA7PXmv7ooF9UoT
eEkkBtCqi365dJle/W7Z7M3jGvVc61I2u84yTQTEZavT+WLysfXGXSsa4lEqzePkt83v5sKCrQ0j
Cfi9Pddi8A5SFtHavrqJ6uXOPXT6ALrj4yhJjpPytTVoqbTRMkW7w8Asxt3czVQF6LIRX2Wu/ypf
/0m2YkNtrIN3mxe89V1ivK0ndxRtrWkJjmnpk1KbbmwYtC2IHrMm6gXbNhl3o2Zhr+NH8hyA+UEy
2d61z+jQEZ5mSo3fOnvpDoJMV/OnWJreY0qiHGFK4lNWxp1feq7Kj9tERQhhVk7xgYoFFUb5YW/P
S3uPvSuLZzLzulSYo6RsCwweCJXribaa+0HElAKRztwadJUsi1dpErjKrUubAU9EglW19GEjdf6h
F9PMfIzk1xBjYh7rcSL601QouyuXrZ3j/PuWPgfIWDaap5AjH+ykGU58zjFbfTD50OgplfZbPqwI
Mu3Ujb2HwsWzeII++t4xj4xehwuR6mK8rYyXKWBLpcJZeDO5wMHBlZ8KN45BLiC7VsaVNgDqtcMN
s/YyPho1DJH9czy5HP0DB7rBcKK3MvBdBFHAkiCopvCP1b2ZqnILIRIuMODBXmyglzLCHg+YWVVT
qHjXExagrJHZHUbTU4MUJs1d1VtP6ZASePGuHoC28J5GRM9YXmbNlNlxPp+as5+pFdFdpQDecsjs
ZUeTIWNTqzqiXjNPXSiHrUmkAXkvZnTFNGI5Na2p45eDaBbeBGnVNsWnb1JZVbMKfAShsWzjAz3m
0bNyHSZu5td7CAqz74b+BIEc7+dxYZIBKVCKOfexOF2fSscWLwqPjmwUv0QTnRTtvYum8NmfCmfB
dKz7Ef2006Rs67lsFdKGRtmSelTUZIWywJ9BOm3FGafu29gj00kYwkTZzz3NALUYFdojPMZJ5egz
/7UVY+dtIdz4pUM0HQfMn+sGMYeGZ0b6YbuUmNaogTuEe72PM18zY6ZzltrzTpKKLPggi157nHEm
/qSrt2S3IpWlcd3r0I6KjZkKTCXJk3w6Jtpw7VAnFfH+LLeQba+qdRuRcr0gzcz7Fdru9DbyjiRv
ZSF3qBmw/icwRA3aozjP1TPybCdIp0AFcWrwNSpGSuRn+iaH+N8zwA62UhsoYykZOnhMhYhASw0F
GznD+nHSduFZ6muLtF56iT8M8AQrIDY+KYfevcQkVoJwV6Z+tl4gBs7aq1X6+BzIzSmlrTeusXLf
u/GA9b1Xo/vRRSx4U9yZNxVuTv/7DBFXIPRwY0GueV/EoxWpjYBKshhahMLL42bS7f52fmmOma7o
S+7BwTaHQCt0ovMqZSHkNO7I9uhH+lVvAhRsBmvrJgM90RiNLIH3/Ll5BhM59FTKSBph4qD3/piE
Ck+X328KZoWuWxZx3mtk+/QAlyiRl/ThvSL7Xjcb4BY2Ix+pUS9UqO335QzwDFaONw3gE6BKu90m
iJoh6y6T+XmRZWukOqS3fOiMutBG9qTIvrdSPEP5Z6laX3DZJodw6uDyqAqQGQ5vz0pPyvS/MSaE
TmNRIxCThco/8uOxIDYbB6UZfGJr9U9niylrZTV66qlFWIi0zhAHQrI4cPe9bL2LErK2tS27WQOk
WnC6KLf1JmjG+VvDt6TmDY1p2WcbpPoOYmRoS1yRVvZAeYR1650z2n9yD32p9z0RldzWchlQD4Rp
tJadC5R30jxf6DcIvNj4nmLbSs+mZwaWmllt0hD4LQA/3AyvTWkjiGcvOBNNWfuVPZa4bEga5p/w
bMglSw570iwJrX0IUS79j1SD5y2TtNtHz8e+w6E1Dg/UCG/TiGqGqqsSGEmBc64mOSOlrRSl9avs
CcFPjtxN9Dmxd4nBZt9VZ9xrh4J5DRfpjxu4lC8LpAEN1sFho3yU7jU1YPlgpYOzJ/OOjfrfnhgH
Tgk0OP/5OJmeUphcpfSAMo1Nc05SG6C7oFrcb1s+DAsor6CIFIY1VP4GGE60ov8gSlOeLeI+T9Ve
JFKVeuf69IroOedVX1INMCaPsxidHNk0l5CJb3/7OfIMhav2b2n0/X4+C+xFpKo7cb5y87UzukoZ
++LMwbToFh+9qF/xJHz+hK4NEoLK0oeHAa2BZpa1DVwC/PP9+zb7KT6pWqp2ywkWNVKIuw8Z1F4n
krCK1eNmvY9fCyHDTGIkcJ2YcOOlbqPMPAxudO+B6RKlxoQoRuYqtQiULen0g1Rudkvx7c5Cobjg
6QZFDuNMoPKRsKojdsxQV8Nbsu2hB3kAm7JfB4zRD8wFLiF2JaR2sQTSVJc+aryxJt+FhxduHfyM
jHA1AFVqF1vuaILxacKPtR4L5YNxXAtnYDaJWwGx0A1GcDSuFSy1uReXYbCv10qzBEIypvCEVKNC
cqoTcsYSa7AINpFREFwRkVBmuoTXcTlPzSxDvntpslyfbWSEaIoLbRCkT1ICb3A8fSFvq7Mcxzu8
d2IN3vcJqf6RDMSKmq6na69jubejihjoETd0JA3Q3Bndn+E1Egekq9l+rL0n7Z4/G5HAQ9NmkmlM
GYuLsR9igdWsVV1av8G1uXoLHhS85dkq/egHPvgg9oSBZ8iBPNEhfnWD/iwElXV/undSrG02AGff
MFCstgdcux05jPcIN/hXS962YyEr26D36zgv2U52s8WSsEObRzg1ClawOePx+/eCjv9C2e7DeEM/
KJ95pPsw2f885GQGkz4OODPbSSFKoJQ2ioBXY5SAKzJpFuCmsrB9Lcs8uouozN+HK03eg27ESLVz
tsNyzAQC5QqWPBWJjtQIUTGn2mKZUTpbs5RbL6R0oaxcT3LdCiezRfsMEWWDQXacFSa3Bc6G6JPv
cACJ1xL3+giAF2XSXXkHP4AD2Tlq63RJa0ZQzKAQEWEKgVWxzuWJCpuito3TjEy9No4Tbwl6Hu9T
ksP4Ze93zw/nAZDtzq6sC0NP25tr73HfLx/KDGf7h3bf5uyxc0tEdqIunpOv1U2dQ6cjQLLMG1CY
cIoKsj5X/ErRXSmAgL+JyugRGx1Aa5wDpE8qQDdRq1IZmgz01LvHJAlF0GzmoeEOb2jY8j6z/M6h
+eDfCimDjwkVfQVekbdmawCSBpX/ulIncxvFJFM2n5S4vxWJ+GnLCncGXXECQxk7tj3339omIhjQ
+eHe6JNww7Olqe9Ec3xyOArbuIxmuUR23UyNVE7pws6X+/1l+JQy76ColrIwzoVuir0LIeYV2knH
6a6JIoE8JbIRwBhE2uXnJBjtwkBOSCt1Um8gc41nKHBOI7ozwupSpy3od44po9CFcBXzDWsd2zvd
sB41qnSoecAk/Rfsqv+3X3XfFsPzZFXu3L3Ee9JK7HaAbY5WrrvhA6ykIW7E4R/ljWw8HqkjJGwM
im9pyUfRLGsmd5R3RC0ZmJleCuFfYjk27/ONn+QhW34WUKNBBPJ3Iu2NoOSwsVYu3LsAHTlzoSrH
xrUswCo+WG/RfekDay6YRc/Eyp4uCA+BpGZffSmTBNqvSGHjEdsZBtsd9gW0dNjN9uoHLOd+C2Lo
qgCTvXqWEGaqwkedYRH11gBpb9eXn+BlOVfQs3ivJSY1PE5bSj6Eh2l5q88Ba0V8ldG3SWol6Syg
FV+d6QCY4GOa6NJQcUPr3Dbqe6Qt+xbUt9sohbutU0u4xuPta216CeSrP/KDtAGN3lXEg1jLa/KU
QTlerd/cv5nJ4/KJHh1lFKH8XegO5D/TkoH8Vc+gNPjEU5ICyAqYqkIp4fl86yaUumxr5sZ2mCc3
CaqeQc/I7tktUIu2J+LnM0TUVWGJLrQdHJ64P5EW9PpgATawNxh0V4f000/q2TvKdr9HnTdDUv/O
/Oc4erSQ+qvwQ17pc5MBQG8JnqKkBahHnR+oAmhMrL7nITBhILDahV3qll/sqFSibR8QRN/cyc9b
kLyJXH4/x/ty3Q1A+RZJ9/zQ4Uionc/9d4kQH3MkCi8oCRb1GGmE1WHRKj1RY8PjWJop45GlhCoX
cDDvhy8CwPLHQ4GLqrj3VaRTlS4bj2R/XK+18zQkyJobc7eD3b5ECwagvGinqbhehHMxSyplj/BR
d3umjge3FDxETmnf1psJ66upthJWJq36362YIsE+WprDIFXQ8RIdmO/pS3g+P3aQYBq61Xux4hq/
A3sQAuhd9q+VCqP45yjIgGEhW623QYrkFmqrzMM2rrnJeBdVkD8ELtSkJO7bDyTMk/ReQRQGspzx
RCt6fBHizX9w+AMdKv5Hy8cu7VWGgfFQsZk3gA0KuKw8CED6PsMfFS4Z1CFN+6DjiyuRux8oNVfH
9hKxKb6rZZN9/k59EkAjeGGq0ivY7vov0LUwhEUQAooKzn+ESna9Lo2YCAJToWAJN2BD/i2z700Y
Kgb6+kh/9kLQOUyK8cLc4MhXJP+QiUQRnQ9bqjRYNFpWo66puXUYpMKr/LUzzixaiaq//1vELoOP
u81oWtUAUkpw8cHavsldXB2pqxQZkkO3myZP6FyV6ZTklMYOUbHXR5ifCGQWxafR2wt5RdWXm+H9
agS/aoP6RWjJaqRjWzC5ymtMX857MfGb3dD0a+ngZkDpwfg+g4WV6eONZzhWmwZ1Tg/NwftihVgY
CyEwUunDHoMRPae//LDApF4edq52499RxxwAMbo1dJCuhWAVh1/cLn64QQLgXffvi/5aq6YNdG2q
29mUt0Bm6BgGtX4rW2WoKUFoagze5kYieZ9v/LwFk5Lcq30En0++tBJwIbLQHSUYK+CVqRgBTTMz
VQhMIrReSq6cFotp+zRPqUt2i+szGnuXIg88cpFEjv0y7OjrK0yXRf1nQb5Dw2SsIRXeGWtLdn6W
foTnlbM/FB3x2fAhczTd8rIFogXcLnUwR4j2QRaqWmuKXRLAVTIL8xw5TmW1H7ICwYaYNhzSma2q
UNYZh9CvkMnln3khzfJ8V4oAx5LFyQvF+rU7/WpfWREaav2NP5ojlKBAVPk3An+P0C25CxJVmZ1t
JWPtOLLH5m/RqgHs0FNe3pn7CvNZ2ufebTbauC88XL7O99+cSVoC7tIrkdi9+nQqru/ZyTdQ09kk
/SmrT0wXtUEmHP3BC66WqM1SzuaRgaSCsN52YZWYLzR3hAV+ZLbI8YNr7DNuBlZ8xt5CNL+SrEeH
BQDCJU9Ki5Uhi7v0m4DP4iVY8OOQXAsPbG/Pct2JigDkNDCVW8OlYTJB7tsGVdDtu3TmJhzIwHN3
btLcgqPiAJy7MIFY8VCwlmwWV4Gm1d4RfUxe4xaxfHoG4UtianbCfQkPnHEl1ooeQfSDIgqBa52A
ma+fOGSKZ8wlSBEPuoHrYPfEbbemHvucKJB0qfDzYKfQIOpbNO8/GLqE672UvPbQhLR6TpzaitmJ
rJIHBT0rlgEI/WTiBxpF3AeZmEu60lhnM2+B2QKkt02EYEVIzso8XXa/kgHX/DXKKUrf3rTf53cA
+4S8zEp4G8Sew/vS2dTOPrRAbbsurWc0wruRGhYCnbZsLh5tBSvrsCzSpdPBTfKGuIgdRcXdZu7U
slqO0W27kqdAS1Hre/w9qQ7K/fa1QziVSjkSsHnf4poHWRnNCRGXndv9LCr3DMGwoDhrtPwqptRf
O2jRRyjWPrceF3bWnk600JUhuWUIbcJKYf2c/ovjFAyd6CjqrRX/IgZWduCIoI33zFToQWFkIxCA
GhT8qdGZ6FUDKxlVODGRIPbI761hqZECCq0qotvJxkv2e5eumkMY7c8X0mAFU/CvMwy7VPsD9wbM
EfZUQuryUdwbUQZv1sz0gtzZvIlQ/7GAG6laTg+X2kTFdkXCSsTy1h987nApvLadRx192+/lI+l3
bAPbcBYOD92DwoMjEES+fM4VEWidUy81bHhbMPScJdsf/LqclVVyYHt3FSU8WYN4Cgn3C+Tr2U2o
7ZCVBDXfcH05xXQq9Hg/L4ETx27zwv0PJen34VWlkiIZvghMrv5UHD7cBMAaYmap0WCTatV8UoVQ
GRfzkXjdGhpsQmakQkG9Zfj7wWjTG4rukC15xeBAixh8dlpggoOVlBNrsCG34yeaSq1mVODF/rg6
wyB6t3OvSSYiQAFjl5DGJNElqGERrMYEnqA1ae6P5SnpwKBwe+AshOBJp1yJzq+8YG7GfJeTAuo+
SNu337By7AjzrCI5XToICk/pLyukkQXPEvrgDVTF/EpQMjsO/l/X1CnXDEZQU0+V5owOHyDWpVoc
nfSSEtDOYETveez/DrN28R68ZSmIoRoArEAxJJ3WKsFhpVCkRouVcmyHuVnJf2GsrBi/7f8e+wzV
z1mZrKlhv2xmQmCDE+Pxew0iAI92MH9v5r1w+XZGdYCPasm+3IrxLpEbpXh2UtJl3lZCp5YPDDhv
B/t77fu18bcwUShK3pMlWpxg4H7C2ZNeqq+HPKO7VsUSxwNEARIfaMIWLJzMkWJJDv3K7dobbPS2
hBmTMm2y7NwYu7OmHZ75WJcuEP977rAkpj/xl9GaPsMAECshdfN32AyTnZfhaiFfxMrWFAccwVWa
4aVJlyS5EyKfIcbf55DiyaptVT+iQIP46me+TPPbwiOj98UbJ8KKXCGNnB/k3aRacdfLWgKEWDCS
ZOcuIigOvsk0mNXIjzCDGzC2LkAWRIEDXIZMx1x8KbyVqG5vIniXyBm8eCz2Iy0a37jqIFLoHGpR
/CNvO9lv2KwX6Xk2NhOaWdzZXEWtqb9kMNMnsCoc7ZMTLSCF5rGsYj9UIi/+HBjD0E9xMtB7Y9nN
bQDbgji4iJVUz6wpM4dysMFepHhbPZPWbuAd6YCfr0afvQeC0ZU00LbNiArMGOsfCL03mmCc0xF2
eYxyItfGHqN6NIM9dJo7qgOcJOkZDdtZ/dH7IItFe2x5oZtqO/5+52WJVetRoHBeY5nkARkQ0Oqd
/J+0y+zHmZ8EikUw6bJtfVx4HCkKP6Ui01vajo7ipiSmZ/ldr97Gi0CcnHPBxEdy40DL+F3vEU7m
hll/WOWAZx2w9aJ1M2J2prFO16eAGpW+Dh/hEc2KbChufUivxAcItp0AR8NMYTnjLC5z7gBTCt8U
tO/wsfQVym3AVNq0BBeIdnP4/KObGXkXrbiM3M7F6jjJDubby5+GpK1OJywzNMvUS1H1rBDvh5lL
fWQopT7kKsKNXYn1ONm4Oo04rEeg6F6RT2KAnxkSW7bGrF8/cvjr4vx3mWgVxPIL4ha4jelOhMnk
ne/gr5dT6KOs7tdjxTkDJ6jhGujxAcXJfXVSZWwENWOlY6ZD5jBTlUfeLS2rFPTytawfNISxrDiw
+Pfbeqg66fkYhUIyVtDQ/+NGfGbd0bdPi3ZR05D/mAPRF0BuQXOZhlnIz3B6S8b6+9uMFEsjUr/i
+FsITdBzkH29/PUeVyfAHHM1xsjeJbj85bN0kbzQIqVfnlgiWjqpubKM03dKwRUDCFp7YMsOXhB5
FmElAStZj5VLLCyEJtetA7jSdNDMof/ETKekPYwzq9nhLwgdOKK/RzaaWOMPUHlEHRSgELoQ2BPd
pUvkKRm3x0dkNssJQFd4qd6m2o82kPU01pU/HuW4qAccFRfgySy2pEDHlHdWW0u8nwirwJjWNnNn
Ei9whjNpwy0YVpnpd1hc/ZIe/mAKYR38NgLdLRCd0b5X43X9pORvFFQwBsQuer69LqyzmxLx20sK
y6ayCsaqlnvY6a+xgtKfxow5Uu0c7uaW8MlQMsNobAF0LMbxIRxXmeYZSKDaE/IkUtvexybFD1tq
BYZChFkmU9Wme9YtqdFh5gtbBTT3qEHaqFh02dbyYID6Kf1UqNskHFVnb9tMR+O+kkMhIUt6yM3t
Dk02tJLkpj8z/gdsjbbj0PEexx1GKTEMiBnePUac6LBERqAtKeTjVq+uXK9O9GQSacZ8tZeXrWjh
mIC/jSwtHgxdI3/UG3GXDNfQr+NR3NAjYfVVwgAuoOcQFVrdfMhoPqAb3B0GlqUrAHqSeD5+bA1f
kjSzyDPimDD3lwYrVNwInlpgEostfohA2YoTvvaFhiPGHpFNuaRnNQc8xtPmkQmdHRz5oq49RWT/
3v97iUDDyA2KAK4I2DP9zQ0u5MEqncKIuxhtbdiofWIrP7QhUOX7J7AB9phS8PIIPA4PGL9mABdc
PbyCkLjivOqzU2dzbn6dUmX60YxxuBINGBcgHGtPQn9Kj9nEZRKLNrQF8PYde6NtDv/KAmjHf4uz
ByAVhTWr4n8hJWBWLw3Tag1WzdzZ5f8Dar4dF5CAiEPMcQfQTabivDk1uLCRcSTwC0ypP8212o+6
5RNnIiIzqhhXAFmC0M1COb7u0q1DcceI62r5Np7ZXpzil6Jz4uderjjzCqW5ydN5OCATKJUwfcpB
DUqXPvGALuJ90rwHmpqGXIT6RX5Zf66/rmlw2uTfMmcgaPw1WlT6VMePCCZK3N5iozrH+0YIe+B2
YU8gu2Ku2HyRnFFFqSMZOtq7SY3N6ayg5QwX2PIFG/PnACuNuI4ifgQ7g3G3KQR3A3VSBBPLhXf9
gbgL65krnEDFEn7qejudfxXNKgMQFh8tT7IjLsAqqOEkqJpqza6dI0DjSRdQkZJew5DHT+U6Xsew
y0AE8z/N5e6RRBii8wfV316gDwO/jMCErbyxiZ3aTzuh4CBytsJm58RDSHa3xFdXDoRlbj/lUcV6
70IDezt1982+VCHgKGnDtOq/w/ap5DeUWKcxQkRSafPT8tZ7jw+IkNQEKzX/VunsARLUfCud9AH2
PfAszanibxdWzk5wTfwy+BuOAfjwa6KEfNy81piy0YKvm3fjCz+JtcEltG5kaStckG5BZX88UKEd
PzSLxAYIrzbk1AO9COjf6zjbz8GYFH4opNQM5CBzNXRQPCt4Z8GWcl2VX4090KaH5WfaV5WDUz0T
rCiwyQ8t3b1t8wMIzmrOpsJOxpQlaVEHfjhSSfw/k21x1WN9qK5kTa6Z9cx1Z3mDwSN4rRt5QRVE
g4+KT4CGDwAGNpj+ve5/N6bp4Rf4ZounvdjR8YW394qskz+Hd4CO5Jh3a51Y5yLP5DaC6NkU9Hba
kySXfRAtZUfWpQVXWbJHWoaha6DJkxGuAytRW2QSi0eVljiNv0Uf4L0pCnGJu9BIF7lJAxN2fXOO
O9HpZqXn7Ss5em7vbgqGp5gCsfmAYmZngbI3dJtQd5xoH6khn+eS0xyBgB54pKnjM4unEW3NG/6u
1V++TkGjnul2iMs85kkTtvy4U/+7TmnOw2jhye53EVBpXSvZMd9J8MBqufyQRkRYPUbuD0rH4fXi
ycLMAe3IU82LGs8n5XU56dXUm4ZZAnt+6uU2+pEduFWlBqvTTXwHPJtLU/aHmJ5Xu77IPP8PSow6
i1+bTiKXySFNhb5mP+iqHvrlf5LE3IGR45FvMsBGQnRlaZ9CAsCuhEdn8zak7dspT379A0Er9Bb5
vxhEQwuZ6V9QateFgnd/j3qvC87SLXaOG7sY4m+2aOHA/CatiOHCp+hoWLleT6JDXB+GgSUjkoU0
I9UNVEkiws5EvuJm1mxmb+jfNdWwmiWHZ4WNEw800DbmvQifwGbamMlOZ8YcMVk8vUH6RJ1V4kvb
UCH0mSJggYAJc1o84T4qc56WTJirmbp5C+Ahy6bKFKCJPUxsicYaI/YHNgti8GDArLGsf3B0pW6t
/DelJNGY619ZS9iLCVdtNB1gHsVwDgjptGPVnA+9dRH9YrqCIagwyFdSeMSxndR/FinJM2jr25P4
CMowtI9uZMPS82YHz4AucQEmLGEMbLT8i2yjOtSzMy1pgkBxI7Nbo8kOgL3h7cX2n4HYZ6sH75UI
WNUAbkTJ1fLa8U59P+FoIJWg4hQSDxLEFV8bg4kgl0F9YXe/K4XdwkNDP6tZxNExboq8DibOZhff
2IFodXv17VVOggp/7PoRI6VCIG3mwn/QEHxzjEE2uRhZ4hJ+Cbxs1Y7Byrxpt4u9eB42bE/hcfeW
x7HkP+UsM2Wvn+3j9WQ2rTk6dneL22ypO5u/BPcj6H2ZTooLAhMASQ7Qd8LO7xsRjbzTOhuWwfhv
rXuRVRNLIb77I8Em75h/uk6AuZt5KRxhVM8R+o0EQZE0UQ7yzWkEHyfazjEy3p7MR82dRfJoWRwY
YioXP1f1M+iKCfT0xJbkJJ3B3pS5h43fVEIL5YUWLeLkCj/CPTwyE+Ix9bUHVKmvYmJ9ApXjqBS+
01Cpgor6bodfSbG5nWuroeGiniz/42r4AD+QEZyVSKIdZYtXD0F4ESNK8iI4jA/ClBIgMmbBabtx
eeQreA/mSHch3BKmTwbBYr0jdcCiivDvHunCjIR3v+nYGed2qtbMhsnIIsAVvqGoCac5OqKUXqOL
temUcFMjTUDp+De4I8kzOwFXRobyNds5iAVYhR7g0Jo691NbdFW1rI/degkCS/lJQtPchvUyNDg9
GUpVd4yGPQqj0watnJGyiPRwy9Wqbq5DUvldFqYZMHNiWq3eW98CQTNMtJgBMgMF5jOkKQ1D8vzb
4D0F7C4YPrSyCjqqF8MU87dLI7O6gvAOG2zscYoUIehTIeYWbMr3MwV5mII8j8JHKi92u+ZQqjD9
cb5gpA7waB+SxNfu42esqH7vu7VJ/Rkos6aO9GkpihYQWYLAI58ZK+Lci1kCA5wgaLXFoyoUeklO
OjCQ7PE6vEDPfoz7teAlDwtDffZv68LxXZnF626E5BnaKDkgXOcPKXF9AS1yXdpO854JOrc0bdSJ
iqkbtrJUTakBYa/qgnMAcwCCuzzErQD5NqohTaPu05rF/m1DrwpCiY/3lar/w7RqRe2o2hm2dn3e
aCbDykh0vPmxVIHbsu2O6+5YoQj9K9y6kM8Y6ZDim/708cMf3Exum/Ex+cZgXb7XhsTbgAeYCU4u
OOnI2Rsbavp5Hgw6a2cvjD3j998+qYGb9YA1J2lrlNXC5pWrhooZkmoiMT2c7BINCmfAcQ37R5qP
dZmMugQz1WO++KYjFyLWRzUU9ElrdCzj/hSkjDJ4HbbdH//o5stgWW2IbImYgBoDZOTnEbdDxc+f
gab6XZ7WdsRYpFDYA9VGARnda3BJ7qYYp8AN/HB6GfsiWX3tbuSg+7oQ/58Cbc9CzqZkdiBcRXPM
oAsXQJGqHHLIUPlt4gppRGUvdpqvOUeE2oVwyMupscFI0mmPn2iKHbl3/fIy1iNRR5+z7LOBnMR2
CEq2webJN4yqT1mPygHJg7ZuvEkWpjFlvZg7m2t4bwCwjwTFxG0Fgkh45e3uNnp8jzVwRhlI+lyt
/tUPZ5tIp8KNkKkQ050yzF0MHc1rwChBZ0dEYEmqGgB0dbYcbyeYnnUxyu9y+pDfbQm9iOHcoRWr
MLUbEySWTMEwkP3l5VRgVNk/doDeiNyBTuU86Y/pO0rFj1uRoafL5u+dgCq4Nwj5TfR1bDnvnWIW
YS8iR2/3N1g81p7LNa7wUMwO4IeYx0lxbAzen1Tp3vTJ5O1QgajJXZHFUbVCCIeMM2EHMt2I8gDO
jyAibd80kBuLCQgYdJWVZi/dcYQJQ/vPrEjuHnDw+oM7EbDzCOVCKn5AEfmS9oWFmOFNMXYsRC9f
Rdnbcc6kRPHgBcRMB/g66xD/z4ew4kPiF1ERDKSugy56Pl9mwKKQmMNqirq8pLwV5iGHJoyAEnPf
GKiBFYQZCHYbyMecNIaJqmcuiQGWAqCczP0spKC/YSvaS8c+ANozxvf31RGqUBVJL6GVgsrw7JHY
f5ughheyQRUSDsGJpMNm9YiU6uDfGWsQzcjW+oN9yXTeFlEFklTKXeFLPx0RLWtJvEnss17/0PIF
2DGuHnek5JRj1MMAk+AVNT/6SbEcZvDiPr4eEoPsH3+TazesazYEnfxU/Qe5pJGNoflJn/12llUs
jcowk7cNhVaYs4P1zVs6EbM2Nk6gGiQTrvVFJvc4Tvd8MWI7Yu0dYMIzLosF/q+Fe8ontRt/HjJ+
pysCyBPybXURpOjU+zuySiTBG710sbJpdWk2YqPkLwbXCnqLvfxI5I61S/YwJGjpjewaw0cA/WNC
RWcZmcqZZOMyj5X/lRkcgFiOlcBICdGKETnLbcU2fluhLPdDhkmSHwdw7MHBAIz9vMKqGqjuOrEM
8O6jWFhQdfUN+vUlgqLsxn86uffOuWCaeHx6JtR39ml0D3aZPzdIUlv5K7s9LU3LDqoxr04RMsKV
SZF1eps84uuA96Ma+MzEhsi97r1w6oR5NkWe1E8dD7Y7LZuu5HnjLHZVXZjMRZ5Z7mEtfuclvmfn
SvtI9SCAUkcmPFnIqv5JnnghIiIJcWhQVxpaCHHQvK8MFgiyDBStLc5hFYGHKzAqBHN2xmJ6VCKR
kE8HD85db4GoEqIiZbhYQv62p/7TNeuI1h5hxcqAy4Bx3oGb0qhqYg6XcH1y6l/LvJB20cMo1zJj
BBl7UuTyOf3DNDXrUmOFKAl3/KyUKHYH6kQ/Wg+13yb0sk6ac309KU/AypoW1rhOxhHlTZHs46zH
9i1NGwrvVTBFck8GlbtXk+A/iC6hPz2+aZ+yNquL39X2ISnQZqne1/sSPiteubCKxqPQQVJ5o05x
M/09vUBeOxLnLutc3Ci/jEBbUKyDRJ2FCdP9IkZ67XK9GODnO6xBZYfapS8NXiH9R7cqEYZOAx3Q
WPN0ZMqjuxu0fpPnNbmoaa0yBqv/1q426N+T28pFuQqIFOn80fVmXoZt8CImmUo5vlKMYvAgTTyC
tEh7dO9IihNqfbnL8WJAcKRVh6S/JAQaaDcb9uL0CjESJCgI/nFBKHtYoo7c5a7APlJKrp5LZRzn
FDcENh6fzuXjvx8drHlq13VGdOK75rk7CDYtOSe2ve1aqMArsfFhbZaJzfHj7Njp9ADwBrX0Qzl4
gEeRheFZ9HYgY+spSMpAxt1rOLeWVeGdenUtga5pSmmh1CNOpcUzmsXeP0ta8OlJ1d2RdAOuPWTv
Kpw4Tl3h/tHoqnJCila7SWpKuNXsqO4Iug3rHw/GUZNC1l50WvYR/34kTAlRGEQxEt9A2bkGxmiT
92nRsNGEZrPsVeR5y4NGtuzEt+os3TzXh7eet4LhVnSjYIlze0ray8SLy2kr7746Dw1zTPYo3pJA
JqhUmcwPMFjdCSBEwecwlT/u1QTWM0Ll+GIB1lyuDsB+b8wHxaftvduHGjlMlBBEFebWR+HBoZ0U
AYjvxwLeXhHxRMpFmBpfQjG2/Auqez3oV0CXUthMp8kcUEy0ApeWsCU3MMCFy2EwgpltxgOmEFcQ
Zn/xh33KeHOq2aPnpfAq12UAmRhlnyfvmqgYhqP/hwAwrqOLeFMOTqdHZ3lRuViX3f6AR2v99ZVs
xjsTpzFpmsOefeW6Cy9+nJWDHF53O3/B5ceGjZrMnNHuGf6gj4dNJM0hKu/UGVxFAQT5I4JtnOdz
NUlMM4B6Yn6Kwr9MQGV0rVVZwzPx9IMygpI1RepiTQTyN9i3HAEEOM7t21mNv1UaIUM7PyyfKx66
FdNvHkV90lDVqVdSH8iT0LtnK0rtqzg9CX3ISO8GonLAEZnDdz8/hdrChCFpTOhPNIrpwmhk5To1
PlRiGjsJ2ErbRt4MfI72HQDJsfgdXq0MpqxywARwnEf8llGwP/1DrclQ+slw0sqgJnnXiaYhadNM
FxewDTuTQXqyJnLFubXjs2hTy6OA9FOWcbRffadx+kVJJ2q7GNM10Z3pIwY1ZkB1PYXdZ2zALQY3
U/meEBcRxY3+oPjMkQJPgSsYWbKNTNEsur3gP8znuUtEWPCSODG+DuPX2wBVGXOePmcy24Qfe2Du
fTRMr9u7k1k1Rrykj+faWsBHRqCM2GN8du5kfuaYzUhrznR4SI3W1YXBxvL6EZrbXfn+J7rfjiJZ
3k9sQVR3qrjd+NfR0NmLNWK7auZoP/vVtZ14Z4zXjL0XTl6VA7DIBksLvAz9QLRgMPrg/On9mmCj
ChxftLhjH1a37ICLwKZyZL9ETZhdzJau/v2r3gJl8bhxVBBWynfL6w+sl0vAz66YSSjyACR8YoIN
tQ25vqSqb++e9dEIM61e2WPEgB4ok8mqcwaC6YtRj31PfA27D2ClO6pz5Kw2KHa0ZTkThVpzuKmI
/WI4WjTR/4FrJlHwa2oMsBvMctFmgX1jO/C6AF9rKdjws1AUZjD8AwyWqgN6kTYCdJzoZVl6m+rW
QA39IAARhb0PcWCGONh1H+fDOt/WaYRFCpsa0iWSEKMojyJMOVc1/vpW+ovp9rUw62K2vjtge5Vw
9NXTLlMFYkStoS/FeuQbTCnp/5UOMMxfu/31OE1OF8A9SKU/gq7p0rDipYsB8i1BecxK5IuZIult
KnZ98lHVLbJhg7QmgfJuSAQeHANrV31iiY/VPCLQANxlDo8rqipcAsseDU//lxuBZ+YrbV/NkGKj
2bxX64dOvBOiuzVUSS/c4xEHmV+hFdInGEkXNpiEXbiPNmAfcYPLJ2aSHw7naDbuambqByzYuLUl
ElCYWYryf7g7R//XxN3GXdqpm0KLLI0UrTJwUeSLS++LyJL5XcZU0GJZrb4R466DeZ8jQBYctZSl
6goqwgLamfNrmi75OGbIiXYywcqqTedCXf05sw0zu2AU4PpfGQ0wyydLgCI8EQfMnD/oIAU30eGl
Onka3S/k+Gclvl4hybMl5PtBODoUHMFNhs/nfyCf55Ng7Q2Gu9DrtZYRJRBF8JV0z0+yTkI3/yNF
zxmbNWplLqUjrXJPS/L/4KDR2W9VvWO6i9i/JRYbPPbsrY434bONCi9F+Bf6t1gnjKpfgi6abw2N
qqc6pBdBurVs/1Y6pMFfZUzpgu2J1bpoVds/U/KLfy8oiBrgRbqmVDrYpcYzS/ARinpRnoW7m4Qi
mwuo0j/nojK7VzEjto0usWq3l4jDO2it2wR+Dp1mU+zSfgzqTVVsrXB2PxudvASwKFVyiyoJs0Jr
ah+AT2d2DFacPi13ZNwQBj/lJ91q4lP8xdINTEW6KS3byzDmCLnx/s5mwRnT3KjrP0eRQsWS4u9n
2bVYAPuWWSaIhNXvj1WOKq+ZUNCNiQNx/EMk6VUvViM7mRdGtgKZqKMAtob7LzFPmWg21Om7zKjv
xi0z0QfUJjkIDYg0W7yZkps+FkD5jv9kU/OvcyYwORoNvY5dFg9C0Rsq46LZ7GG38FoiTjnnJdGp
x5H9RMinNP2bB6LE1zB2d2WDez8gZiBtDWC3O72SlXVH5lolOFSwRpSycvzjIX8JwfKR5IS24c8f
VXJGTBMPK3H6XsrZ3VVxitAjNCXPfEqUcMeUuQ/MA3NHSKYtcm9ztMAir/Ul4+ohfp5CbgXpYGmQ
cy12e2FBCaj86cIMdIXBA/+Xtoj95LQkTQHLietzBzBncJw8kaxYxWuWNA9XxmFKdf91hvQYWpEH
zUYD9xBw6BhlCm5ajkBoqBsDf6NiZD12DYG5Z0WwR9XhwDBecTo54KXAZEDijZ/Ipxis4p7sB3NG
EE9nyirxIXy08tPCKg7Ywt8Kp3EOQMLnCq3ZItD56pReZenxpQoU7+USdvH/jqqBvdlsr7TbCAu1
L2VGOdxDxOf5aLpAQc463xCNFLP3rCuO0+r/zuRQNf0wmWuQerNfzb/hsW+tLELmzqlwjrWkgGeN
f211ZU4LYKSkzVaWpL9gqCp2hu1gJNyi6F/pZhXtPeSwuvLsizB9e1cFodyJiucJuGS8WO24u2rg
8Q2jbgfRFjZnQSSDTiKwt79I2VOUb8ZwK88Zoz17eyFmZvijAAtQE0D0z7g60iN3OIXmPnap7Nmr
LXejIi9xm0nYg7Pi7eIyIaS/m2j3570fDzSoPfxgf0d8cNSvw97/uKhO0ckFrXCvKuvJ7FB/Ebts
Z0UO2A50BoFC6PudTDpMHBt/Rr4O0N49zFcMWYcdomGLHiT7UfiXbZSPVVYjBApV1wNmnkTsLd5R
SMr0u1XZ7yPNAF9Y9gaLpreBthtIqCTPfHZBn6Y/tWqKSHkX1ETmuMeMC9Nqv4WKXWxluiXEK8JY
dN6ZxC6d5j0NCATc57hs2KrvsAqgHrN8APYjY23gNUEOdfcxAYVr53nNT6QipBDiKEfEur4vQNsS
o90EvP78uddIAHWuZtvmEbd8NzK+sAumOflf7rYsilnivg8jCXhAI10yE3c2/cEaVtExx2x3EtZK
kAP9aszKR2xyy+NROQebErvrZ17khEZvb+5ooB6b1ghWUm6zzRoOf9UPQWchp+5BZEEcBKNR95p/
9kort7dugOS6Z8G0JfUDP5MHqnfSwwVswm/7ZceBd92cXksJsaQ+RuV1jKIGhpSxT+cSK3NopMcq
VGhP3twfB9wKmetcm0pfoCU41l9411YGbXgUShXKRwW0jJNpcBpx6kgpDcNKbcWN6bEgyuN4u0WI
qdm0X++/gvZlWjM3VGzzVlt53WSrwB+xon5fhqPkQj2OgxVoIbqTM7HatTibWGBSca1pXlQspl9I
sA1Sl7osqozu/rexEShzy3khARwgyk6QW7xnR2MPocPnvYajUMBos3ETDA0HUXL3m2pfXyTzC5AR
+sButoKM4MtO1Jcnd0RIvNyE27GwWqsNWvSdRdeQQ1wu+d9MDdanb3C94ukDo20q6WzuqoQ4PCs7
VHow98iqeytONia1gD/aCeA82vUwhSDx4FKgC/72Nyc7SJ1w3PRzIrh4P5d8ghW1kYpGLKVphgwK
jRAG1l8s7MwTqYDSodDdP6eUojMwXIIeuGXD7vhclP4zKcAruPMRtgviudBkIxfge10DUwDZctgt
7npcTxiXhyBdc64/gB6QWDoIyDvD6DDt8oMxHgtH1z8Y6YTwNPWjIhg4F9Yfi4ulhfzLyNnioLeE
UZnda5OwHHlPsaLOwWawftRH5lZz4TOUI7YL1xaqHhs4mbF+ADpAknBdWU5zDBZgKx7b6VAFJUBc
QNkXDAnqrCc3GzR6J5zUddNhCbwXxu11SDRE8rC6tGRGNOKCD6OXL3oa2bYgfBp2r8NAmCHYX+IS
L2N0blYUzPUcmknYIScSyLktNd6AMQUWAmE5LwxwjahK4xCrx11gaEspCT9G75JwT9J7Fma9wvfL
R1Le5vf4zba3O9QKu8Zj1iAPlx+RNkAigezYSKSrasv5WQ6PzKpMjcDngE/FGOXLRgjSS+3FRjmq
7q2bRUcNNeBVIgrQwqJ9m3Y+141Nq+U3aFsI1RpnByeW8tMf5cFwlMiQe9B5R6jmHB3FnvSOIaPy
IhJQBUG6faRoOfXOU3j6xBlX8rP/G/gz7+ss9MmqMLA7RZdW8uirZX/nmsQEOXeoidsNOP0JyjEb
XNoUSV13S9Y/1stmLw6oot8JDj0AGp4VgQXwLo2QRUjA3ORW/EEg6zbVhq/T5b54Y8CBGcWl/s0r
ByNC4I6DSOv5fZt6ifE9hDqbVs1AeI88TkWXJdKetQVCIgLmvATZHQM59kYlXmMK4o7FO7PmqIn3
9nPRO0uy/vL5SUzc9722v/zYkIq7soXh/uJRbHa1/82+tKe4JqfkUXSqk4M6AbfrB/q31GJquAhf
SNhJgFuu/bUtCsWGcv25WJD2hc3kYJUA3lbgzw1JQmhvDETRRtvbMDUv2TqBPvf5LD6+PgI7AO1x
nYsLSiQEIkCToU9hh2DY6nLWmRMoI8L+VZwIRA9yvHRjVJ/o8m2p1plIHn4aYHbvq7E7zp6BrDMM
5jeoO8edD2qWQyPYh4lcbKKKRPkxomtjZ5ir/FRN5zxKruWS4d4f+JqIIxhF94RKVx3w6hxHEelv
GpgRSeUUf8FgS9mUt9a5EmiC2IkCXvE8dVJS2lCQHEWVU4ZMSNLXR8zaTMwj9i70KcXIWxPZiDIV
1ZJqLaWA0d8D+8lM9PzKmu9npE4CkZKXiLx26EO63i3ito7293dIy2dLBFS27zINYZ7TaRaxOyMA
ZKQm4j5hYDR8y8nnR/nYC7KOnOcKTvGSrCeKv9xbn/Zg9BnIzaE8Ay4NqJwGEZVsAuCPu/qELXff
6t+i2Cxh9aGwogwFrnzNZca86dCDMpTYU1udUQHEl68apZI48wvF0pkQ1FIREoXwfjj3uuND/liE
6cmYNzG2qrolx4HRU6XR9gsu60OLsQbCvsn1QLqWRO365ka667pUaOinCpfgI1UXm5jcZXA0Tf7H
wtx40STwcmwLOrFQaJVv0wYI4jx009DOjAH76t/LBplubBrEHATLaZa3W+h59Z54LvzT3yAd1pPc
lS0cN1ifbvjdQRvXa/mYNm3V/sWzkdT5jaftnXfWhawAhrg26gSRYYbMaS4ozra6KTtxlZH4PO8v
j7ygWTltCqJaMT5phzxJh6Oofrl4jCtoDU6Uc+4Ex9SF5j5WmeH/o8MWWWa71cmaIM6Ipq7L5BXb
3ULNXhi7mdVL5bNnfa6E/Rj/oMN6uHDl1daCrZlE0ZFOveiUnjJ2zw4NXe0Ua8+1Wek+defc5us3
IWMUg167Yom6/kKQSt3MSCeIMkc9vXDFtj0NC4RcjVZrctx9TYVvvPCxmE+vqkXegZDUzJoBLyjS
p+arRxUYUf9hjJVT1y7XPkGwg6cVHkCqRsSrqQO1SKXT1zj7FYbhZFXGOZ3Z2YMlvlNJDqXRIyR/
NnHRi6+dQDE3SFinxpZxXW5HkOC9etO8HRTIJ0ewqLw44VUprS/ylS6YCOUy0l1DPd4lNs+54wLT
2xsuuNRI/aUKNRBmDqx0NDo1FqAbMtQ+zeF9utfengginP2L2y0qCmR85KgoF9JMF/MAP4o+Ko5G
mUmn0JPMgeCZ4PFAeHVF7XEWMH8cY3CWKnCc02mr9HCEmV65YI6wZcBMHj5dvLW9tyUj/PVi7MDQ
a5d+JFnAOXKbQqHkUCB5f+LPMNyb6PzabHEVtEdK7aQ1ZMdIz8mqTppU/eI7hE+jnkAmOCG6ADYK
8KPh2yFOCupnvKY89n7I2FyBOmpRdk7sZIJP4lvYxQUjFV+SqogImmlNnbPTc7SCqnZeCAwdyu02
h1QfocVlfWsLbWPs+fRzWcsHp0myFV+SJ4yaZ89ITZ2IHU0JdYjh3JtmouN8z81kfXm7eiCIHRa3
V/5GDhJNP6LEzL0bc3Vdv2W/sjHloCe9txS6+2Tt0OSP3jqel7Pun7XQcR+zpj+n03OMBbaGRH7A
bTTIZtYWtU28i59HZYdEq/4t+yzcE+ZXzO27Y29dozFON5G1eJGRAlXU1uZvldedzaDFVcIZHBuM
+2g/KaIz3KoEtrQkTinp4vRneqoEFcFPIyf/KYYWqkaKkWpqMSg7NyMWXaEOxBMU867xV3jTZUVO
3dqHDKqzuWZ/9pD8alr45GzIO6M+Y9L4RgBvkCBa3hcWUXdxKBl1exQD91XlcM1S3M9/mp6RMtYO
8WtM35KgKQuRgcXfXWVxBROEqD2aIhcEmSymWXVqPgn0aooLrbgudV7SvFLmYpPFKRzCeuB5O6Nw
wbUrAMCppg/cj6S3TYk92hZwIaTCLcbTryYCu3d/4f98A4uVEvtiU/cuWeLN5flM6/iZ56IBYw5M
eQNGzN/FG/Bbx3ddbYQahnMGCmEF6UTVyiLz/mGs4qp0b6VmcXYyKUBvS+JhHDwqVd9X86PCty5S
Iq/Z3pHQMnViKO6me3Amq2XjSf3NX3Zpt5OKa3CUN9uy4j5IF4WrHEy+ESf6kXf3pXkVEkslttBJ
RD7aY54ARXPoztSqPNggNciuwVOuwpOFKvYU91RQ/RVVgj8U0H6R7N/2zKt8f69rE+1ACxYc6BzX
iz0QIA0OVxiIgzZiG4uOZ6KhNDmHlJLKmEn7VNJu8Y494xeKHHgr/9bDI4AI9RNQyiiTI1QzvvXe
9LtzLe7eT/PVOh0SxIZmkYbCIXI3YxAywUwQVF/QKoE7KpM+Bkx77YPpCdG1uMJDvFgmY2Zk/86G
wsJQXEvasmpbuDs4bZfU1Aud1qUnrg6+6mULgAPJfJDM3QiphBrLIKMDNN92rvGPYR86U6Ct93O0
6BEvTwmi7VsRyYs4AqKlG94I3K2TuaBtGKN/M39Cvr19hFgFNzjlrYIN+MgyP/m9RIMZuQgN2neV
sKTXUKBDJZjUeoUf+rE17hko03EB5/jijBB69k3b00lFpD1oQy4ezP5NLfipLbnwS9X+7gZoM0XM
whu+GCEoywvy76tLDUlu/hIHZHjMtoSnSEBRPgVO1AWAlqAUinjb0T22qI4RLM7HLiJE0F4PuOyO
c5m0Ak1TVnnko53DCiiYiseI+yt0SL75tMwm+umuZzdavFQXx+ydziqi0mrT/C5r8WLilF5EDIbO
IxUc684s/3D8GuyxAe2MHk249IqccGkRylQMQWpSnUO/5668c5r5GN19rg1bNyH9IP5kn+aUPHS8
7vjIk75KO0qyXfDzT0rKIgdHkhjQSV5pTKE2y9LZuP1SRqhGtG92S6KPu4DpU6JMdJ8Y9OE8uaOU
YaLfk0ypWcNC76cwcSHVWWca1CqEkuZJryOzmJbd7Z6NYBvAO2MXN212Rw4d9a5+pxfiu0MntUB5
ta6IA6O3o9MD3xKDdi1Y4kUzl8Ow6DMhK9XRHNiAN9ZuH5ZJueJ3qmPaoauVPPy690Sf/8u8V8wo
EPfgfwImuF2/XWbrUQ7t7xtPcILQkpLhHEFlaRZ94bgQcPPtZYndYVAdsNkKsGpkkhiOFnPgNVaa
QApVzgBZ8b+xOUkX2PJmcV/ET2YzkFabNKnQ5Poze9Az3k9waLnJQf/urGHzpbZiS4sPniBkGk6E
Atm4r5330UvPOwjqP0aHGuWcD9OU+egHvngeRU2sjwEPHrGp4QX0/TA5Z92EuwGuyKB9RU2QYzQE
lKs8+S9k4kNYv5gT7SiowVzt3xfW4jL3j/JhwkldwLMZm7/RSE4KddcGcwFvgT3hmI0jHcEvpYBV
er4x8IIjQUlJMRlAQJaXxZiSWYEoY2ctsvyHzegCNDAGz2FIo/u2TaJZEGtoUkw9jNKEeWfH7DhY
ioGYT70U98KyUXtZ3njhSEM6qDHN3P1xFv6pdDJWoSYu/S3nVKVj8FcHvUFXGT19ZzLeFT2Bn5Nb
LCwFwonvgws3DdOPaxeNJwQfQbGXbj4d7VOa50OIXOuFsE8F7jrrjGe5Yhxz5PvjLp8gNcBkJBwg
HO7CbcmbXyz018akjnD+uWat4z0BMnLmGk1s0rwEYZs/qzIgVzrMs2c3/IWQb2roEEo3oVeJFiAQ
ktbjLquxqLFyhkREpfPDwBrLPwp9yxaJuHxEgBVzrGseboIN+7tT1FwbMg/wuqoFcbdxwPgO9tNw
Dm9NZXAnoKNjGJ1Q8d7gXpYicKKZO7OIsZjV3uOOKFOk1/snRi0UQndgiacWhyVHJ0CCGiRHQjyO
nM2zdS9WR03yU3znYiKV+qHys73fwftUx8c34ZobPjz2RR4XRQk1Q4K5lPQy4Plhgel/7gaaRQK9
6V/O5cLmKhsVn9tk7vVc656hFJR4tFP+s3OqrTPFI8nzCZAPmDUtXAKM/W9Fx4gCz5dZ1V2dXTmV
B/R+Y2ZLnggEe8PgNZl7myNaAHNezsK5LtgkVc8VnMfa9m/X36AY6eCTsETYouDPyVAoo9dx5wci
8zej+mSqUYy42vNKPc095zblg4DMgSxpsbPjQ/KuO79RTw7ne5MKklx67YNJ4602JxIbSu7eAf1B
CjSPHCzTnILdKcMlh5J66RHHNuY0B34CA6PQ7mjrljBDpudWJmmY5k0roJ4nsm1aKohB84Z+Oc3h
C2gyIsw9x76qhl+6RHZ/a6ZNFVuaae2t+Pk/Y3EreBjxkDcxJKFKkCnegGSrsH2LPqKcIuC60Lx1
2hQ5n6F3uIoRAgAvTmlEVzioDe81pblk5xBM22x8qevFLIdkJNFkd7kiwzJMBV046kDjkEbUTXIU
GHcsRvhmmJJa/PA2CHBP62ni/sIl30fQcxjfdBAOsWSXs2k39sIVdZTSFa5EhOBXkNFr+JlOU2pL
Lhx6S3n+b7KF4qVoHYeD06l4tvywUsFZd/p/ddXHB+rsvZxuFuLrqjJp6AEFyXMQvqI3RxYu1HcZ
lgkaiAbb0DDgiCJec2Bc5E8PijUNxnQ6ikhDRL2dgui2xxkZO1/sc69FACsLnXkw9OHhHpsDpz2z
qVsIebp/86Qr2Qh4o81x8x83VX4eDQXaY07BoYFgsS+eu+rTw3RKjsklt0+9ycQ3kzA4QPKN3D5H
NCPgpLZC+Q9o4Vjsf8bK81MKNZDyqOVoHxFI2FZXndl1KhaYFkt+HG8SL14LkMfAdItjFPdnmRsV
Mlxf3Efid6+K7LKOSuxI9b9WX2iZa+QShF2GiX7EIXlJA9usMXi76HHDk51Yzlhs6mAU/rwZqQa/
4m5YG5CYfZFQkJdD2nCFzY9dn5wGR5h9NoowDNBp8rFlt2wKj9lwHwKu16xYRhdR7PVRlARUxetk
up4UTQoLtNVPYBBtZRWpE5DtA+QKwB+I06NjwgKdvSgrQV/iaLhJizG91p2IvqyJTrMFDZ1RtCc3
1va6PVNWrqny4LZXvmZd8+42jos5cUf86xTFPUKrsIscXmd28eGqW8xshkzWw5g8x1OF6rglY6EP
YWi94rjWh5R2z4e6tKBnlQRvL5cPnUPoD4IVaLs+xbHTF2nTEhLRIsVNw/5c4DqobFqlkyX20lSD
qxvSeBimhY4F7Sg0abuZ9TZfrOMtHkOJ2pIZGfP/UjmxhFBo+Tii/u4+qZQnvdZvLuMGEJhMtUZk
KBcJlTtYqRdwRDcAHRek8X1Y94ENs3RRLal4MMw9IbtvEG0PRqPT4Yj7kKj+LLYrZaxxLjjz4cW4
4YNnGhiiDULZcUJZGfCYz8Merrfey2ejx4YDdfT37vQCvQg8lXSPWDPsOs+SBNqAUiOTTXxuq9Hl
N7kKaFSyAJgqDPztCGYvsihal1pDnpb+cl76MlrCy+8k9rQDd6xDof2JckFRgv4/OwHOmov3bJ27
YEhvwrC+sAiMpO/fL7Ef6HwsVtQNoFL4858OPvfPnR2X1lR77cdGD+0TJa5XTu72acxCK0OI7iax
HXOrhbnQcFCbu8DRimc5zEDUwo4RyxBDzdb9UGK1dee/lEj4amRzK6Fn8A9OFXTmciYqEKZf7Vll
BjkJKp4MotSqwtXIpkjANS+rpfp8XduMPa+zAu87ePKXgItk5VyhNjEBFVdENadfoH0Dx9vTrLUf
1wBtaCaRp++t73ioW8IWefkj1T+AHpWWqXH6qgjbXpPat7G8coAx1S82JuuvasepKrkclYMKwu4+
mIw+SLyOVyEvvCyfhZNd/5Xk/y9S0d2y16qbMBDHfY0YzF/OI2m6ekQ8dOCn8mb/KjiihXkIK8nh
GwounfoNE0QJ4W1eL/RWVFpaLCESK6vQCcZcpCim1q5mJguSZWT4Bsh7vvG/fJMf+2D4Uaz6/GTC
J8Z5GMhwzPBl81+XRoPFNJFwgYGIZvMA5H+6cu8ABuTuLyO1pY2pBqu8AVTyQQknWa7qnyqN1o/B
AeLhBcK0Up2YAWw8FA+7OGBp5ztsx63N/bU1VwQf+tK0nAlFD6rNzXMlPS+dOtLnZhYymrx3ra8y
Tmtju1IE3rcB+FbFDov01Npl22nZJRNda6/RnVEaX4vlL/bp8iLlM3g1+zC+lzWfe6Cp1rI1OaAS
Vp7FH6Z149PY1iQC1T/LlJ3uABOXocsJuVbzxq1aDU1sfv7H7W5n2I5cw6N7bR7KrJB03NPfC0ge
bh1+M26+J4VssRV2jfeWd7RSfVMdBItdYxzLpvDiS7L2xA+dySHAnYABD4H5fvkTLyOohhb/AHXN
9zbfuSKT3HXRN1/ML+QubnYG7vmQU3NXAra4xEDK6kz0bi3Jj65utCVA84+O0Y2hPHPFle8w+vwA
jHXln++Gg71oVdIK1MwgH8opprLASuEQhVCWdDb+Xc6J/jkvBurVkZeMQpBv9aEEkYNFW11yfoFZ
h5Qv5tsPLQYTNF0OzftwBUUbezLwWaxBe3zD3dePbP8jMco3DlB4MFmC1R8+OTpXc7AtbzA2HwwX
IPceYcCJuv5Y+X1jrImnSs1Y1y1F6G/PraITTN8hhf4ZvBjVe9bE6hv4HiKY7hPqYa9xJ6XFfOl+
QQEN1WOcBefqbIDcjlZped6RBPThAEmoTz85pvbhDER1unBJs4ou2iuHSE5rhaVdmBxD7ovYvbqM
efSp9rYEMhJjYv0txRK2/KBT3xDY7USsftc8W8b4BvXQ4KCTwd+b9vgaLo5WVCrknG3mrHwi6QIH
82aSw4+/WkrlEHz+kJ84oi9DyjMKwcfKXdqFSdmtrvoJ5zJxmALipQ+NhmLbQLqiIiGee7abTDSY
fhrrFWHH0KI/GjSIgzNhsU4bevfvgUncZcnc0GIEplCmMifbXp3E5uEllpR+Rr8/uDboqSYPuZo6
cvmB1zOQiyRtDS+cfV9cVv9aM6wbnPcxmxzHTuWFX22OkLDTqNWaAqtX0t9mKakJHUvKQ4wP+UYW
UfmLqjgppjuNYWEmybpqbdvgJ21j7018PIFuHHRjvbLoFACKWR44ZCzAbdYs3whoviiBmZsFt8sj
pJ63efbvQGiSxtipyWhqbpivrQwDS3RK2mkL80kGU/mdX5DMWartYl7VZ52WeU76buP5u+FuSsn3
yCbdLkZZoMDVFOCF9si8C4Lnueljo89gXHw9dWMkf5yMOdDXiY7O3esxPkoQzWVNKfUMJIcBzrES
lmZ5/XAzhMGee4r6wHVroHGQqzyML9JabEc5CJe3yofjzaO+2S7/Z0aNMuUT08mk1CqIrz6BrKlB
A7NV5XnWSvUMjxn8LHrunB16TXw3an7ov0bYsHVVDQ67nKT3QeA0b8a8Xpzv81St0p3fm6u/gzD8
+OqpXhW2TGc31+gVcNJDy6cLoOGIS05CtVh2BXZ+VdJQ7YqP8GcmKH0+lccJmgYbz8W5win7GOfL
cqJjQ+tgA1fhYRllcPDQJceGwnJFyZLLtvUkknzrP6x3TcuntK/cuctKP1B6LPnBi8KKgTkHslq1
SytNxJq8GRkZY9/942iCXTw0gmKFl3Pta2h7A7r5hrZDDXyzsq9mUFFoyDDmvFeBrOBoL9fV6K1z
z04o7fPmrj1KL15DekuTi97MoeKNwZvnAF8waRj2Iek0tx9UV9J6xDS2GidEYpu+adtd/6+fXePY
QxLSQ+ohoY38v80vDfwWIt//o4pSR3Mz7ISzL7y5hYgw8QoK4LEeBN+SIonuNL/dWHQz+D46UxoE
CLBnl9yn5WiRD1phvHSojGwFVu3DNgg6YP4yFRrJc69nTnb9JNuudpfU1PWLMVfMjkq8+wA1cnVD
BdSxMwVGtK1fW/oD3eZ6umQi6DzRAQ5i5kQiFiLzI9hDMi/h3pyWArAkTml4Azpqcwrzq0YBDS86
cFlkxi1B43t4s2+NViKkmw82EkNoudNVOlkMQcFYQQzlt2ptxEzBXNDFOcNIm6QEpLYjyWTfQdyJ
vGpO76GDakFrKrFXxvoddhQvdCf2lvl5T7haJNv/ZNJY2HxZnMhWRt5Ab+6YOJRCfvDcXpYu3PuB
hzLJzD0Qc2plplew/Aje5+XC9f0HtXyHv2lE1LUrawc2829LMn5ZD+51yUInOx7uZCyGiNjEHVVk
FRCqm297uUvbV3zOOP7xzWeisLtH9H6Zfv7FRE2lhFij0wnRI9M4wOUIwK2QsBmwIsXFEvrBrjCR
BJTMd064qdb7agQvAEJF5qA6UTCfXOkKkTKGlStjF1LyKGBhJe0vKStFnBP7oLApdbNZDKLIouVr
aO8xGZAG1uJb4eyK+rQcb1rI2KCpnjaJ32VaJRGPz1VkWmIJWlvOEsg3MPqje6/uJ43Tp67Kmd04
BaJ8dDSorCZE7WHs6dQtQ0UDpmcVL7gObnshLIRJnBguPNqW4QEO3Ba9ZSq0BUCoZfF7sV4EgpVg
0163bk8UEnU6ZrxtuhUZ6nwZtbr67rcqdqDEDcrTURs0+Z5WpSRbmKorRxbkzCGbx2x6VXaAS2m9
FohPV2WCQa59FZxT2gEqAj0DDgawBs8+mz8onRPylvnX8YtXjlZXyGV11J2NCw70M6J0yYa5qu91
pC6eRjYTpkH2+n62tqZsUPx1mBXe2fe6HEXf7A4ersnXO45DL7vjDmSf2ZZUqOQ6Qn7J/Wtgo2UG
BjetAE/bsDfKKtO0VnsCp3++OjIiYKm90aKwXb28olVt7Ygn2yCk2ijff5A9tDb/e5WqTtW4oXMs
eh79Gsx59CBPc3DcJIk68Dzxr6tH/To5qzCDo6031T9BjsdFYphhWRIeqGOEVo0Jh/IaMecCE5oN
O4FIiuIdVhFDlJ8Fkcaov4uurDas9/h/o/xDerYlY5WTaOnDdRqnq9FLb6GYOHVjj7Wocbfxl/b/
lKyyGYMJ5ioYyGccWZsU8g+KucjlzT+0SokmVKUiYy0JCES2zEkeKko2fTjunfI2A2lXLDF2T/nR
/lLbXSr9n4I06GSb6me5jjZo05tMGkMQijS1HPqVIuVjSCxP7YRJoJuM+CEDW9++whHismfu7UVe
mGfdC+YUsr7FEUmoAfi2th3spH4S0zA5F/Pq5D7xXpsSgJ0micMKX/GYjco5Uw8ElhpmgUfa9FHK
tmYhorBj2rawVI6pm4K6pnGNeyDLbGmlM1DPGTAztO9td0aUzlGG3Bns/gj607aywMsakYZXYj8/
tFKU8ryQpt7eGxPP1eSrRExfQGeqgl98Ca9QaXHZFWtwHwX0mytXTHUFTXr3NDZzW5rQAxuDYYPH
E2BcPwItIwehHFqMXJmDbvma+IsKuRleJeOtYgznPWeD0uRM3Y2bgGieDMJrAvfiLHooIz158pAS
nA5woZjBil33RASOErGzUzMLQCnRpvN8qsM8mS85o7rWs6ZqOVQz/8d5MumOz5dqTByEoA1Q5lga
O+1i/QI+wGZhUBAENAlHbokJ1P2C/8fV0eFPbjISJRD6yA5X6AE7mmxXUhy3BIV7YGhufQ2i5xdJ
lXthwWl4yMIXPVnz40L0RvBh9PNeKE7vcb4SvDR2y1wK2TlJQFnPedWhp7TKCepFBkcr8/eMptg/
aI250U2+vg8LTvn9YMyG4yfZp6SgiWCtDc4lsR525lXou7cUheFtd8d8CNxmXvu0XdNXpjlijOlI
O1u9JJKj+10J6cIcZiLiSfoEug5kq9QpkzfXvj4g/4qb/kjmkkPrwRimqJbckPfGDLFg/kmyZ6ZB
MtMGO+FSEihRXWtl121xQO7fglxSObrH1QVssrPei9VRi+9jFBhHRQv3k1Emkecx2ao7FtC3SK3/
P+ApE4bHT+GbaKgJUQlLvwfgOHY9p/xgoamP7RqhXj3TGR/eGypV9j/pxPlfO8BV4hPnREUTpww8
HAh86sR9P7oAhAlmdqViENYEMHJTZO4IcocpYJUCQdL0n9y+CeuSGPI+oVKVTFNg0qbmDceQFlDg
Uq4TCcc66NeACnlEMNCTW2tpZiUi1OZ9zvC7AEnXy1SYINfRZxdFcrUNVQvN4gQM1hx/GCzoN8l0
0NI/pGMwnL0+L28iFiizFBdKZ3vG1aufq/T03SLXhEWdNvxjQu7OISB9C+ll66w5brmndnxeQAVx
bl8nwYW/A7j2PzYX/bshuiEposU0PmtUh7eYcnp6MAarZSLcqVD2lTxgByZbrGynn4/WtRexiYeQ
SJeCCxw6hv/jQNEwgUW8Is65zTkOwEAPQOWS0tjylNlHgnjQoVLlNs70fd7d/XPU3cAeizNQ68F+
Gqzm8Cam5WBlP714pkbSCfmzo5E4CH2bRxHbSfH83+8Wlpa+1Wwtt0JlxZX+oS0JAVuTj1XLJxWU
xEFD0xE7LWK+H1n4MCFM5gw5lwnckcyR7MUKYbGQouQhaowQWMSdMz5KN2GxoWOhmJEC6l2RngbS
EfLptGpOjtV9Dxf68gI0jdTpoj6esM+t0hjVIWHYkpFkarwX3J85AijzWRFJ7zPi86WpiZc83w76
Y2cH14vWquw63LJ2d7caMjKCFJs1MAfTPntFZkb8IeTBZn9gZ11MkiKERiHt8gGRnnHkCp2+ZkWp
T/CK5FzzfXAuiRRiOzQ+7E8GIKrGOZCCiCqn/6rEMKAtaGSPIWDcAH9A/zb3rdAWAmYzBIJhpEPY
6QrEqlqfa1SEb+ZVyHct6iQ/lmH9oBHnOGbIG2QziOL+xn9CQ7pVk0zTtUUrEJ4oajWQFmYhG94Q
7Y8KqvWDawD5X24Mu/1yjxm7ImsI+k7nykvNkkhOeaChZnJu6hALrGk6tIgyWNENASXUEUgICfL7
ET6KwYBda5OLjI7gV69e++Ikrjf7D6aKy7gLcI0aO1GGbyoC+p9gMXaFVS9xULbH+bSL1pn63aQk
I0PqzHGKX1CbaYhC1JLtReLGLqYqiRqfxM0DHjlQxy4RhpJX2wst2S2By8VFtJJ5fz7Dz87GPW6L
2t4b1Ti9i8k0FgkKbuW1Qwo9Yc0fXClJNsWDuy1+vso3JIogCm4g4OS425A4pg91mJVf8g2GTj5u
y2GJ2O9+SQ7RxKbuRjGqimNs7eZj+WBrxGJnWEN150cRoLutgb3yKgv32jSaIq1idq3VsX7Ji9FV
Uf/I2379feCKw15WnlDmaCHdBTREcI6pqeT6xNv6/35Pd4BuLPw1/ARGPU1bLtisHzsWGbzPaU7o
RONRo2SxsCWTR2DByPwIj8Skkn2U/DOUxOJ2Qz/Dr9niIGhKis/1Ypox4RrakkapCWqWwtvkGMLS
vKtj8PT6V2QBM4FqNnPQnZJBigLVWwo0k59+sSRXCyv57vijabGo/trtTjeCIKRPiJ0TTids4qkM
HBM3A8Dgcj5jj6TwkUfOtxPuF3LzRXRqQsGILGiqR/fUmCHWVDbFIYdh7aklIFQ95WWQOz4AwAOP
X9bGNrbmPiOXo3BMG0h5NuS4ukC1DNJb7lOb6YF+Y+8xj8ch77I/r5UkMFsSrRYz/nmFUXnq2gWC
ggHz9BBh/UUe8XALzMa19v2EeCjQai45oUgYEGSC6VZ3V+bk0EcdjAt3rFSE6nZ/aG01TTh+3XIx
DdtEbSDVt7KmaDt3E548ELjmq5lMSkcSm7Q9Io+yRxYzifyZnZG5o5oEaeaJh9y53Atp3UbTVgQM
o8RmjP/YzqnlG6iALldW+uOLdwMqiARnX51hqdcVrjXfqQBcYWjjndSCs6DjUPCzvj03y6E3nOHJ
A2tCov0oc3L7ZGYlXCk8xBQynENTL8S7EHUmbcqBT64C1BKmaCyAcIsTYVSECR4wv4DLP7CwHQr2
DjB7yuGwNvbwFk+dtlMXmVvb6Z6DyJBHL4UFkTgPuqwjavphbxtbdgFjN3JlcHlDBOptThh9v1mx
syVuJqqoMLZbTirZdUCc8odDd2/NSb50HE/E0yvL/ZCGuD1qdJG52rEU/ATwMBQ3oUcu+ApdA7gY
x2C9Nxz4hjD/f32b6lyqV1rGoq78iIrwselU1TjtBaus23ZgsjbJpP46msjYriDAc2nMxwDXGyB1
ZdmAMI1BCAd7wPEALhg7eU3tqG3qz2PeGMhy8RPG57P/aa1QhL2HyL6wV3o/3T7STxtTSH01ReGU
J4bjSdseXKFYD+m319YwUanoQmYsLyuAfMBtnkI5URK03ReT7pUMeH3b9cdKivcz2Ya3O0ZI6B6G
HCZIiJMbWX1VagsIOypkFO/WTfpHY/4E7I5NQGoK52UDxjE4uDSef1R5FGndwNqsq2fY6iChAwRe
KqQgVjFSPi+N2z4QRfFgE4i3jIa/xv2GYRmHN3RhjNtYtQ4emyKIBfWX281bE8R1ZP3pNlqtZtKg
IMopxZM3d1aQLztO4cDl3Czaqu8lxtpyDzGIJcj/ATC8WpIKJUmZTl0IQ9BskXwZrsaZNC+k55CD
lmQbmn5BKkyasMsogx+OUwcQbAk7KdMqSczVO1p3or5qc1oddUEaYp9B7T1vN2/lA8ibxEbY+7yE
KDRaEQml08YyqjAE1hA/opKCdYB8oSh0nb+ZLpZ5WCHjOcQVqUuGd3idCtlkwA3hwfqr354XAIXP
GLE7WE72YgxSp54EM3Yaz4viQ6WDgZ8d9AxxCeIIGU/w1xCGUB9BwRPycKaWzF68Zb5NN3Vy3eLv
iK0GUSRU3PQBESRZnDBOuqYFmEJahig8dvrGrLOurXGrhzyR4PY6lQNRGmvAs9ZHl+IOR7nkuwrP
rcYGGetDyXARLPbvb6NffnTPZyadzD8B8A4jk1/s4UeQJiA4zAMJXy0lXk/BkcGEhzLKbekjZPqB
+T0W6DjGknMwGAjLmtntFu1mZscojQ2b3Ur7hQUwDLBWK/FEiqD6KsivLQMrwD8nZ2MrIQQEugAe
qHCLQrbH5uTt8A4Zp7I2bvdZ2bxNvQ5zQmb2BlEk6SjcUYE/Jps+cVYuc/1tKVLna+ATqdaLYtmn
p0vZuevUGwlC8879mmcGgPazhgyGR3e88Xc69l8Z0HVp12CIlZ1KHnFRTmAHxTeiq4B1E9mE60am
67a3JHdx3HAbShNx6CJmwRToK+fEsa6b95JiPcsSlZ2LPJfseb6dTlc2xiI6y/Tm1z7w+WyCdcMw
rJ8q685m5ckW1rBabFaTUXZnYDFCmh9L3s78ZPwjlJPMANM3Pm6Ow4leYSIPfWhuwX7Mfd3NDGqB
cMTAfhOLIWWM+SRf38+0YhE5aNvoR2novg2TGATo1m4JY5ZSFA0aTCOt8LRks6EjkIhe0oH/vL4p
nRh0NEB73otmHlu2LRV7cdxRTWI3203ECDxxgoE0/CrQ9MYCVKKdl8oFX/qp8dOnKSkcBaXJw3va
NNr9XmFT8k6GEf1ZzYKyY4JPuQ0Y7k9CWOBM9JGF9CV/kr442Cc102BsOYJhLUSUOZR1FmxO6thT
avTuF9IJUuGY2OYYGjduKkbOWVuGQjbTjTc0+j7jwIYIhVi/teQihsYl71lRt/T+X79/MUGlIRh+
OKgys1+aqpwrUv/HtLctJUKAaHndtbqH5AG1Ff+fnW/4/pBz9CRHztn9Z8yF5K4mzbczYCP7FIzB
u1SE/1jJz3KNdkxRTS6gI+wOgjcTirNgwMjo7+WBATVZLxDpvvWbXJSR/hh9DklALWEn91rWqYup
/UYMo37/nDiK8/aZKqHshbpgjAh5w7jkY1urgwDynqkjSYa/yyIuFOPQeZOWeVIM0G1VZyoVf0EN
+wZfc4Fs7KqAkVXva9EyEDYlKDaeW9nDsee54E8TnmTpUR9n+zxl3bPKbvS1tsxi2TFLdB9Udd+/
8KxLVsUFqDLv8ww8as26TC8qvRIhPDA7Vq1+8kpn2zXmpnBNA94RgP/3p913CfI0W+ZNqCpiaJYf
NOeQtw+JGpNjnCib0TRnyS8XqtPyahWtYoZdwx58e/33Gv9ukMTqbzESlzoTTKRtKT5fz5shAGrS
/gtrQgDWQMpgn60ML1t5Rk+Dkyfvwo+j8EvEOn0I34Lux7mKCrdqgsmDkMnqvDGx5QeUyNUQFijx
02mhPSp05b6lB/OBMqxnQ0Ikj7ro9dLKyUihiDGNnDUct+8MG1KTKEbLdsC6MSULgw0CvEwK9lg7
YTf+vrRgJcNaTgYRtqQ6EX5dJ5c+Xrjh2EiknTdfSZ4ipdtXWWPoDcJgz/VtGH0zBJAA1wwWbuPV
lDwm7vEitN/05TtonSnRqTnAInNlC/PhVPqo4npDyk5b7cOpa+a89o/p6TAvzrUBs0jjs0/cUoxu
B1kD0294qnSv+bEkerK08ECG7HyWMWM6Vcrz0oCYWWKtNkYtjuvVoqOdMqvshKYrsSBvhvcqovnl
iBpAJPDE/chYS0OcbMK5xDwbm1Ga53CBPNxgBMMsSQQ5XJIWW1Tnfv1Xl0NpLedy05Pz9csdwu3J
owSEXtSbV5w4ZIHqDTkxHMldVzetq00hVdD5L/Gaoco4/KMu/JeTqoi0X6nT01m0EIegxdevGDD8
b7Mrc4e4L6HdJaSOqe+Plc/yvigbcpp75Qo37ZCuonSIVH/CeGUIH2zvIxI9TMKa+lnveKzFXRx1
e2rWrWhSprXi7UPyviY8scjJLJZ0sYzq07Bd6iob4khJ/ePpRsXHWt7kipFJU7TMRQXC4szK9VYi
fDoL9yMDPM1q/+h7k8y/5jtxoP5jopENp/MreKRlT/M2tMfYnpsXK/6+C7L3ZScATLblWHobX2s9
EQQbfzzKJdE6GrvfgsD1vbDayk+gejHHm6kyIcYr4qE+6flaC2Hy12O376h0xzDkiM2vIWyKMdLE
kvra7Kc/z4jFEY7dOjev5vl7waW2CtDNuN/W785XO11NKhDA9uI8Zygd6zxCRH4bWKA6L2ClYQnG
d4DQfpewwyLhH09LDsNMoGaVMjDwWOK93UmPfGRSJiJz68mQTXOv8ZL4QC5TZe9evoAvk1hEauE4
nSDWkbk2346pyw6a0hT4pah6LKJXlTkUdq9VZ4ZOw20R42BBzpAgA8Ay6QOPijPfhO6wf3V2Tet+
a/yHL6ypo5MrvThl3pmGtcU5sRsAMP0+gvOc6ZAorPDhHXdNkl7fwXD3UI3U6vKBwlZG2utWc7Q3
QM7DWf4cvupIOpBFgYlmloFbB2odezi4SuniHwueMMya0C3+iKQcySGOvczWgbUOev7UE58gcBbN
E/nwS7Vk1OzcvItWWktq2pqMDZ5rUTSqQZd4SmItuFNh8c64PuuYlIhA5XU3xA9GYVJfnZsRxL7x
qqJImHDeONNoSiJuGhYR1FTXvwPAOm/2m712XXLOTJezfDvAU71zfgIyjgXvMlJSXr59nYgdQzo5
I6hxsbcnRhNA22T/4vtEMzmMkym0+m/K/0c4xeKs5VeNbiwpsYtDAQlnDQILtD/7ELe/y2bDOkqC
b03f0DTYrC8Qfg03EGTy2V6sosfB/br5TkZ0GDF/KsW952Zt0Qxu490htP9IoT/0NWm8UXYcELLW
3C2tdyk07C+AkxHolN/iawIjLJ+EsO19KNsnXrTbTR1NIYwJw7mPW/gcaIFn4BGGnQPPljcIr8Is
RgrX6yweTKH9mhesn7Hs8qIC8axP8YDpDfwJtKPAayS7saT3iEG0koPC9XoFu2IVknqp8miFvrs8
xCDNjdxEKdbX111vm0kX9iOghQhRaXdMUi2csKhtcOvqIssdeVDYxjcbPX7bz5Ze+a3x+secW19W
mIwin++Cd4a9iM6pQTSczBSQzSeYCD52tlyhG4EkShGab4u6cfeogEk9uNj9lAdtggaRXh8/1XJv
3BxDQCz8wPQBAA/HBLjaiaYw7XFzbtRoR4bqSduIcjBK00RkSXrLvdhBSmN2PhJ9mE6z1nsGcKJ9
cxdrBNDccSF/7sHms2JXP6PAC5xU7997tlCecQT9wqIyIM+kJqm51i5Dc5lAn/4hCBQtnRApKirg
24qocdrWepuXoR1/tmYxjCw9pgT0vui1mrJDRawy8OZoBt9f5K1IHp5G9PzeDzUmQdx1ffcQkw/V
PkqNESavtNSw9JAX8a7qfzsZVmF6tboHS7rhsVfaAam9/RKqI72f+E85vi2uibd98eQBl/bb3y14
4hKv+DdI7GDZmRmbLSA6nQvMv2tVrijgdCIqEeLqvFw1LimxjKp/Sk/uMFKsJg3GafnoEWk6eyLa
h1iw+Ye3q3U/gH0sY4dPtnT/br0MRTmPhEx1sb0ffSWE9oiX4w7KKN0WlV1KYdEoBLkWaeiHAm4j
GWpRqhjUzWE97OZPUDEvvK20D8AW57FasTsV1XfKWwATWQUIWRLKYVk/RSR88CjBoEOtHDObGRMp
Ar4uWw0KBkPDTuIg2jQMJPWzrmJvdl/MSqNmkJMG54d29tS+6f4fH8gzdgDza5EhRh5nwtvoQST0
BwqphFFnzAdlJVoWIhq1yjJwocuz7oMecIvN7N2g7Fp3ghMeGv/JbHMnEBSqoOoCr6S24pD1CkLh
8mF4gVIxadCeeNheBOAk5q02Ea/FbPYIRs6saqtVUkN0hhUlkudvAMXHMNBSFfsLjp4ZmkW7KQsC
gP5Sfvgin89hFUm1uhzF7R5WtZ9OVMdDSlRG6YPjewZySpbMVyFgvSnGpBCS5ud/+I7glCp2Nqp/
48716X4HUos5GUEZhgNwsuF2Id33S1k1aPVoCrLDpQdjRS+QLOHctbIrtxG+gKT9eXm/7u62vpCg
HzJdvyWT3cfxnLJSvxUvro3SBA8XkfyOFQGeKSfkIEBW/QUxiZamqr+8r7hEktQXYjx2hWk80XUX
czyP20ypsCFLOrvu7waDeKD1MP51G4+EDcMD7vgtEd9Lu0pHUNXVN4sb5AiBoLh/hd2/4myf3F10
6g6GgJqPbzQ9FTzUGIFWCSUL1cEznp3+UI0fUEk+MdMrVVWidWqhy1NmXeeQIwxoo17BWYeUCFtr
1c6DsKFjnkQgULxd/EIlatp/2rquFkVbuOq72X8a0SetmZKqpPTBIOtJmez2VY45uvh6blZb5Wjd
JWx/KIippfg50K4LsyZHczQwB1JFJNrb0IzV3I/068abqHllzsYQHv8Sd4MYaRVkg0R5ysXsmpFb
D2thS4yDbYPbMUG82fiPuEBxrVnK70OxZYDNE/xn5QQK8i1gm8kh2dLhz3cFpXQoeb7/mzks7Ko/
btrJbnKKRRlmRXNTBBMuWWlF1RwZC4BPawSO0gLaF6wVoxfCbqfyT79+nOlt4o6THlm69bzHNbis
dsj3xIAvESMGqYOcH6ftNor0qaRvV6hZ/D6t80sUuqxQumTdxrnMv39S8hE7YMyxMaQCc8sfQ2YI
XiEee/0Q2q2gYa8xfnZO7N8HDXYqT3uJFfATAGUEWQCNs5rpswelqpGL5QusVZ1mzdrX3ykl+z35
6Vez+8342gFrHYqe21gAeTFSgwFWtjctZefNvNxayq12T9GLjXx42IyF9qV3qBDG59o0Zer70H92
jrFDD779NRrfcob1DuQ1j6z/wB6IXjVEOlN9+QLqtDQ4dskqcztXuxygBOFqVy+EK1DL9Fe8vtvS
5x0D4M+vDLnuB9WgGZ7j8GIUXZqhlaVGw1rpv3NoQclTzxobLtJQOtYv2gmhdozI6eno/uEepyfA
e17Y9E4JuWtg6hOnhfcZTb2VItp/HhRcydr2NBvtZcBT4V3K8yNh6lmZe71QyeRKnhC3T51+tKgX
k43cUJHLkW1+tUIOSbUOtqB3XynSAq96L2zPr3s1xKTMXGyCQcWCPwUDaTclnZLYcVDYJ8mIZDTo
7yVZMWwt7XZlY9gB9Tk3fgVKfbZMk0uIC7JQXEuIR9NytK6cHxgq9jl03U/ZsmDp9QJRv0RXAc56
uIJ0okB5B3NiczNDrRU7aIUwLXa6zY79/0KmIf88i0SV+IUlDNTgTeajppd/PM47XCGoxylgY9lA
kRGrG894rYhFea7LK1HCfL4/G8OaJfmOZTa5wekNJQgVFvcndZxZf5BU2LSouDDkuVWcWuXalFUb
Lx6iHEo6f1RWwgvbJSF/bFtCKEtxYc5uYMMUS3pe5FZWysBOXCRrOXYCIcAurrrlUIdQ3hzWt8S1
wi75otgFWqbMyiSsLPEHgcGECY5HME3FqvV1wvlw6qba95JxQjZDx5QvFbCrohfdfhr71YXSVYMc
TRCIoAqXBYFMTS/YlE3r4BiO0VehJDnot2WvXzF7kAtsK6HNnVaVSl2Af8adYNRVqbi4hGyXEVzv
EgOpOCdx9CBlau50ueUuSca/FsTRcEmw6WLt/kcXLP8jv2q8WrP+sdzgKk0kgKIFo/r8vTtxEyrd
YA76RidNEC/3f3l0riZxGoX7DLf1YKI9qVRiCK9i598Uv9ipZgWUn+vXqQw950D6fNrS+E8YrCkY
zSeHLn6ubBY0ysnD49Iw0gpg9tEk2/fo4vwTQ2Poy1s1JLGPlDnLwLz5TxlFu1ASQjywTmKmEGS2
pmV53AlZIYjeDSUjckzxfNYK1keX8L9tH1qr+zAZm548TgOO7WNHEIxMz+MG1D+udZbhekVuhGUE
LooT89gq3M6ZVRxVLmViNiF4iSZnB5DgzTZ1/3eBrBS0fDgIMtNjb30rdyjfvGPJtArN8C68J9iw
k8pEdxkW4U7ICXrfJ1rWSqRzIg5Wv4dYCUw7Uv5FvUXknUPCdBzztM7+Np6jGONMR9WqDGEP3gYQ
4Xq+6LmePdvFt1AxikbOKIhTgUICfoXSWMco/TaRFEvCvJsUeIQWB0nuryfcaX35rRHkKHTqer82
GAuHwNbj9/8L/UsxuXiMFYwULwlJzhazXyNFF91PzrzAXjvwDBaeRbBZ3sBaorwrmgcZ5JeD/jVU
e/XlMrbv6hOj2totyL4eSWfD4Zf9HbQNFcpJcu/bGNSgJrFBN3V9Id/a/cP9XaLn/WghQ+QZIppL
2jFH87se84nGtKfCQxP+JjbzaGOzA6CmNds2aCYiXYj1AhH7F7rh2ANBXcxxLbQAZ0eSB3Useh5M
XIVWrkztsyOdGsVolS46B5+zmhWSeMHI40vy9Ypuzfgn5bIHca4hAyeP2vie9I7DyKgUjgmW0eeC
7re+RhI6chU7qglFenQqWtPnpT5e56RmOEf3ZZ+IsuwQjD490STFVRsALiFpVSwSSIhs4s83TR+y
Efh+c67UNyLrF+c+pmpAtmnAOfsmu4Hc6QjqrBZE17C0/sTK6BnoA55AgQhqgNId/SVjMWDqs9hG
rWZBO9XjsQgpQrdtJOdLqX+cztgaa72BMnWgcky6Jtrdgfv3GNn/oIHx3cDQn6Sjcd2xvtcxR8qd
2ptSNHUZWZBMklcWhdDS30ba/7IeqlsnlYS7O+l6QHbLeF0G/Dg71lu7PRuEK0/hcQ+chOTTgx3Q
P0oRwcZwcJq90pLGnZDh3W7v91uB1snRfQWhbx2HrfR6xDZw97PQjJ3MiOC/O3p6AW0NI5maAPvF
jOcmpH3Np5o+ZqQgsG2axx99+FCXsk5bs0v5kdoyGmmK+vmizO3zomDIPZ9oo0929umHAKtVziZZ
eSV696Lti0JBhreoM9hUmGCd44cszlxn7uuZkp0Mlv7GcgLvGjUu+0vWk4HrV84utyulnRP3c8zb
7QWdfnf1KMMDDudaJeHAgaTXjEUCe+sBkPQlV6sy6btEDH82D5N+nEbghZZ63AADnqysmUpkoRL6
qypMUvbaHB0TyMXQMbijhiCqJwv/sBYfxBIQdWlmrnpzfoKnWzYbWWdao6VLDR5P5A5gTyi8vi9T
Nyx2dxH5C3PgAdy0bAqwhJKCnuID8RRJXvvLByJWXLiAwDInrcs6eQN1ue+vFb2sfkwbJCCo7CnJ
a0CuInmrNBaFYXco9lfqzdUD7h5HmD822MzjVDyZ5FqEGBrc3kl8DSl0HafmpwP8WL/1V1vy9h9J
BoKoPrh4cuoxpwsRmBQsfp6kg9FxDBXbF+53OrlT0+ut2DgSbrc0l/6B64mGad7M5l/ucj3Xb9mx
qy9mRjoVqsCoEwEzbPV4nDMKFnF919kjfjW5Fbsn5kykjsfuaHCqZ3T7NmKbGVTA1yIsMaSR+6nD
+idEUClIlC6Jce/VmQrpm4r/vvzCenGGq95HNogD8or7QdFpL6u5M0NQivzYXJOuoAy/DMPpFqgt
vZW6M2QJQ3/tqgwkUYcav+o6ebNYnbpt/6ACQ/m/6N7ypzcEP+rruL9Re3VJnTb1BASGtwrzQN32
F6UEZvhNrtQHFFIWZZFfN+xVFVX/DTTnnxKihDZ+mpdzBltTaqbGR/IqRri6xIYBSC3yhlJEnVyv
ajT5lMv7IfIidj3bNzEsN1iqnKa0HjXLFIs5gXf5PJoSvEb3WlrJ+0AyLpll+siE/02hjgO8300Y
sXTZGe0ePzrc0oAVgcaK11A5UG8DgREob2L8B943PxTdOcTjbFjFJF9yZ4WnuIDzOileHomAnuGZ
W8MEKrPUQo3Gm89MHQwZoKOmHeW9ri/CubbJgd4qnEfdUfnVA0oJKYB970e1iurAUsGzPEKqaCIE
LPqbRaHIFKd4NR5Uo7xf+Pf7ZyjgU7xu15keN00Mntw3i+nx9bUFFJsuGmNum6V/QAnZCJDBuEG8
B0/uZYTrYODMypim19jxmSujvqm646d5j5ZcUXTFnkg5ATLJdqjJlCEKrTp98GxdaMQJ9b8mgTjT
5LEoaIjWAPJ+KII70QkjlnNvT10lDm9LlBKkAY7j3/kMJ2jpswjaylGKQsaPwL+uU65zkMSXeUhC
tetq7E3XTRMHxlYyHUFy6lUihLP7LZMZ+sr0lk/85OzsmYR0t8vAPMJybZOZC8IqbI5da5roaol/
0ko5DIM1d00w6P9CbA6ReBWdzPlofJ1RKtr+2EIzhwqNhsCao5YasOnqgysLWns8MMP9dubq45Cq
qNjMjFtZbsYzIqlcP7H602b6zeyH/t8SFCTbw17PfPG+5r+8b0K+FiWd27MmJ6wFl2ZTo2dCAzWZ
8im2xtolYURGvYNpQM+jCEn73EgFoIcYXikLY8KfMndrcl4fA9UmiLDkr6CMSixZ8Q7qUGOCbrv0
79y/+X6onsNk9ME/m36K+KQ+ZIcAM+RKYjcoGVRqKpiUkBk7O0SoBnUgF5BhIpx0P+9zyqiSAkjn
Hq7Vr29u/6K/AQPALqsVgKQvPePGYWzy+IlUi4SQqJ7M374j0v3a+fw1J7H/SxDtCTZsxBbp4TZW
H0pvPc1j4zMs09srMoqqpp1CBa9ZJoDewlIjc/rHAv0K+dg1aaraxEcP17fnBaQwIhDKDO5gb54l
xSrrAqttlMdsffdq88EPmgJlvZ/y8IFUAKCVrydrHnYcXvPiGpM02+vDBVEerq+6phwRh4SiD38q
+aHbfikgtRoA5xbGvCV/J6QLw2zBe2cjhijrV81yj6KUE/Jk0qNxc4en2KwynwphVObE9atM+htN
41FFtGWaqi5le9st88c1zY6F2S36/LZQ5EWddbuDWZqY/FADkV5NlYQsXcPfVjouZFePFQ887j6C
+f3ePMHq15J1JeGjiCPqUqDzKerfp242KOn/tuDSfzT4/wRSE47zLV/ciLDpS/g3GJ4U8LXTPBpo
Ua3usRbpsnzYp2jG7/dU90G/6Q4V8cAHcFPpyuu0fFpLxKK2ZVJluFiNwwIWlT9Szj7oAVTG3ps5
bX+KctQBm5FqPNJ/us705gh5DBzX1Q5QaAkH1wyqq3LeX/4/hxZUSPOeGj9zpuE6IWErYWM4xsPC
dW36is5yHTLgVgnsH73HwexkjCpwrkfmSQf3PPaQQIK9+uqGZ2cf+EKBohxTtRnaccJOMCs3wWlg
AhJ7oci/9QnN9QdZIK/EQSAUn/t637iH+TxufFhXAlFdRG5RABbgWGgoFLThF45fWkqVfPicG2e+
EIf0NoM7lBo6DNCKlxtbX+CumKJjSnVJPa4h6QF3ZYDpKb0uG4ufW0GpgCaMTlXFVgWcHetJ3KD1
l+XuKorIs3AthW09H4dEBmbu9fMI0dzS84+lCmYnzvsJO9w19/afF69GJbNngpLpdWo01JWUOBZB
TLvWC9GIJsVOIBcEcpc7aqa3puG3spKD5v6DIc2YJ4jEOFp3ChlE2RzQITFaPe9w41tkMELq0wcg
p7/HCijO4HnoFHJmA2uin4nl8vW7xuOSBymnMpMDxtMXZnqqVOtH0u8MqHUXYGYgRBSpYFJFknE0
wtVH9fkJA/WnrvhLiXc1T56cmKLp0TIUMH1bvOiATs9duY8PsA/zqkyMXlJ7DdYFqYRbjFZ/hreX
XRFOTwzCU1Pw712mD57fBWl8pWBiMsUKmjmN17QcJ1zZX4fKs0TEmvWQAcqfDBr6w/+yF8zFLyBc
jNJ2S1bfMXZZOAU9UCIVtLSGxTOaR86KUkOeDtViLRwbNBD10jAExA5IHC7kro1+7AHKscoTQYIj
idJJwGInZ02zfS27Cx1TiF/O79Pkh8RpFH0IhXJ2QE29QoT4xotz/KE4seAbT4uuGwepcIEuIL6E
/AK8SvcHiE7GYVPZxk+zZMtC4QAx3ci9VZOvWVLCSq1Pxc8cmZo5E3THgqrL07+ugcjAWNDj/IHF
ESfjUZJpkERpcgFb+5bQ0xn86MSUAMlA9cIgE8MynIsIg8aTEGtwe2rgL7/K/zgDYGRQ7oEkN1UI
eVqLAy4xCp8fEzlqghdjfdRFmtSZ5d1H1AhD52omZDpLac3dWD3WKbK6izSRv6DeV1nZGY0Nh1+w
nr5jfdk88qEPHG0zyvUjEI02GDKEMsEnUq3zP7cSTt1qKbsEdfhgkBLM4QtU0mqRRDOX3JFMhnGq
GYigeCxNdt9D+QKZikVIrjJj1lDzUHUaf1j3pkoHIxlKDxXYPsXi/kVFEHcNruc0BOeYNi6QfiIP
sUtXvEUpJwdhgGVZiHaAdRUWM65jK/ly6zcRhYGnGbE6wGCmQwK+MGwBnU+zqPce3z/xkDO4b83W
LRuxRCsVGwSnnDp7cK0IJ6JJ/12/yPbH58MNicws+TOSgq5qKYGoLxbLA6MagLPDL4IXHzspnJxg
JQj0Rocul+HP2CmMg0Rr3dgTxdySJPbP1/S4kSiIf5+kKd9pBtl5ZZWXZ+vgZtN4XAx8V7um3gNQ
Rnv0sLqhilnF3kzjk56KGv4+cBgjeKoPB95RBVcP2NGu8NZdob3pbzLMLD5M9mqTPvBMvlOmMDXn
jeIZtG59f2AfTLwOwqvDirQAvjQH2/VTYIR6gwCAsBMjkzBKZyfFY1ls7Z0j99wiH215zo8tAiao
nP3TfJ8VOVpwq3jgNWNFnfrFZWZE177/bbrarUKy/l6ZpwDJKTBMY5QJ+tbX3ceLfdKSl2Z9xm12
7PXfsFsJV5AZRPhydkQHqFImlJKwQZC8ORtGJVFboMflnZRsOvwlQSZIzjKxAi1NwqCm2pQmJ85q
PVXT5ec3JmDTloRnao7Fnt3/upXNaYo5XsLa5gA/P8SqyvMFUYs2gzJ99YA7SCZRBrQY0jxjaRqA
4BOE5j5sk4aMmmqRs7ptGJIKpexEjuEI+AECCM7If7nDcNjILuTjWeomNVOgfgoIvL7ujlXCVva4
zD525tK75/84Y8onELQT9PlDi7y16M4vxQN4xP39lzzQTr9iAkw3/jJFhecr0dYrOU1Y0TRwVNLO
Th8bNziojudXraRuc7DZkcwBn5bDtKbDHloHNXo+1HeLrakMtAywviwktDILWV/Kd3LGJz4GPsxT
CHMLJiAIrdrP1aS6UOWIj3Wf8AWCTol3WVOhNNmPsM6bk6bU2ihCusxNlbatb+Fx/VDjepfprFuv
j/zH/SLEYeC+huqhlui0JQNhOuapAe8vWAvE79bFKcO14MTJhvyIb5d7COyVIj7DZrHOJCgiUlEb
Bzp39hhpY3hBBBWxB0LIpd+nysDraGOetkVbNqTSriBgqJcs52Mvgj47NULa3PfuZM2CX4JCs5/B
thEBzvxPUrIUt/A33Y/7WcW3SZJec+aBLIH/Ku/BUtfuRqO/vPNnZYtBhQnjltsDVeYDdtvpO2Eg
XeLrW0+hhuYd/SwmVq4jiOKaMIZ+8cjvGNQglfCn2NxfY/tJCa6uYd6pP7o566a12FhZOVdBiP2a
j6IZpFt6ZM7Y/FacM4E1mMzgaYYv53p3XCBTRKBNIzEwaahLKza0LUAXkHQysDt1x/gGy1pX04mQ
u7on60raq2bJtSKQLqYQsz2s7EhnXLKx/Pa4iDDwyngjCpNAgnEsdXTRl50P+oC56kouuSC2g7Py
BR+PpW4U//w58AQTdTy8YXKVTET2IUMME5gSXZ0EOyWXiw9XtMr74vDfPe0Oi09z/m/VOi/rwkY8
g6I3G/dspg4xq1sMw+Y+JPn1QCVzwWjYpMKQsyq1it/4659DeWqRc7SL3neSIZZkXmAsxtaeTG+g
Rh3Cs5zo7o8N4ERIt/QVitlt0OzSL2bW3YbxN46ZvCGuecIzUZE+ToOY31hJOfq3mBh28g9fh0EH
P9itWMLKg18sU9OVP0GMxer4wLSjUkZr9s07QJgHrpqdLTUfnAgl7XPlcmYkWMsz/Ky55DDMpBI7
XRW6RLdtmBGO/tRSulexP94TAtzXrAuWU+z1cprJbwX3xyqA/JoKjCJmaTDbDspfVSoDb8GAZVzJ
lLHWHKHxcPO+tCjdnDsiorpe3680uxyqkTIx1dwWodpepDcjjIGEx1kWm0pg9OveWfCqGB5CNwyU
Pd8bSqSDvkOVeTp8HGfKYL8L/O6taue5bh4AvRCQUiXf5UwA2CnOBHS5ugbPEc+O2r73q1UcUcaj
N4OK3YUbf6YWn+W+ZLaz4mbnQxTuy61YWaz1QTR+sbgTID1F51RfFyRBpgkCa2QChZ64EmIZBQK9
IgMf9z2MIcA+pZ56xzLnlnxVTlP8CcKbMtL/pah4YacSVWUBqFFx0QvUJBZ3C/1IZ2k6iYzAmwnE
3VJuk4GcCjmd38UjY10To9f9jbp0AgjfivgXmicruT7zmcynBlwJRorSvGSWITXLszPXzCVhHx1U
oNsdzRUU7b5WEnUe/HIOKWwdODPwgflL4l8nYeEzzKx3kFVoDaCI+yZBw2u7sqawQUNsC/gtlv15
+QqO7D3gMpxKAK6ie2c5TmxAw5ySY/ZLzhPWpknHljspsHf0onz1Dg033RkT/nwKAtSfLkb25pqn
+0OVykfEQJxk4RsKeCCHxbPooIvQPshtqBj33fBSlffegYNfT2JJ986zF3pBWTpTbkY+XhVkOWNQ
laUhuIyWoOux6ZkERvGw4RjA1hv+5KKOTLCuqgYzTosPkrmzTbX8BSuSAwNi+Huz9RhzejdYPsVd
SPtZ93bciLFtb5mzz97XiREfWZRks3YO8dMbKKYd2FTi13rioFhBm5+ASnwFNNNpb1WwB98QigVA
PjZirM53QZOzAVKaQ196Iq+5fE78CptbMtk3hLj6npMwKhhkDSMEtcgUEWLFqQddoc8eStUH3FyF
bn/W+/uRaKrnZlCKnOKvV/88K7GeUsG/3hRs5Wu6ifYPGJDF/u8HKIjEnoOXUxj+kEEIjS+3yd34
STmrB7/G6hNP5l8o+Zejk6ij7rs32a3+UDJRKHxMmddGvJ8rb24IAms8zsqL/9lm0x3BxTtqpBc/
O54t/RAc/ZvlDnL7Rj/UoYXMJCWZXMegBmgU1ilfPrLyT1nUHLqMqAuEIx0NKxVID6KL1W67P5Cp
mySZvawowLH37P4cphUIZ+lXfQtZpU8xk0vuK4OJtFPL7VIXwCuEIwdgbdTCatrnhentQTNaqJ00
w6zZFPolflX21FogqSCShZkDvjic9MWQBXWXGgokpgEt+qEC1sv2eOC7WiSQMhOHuaxJzqf32dAi
YGfgxxngLr8044+RIYZthYGkogu5DvqQ9SmaRwwv6lQgkPPvMJCmVolJajNXKTtSLJVf5GNGsLTT
UlBAI69P75FNpK/8LnR8e+16meWuoWUpjOIR2sOXPXN2fGa7HjsypxY6qffX8QSl68U/V3VhIerq
NfEDjQsE6kTT6VF6DV5+33M+0gWulipOOo/o+UlLFpmd+4G5dA3rhWTcKql/D96UQAMEI21WDtjf
sMduwTmZ1xejuJnYG0A/pDf1avoE9k3nxSiXle6yrDiwbevSrOFzFqFD3v5AfUnFknD7EWp1s1OS
TVrpt+3M2wqTEw+7hwcAhKbNbPrrfUIVA4VLQWlkry9+FX8f5qLi8aKRLom77Iv1vbJo2O1G6OCs
cs/fA4zxfeXpLBF4mDxGYKrw7ebBL/JzDLgWXfxCq+06PsCOcQ6URoWKV9KfvcwttpLNF9bicxTK
jKDnZTCZTvRlrUMU4g0/klKN7e9IBjuIpro18KOlWupyxC/tZSzL/FA/edRIdNMY32+JKjkGuJRe
1KWaXXJylldmLYwsBKyly8o1XWu3GLZuQbndgYkj64I/Rmq+njthP8D9CwsAktwprlPcUhdbIdBC
wA+wkX0xuZYyPxrTcpoOHxe2GfN0FtTt3lSvQp641MSD6F6T0S8pRP0yhNlc/Yp7uDrkGXEF8d1f
TRHoAwAQr8vnNNlky7A6L1wgIcyn2FoTQ2lW9tIqfkc9w2CFqtPC8YWZFnoH9dLU5g0UNuah+Cd/
Y/RZoz3EdDamwTF3JQH2SQb5LHr1V0xqZyBJKtBlOlDyn/f7+hABLMd4r7J3tCzFPGSTZnSkK7hd
cZXDOf3Mh2WTyGnbG5koGnp7da+Y6h0TMME+RJjsu0PaDDQe+zLRFC2rNhHPBPtbyKsLQAA6EjwG
/7GXLu0vgh0TG1Zm1oQlIiAAKQ7ETVtyRE9xh8DMuxBrI7iIL4c1LP//hBE/kdSr3YSDtBGAH9QH
mKwsNBdLxdVgk+1ZaZAckJPLQ3EPm2flNHEpadOW2lHOfpH1APNJwdm0LRVlLGL/QRjH+3OkwM55
XEZQ4DwDeWAfSxIdyfP5p43vYDPcJlydX6WAaONn3HFcnwalVFem2r+pZq74dpSjmfdOCNMYVyH7
sxbPlez6Bq3Pih+Ppd3RDaEOEzPOcLeDhWb8pjs9zKD0S6+E4B3wTsSDBD0X4OaGIz1rnovowoDi
Mux6u/kzMwdtr88W43yIdSTmCLHIcIWQm7Ij68V2Cqnpe6uZnUWWaAfFIWpdpQ6tdSs9G6w/mpSm
7XiYSB2u7g2ZEAeWP5auKqHgs+D038x+D2n3/maq5gm6N9+kQdycw6GWiH/FiA3neelAf1S+UASz
WgV6X86BjjMF4eeOs1eVZojqAzMkOGTNIC5FhvTpmYt09mNeniEDSjz3rYjDlq1nAWMiObY5gLX6
5MGV7n16SJuHvbuLwsdnyuRTI+6iyWLNEG9DElQozFC0kvcYt+8lVURZ2DYepDLuycjHYd3InKWq
NUzSBhkAdlxb9VEDifzW7CzjkMSwKkP3BJy6uwgEIGfSPwC2peHrkWkCQG65ddHwVz1Lg2YrsqUe
Zoew3dw2bjOxluCdiyHMtdKLOO0r0gUs0HK1DROWY1bExGz/4JBVAl5tFwxPnhZtlTIFMZ2LxKmW
Idv2EnM857mcW+o+PuBEI5uhP9ARaVzRfyqFX5Z06ct8rissNDC6zspENFqPK4tMLq9SNAVjn1Jt
FBJXnBrqixEkgl1gS2D9PoEyKs4QuxMkDhOjNn4fUyLovw2pJ+CoXezvxDrFHQ0IfCUr6NYM6BsB
GyqC5cK0Ks7rzTgTmgw163FI0hJDW7PSODIW/Ecejp7asz0OsrH46uZt/j3Up63G9i/dmoqAXZeQ
BptZpapLTux5NC31vxgxSrIPdEVcE8CIPM1V1WzuNPPAGkDrGse7wEnpUI0dxVpMni+yCapgi0v4
BEFIIrDjrz3ZGHLucczsWYCIWfdG8jXKKmCw3gS+OrZTgxZP3VXDq2Sk5xgXBL0aXJJ5+Mu+y/Rx
RJsF9lbYpydG5RqsnJsT6f6fnbbwIjBJV3wZSkwjanswhLonGrMjUpfj49JjnOKCIlCTie01Gl/r
FafMRKbdv4EFu2Rpt/2WrNp+k26yrHbvrfi401n5mKysfSHcutK5rxcjSIz38Ke86qL/8UEIJ+dh
qRiy3PS8DAcWhryCP+N/q47i+o2aVs7yW0AZdDa62qqHaiYmwwVO3HFdE9FESq0a6bTyA3Zo9f4m
w9q4T+JsbeZ75wGglxuv5BSbf/fFBdwpYXV/zhRpLa2RuLdMUO1niTqstKfBIriX43tOy31ms7l0
Cn3lQPQYDXkne4L1FW0hKD6DAv1ksvAK/OJs2psmDWWmM5913gFXK0qyLlT/lF/SRp/5Otm5+JIx
aWxTWJ9frrxPuOi0E1x/tg5HxtKlxGxBJsBwVdat3sjD2LVEylPO10NgDWMLc7D5t9Fjme24Z0Vy
UE2tnxw5fL8aZ12NBmJZz20jtTKglt946fI3Qz9QGybt5d+V35BBncT3PmUJ/AJePG2+LFCSvqBn
O4sAhtencwsOwtieUMkahHnXhOX3LB0k6rguVFyXKtpOnYa7HTpj494snAR0S0ZVxZZtzaha5DIu
TAx9QbtSogGuo/RXd6HdVru2Y90dNVNDcp9Vlp18n3ZsXfiasyw+TdY9cBfHuNogdoxr/24aqVjp
oeXDYR92JNEWmHLGiaPlxE4FpecqEGOiAQfWGbN4BmUXkjHKGV5bYR9RJBI1SS4UEr4H1XioYiKj
d7QDCS98v25zzFpIhngIg7AWOdCFSZbV804md+L8yisqtT/k1wu08fz7htpyJuI0mIIXQFov3Qxn
naQdzXOcABWLtWiUnKYNWBBqAWDkO16F3QHkyeY9Fi7Lpd8GtlM5yi6fJowg4ZN363dFgwX1SidU
WfHfEUUrk6VBE/fwWKv5UAMDMO/2Za+P5PITKBIbsEwrsPmhxht8ulIzoXDzvWHY2rvueqjRwRzP
bFj9IgrX0sNLqUJAXgcZveXOmlj72lojziPKZIhgl+QWEkcJacUmdLJUcp3eW7VqTqnVmETqS0jI
qU/NE2+LkIVCDgi9G4w14QeXo6rKa9DxnRmHiAs0FD0YeHiBKWzCj++fL3rN3w6p2A6mENv+fUCD
3KDY3o2oaWlzpPYfEeyLzvFO4nCJBG9qTkRrRq8W/L77vl9hRhv4TeqlC/TMEhGbcem4r2F+qEuo
F2sdINLJctfbkl2Kypp04FnIUUAvutDTLasQKbZ3ukVKLluIDJ/QgQtjgOa53tLQxP5bYSdyEbZP
w/etVbwHaId+uvNMuCDm+zAxCHKq5f3vFjQ73GVQ/uHu8fiZkJekPyRE3VOkCd0uQg6blJhSh059
F9rzkAKByJgQLlFowXEV7kqK+Dxf77yNA+dIp5koPAADAc3syq5xr6sazrQr2Vbs3gKmNzRD/Gpw
opLSmMy/w4gzldFUEq6kdNdDrBAo+Q38ZWJoqdVselcZvB5M8ti5z51aruVzqdsquTBAJwHO+3lV
yCibzEP+QadjudsAL8yneBCkeTAZZz5Gv+U6EDFZqUmpXNOdodSK9faF6no7Ilx7xEHqEQUdjPKc
abjT6Pua8TdJd2M3G2i0A0Eb1LFXcEjlHMHBfG49m+/v4/cTTfOe1D8yt5L/Zp4fI1/SGyPhk78f
RiGH21xtQ6mVPJS90SfXN1+pvr+ow3D/pawgPnzBklyxzn+CESzCsEtIbXWpZpBEl92k5tkPmqzU
Tgt+rdJRz6c6DcciR4QnHsMgpCgl5EEyx9a/Vb6mdfiZPsa+w5x/Tv2u//n8sKAuDeW9UomlDVr5
ZAVC6Hn6H8/TpiO/46CX/YTv07O13+L/IPukbzgtXhPqXtsUg1Rmm7VKfs0Af2hNWZmDFWICIKZG
hF/4piKnhoLjR28Ok1+DSb8tgrF7VpgJgSPeHAFilRs7kcq2gU7oqxRRlj9Ta0Hzlcs7SAkdILwT
PP2D/JZKJaAHaRuw548pXngM8G3X1KYyV2qzaw1CCZQyr0cNSjKNM2u8WAUfjZ4jMcv3esnOJoKL
cIMPhQ8We9hQdmJ68WBLfWCriQDgpKAqkIV9I/wE5HsIlznTWuve0Qjp898dW2SPRGhpIa54y8t0
ec4nb6XK4Xz808vk0xnG4aSb57WCJJXnYmX4DMMusu49XDOzxYJKUEiq0tJIYG5BgNL7ypeG0ZIC
M+cMgV8M1NUJG7zga7HKGqGCWxzCSUK7w4x9vdWejSIAmyM80F5MqvnGqir64ILsrjJbNwKnywzh
QH8WKsPEzo5YUbpWUwD/jTdWvG9GqI4IarfiRcniyO2hp8XNtjKTaYaUu6huwM26FmmrU9zNk+Cy
P7YcccFiPL2TD1dgXCggwAj9R0vfa18FFuq4Yo2GvYvq7t1vri29A0h4+BRxxNRd1mOFxjm4JtDv
csHnN2Ll455ttpi1tJ1+pC+xByhhALUPWRSYJw9Wh5OXkZR2CeeYtCycmo+cXafTktZB8huuXjtO
P0LMqjkU3ysrDDCvoyl5DC3jN8zfCoZlnmxsXyhv4q3q8mgipXhSwZGvM/Gspy/QdTvcw2J83nMK
jyxXLlvCLSEXWCHKquIPTlZpPNzs8tsOtZbj3JdlCrsqiU8VsRYr0E3yeOIaCQVs0KI3WUU1dvw1
eja2tfMrw4VL9HRPwkYdNj2KTlNX1HgkZj7R6VmLPqf56sRsqre8DA61zDU/xMbh9qfQyD4P2ZNw
bG9rsJux8HRnoLSRr7lStoGnchEX2FG1nGqjHoshtJfuvWOvRrYUJi+KyFcwNu9lG2rrSkEvJ/AZ
nI6Ra1VMgcw9vP2EY3qqlZpRU28dIlX3Bj+42JFRvFSJjb8jG6myNb9XHCXpVdur0seXipFWwCd5
ZVyzc0xMlOnWVciM+2GvMyZ6HI1INTbWAle7vz2XB8fvFm252DRedpN5tykw5dGkEyXHvGcmysnE
yWZjL1cid00VPG89n8UxVvrKx52XcX3W9DREmh7Had76Al3/dY7J2vlGLeR27LE/g9qZ/fdCsHXU
C4bEHSeIztJDTSUf9TPOjraVtBBB3zgP9cirAB8om1+1Z9TO2cgdJfQPAJTEzCBvwCJRH45Tkti6
JOsBhlhxObhviWsQcTyd+j317+3gIAu65X0AIIt2SR/GOah69gV1qPY3+xxZ+WDM3PBNLWTOUSZO
Q+lWcgzrz3xMno+7uhVwunSDUPfK6bc7xv28LEu8/PvzEAdAuc9rs2xai32Qc0AVE44DHAzmhPAV
/O5atUD5QyXqtOXA//hjuXsXvei/pTzZNN1J1HjJbn81kTfTS8FpgV4l/xFMYkhKLmmBRX8rWFz3
1oYzJeoSfyT72EeY6kf6BCckhxzl5klMnh/LM/d14z2F+Ua5LyYtsSzFIPcvYBh78A5QanflPYeo
njVqt22cO0GsXCghlv4SGRnzW7b1lIi4QGvtA2EJG2MsmfyJdjWEdtYjPk+K9Rgm0qcYmz1Nc+ok
s4ZuA2750ErP2+A5nZifLVwiQncrSFrGvBA9+Zt/SzT9pvf7uTImXdJNWugjtY3aOo52/waBPF3q
/OK0e8R+CPUYUj8vLQuU8/2NBzj5YjDFfOXVMb+pEMCszmFeqscK5hEITwKzpirhjQOvcsdHbupP
VTjSt7hLAXwADbnDYA4m5mvkdRhTJqVqgR7JdImqbnsNku9+QCGcRuEbhIbZCV727g87BPjLFD8D
4V63hFJfZFGzIsbkg5WL/p6XxM5ZJ1XYEPZ76N4TznWGGmdsGE0Ns2ClGGTS/2RHh0SWQXFwkHdm
+nuYLnDsKJ1liLb0wrBLUTE3SGEyBVyIDvT1sICubCrOTDP8W0XMBbYI0/Bcpt8F7pbeqWQINono
d+B58vjDIzZlQC7tlOtaNN42fYxymQS1Zs0N/p8c0sMAbsENPnncY+IYfR0wCWdBnuPfypJVfOBb
3vVsCHVxujF7tEgOmxrxXoymo14WKZd0uPMvoe89vawZ7jf6NrFNDte+B68Bz+xzXHANDIaIimn4
Bg+UWZyO9tLUjJlvPyABiDqJRjQEG7eyeGnibSXnJBCekLov4FjKiQQj68d8jEsj/4GMGkSc7OXE
ZDX5Rw23V2fy5kADq4cHO3IalwERFG9bK3Fktkpszlha7yXmUxRIccUIjVJqWpGDlSBjHbWqTTs/
D/mDwwt/vU+HBpCbiiQrLe5EucDgqqmZ189Q/9QOhV2YihyfsJoPbWc+WcFxOr1zL10br18rP2gH
It9jbD80SLShQGgDpUqbS+QOqDN6lU7vN+oYE0ANnYzwNpkv+ZqLUqDFx+l5MkZEOk1f+1bab6rY
qvG3aGXcMrQKBu1pzfOm7AUuPRUEToWuHQ6kbV4u6Y3FccVSFfh+oxaq3IlsrZ4/oe7lenbEWxPb
wdP+/JwcYYNFaoypl/jqPlowkiitVrUY7jwl4UHwgWSjMM3PAghp8rRH+fJVZrkRN1W/QcGutDLc
Rsi+QnPZ/HlpV9dlOfOaxcYk9YVHAACF6oLd34thjapTN9E1YSGls+vefM4fNtBhxw7fEKiIcP3P
34y4tf4/7rcQfbQtu6FpeOeS3ElxYnE7Oejr0xzCRtdfzTYOpIWul5Kb3Z1KfrlJcozYWgAGOZ72
mgJxEhjx0P7gSTuFyIdiYo6PZEvYpSYBkH1TnfnvXJWUM+Bv7s8ljZMrzlcekMKNw+g8V8GC90uH
3nTwE6FsmgOc3gjPGniw+bHG8uklwoOwy1c29YJxQ3FgsJH/2CAD4JCK5QUC4QqbPZV9JvWkxb3Y
G78WTTszbmIysyxf4thWftMZ06tIHqD0wDsdSf9MoD4KndhqdAUBpsF1J2p0NYWAMsGE+GO9ykLm
vSUsmrz3fS44j1n1O1drRHnwoaeF5OwQcuCdIy50XQxEev3HZU1NfAiS7nnW1De21WJc81o/BQnf
U4/tlotp9CBJKLX2F7k1qmcMfhu94qD0n/E34vtQF7EINLLJrjderTHXmRRO4XeKS27SBvnWh76K
zEsySxa2riOkmshbextvThiGzCEgjx74Gp6n6YvJcjN0QYdIUAeIkQC0ucC0EyeMcvAs/vCXe7h/
rzCnqZtHeM3KaH8fLkZ2HP3sRggmzm74Uo/v013A+kWuuwyI8asq7AmlOZPFDD8f18WEkLqT3aH5
FMMpMLTZ0ZPmgIlFZXRPW4T3s2gYmrr3rwWnV8T8rWv+XVQvrvBAJDJCDUMy1zWz9Dmcqq2RNnPJ
7eWZPXGiYnbU1PlfbA6YBYCpoK00AHnl5xh2320k1NlyQ1K80ZrvMZJsg0lititzQMRz/ot8wEos
UViX87k8GStBx3mcyLfgIqlGjkqEgbDe/p06oUQuKY1JqF1/SdoOd2b+EhcJSj0nH4fSS+SvZ82k
+E+hv3F60JGDxj8vgHHnBmcaGhKzvRqUxuPmrUdrlmpFbcnmz6QWF6yAHGWS/aFzNOpdJoXppJ7N
HQBkYtA3/ZoE46WgpMEHRjbNcu2EmcKRlmyveMlSLymu0qdELUG9z+DAn2V0UF4BPTHg6z3FA3pI
AtP/7lDCYDomyzTHp3FgRS9iuP5CdOgwyFU/RXaR9/x8/l8ILvYiVrCD5qfakVBD0Y3D7UTr+jm4
EPdtX1hoV+XO+/3hTEdm+tW1cbEn0R8gbDneJ+9q+a74vZpkikjpA5bykTXwuEjBozFRoJwfT0HL
M79U1H4uRQi3JlXb2HK4CFqfSIM+/6kOOkbiPHc8e+bXZGKlbGIvldFv8+zUcUnj5qN9qSk70p2+
brbLt2ArgXiOxcs0eoymuwfhYxLbzsZUFDLUdIJZh86LWnqH0CwfZxQsDj6JSF9e1hfM3nyrRX8S
2w/qFvWuSYm7PasTPDUi3Q/ORnWEvlNUlCFghkjUT3WNbHO21+zyOjuoNE1dBLVq5tMdvktbIA9Q
PiL4mXNCdkxKXtTbf9maGsXcKmokZxw/aNB4ImOc50hUCFiRevGr+RWoXf3s+ZohOiyh8lFL+D6s
dw8MzvMtWTg5hW7gbkBulXjqwu65UHN6L/U4kpqjsFtm0Nm1/oFDmGhTDsWitIBc2xUfJ3v94Cbi
KpT0xa904cWBUJer3/bG/iYU/QLAQwkJVmjO3UvqKMQJbImbtc4wbqCnGzETBENyuooEcphpAnMu
JYHpcb/EeOIDgx49x14FMWYj07GKvTvEo2kEEN/sQ3iCe4z2FnKeAot0EjQCzy1Ye1X6eWRpm3fr
uzXpc35bJvABCUtgU6NjMU8JuGEr9y8gDTcHy59FNb7AGEVk0/Mam6F9ZSkPFL5msRk3DPydtyD3
l4XjwcTHb4aMP3LFVN5dq5zGHxd7CCe1n6JesrXt2hFLLsNZU9oDeDvmF3t9wDmtgaP4i+IYSVEe
+Fajzw5llkFZKN/s1uvi8Ak62piz4qG2swfTTUyTusWZstw1pSStoJJ0UZkpZw2XVPntuJGYlhMI
PlIs5t7t4Rt9iFZkZGRZHoUB5Plnmct7Ept/QPKaNt7WPSO1RbOOLMMRvfcSXq5/6iM0OGv602hL
xQuNvi2eAH/zGRaFZQTJQbIEAkdFE7dRX7gPTWTff2ZCP3dg45R6HUF4ie/XMjwYfvenz5nBNoSp
BEffEd92n/uC64x2w2XZWn9rBT2BpQeddd9Gf64TOJiZtRqwf4bB4XjjCjuVdPtasmKcQk1yWV6o
fssnDhjNDSJl9Ql+FrZEUGYTKrQ45NReM4gL4FjUdoHH9VOjjpz3Aui2oqtDYGm/Ir2PvX+JoQOY
5SwWxZsOhpTED03Vp5JN5H8ZGt+6wyYKrLaT/4FterysyOv/RkdX4R3WEfvB670eSH36Ej3jCbIG
d9htEagyyIanJG0k9F+0w+xhXEtiefOv27X8yrZzq3dsqnRg8tnCpZuigukkVgbF1P5GdH/CQtZD
bLeLLFQdOwOF68e4oJJS7XslguIjVAU9nFczN+HF+SMLHPY2xBa5SkZp9+N9kDM+zdw5gJBQPPll
3uumWcTJWFtPDFB7pwg2P367oMV32d7YbgQurTFEkcTrUYqWicmq5SpIByeV1E2Z82a5oiZjl1jk
Ocgg9K6XrAlmydS4q/2yux0utsJNmT5zSHKZz/Uy/Dt/5QhsO7cdI13vOAPRllkteeFQHWpMd4Mk
DqTtWpc6B8fXYn/UZ12YVHWQIG75INwMr7y9cpbuUjTFx8iJZf/Ic8T09pqR2rQiem2wYq91LMlc
VUhWqMsa3yttbTYkfeg00SrNaS2pSSdWWKMJT0F2ZpqfONL5eYREaOAhWWu/As+WNgZZubWOPm+s
PyRTVFUakbYMwZjBbilXJLojflgEXx88yHAa2LoiU1KqiHCuDhMVUZZrHljIhbND4kCPZEm4GSjO
UbR0cMsxG5zJRRqe8ZhFnVuYV5tFhR2l2P8GrbIasH41edCHGNrbyk8KhTvbOGSMXIY7NUQ83/ZY
GbrxnDjgcF8JgSIBCW3fTEZD3tt05Y/y+AmDicg123DVSIBjGLMLf4mc7PhNNwRNx6zCTaT8FUT/
WwHFl0lQSDz8MrFEAeMJyM0kWzV/qKRUFpBisoocUGPbsggbYeSxISd4q0+P+ejMCcBSPKBooroV
gCGZH1qQC4f/u++aH6n7DsnxzmL2gC/DDMBCE+2CWIGYQJz6ojetjMqTs57Jrd9U2ATzAbf04K9D
9zYpDGPpYOVF8BccgX1YR5qc4/tUuGg0fR8yUbLgHBmLmWRnlm0Y/DZ/KDY9QCRqSltqPBJF337B
Xy+WL9/aR2pyXCi21wWU2eKqKPYJ+3WuN2TQ5+zc04FhRzZKBPZa9rLFqcPHCz2hMZ9+SDHIfW6z
OtSKb45fBTtROocBozacuSELMAUvLRL2b5D8HxKC99Z6FOW05Htaj9ZFQiYK97jg2s22XhH5r/1E
waxNTAqkIk3dVSIGQLvDFCO49iwB5wfv+7A4pS28e4SGWbr194UmOGJDahjs2MDxqLyrYZbF1xX8
nv+4QJbIx5Z1ZuGPL3PGQIE1dzwRKpzupvSJ9fyt5SxhfV3hfMWINFF0C5MkMySfSBuEXcJP6YS4
5euz471A4CwCb15XjzB6FV08T+0KUum4AreK3lr9heVimzqScCpIti2yjNgy1WBRnDbb1rLt8QGJ
FgVVbpnsKxL9WEyqY5w+bADrhMqbU45Y7y9gfRJoPmwGjWQ8QtTRJOBZtjBZ8+ZLx0Uc0q50ugIu
CKNSQSCjQB560hILazt1yTQn3kBk5GFkeKsoqOv9hyvSnljo5417yeqea7M23R3QwCsQzf6N+YD4
U+cWKnCW9JJehgTKxaXTnqk/w+tg+70Svg4uuWIPyK6xXjaTkYMWMlWxTiaduvGS73U3KJT/HEER
ZjJa/ZnjmKdKhvaVoHfvX70mXnZrdY12mlZegFxxITYusGq0qmSozF25ultReq925IV2ewc2drWr
TBS0WBgKJWs8GrlxCChW7Sggmh6cq2zrNGR3ZiJqNnSUUIn2z7VErjsiO3ULIRRSjU6D8VfQ2Cr0
n9mm+nvTQ2AAJ0MNRbvQ07iPdGIkKgT8oFm7pjIYrQeneS2sgqy9ZLT5sAttfnGIgXEVh/jr50Ig
HS+i93FvsA+XvU2b0aEPJZYvZRiw4uqGuzXnJZ8ATMEXd/7XPc0Zh0K3bw2ZErCV7yxPQmkdDYaL
EWClH29jaVfSz7RQ//Eilkx06zJ1MvI/JQ0b5DVhPF7zW5wIAYssde8xijmw6XvZUjFdLAIEcQ3D
orM9c6pEj2Acroywlt4SSKstCnjbLvJoaWXxp9XRjfe4tuJAwfzm7ziGQS3PKsOX2wGoPkkjc4Yp
gmBMhJhGSKu7NyNGiy6cDlDXS24Go0U05PZ7/qICp6yAEKPFs5kaBxEMkdubAPIyVdCG1F9U426S
k85mxk9JbnHwsKdyXbGQ/ttiFFqJevN5jg7aXWgs/b4I/hje0MK4zZ4dsT/dDEbkWUvL98SkB5KE
ADUGJShD0AWAfmJfKXC/OSXd1CCbMCGP5MCki9Z6C/8TnAe+OJ8KViQNE9oCKGnelBvTykrrS8nU
91i4C6MqPY8JAdxrSfFwbhZTg/TiR/2tYTV656kZTnw9kQImAzLD5kM9pjK+b8tqNKUbq0xIVblQ
/VtwNTA1sxR2ox5DC5nYM4vPjiJS4NpbT0AGTwJATyLLHLlri/YBA8Jevf0c1gU7mldMnWC0XWHi
94yz4dGhcx4dfaZyrj5JiJYQQltM30UiLLa+K5Vloae5vCUW4UQh/DRquen8jjq1gCPkMlYAOP5b
PAopG1lMeJYnFu+7sFkh+i6rqdISVyP3xKCeqaLb7awdngkP/eZv6GUfaZoVtA3JEQFLUmjp/Mfl
mVi1TD+ZD5zs2/IOJFCgQMTjuZRD4tOtaG4m/dKUrsmPLJ7BVRwgj+Y/6tfcInqdy1Fuqc3tpIYA
lO84Bek3gvfm4fZxob8vxcTaE4tTFQO2wZDk7Mluvcf31gHoOwxyisFym/stYsbhKdxY9dvIzB0v
y2AHd5CbHAMeSytdv/q3dmftszBXOMrGA2XUyOFiKPvl+nGA/7WmMoXhTgg35nd5WjQByaguzpym
DVcgCaHx75ueidQfgc96c5MhUuHAwfFLAw8yPf4UO8gS9/EArzXUw+6lBUEOpy/BoxN1H5ErP46E
JgN4muIQSO48pLFSycx1mFVS8TCHHkRxM/liESN88dwt20O0TNZZ6xRfomZAoP1EhXRex60/zeOj
lpTc/vKMFwJKDzJkZ5WFWTD5xbYHXOwRuYggCbXpUXHvlNSUlpNqljfthFdo9HmZCI+fAGclA2N0
Ii+qnoNgfZunWA2HL8/2wZmzaWzhugyV1BnvPPs7K+VNMJyV5aSLvUwHvfAixNCO/Z0nm/Pifv43
jj5NXGGsj+exjrrPoNeo7kUNsuaWYn5RONqhSxrEi2fQ9JsG67eyLf4whnK+UkW8KJ1dYDZhr+Jd
32bZj1sYNYvAFUQoFuloeev3tUZ/ABqihHLzrzFI5/w9AAkuW9AnW82XotPdyMdeVNUHiD12auqa
ba3mUCGP9EmAHKNyfHRZj8r0wQX3BlcOHYQEYbouF8tkxJEGOBNiDMVRW8YXErC6Xn0kixFC9AZJ
3FaIyDaWLAtjXIubcvKgp/hiT5A1DCQnKRAAemDdi2JSD8qKz56BsfxR/YOGJcy6jiH7Pb7tI+IN
IiwceDrRbShELU4JKAI77CCsSUxDTXVmct1CxwemPQNf0sv0/2NwWmHDf4ICqgAb8bFhZ4VMCWbm
wdUUV8Kzy52kLA2ofU2XTp9l8Ga/LSRCAptZzyOl6cWp9BYIyP/CtokgIhU+UecKHV74xZ7I++iJ
RVMj0ho1iS8B1Avesl+AxvP9+VWqbqSiQaVOmLlOqcVFoG6FqM2jTsxiqG0tncGapRrBvmiRz0KI
G54kCVe9XjC1mnk2v+z/ClvnB66XS9XxbQDq9JsFXUizEBOeqTbpX6iDy+3bTXcXozXe0uxU4qb4
bj6UucVZ/eLeiVJxgODdJ8G/rQlxG34wvjz4V16DzuKiCBGre1zj4Px8uZTJ05s9EJBIzDl/InHm
zCuQulEVQ8u8P+FzpOnVNFpCzb2rBZzxyYF07zj1FBIVQDOpDSE9NcrDAwCHtEQd809p9XZDq3y0
F5d9ioyu8MjkDjW2CLNzSjx+ljztS9kf3XCNucl4lOpbHY6sixlKogNIOUOtXx6YyPbWCK/tgD6W
2520BjrkW1FYmlxLBNF/rf6Kk2oCSSkOh/dMD0pVCJc8810/ZetcLhekHhaaJmvponpEc53UcCKL
/u/YLRi+2nCJsZ8L6oWvM2taAaNQLprmWisnxlCnUnNY0lbJt3//llTY2D8sG1HDPI/jNaFFQQt8
gdCzBvrLuJdLOONU1OCfCPeA4VKBQNBianMhZ4hTMMnCHlukHbkijRtD84GI2k9dEAkE3r0mQ5v2
TLADve56hTv2W41+QNw8kpHMbQ8v43BiiE8v0CzWnDVDM5DaiWZZSQPOeDR3zXZ6QulYIuD2tXL3
c8Z/oYZXZdUUI7RTd8wPRa5+2Qh+eBXROD2Ufqq23TPzPdC5J1qFzxv/MfysRq6q06CkktPiXV8a
f3k8zwxZj4Dt1nmCFWNGbSo3Yts1bp/58zhIRjy+Cjb2gt6FBVmhgYl4k+ov+2dgthiRzwTRuA12
/WFSLc/ErvCtHLHe7t2x2HTzJymYM3GdzsAIcvmjonC3uUQ/Wl4tJQi8W/pGvzAW5121Jc2Kbkz6
NG8G47RwXGomFu3ZJAuqs5uxGu+hgTeptqnHXtRgBMKzjXdx+gmqlWOwuLTU+Z291mHQuP7yAxeh
ojUHKUvnylyeicCazRcXxTBXIsP/tNYpaIA1lx4GYdJvD2EwG8WQKZnnUuP7h4lChWuwEGfALjF5
g9lQkuY5H7FLQAbfxetAU7c9nd8dNIBZ1z9gVdDVIvaSSaRU2XWUrZxDgbxg0Ug0aDawPkNjQW6H
FdIu08rs4bS/N9VRu18mlM+Ty9m7OLQMFQt0XYb+rgJZ24YS4egahiV71hqSG01+qFx+TIHhNXsp
0HfA70stuc1KnclcM2RKFdXHINnLwAaPLPSAHm+70qq58/OwFU0Kp18ZTYtPJ5d43GrIBmqAhSH8
VuyoPIWz7snl1NNQJrsCYQ5zSKiH1j8LD+O3I0LvmFyR1d4ZLItjd5bYjBGGYEhOauqkmVrP8Oxu
l/eSe281f34C1SdfEGwYG26VvvHiQfBWLxj7zFV212Xb++ujJYXVTiD7xZ62HWqqI018duXB6XFc
pkZdMI+E04zzjdwibJMHA621ZiV/kfEAPrArr60fzh3WqhA82OvouWz1EQ/MqVFbqGIAjBMy2vrN
g8F4KMpANNn+JaKN4C1H6DMRdL76zqdNkHfkqdxC5Q97mi/BT5NBEHy5ejYbq3m7ybVTR7imVx4s
v7CZcdEsaVhGEnXOZjIxqHboVuYFI91nqZzVbDsv05v2zZCCNMnN+NiBIThcNKet6MlRYhoyIIqA
72jjE5zZeMlk1a4mXex5ag4rnQ2lSYvKA1gUMfhPUmrdgTAw0fvxPIsWuvzhSZ1Py3D16Lo5iub/
VcGFR+F8ImiJ/T44yAX+P7T9lU91YoG66GHnTyeotIINyqI6hkN0CPqzTIhbBYABB9hTWkRnGg9p
ipbpk1agodPugvCwR6JqAYtUZ548g8bNXGl3D7uEwkVn3xojmpyvxIP1rxL4a4pFOEGIfnX3LS5b
eK2Wq0mOEaMm6zrROM5iHTdbSKYhUZqMxGbgR46orvdB5wICN4RiTdoD0SoJgkRM5bD7OTNTf3BY
9h6Dq6B+w3+21+cZKDU7KVQZOG8LchJrLzPmFIqCVDGSdi5EwKWBC4Oz9uDeUHFdqx3pLGvCAjOe
rQFXTK3NwljpZ11yaZAI3F0oegU0JW/lwv4Q0+nUY6ON0txRpjQzJsivLWMOavPdFFfDd8wx+mRs
CzqMQzj3ct+HW5kNguMEUILo+UVRpDn+RcJ9CXip7d66DE3eTVvMmIbnwuODFBVHulhkXEho+JTK
a6s85TtaJ2I0UQZmZoOuy6ti83Io4aM904DHzZL8p8MHzqiG3bg239b+9zkkb0Go/37uzDPtVocj
U9E5zhLFK2RnevWTm1Z5jB6XCuOZuIpdN5aZOaJw/TBTCNGXl/pE01QI1hM4Zt1FzRCUMhP6MSNR
naUlDkBxutuv62xJbd2sMsUyHmLpuXq6HZozL2fo7YuXOQiiZ59I+9FYA4+yqjC7rKdKTW2HIO0A
JajPnmzh79Row2ZGQJ/uVhnvY+7q7a49biHR2Noe/gGSorQmL5Bn5rnj2ZbXjBgjN8IvFYMTNeH8
fiJkOnj9l7b5to4KLuKzooUIp6RxfTra3UyAtQE7SFlIXMlqaFdpzGeG1uAqy69QfZ2f77/bUWdI
GvtueqJ0x4xon21mgSLNHMglUzCwBxr/xsCcwnPFHwVobxlAKjE07Y9WFizmwVUC5QaAQK6Y3GUT
hCgYykr9iNptIMpWufwt1Q5ELmw0ONUPU2OcaXCkmFMFFKFolUiTQgo1Asg7IvwcsB1Q5W0wqt7r
EfEdbBTDvbvrp3oU8tL/Rh8jGTGOyFQ9VtWJUmU+g2xBM0f5ZkIH1QYtl5mJLGvHEaTRsRzI+kIG
Lot+ngPyXm6w6FcS6/SDeG8ogr7leZwDNmHRUT7K35tqDfiB6Gd6Lb1b5JIx1pBf0JCgr9n00HTy
l162kQXRN/KEEW8ckkG+W55o5ojVXDm9f2XcYjp7yHoeEQT8R70AIkGqwgsEw6AGLASRrLLSdPuu
TyArJD5ySeV5OXdbxXXiwzZxNaOHq/y9kUWuDIzVzIVp7jgGJbopkKcZM9KezKXdhEe9Qvbau5Ax
zqWS2S17sfd2cLb5KWnpcFrNLB+43FKxkT3amxkNALA+icZla5xZ8QsUlU23Xy/J3l6bSMa0TWkz
KHOoSKAWy+UVTrVM8nFHUNuDI56DtYUo+kQkw7H71u5bo8iXLnSAgMfjVaE87s7rgrLeRIoROHQa
9CQ+9Im6J5VZALgfLphQuQZJDFqU38xJgcDBSGBs1qO5dOCSg0Tk7fQMJ6Q2cLICYXTWaPhYsyrW
laBO/8Wti/YEljNNbHtyJwR8qfwcTJZW7CWuYFs22UZwGl7AuNQ816hjzNNUto+S+JC6ZnsXMnep
n0QLrnlIAm09s60mpPVFUkYECPK3KEN5aV4Yus6J/AD13XHe1fiGX2CT4WMwYi3M0jVr+MD0Byp6
wV26Oqbp4KVWBLA53nKNLwsEFnkjTcJOtTLWXZaEsDqwYf19M9asJw1FKpSDfJ80MB9HvT6H/F27
Nn5bBJhR6O+DFeFl5qmChMeiwT7fLSzw3LNixx5gwQI2/DuH7sxQ9O0aWxRyx+4mU2LxWNZDRZL6
+Wx7G+89zbWfKKQMcd9ESN+9bk8ZtH0Yx5jeNhOt0gpN+gkAJtzbxCApeyKbAOGvIbLyVqCwPIe+
8Wj7isfooCGR7qma5s1wZ2CSJBK6ABaBcLoV4OEZRW2YyvG4u51+w5h9blKE5+NdpBgysLnQRCfX
Q5cApeLqDBQjXvFLinQHhPGcNOgJoFqPmxNADixdal5NzD4dVsIjPYNkEY24E6mQ5kwRYvKyNv5F
1Q93UzwSdT0UHl3UIEmGQz0LpIFYVGYrGtF1hpP3A0Az2kePos1lDTL5Ib/aLB/1HZPwetYKyCHE
S2IJIDtGL61g/IKt5K1ve/5ulnM80PxT+zmE9NEKBeVuJQp7PwuzZU4IwtZq8OFiwCpsTDM7EH8f
xK2SciydPpBAKfCqJjXyR6QNjYXanRtPBThH3A2yU50HxEnYjOAnVhmw7J/TmhDTmCTbMfjjaFaR
WSgAkWvOVErnBGtnwuPoX9wnw6RoVYHR5VkWfzSdq++fhQiLXcgcAVmBj1mqco3s07o4QmCLRfJK
VjVXbEyDrPuiqjyYsjqteSZJPwzRstuof808bb62Kl4NdMJjcuvNBz/dwKLf1YRMCPFH5rPXTfC6
byj9LAWiNWS+lQKhmtIB8o2ePCeRTSUyVlDkdl5/7fekk6Aig/+NGnEE/minYMnasSf1VUFyF32P
Tb+Wo6lISpz6Egn4EV/1m6CyWn7Vhi6Tk3L91nNn0puFwHhLBD/FecPAVTfeKCl2QoYgfZx+YmU5
648Y0CacZsNo3vHXMRoUwFS8sMnRzILnA04/Gyu47aRzmrEX1O2Kt/T6hfqQpMo4yOPow08IgSRJ
3YK49EpYt0C0+iieZcHA8JstF7LqGL883sF/31C5yThEtoPp0LAkUTyIrbDtD99txazS9CAGyDN9
KVqdMMquL/iFdHgrz+JWwzWDgNijWzA6PoVqa/0wwtcgyKouCxJGGX7wl1cYUFZwrLcHwVJ6DGxw
xpnofJ+K5KGjFCWGz7MU/8MmyqbYXomJXLQXOFTo2tTqRsTUrsvTcyYihI0I5T8zr7ksMZxtNGUo
+A91bTnUHg9HTw8EJqz9hgqB4XQb6TdnhbHAG71tkXU0dBJtKvQar584mlLI6d1BosKb2zoTS7Mu
XdEQtE5pbYklMGqoQNIP59P2kClB2Tfdp9c2N+8Y4ANjKgjjhVqoJJO/Ble7RJFpIxRI4ItkBWZ4
FQ0q+mqPDZ4aRZlqvOpnJW1YxAgCzc2DZoC4BXvb8xo9WieMweLOaTnhP1AY1FQmB1wkJcPTRFMn
mhfc7jLL4HUiwseazg5xYM16dBR02P4NgdJRyDdgzb683ShtNMkjFSoQ3dADE08W20NeugWJyeqq
Xeb2pWAA9bhiYFmNVJbZA6rLir4JBYHQ+veoZzwR1RS7sbEAjjE6oy9UmYfIuqvzubhFS6hv1VDl
8epHsr3PMQE+x+zRaEB7px7u5/lY2+yzxZTuyjnnIKVwjegntgHVI5XiNcHtjKOcrnoLLJ9jvRSs
qzHJB+G6+xnoCXeD07cimWS/iZ56WKKq3dqdba9T6Md/6AH9M5c+q8DqOuP2yRqVQpnZ7nC9KIoh
WLxgwp7/+7RdWj3BWBvU3MEXhsxSamAuzvuDLmUVTktV+T1ECZpWDny+xuGHWQpYLYLpeF9b7kjI
Q6oB3q7FGuKWpEMduc01aIJc8HxpisSGsYDiGOf6QyyNeMvpGAD04/C3DNDpHftxLYGS2XBEwGj4
Nz0KIsjM6zhDdiwuAji9+Z4BNzCTnlgUlWEoaMGsZF8/h/p7xjT3iAIGRWeK0FOfNUy9aT1OAPdt
GWKPymvHK3fy52XhR7O/thH9IPx/SDeY+TrjLQUVlQv+DSnYH407cqHRZf4bzK76tT9GMBe0lYFh
0hYCjvb1ubPdHPgxCRdHVebYslziZVVWo+6D6qET6oEd22Fwj/5izharV158WUhLDY/AogRI4R37
1Br5NrMBcyspfDlGoIVPZYj7HuKhnifrb9IrjyTmQnfBvcBc8GBcN+r2i84hSklghgOR8M/TUqyN
sK3JZr/R2ATeBHvNTMShdAcdi7bk6XdP3XvStRDqQxisQMp84QhZb/Tp01LQY0wAkafnyOV8dVQK
uLxP1qd267uFALEqaqlhOAuJgUl1OZvP1O8WSxbyHAe08vD6uFV931RuYhx8iFX80xb6iLCmmmM+
EkUsRFBdhOxjGZCws/Q8xr6SiXwR/i0ChAS3CNXMMfBzAPPB/5O3XYrbJJS/oayblZaaSHZVesff
IwiGAopDn7F45wX6E1TaUxoc+JfWcR1CVsjzYtTIjPf/3PhOYYcPSNjPkdzQUpEWxn2KA9ddGpKU
sCOHmoHH4KYsikH0GoNM6jZHeiKDdHwuYgEL0y9AjsC+tQWCMTYz1Cl7Q8gNd5nCwvrWzQroMJNC
btOgtty48HKTsCEUp8MSL/6q1SXyCj7XL1XpEmT1DpUGPcLzAQAKT3cRapPNipCzcBdDARVSzwg6
aqYGbgwxKdWlF/+8AeR4gptjqqVTAscXTA6ciNJMymtJJuiAHKc6DuE3ci/GK8Bt+DpHIas6OyU7
+sHjDx/N9PNXJZyr+ynj17DE+gtiTtmEdSFrE20eeXnslvf81BO2muOHJUbKPayEA5xIwyJEacpi
PKhnziZ9DsDKYvbpF4/OfbLMJAqyIm4wiioymGoUBF5OCoUEGm+D0A0QCDYJF25jXjM1mJT30oBV
6SS+yVPiE0ikxGb3++8AaEFN/2Z46KdhwwVwRKFlLua0YyBIEOp8D1/ZvhVBvslg3AgHEAB7BH53
NMjouqUFQedC8PRTzfxX21uBXgJqwQf/wtFvlbmVd3F0OfRvI4BI7Cd4NUmkqn6j3ARoFpnyyBf8
ZgiEMfmr2GlBKWYmfsQ6+c+s/xO3Hvbt2kfRkrnvvHZ0E27+sqKHh0BijIrhOVPTHx82WkacrWp5
0vK35a9WHPYwz76Ms3RDlYwTbkMgzTq/q9aPeW8Emikz4x1angZ2unHIdkQzZpzIjf/2qFI7XFuB
TYruTCwfRSKT0aFcBrmJRcdvt5SWRrzQnNgcf5SiuIP+QAjm2u5ID39lhm5tbKYq2qlcjquvkgRu
51XgUgnO13Brtn8JVtNxm0G2muj8IMoQIgaydI9dNeESYzV/3KJKTxc0cU/mvl36ZBD7r6T97XyA
wrEdE4oXVUuBhX1gcxRVKdZO7NfsY462rH6UcSHbnGaWpf6/rlHByNz/ftWdmNpgDtlFS3dcGCmT
1MgPYJuMsCUVupCpvtBl5MnDIxRFq22L0H/qCrbn1dO52V3dzxr+8uIOxKAEi3TYZlKIRPD86TNB
pLE4rlq5OKVKBUn1v3kmIGgi8ye+Hplm8g/JRus+Mk5OhHdC8OBVud03qTnFn6gpqVgWDXpAD76+
1QJnyFDSXzx9Tqik4bzSokjKqpVpPVVQThK/4/lxUlkmfDQthNfiVlcCRAcDRIfxSavQQp+MC9SW
3DNoIM6buQ3aeJzVaxGerCifdLwgy3MUlvWNc6oOPmfHu5sSnwykkXjrsRSC1KXMDDtNjrNUtXPh
lvcE3cDhGHpBgY/zrxx95HV23lIHjPP15sG6RLjLopVvkEQ/bXPIYLEIp+IoVdmGPFpW4xex25Ep
Vrwwp+A3qHUSxnm9eO2XGUp5yUalVlEKd+pB3HTJ/RnMg11BvmjWOfCNdxBRGWy4OazBNeFY2EBH
SLGSxTFpb1HoJBIQtLlcFqxTDBpLTL+7Iuw8SQCAVX0wvTwzv8eZBe7os6h/Yyjj53n6bdxeeogy
r9bUSc1GofVY3HLUuCcSWIXHH0/c9VZRZu8ShkU1SO6xOk9rZ5nokFskj6YM0XSJNyVZR1kZxGWW
wA2nOEXYbuLMsWKTQlYaSFxqqwlR/nmigIuitQpvMDEddiUrkEaPh5qm4cwjMGZWwlQ6aSe3dWde
XLZv8PS4rxZ8K7t5ismVrzeI9bvDmXG8wAcMGREneHqcC9BQ50mkaWedJbrYjahNjoRm2AZKfI1q
uguOEumzyGUZM8PxatAopZlAZFo8Zd0oEbD5gSl5gIBYO3tRNey3rVvJf87X3g0j4wTb0G7Gyxx/
HqoW3Vk4CjjryuPSFm2gTzScekrfxVhv425JMgTkusBFj94Jzbfcx1P0fXUepHwGyFIY1thGwxgX
YayArIbMvneOjrLKWV4MKSxvOY7Il7EHjFwMucmf5llxTjh6M91jg+GRoDDj9HiZsJGxf8Bk5daf
I4RNuKq73/WGgd5Z7Zu7fFdHb+lr0B1X9QbYJXeF72kCQ6dVdJpEpvB94AsMwk2636J4HtCy8XEj
Ymau9M32/79dfvroStrisfJUkHgKE56yOpyPq8eJprvQZcDvcUirUWAWE4lVdyiurepNQFG65W2q
uqK0hMEiYs7MvNoUELbUUNMj9curEcVcOyJIehWCyUCP7wq5YThp4kP7FjtZr80I4Rs2cior0Rxj
kjm+PCYM9FHwR7LOxFWa3WSU35DzYY1ljs60QWE9IHAzjndZvS9R51Ih3MZ8Il7UIyCV33yq92br
09vnrKD3bPlOwM2kb+8C5M34DvPrMQ1VR0njiH1x2zMkxC0gi8i7F8xt/C6FLDuMjmS6Hf83c8C/
0s9o9U91v4Qod3Sv6Glcj1OSzmfWHN43NYuZmJ20tiwSxJw6Ml4KZ21HZH6WSpx/Rb05N9rlIoS9
YBin2XXku6sPJ5ILVs0donZPI5dqEsES20IAqabxRQnC7w6fCAfRCOeRj/eWLSYFipjbp0VE+Pox
KzsCoRittVRXEVKrYw+MP+YFAeWlgIdtpHwYKb67ePl6/FjCrgosYjVQhK262KtQcw4/pRfKUX18
hfyq3O+XQ+Qzdq4beqn9Rovd3041mDlXRXCgMEVy7CVECu28k9eMVYqQOx5r1SdUW0sNGDbaplm3
uJZr/hZeVSkdB85DSx9yzwuSijeCAuY6eSQRpqxq8tUI1H1hItwe7F0BwjpnOUR4HrcwDaP5sR0q
YX5XhQVR2Xcya/6l4TXVTg3RNanDOQrNPxNjXdJi2RPmOUuR4Vh88ukrNRwSBK+ahM52JNY5Y3kk
d+aSRmKd3G9NMTB9VEFEfke6SI/0h9LdAsONSSSZCqLtNZGASXT9LYCCphQ9/xYkL8gesaAIPyg2
7XDcMVc1r/aoRkcQN0OqAuy3eHug0Vu3kIfX0bfetyQ+O3W3y2Nh8KzVWNVwnaY8sbAgF5jL4som
/N+riiNX+7YzirMCH5cKTj6QLMsWAsuivAFETZrNw8F51kNyvwX+P3rfmEwctaAx3vwyx2zWPZs2
XhQDn23XRTw8OLg8XqcsmF2DtzZJGmr8vOXfC3hPGFcyt4hbwXsGSLVlHtl15pcFREIdNqeIE2y8
hzd1wZxjlPf8fQdvq6YbE7U5H/9LcmaPDZV58NmR1+UncYZDoi975lstYwYM9joNITviZ5LzOFBN
q2BKLzR2HTQnRANiR8RWXd4a/i0s+gVU3SJN39ksXISYvdBNCMgbug7RYlua91cRcmFTqhlE7IKd
0HLIfZCjiDQcdmDAjmiZXCg11cTEY39VrbIrBGWKT13TkD5ts3VXNj4/VZumq7oMvY9ymRnj5/FN
YXLBk7hOpcYB7qB3t8HbExscU0+AbK52jvn9EoAVttYp7S+qymLnysNolfg+o10AtxhangXnNzzm
1KfhTC+LBtl1KmcFcqKsMrZfMbHhm6IM1D/fiFScIgAns+csjVARS8uM7w7YpdWWPjXOMAapbD4L
rqwjYR91lU8LHRJqiJF6X1mNTIa+M/CS50d9GmflvXs9t/EaoRycVuktK3gPyaKy4zOVigFvlKTG
jiAjekFGz/tKesPoFRHCLjD+jKnen0J9dP9NbpkR0Jl1Fl+iKWRJdx4PVxiscTb7WLk73g2BXFZR
5LclOUhK27lGCq4bqSes3g09KscL9y7oU0XQmJz2MvBE2krZhNCqGzARg4YqnFO6sZYcUDKW9w7E
lC3rZe6gelfwOj069+npTlJiAL8eq6hFfInozJ3Thd959mv9TwU3jT1mHe4i35vSWTf8UKA0zY2c
k2CDHv68tfv4dI4emvZQZMIlOrnfN/f6BRppssAsArH6ti2jMfSY04EWOHKqA4jsOd0E9r29V0iH
W9wEGQsB6hRtW0S5B6Rl2iZAseN84m/qscJiliZHhUje0b6JlFsgJduMUsF29XK0QD5/IgOxHhon
mY9L3wemG41JGIWjxgl0fEpm0SsEPTmexQNv/EftDddRCOAFvS8qc2pJdOSJ6qeMV2vymcEeBk4v
Vj+DXDooYuvmuJZ4ErLHZfK/Wae/1uKn+ByiqUuiAzJu8/b1lIhbKIsJn9N5pWTIXux6ChKf2m7Y
vsbpnBc0gD807omSQN7ys50aG9G01q8NB4yEht1SIxNVKhmvnGGE3I+c0qXZ0JNz45JPe0XyDMji
RIQiuAb5Ef5L48ciIb8xrTFNWYta32Oxqc5l0LLBGx2oCZsxbuV+2wD7HjS9srpSvezDwRjlvjad
A6zjvb5+JBcOY5AIJby8ZnATbtLzi4+UZmRySYuc90PDwXAxGrXC8zOYNcNk2Akb6GvPQghdXdLd
o+H4orbNJfs1BgoYg1dtM35HfghnawX6PI0K6gGKtsbx3b/LmbT/1GwtxbA6KtdkzpSFnMziz4p5
33Z87hd/I2ubsNsBoWFiaTdKHDKP8/Gl5vHrM29lmQxgqHJUARbHiw7XOGGMN17B1ta/BowPYf3B
jADUp7vfotV/o1IE353Tf7W3hg4OOeLqKqfHJITnwayYbLDivTz2756+W9Phhe60zZjyV21M0wFn
Fidrpf1XZE75H6mtb+mdUkGbfaOmdSwiM3HH4MXUnq6P34hlBEDXeS2dIC0mn+ltPPQMF6i9C65W
Z/mDmlQeSLE0C7SFKCo6dcFWL7BSkxz7B682BioHqe2ZIonKeWA68Kokby8Nulyj8FICmhCAa1Gc
gpaKYE76AKKP5+FB8Z1VO6GbOAnnD6qv24tn7PMq2tBRoMeoTvIr3689qX97ZkK405wgydscEldK
rfYUuJcZoNuGNg0ixNc3PP0vjkG/t+Y38EJqbM0p/JkcyoLjxlP040uIZtic3fsZctwPwxSyorTc
ZSgqUmwFrokgOLP/2G1rIiZgJ5bDNwObn5gYY+M0f+gNRN7yocxHyVteu5Io02ITllmlT7fhq+OT
TahrhMQn/6zqvtaOw9Yi+2njiRQ6GWEazDQTK0KmZJkD5Ir2Wb0RowEdM6Hd7D4+kpwWIgH/W2Xl
nCS0RaSl14t7G1Qo0nLYXqOhF1jY3csg0QHH/rZZMApUodViSIZITGLtKELMY13ODpYHByrFSmRa
JOEHs0YkqayQQc2u9vYH6gH9/9q27G98CVfouxGe9wf9ILdRYjRbtUckwBcDG/T3p59J1WOYHIEh
8yW8DVehke8waT6T3SD2vEXwIZ+TLoJ8ueNEwdZIIMw3p2ygdinE6S4PyZjHZYR2HLZSh02IGI4J
dw6j5pSZQuZL0h2NiUOzvWGWOoM33jVldvBGonAqnaPyHuUQ8y85eD1iw+gnzoMc0gJEQxSIlsOm
YE2HshhkPtdhfER0UIRJCkUcguoBmi2tAo4Gc6/rZ8x6kKGGpGBe7WgfF6WEoEAxxY2/j7mNalQL
Miw/ebEkc+z3qYb8u7Dzob+2pPuJgUMrXXw1GJu6nzaEHeBl4MzZVkOWW2l9nw/Y+Nzmv7H6qGyL
obv4ZesMiBZ+8pnQ5CVOJJESCkj7vXLAfIv1oUHrxgHn5G4PLbMlul9LFm+8HpROgj6ad1WkzIfd
Y/q9ysUkvDWZ+8IHMUMR3uff33gnzIcoSrvAo8xOll6OfnVOd7YXqEpqlcHwS6k9f6dP/LeCwcsj
PVqhNHz4VziljMb0M6C28vUgl4NO8gzoF9ezsBHEKZDIaOMXX5rUxmsgDgTG/0ORv93wifTVhZLG
0Qa68f3uno5x4W4Xs1ZwpRGWyHL7dbDMUk+cLaakVenG/TscgB9YStfpmRO+WIn62zIKVA1fTVt2
xZzh7FbyfAq+dVXECyuaG8qdw7U41GqAZtnv7bRVkgLrEtvNeeGVsFtoMFu5C0iis5g7GWpKZKjP
D7zVg3SULJdVoMZrHxbppj11M67Vgl2oogXNnBqeXYzpkKvyqWopsQKsMYmHOnodNC3IwFXzCBit
whNfZpozfSTa3QYKncVVA8o6+DkTTOAn22nuHqGMzqpGHk+TSZgbSHJOmdCMxbPKaP7xuqV/ETcr
VlLsdCg3mHli0UF/MdIrMoHoO4eXyDxV8gCYPooVMSENLy+2rvbHfRbi+4VlrdS8XkfcztFfxi7m
eQk5bL2TKvFnVf+NRQ36cXRqmZGBTOhOvy1pUdyAw6PJGjymua9qMUCy2k05c2PM1bCOvIGrBSFC
ON68sz46Biks9Rs/tnl0qNpntEtRMVaOqSpQ+hlgOYwr+qREQIXzkalC9c/FlJMPjG6ewMcHTXnJ
jxAayn3aUrdfRwdUBQhomI/E9PwbMxXx7R+Nbogshd5wW4YjY7n20PkZ+lwkAMyqhtGDB3frUD6X
J1Ha1PZ1ZFVq2+kE9PvXhO2ddZUtglMSQBb4dkAaF+WV4MqFjOVA7V69m+IUX2qA2SdC0Xp2rfKH
/duD310VOshrWRXq0RaNDzLUqgILm5dZ7tp0/rYGBGl+asMDSu7xKJ0EaIkSDBI1aimkzlp6yfQX
DoRAfJUXTMAB+ZioiMAC3z0sgH/dWwZZzYbLKQ7tUTQbJf5R1j6mbiVsO+KNGXW+vtiQ636pOlNb
aquu+yaOsj9w5cEGckfs3EUAXQTcHrPh2kiA/bfPX51g8NGEcxooZMjAqUg4TPYIA+W5EIr5RNmn
buDKa973KFKXCsmocPKsVRTTvY3+eJomlITBUnX5r8O+ELb60HsCjAM7RswkAsTThOBG4nTWJgAR
jlzIWjUEi2Wyc/iiZfrjINU8RU99G8gCR3cvINIk29NzXh+pH4ditOHA1dqwSa3sImmsBKOKroOM
GLabDGs3WK9WKtuYVfoMH4AydsF69omwzMlJU475Rc/mQVTmt+c+pPGeGzfdFT95gz6mJBLcNTBD
pnHLxg+VWTzOFa4EwElvwge2MGa01GxdaIgC5KvgCDuSITESu25rDw/acIpgtjSMhI55zD/O+Gmh
+Spre1MJHrl18jAx72O9d+nlPZVeyPQAEXPWHRASvcC2BshXYULxzcyzpAhFbno9Jmot3GVlAs2N
bajoUbxlLlLzasnr5iwXRgcG5hzwjcV83xbLqzPZ6UlYTWwzaAOXYnglWii4UKOrORIjnH6Cg05D
iSIbaJd/YM24c3m/n+j/CAFtZK1pebWZNIYRxyttfumrrc5V01OSsIAZs4KbkcD1Res3M5Db7Y+/
kdrqDyQtMpg9a/5c7eV5cYZ8HInK17mso9BLlNJPvwYNDjgXsa5/1Ui0+Liv6zUl3zQ7MrppRGNQ
+zjFe/MKcaPPQqXpY9ckaWtqsO/oPkDQZspcehqW8S5o+pmgv9DLshPtjp8flx2taeqC+yCCw0et
2HBpWZDN2HZ102QPi4zIo64i/j+lHEjE7sbJL6RSH0Veohrx7CrXqiANNbRfSPXxzLXFg1xEvhrD
naMo0S4jVd+3MUK7OHaXdofiUFijdfMgns3846BAHGvOmSdqCpoFq78xW7dbcO7IycIuMAeu5OOi
4xV+2aaQinaGMDhne/DLmX1kHjGQwERxi4quVoYabPzbjmM8RlZ4Q/D653ud9zrYtKdfNpBnXbb4
+w2g2WlutBfaCgDO/xbZbMY2M2kFIDJxsfvb9anHj5+Bxuhnxd7NjPaj/N7tx2OQTn4O0TIJy2/8
8CyhEUr500wzRjsSyLq3W8TNLeW5o3Vr+CQHBd1sou/e8Q053DerQb+7wvmchgqazrfN0uVNskrF
gwgEHLBC9IXH8PxGqTTtHTIn1aQLd44LIoGai0TT5I6EWPkT3d2iDMA1XBHDkK/d66REblwupnp9
aiPjIgTdqbFpKhiS3p1C+RMytlSO/EGxnb675aqyr4eXUKJ6nEcXVWheOprGscXdlsJK+/4lIHVU
JlDR+G7+5rjD9rQkQFBdXouBxbkhvfYLsnE4DkvH2Fxth8NmoH2oAphvMlZt9hU1U98uJIUgtjG4
5gmuigUM7S8nObomFAvp/WCaU7JK0PBT/FKF2FrJiDROclurpFSvlLNUy1IbizGapmbAvLZJxuRR
WnbfLwZgskmyCebNk0VIKX/8tFrxCmRc0rdEJahFs9KN2TlUJ0jP/orUSfbur4WLIN8yBCLCG/+6
5lupJKHeJnbRpRcGMlL+lXs6HB7+lBzQSq0MkQpDIEvnUH5GvxMzNVP8wZoUzWlUFrneIlPMY8cn
4FW0TVpnJHNld+Jvj7Fzj4Xf2yU1W9LqCS4tGFuYsUtAb9b+StEu+WrOSTLF6Dor8Ek2MWn/hAVk
cL0PYzuNgZen9qzZfwWzLyR8D1EH2pSW4LLsLLNmJqEX/QzS7u0h0bcQSQd6httjJjv7bwRncLLS
bTRM1ul+/6kListzlpoETyR1qdLtSVouvVsPT7wJmv+Uin42nzHsBaB45JqiMWFUzIR1mTJu9YBu
Mg9FXiVag5pxVLrRL0cEjmDwzqz1LKKvjKytDQSzT0XVIP/fiTe27Hq4JCQhJAGOO3uJ+Vn0XH46
QFHl1NqIdeLrYw7XdeT/L+2fYBwJYlhTWC2NvSbT23tqZvLVUGJj/QGi1L+DBqoWg6JOn/TutUxp
YXCMCA+E/LYTVTmVS5qZ0ZlKrfSB3LD0vCJcwAAmXuXWzqKqFWisH/hz2YavEl0RGK5S+bgETPiU
T6E+gkD33NGRIrmzWtdF5neb2zcZWH7VzmIGLDGx18BPj5RPaJE6wZJF0W83HP+0NaayBLzIeTJr
ac1wvElRjOMBmkAJFavtA/tMYkO6zZgBOBaEIE12DL4xLuv4LIldmhp2ZZiMHdqTrAiRzGzIFZNd
zm1uOy1YTdA2CClokJDifk5d3vzm1gzLFozBpqbyoM/CwZAjY6hOhyHFB2D2AX5/Q+gHkWMtr2wy
C1/xJRLEEYDERX6B/3ZvzEyazn4R64WOTis2YA8gEaDaEs0x8/cQ6aJedHG3Agv0B00yoewrWG5H
bpbHGH3yIbsaevkpqiiRwGyiDz4TQbLFKvzDYY8x64BebsZLYh3CxivFBVS9VdeI0Ux3gIz6xlWq
2o0or0Aeb+FaTWVOkO3br77ZT+2R3o/Eg/nmkXsWLPZEwgp4QpxGNoAr3eCh8i2KAQ84IOB5cZMg
LmNAeu5nNKVv/pwB89e8UlSq5GrHfjey/RoqvDoTDxM6K+oQQeD/+6mGr4qWxXzc+Cc98dok6NDz
Kq4J4hif5O2zO6PVOtoKHZ2Pzm9erU0HPti2KBJ+rZNI5DXDPf6lG9lE/PkYFWX++FF029egt02j
JuSZ5Rl8I7Ncqqg3ZVF44Tr4HSBScfI+AC9Q8BCxk6TabjZXlXjO8Lskk+uSrcBHAppO+Tli69R1
QMQAMO+gV5W1nNoXEWm5VZPt86NOQvflWL7NthnFP5b3YXF9smVTzIVuYW7NiE+Vbepz7mViWxKl
iP/xz+MpyQ9XNF3iy7ToMaRE1rqCzHEAHmThkVGVZUif3N6KGyO98lfiG//yzTxIQsVleVEwmKBh
KkgteHSjtgDNvNfsslGMu+E8yh7uLo2JOLfeBhUREiJUKeavNal3j1DBws0CFR/UeWlzaG+9GEjb
yPN0iLU7+36VK4Rz8e6MqdlzshLuWJISwwgDTmP9wc8ViAAgSBMcL21+ObRsL8Y1TDsJZmGlvQBt
ETMhoCPNZcCcek+71LWDEzYp6LmI1BFx3Dil0fEhpSF9tFqMBE59HODgr4VpOcf1eTCKp9k2UfxZ
S9ayQyzkHDMxY50xHyLuNUBFfgX6HYYHAxicw5wPjCA1A8NnH/+3Ix0RdIndUugT41wycZTHWWtm
EZwJlHI8wo5ZP3NLHL0kspoCNmSp1up/Zab4mKgYEQudGpdgrbHswkbYJ6oxhC5hamYSVNt27jso
t14Gye4MFU7piadvFuGjCZH8a6J2qzE766HKdtMBBe5oGfGnTGqAYGbbVn4uaih4QnxY/4LdmkFe
Jii+1Fh74s7re/f9N6w3yMaBcw6eQ1GkSVwocVNjT6yIVEuaLrpzwCNJ+wlxx0n/9wsHXAdFlyP3
i3hDR9Mo6dyIwnKwe5C2WXHGo8FvJb3t4pWSEEwWVY3dESQ8qX/zv/GbrkaT522j7ahnrcr3Qoli
RwanCCgv46UvQ4jT46Z7Og452GFiiei4Mnd5w8cdm/UK5auThuwAc/c0ALa/bOBXAg+agXyG28O8
8lBvjYQ1qNE6hyyasOyaP+CySvQycTu2Rhr6xxni79T2aEJiL4Kv5vbXY4ECPGqFVn7McEEbuBZ2
OUpVWGFNGKXjE+buXzyEiyrlLVSlWAnizSp6UdHCJ4kXe9m/mL0gM/RGTouoLUJ8ve1Jq0V7pqSr
hh0GNwf7X+HAZKFQ+pwfUHyg7ynqCFZ0ygHR90BFLLc7az7DRokl0dCc0MGDGFArKGCNrBKxjaP5
GwpkoZ2RL60PJTQxbpxSaDd1/YSMIjn3HxGtEoT5bgiz1aXGya8mKrA+UuxBzQgKiKORQQH0FEdL
SM4HIeuggvzTfx1JM6fQ2MJlYubA7tZPxGjRp/qEXHLQ9kZ7kiysPxtkcR/SuiHkuD5dgSsqEU2p
wTc5HVqiA1m1YgIai6lEcb0j5CtUdGUTHqsB0poTKROWAoZB9trrSOx/bbv+1ZPZ7HQYDv6tjoFR
qOSPYJmvmtx/paV/fCo37BQDZrEsk4Ev41Wsfq5UCcyv8J4rklzmTeEg0oksPamJwjB3+Y+tkTh0
N4BvRnQ3WmAmNHcNSwDpeDz8Vp5k00528CJP6lqoqiTEDfYrxCg4HcSkPYxpwYzZKxtGW5hMHdfP
rM5QlxvN7yNAI6e0xrQep78084aJucB+rz6V8ROCsy8o8VjfMo22QVzKcOa+kyeNwRRDxTbDtQhI
lrQ4Fv6eg7R9IMjhfU3QJLM1gCNuWxIvd0NpeQPQ0+NiF77bsUvVRJVd6S4C0UJi6dt3Q+Zokshq
GXUe6hxHLZmiOCSWtZY9ndxu+fAEf+E3a4IuHKmkvpTwMBgUl3ic8UaVjOKBsVJQY0HAdMu3tP1R
kyXboiA2ztimB6GbbWCBCSH6FXS+ZJfXoVv3n/qMA+wD6Tm638pMNlKXO4pKkNCGpBdufXeoKAnR
s0Ac4giaHfLyZ8BraKfm4SVh1MdzaMB5x8zS9viqRboGH0wBTJrHQXbjLxJglHjtdYFk97LlEIg6
s7Is/nVn1ZsOLbz6NVZklw2vVHc9xnNP/zeO0mApgf2rmRvXFnqK3MDx0+66nEf10DmCGhK4Yhfy
sWZcyC0WRq7NC+yELHQtoTGgFMYdXeWeo7HytvRXhWVHGDCXkouqAzRW8YGRKVHWjbBmrYHiD2pc
uqV10ILqniyfc1775ko//hONvrts0OQ3PGXNJ1QBuZ0QnuyOy93g4qn2x/iFGclkGquM0HrUPT3e
0jsHtrT8C3P+PAHjY4JXYE9Pb/lc6gUd31Fk1KetilB9V2PISPLqzZKbKEhJrTHXvUzRGqwK6lHo
CNEvexEJ3aL49pFrW4UAfY1BXXPr6eHdZ3Ofi80IIdMrjiCVYHOZCCkDZn+8XKWplSNp6IQEnIup
TqBMf5I1rWP6cD1KFtN7xvACG+p6BRsJRDv4LsTF9H3pGpiTxsvrZxdGOEkdygKcpBZoAm3kClXF
m/Kk3XLMadmdf97C7FybtZosaUGh7fdKMlHvtSywBoGTJnursEEURY9bKdpQlHkn2TPatZTArWCr
kNkUwfvQ5aytaJ64WGk3fL0bylcZVAjDzkMQrE7qyDMxEdnx8lrE63vaLx3/PJ04zoZSta3fzuHk
z/qX+vpVgLJN9f0n4F0Kan7G1RM6H18sdzAKjq/UUXztV/H8v+/YroK0SaGKTgRa/vzGf22A4LNu
zN0TecolE3ckkKkqvU6LEkrdmSyYQgcCFmg//65bFo2IPKY8GPAEN7G+UxNrTPmmPkhZVraMufHX
WEeXQgBK5zZCafFxM06GoouEtLDWEMWmfBfHRN1EL/8aYYruwXaSGArtfI9tA/KbTaNGXXhlhUJ6
3rhX6TO+AtMaub8bikA9QJsVIXBN2L4wyHKS7gqi4hKWYVvPtwY69Ws4NQtb9h+yns18SdnwxyJK
GYm7sunyXJJT5bHl8d8ogDfz8rpyNfFFp77Kg3EkqAKiuBEiBoUagT7V8ICduRX6xvJ9JI7a5GDt
bIt7cgDOesqlYL7nOZEJUcCO4V/k8avfxWIRKDZSngFX2MWijpvuSnkPbjbfLHw+qo7XGf7a9m1g
6+EAuEMGcK3KlFFFzhbAAXfSLe1It4TAB+mZCVrGFOgYb/Ef3HMXPlGRceD8/c6DXl0LIE3xGtAW
fqppG9f9GlGxQO3AN7217r36LuA1Dzi8CPql8RySneoFxuGICf9MFO6laHSmgIa7O4pcvNdGlp5z
j8TR25krvFckGXM0lYYqw2hnMSAsqj/vvPSmlP1pMDENTCHyaxo8mhoP5RWe/07y+y+1Q+0A+Iu4
N3ygn36B610M1otzQi9HX81alvE24oC4BO26O7uoZS/bS4KZHKt/kTJVlbHW3iVZpUUfihVMf8Vf
Bw3wHvCb9i+YL+4Tn71/uo8xtIRkJ4RSVyYRliPgQThFwL4Q2lFL7k9McSsATgeQEtgRGUMQG3dz
nTi5VzOPQ3UrPQD/LraOmUy3ifreinWHFJZXAUt1yMiEqIO8C3XpDXHuu76BjVcg+JYo3frzZ2pF
U/gaHGaL7iUnZaUeGORMpwwJECpotG1zHSzutRDQEz4cANIrzP6sVOIi4LGoITzl1o8hVL02NnSA
qySETCYvRIbs/h95XHN2+fsxUgrxGqxI8pjShQf0s53gQHn/PITYKi0B8IB/WJEXlziMniQpWFhp
PYnr/YLk857WifGCOFujAcYTKfsct4PHVgku9pw01eeYtg/gvdNVHrTiRPetappvQs2TJnuBAzyn
w4xRSpyNyMjMrCXuexKO0nZu90cjvx7CnourcqjwPhkBJw4WcswMMBV0pfQyRcyTzZ3Ass2IWZqz
dGQWCNIq0VZi9XOnkIOWqJeyNQoecotsfJaSKEJe9K7cgI8UnO9hXWUoXGy93TjkIz84FMOiMJ8a
EkX40h+Ex3mWU55CH7twwHaEbYH4zW8ai6nxWAJUa5XBl6XYrRCGojIl9xRl4MMqWNwuHuQuNAF1
Jp0RHBD7VvVdp79F9BkeMTT5bADoj9CkWzCEeEKTfUOCCbVs2gPRmypC/KCukyeyhh+vAGe+qLbH
eW7oCVh9KiIX5dVTDkT39nIoJw6LZfzgW8oYxpMLcQu5gcpsNGcGdq0RA/cV6kSusjy3akzPZjYu
YOjLuWeXcj/X5BLvPlX9JZqmLk+d8p9G5+tTPPO/NRaPtfo2SmIG6xHds6rS+z9WNJ4O3J50kFqq
gvqk8+bcbYK7suD/TVeO6+A9J2/dtx47CQEP/bq3NWC8rEkfc4zhEh8XyNQawWhCZyM91lNmsFxG
Mjz0OXaua/Mtl9aJhv2EBBehX/4KkKNhW8qSL1Y1xtFWpAbwglhgJt/FGUMd3scv1NNkO1R447tA
J3ToeTSJHeb5XaRjJkp91rrl6ajmkA2zqJTD/+nqXZGDW0QXx/n7VGcGKAhwNTjTGbiAzPyiD1cl
scBd1vUyI6AXlDVYBveqU7axVozxJ4cU3acuyr84XWV9Qe84Rq9zrpB5rXbq2swjUE5skFzxchq9
mHFfgnkSs2YfQMWEBSk309BeEl+9PBlVqNEb4jRjoIOfgb8L0+bAPzPfFQvKbkrgLAPtnrrehY4i
4p6IJSg7WM5yRiFiWh1ZPIzTn95MlAuNyuu55+WZPqPNa1hGTiDeTJizLgwUKl27D2W0mak4pmX1
vY3i6qI3mc/povBLgKwSw448hyQhgdenIK1pXA/xFdLaFcY94PNkTcnigCw+62XfVGr6FB0I7GB9
fKTMGO0lEECh4BU5hnzdn/T/lGkPd4gQK9mTHCb+hh6ecVe8ac6JpByxeZEhjvUj6fKxdmqkS6np
2GwJEoXqEKsDWa1JcJMG49uVRAlLStGjVjDo3P9EXsDB9irrKrMl2os2qdmOKpYICi+UmhO1vNnr
w69mhUYKbNyaXrgruC3RfMkL0ZR3MTU3M+83OJ43ivCv+QKAqBRcBwn1MyuAD/pFu4CPtk0k8m03
kB009ehnHFv54PZuc6sNdlMKDNOL69pI0PNmTgYgoRlOU2vEQln3/hklynirIQEpTClwtW0lTqiI
3MLqpowcRSiA8UntOJSy1VxiQvJCaeCFRn2Lz+36UombBRgqWmkR8biT4wJa/OGENxchYUUBJaik
XawOdQEIZ8tr+j1JOMYJGiaqQM9KUrfYkoduzEl0UZ3bcrgfhrUOTg1snxZaB2b7bsgRATB/zXx5
tspyOPpcslFpV4SSRCVWe9+Xo8Cx3tTP4K/93gt2RaXx/k9lCnRbYsYI0NQoJo1cR8Bz4AOn9tEq
ySNrgytCPIb3PQpKehQSNhgobm3j04DGTnClAjF1fb/aAV+9v+cg+XTj8llxY736ceBF4UeErcik
QM0OTL/Ixxxq/9SCH5+L1ygUT++GVral9HRaQYmVGRS51KbSt+4FYNCB7W0uFixnZ/tFQ1jq9Bds
JM88wCkfyDt0HKpfrKqWYqBzWNId0tFK/e14Nh+qCWAZxcN6zGl2fsnDyW+BYCwhpE/Amx9emb4n
bnGJHexSY6Q+tkcivBy7ueI37JQgJzhzuGr34sJ05Ol6A4bebxa4TI76S7V0nIrl7AMj2wAmdoKj
4sxTYGdApFrswNVw4hjfNHvQn8UbQd6ZfHi1Yl8bblq+o2FGf2pBJJbD0A3hr8xjj5z95PhYnePZ
J6KpgVzNL15sOxOc7dq4A/AIjVwUOe3BJX2irGx7Fl45JYPfbeceJv60N7PJrbwL/NreOzt/rIoo
5J9WaQkz5ShLiFz1BcPJ4iFlWboesw8Ctfipye+Ho4t9CnUItWFSuQflcQ5+MPNDQRjLnFzkTpkD
iWrG8YDAEHUYuytUdDqlxlboEHujlAy3Gm0qzFas1lFW7RccgW1RQYIOy423MoriZOB/ehvGyqle
JKYzIRm3+45Rt5TNCbSLT4t7gChKRAzEz5tkx/t//hBR9kY0K8zhurhH1NftrMf4YVeMo2tbSsIQ
t6QeTEr2GdPLA4yte80KjWsFeCp60tZEktnAOjlNA1vwiqGXsDSHrgEAu3Q2JaYd39yGfcrJvTKs
p8/Te6G0qFkNCnwcU7c2o7uG7E4EniXd0lPqf6s7BZUCjBaVeir8fgKVLRk/QQKLjC+B4rJc2IyS
/8JQWCc4fqcpYWM6dvSqF372LHFulXxgXKg/2E5b6CjYF6U8W2RbDbzXLjXzNwWsaYNK5Nsbzq7U
OJGOV/iFuGCDq9JuDm7jPgT6LdN7wnb1oI8pMrVwCfCVqoDkqvCkoa92BdHYarIxxsZFEFkCHXoE
x6Zgkm7zwmS76doD4qXJx/jaRzL8DdYs0HQ1N6JiLSbAFJNAtPMy1kRV9Xll1fEeNSeXc2u+Ukh7
KIzFJfHy1I84KR188FTqn+fcRTJPGFFCqOGvkQHwiW7SOb8YEx0lVI+9jq1aA+41to6DT+yWn2Wb
h41Tp9L5wCcclwkh0nKA4Y3yQBn7lXEYYnHPd41AXlkZaARDT4/mLvObQXvTVunkpAFgK4bMQEF0
gvkasHITmDM7jJW9+5ULee+H/GX2ddeB3f95uYSu+WPGCCjQVVapIy1FIsPjibm3sAqBsY1yH5u9
/D8D4mzasRzYIMW0ZXleZIPrDGoHkGa+tEWZ3E8/P89kIHp0ctOZcMYYfQpZnv2D4aX/TC3ThPsB
+E3/+D5JVheBJw92TiRhhI367pzsYaB0qVA+eIOpPiQg/qhtJ4KZmN061VRUjbNMr9ArbfOAOxtg
SLxSvJdO7a4RkjUtbdOqK3u3lrdn6aM7yuB6SLFMY4YhqIZQyd29HsWooOHoP2zuGzV1D4aCX7FY
7QjTxhkN6uC04leKaL6V9owXWBp7HTuo2NFvqOoOE04jbTT5kD6v0G8tdbCgxH1T1A97JE3wXKtS
RD/YsUVseNImhPF6FrfX9hak2x4M9GUkDkV9P3KQRbqv7ddzwa38fjPacLs9AmAOCkkiPeHrrwac
Q33XLWUZFAxlo0JPrA//LBAELGqgk6Ro2du/LfggHUAjRyfGXRGJfcXf8rZpsoi9f3YETnCUeqZS
jPk/VABAW7+uJvyh4UJp2+NgVTSu3L9Cp2J38+8TRCe9KuPCwT6JAW924laTzOd+EmnzOq6WjFX0
jNx1vlDmnpIU2A1ImLSZGtCPxYziODgKZVNSjxVPEpSA7qfrg91nA9ff7aZjW50flzq1OPOzI9qS
OkFe40wRXi3xTUUCWzxntABnWcCXmkULREm5FTtBUa4i4dgFrZvLIlUrwWn/3DMjKYXQM+ihsInw
JvDJa3pxBE3qBU4QOp8YsB4YFiWBovjKszrlvcXnGqrb4e3PqHy0xnwH5CwpYmt9eEcddgxHaiUt
rPq5qGn/3wCMUKBtxtM+uV+Qy7OVXtY6/TdQGGN1OzCzMiic/aycox0mw3VCVB1J3X9vvhYf54y/
agm8MSaUAkfO9l+rKsXWz1VNNw17BrhTxnWeYzzr6BCdXZ1P2vGy9CFrge74Cpr4LxyQI9IdHFJv
Hh7HYdXgV/nyZVhX6D2xmVJnqc501M7j3Zt+GufglHrhMSDJQ1MaxaJEl+PKIsdtpdUzlwsej1M8
SrLKwVAJXLkchRm2g4SiqVESfCK+qDxe3YaKa7vBSttMY4pUYedLFDP08/FspwHxFMCl26sVuXYq
XNtuOEvO3dGegO1byvO9D/w5f+zwGP4oD7yegQs05iio2v0ePRptdSR8gwhuEqTKmESL2TN1hfL8
BxYsL6GkaVPJRPbJZRgXDKXftmhpKivu/SzJVzn6IER1aP0gCXL+GKZRdB68Ud0GpGgEFMc4ba+j
FxfKZ++TNEWfKtLDe5/P3yAN7aeqQky/u8UIEBMt1gk2nrp1VHXmxieow1gvh/abTbOOxxPe8atP
CgyYMyvHlplKlkfrqd221UXspWgp9+P/FJ4aoDHxyF5ras9b3kEjOB3+ZrjH1Wx13OpjRHjh/Jsl
nqsgMP9eeHHtXdpBEtvrN1379H87kflwMsAkp16ORd3vti9sSuASneO80eM8IkAZB6b5L9RRT18q
ngYeagAakzVFKgonIXyrrPlzfG5xsUGMAZ1/0eFl9/cGO3IGMqDRpO1OWJ+zdYWzTFcgq/yNPfvQ
HHtyIoXmO44lg8BPJTaA0vIAmfanGCL7Ha5A2bCgKgjrqqtsqQI1xZEiduoU+XYvjPJHzMFRnXSJ
Zvy12G4KGD/DCoco4p54IctiHMwbcp34EyCm2Jpasgn21r1DOINkkTsJ+gKUeLNjSpqJpPjC+HLN
M7GapyB0aNwSiPxFI+K/Aj3h45DvHewg9+aFxplIovSri8Oj8wxYfGAQwnE4/qW0Mh5KJfzi7gbK
X1mGaV/ZWJHm863ReGWsnAeQOkHbTZgRCXVF/2Ud1nOeQhG1/uoPnNtvN0Kv/3cziY+4VdKDGQVP
E9oP7sIx20/z+JKdl1gGovSIXAI+Retwk49EDNWVYCqSHmJT2WS/8JawygyeqPQU69C71DCckghf
DHDR0D/TPHABTWFo1CJZbKz8OJmmsWhQBGzYrE8eVTOvehFJDSLhfq0GNOAN64XI1jlZlubMaxas
6ViU43sCG8W/L6+jOKE06STemuzM0mBP3qtIevYVangp1jGB72JWAE4BbRr3TdzpW2UuLu/LZUkI
E+dDUsiuXuZD6+smeDBl8ildFWVkcDK6V+qfKp/Bfqh498xCGCcXF/ZNARKk8Gj+HNaR0MoTJZZC
cWhfHtNHGj8rLZHzipWDIkvRqs3IFGDwETe6pkM4AB2nPx6wg3yqst0/cJsOh6B8cRhCTOeJdU3J
jSfH4OLlqAqyx8cSpmojw/aN6SBQH2GNDGV1N/K27LyncUsDyWuqqMCc/3TKdAXinN6/ikl//y6p
O3o5C14qBhdFRplXLWr/IpzkXPPEm/fh46axr0CclMSwGwIANhlHZYAz0c3G+/ARJFQsUfW7Rl2g
jNKwhS/l8RgMs5Rg1x6lChSuF0kgrciRHxs5Kbc+wRm3Zix6BH6IYFbTEV/1iXDQ1dKGIoNADxTi
ZmhghuyhHCZ3hIO5aCfsyplt3fLNdI4QgqwucUYD0XF0v4LeSno1uFhIwJeDhV4ymG46Fr2k4x1Z
HFJ245onTk5mquAmycLxa0AWH15blPugXtEXaylUvF+Lux81OMguvhkQjhKnOeU8xcDd6GHHbLrV
1oKcnx3nsHvzEETypGpRLkA3FWi05nCZKzqtXdf0LFTrdfAfPl/80UhKz8n90BzPWXl52KEbwTSi
Qn2+FNEN4LAnf1IYh8xa8+Y0s+scgQxJ9fyuB2tL9tR+5ltARVpZmf/LoEdth4RWhyDWacrObSho
N6C1IgZqThm2JECbB7hOPPnsUkVkIjqiQ+oW0JOHAYp3S5xLO0EwRniR2m2UNMwFWrSGD2lF9GPZ
fjGv6tTu7qHzorvR7lSTdbmsfgvPhR3ei3STsrAUASgvDgtZukbCwJt8JyX/bGJdbDKUgBfp29CT
P9qxGqnkWd6sKh7iVXo7Xs+irZ7xoA0U6izWusjCcJCMP3WO/iYX/6XYWHwF/9WvxHVQwku8tyC1
Bxnv17j5tnGqYInqmOq3wRHBCDY8XjOjUbJLd2d7pPVhp5AQCvDv2U4oJxBF06h2G3OVkhWm3MnL
WGRu9zFJSCgM7v57LGn9qC/mtJswDpz0NZvrzlxjfucXY6eOB9Qc2oKjYZQikBGFRpZVp+0ZTsfU
g+oMEGfrF+MZ3ZsksbcTFmfOI1UpuripF1AEAGksJX0rRR5K9ApR2Nk2SC5ADFg1DujOTKw9tObo
OrLw83IG71Fst+Hiecd9O76UjBntgptO/480k86/y3jU8b9hagru+Z18T39+tXND2eI+SmZWmf1s
AIonYMCkj3bDTV30fiAUI3vcE+f/ySo3nJtPm4DLIalUsTtjV1H5k2hIl8koU162w5Lplqr458i7
OXIMAUbmq6uFbpVxS0ppRzT8AdmQxZMzgjuxGmUueDCzeNi5oh0anbLu4yP0Oyj3SymKvDovlBnf
LEIwuVSBfRTImQhe7vFJuKwtX2ngZlGuUVbZ3fAp1/rP08KlB4oaUwZJjhYQL7TLwEQFflW4OD2k
4tywFqB5GkaA0+4USt2R+I4iuehCpLMuCWVJs9OkCXurhTG/8dUwFprqu3pzWH/mvrtaFlvHDg6X
SWLOrpKvmZGRx6xeoMI8JwpWNzqBS/bxBOcuFoHI42kude3eeGpNVBxYIGmdOYTd05o5eLpgHBZF
Mu55Jp5QesvCITK4xmEjChQsRLi6FOB/Cm+CpXwvUp1EmWpGc7OKYrRsJe0njljjAaoLJVHClUeZ
rwrIympRTqKe4EfdsYNBNS1qnLUpO3yhoGLSWwsa2pzEf8Mf0BueidZGuaP9pcEBO0JREm00h5ov
FWN2PeI4WO2izi0pBUzdubR2jIZGDnOGhDeej2XV4qTHXzg4JSFYc8JcvxSpe3Ixms+1hC6iXxoU
QhE/nWZ5J+ryotlXMCm0lyyntSXe5L4KXlIuJmLw2gs2cb6kOg1k1CrSkfnTd95Xgd+1/+PNmn7f
L0iy7f3Mse8z/XkdAGjkKubz4Ql9BCjDcJFcJYGWyh4lEqsYObUrCdLvZirC1REP8hXbXzVwGjtv
idCqxDtPTENvxjyO3r+dkAJ+yUt+mfc4zwvYqvMO9tlEJIgLINvPsUhCLxEwCWAY15AOiMUrknlP
9yHIERAPzCx6HPjMWTQJ8lD2Vcrriwx6mWts5+gT9qx+8aRLbyW249luU835CNCWrH0f6Sbw01fg
vVdgwhdjUR1cOquLn5xJBoqSwlWhBZfUFVRPq9+EibgtFnQg9wIfVTfuTftptNfqtNWXXZGCpz8P
zj3T8T7F9nvFChB/pDUxEbcrnkiC8ynhiQ26pKk/o7QDBxUnnSUk7wKy6O0xsEM5ra6s89PWlIJ5
3MoVNPSWBPrC5aJqRHGX/ofr7Q5qXzXqfvkAIH+vZxM/WkebnIOIgcC+BS0CvaqQTQW3p1bPIyWc
V5SYt6bCveTLHIEnJbSYlICA1wiQxOEDCg1AMHw3cvCkwoodSvNK8IbKAWYB4GEjYsszKutAlG79
9pjvjs9GLc0nRUJWneSI0iICrpdlA7FcMSsFOuU4hbrnUZ/YZnaHPM28+3khQZO6HU1tTn0R1kwj
uHNsJxfjxy8zE8qM0mOv7Ug/klztgIHqsYtkNRHSCU/SmdvvPxM8xuI68Zbtr5+vC5z30+jodzYm
PMDlpz91zDiH9ZfrZSMVsmMPZuJzFmj5ELqkDnqir8vzJpIBmzZik9fgjB/Y4U0jr4kCgd7abjfN
hf41z0/Or4IaW34DDO2t0eFoVR4iYEQn8wacEURl3NhL4qrYcf88mMtpaMjKxP/VGbSZtlKUFuQb
Bat2/wOe771PCaPc/aFuPuKEBJ2EM1sPf0tObt19itm4z+t/D2hFSx6Tf+txFggjq7mHVuPOznK7
r94fOr7KKw3j3f7oPeUWTn0RXLcfe7+U8HvKvwYs8Nf/IZViw1ZJnrnEV5ogMxMa4kfSPNmbAHnW
Jgc+GsHMr/8iu8LNqUgYdM+tqJxMeHOE1wnqZvemqiPS3V9k3UghiNkA3AM5SOR4VYYtksG/p/fk
DSDzcYPvRIFiLljkq4G/nKb4WUI904oiU8Z4izfS5Pw064VC3r6DoR4tuSthG8zX0/Sw+9UK8ths
XNUC1ePmqKHasnu8QIJQEmuU0nPtO0l5arRM4NurG53Xg8kVhm/YDAu2QVKkdjSyS543r3we0r4a
o+nAEc563ae4xCG6r25bCGDeCktsLoJULtTAdEzeoxvluJexbHhMduKQ4g9lRkMFaA+2ggqZ/+kb
uzC2fnOuPB0KXL7t9LTo6vriGS1rPQMt6ArUcSoTYyBiCYacutbmkFZlFUzETzi32eDkOJAevMH3
X+kQSSYpmuv+HkabeMTo6iOMJZ6D7D+pfiXfmZ7fHbCp45HKa10GReg0YC3mqnkSg682Sid0ZTpv
mV39i41AVqAYC+lEDe0F+VNafw6I5WDSpeGhtayAuEFSEzGLV2Hwkgi6jLh5/19PgGfVv0Br9XmG
vlKt8GbBmKcC5S2CtgtyZqqkbDLOTh/AGR1AUwyPjrtOTdK+EptAjXWoZjWyVnMAeSAkeV6B54/X
Ya7tA20cSPmApwVZFzww4gwKwW8R/PhJNjgWzarPyt8ACaZ1YtnKH41eKJiffWaajpzkWbEWhaab
5Ak+qdwr3I0784wpUV7HzQzpyStFiaRFjIFM7JG7UqVhxAm/xiFx/CN7LozAtPERcgvmPyF/baxG
fxuwLVPvZbvxVu4ZwrfsCE4uVOsZ0Jhr982sBQugn6h/7pJgV4ecZIy03RxnrLy/Zrkm2Zi4biGo
CfRX8166MrR2O8PbHa5C094lg5oyNrcEtDQAlAOOTG4geak0EPScZLgFJ5SmUfgTzt04S1W2D5k9
gW+pNFsax7Ptq+IDBJ6/MqpB4dlU/8s7TqBVWiIHflTrwDeyPKE4zEJ8h2PalQtpHHIzWUddH/T0
IlVn4Umgm6EtQaIwYYXRsVq6cgAV3OAVpyOwclN+E4jHcVwzqno9iXkCbnuZhB3XjsPqdtzkrgSb
i6ip1ylIU0F6qJP0TepiWutFjMHnHtQ5Bb0i3at2M9Sfb64oWzSqnTBsYNzi4WyD4nA/chF29vEA
s4dFzYAQ3FHWUYzdL5PFG1JT5/L2gyC7e/Z4FG4yavTV3NlFguhuq7qwRkPDa9Mgee9xdrZnoEAH
d1eJTyVBdJq//7MKAgCI78x+SkOIGDDKHe07TIMePJzGK0sVWOdSLIR6Sq5HgDRSjNnVZ+8fOSRP
PN2scxpecVHHlUQTOALlgLn7PDBU9AiGh0OdKUnkcT50pIkWj1wiF1/XX4019q9LJAS3yZ3rsWJy
7xs5FPe1aMIvwhFsYEpO7Y47ULDwclxakyQWt9MHhlgkK/sgQO1pQ3O6IsUt3bnFmYalRsBY3srV
PyW4jdpLS7F9t/ntv5iCHkZG1H57Et2hybWwBP58sduAo915s0x+ahLjvLTdb162mzoaqT/jEE79
AWbNzJL1Gw3YKbItksB6Q3bCWPduBQ6+Wq3DPgQKgRbMcUh/dkTIUIk5bMTCcAQSx+ZaNnCyeg6q
raSEEYAmmckq4h/qJxUrPDQMli/BDFrA0J7d/laBkEmO41pGhrscFnTyobKtvjSb2xyvOEnUi0dN
fPM3r3lC3V7D3uf0gAZHfWv6jQCA/G+VoDpQFtnewuwz3a+GMibNBL89B4X+59N0ZjPDz5DT67Fb
xwwjc4Stmgxx1nTZCq6hEkSMQPcmjr5czwgJ4hxzj1qIMc8orooI/CQRqabzyCtXPdDDaZb4+ZdD
2zVhnbJ0RBAyLnI//vaUOXW/TI87DHbZpcDp1BJbFtz2BaHdnY5xEVBZPL6ltOek0lKeGE/K68WW
zD1NfTUvhRV5DsCcKwr/L1X9QVCfqFFWU1AWTGylKZccEXiAKfvHSqm7L/4MgnlJX+9zAp2MrhwT
ciyDPW6s/pQYge/uLZEOIK4dk+o9VR/BcPWCx1V+gw0peqbJ7RX82N+l2ETklDa38QQMoXZ7inuF
bPdYm7DLDBytLs5TNUoVhS8v0QtY15TnWmrOnkJ9SIRf//3CXF2p0cIkrn95U6LEKip/NE0Xyl4r
3ko1tvBfvMeESDFfAFGhpYz5V09IbBlnxNjmseojkSHyIE+py2qvbXCyhc3i2WLcSME1kwg/8dzI
izsX+ExDBnf4lxZCvB3TlOLM5yM6z/6KbiL8SbA+cKgkryz9Wlqitnf3MSuF396EVL1dF5+hYU53
oRUNKw1/6qzcVEEvM1k9ECpBwyc80Yi6eFnAvwdFqw9gP0s/hM7CIMw/ZVgbM/ow/SRgNWfJQh1d
N2Uo7IdB9+iaJrnAJ1t9XzCRAUMKCsTd0QjIsyjB3rKCcDEcHvkPGj4PV8xBa2qjvZrpJRwd2i2j
F9PSg4t4/xPwY0S4yIgHPoAblh6cjQ5M7KZPNmixO7Yw0RQepgQWZZ+lDsb/R/t3SnFpNPwFzim4
l2mj2fGaSMlZaDg2pcxKiPQOaJmVg2IP0DtRoUy2cnPPTQnei1E5MhbgZqjScvsXGoCS/8iKN4qJ
UTvTAE7DeGIfgXyWv6YgA2QwjhDWhBqS33lhozHjx/IKuDiP/Pqpi1GJIsgQYtK4eyJXxvDyyfLN
hPLXzgRMHXIaR7wFnFOMUNyywkPoXTr0re2AtGWrr/ZqL6BPTDvX0dQv6vMeV2wwMBL0bHAQ4qvh
5Q8MMDX+eVvs+ZPml+IN/KziPFfK/Yl0fl+Ov5dqyQE8quYmvazITGpxkLuGwyAoheRqTzuH2ips
gJ7DEPuoX3a6EWpgha9j8OojszksiL78ksDOyPBf+BuORkDTzFwb3Z8sNivrNuL/vEx2SXMtbssX
fkoDf2m4522xrB1tJoXL1FSQDs8d7kKAcob5Pxki5K7PRIc0L1Qd+hWiAfoAJfmO8Mz70Npex5TD
zu4ZM24r0fJ5TiL+ujSxzx5OXCaB6xmYbJF2PC4DWcp7jzNdzLxG8SBD1NuGj35AcdFQKUQOPEJr
Wa/pDqNudF7/1fYIa5MlbWRtZw64c30hkJMmqFnLsmkREOluQaZSIFqVvsCk8RH2YfQjYntqvjZ5
9hylOlQKVKw6VLWjJdx8L629M29TZuAi0xRyn2YWWiqZHPPsHKki3nNclMpC73af2zXdGOlGCCN3
4Xoe0vc2Qpd3zWwvVPiyDqrIheOLS4V3q9lrUp1z05Ur7un1J/GsYemWQHXp/j5d3FM425rJwwAt
wcfn7FsjtD+UwjUlvmWSCw36hDY6EPzTGt8YnLb7ijclHR0iExIJjaCNrUeBBE39w9fOe+0BKzC4
68iq77qPRSWQcadRLersaMvMzcYYMz69kAsMyaxBwKPSnfE4B0NVwdGNglOiHPDJ08pj9uiJofsw
n5nlzwS5TxJblhlqE5AUHgzI/IXiKWKZ1rx3MPP3aahydu7Rafk7HvZwZeLXxma4gyNQrzOzbImf
iZ+9muGH8OH95KYh9A3EY0Ai9LLQJ0EWhRGiInP0WOSzZTJCWTkyrviot04p/TR3jk+FwCWx9Ykn
zU6xH7uGFXpMlYnNKPlpEHXtpkXJlZ7NJ+EBz4H9sUIKB8gLthMBvB9Qcgc201nzTrLNwYi2C6yh
AjWgOGzHPHd7NOxvqe5k/AnC7T9soBcf80iaoc1voxYSDKEd1Hm7wugbPhMyi5t5s+BrvMjURqAm
ixIMJS12nvD0bPxrD5KmnUZONLpBN2EI8HwbdILq8oDojhVtWvjjIAyKj+cLdNagUofGYSd9Y1SX
YUJFfKtU22lyjUMxUlTeMv1FToJwV+fWBcWgLpn3gS8uQrNcnQxae/I80fRVCzOu2f79WpEAWDAZ
kjGU2o9S2vfOOauBXleDtiVGsiS8VwFPwmTodr/2tr2oopuP5F3xwwtjnPQ3imzyGIv++DRQJvf7
DBAwIQaXmrE0I1u8gCK5HYwLygqnka+jk3wZdxl+wNFIo5oiPmLQmaNQDugiKdMqIHJ57BAbtfQD
N1uv9vl05MQE7mbCH0EaCPqXnSCfLsnutCCeMYs2lNJGtrQ3wF1nchN+hTOmbazutjE7N2JhLEXc
QRzBFZYaB61NJA/jDgXV5DS+4OnsotCGeOwl8qHshfr6wFjobloDn3LVfbu9IJnVHm+MLwf/72qv
k/RMUELcEi4cs9q58ZdAscU/41DT6pdyZhrJAQWcndYzkJQZ8LIkPCg5RCQSWAgaASGwo136dEq+
EHaEFK3QKS+D3Lo7GP0YZ6cu+y7mM8kmJChjeefF4IfU9BMpR+ld6y7A62C+3xLTToJbEc4D1Cmj
b/QEJLUZGnX1qEA2zshITbsyHhWs+najIbcPdtugbgLNIwkF3CZcDM9U1SmszA3RIYV64JnJo1VB
DwpxOnVsosMG/EMOIR6zHRVIgDFf8sRD41u7xNgt5zWiFRJNedvP/ijDAHFRYFjpmX8MhDKSI/1M
UAZKKFMnmNQUc7yKYE6teb0+crlLTm0cLhSL+ypSPPKjYbBmBROOfsdg5yhgaps185TY6kpPLtTl
VyHLhU2yD/7tF+vyx9SyXeSTJn9zhyqucGK0dqUV4vClkHG+KJHOZ6cdYUW9oqZ0OkryEfqs0Kdb
gRlciwme1nreU6mGkVSzyRifIWHjtiW49OF4nErUv8HzVhnx4FFRD0VABZmmuVFIn/+QWuNo/2Ap
2NrDRGlzLGhxuEcSx4nMDYsWNL4vC8NCjKZIieR04HE7j/+3mVejvJ64kp6KfmkuN0QoLStjFgS8
WvG3AJA+kxUyIjhaS/QWI3xeWIOo/OE675wuL4mTezMHJZiwCpqgML8mML+FRgwHDVrF50WWCmJ8
mssQj+pNpGyZ11z6SPFNGzP8viaQMF8CN6RONISPf/mqsRnYoSxu+v/uUPc48zw2St/KVKhQkKcB
tj8VfFfWD9GBDjK9LATWFNi19dVaA4MxeJEKzR+nDr6BMBaon4RIkKxErIHsZ7fItEIT8vwTygom
WYT3Si/NENSVgBjTJrNOBDW31AADXbH36n1ujp/btUXUeMwkxinf9/+YoqguLOZWiDKX7k7GNnzq
3NMrcmonQL0v+P+jCHiUS89RhpIPxTxfGojBWhLbcN6voHtG1SAocaMi6xRynr54UxVLyAKNMveC
NjjvNbEY5DFZJTLxA8DCULJqJpU67A+BQ6dkydZELS45nsnwi63pA2O7mYpRnfe/f1yv/PIDXMBO
0+iOrxlzjcUyseRdcWHhq9UoevVrpy+h86rmr6W6PuPeIo771iKMRw1wIaYk0KhJdq9P17ZLiRe7
AWB8p/qpVw/x7/Gay1/GUYOQi0CieVQMyYMTvT5W96+qDdu3GKmjaCZ3YLLhCPGv4tgmnNE5LfCz
gRUBdv9AxptMeBNlPU9J/CYoTtupML8L4aQ8esIwKwOgKaFOFD4AiO5wW7ehH9zrTOEy/Qp/HTd4
CIJz/dqqfD13MGZZjU5LQahZEhHygyx1XnTJPuGOis37mayrNHAJEf6qsAPabvJqP/UlTntSDE+T
n5RHw6y0E1ZTjGn77qPMOETF3ka/CMAdNVb67HAMK9FE/ob2l0ECNWzFLS2EChSB2Z6inSPOk8B2
DJ6wp9DE8/hsHPRKA+0ADJ73zbCw0k5wj89tJIvwnn93PmQqYtH0YXJG0Z89xil6N/bosOf7DO0X
xTDbkaM4CT2z6TQ9tMcbwXVs0rYyrR+joJpsml42Audrw9XLCkZkAmnyHjN1T7R/6yR8+iKqwkPK
6/z13+XqJL4G9q3l2+X2h1eVEQPZ2pidR/rRLkLAdFAyTfupOFyjR4sWRyjbBPO35MNvC7w3PXk5
WWv0YAv3uC3uluy/NdYCzTh5QPzxpXWe2v/3T9Ow3laDiGW/ope+RmoJsv5IJbhaWqDsq/Vy4AuO
yC8eQqHMaRTRPj/X6R6n+VslvrLsx131wbuMzHcu1FWQxviUvEgcXhQQjr4ecNzfAwMmYPKXafR+
x7km9oonB2Fbprv1fyX/zzm1ICeceYaHkjMfQ+ca7Lt8GWD3lR9Hdg9xs9Fmzc2tLYsc0ur3TIgn
xnsqax5Bs+8e9wqdsTLe9fM1CzHFXC61WvYolyNXpo9ubmHqKlkP6DQ/fxi9k6rjGwiatKLICSAA
zN0oiqy1rOp0rXKmKgbrc58vKkzofMsw8YExTkun3qTDV0+YhCaiNUan/IjRjJtq9fCBJk3rSCpL
bK1orxdf9WKjalZvDm1xIgahNXe7f9Ggl1EgGSt08tUDUXvWPR2R8h+Ulf3ZwCweH2iQCsepFpCq
Wrzb+qOlA11WcHOcMUektUy2I59syYFykpv85/NnZPCiTWJh9dUMFI5L19jHOdF4sRrpB0Ussv0k
R1a5AASfv9JPQzDm4AM5YKH6dekLTbXYW8VmzxceAnF17DAlkE+AKjhXiLFZ4J91NLIfT4GDNOA/
7P22PYGA11B6Ai5a4rZjPBpiYSWiGc8+KJV3ZDlODdm2LPHpDtpPCvyzuObBNNcI9p8HrXIYGbPH
fu/fW5SWZoFHRq4fVkFttON7ZfBEVVlV5Pfm7P8SCis1lmIOLRFW8ULkMWhllMrRlYvet8Gy2vzC
miQJ38EtgtJivBSYmCxkGHUtrhiOa/pg5mgfUzRH5koyfkh8cev1PmPlTpP9kHNS/19BosHZL0Ph
ZXA8uCDhiVbyEeT7wrgObG5dfFyzFYNBk53tdEoQCFh4hisrz+QElIv4yk74pD83frBGYV/hPkYi
U6NfK61iSCX56D3GEdQBWmMRWHdrqwO2MzyXfxrw+svGw+ggr4phLdRIzpGJ3xc2z6UzANdJdjE5
o6YRwjQMv+ytl3fkZ3u+Yv+7/gSfKxbYQaBcSjHXgtCDqUHotibnLz4XBXm9VLC6JnfE8dSmAqgq
tCcV3/gqaMh48qjwsNslS+7QUG38hLVhG0WElH5eYkgT2rfu3a4meNTZAb4Z8Lhrc3QwDb91Wa8i
Jbl75EEBsmHuvX6jmG6lgcUJ5Oo0GfImNdd69Dn+nneHFpnTJ18ZamjYLxjvH1JB7B39Z6Bta43C
Xi1mCTCJPNKpFZ0uLoXHbgB9wQ0swg4TDiQAXjVqZu30VzN6CZsJh5UfIvZVLWH5qZYxUJ+3kBXq
LYJXjaILK5GcPtN1dc3Zd7lwFZLJMN9QgwQVFzwUU6qCDmrNHKeT5wBjTX1nAUoEN9AvZOTZnHIy
htqICyIMwWxKBu/6D53EWunzyf3DOOlbVL3NIo9HHNYDvqN4EclwEI93QbyzTSzusSn2fGuRTLkY
SwDBjQ73UDEmjWh5J+sBpKoZHR2HzW06DRlGBHS5Jsxhurxal0wuW2duwKsth7BKcKjHpvJasC1b
z+c40CoJNE5N+XAEyHTdPg70o/zQQ0gXi2RBDYT1LZqSuMLHvLFAF+KB7MsARG39w4EFdc3GozXX
d/S38pyf6WDPYJei2yn4+i4QUsyllHyp/Az4wPSwT2eCSqpEdf1cKXuwDhdzqatr6K6rcot7KFFo
PtOYW2zO0EQKZfGu6bc5mvPUV8SykoGvVaRyg4reyiHzhjpnSJLAuGY93PUz3c4yMuyKucPb6moJ
9qy89gyETARMQLcKteG22maEjfpTGYUKnNvjVOsIhJNiHdzGZD2GUFEJJ2lEG6u3F2ym5U07A3W6
orcj8qSb30XwIgNJXwdBlqFXVZPOTOAuFLgMzTdGbl/3h6K6rk1nV70di84NIEaS25kfgfdhqyOj
zTG8jnVca+g0dK8VBI/ZjdDgvdpRiFpcdWCFAVF3XuxZ1mi7zMR0C1Bk2mFRbbczKeR9JZmQjM70
h2/UdfOd5b+aeu19c9DanDif1kML6NAXyOiJop4gCzZGsGn0Hx1eLKzul98AuCc9Om2wsrOuVyxp
xhLt+VmkCSsfQJ/PhZWTXPupjEpcAVgfro1ILo2XMrs08g3OyTZ8dzQ0A0hsiVguYEcNG2lRPB5k
TooCP1IFUK1dceY1LhKrmx7E15QPAWgv4N2yQJxms/G0rIKzqx5y/UcVkC/uyhVkHeuXxawGpVo7
4S0ylDCweVn22Q0i6jKdDMy/D+xM/kffQJ7klO6VXTc8CdsImkdgjCEZZnbIKjXQPxE4Ljqf2ely
0bF4zKx4mKfhh13yV9gH76wZcPeTBRBjvad+FKWRgVwgBhKH1q6QrQw3QafLmM4u/yUH62JoYFwJ
dbmWc0N6IOf9Gv6Qq0SnXKxJG2TmK8oLIOvjeM8la58UEwqEh5XCMQHHFSWoc4Nt0YTtvhQaZMGO
ca/gZQCSZsLf+iYmaP8zv3uECO6/FgFMnbCU5R7Ufs9BCoeYyM5xw4yLP0RLRS/mu2OHWJGvToQZ
iY/HgdsqiOPTRyz8ikWRllJWdevBKTdfxRh3FoDpI3cnescuwE+odimIW1P5RK51ndg3G5EnzqPX
Q8duy1MITkMx8Flg7Ea87pROxI086aRSzkOI/xIcBcj9dRJrCCAXQ1jfmo2TBotabJgXRqnm1Ui9
IOgvKDE4UdbDnMp4hqzC0BB4nvrLjAkT30Jk9zKe26at9D4pPyvbK+ty5rmi5testzEHtQrnB1TQ
NlhtR+/2Lk25+MQVQMcFp4WBIjwZkZ7YDiyThV5clTAS40QK0DmLXBENdvDJlUEEtMClmL1TGCGY
3OrwqDsrXmY2HUkZA9Z+DLJt5awmaIGVTTKV4rAWX3TpuXX9WZJDWqrMbpYwa4hrFSy+eEoA/Wx+
xVSGVpvS5RasDuX1Rogud4jFHA3jEC+2T/EOi0ZHhAfsREsM5dax7+6bz+1VNQ6uKzxB4bU3pooT
WhqOM3NGniQtnoCy4gAzrX/d64pS9vdwtPCuo3XKS3KnIxMas2G97myhE9r+8nLnWyWFoKuynwon
VaCXTeTruoAenEWgvTqUjGOziQAVAIwVWDwEbQCfDG9JnBAlvMNtxl1I1hWS+seQe69Z2pPcsmQo
fWq6k4sokmFFYdPy4AAHczNrBHmycwAPyryOza7tpTyF3boIsP94RSap99PwMdiFaAfSmS4wCWPL
6TaoXkRXdA+a41uIkJMVhsG5KDLc47p8mTt1E63HcAoMqTYw+mM1HkE1CuwnZ9dmy8XPOFcNPmz9
OvLoiVD7JKYfyokWt+8Q9kdAZmeUKJGIWO9c/Jcx1w6DMcddJ9NNEVBjzyKxptkEluMCtBFt2+Ov
wls17J0S93p11xF5qs7tfhHfjlMA0Pg/0BmZpgYDzjsyK6I2jYXwrhTw+Z/KiMtY3LJ24WRXJc0U
alOkRlW5el4DqLH1BQOKI2mt+sVswUMDXo8D5aIedbQVYoa+l9/hpUEyFyCrB1T7TDVjhDcTtmEG
OJ03g8up4ILLrf+PrL/b5YEQw0OTdUou5gRsKzckCHoEhtn9aspmhMOJxery4MwAkV0YB/eEW5Es
PS2GfumUO9YDfqND4ogG1P7dqZeFrcji1i7Akbr75AiS3dkP3abbwJEiZ0riyGsLeKSJEoFRwBML
R13wBEFqGpcHkRrtyKCtAD38s3gyzfYe8lh+ProNxHmu+WF7ECi8BRkF7likFZNkcK4fqTL00Evd
VCOU6trkSqtgLWL6GL2cnGaQTzbAekZVDLMFUbZtpAHW3Q7zoUs0U22pWhltLq1O2+nPo67+YXIX
BrgvPt4dAPelDigomi9OKLwIBvHOMrAbR5I/dZ5hJIB5BIqy0brCme5tXVwXFWXjGFu2uPVLQbZe
Q2JQgNYOvuMW1paxXz+yP6N11PT18630vjZa0DwTTYBU2EAbxBzvY/16AlHhjxHowyCpdAFTAoky
8Kk/sgd9vhugYxQmhGE66fPsJJidKB/sa3XabGuZd7kue2mj+a2UPswS6FZRAK4ZOwGRqocUb4hV
U6kV1puhoJaiMvzhbtq+nJjgQHW/b/OIck9K22FsVgc6W6UNAd+2ErWOawSpAAbqSb1LONVrUNJy
Z74CWPCpKRu+jDFfQ3iHDfy7+Z+8rYYUULNpHbunv/o0l4+Y6eB5d5nFS+S7GVHeZostDgKzmcRJ
UARJSoqcAD6mXVmJbyc0Hujr/JiRz3YjwRtoG/IajxbfaGk17Owgt7oUVasgF1ujU+L5zizRhizo
nQOpZNhbk2qEIv9l8x0VyX0HMceSSUw6oh8EzcLHcb3kIAxWKHFxd+Bd3ywI46Ix/ke0NFM9v4+p
Kyz4h5XEvhQOQz0lmfx3AJwhpWCnvT4xyqoj2LauBl8uKkKVGNXVHeMXIxgczXalQcZc5SlB+1mP
bJAZ58S050W9Oazc/CoMbU+K3fczTE4uRNER4fohfAxb3vNJyBALJedxQubr7FrGi9O5XpjIG/FJ
1zrD6amtF1/BK1G5IE9rWow14QFh5SfyHeAxQbF7Kd1NTudCsgU86Aug9udOj0a0B9A+757E+tz3
zb+b16xlwpfYUIEchGhM3jhpk0dcxunb+kNxrY2V6JKKcQj/aTcILXiTwqB86D3/GpnVkE/8U7AC
cKPHqBuEYsVWb1L1DRXuw+gB0RKAJVmXGY08o9WMwf1jqSM2IVXFtAsQKG0AKNFAnMpDwN+kjtRU
ApgN49Fmg48HV24QiJjG7rK004Gs0FTLE/DC4VAmpWBVD0G3zl6uGVsyhhEp6bt45+7H4PDdZ0mx
4h5EIyHXEil6USnt+7WGdXwMwJz44ynlijLXlKcMTRRIY++IiXIzta/yTCxzRNRBLx1/gb6QOz61
frX9Q/aC0+KS3RoRAI5TZo3qFT/hHcrI63yDPbXnp0XPZ7ulVI5YQJAjQHFpAvWlZtliS61kMvw/
zLlvNvj7dFa8lfTHl8ePZHb+t3dorCnQhyw/nFry9TzDshcbywrXd5Dkz/yBBqFZai15U0lEnEFc
MWYKZKaMZSb4Sd22I8+ECq3LTRLG1mOHRP0VGijk26shO6CGHvzgmkFI4oGyMA7gmAwqzafUepY5
97z6K4cUVrPMZiG/ZTZegSbmx4APZKMzprDgfYm5HG5SUSNQeWmDpSwc4MYzdoBYU5tiPbcuMWVp
J/edbygkgdbeCQhTc1/gxVIdCfVUaMMPkI0TrllDdx1s+RFW/41ljL8WnJ7rrbtji37B96dUjYjq
xQWt1zNwU/dpGQiYdERIBs2A9kF5SgJRZXZxg6OVX4OyYxOqhuYfbO0EY0qi8tkzY6mh+lE/I9T3
JWuiVFFsq/KSaay55IsD1BYqQyEtOct5NGUCOr27CiWT6f8ZU70V/HG2mHSLgI2gdVAvnYmoY+MV
/J8tDr5NueCoeVKW4vtd8dXkod9c9KSjBmjzYKy/zO1Npes2ViBfLUDo9GI74lAWvF6t137lFOeN
qg8mtZjR08lLy0I/hokx9UMbXm9Xo/57bnIOjitZpOFMAd+VDBCAFhLfkPZIMj2eGFGCqof8FvvZ
lexQuYW9KiOT9x7+Ey1wKYTEOL3z4bRtCLsXYGgqjsSxEt2NdPyHXlTcRM4xsG2xAWeYvzBGk71h
gKvlwm5dsP5gH/LrkSJ+Yltv2cCmINh7vXvYq2K8woMmCOjOb5qk55eTkHtT96MSvSz1yVTau1ZG
CqfL5zCiuXoEh2Niw0VqtJV2mp/OMAupM/tOYKoxuM85gTSd3bPlHJU60SNsMoxyvxFyqpypXHxT
gtxx/lK1a2cfkX6fqtW4i9PULf2gDQM03q1Lc/Xu5IF2OtsnN7WQ28frsP2HF5giuQPbPVEGs4S1
6otQ2QrywuRuxhgyxdtVgSetayins0nWFx/s3Oc3d+7J09afNBpr/TVWiJ8XwJ8GAIDlTUvotMe0
3YVqZLX2y9Tu6AXHm6FqnPkoxPQ1mUg80h8JVXLWWB0FO2PIdVDWtwC6N28sRqFPuUpLygV09awq
ZnV12ooB1atsOKm8DittN5rz/OitWY3bX1BBgny4INKDF8UEUtykRRIwdEqlobTEwD975DmxGTpi
sYWn0mOY/nxt3B2/1r6fWrWJKrcVzZp2MWngMqrPCPWOtIIsgjVQ2LLH4R5ARnRLe+jY5POASzZ6
MG2/MAevfd2XbpxDxHpfNGhxgBmDoxsGVY7IsZg0pVY6+X0AIhwgq/V3Pej9n+OJmnPoZ6Hc3sAZ
MEXMcLxOeNVoTRd/v8jkt5yHCqSxKHZNFF+U9I93dxa7SJTaJCntMS6NMXtHqTMN7v6DP1ecdh8P
vAsMR0+ogWJRfr5Ny8xvSsCggyoyNpB513o8pX7Nle0fbtyPmZMOrRvOUPaod/dp6pgzzxlaeQX9
YyBSe52xiG6iWa+zr5vsayQNzsyLQtK/aayi9DF9NjK7GlSmcUeakYILOpWYyXHgJQQOu7EkW/mQ
TBkXt4CDVXKaFz4YFHK6FzMp/Cc4iQmYA/yT3WblZ6VY2oxoHMmprFSPvjJ0RqwSOfMgGoecYlnm
jwdcNYsEt0W6ZOGQ5HD6Wlz8W5Nzry//ymiHHzgOFA2AtnHSS9pVwfBwa/JNshL/mZjKneqRCzny
CI3OP5XjiVF0RW43NmofAz1hEmdyJSQGD54Sqg8UqOmV3XlcCf4NR8HViayrRDDufvQ1BLIZJwA3
pEhtK6XqgblDS6jXNFHv2eLTfYRXxKjU/r961yk8gSz/RU2D3+INhJOhd+O6UpSg2ofrpbq/Z1yE
F2hb5DYqsEB+lR2yGKrGND9jdE0+CE/Jhmro0IR2ifnwWcQ21jvnx3AB88JoKeb9qrcNKlUEBt47
vJJUf1PSWlv4XMFIMdoPtyCIYk3/k5cQW5S3W1E/yo7IPeYkMKIiLH59ncj11bzwQC6sLAglTfk5
vBou7tsNqCeg4ZRQ2RPc6LymWCoHUWjYmJIMYSww1J4nf1iH8FtkWqjUCSrZcuXQIy/Z24F/dTeY
uLyRE5c+Qvu3zm+ufJDIQqh/zL7vX5ISAfUrdIn3xuQ5fWzvdefRSC07T5REZfN3apkA7gmAtz5G
A1M0+Nxs4lOBVLQam9I686hTPT9b5t6ZkMrVjqFo4dIEeiWhp8Rt/uShTxTYJqKf9Zes/VE/qITk
zERuoPeTd4LAXH4u6qxk6BpeXa6gQPKByIIYcqYawMoOnGfGxBMWWKdQJjgUWIjZkJsPPK883WMZ
+ThRWctRKXFTPxr3kUNYMsybv1NvlYLHqAMbi9omTA4VeQ2elwpSqGWORmXN4tGT6Zaiukwo/K0m
TUsEGUk0RpToJ++JjQfgrMswQMBZO0CCxjLofyZKyWs2BA90gp35Yn+ftnKb1S+Ua41CvyaG73v6
FY5mCVodGKv4H4EBnF6ofB2bMKdtmFovSBOrA6B4iEYU5+8CSr0+3sGxKAQXwG+rnIuIzS3pJKIr
dlfxExlKwDYxgHFUCDtAqk7Srk+guMcZ88mt3OxdzCeXTCFFxQi6ZtXb7rn6PRgCPNQBpelzosun
EtGWPOS9apkxgR6cr6vPPD+LZgCI+lDuggWSNM9IqWSM4+yIDmRmrW/16GxEKd5JTm8HUiGtI9/u
tznuVdrtnmePTaeabGEn0HsTLzurkQT08Mt2YuudSbGnSB8tvOe1aUKq8GH36I4oxJcpBLJp0dca
98wKJE8gHKpveLnkKjCBvVhQNkoFpdmGlWpkYw/TBhR5syolxonTxXFCJuTDh+p3tjfFUvl8nxgT
CAMlSuJ1m3z7CXsJtVDq158N/duMnIlut13bNoCXM2CJh/Npf3KnOfMjrSMdLhHbNHA4lc7WzIs5
wo8Yobsn3UHvX2i9osrgYuzUb7gPCRC471BaWk74Lh5jM0UmxYZlJfnWt+fDfUbPQYV7bIIjVRSA
OZgGnKWaQycZO9YUgfQstU1dpBrilltwOI4+/Er8F8QLrPJcrO6ULui+wB/x0PXiiiztEUMaecd+
wALR5p2Y754f0DtestvITIs1rBtp9tneZSBysmYCBAH+o8LzG1065HTILwnhE8szdcyW+RB9yPPw
yGORNIyadJPCQ+bMtuCTJhJfwJsgwRHbHS9Z1ptMLQ4PW7DN29DI7Wohc10zH+QLX+9JC/6n6lx3
mDR9FJvXRTTOsit49YiAIMd3pW5KP5x4/0QhB1tJwKwyYHUD4HyOZrMd+tcCUNmyDAitOy3xVdif
KN2HGwaqJHSpzl2c3T2bgayoebSk75Eh5rxtgOK3/fEbRnAmgVwQovq/TMd9VuCop7kJ/ys14016
F4ULvhAkcuZQS4EteNO2RbIghaCSkYlw9B59BFWcal7AJdfpyyd/ltMu9uJFv73BWWqAvdOXlr1U
eXn/1BcYPSViGzaLTbSFppMztgO3ka4rADp8F6+coOnxI+Gef4zIk3uXgZnu0+LDGC5DGP70x8gK
QNbpps7IcsmAH2hem5DIgQ+jjjN53FTEwH7yXj//vqva0jARJcoEF7IMioasuGuZyOBiR4jfOpdu
hUl8eYDN8fYHzD6OnG58YfbHvHS2QSwk9LiH33w1pHDDjzC12Yg3KWJWslZpMO6ShDu2XzNyH3HA
3YrdBjBAKUT2CmfukKWDYKLhVnznuDUpz+9l8kfGa+6e2LJcDpRUfJE8+xUAWsRr+EiXlLnHiHne
vdRNg+EqDVLWxVZSKrY5Re5IQt1DFTcjJIVZ7qRXDBfNNJs/aXM1oXN9/3iZrAJVp6GrhUlYpLud
nHCX4bMPy8YB08Q68/hVRxiT1xRs1l+/a/Dj0B5l9bFmoDllt13l8UdW4bIFc3PvTV/vPb9dy54q
/LL30t+yTb8YIpZ7n2jLEls4SaRIJV2x2cVsyonfGA5059rAAxX8lU0KVqYvcSLXW/4gbHEIKmdi
qcNacvihhs6nOZOObphSNezIlar44WzmXJow/Fa6e83Lj8msEPUMXHUTzMgNySbX4iKJdc26SK88
Ia4ZxJQO1tlbPCtAapKSms1o4RKuuRkuCcrtkyH0C/JQzWml8av3xqBy38TjTGxAsuzDBWO6JLr4
jtB7RrpXWEz1+76Iz4gEL21NF9Nyd+lqkYyqmOJkebDCP0mZSmCGEZoGYETMZ2gsBeQe3rPK8KAC
LIZJMTawpPRsylgubgM2KK6zV5vXUJYvwOLFj2b6tyKZ+CIAYLwz10hQn7CCNK2wJsCc7GNhLu9J
pqsaLndjOBUudhIWuZcCPtuDurEh7u/oeYev5lEfBA5WXSTDqu+ayYpDrIk/JYuvGFHhZeNhy8FR
HtgaV7ybVSnI0XlKCZFAsDLC4IabgX4dQ53Q3oUlv4wdUzoxgZY0xa1oeZ+/tyFJ5MTDX48OQ4o3
8SSmuXdPKWz9JjSCeUsmhBe3KXOiGqJP+Wmn2l4AjFUM67Pi48mlSlFcFCx6PZLJERunB0ztKdQC
TWRZWqcLwt52Sye9yWvguBl4Uq4SKV+LsWXWbYKv3jt+cLYgrmtMa8GAR8lVRmccb31gkm1hSumu
L47HijZedfbaYCGGdopxDl3WLgRAmly6tjAYLFM1p5kkHtvY6lmspj7XqX6PEJ3ZP9Zy3YYc5hwV
9ImYE1dXO8v7lUWmPKpMPA2quodlo9wFJZ1+8VH0uwKh/zTvHMPC9FVxCU6VRjWt0GThLJKqG/zk
hjapEZp0jui0dOKXgVjvEZkFTNaNQX/wOkLRawBIVY6UWRs3K7wYwfeTbo9KFaRdHDzBswkjg64f
L7L1Fmpdv3Aqt4DcOQH5sm02YLMK56mxfirVQRj4gZldZmwF1K117smzTNCtup8Ocp35FK2hl6FS
YeHz/S3i8pHEO4ZlDrY8NXDPMR1m9YI9F6wpKuc0QDHSEFW7IPVIxhtLE/KmICx+t08IFc0ZiFWL
hyGJ/rZGt7uGKYIz0i73Bg2Oan1OWDI5iZtAA88ZEdRktKgkS93DWq7SA7+01jrvUosQ3kVz77So
eW0/MdAUnRdp/kiK/70nw5+0c8sRu8/K3Em12HKFnBOT5KNDWa8RA14aTOxLz0elhHib499Xgy2k
zXDteNp6TBuciFxI8B+3q9CjICl+6jrvNn4MD+eQcio3mURJA8y6CkGfEDY9Su/btw5W24ewDKXm
IYGbbMX6p811OfxUEovJJKs3RA85yEpo9ucExBEYQctHbRmTnBD4MuORkoAbKdAH28hSyjq2QoE9
0Oy21Xg1KnjCPD4ZBPm453acxX6QCxxbB/vyx4kX5mVIw3vH/mG1MXRJauR0PT68/TfOGmTc/dN4
L09Txsc7dJITaeE2f2hPe21S1KF287tx7wQ6k5P6CgUg4jTH+G60JszVDPrnaOC/3eh6TAMiDZV5
dkDsRUtHT28E2TgGsP6plicIkjkC+6VVU0XsA86wO5JyE1rZaYbifle8Wn8YEorDouNkNo+yI5ZD
wSDAdKLGo3pSvnZvt4cf1XbXMvRGsMHJFMtp1FL2QQM7VG0h70WqNFYnSZQ286N3F+CYGR5JfgPi
9o2/9DmFRyTn5jRNlSsMHWBFqoBRjWAC8CVQw0d/ZbUn9tK6ssr38aayj7s/aAq43uB1x93ohded
m2ubWsaVdTu/eExgR/X5ZRufRqFKHfT6ESn7lA6tQrpUudByh57Q20TyVtxlNzqo880pU9en3f8A
ECW3nGMRYnAKRxA+0AuoKkERfVNNwNpVZ0F36mp6JRNjlrkOZtzIKkWtg9IF9T2vat0Wy3X2dowH
6IvuBB5Og5Zsgc0x4Esah3qL/VxQd1u3QUnnthpjkEmwvdoVirMZd3L6u7+P8hfyTu3pcpGSvxBX
oOwfAaevGPFz4ajvxJZ4+mR1OSdePhLU1IjwgV7AABT9EdTUYy73pNe2+5JIr4FDv+oUF1vAwpr9
K4OosjtIbij8pFIxQxXIqBsfrvPNRaCweuAeWLfg6qqfAtYwtX/1l15rxQddIzLvbxFYJKcxgbGA
zwkLk/vr6y+7mRAlBRHbw7Du0Sly/n2l3gEInf5IbD4+Jp6kKwfg3+8ECfqn6j4Mx2xl/5ereNsk
oE9M0BfviBpFsYR6e8eUMMi9sV2fbNaIvMG+HDEzNZRb3ZL6EaBzkKMs9aIY4Wfsv7Ix7sYxFwNq
8npvWn0TIXGzSk5dnzxPTqsq/BUhJcJcmm1khp6kqGRxxvTBgySkUDyLBYDAJj3iYvAYew11OAUS
P1x9AEAW0RCKY+qG+EqYsHi39Z+ne+ezP4VQpjOmreoCS81O9pHtnag8vTkeY/j8RmGGm/geJd92
8VqIr4nfHs8WFXUlUPghjLgE+YMdnfjkHPEx63INYMl+LjPE51Fe3sXK7iciEqEJSS/kc82VY9GR
VD5Uy0XCZnnaM2ZBst4FBB25UAa3xHkrzW8EkPb8/zJ632cKyxg0Pe0oCuJc4kIyroHuyEZVKrd5
GGyD6aqD+ih8EIfVnfDL+1eiZC3E+t0CDhMylxj5JRVTkhjsg5x9irb5VFYmNf+ADfg6/4sWdS0s
OEgv7sciPWZwiO1lGKK44SHwzDAuV7gQcxqUopqJmMsKLfYsVq5DQseE7z8AOKlK8/QpRlkvH/mz
NNF1JIPIVlTJ/Csl3kZLJ3P6ThF5qLhXqnjaxP7naiY8xLO79lfSRRz6VOwjb5A27+iXKBNmEpR5
ZdQ0xTjwFQuNssaUYMi8d7wJiHnXekMYEfWWC4vGh9pKGWsKWYw0f0wFvobey/4gm9VnealhI2uB
jSw+nM/tp4Moenap6xqT0YCl+dvcalcdgbHSSAa4TM/wKyzKKnITnIDeO+ZggFV3uh2Og3n0kLIS
aKidQmVLturbiQf7DZWrAMrMw/qFVib6B2v+4VZgouOTWRORUNl5D47nt+d3pBZ4RGWwGKS2XPPN
bS+YpeuYXSqpPyUC72wYg9mwpf+t4oTFKvhv5PI4NX4vfdSdkDKgB2IBAaKC6GmgiyAFn2XnVQj/
T//g8oBARBzTddP03a3BoMEUzQAU3enEv/PRFGWn9EEN17WjOSETfgegrKU/pB+80mWZAWXGvFUP
WzfvebvBg2W2GEMz98KBgqjkjAE41cmmjUx8U/RtHsuc5wRem6/ePuHmbYq5JNyTZ4kUc4kFMcDB
DGkdeErVtM4M4bSrlJYDo9WqsVuVDdpPh7pZKhdnN267/0/T2aoe/zGCPa76qki9gYJM8o0wbmRb
ktIda7N3CZ9fN/A9/WrPkXCDe2Os0Lcvkl1W5XEcOryXtdq4R7dTVpPwEiLxs02SKZZZ8MdSmFI6
InFq+N/S337eD0lox5d26hhcIULaIGStbqwymnvTT2X5AODo6OFoX/7s4Sxkg7BaRr5DYj+EJcCu
XsOR5bCXxeSWta/etBWlo/KL6sqzQ8rNvPoKuOL1mWj6tX5/ouLCgOSpBX3keGz9fyoJtIX/K3dc
tKe8HRIMt26WUqqFGKP4rKj1e4DbuaIyZxKcXfL7LGjTJqZgapm8AFbbIlbp/V3D8WmoADmIur47
NU+W5E3wULoWU6A514Y8Xnz4n3tqTSx80fns2TRExfgc+W7B1+5Hb06e+UHlGS1yEQ3kB7opax9O
uOf+28YCzSj+htHqI+nmRPbbey8/MZu7WIPPLzM5VfIlIj06UlBtZZaMM+k1ppys9xLybioEK43a
LSTI2pOHAjSQgP+SK8ucdYNVNepzK5RvPNO4PaIWlXI4jHXgMCu4w3Xp4F8i5PRm9aLokZKyI5n+
EcWsrc4ubTLpzYlMZ21F8Swp/wPQ8DdZOLAfT1TogLcQmfVCwLmrDInUTRrltcNTkahS6niSZGIi
8IB9qjz/DjuG2uZnhzyxQMuZJsQq0uO9MERLC9NEnouYJPaDUsTrCHhqea/wnG/OrXKjvvIE23jr
9xrrp4rAyAOA+k78AS81t2kDymksKNO2Ng+5dOpIEmjzlEVYsvtk0Wsm5ldOLCbKuK9V1SqbeywY
0v95ovXibKKu39KmjG2nxoTZXUDJyJuPxR/uC1D9uLL05/x/D69TbPClfHJ8k9x4IiwAI0RSHueT
hKsqsCR/mDygxbyUNVjDurLiEMooEp0X5XqRb3zbBqIW8IkqelvbN8zB73nLxSYs1HPQ1pRseRF4
DYUOSqxseh6QGN+GQS0nP3FcKUHa4o1GrRotnv+fOJjZt35J9xcnusFU8frbIKvLkzRAiTdvIbyv
k9GJuCUTTbjEmAJBb6u0AFZoemQlhwlm4G74VroT7x7RnvX5jPhszoZ6FmzA33L4RroaFtrOyUSt
XJ2MLjUljHQi3Ek01P+6uhfjxLA+IT26fYYstqDogp30uycGsPI8m3sugT27xscRRWkVsooGK1t7
w2m06x3a35Za6Asj4XTb996MjjAMithsJtnqOa542bwBOF6utP/mnwdeqAchOviJOW7LsW7rLQRa
LGtAZjeb9/a+RF85WN/egbD1Y8U1ZJrMr4X16vFUnA9Hn6dq8OQOVt+4iHWrFc0oV42h3rViKhMv
7T8r0D/WJffYN5nnAYEaG49m5UF1Z7vFOcX8saoLg0d3F3oYuicC9bURz8lRTwv9ePFaOIbc/H5T
4DRBnItP1Mg8AD6JpGkISPLnyJZchwqr8XO+JiVvQovZsX8IsbLvTcMeaNmUI3czuDqJFBlrkh62
3D6KBU68Nueo0kgL78fwiNqX7jEtNCb+0HOJNajLf6NWcykUsy9zE9FDSDok0Lnkr9hyLoRUOOPR
packEXR3iaPOMqT8AWlxg66IpkcERMB3OVwlxoIfqYTTt71Cpffxi942BGSU/cBrUipZAZF/SCwt
7zp8kSKUaHcsRp5b5Rx/bKVQG+1hvg1b4xzTeA+Elwc24VApSmP1J9NYPFvKucO9PGgrtpAwHSnq
HWJKs3KaHf6EkKBbNdqgJbfK9QSJtjaobQ7QOs+MWmcU4lSCb1Zj9vLhI6m9HYfrEmqU9tw7bNZn
vG0N9pn+Q+egNOPu+UN8zmrzc24l3klsRTKjsv/8dtXhwxamqYxEA6/neYyCu0ZjwffjA9h29NpW
YGbjkqRbWYBxL6CJBO9HYRa1NKsOwNJXtDXo7f4OUJdeWc3AE1nQuQGtysc3/EH+HGWaKKB+pByx
CeNp2izccdFOOScK4fe578rG4lfPuobWG8EJMRbCUN92COoo/jXMVj+JCJbQxGpl5lsSkUtpqtf1
RyIfYvrv0OutIfp7TpH8dsqhjAo1/zXvAxY6aAoAjxAsDKqqv+vZ/b8aKdw8U9dB0YZlWFE4is/Q
jJHcHLBc522aJOKXW0iOs6zKnFcihbWQh77L0lVaSBf/XCtdZcFKTQjhtCbDKl9EA12MEt9LM8W+
tDeyUmIzI5oyxXamRt44yw7jMvn7+fPGtvDwV53oulptGPRYS+AlLb819/aKy4+9db/GE4Vyc8V4
jsDYoxYNbXYgJmWnpJEmjEpOygDjsxeU3geOyvMPPn2M5PviGLG57h3BDKYkSl56UvsnFvGiMqEC
/mspvuO4wUkxKpbvGluDvjJCQ9rw0IjU5g4+GH9AjrRc5HfYdjR9OmD1EHOjo8CrAW5Fff4cClKV
O9oDVp1UF6GZrjZ+YVbjEgwNWYs564vvNr9We1o36qs2GmRdCyJpLoiLRJKPINgoxggZ8FtGbJWW
7H+8WCFi4GVQi2RjJRaFMzAzgYRzqhwf5BTxFa25nrxDDUxg3PheR7gFO/EztRRcVODFjzce+V5d
A82lAbE3Ugm2fwyVXSt4uDk6qSW3SekUZD7W1qXa0FvIxBBWLRwYhiU/TAZ9JoYcsRd5gObn0eUF
qT43sGyiBu0Mk2P6HYf4/Hx8E9NvWIBkTEGuNPfCXPzMCcyaMM8VRzlbJ8mDKn8fyNStTi+AQFjy
DoTP+vRWOgAWIv3a/lk5S37pRglN04sHzv/ZMdUJq7QRthPwsxAXXgVfeG8lkV4xsYGdZXSgNrYA
x+j+zJUEUmlh3D3VfvjHT5HuM7qSGAk0nHAOUjduODYw2JoQO4wHabRLCa/+fCT43ZV85VZ2Exmg
j5oCBgEhR1t74Xewhm3D6bg8xe21LNIMugw2mcnioQ0v5wLPMuMEY9Y1sEf+aKzhb2EmrhxenEHf
xYkdcE9fZHd8upB44xpQINHaULVXF2VlosEcw7Ly26KASvqgRJYObsSpjNirD8Ot+52JUJsr3pDn
UJEs/l1c/y8PMSPyszr5haRzcvnZJxCVxAxPYY75ya56+1Qzmcj/vAPu6PMb4zSVMNt6Ol1siJxc
2Cmx992upK7cMeTCJcWkqQqws+pQKYpQPh0bstvn+ahEXPYcMik4OZTNQnuqW1ZoUHpsTzJ78MPn
t6DlBcHFIk8KArzFmIhHGw6DtsiweP91YcK45g3m9E/N0EiGAkpaAkPGjMF24w2gjVB1+CWi07i1
Zn4cCvuuPNUS4ZiYg3E8k9lIYThAcXrAvDXq74bS5d9a1H0qmcRcHiNnBz8rKkhTDz+qui1eyVUd
8bVcg65YDvBVBm5MquMeb3stDmUmIpZFfJcwEYDK3XHzEm8YmufYcTZf8nOxR0TCa5aGezkcJD20
fSJHK9RmuKA+wbffiYWnwxgC8Ny9JeUkj+SzgYM+wVf6x+0yfjrrAwRCT/cdpxR6YaLbz/yPaMqB
SwiVMj4A7IykCwdLbCATC8SdLOyxz92zgBS4JpGfEZ4PPGwtDTBr/kwwiGZPEgBc4NpIy5eeMuXQ
+HdY+owOckQBEqCKMn1fwhqceTZZj5lnQ6xulI9+of/zBl/TVQJ+UFv9EOdTEF4+pDn5bcIiqwXZ
8g3ErImIZUMtW2AqaK5AFEW9+5/44ofHvrbvWbhIrmFpsjOGidP1cLhh7KIQ00TShPOSLxDlpYP9
KMeFpIZCNSnwWIjohSUQcdHZbniFmzNN1+jzgmJheZtjbdr+5WIXZbgF6vdenKtuvrjIHbamoQTn
294eHvYMHU/CP7Cqg/ykWY9zvcN2nNCM6Di8oeKb5N7r300Mc1Cjnf0j7PdaNDl2jErGgm6ocR6S
2CrNdLFqiPJ1spn2y372xd/UxJQOeMGcBWKFZznJLuJ8xeypGDoszwQbCusqKqksUgRsioSCaYew
QvmGXYaSqOTmRZ+ODhGzpCqykJ7A1mfSL05hFuJwusrnCdTbtDjuY0sZz3enHyd7p6uTZLRbSp7A
rfg+3mbccn7oq+7O77JedaGdJMYgU6Q6yJLBWknme0R0l1nJ2+fvNtRLMW4wkOYzNvHnReffG2j1
Z4SSELvtGVby+EipksAM2g9clAQsnuxwgCaiFILtJvQrrMQfCrNipEWupRG3+d2X2J1YS0CE+Tej
UeHCh3UfOYO1P9gW4ZG3v103K29eTy3m/A4ZIFLFFdgM2du84Uw87OY1wnc6H1se/XbTA544uzD1
XHrUIxy7a4GmLTzs138a2RyMIq8n/P77WvJZ1QZlzojE/dCZ42m7VKTnCMCWPszeFdTIyaEH7/wn
Y1z5x51rgcQonROv2jNcmvtRYWIh9b0VdJWy7SyEpQtpIydX6UNDJfc2NsmNryja//Db4NhRvqRO
bheMlj9Hs4Ugpg758Vj6tlJEooYweoIkal73HUR9KnJLYIXNrM7eL6S4ZXD75mrQSmQLSKb1bmMZ
Jd5TQJTj2+auWwPXbBPV6P7JiYlTJmO+DMBJKGVWATJTXM2Yri+l0I3CPNGPAE7XDEJco2R1d8Z0
laNIjUt+EdKBGTIkkOKSU1toioO6m2ywm9BQXfw8QdSXVpQyasOACz61KIHoE0d2g56BTGLwV9yd
U2kBmmkm11uPMZKMW7OPLQ/ET55GPvNXbCVOjvtZED5YtmMNNdOEvYn1Z0C6UKlbEKNfKdnERc0N
IMIxd8ugpNbQT6lPX/Zbf4vAA2yCfh4sL5h+lIMsFHiGiiyP9Oe24CPI8HdSf33uTIfn/4Q0KyGq
tqJWsmEvRReXhUCPppJIoH9WIWjoGw/OPjZ0QwpXV7uWQzqYesio4XMT8opMfElgYSNaYGsuQ4PR
86Zz4ZhMRyemf52GHFyaxVA9Bapy+ZZJxWvXkMLBDEnZ4VnbAZyQ3uPOCxZyMaVvyE6OZZ5tgD1R
PqS+qba0sCNf/iqHR60YU949CJnaZhmLoc3qAOoGoRE3sieK0B4jdWbzqwa5WtINRR3f+aKdKZh3
MWRxnzoPTzJLkYduvdbwWhJzxhEvlusOtVJMebHsLgVSR/B+bK1bCZmDKngmOnBowBwH60pSWR2f
JJuqP+tU/FJf3CkUW0Olsv9DzvUjcDfsCbGRv/rL2kgB/2iU5iMMxr4Pafe5cvgREyZPdXhNOSWi
75Cs+cVE4V8kpxBd+eMYLU6MkDByGRa8rlLD+isZwuocuXJcB6HtQY5uZSmxCfyVsD2o7a0Ut5xt
FS+nBp2oCMSfvk+O2snx2W59WjEukfTupf0csJg5t40H/zcHgAvQlqSOfWfVwBa8iomjem+0bWuH
1D9aQPrI3nTMkPDEyIL1TtVp292WruKhyVKyIME3fQT0rUuD2ClyO2JN6IYAsebtB2nSmaRNTZOb
ERwl4eybeq37IJ2G6l4eujk+9xgwbVgtXsSBmvE/GPoEwJC1dFcHKvivpv3yKQSsHNFz3yi1cLdc
Vh2fnRtZ2dCWm15XUwNdC8FZTkAvQc0K7yLb39rK00mpizMLXIkJqJjMfCHxoY3LQK32WPf2PFdW
EhW5vYuIylZHc0TgWOo5b3M85LI7VRz272RxyVCXbs8B28auiQYIevwWrN4xpt52/eOcXEiYNfNF
SXAP1IrgqJW9bb8ndtBSJNoqXAEwmqRb/RcSRWbnQCVR7WtMAvMvyS1MjcvtjYxZIgwxlkupaMVX
yaIyFRUI4tNIghQqAzL0r2ollnXIqyKMfXLa0TzszYGk7FGqpY1L3dZmO6CQdzrrvSzgpH6wYejg
JY6Bzp7ooFo7U7DPK/chfbG+u1x3ql5AlO/S5x4pAglXVSTpbME9BNDGIYf6TatAAjKSJu7zX0Y/
yseeEgSiOSXKJB3d4A2OiSuuIPbTPe+i/3m7zBU/Hi+vnAYI6SvldrFPzdPNwb3BuSOUx9tAUoF3
dFPaCeFanGwvpZc33SNa6s9bInDBjrkAxPWlnsBI9MuK90IGBPGrgBVLVGrigmLPFZ2yycmbTok1
w8Q9HItlvpc0ECS3GBBn65BQDyQ/1C5UfMQ7ZZHS8+bdIJpgREGa9GrSw5UtNg7JT4qAiCvTNQoI
fGahDcpMGTtklFn8FCvxGl3WMH1IfAYPQFkgKYy2GKT2J0jnh4Ubte31HFMBevpZPYrN5sI1kwIx
2Ifj3mo5J7BA8Bc3SqsGnwkWVKqMSOFoOFAXVMmt+SGegKzKvnRW1WuU6odcv77+O5va2AXvzw1n
rZP2D80JftYiOh24wUSuT9v9smKO+LtStWZomPROpxaZnU7IXy61HaqxdgKXdxdyHnbxw0fQZgh2
0naQBwr80W5IRvpbntslB3E9s2TRPCKAFQApaN0OwpBQ62ycMQyQ31IrGobB2yoo4w2mfaPlyYWe
MEZ5O3JcAC+1eP5Fi/IjpauA6lNIdaWOmkF73hnYOLbBMjAPKRyEMilfCSIwN6z3dx+e5e3qtjYm
kW1EXhzkKLf0N5WOEWnNLx+o5Xq/xdpQOFEZmTvIUBrGlO4t7SYKqpMxWGqPLKYk53igo/QERoQq
XtOJYfghpe2mq6OnD6y1gbY1MVHrc4m67JKjCa/WHPvHqpP4wpUeGWQBO/BYBCYR9lypHidxx7zr
bGnN+dGpYphSIgZXIkiGQ3g0rWM8ngSXItVxcbBrekJpfmDQbJFqZx7SvwMrDrRqF8ifTSoQyNz5
q3rUxjUdXqNrpYaOXyuRIg4At+KaHF5tWqQH7fVnkyIPp8P0QscUI/Bjl7qIGlp/bKl2KtDtXEZc
KGeKoFvkudAnVf2NTpvrUifJ4ahg/yUxWBA6I0X4jDkIXr/yIV3+liWD/EUHfFfbHo3WkGcpzmlS
MduX4BN+Q6brRmyst7v2grJDfEuj1HOI/Ns43WVgYnW5ZDrEMYi/qRlj260SE0EfylmbPpmwbA6z
FhWNa2zfAk7yyErFGKUB4DoLpwsdk7TPfUBt4nvfBov4vd75amBJbw518FFWiEikMsium0oBVdGt
dc2xT88lIQQl8V3p//K3QC9aL0Y2O/2hrpvy27JGbUcF8fJ2M7XQhyDWOLj+LdyNNkwS7FRYuQ9P
Xh9in3Qsti3h5/BKRhE7q3dK4MHeRCpK+wcbrirXeIxa5oTFavIaehYkj8LjFhoQgeVncz9ED9C+
uKaNpGeHWFX7XzxMO0YdeCGHcAPb8PsCxc60bbgk82AIEwOhB1jzD1xsKGqzITN8IBZF2Gj250sS
vXy2sfIObQGed7YOGGu2iPQ4CqVcR3cv5ngxdaK5Fz4NCGnFyl74tq7AyFbzMmSmf/gw2x7g4eg7
rfOeH5ZEarnWmP4NPvZLur0nGnV5Nvyxr28D+KQn1ZJ4XH1sfVZqwEaFPZupK/+h4V3bQX2fCUVC
t+ijzmegpfxyV6oL5nOg4pJAeVLyTZULK7Rc01TLh3GVg/S6rb4wf6mzdQd02ibAUwa9p3dZ8sX9
7qW4fw4mCGnqfOgg4pimPRBxUt3EhXT1UBaBol6LHbH2DzWhJqHmN1yaeCsNFr0A3o55kxOM/YXz
vuF+FAhsWMCo3LeEjV6MgEtpdipkH8hVQsbBTcaniloqOqKskykNL4sD5OJQqDUMiN/yHyYZLOSZ
xSpYCKlf84nB+4vKh83kcY97imVxOkuih/1Jf8/LrNXx/23SmjNKUxUgVa0jwMw5K0b1NKpMBuaq
AA2aaJ7MIkyMEZp36nkhbqfeR23g9wifqakmYE+shGnFUKSmxMs7Bh/Y/08BTqmScWwlIoYy8FGQ
6UUss8yBXmRwK88u7EUZ++QPyY5cLnuj1Y2WIY1VhcY8AJDeguwfljOFK6mrMVjjnnapgS4ArM2g
fdz76BQS83ghfq5jrMkJXzqHnpYfmCryyjK7QPYzrYDN8VG12s1SQsxyzBm0gNH63hLrov46QmBL
InDp1FyRmPyihKftzTwZqogTcTOUp7mGNq8d/yd2SRZUyyrzSvQgbRKUApySRRseSrOavNJB4NfN
1nOFbqegWwcFn8lGl9FW8kcaA1UwNHPtOIKdMWTD1d1hVKDu098Rq4tD0FeU33Z2xduFz4H6PKvx
8h/0EeA67QzBmKaxoDiDU8+RCoQCVt0ISAcWO/PG0dWYTauvX+vzm2aD5GDb9WcOzUlbrwPNy2UA
YkIUejpASsZe15qJOFhyG3sFd7VVs+8rpSoU2KyVwX+5YuT80EZsPDNI3SDgK9hvUy0qgDHTjVXA
s4QzGv0J9nJW+TmlDO6qxkR7VL1UyBZ8cpGRCiINdYZsREGvx799IbRnhuBu6zhgdQj4zrZdT6HI
jx+hDsUvxzFpyptkUf9gARZuhGX6XchaxKS3ZS/jvr4pBe1e7fg+aEwOs/PLP6lJ2EbmyrFASF0j
G6wof2Z8h0yRrT8DMGJkuRdrGFAxHlTmKydFEP+kVaxGsICuHGv3hnUOQEKJX79UIm5l/j4X+f5y
mfHA+ymzfBqAz+8nJXPUMSLN56tnx6Vlo5PKLAt0S4oquUhfo1AbuR+L0036Bhdhvd+L+FeS6xPH
Avgt2y3/BNqoX37QUcEQzishIEviD6mLrfIedmpO6LDO/9Z022iQe1SXoee1aRVk6cRGTH9H9WHe
O/ZGm5iwrWm5bRVDJFX2Xr654RbBVfc68MahBWqlbTUF/l9/ldUN11GpObbWY6jD77Tvv2FRc4gH
gFV1SHw+RlcJgPatZ7W7JbEeUctgu8Kx5t2/rtyOKUIqR5zQvtCq6n444w6cQmryXlTm5Kip/Hy/
9lzIFwyQdGdLJ/qcOpdg0tm9s6yrhUaJU4jfbCl3Zbej3e6UoW9g6LYrPLdHshwYSfHyTY1AwHbw
mSpWe8dDYd7RQ3Fxq8Oebm8bappaAj14CmfsZ0+qKz0HjZCPDVOTg/GBIy/6n+e4b2YavYp5yzFE
F7gsjejPvbXaUpBEKXZve+c7KPPyQmVZWzbewAeVlmCv3gXZNGK4WPlxnI8L6fN5XhMH44Mnstrf
HBxleMRMYDR0a2rN4N7DMITdx/GgmX2SZ7MjTXCEPkH9UEnZmNOboPKylUIpfGrnWfLABEh6QfLX
MUNCnFfcJHus4jVJkymJ/gpah/dAHiXRWS90QYs8CZEY9GqQuyUxGXydQiCWI+acQwmcuUVTGeTT
SR0zF5Pp4mrjef/xD0ZrOeZzPZ+7R7ValJfYmE6dmZM7eI8CAHilDTbpBxWf7HM+OJ7b4dYt99Uj
muWhG949+zj/QaT9MidRQV1ps1L29qoZ4VZHb+WxyqnMy7IBC3CZgM9RFcnJdpFPeVzYqpJAblLc
V424T61NkQ9mUqTdlrkefnxLxID6iXo1/x9iXq3bQWYE1f0fsZbyXuMOV7ZDrHPxjWd9KLYhFVh6
CVW5GuzXhOhnlHOwrNa8M3CCbmdbJmAvWsjkN9ZOh6kymGBS3kqehmhT4IlfqpeVIVJY23JPvkFO
d1qVYYfQ5ZB2NAyj95JV42Q2wjx8SCC5G0wGdjlP4Fw6VrP6mskwNvguik8N2H1aMNfkOJQSn+2I
TTHB6dhHR9Kw6Qqs8y9oVSUAqKY5fYxcWYGuu5fj9uHY9shwS0piwkd2Fz1q45T6LypemVBf+D3D
fi5pR6HMQ6G0PahwutOMWV8pjXGAaqw9J2ok3ArCNnJ5X5JndPiPFumzlsqUnU2cOh5qyDenPQQ4
IkhA/EzmUFSa8MwO/5Llrj7kTkOfydmaM9aG2z4lofX78UcmZ4W6a00+wp+/WNF/56Z/qcJfOt/c
9pEw44cfiBKLcRUp70eq9f2XwLpkTbJzUxR/WxMZaS8H/xX4Ug57Bp8Aw8c7KZfdfEQxKkx6I7Ig
xQF/fzXDV9xDlaYacSd5tZTJ0JJtr++c+/j4HIG76+j6w1NojYOSxhORfiq63GNlwGuMTqAA4eC7
IIshTVUNC5PDQriByH3NAdBIidWekMNPoHKbNFfy1dAlZuDpiWSEbG16ieXZNuVJLPrWZtTja5hS
xDClS4aIiI+2T8Y0WNuOio2zXIHHGlO3LAemI8njCRBrtx/T9kBNW37eGbH80FZVaaad1YjCJpbw
ZnfdzzYxiM6rI1ycHUtTy/yNNPPFUSMlqhPp9n8KxokRNZ5nvLeJqdwBZm3fEmvWj9kjZsSprgNW
fI5IlUvE7ZSQZdzBU01B6sSY4cRUZEfCsmBiZajkNYSWIljBZaGJNiM7rnTluu4bx/1PZcFPStr/
U/tnu+N8IbMWn6X8s3uHYPoROP5gifuMRGhpggW5W5eVHCTfK47zBue3UYXHY7tInxrf8bFwhwR/
uwz1q5UKyXXDfAWECFR5h3kiFbw7bKlo3hNPiGK51SpHcAWrGlpNRyxuIoqa8dx0Fq4z2Akl+OvF
V8SoVaW9j29RksKfjbRii/XHHl0m3XeB1nBjlgjiASrhO8Y2z5CAp+/Bpur161+YjWv0uHHARd5Z
gFBSbYsMRJTNlOKoU5EGqayVIepZ4lZOkm6ussbS8e/A8JN3QoEDh95iH/lnjAK7NtLrqRJB6u4m
gN56Ef9FzWFFDWKsVL8pQmCAWoWdVk1XjssfSWvyvshOINIMc1ea5dvpc1HsJIZ0voHKH/bjr0GF
flDq0rtfZA1L1AY3ukNptFN0bXFtAegxcvsr7z/XRKctz9dSIevwWYI7WdL4oJkUL5HRTXTVR4EL
yXk4c35JWBWUpkBPgmkHdbckzQtdsXK3lZxGSS/+JXJMv3juvu5zprrwrJIFrDd9JqgARgLSHKFy
hkkcn02O4H6HaOPCIevUK3uom/rvVC2a/VNLcEMW8VnXZUjJ/Kz/MIi9WKuCoJioKuNiDCo9kBF5
cKVjGW8DCLPudeUBVng9ZgtMxfygK8rCJqk1pm5J6LKPB3ElO7iFuMZu0hUeb35noQ6HqdONCnlX
5a5SFVT64njcjuhDhhFJZKGQ1dGtQ99aMViyRKnbho0WrDgZrraVeeS75i768gfe8V50VyUaumpu
ImSOZRA8KtnycIqN1sHQBZPTTdHIvZbGQzmdhz+XzpG0DfqMQ7rhsc5ONv6yVIVzHUpVKG/iR/+W
V7R91Om+wDZm9tlWgk8StLS8enEOcyUqJITXISnDpWsKSjJzAsdllu/TKb8yZzs+71hXCJ4XaDTD
7YpOUMGiAdmXPM1L1Wa3WlmpgYN+Yy6XsCT/+/e6Sp6CneIUWWuFyAfd9SZGFNqE7JPwlW93pNof
BK0REetPE0Z+xxesUxXTaOlIQ9MFH8hWakqB5PCtPFXSwFzvjlRGvwzJTy9JITt8LqNMHEU7j1hk
/2hdBv+LYJyfjm1lXdGuuARPxcMRh8Sr479rTUzByhJ2vRvy20+s/l41iV+hLXYw159/z7aHxmGk
u76GpReC2jxqlXqceUhr9bfFQNEK2A0VZLGJDddmnulMz/inX1oW9G8A1Da0JUl+nveVZHMPLy9M
pTAlhV/85FXMOUAAr+7vAO4mFvp86ye1TRAkodT6Ygm5QtHIwBmD9LrWmE+jQKLUQJPUk+Snqm/L
YEUCCpWgYnqLx+bIg9jFAxuV7dwtiqXzeoLjkjye7HEpRBia9eGR1OTJ+CloOCj/Wppo4sAcxgoW
X/aFjTGR0oinm+uLCHJiwF4Fi1ZqH+ubT8DEewNuPbV7TE+uG8nYwoN1y6GNmss+G2LAOUt9/BAd
6e5ScynQqWAky3SJXCNpxaNlO2+O2KxNA1yo3TgWHIn8mQhJL9w+hOR7oK99m8N9cO2d9OlikK2B
gRGsWhehudoZ7IwJxj589n2ibUS3rriDQ8LODflDZk/vOBdile7EVe4Wmfq9V2bEJ2eOKbzEk4wE
BE5hoabbPdSxrLEuCeyEYGUG9JdDjISkymdVGqOP1JZpugVAF5sdN7RsLfMBPbDXvCPzGWda1wfM
j3r+0qLRcYF5Ek4P7nDl7EEWk6Z3yx5h2MtSmVD/VoBZYVw37rSdE08W65EUUpScqbiTxNkfVKly
stuo7Kd9D1MEjnVezV8NIWYl4ftCXrb4arXvshxw1yaR5VBN1dKKE56Q/+fVbKDNRZOG3Ta+nIrv
Y1WTUm3s/leGoOsRY5cxEj9Nk2j3h+FvUFPaqYGpuTAzBwVtoQbwqtiwqJFFbASQ+TzhG56J/Qur
tNTaOiu/OZ3qECWzGe00ASiu4ySl0L43LBBmnr4Ku8w7n+njplqsGwhggT0A5oHYl1lShAoAkd9G
1kMostMeazdM2dg+gj1vKZgWByIF8S5PB31U8XZ9zFroWBsMJrRWjYqvdncw/YhIc2WLo7adYFtt
Q+RUiSPzq8SZ+NFfPJWTT6kkCToUcFuhW/arFKcn6TZynjNYLUW5bXnyRUuXD+4PupF3Y1vuUYqa
vNfSwJtbKavnlpJdKUCl/cdZaNBWzFmc2PSXKKLTMz85UtxeRb5IRJFD4TFacEHjiGKXkTeONla9
HreyfCFyPTJcvH30c25fmVD+29rZgwFl3g/MIJ14duoxhnlGvAs8Bs8+pkih2wxZmcTN17ceuFyE
L+csPZsTuexE+R88T67zGwNvNpSzykJJXh691pPu8oLZ8sgodfoKTjX/e4XJJWOazc9bLYD3A1vB
ysgGCf+c82lRli9Yr3vC5U4MQhZwiffBwkuRx5rBp0+1VRWgWxoMcpVUXED18ZPE/O6VrIxh7EUx
KwdwJQTUMbJfg+P4eOmiTqe8aREJMUcCR0BtZ5DEbOznO+5cIhip7wWaJVjQ8ZEZdF8htbXz1gJB
g2tvK7p+wo7HE9vp0pneiL4ArNw8+2bXl184x8bAwSVTEfPwaobgewQhYpn/voCiVeN5v0AqFOj+
MDx7H51/SqeF6L+m80CqEoL9kH5Tv2HFu4TyIoLEaCpq1uy3i3jD8rsrZmXkGufii2w3CGfhU53c
By62igX0HgUDcXjdh+z65gqmuvanD/xfiEZxpmoWlhRDIFo3xZheC3J4BGCj3TSg3QNR2/VTjBPG
864f8fgNtc4iiy5n9Sx8tl+yJuhL/L6MgrCcZMHT08vq4VKO8WW6LRvFMqgmqTCoHeyHiJBWuDgj
yqIXgiP8actj9iaKi9lsdW+wdvJZmMUX0y+7apaGQMlaMNclv38MKdb4AwHh4B+FHKbQUB5du2YO
2BTCRivVwg6mnVvT1CLYF81RVcOWQxf7sxil3UERWe/xN0AqyJaf4cY0k4483IUpq5RVXnJnbZgO
aqJkcyVFPAmbDuVkotH4voLZ6G8gJWII1LsbKP4/Wk5xlV+PiJYscZxYFAvU4hsSS0sKloshvJ47
O12PA5fyIiH55GGRz+IWgX1zCayxvk9qqDD1QOYEdDifDJY2M5QiavncpnH/V4e6AxIUGLs7Dxgl
0h2dLSsRuyW5Ttq1+0BV+2sORVphwPfdn0XQcflO2B1wWQUaDxa72UF8iihZy9NX1DOjgbvCy1T1
sAUUVUsICQWPGXguFrqQ1tCN8A6wLfnMyM+s2C6ItOdRuQT9hHXIaD5fCu0QyiiGvb9OiGrEzC4F
EPe7K2niN8pkMWi2iJ+yGE7YSIMpFoDjV+4jbVaSZpIPMtX/Hy2WEbv9hQ22zK7PstbwumZyiMOU
LMbKnRxVWD79ThxNTU3bbqpQ5MqJH7LdBIwZArg4ndaeFLcwdGhYUk2/0T3LPWnoxG4zxmju5UVs
HvSELFKyg7CXzJkN4pc9JV4suaJ2xXeQi0n3NnMGA2VSqHLm+R7+jFPJMtOjJSHwNb2eWpCwqAGO
2J44mkKL5W0fYimFlphLaXH07fZngMsgBzuIBcqajWI2YtnpP0ap2qdb0vd8Nq+reQsxgaJtgY3T
Rhs/caFCCXmL2euJM3u0bjgkygRtcv4qE8NP8k5alcRMWjnGqDfN1xfev9nqP9dtUU3K7H/NhSNE
h835OJjh/VyzHQNX2ilndCkLmeRSCF/V1A2f4cwUm6AkQnilJDciv5pCLahXJaQhNT9djXYFaMos
Lqfy+RUiSSWS4uqJt1ChD3jjb0dYA6mrN/kooW/L8rpFJuxWjmViv13d11/i38GK0AE7/JXqkI9w
tFTBA+5u+UFfiASBLMSnfVoH/oSrYEycY7W159L+MOxHF9U8t66dUK1b8UHK6ED2kexfSQ475BGp
+1a9LsSvxNg0rJymWn7BEWxk8izLdU4Gu8IlmeueodNLvXOc4eU0oL5Bq5U5aUdcCjCygLYERNTF
IWjS5hqNKAXtCC57Z3yOqppO8lBfdUdxM7LeS2DbLrx4E9ODmKRJbyBlHy4qaNku6EmjUZlXeAGz
N6s7w0zUqUXjqPhv15fB2hNySAeJ+vEvDs6Y6zWLFGarTEysHBCih4SVf2tLAyw8L0zX0XHFP6ar
pRN9Je08xRjloA2YORqepAO2Mx5igZsYrE3b4nAyasyw1vc2t8LDYMJlWW7f611P/HCdg0Rvb9MV
/HKA5L27LMEwjH86gNGxyR/LKQ5AkMl8ijldlFgQafWBLyfXMRz3KZbvUDh6pDgnms+LZWrqRgKG
cXdD7fULpdBUSRKCyU3bVowlLweGih0DELTKEE1NO5b7StgJZgD+MBnkq6eHJzp6+yA0p3NvalfY
UfNyDJRsF0tAwA/hQlPonb/hzYW7I1Amq33fsukzoYcE3fWDjlQdEa96bObH8N4kiTET+YWHPNiU
HuIz53EyJXAjjJh9rE8rFohYqmEtz3UPoYDWaq8v3jfzLDAPIv2YeQ2lwvQCU58a3cF1fhBWBNTM
fUL0vUq0QCsTgozCetJOP784JH2YUt+j85fTJTTo4VFIbClBHJDui8GT3GxnkxRt297C3xvQv3L/
4Ntis2P/Z/9479mx0Iv+WnifQLZmF9QQk/8iNnS6/69Ms7I8Pf5EGYFwVamUS/MPd67DQRxJq5h7
XlPnwP1e8/Yh32DjhW5Nu9XrdTu8AvW4U2qWvidZGz7r6MGT+lPMUIicLfVBARJlLXdmrguY9V2/
HsqJHecDj25Yk3vDGykvKsgbYliHGW0NK8wNKqp/u/r8pTzziHVPh67Z0+3wdGMGinQgSZcPuIO7
sqrS3ScWassnvMpzc9cCoNx1Bvt4kFTsa5vepJAF58nx8u+mAoG9P3RvioifEsHm+LKB0s90dKB4
iNoWJd8NjhWsIRAmmmGA9t9Gl55QyIXvJuJHNRb6UR/YZDScPr3AZErIh/apKU+qNlSeta8PABwS
5YrQ0T5pWTvdTwLjDSAvCA2kPo8el0+Nw9lwis45TG7GcwcD6KaIo0XgTwRjyuIj0iQ+XL8Mc2qq
WKKTEXmzIoAePERxRKoEf22qBXa/+uC6OMkEFP5hZJRV8ov+qCKdajP4jmMARrPgT+JzguhoLpTY
mHxJFsUssrepBpFP+lWLofF+8QlQIl5z2dx3Rk1s8/92crQf5Dui1YsvrrB/R9hqEFt/rznLcO5N
xRmL/vCZ86paDUItytRtPJv0fH/twi+Y5XXSVolNQ6aNJxr1J8VGJKLMPnpj+T1jShzQVO+fCL7x
UbDjoWafC9+s+ZStVz8B7VV5x1ZImvxoGhaBAVQw1NoqXeekfs9Jj7g+XvhwuARQW8XBv4oH9rpj
ALEXKfdJi2AKnXzM1gBOGC8mZ7m+EBf4QsYqHXET6F4Hi0mYJS0zJTEPKzSDCnKnwqOGwCaMS+KL
aLmeaR3XzioHVammaDhwqLigManX8X5XGDURfe0Go/h7K8okixZ3/3Vk+WM64rMIZ12UvmLDZlII
qyRi1+r846bNIUFQRn91Sy/ND7pbSpqi14fJkJwtWOk8SW98OYcUhlEJ7/HmmK5bW2QsEnIDNynH
uOHVcsUjkiKHsdDy/p5ZFUM2af0KyeXMVNpG2VbBDmCZweUDFLqbDzP8lNkERMOC5trXx/YVCAM5
rvpZAFrDbvrvMLd1lqpmTwEugE0uDnM1fBT0nTYqAdtgmAjVR+LDpju1rnj68hP9GjGtw3r3s1dp
8tkFW+/3OuuvmOiCeXZpgQfMdpqPjt9jjlR/ibqRq8Zij3rflHcXYrtMFQo5QM3hxSQYoC4VtdlK
gaHOMLY1AxSS/91wO6vjcOfhQuIpHbwbTio6fglDwVm5A2QWfgkqf6oWX0S76wH3SnhwsRcRbotO
6WUSIlgQds+cIXM16lQfEAc2sH2B0k8HZMRVLMrnxbO/aWEUJWaczecpRQk9slDxa9e2U5TDz0jC
YmWPopT1SSESJKOC8wTu4AWch0XkUOVAFttnbizKPNaz03NNOaiVSWnEVNi4lwMqnT9cJSj9otp/
Bk1I1rmExukO4sdt9XZgoDmH1xDXGtSQ/84c0Gq0WZ0IyyH92jUMoU03nyCN6kbWx9dYkL9+VMmK
j66jQlzFRo+ontQrKIm5pYTfnf5KUlsIOr1f0QWoTnhNs638WA5d8sjAyvQ7UaEqRRUID8KyHv/a
YsPqmJ2qy48cqhxMUeWiQLVqtOvL8ff+fmGwSdOCg+yDOPXkg5GuVRhzA8WnEWr7nBdr4K9YNAdp
4YtiEMAD1L+HHqCKSC3Xui+3tgW3RM+OIztE+1HaY8Lz7Di9X53VfsSkSqcaRBPbqYw3l1VM8voa
h5tbUEJREYrZdzpffN6Y4lv4cNK1ZTE9zg3Yt3MeT0g0ec6pPUUBynxt6mbD5Xsa6c5eR1cDm7zH
XMANzEsIDe00Q5Rs8RvnGT5SUkiFQg+WvtAa8m/PW7wt6lC53ijSphshJcw/kqnuTd8klHdvIPxl
hClLvu8vRFANsb9+GdiZibxa6t0mCI5rLZN3hFcAj9fZYpFzQKBsZMDtDQ0vmRvcAh7zNWjk6r2K
oCkQcp35pwPeUdxRLXanyWqjW+V4vpQc8XpW1Zq1sBShqokyiHf9GWfb0dW/rVDMXb+/OUKsW5e7
rFmkIVEbqtmdlyfcd7vtIHrdgbu5jFWkaU0XyLPvX/+k3MnBzJrfzwIynY8NTOHAnBWqDfX0Qkkm
UwAFffvgGAUil/48z/iL9bYPXiQ4OLKzAJz/ebS61kA0rJaOtWBd5IoUCaQ4Hfv099Kg8mhwOnVO
qiGCG+TS2KgexU0N+8c8pYSexgePmPqdOlkxxnLfR8E8JZ3exFV3zt00XNMtJJMYknhMKdgWyJ/P
ofynRhLnOJBJIbhQuNzZxxffHSArhIDvTqcg1UMw81w1v9oFge3+BvgDymzoV5Elm8IGFq2npXcl
7u6s/wWEDxVENxTvL8wQOwpvIGj1IMv2HXgYxZBvBnCH60SXr+LCWjLVIy2LcElJjJHDKwMD5l+A
l4zfbUI9l2DDTQowLiEUzd2uWfqwY0eGhZd3fc9AR+vJW3Q5nXNnNWUYjmHNiWEJ7tx4VIa676Zk
nwQPB3RPwL8laJUPCFMaWmqvRaJqTXO+vWlWKwrCRJ6VYrlEi8mNXJMqpPvmkIwgEBdjEEY6RLG2
zli4shUsAUW1c8DsmspK8dKxjpyu2moxYLSvknuJemSp3Xbi3p1MbsrjY/6o7wDJYd1mhzwGgNE3
arYCbxrClvg1zeAjDphtwfZWIc/hax87D+udaB6AI9vsjjHrp3CQHSfvPudVazX+1f9gAi/8tSwE
c3uhG30sFB9NSudXNSG9KOSfzvbRfrenf0+GqN3anZn7m00ooesSMagNYQHhs4ScsDDKmYT5DsHE
lgwB8TcNWEJ8k8BSc0a4o/o0XvLFiMhHEnQxPDKGm3BQHAtSdNx7/OzWSOLH9kN0RqsGrtqKWyzC
OhjuKQjQlEi0UJp/1ygtcuFxO3Z+WagWTsQf0R9V5GFVlPISMjz/Xkd9NRZHjGvSi4m+VuhiCi0t
EEh7Sk/BuqNMZ4+VMsjitV8KZUpIhiRl/OdI9C5zok0t3FgKb3G7CzLco0Pmp9NzWiZ2TBKVJHOD
5G6hzh7Li/K4fGIcyzaTVQdNSCbfQC+X1vFhm7+7pCqxWLiUMeXLZWP1anY3kz0dueKog571ryg8
3BClGKyUPpqZlOaE9bxeqrzHeXTfoox5sWHncNMC3589msQPb1Rf7pmXrFJB6jMJL6n9EEZATVFf
MIp5yyk6g7Ifw88KmnUJi966EQW0p4r1HqX6K6jxBkuKUgHY4omOn4tBkiKjr3GA2cV+qlF+PPCH
0IjY5IMzBe6R12V1473vkcCjTd2ZRc109LEVmu6Y8aJp9l8QvLdFGqYYHbwO9JjVG7fGoAhn/D+w
sViRs6/qFw/sKgp/S7bEq9/kEe87XnJDro3rhq1cA3CmOnOMCfd7dY+vt1jA90eIdorqeMjbpGtM
DxHp1xGzFkjPZNTkpugLfJYhL2gnu3c/3F/7cmQg6ET6FFe/8OqKkN6YDKG1wloE904smOTe/RS0
17XxSro7YL34Ps0oOlJC8wvb3jiaecGxKcsIrlCuM/dORMAjbl2RASQl7dCQxGIEIUKstYcjH0z6
Fj57CVAfdRVccV53zoj3cd/xxcwMIZEKKr+oKWG7uv7RNGf/qN76HDb+PKCL+KlgbklKgxhIxMlO
eqawqPkK2XcQ8GwW/SqShc7MRvLmAfZlNqHZOaUZd/KHDyPdhg1EpYjNKr3kpBScrkMiWUPu5Qjd
ilEUFhkLkN35GmgFs3H7wQTvqTDs9+uvyvvz0F9pT7dt34Jrqo0OWWqXZkzvTB6xyXSTuvKNC2eT
lzYxCygDJ4BhZGkVU7SPeXNoiNL+8D13qyg7AYY+RThevL8W1FrFo2lBs7+41gKWq0x6246FzKkw
iEYxswTFzSOTIBh7A9gakBOVjbAHRsIOlpZKJDXf6eUuFamkKM86fkAUHM/lxc72RHnUZw/Ggnyj
ykElfixKsj1KfvuTm+LV/7CYpg4UBC6wtAEGHdCyClf46bPW3t2IKmlEb6bEWLWQwjcoIt6eSC3B
U8/QwZmsAn8KVR4XZuph5amJFRxy2qDW2/70O0lKzafQ+1BGcY/XfjsxS8Eh8+rCB7D8JtNdaBjq
woVKK4KE6AmcPhaDJtzMZZ5VTGMhpdIzNy4dZJSBB5DWjY4XbEJh8Q86h42vn968eoo9UHM8pFQi
UVZOxXsyIchsl5jJuqxlTuG7qW7Eb6GBcDPfyN9GVIdD2u/Btmy6vJD/XCQ45bTfdt14XJvYLwdL
w9qK1bkisyEiC+XROhbDtIZjhBhlpCXbxhKb+thktboIV3vSc4pNhxXFSy0Z2GV725W+hC/FNonp
fqeHdietKyCnTZ6QsPlUNhh1nogzfgbDYXnwY4ij76DSMBPU3mWUTEWuAxw0SDIeJVOAwgchVGGU
ShIr75GoIqq9x5hYeXgTzFraFxrxj+SHhpR58eOTrhqpXGIoG7khEP0A0Jzmy+92/g1ybutT5Jpq
6edt96SGWTEb7drY+zA4kPISWkbrcZLcJZvD4YCajGVggG/fQYKbiipzj2MUuT5byRPDuM59Fgcd
+lRZRPq39hSljy2e7ubPO1kkfz/I38N40+vEdnWK1SMORvhPcdi9cu6rPZGXDTdcWsh1z48/oqVe
c1XlzDJdEJXeea3N7x8kkEu8OuPMLvs6uwC02P/QUrZkscHZ430CgYjKgaADKXSv2FEzcIph5LYg
SFtHeDVMNOsxUC+lYQHe9NAg+636kZdH2lnG4o38R/CC7vJFqDW7sO6ZKKpByQttxM00biGgK7q1
Uvmma1mWLL7TaCykG+iQ0aUHpDn6znOjpWsnSTrZdRUXTL/NW5dQ6MmVba6mkVGSe7dJ6OgqGzzr
JBYOWogj5snKOLzLQZZKubgh5dk6rw1D0NhqL+BFgC4ejYjz/SHAaqjakIzuAbeARkPiWppHQv+W
iULvL/nuxsaQsBmQ6ykeXAci8dLfu0Uh1Re/7GYMTANMusH+LuvA7aLdbnYW8nOlTI7fpeBwOs2y
5Nlzk3psFtJLtmJXZCSeSQvqdMK6FexDunZoy3oTQ8ODEEwxyHEs2H52cCGQ1vyGUvWOEeV12iLH
ydzMmcaxsAtKA5sLpnd7Ef0+j9REpOl6Ltg14SltxibBiLXg2CbqgA01UUnko23K2Zb0cFjzhueb
k8qnOB1P0AK6EBBzB2HWrlX0gZ4W8LXcftp86fQV5iaJlel4pU3uU9zzUJhaLmIYPBWxGOxXWkjS
c2V25BTjuMzDUQvf2kBLDdmNIkaUHjOdxFRPgOfcQ4sbpsQoqvUB5fUGYnPx4mhT3P+IhaAhebZT
RUsheahnkP1Qej7wB9BNkrfm4GqRAYgxqIIeosqJhVhCdZVA4/Yc37m1O3IRwFFfR4D/GZcxWpuM
b6Q+RjGBUwqwFkd/BvGqZm0k3kIRlW6T5bv6MsnvxO1KGIHnDH1NMklGLpn+99PjvlP/ZMDzryGA
qupChJQ2iUYAZpCHw6qecHEpEy8hG2iLjmazl7LVQxpUyxEIuudyej4oI6Cx6rQNr6EL4cTYvujL
TfhD2kZPCtuvxJMOK0bc00OTckMUy1HdNMrOxkrbBXzMSrKYlPeRNAqNFbOORu/Niw7hRJAUE0FO
7hEU9sEeN+llicUPQ9f0MA3D1L9ugzVs8khrvlz0QLBOFbb/BI4JVX8ft0rHF6pBJQU8mjegmXQa
gSrETKPFv7UYBZenh57BOSZHcMiAgunI43Uvcmpo/v6EF/8I/0UYbNUuapQNYm1Y1kW/FqBaFrSH
tiGrgX175jHW1511YxuYvrDsbMUaiqYml9o9Kriyc/SUxxg3pP7n9Kt03E4j1NRbWngXK1WLOD1T
7lSO2BFicY23R2UINZZOratz8T4wdyoMB+Dter6qG8HBPy+aFG2di/pBS8C5tK0YeFppuL8HG79r
TCYvTCAJyJWdygCB0pxudAfPqdhwczQrM2BKC5oxfbCRQ4P3eLFf7SVD+fP7H8/UsK07af233IWQ
r4yd1NDqLpohwuubgqLeM+SbckyvYhrbnPJY0d9CH+I8AIlGTAEen6PLqG0moodpks3z8z6Sf/dq
3nTqKe4DfdoQ9YUeiOaC2fAmCG/AVD7vWJtnlbpvj+JV2KNtCFfIGGbxBVj2an0RaRUenvB2Nu1o
MVffb2oHp2I3rJB8fp6TcHvTCkxrDhJErXnIn6wUbSXj6rKnWPTq/PeZMPBZnMcR/ojpeQMCHPWJ
zAr8Hsv7mq+PX+j4m0lCHn3Ox71duOfXtDzpRYvPD55nYNGxLoIyEK9Q+mDORlnkPU13kGCEl/Un
DUH5eB/eRc+M6V+6fZKan4bViIiNKlQJkXQeg+gPSRrU7l97uiqruMShpImCWrtrCMfpun4roLI4
wdxbQytGW9KxbPCpy5X3waqqCAgtkk41uP3UJxF+2KdhD56VpPd2EPdUhB7MUZkGGo/eoAiHeTCe
fSFuxUyCEVZnwQzkapjst0kJPqANIJf2CC49grjBngSekwJ5EKYv58mzwMitsZDzkH7AaCK3l5eM
wv0O2KS9quY51WoyrHTjHI3Ugy1UpItDENipEY8vZrQ5QWG8RblGNNLeyjDMsWaykVW0j96EFWmW
rbhDFD8EwjXpybDhlH0VCNnuSrYnis0Jxb4JLTvDO7jQdlCBOh1gYGyYLkMpMu7bI65+PQFnt6nb
O4tAJeDPUwpfyjA9EDeMeEX+yQb+5czrvtcELz8qzXZnqEGVOeckdCL/TF10O5pdFVsunQm+5ojF
QY9Lu4L0ssFZHLBG4jeX2qhRgEsfr86K17noa/WMOiNCDw+WrUQdnagPRjm7itCUvAzHczTdItkP
FdEvcbJbkEr272MoM1b9OSd5AAJvVczENcdaxnxrw9+Os7My2vQxBhVWPQHu+N+79gxYl3nVFtPx
BgEiDAJg3RxBzPDlzrvC66M0Smc7Yk/UeA0TSdW6Yfnxy8/0gxukfXKgNjU+HOfPcTPnIHr+Ehie
om3BssZigL0fuie6ZkWos0laJolwdz/cZNZuPcmxRT8IM+yfRi4+3YEPQV5bAnSWXziup+MwGWFS
aVlz62Hn4iu6fPwO+3cuhHWyuPrHf0xcpQukGeGooG+gMLvnOLoWDGEiYQWFpXTIB+SzmfO8CBfL
S5G+roYZjvP3O5RRj6o7hgcQWq0ej5/Mcr7BLxUT4k44zOQbZFMCuePI5w74PrD+7wfFxKKJbzBj
zgpPSaLN0k2+ic201pGo+s89uCcqsy2sgtluGscF4rAX/jWe3MHM5PJM5PBfDzhRfBRrd8fmLpw9
HScSq3A2A0bYSdhm1nLKqpv0i7uJs62Js7m5jfw7SYjBMaVEWCw9eFYmKN+nvKfkc418EtRqcYGr
yN5pKvSWaWJcnkeuCiNHUdaAnjgmVM229MXAxFARMfjXsuVWPiKU9tbCyurIP9zyHVNx7/tsvPI0
Wvb/VACqvFKb9n/POTo5bRbjyaPPDXGGYmLu/5XNXcmLfyoMO/5UEzVNVBkMcahMq4p8HNb6Ythi
/bl4KIx4Z5Iffj6clDfVBaNu5sOAkRbzu1hugsRwP6CUqymfTpRRdFX66TQRPexCsLeadN2SXQwh
oTwYzBJ74cZgMSfOYRa6DQa7gYMakGyVN1j8vtIAKdHZ4Q9tRLmN/RyVhnKVgSvNHX1b+/CRXY5u
K8Zm3Ptq748XSC4EcOiec2boQ1LdC9uZBfACIqfmkppDiiHhtBjYXR4XKrrfAcnnBkWcPUQf3IUd
TbBKLWYqxyOsuW2Giq/8qmeVzfxoJi1W/NuPUEj7LOIWZe8Y8FcNc/0an31AP4Neyp2dmVP5H073
VemsdPUqBCa23o1dEOJd8jr+rF8svAOzLzgfZMFxuhksANxD8CQuzGB67egJ8ywukU53UrHC5uiI
7wJYPk71vi/nUgq8SILhwKzsXN6o/hkqcSvSLgn6mwUKXDGRh5tpGdJPsrvEy+pzfKv56cxAPgIJ
GgDZEmV8PdMvlDl6qAPX8QqGru08V7q2grneV7d9DDziUrp56HSqe5hg0+9AMRcH0bTXMeCgmIwK
eExOW5mqjBqBNp88qPHPfW22+tpDMsz04aBcrqXZnQyARaqqfVzvB6Xx35I9cNh9CCo28TW74XwK
gXlFBk6irqkA64cUthhk4ZY8rfHjwfesS50dB1Qs/HaBuxe9dF18H05ewL78G3aMzwxxaogh7FeS
Kgv3D5E9vWZa5exu6RAcQUSua6xooAm84ZkKf2zQ8pSi5oJpdIfEd+VzAzF9M98W+RaJIrouOaTD
65/WCD/L9Xvp7qHqEP958hl/R1J2erv6b7PQ7j+ntmaLHhHrmtj4yQRZskAaMLDgLFe1c4+xMu/p
tJYuVif44Q2CwsWETsyjmmcyTjz79SDR/zWM53ZOPigsGN8g7jaZvpZ5FhMn78dAPDE0HJ6usBIF
2z/EbDitdE9KseoMDTJjOgl8Z+yOSNhLMT/3Sd7h1uCL91Fz3zjJeX0byK/Fxu/l31vdr44japQr
qRKDLR6YnwnK6aY39H89rJ7eYWbFVmegUh4perjeYCZex9rM44+t4os7Ohp1jwLIMKYgfpqVNZen
ULA5STqAvUe3iWnsH8T+xt3vDEsZ46jh7ReYFRB1QlLM96PZExIU0SeBAl0y/cbcCNo9lB8jh2fT
1lmjp20XfezWSBq35B6KIBYE9W/kNlMbN+gmf3uycbhWgsC2cZplhQGntBY8NFkdN4c7AhKSFzRs
HJR2ezay7Tb8pXczIb5KJNv4ODq5NuH7b6cKG9sSLc6ux8Vnk/ACDzjdChlMaxJzhWeqs/a+oa8p
lEbyW7QrQwkyipocq+92fIWSGmdyN8jLjcOYYe4c2wyo15I6t6PbMDN+pZU5oFddgTWgl9OhnQsz
Z2EBV2R3s4a14WuHwgnif5LhnqyqMst8b0mxeQezQWN6QxPYcnYJoDS2/ONy1OyxDI1eYxLoOKHk
eSGzQpPTcp4xVX7djKm10M0vPIxujw5ZuEZlpJDR0a7v1hS7GNjSad7FNUrVupwOXKWwwpQ2EIqj
FFtg5GdH0UU4iQkApbzDu/5JOS9l6ijpUYF1tEo0CWSl3TsB69nDuTapgLY77QaSPtYVwVMGb6sl
Gp/v/Kq0krw8rQp14YySX0mhr6Zm+ISJWopUcBDcTHhd1YqTe22g3niyfpKbgoBKDeILunPKXm8w
Yshsl2xRfXUJe9C/SG3XVOSUESpAX4y3CJT2mbhJnRtTxG/ghXqmDPYNxzEInrn/UkSsQRYpyj2S
/PMgDHVMzmNGxNLFgfFETUDZLi+ow0dSpfTHA/qj9R3JdRskVF5AQmO6B2XSzZNOcKPg6uAVO8K5
rgGPV3FKOypzVEumzKOimSZUQTJ8+ytoxc5el1bhJmNuFQjPAYGb5P1DI2HPOAEPyVq1wdsLjM0V
OHIG3TAQoi4y48mM0SHbOTGwHxF0Gzs6z16C9hD4UaQTiqXSbR0/K1YjaXXK1kxM+JsWexDDq7ZM
TnDNbObBPE+rWeTEip7mm0B60HgPn7V0oZkQOY+F6CpzL8L5j/MSI1/93fJE7cq+/CIQtSYatSQ6
chfdH6UGmsr9aTCpQuyiR2M2GA3/Ca1qrhx6W3ebTh1Sh8PEuiP6n4khzsgPhiWc2E9g4Y8Ae3Ii
pzPAiLQiBNtUg/OeYcOlV2dnal2BXx4Uu25hEB7fL+x3VlrarBe8W88aLZmvvnNfK/Z4a6HDtXpC
XTG8BeAflK+yDiPwiW1xg9OKoonZGP7G36VVRNIOP8vy4rJ5zBoGXZlRb+Zv2KkMCXWEe5pB/Qhe
ERYkWBU1+85DrjE8WaTfrMhmb0nP3ALZetRcTt+oa5aYjXS0FsQiXT3KF6oCB92G1l6kDZqESOd5
xvl7qcZ7JgMNLWCzU2PXKrnKd3PEFcNUCXfzjNwleZYfy2/FZfLENMjrT7sc7FQrgBgVB/rsBxRC
qiUPXLJNsyR8zBKB2W3g53zvbU1tC19gXARvlKDXoxCkZeK2867AXwdu8vvNZiFsMB/iayDEHLMz
TMF52LhiW2i8ZntnzPmWt0fq4jfyw3hO7SJDHbt1rZcgnG4w5iQ334D9ObrztJHfcNYzCAx6/Ahn
exVdXNpPhQ25xT3BaHDK+Rnma2jOAmAUBPNpuMneF/bF1xpGMBlU67IB5C4wJhn4wvLawYlA6ecA
LoaxhZQvBNgzUBWOHin1GOfL09aG1TYtK3w0Qnhe0vLtVM5469ZEicM5ut77GpZhJuoAL8g7KFdc
+03Wog2pIsWjnjokIK7zelZx++7IGggjfcdUqIUvuAlsiVsLLqK6QT0EP3Dri8jPogiNa0cC2z0x
NeqMwPd4/+UukIwVVdZE9IzNau4v6DteigDNDnf/G9RDdHc5HcUoyeDMBYGC/1Ejw4easr4eg9hk
OSl1j9i0Vn/Qh33+2WatdFJpxwPZPKfVOn5oK2bGN2wah5v4cN2AGT3Ny/l2Jzx1wiL6Qkdd5iN3
xZ3L2Iykgwdm1qQhET6z3jE6RApbQAUbb7u1XgHUJCzmsVJ67KwUQpIABUeunJZ9Yr2t80n1YwxU
ub7WM2vHo8uXUfPT8+6uv9ekxAn1Zoc1X/JVuPPJRNxS1JtSSGksKLfw0dJzDKBW/+51LWpInrYY
CYBFWhkkyxWbBgYQpxuXagEy23qGq+8ZgNCyD6EiGXuNKYE4xP/Kr/UvWS5rNvlLrabWnTN7Fdv7
cGbe7xMyExiddadmIE6h34NIjlXKVClwPZ9LCh7ZnbqsNk4ZS+FkiUnr8ambZXC+kLw+DyhGKiZr
1Xff09tp0CKoZE2JETdaKs0C7lYY2U5P5QbPuXQCO+vs6wNwqB9nsbXLafZvvGAx796cyjVE5q+p
QBLWzharr2E9/glyJEJ5EgjEbHnR3KSlnjz8nx/4xSs63kBvyvR8hZGbUCSVhNT8B6g5tfJS9+j3
vsj3FU1PT3fr3gc/akka98lZv2qeZjo5dDkUKjQRpcd9NrX7mG/KPFHHiLcZzW9cBNsOS9HpTwVB
UT8KhTKhRugIfmPoo5t4ZNVGwgrDFo0+3zEWCUYgiUFV4XBHij7X0F0kAMEZLavp+UU+UsFiPE9R
onwX0CB64U+YN1WSKTH0QiKvty3qJsVerl3Qxw3CQH1nqYwHxjzvwaZflGwrpVJz1YFdVHK44TPv
1CQpWlBMr1dtJytDtiuUFdMfKF8f2fwNhQkY5LMKpUW1N2j6cZTVks19fNTr+HKVUgAtS0vDkr07
JFbKnvx7oTmLd86bbDoz+Wkz/iQD/LcDiQs2YUYQlPGAs7tcfUgGHmOX8yFRC5q8nFIC4YVZ5hSu
LOtTadUUKRJg0OjITBV4JZGKiR/RQ2UnNK6Pdoik3z/1/8Ml9AqBa42Xi7JB3cAkGW5nC9HRgBe3
mZRVlGnTweLf3VKp53tEdaaJzPJ8kfa8bzQ8Hqe/CTqd5qoGPIJ6qjmS/2RcH5L7HaRTibyxTmTz
cRS4lWXlUfItXZgr/VFZxPGYCeR8WOreNz03jdTKw1v/SKHsUgo8PBlyVSC3qkkANRKDWNtQU+C8
/2GFdnZhhBfM/aAMi0aYhnHkd0Vl/7tofBHPtnh5xW0jT2XYXFnRTovhkhutot+H9Yd6Eb9/kDxo
R3BtEVdGVYksX4ggSglBsJOM7INBrXi/XJ1tYtEpHwrvqpTMd4YcFEPabxuLIQbeWo79z9+zGNu4
8Z1+v5enyLwXBmggmRvv163ONL046z1Ve6BMYmUBtTgszY+ChFWmpcWpChrpF9VuvuksjpCZ0Qd7
F453Z1PJ9Djr/GVrcYaRq7ou1KnmCIKV7iMB4oXkyMmAUiMr6pxKHaOupIcMtcRYncfydoCvBkTi
Yzo/ksosj745xA+rzbbDss5JGhi+jTurBJ6BcpDD/6uKc6FPkEjsiZ7aYUZ5O+lh+X93umj85+FC
M/ZPGx9Iw8Fy0Kn5vOrtA6Ly18eADvmQmzElSOdX3tvWk75iX2agZhir/0vHmbXRdi+S7XodiLUA
jHZKiAQNMToG5JXhRdm5ZxyeRpLcJ/sd5UjPvAK8cSzPJLwN/wjRotJHIgJ3p1Iwjkj/w0ggWJGJ
viZPztmSyY2PGJzp6aHN4HwpEGFDdVaEGsjhgbqZGBp2b17Ej2pkPLSZqKuigQantLvzNtyXH/US
D/OJKy0wdNGFzCdtTF+c7z9tjYt7aU2dGpFJpdgO8JfsR1RAa288T5UCqergCJDFFQtq/w8eXDXC
fdX88U/xcHhwoFn1hFlbKYKUxH9Z9wE7vg9gZ7KkYrAKGpNeVAwmcx2tPFkEwL3X9+9FaUQX1JXK
/Z3rjXx/Q5PMH7OcoSLlO/GlxPSCzU2NdoS2ZzmADriFIQNE+oRzd1Qz9NU1Yg5juO527yXNaYes
aUOzI3jrHjWrG0pK3qlDZhww4P2fOSZFYMIz/v6Mj09r3ZeHOHaysYCHusiaEuUyEo+WCwjXj0ix
tQVMx16/f7Mo+tC9/w0r1irXYxSlS51VUSgXoQWJtEWIaYT2tX6yYiGq5legnxwvMf0bdKlgCbWo
OGKv5IHjtnGpgFOUvccr04eRctK9EvmIXspbO/EYXl6lSFUjYEDjTv4R/CUG1Eu1Wg7p8Tx+wLaL
527xsyQoozVCtYFQif0WJZeO1S3iy8/5VIOV1VpmFV/yKnURABqV9lu7S1scsXvXvHZ3waM1LYNc
nRtpWvO5yN99rP3IEmgim8SPOUGkgQJroVR8zQgO+TT5OHiVgsug1d0Q4/WS8lVdWU5YbUGDgmjY
C9ZQJZ3ECdZIqILllJcjlV50fXZMp/EWeNRfYeRoQQQW79ObF3RwPRTFI64nZuTFtLm4aZyGJr+S
N6v9hfFVcKEEVy8CNy4cjM3zwfRtm2hfSKHIdnh4Rm70GfEpVhmpe/ZgIRQHWgX9JmzJtJjObNTA
pDxRXAVXwNzrAluQRknP7gqYN8ZoFr3aF/6mSTUIzeYk/PZgS/OsYUKFYZmSHB9kC80JFxP2GnOd
/ZfqS6xoni8q3tGIu0+1lmgmjFoE14wXJwkFQ2fCKrd1kqR1XE9NncpwxF2xeSND9BAis52VjTdI
ypphQto+q5avsoQMj1g4KFnJPQZ5x5zn3htHV3l8j4kYBUb6/N2ZePFVSWcx8ztXfSt9E6mnIbZV
LZyXzoyulQkChod86OZTfjSRi+FK3FVM4+PoIgJriNbByX4v0csbmwuDP53KGb98l/VuY3MNx68d
H/7V11TQwC0asdUp9rOhgvdmkui2ZNfG47tXzJ58rgKMPfpYGPJLYE41SBBXpavJDMCj79Y5fh/3
6J770gt0I+ZknJujkj2Pg5clsf5ZQImq+efO+C8SVG+Kay9Y8YzIWA1zNa4S5bctu2gPtCB52Clq
9jq8FbQivQL3wY+vIMhXP6gDNrwFPrwr4ahIOewpPNN5/mabyF81mXl+EV6DsrgiVGHQ34a9ZdAU
zIkrtawxv+MY2iUS452lpUFP6zk1Zt1IIl57H3fD7YE+kqwn6t+tkBiJmupuUqnu58ya6c3Y2NKa
GYpkBAlFzENyS9U5m8pH8k+91H96QB+ndRgr67KMeKGQUbSiC94+LolQ18jFLd5owZz7CSo8yR9m
NB1gRL2Kx4kw25MCgjSeiT0DnaA9uchONLYsnEWBhlyiPYiVUcStZkyXK7TOyZI7Uha2SNFEY3ok
XNkYcmKq3YNQ1Hb9oN+1RDuBsJ6oPmAy+cOeXV8WJ7KAkUkQpvYCkz5rRzPqDo8i/HVP1/Q8nsjv
tSyGDC112EGWmOVrQkgGUx3nccIjIY/+yhzMrJcLw+Y9boNt304T4GfKuqOCbuCWg5MUMWayboM4
yuiHHNz5a1qrl+2qYnBzsFbbrLH7zp/LRa8VAGt2ySb96ebdUbsXZErVBQDKMsiCb/2Qa43UYDev
/lnVpKPWA8XY/e33+NTkzXJXql1KfuPKyqRF0PLlY5/DzrfThGbR1k9Cb2G5/bQVk6mZmtZcqpcd
Mev6zF2jOyqwrfVgGBRhOvTXGqrA6FxhKSSvunioiVetj+SJRValoRP5YbIcHySI6mjSaCr6YICP
jMPuqnK7OscgPopSwzvHO4tRe2HuT1ieeBAIic6TqhQgH0ZH88bYJzxk9iarKREy4aO0pCWoEhM7
yFFKrxUaVdlXxU4FMS1pa6U9vi8Kw1WeUDeN/DF/twnZJqYPKRa3HHnnWDMarvhJ9JXxBJFKBLa5
n319ZxNuQQLE4ECa9J3qXFYByCa9HJ6SzyjL8rrYUP/m1WDkQKHTcO6u4NQizbHoZoqRr0WSYOl1
Ke4GtAxrU3ScOGlodk5Q9F3oLuS7jwdlu9F0mjjhyx1hs2vHkclOBaJVougcrNwYtL12/XjRmC+D
gcY8o3CFpVGjrwH6+2qQgmgL1jhDdfbedYgu8tiLB2VGdJoB6R7AXEX7rVWwReFbCUGcnLE1P3pS
EOAGX55ak6muj4N5gAzxX14zDPgpA1JrvWcAQTMrZ+yZ00jEElygk9SNTA5MYYFYUSFpzT4OulmT
JmU7Fv6g/Ds5fADDBSj3/YHKzltE+wOOVZ+qaogez0hQhj9Lr7R4HSnt6aDRYCKrhtNxINryh5h/
nW1Hui6Cr8Y0LZUaaacG1J7HqCkMEoZMgB3Jt3txNswIvjqO7WoMdwjQCVx2PiWntfjTEsTxgUF/
KtJB/Tq3hUY4Ko2wjEGL6pfUhlCF+UAxMDQl2C5B9D0fvxiWnrHCT/2nBw1oU3JEgphatuYwPxYB
wRma/Ant/tYU6k0pq98qx6XvagV9ULds3W2CfSAWJhyKpAxzaTxTTkW+dPI2ZYKSbZ3Ik97qhcrp
Rckpn4cTUYgLN/TsFq5yqfhL31FZ+/QLIhuoi2CmkddLDbrc+85Tgx1e8LYzn/wxpim4m/acYm8Z
QZ6VmXv9tM1+jf+bQfvtYx8HE99a2mnsSaQL/HeKIrtsC6ctLGuIDIb2gPxd6TnmS+SP/T3z8qCa
hPLN2wD7rBG8FUtCho3H+y/+MZ+DtTp3jOE6s/Eg6gobPC7vcJLJ9plKY/a2OB1k0l8CmLkeVzJt
Fia5n2f8Nix9Ss2HGfioQP7wiKmxGs7zgqBbFXMXhy+cIOfR4aXJkIHKXRUh0Wf9QyhG497b16YM
qJXIKc0tskAwJXJxh4op72AR1tWUSevJZ18h6MOrxJKtoYGCZVupN5WR9z+nBLwv+gZSppszcQoo
U+IUGWvwxMt9RPJyjntkaD4fnUYoIxjxaAmcB0R38EzQHHs0l5fnzFLWGVVCNh1xNzNG8kY8omYE
4KVXE2cOMb4mi8hQfmgulAlqFBnP0MmUPeM3NwlvVA7v5be0oDHPmznnyYKr7Mp9kCRBrpnwruaM
+tcpvYb43GMgvl1g5lyiR+b4hlCMlZX8m1s3QnUkYXEKrvPeabpJgaCIx7gl91pCduj8L0fMi0Xl
a9tqAqV8YFrzehdvjQfpgId6Ds5tPNgTRUcGvZjf+QUE4EVpzpjtBJEPPTTlkem3ljVZzhDLxc00
zAXmHsA68oiIoAb02stVOYDa9ymg/05DikzMPQDAdp0pKkZzWe69F+dyQtax78fvxRg7f2F6ZhS3
BnE4toOea6gvVMqSP12b1savmaHeVVAA+e7XbPl4btiHF4BUNFePoCDVUde4ylwr2hT6l58ZyXu9
7SdwnfUc0yjzteobW3E6q97Ol7Z5VW8A7q4D51dLIXvHBmofTkEJGRG1ZgKBTpsJoOC6f5brMU4x
W617YQPWgj/egEORbNCHKua7Fievbm1NVOPq5cWtCjXZOKj8sDmT73f/FPtjMbf7cnCkflgkApwF
StX60TTdL9b9SsXqd8uWjfSXP66MCVKkKgXOrDik0YEMr3QmuO3jUyRjrf1kjesosSnswfI8IeX4
0ySB+J6hcZNTnh/fRv11WCRFTD3N7wWSgnNmuyIMIuy0hFNejHBbO8peErqIKi0OzA9vIndsTglq
gAwRkT4FRu0Ot0dmOTQ+o/OeAoQEGhGbj69hVPhTk1wdbdPCv30BhZtPzTcQcwcl1MuoAMFx02Cm
KGKk9LxkrIDDPNZvNVDYGtgHYyWLdKiwo90+Yc7SCZAt40dJ7wqSisIjuuyVVIMeCm7jOAHTJq4Y
7ipl/BADG/xebimKpUpdM2mnwHos1TdT5ntP0tLW8hGM5BRPuUlrejKEFHyuAaXK/Rzjhlc156xO
JOM83g5vCM5BZ2Mt36feeid7qIy2hvD/mdGI0hyg/dyp8e4pKFCtQA+NKuw31IGIUbzankvB1Lsm
wNpkkENmjxCIsQQsClHz9zlnCBYRCYNCCBwAblZAD15duAVdmiGOHjyhC8iKl0ec0UrBHcGk1bWi
5ZQU5pLrNyzwdKVJpWTd90tvGPPDK9mi5oGWJ+ugiDflrV5jyBy+Ac1fsRmlF+7pCVVq64jDyeiK
ZTU4M1rl+vbkrZv+axufaZwLsEjpxgeiogZJ4DUDBnna20HwD15Kb5gW3g4lSpheGQC5OjnRkfyF
7tAdo6X+uO33pz7MfkY5FwzCIJV12NKuD+66oPZG5kMYuj4MzuHp+CDTtQQJwII7fV+b2D0bZczA
x//dtgd6Pxs/Q6KpfnXXKumfAt34FCSfLaHpOAXAzIVr60LJ3x+Eh0fG9/5nSuw+DehrgsWgbd+J
8jcrlZnTcVQKstz5XA0SsrSThz/D5SjyHWgcMNrny12Hdw6Li/3YaP7a67T9kewy/2YVeFhZwFWg
gwHabWsmbAIRZyr1jG+0fMcNeBxmeW7nTI6PSsgtafHT6yNpP/z3Lwv0wwAnLkrCOLGPJfQhy+fP
RoD9VUYDxS3mMDnPRSSIFrzENHKcqYfHXzF30HTVQ6bEu+PrrZflYWpbamuORNkm5NkpyInb6onC
8JeXujgVJ4QJPNQvLL26u0lOsKsOzHOdNlhZX95uSrZMXd25myfWPjpfjpdBMMJOWRxWt18gfZGq
1Dg/elnZfmVcD+LOw/WqytaDtaa4cjVlx+lL2XNw5qAaeOEN5INny1Q2iRzzSgSx0ff6ejiZEmNR
VbQMfLq+A92rUbofjvTik6K+9/oMY4i9W+aYUWAurVa9jQkg7YLe44ayRy7ou/kXjqRN8jN2pB25
u4WnrF1gAo29bH9RWG6LID12ZK12tQcbD33AwaAXKOTd6A/kpHrbG07Wjx1Ik5YMEfLcOvvdoBgE
bRasMXmsS4t4zSeiB6YLUCWc3NTi03uSxSVMJR9yVYyUpfvS22sZxf15jw3sXYRANmem5c/6LlOA
FK/5eEZodL5pKDm9ajWgLtyoVvOnjj9XDSE81L3FjgLB718mKsD0UMibYhvocnhsvCwCIZjyC13q
FbfADderFZf6Ik/XsKXPVPz1LGIJ/XMmW+uf6aq2gmFLdoyYoagFEDc1NSYaEKbDZU3jMO3HwzOW
W7JAVvA1MG5+3JxRD19d+o7LrOUIy4s9wK8Gnq8+Qy9VqIJqZhPrCYVE6f45HJqxW8BBOk9NKDWm
M4jaqRb1NKnrDd/q3zwg0i/if+VNVKgeuCNTW2ptSicOXqDxJCZ5yAuMMy7o7a2umbYtg0gvZcUT
mHanJgiRzxeCBCGk3XzUimcs1FsJk3fc9DxJtH2UccgtBaDHXFSE47J4PgqjVVMxhNA2EIDqgb1e
cHwh5e2JQN7uOYfugunYZocxhQjQQuQpDjapxwg5r8JWArQgynPcFs3ltbI/Gdhm4ucxMveifhvY
0aCp5GimXDSalnEsKUoEPRHIhKaraXm7YImSyaIZ35w+nPzl9R8fbgzz9muDC0B9SXQCw0kovJQm
lBO8hXxmtOTkf/MnNECJAyM5K+S1yvA6TFAch2GkUuLcUYgTSr81W5MYM3QwNCFJJIAArcOR5EAJ
Oi7jK1XZN4sbpoOBJuQU3p2ESRwoO9mtDheBHFhu81llvoSdiZRnynfAIUWi+64X8QlQqHPZkFzz
HyW16yl6ZEOlhbfR0W0CjWeuL6/S7vhtt/M0tjssXpvJM0FsE684OraJhvw1s0LJ0b5mStZQeX9/
N2spX6i1Myd7/HfH3lW8LW0TSCZTUPqlxrEJ5aB4j4D1CWQYHFSi8YkFocputD8+ZPH3OhO/yN5s
UvqD00k3a80Ga6ZBXeHdU18ezwBmFIQFf0DuWsN00wY39H1m/0cDkU3JMXj96+whts7UXazjJFNq
2eOdGMDkSHHNwAe9dID0SA6G8sTtPJIgsdVYYVdRuDcMWoKO383XmlqQ/ruTJfTBWJSNqYp/4tEq
nlnUs7AEQgJUXtoX91LhmF6IXYhKZriT3GpJqNpIHeBS8TZi0qTzAjpjgvSsH+sq2DWRrVi8PWNU
O+t57ChuZjdKJwVLoKEtZaoDpkM1z8DlZOmkhK5s3gKdgODIkze2jQZjGJKm5wNLrZz9MJVORXAC
viHDvIVAyfE6dGMrUbjciNjxUWshK6gGwrrM61o8rsXNiMdtA2XUNtPG3vfKqmPmWqnDLRWdHI3V
ZC1hGSEaX1Ky1Wo+vvxbN71lwZ47eo8dFuzhLWOhE14ZnTEUPb8Qw3sIpQlP0kUvKZQ16CZGHEto
dnmNutK6JjevoVaUdyW/lGFuAJp2PEgJ21rBdmMso14THkqv5WPHMPhuyficuc4LwK8cZImM/p5w
Ou5bUwDwLu3x8uIMZe8+icVQhrFlwyvjw+nwy0vLjow7hbIUrSki6L9z8utURQphJsjieFpA6QMV
vf2XhJlQlU+OL0zwN3WQlmoe2j/MFS9A0sF68LD9F81Lr56JCw2Ah4GxuQsNJYXDlLheJGznVjyX
ClCRLLFZKVQM/1Gz5pJ7Dbv885VMSIq+oBuccs/OTsVyDPqtxBkuEmEHlSkCkz1LVdO2h7NLIqoi
IBCDS+QDKpmk52ThVfkJrxPPfwDlDqZJU+gAS3qyso9+Sm1qt3Q1wWV0x7q9yK7XsQR3MuqaQ/Od
nBA98Phor1UglO03O2zEm9Vn4D6tONQBW8EYVAE5Ue+S3BngeVQdDifHqmNSgPrkP9zURt4w/LcO
i/KM1My84ZZN9tiKdIHEyEJr9/lEm4oJuMb7t6DLV9yEAFn4oZD3J3fPyMXxqAIvqOSFG9kvDMS3
GIKEiG5bICJH9X8LR6nFdpJvZjmRS6tW6F43j6nR/z3Mp/vZ3ozERdBNalJdwMWV7oOVZTcu/vbd
wHu6uoUURZkBhWX7BFh7DOGWimDpBoZlJ/2HiP1z7e9ek1f1dpgkI9q8BOLzY7D/xKycrG9WRR4a
QbHF8sg+iQDnnU5mw9rlj3EpI9tWs4amOdSN1Kw14csT4cGY/PQpXnmKA50n6Xhuh3IhJlzP3wQk
GePcRBTvcdGOrFMU51JBBV940APUSWs8icbat9I8iVjbB/0VY+7ZRnt/VZCjm0z5zGQNSnbtw3RK
dY8OAFxIehMNECLdKwkMRBEVqCPzQBe26rxSu5v+a+N/RyzkMvIZUYt5a56dVXwjFW8rHw6VDU6b
nVdb5+v6Wmz1DEMMcjMvKFfPqNuY9UJBZcUs1fD1tW4aI3QTFa5SZtbBxesl4/5n9PgSmqec686D
yZKV9cX6wSEaNNU9OKuYvKvZlORr4/oUV5RNVW7IN6gQLyvZ6YL94Dd4a1rM5tGbI5BChV4XrrFb
Zh44jez1X436eTmy6lmjmQr3e2BzGcdrap68lhdzevZTsy5+8n3EpJQzPlAq0lI5jLIKdAJsutfr
xKhht3swBKuqsvCe7iYQn+61vN+ZqeBSj/v7sychrRDF06FpCNka7fQfGkyn+XB1D/pyiso8gz/1
LI+8WeK2uF4q8syfnzV5K0/D12GffYJarMteQmluH1oM3ZN5ZvDNXM3bceO7TWNfuuKtLrvtgAxR
Ed5XG32+IhGy6ljm+nV5cQeQ0L6wO5TEtWj4fR4uEuuHPNgsKN5GhYD2SDQWv03YvvIVMW1vAkDV
noPa/Un2uAENtE1TjtSKWUJDPWUrWk5R8ockoUvb7LQBGzR6cDNqscrJWwDwuPxhEOFh+850P/Nw
OrF0W2rtKBlTX9SLwFMD36/drIpaVQS1yDLkaxFCOo0S+RSezQD2PHESwuVUyCKS6tbEVPCiRj3R
ebWwAhYrgQnxhnbgLL5L4GRWKf12qS/fNVxKAlg5acnf1tXKp4aNGbj3ruANFZ8v28ZcvpR9lm2/
JBLFszmFg+LO6Gcql5gtvzsg+w8IcL+MWBHJxYViKw8/t61F3ob6NjlqTD3ybHMb2SlAqXms5MZQ
7yRdy/Ol43BrKCwl7ilslXCJuwlbIXiI2LdHFAkCGyO8p5ReDogIegyxGqLHAgVxQyOdSuNQtoxG
tyB0K90Ec0hQvjS4zNn5ZAmpWubfIVzCNjWAPuySjEvP6VJrfWOYdepZsni8t+yArsMTMmjvga/2
9s2lKtfhaWIVQ20nbQDXct5VNFIBSRqcWRztxD6FPuYftrDB2PfFE7ghw9dZCqYX37upsS4Yd6i/
HIF6n4RBvERM125cM12U+l4riN5asS+p40pU43pHH7Rg+KZv/Tvb8uKDj4S3g8cp2M65MG5qxlDz
3Wv7b5MKir0F8nMl+VTh4gLaBcNstkYeIWw/BiXirAC+5xAdCfuZ+Rz4NIx3PTX1w1AqbEnTuHVo
MAvoKD2RecYzcob4Yv2PkS8dyWh3715434r1FnHwhZqkJzHci3S6iYbtNR02yJu6KRtduZ+OJ59l
P5L/zicGFAsgZr/k0kscnniR31ZMquRfx9vm25EdNocvwgPDYVNKaxYedMsa0fdPMn7PLOxzR2dC
OcIbrx2CTSNg4CJobro2ISWYJzmria/QGnwiyrWnO85rcpKMn1JouHP5QoFOeT7+Z/Hir3jVBIY6
z1P1JomdA/9DjE03LpBePWcxnZHclixtvdkAHq8SVl3fOJtvyRKcvp77TV2iRqVji5FF164fQ+Oo
FKSSaP/t7hhKNW7BnHDHdIgROMml5S7zxSgM11aRZittmEzhHajUMSSSSdAGDXNcN//YwtwRosvW
ELwOWjbZc/kBQ76a6WFqPs49z1akcwk8rNN4ILzwSxiWktgzUWSbJE993dNzke7mQjQwaqOAnnPs
FdPr5nZBa5wKlYAaDw3v4UBwzsxREOSpzbFBiUl4NS7QDg+XlBqBgMhjDYroGIgni1bUARxaMabL
Cpk0VDt9NL88fw3RJE7iiVVcgK6zpJv02jQuCvCm+4prXx8raxeq4seakQVUqKTPc5MXoqeHqh5y
N+KvBqDHDDfL6adZg38mdWL0DSGXp9wNfVPq8mHBkqCyH60LqlPyXR2Fi1Y3rCCrHc5Iv5zah10X
Hu4Oy2ruqJvR2OfqBTA1Ds5r1V1nVpbalelrGCRuv216blH4D+Ck2/6z1KSuxeETSVtHHJ9UKZI7
1u5gUJharjqAqGC4NDAmfKf5+UUQBSmO/BfeJnt+ZM44gtp9JPTB+n2EQHHgL2JKl8si72qGYBiY
pUaSAYFNT+3me1KAuMeY7KlnzUecCkqI8c4LVmLhy6uyLtto5crNL8wUQbx4pDRr/Yl3TdXGD+eP
WX5QmvRoLqqX66EMdkMvW40JrMTXRRRT1PGNbED5YYlA7DbZDhA2W27sejE3U28g2SWQFp/RA6jr
XBTaEe/QH2bmIoDmaoN9+J7KnE1vKy2rfteTMHCMxZoAtB6N0WroImrHgp3JmVAE1m5vwlOj0Qux
loyqLoYDXBXwLVtAGqIK3z6O1wVY3I/NJnuSkPnSge0ykHtI+LbBrP0TRS8Bj/C8UNLkn+48Wg6Y
XoocXAgfUW4jwsnhT6j7xOatMTFG4q3OnxpCs5LPVj7Dh/Dft5NE9qmvKkQTDh2oa1MR7DzSop/T
UKWEXKQ2frswxJ3iKtX5Kr2MvGlxnlMEZs1mg8luOG5wTUw5nD3mzpoY/V59DW/W54h8/vxvKx0o
hFsjoGC2J4brZmufPaBwOgnsxSj1QyHthPHUbKa0ROVeZzsHL/4QbYY9l3zRdDSZfLs01alCx4xs
fjippS0sMU5TTX02qkUxwgxVcoRcclf5t39Us41fFURR1G1Z6xF8HWuRLilvYr7dZ9WBwYJ2RHpm
dcVmWcIjVEO9IaPS5I6Gu4gNE6pjtDILUdBwdF/vwTz2ocF8Y/HPAmBo7gqENg/CyBWRPCTb68dU
R5bPg8WuE2q0GVFXtqVaI3V5H904HscLRz6tZaUkFsR6MZfZiMR5/ZxbR43TzEtjF8aDwjOUKwSM
I6D1FzXRS7RsLZp0FhCRpuje8KmcbHrwFNWX1Kn9nV0X0zvttcgVJerkLENgn/EqAAa2wzqa6pal
ZiLAtHHH/ROsoLUunM54j5FMbpkDTWmUQSxm97A+Mo9zwuu0x+Ac/Nva0N2nTEsrO4DjHMeRzNe0
d34Om8BvxiZ0oo6E90JfWd5RzdiBUiYtZCM9A1LkaGh81gscg5lQnQ1b1J77tAmnzhtpHjq7ldT9
XLebKbRuz0tAp44ulFnqnAz1Eu/UrikRXTvU+/ZZgGTrkweL/GnPixnCetcBhuAx7fwprhbU0s7z
P4WHb2JWJb8ywBl72wG/lJAzbyOE6uNf0Y7U+cr88cS13EsYsVfyO8yujfBF3imKY/V26Jb2RxkJ
QlBPV3zxc4ustGpz9Rqn4BNQbqGRcuKuVMxyjHAEOlbEN5rEG/rIMp/Ol87ZorY0M1ABnVsBsDpY
fAEbOHeax60zFlj563PPvwTvDunBHV1QGZOeQiZFOnv4zoMp9MQV+EbPOD0Pwt5Jb24BbJckDBqs
N1joUStTdveoSmuzxfxgeFD9KyrgiYv8kSMlF/3TsLvZOfEhC64+QCu1RMR1/MwIaJcSpwXWVliT
QFXMkJ6Qny3eAjaARCNFt6q1vA2J2P2UnvQVNGODQIFPFdHzIUYaiqmdlv02jaeCwPzFQI/Yt7jS
c4GsYhHfMoNxt+xBgFEf3uOi/hd6OnjH7cEwru7DULwwK9ZWtCIA3sgcilfEop73w7OwNH5WiJP4
qy+DufelfvOFfUg7426+ZRuSXHAQ2ADmqgSsHT+jOF3gqwoXlt7GuuQcNBJ/gYuS1VbMrl6CA/XN
WVHdRApkzKAF3Iq8ziEBJjgEQPBTfT3aXJpzwP6ch0FDuvzEk9h2LOHBBPiWR+P5ur7ehbHXtuLb
cQMNwwCwnuxVwC3ZidUYG6XdJWkQM/pp8hKp+t2u4aWY3wCaq4M6QWMSC2y6jClWxxEFmWUgpzFq
T6kParc4/4v/vNC5W9H4iW989XxQz//fkOHAXcrIwkfyIo50mHkI6fXVs8rTqnN5gZZQXbibbK/A
wIJEemb4+TA0U2jEQ+VYla+s924fOVB5bn2e7d5oBLAa1NulynzVvzv0nQWMWiAQV97bqOEDfGOx
QTaGtTVpcslFJ/JXndh+YKGeJKZ3NAZpjm6Nltim4UxDFwkQUyv+kbS/9cMxXiVJfUAJ3FFyddzM
HVn2PwjmycujVxZP6joVl3Zrag01anh0uDlnJQpvJgL3XgTZ0Lc1KlZQQKil38k9AjcN/lbsEeYG
LiX2bvo+7mHadGpr59McqFmdJavNL5L8vboO8sZzrVk4adwAUSma0JZL7zSAj1Ft1ChOoApDZjcM
UZ8u/9XqMFKcipunAUHBPX2V01hqd87BnZwVr2COqzfU9tfJ76lqEhU8QCgr7DQLetF2n7WOJ3Kl
pUV29dvOQdDEtmQJw4e55B1w3+K1fZdHcYsCbxN4USbPJ0UGsBXvgMVAN2t0Zl+z2b0tJxkicftk
jkHQQs9UOvzCgU/ogPsf5Z0df8Q4/wyT9lZoVSkCstx8DGDdDogSiTRVQncddXlWQOmOQvXnHB7r
ApgbxaT8oRyaXq63IaoQ6Ag0ziMV9eo3ULzF37LcvQ+tbGkjIvq8Aq+leO5fvDTZDmYmM8raDGkG
SjLVh+RMw+QagqZhbtqNKcvzpcEH3VJDCjWQGVEjxcrHLDLLKmXAN7wZ0p6nBrk+zUvHU+THPMUo
OO4P2hTfu5tVcIbw6W1NSwL68R5oQuo4nuCI8zkYfrmP6TSVtl1O6lQvdbstXE/zSHaMhQp5bwb6
IhITuhBVopQOC5X2BqJF9vTUv7hbWiSoUD7hsL++Wsx7YxCc8QS++5nPBg0hMIqS+dAqDtIGR99Z
JCccdYOAp3zMVlLBl4sWCUpkfg5CxOZEp415jJtoZeaqg/pa7zRyid61KFTk0/FaUe8LSOYeG+ib
FQ78gG7YbAlEJMwrUdfMMDJD9izETlGkkcDO9DhmOGsbTuqMNfBs57Q2o9lk2hoa1HZCpD1y+ri3
UG9w4qc73JQzT0kK6bsidwQTn7nn1NgjSHAS77bp1ZRpMYw1ha6UXCUiO9UiBqWXPj2mbygbUB/s
MnbDl1rJMZBiluIweajH8tGZmddgfbR5nrE41EXFReuifmyx2yGOqghidmvkoUFcL/GKdp7Q6Ggb
iv8HT6wfLYKCEopdC8Ez2ASSiyRv/4Lfjbi7I2dAN94EPXllkmecJXOYhLHlNVgJtOGRm0B+hIun
6GcUbxDFCtzEM1HePdt4kNvn6Qft41VKxGw1VCFUQUFkO0YFuPRt/ChC70KdAeVQE8+ycXdjFads
EB/I+m5JEoDljdsJlNkZQnPiaqOrgtgL7a7uHBEY5DDhD2AxTSuzBEO9RKWagSzVc4lULeEHjtgh
yo3AbVikkVx0ufsh11Rx2E979xsXUdNHu3wxRIkWoSTEMATUIw2et5+y92cVSMTbprIpFz0EUhQv
YI2yANYLSiJgYp5tdV+c87TLwtcE9sp2V7pLkwAhsXmfZ1iNK2H/0oZBAI59d91o/4sUyD7jdc33
rYQZkOfrFfLvrblfGzsCtTv0s4r9nhyvSrJPdOM+J+kcXEXWSBiAStp5gX3xLMv/eby3IEynBmI6
YXQ1f1OnqhbJuAUzP6YvGlp8JqcspljrHY9ATyY6owh8JmqOeI7WAL8SFh31LwLQakl5IPt0gUM0
y/auGMx8DZmoaAT/Ac+RlDrYfp3/Ds103O7/XfsT5Ox5dCOMm/x5TwKu3Ouh6fST6QqwfbgfB0gl
U62bzfu303f8RWlW4psXOV/wbjSO3tuhfyBkZvHoWLS+uyaITB8EYVtb5whXmqMDGOOX1jWUjnUy
pK3Jx1NrOpUk1FmWnLKOptbPa3WWgfPxOK5ogKEGZsC93EVaF4cZo6WdC8P+q92irZ7GzuESowD2
MrBGNt6+HlNRh0pQiXnfIv3bpxcpGaUnuCI84sWCKJydVh/ILgt6qRCVIpQMq1xT1+PZtDSgfeHR
ERVgM3om2GKVrHlh7blA+qgK3l7PO5Q7QdV7XE3fMgM9TGb7Ixe1Y6D/Ul31u/HnmuM6gEZeJ5do
XOu0WYnZebm8yyDY2lqvWoEQvJnZd8m//yMhTrb4JgqN8TZ20ZuRCt4+VZ6Y/7SAeY+X+Ka9ao/C
NN+IrlitVgxzvyKZ2nSFQutkAqO7ABElyj+b1dIQbIT30YEaFMx+rA0WTpFL5DW2qBTwhoBOmV/Q
Xok7wLMo0DuK1a2uGOqUSEiz6M8xT8PoAZqjGl2Grv491rTFqUB+weJhdgev2KwoM1wBhGvjXa3I
wiJRTbyKd4NwgvwOmXExjIEzmC6zmXB/SJTP1odAktsnj2emUw5sF30Urh9iSLAHaQA1f8o7WRox
0oKYdddhofsb3RIXeuJutNeMw5OY2qCMQqgAKTFPPuiUchLYX4ObjGYYoGwZFje5s710U9Gcm4Vf
mqXZulGO4KTnjYxBdC0ltuNoMRicnF0tl975wLKuQixtTD9yekW6ZHO552zSvPrtMmjlCJI8Axvl
2k75Oytkn31liJaYh5stHNJcmEcItdCtog7vP7MbNtj5HpmnMg9qDbdeKifALcLL1CupYWjdZ/SV
JCNbOyQ9lnaSCf2SHl3G/KUFDtuzPz/zOP0XzRY1YVZTfBTOdT4BF9hZhW+rpa06/lIJxeepsP2i
flpQkCYlW53VBr00uhoGnIzXN/VPLDkEY46xK9t/bOsdoENlbdLGRvc6AorkZ8+luOmTxx/v0znw
arm6jgow4eCBdSr53RppijH3JAcanFhRE9/iVXOu/0HKbi1x9EBRMTcGwlmg5V2XvAu0S03g7ydr
huW1z1fZ1xWbRTBf3csFuUqZoNW3OI2cSnjoFGTaKJmQryitWvp9DG6O1iv4u7Z/rWTf0dYJxYd/
avzUcXuBC2G3u3QimD3i9h+0IPbj8SZGo83rwUghPPqnODC9+P+WxaVjrdLjbsfAObHQ6amY8i4e
f/N26t7OAaYDA1rikhEkNS85n27W9j/goRp+R+bw9fin0qd7REY+queeRwTtioOAtnyNqsnjsow5
ZX8sgtQ3c/FHZWwrWB2UbDsCwLGh0qNrheTEOV0E3AVyVsUmT0W9QPKNyrpqiCvBXXMLnI3Ud59i
tN4g20jtPJ8DufDWS4NEbvB61Hd/T5GOa1j8AdDVZCMoHL71MOjqBV4DYcrxLYkIEzj9CTT27UTL
PKoD2CF3rAu1w0F6aw9Mt3VnV0ObEz5CFeCbBGUmqUlkttv8Y4lVhuFAdwZCaDvRmdU8Ro9yIBkl
sTC4s01ijMauhIJkHPCI0CcdU8gdo2QUz0LcbaWtspVHr8/r/PuHST4oDIh9ormQy+sTCacZizL2
kYj0nba2s4JPx3et/7PcjGIp4fLgZrxXS+l4oBXccNpRd4iZTHLE3m7/UM/wf9gmbELUK/2w0N1z
EDYx3FR8CrWQt0HRugKwjGLexshD5pvEDx7rMzNswdN2Zb2f1uIJ2idlG3VetCBiVgSRQunnV8yl
DMXZDgqMlHCeABBajhEXAFj6NHmBHYEgyBYR2656RYeZtfbbpIaN/hu1KWQ/YEjDoMi0UtfviWBR
IEj3pt2kWArJFwSrgQaCSnclRYEdd1nI9350xxqm96xwsz2W91f32pzpJTSJFAyGog9X/IpYJyM6
qaaiPTpw463pj6mhks8ljjOngmM4oNvI0X8O1adQ4V3WaPzX8M8tvIf7kayXiD79AIAJ9BDCheEg
kDjWiTKGmuKgbUa6CnEAUgKnVWXnO8vsX/cCrRM5+MVOAbP2Y7qcOug2TLBkm2lSWqUXhGuyMKUq
uGmf1noWZgk5E6IMgWQq85pO7mN0rwIt8VdGPQOh5peGQUAWo3oqbQ6+2pBv0ZvFI4yKbJzcHYt5
zob2KHBbZCmKsI/5dut7FKGAELJaSb9mIbQhXvjzA+r5zQowJ839ag+1K1KpDRlZ0GIxAjdlDfrx
v/fGJXydLiCZl9jFBFO6o6BL3F3IU9kq3iTUjy9vHX4jABJdaqVhAB12IGb7/YSgWYBEsOxO/hgu
i4nmIxDSO2adCuIRBqnY4uXpUHhcEDmLvWU5AEfB2NJS8zJMlrNGsD9SqIVuzqlcsxAcik9/pZ/o
RR6oWiabGmePlp+fKlTSLulidw7u+ZHe7j15RUO5bOycxOkr7ydrM4VrBTcScvhAna3woXUwiscz
g44BKJe9xmBC7zZR7jf6o1hLnB+cIaVIJkhdWbdJwduJXrxOiL2DBcTsNaXH8wMs65eZ6QY6gSa1
T3wDFe7s+t3+tFXEGJh6AGx7kKxsJiANuADX+U3IJbTvgBI57cnRtE1sZ4TiDz/5gGO3DMrHkdfW
rF1UlnYpWvTqycksqAFaI9D1W6attHu5iP7PYQm7CBQyfVlfgyTIbdboNt7djXEleTBh0ktroJ/v
UCOl4PBH+Iy2/TRLMPCpsMNdGoC+GiBjEf0mSaZt3sM11/NuLJZ9ogv4JHaC0OaKcWDwN0cQp6TR
nfEvTP5XXTBZTBuOnfBhkK87IR3PTVe9T9hAZcrA0GG0/yarY0oCwfR4HDPIm5YbSYGr6pImZwZN
eT5vVYHYq7yauh2M2sdWJaKFHMhbU3AOEP9TXGlvKiXFheVKQBa5ee6Ckug3JvqtZD5bYjx2EeO4
Q5chfNlRfwxD10kzanlRoQEyGtgiSt6wOK8d+djAF/ASNjGPYv1s5dF7jj8KUEzmsTHPrS+fM8WC
3OAJP1q2w3+93qMfax3Y7FXNwZ7iJvWe8lJNPuQsT0WonWJ3mauuwx3O8O/wwmYHjX/9mYx70C3P
FSbX/W//2KKFD4kspQeoTWlLbVNWf9DKc2NyI9dggFUomrQAGiTvZEAejax2byXVYdD4y/fEzoa2
hc3euzJrHOtp5BjuQPqcWzg/mI4yAZD1Q9fRJ/r/hwQEV2THNppErOO1UrnxngitOKj5pMBUdvty
/YtC05yavEj6CZteKwNUFXAaCLi84gA+suZgBZ31c2m9zEgX7YafO5mYxFoSV55m7u4vN4OVdhzp
CsjToBVH4xL9kwSFekZJdbkU1s2JVw1XY9AfliEo5rzyboEgbzYqwforareRKu8tRYgXkhXDvDyE
qcshsto8xYjJauoILsLsptlmzs+juD2imw3M8sqOxnheKcZKVphCdRCkrD+x7JxEjMrvU2F4j2bz
QbOp1T0IJvRB3xC+oriByA+HJhVR5DBAizvbXs0lTMfeFAvsGgYsggdTKSWzxPVAG0DI5EevDa4r
LzWCqKoHkn8pIhiqEcDTeWfLWtLvjbO7SY1PKyzrvWX4M9joEff6C7WL6OO18ebYwqoIdjO12IV1
QlFl3zaCSx0VOg/8qvTQIDu03/MwL/XDyRGRxGd4Bb/qt6BwM4Vv2KhlBJ6D48lQ3DDPdmRZuRZA
yIcY2urE6/m76BaoGbLhHmovUZ4CCPtFRwmAGV/kJhwLvlXA/dCwGCeGSxKL2VIvY3+nslIeP5Xi
JA1ekG/o1SHEy/1sSgJZ4pVYrksr2s/4Ye5Pab/SCo08mi+bUqS192ZkxKYyawZReNim/fZCSMfj
XDwLB6uDmooO1cHIPrP0use2SlysfCCoonb9qlCo3UjqsD2D8aB7FGKF5Sa4WGhcw4IHBTZJS1Jj
RwYPldyOMfLRj+VQ0o6SDcY56biR2h7g8YUGGNu53NjO6hqjA+Y0t2kqW9HaZ0DowKSq+oWie8Wp
DgISKPCZbQwuk9F6zOMWKmUYVfnRGn+MU4Zni4f9tRCN2I9yywgJPeWzivhysAbWH7N50Wda6UKM
Yk26NB54zORW7lPj1X7DKt7iZycH2N7RdnCFnSvUGD1KAiXi9odvNyhGLp/FiL1lxuYaMfQ6taEw
SlK8irtdDKW57AN9o0iMH7YRsDLjR1PHWezWYfHJhVYn2BQWmEdzwcZzac4KKoT2+TR9tn4kdL+Z
pBNydeTxsshOKdxiJvgfXe7/ZO1tVAhivEJrI778csCY12CKYit2nmwEwn/iroLFVMbl0aasFoja
byIA55/S6R7K747qARDd6wIKugQtm/2moVD/Ycbl1x28NwEdzsC8WN+0CYUGPvwe9Qs3cQTsxpdW
05zm9Z5XSQ1sif+ido1Kjbxjx4sgZaDV/wrtuwJenE4PeTwqvn64UHEuzY9DfeBHZ3TYg75T4VV4
IPbQn3XBmOtzxoyGJ6OFGmwfOQmPSzG4zMWBmhkqIH8UHf5XLu1E35xGvICouwi1dz1jp+nuvQsL
mhI5PQRHJVFpYmcm1OFS7IcOVYC2DdltEpFZ6cEo/TKoqoK/awgvX4Cwy25pfeGZ8inDpG2iClRK
U/T9daIuTy/7AU8PLa1GNchjeUheyzxJ6gi3XDvgqlKQXWG11Ij+04ZA9cYolH/u2quv4slTwHBy
UtNnxa6G18ryUQ+SsY1jmLgFUnbYmHB504SRpCBHkk08+6g36zvDAqG7eKIo6PKslhqRR/NzUlFn
femXitYJ42FYQCW4mDaUce2f9iLCCMYXayPrvDqFO7TivzUpRhZJ1N0rGgodLelCxpUWzrlTfCan
K0TU0nuSWoA7aX3q0gkNG+dWBV09dn7u7dwlCFUnvy33Ksh3qcwX3ny5xVUNRzRZWJkVL2ldtGnX
W45qTje8Mms7JZk2izxl5BeSWYzu4fhnyjANnM6qequZRv3gFIuMR/6MmdiukOxCUppRhD8XY43u
rkUECIRRHSttg+bK+ousxJK1sFioUGW0O7pWxt+SEuz8rqsNZdMVNF8niaeX7e0g2eadeAhzuiRK
r6Gv1lHvKq/A/CipWtaAhedYGmgUyxU9+/eFZc93LfYTdYUtx1ga2a6yk1T1jKz8XsyNavf46cB6
1/TNk1TJRRQfX5cbBfdY8eaIMyy4nkZ/SR83KBjWgvZt4cLGKtqBJMB/u1X2E8qwbG7YN8EkLw10
6mYWOte9HPkuA1GA+a3xKJhH2Ge7IniOxEiTdPY8GeIfbL7oDEAnbbpt4VIZIRrN87XuFYN72u3A
ky1+japGHoqueFNlHVAchdSmmKwiLEekeRqlg/mZ7rreF+tPWnBfwiO9LNtVbxlDqv0Giay6xzwV
A00wQXnwQH5ooRRA3h7lejlJUOqAMN3J/Eee29li8CAmoOzwl3JIUshQMddGnegikjdqqOwVVJR2
03pAdeHex6ZxGy1xtjtbI/YzfWT+b/egwXB4hr+A7jVLTzo5MX8zA+6jDx30GIjG2DGd6azozH8H
gCBceJZZ04gc6ct7vmnNX8AAMGHPGGvKlba1GxUoiSI7xW2H3dS+V+FM5M6BuYNN9QCadjOamQ9+
P9/089IfodNeRqXl0ipgm2BtOBoMzcJThZlxH+yegYE9LG9knDtvFfnb/mLt+bYQJvQ/+TTJsyYy
aV5ZwQ91N8xF/JPC9FcovnSibaMMvDoKnXI0NkMMwkn5VSUsS2P1XS7JtlSyAa9F2nSXoFmoz097
hdrk0td3gRNO0WZe3KyR49AK+xsB+bPs2A4iV5dLt3JndWzg4Gr5ghPxbc8gY5m3og/Ukunh+PX2
0VxV1AHO2Cy4qyg5Yzs1LLP8N5azvXRH93v2jf9vwqM6G5CWxvqyAEn74l0QfayISo7Hwhr9Edk3
JSUyUT8dFsrJyDbMTURyWiI/KnoZMbtAaV/8qauXguyZupzFGvR621+8aric4z9pdQIpdSiJ2xdP
f0qDqSVfVQEyuYv+FajukOfRTDXvup0d77lU1OgYm1ODRlg/FNGOUbBvuRdf4rIlaEtJIutUdWZf
RVoHnKcWMFT88tLal4XbJEKXhrfnKNtyQrdjgly0i5tmb1QgXed0P1anQEzUWS1nqFuaeGoCkoqJ
CT+3GFguULXijortXPYG42kMfw6kqofH4SoYrwVYT7oiz42tnIa2ewrOEHLcAFvPrTKi5cLgzM4m
pbpKSrNmDi3IYQjSteoaI9I2vndQpjxXpaEgCRRBqb39eOwp44ZJroXMtsBMbUpAhbfwDHc1VzTA
+1of/RiZBoAMNHkBWz6UMoLWPYlbC1M7XMKKO6/phydvIIW/3WzRejx4/+EVCAB3hfONHW+UDUwl
aCThx7FH66tnGChfr1nbkbT+nfYxfMafcxalsy3gDIJ3GxJxTFjczrf4oL+lgExOrjwT3BLG14qB
Ldrt7vY0pOJslSm5I5PeBqGkBS10CKRw5Xb0RuAwlc9Gf4qF0AFG7RH6ly2mQ5KYwULZYAkbjM87
pOHuTfDRTbmd+ucaqpzqxdGdRf6hlXnvSBBikpGkP0Fl8w4mnO+RFZnqjfrb8aGj5aaEai5UZi5/
b2gh4S81Xdb0xemVSsgZaY2Ip4uV5QJLpwBH8PAoMofOsdo4yG/CeqKKtlYuT/aZfvdTOAnmMnQM
PexXwA5iUHQXzANPCNxCqJsx403inlXgUBOzsPYXgKbDpBS9nBjpq0JvYpfsZmCnmqtzmr63V6Xz
MDe/NDn8vYTM70foohs9B3+sTY5qNUYybVK/6OOvmQl6/QhkCVQ564AlmCr5YGbknUjz4LT+z4FC
PX6RZHSIsLIG5tG8oz/vHsOL0MzdHW5Btuix+LdefzPOtNzb1cHN09pmyr6YALVPyoPGvEHTYSmP
un/4Ys4dBh3iowK9KOn5o6CkFyHoLo6jw/Sq8z1iElDHcrVDIAfgXf9EXt2o7GULE5MR3/Dr47WQ
ycSsWZUNABg3bckUFBgQAcyNYnhLaKaD0zr59AXHAs9WI0l7UwlVe8gAQtdygOzsP7OY7jB9h7ws
wUSj53OPF0pazlciwqAh1g/MBrbVSzJZ5nXd5aMY+MhtQs1jLlNKKj2chPNN6f/OxrkNE5mc7a0r
oXCzkq7GXbrr2v+yB4ZNcC5uK0yBUEbLlxbugVxy6jQHTJNQ3cQ3r4g2NxVYq5FKCEAt91PcTV+9
Ls+/G1OStIjfzLvKQjHVCMeOtccFHBNJIlaIj5Ki2G+27wmD9UBY8W5GY91Kw59csnIB3G/R2WGA
dvLE9NSkQdbFS7l3Gte3d3qQCxZjTrwnrJ25K/hainmdCSpxBkxOFXMov0xkXXCpaKz6YhRRXdLV
z2edk/c1pcJmfRcXPFvO1NioCrZVzQJh561AMxESlZg+SMsfeiKUlHLxkdS5U6J/un8mbchOSeCp
D5QDfe4tjFjJCrhkjvzGWxulzOzoHBpgtoWCdN8WOHWDUOwJf2Pc2VyzPXanMUPJh16k2a/anp0S
jlcSXuV3hid9kJvvNTHaN/j0yduoZAtkTldKitO90Sep9Vm2PAFTue+PdqM4QHPFz4DS9E+HJ2Rh
SRlAETLAkeIxR89/TzE4jjiBcx2v6BuACV7HaQY1ti4t+JE9gUOT+0IUugabFOWfLILeEhyFkHrI
uuqV2bathZoJSQHMC2y9bM39A1QClrOMBEgVTtJp+aufYfr0XAW6sxK0i9JjWZJtT99R7GIYpnRH
M8xa4Ba4zI3ChsatxU7bniSv0RgWMrg3yHewbZ+yjMp3H22lCTsOxXWF8tlAP5eR0QiUTxqaqMiH
eX5foyQpX7+yxhXkdvhQ6jt5sug4IHD7ZlK70Tli9e43szjRXxQTiX6TbFxqNHTn2P7DkPVV3hCM
P1+d5ftjUyKgYecKr05eAut5sV2HqmUv3MskhPBf2I8v5dAfgahRZZuOA7UUIKhjeTcVK1uUmtaW
834CoIpCYt5DJHda3nlS0C72r7BoAiaKLahUuMG7BjJf9GVjdM7G/j0r0X3XHGXOMgJ9kn3c9Lg9
OZlStGBg5xv5HfPrqZV4u8ni2Mob9BY6vgnCSJT368W4u6yhq22yQ1nW/OPSf3ScI/r+OTDzqIh1
tq150jj1DnwJ7d9xbyUJ58XgHXOg3SBydEB2FUr35uxI7cZ77O9g/CGdj6sMtaXnivAQ0B3Z4f1T
CAS6f82W1tpmvQ2KCNWkfBCV1ziJwYoUTCx6LjWYNGDBJSl1hW8qD+Pgk+MaIykF/ftkdUtai4GV
KUFsn6+/aoRsJ9PgYyIBrS8LyNxHzTCOhKjHIL0QWBY8VsGiLVqfqwr7tKcHCsKQZuxFJzOEnvvn
AZ3FrLfdEqq+kOqSl6YpQDcMHqS6WoDAQaOyS21aaxu/YymRcT0EZ7zTrBMfGaQNswZ4AELVv2+N
2WDkhmzgpd5OQe6oW/5dodN9lohsyVOioDBJfOXTkISJqX6mD1YXu1PEOXEo4NbYFSh90euQc70F
NCwvPcrYz89nitqlqN+xEgfjM3Y64otm7D7O4l7bR0Hlko2xI63TxfA3dJv5WZ9x+NsuC5DXtU5F
1KPChss5+ujmjrL5FyBoRtdlOAXDY4RHBfjpAtNgJJzxeNGW6z6Z0L2qemjA/rfULNbb0iKCglyK
BQnDA+TWFJJ5VG2KmPtOzdUbBHqNWES5jE1W0Yd4oA9wKdHyIhhfrYoNFiGMU45sfg7t0kuxLNtB
VcDUqL+OGJLLcpey26TE6IXZzGzFulD1usiHyN0mmphVuMHjJBgs5oOhNX/0c/B4wzC899z6auxH
frJwKXSlH/EKZj+SCikRZJJzAgqdFthUv5jd4AhVwEryulxjWP9lKzeCxgTILUx3+7aePQm+GfA5
4IujWfHGoy+4iTjgs25cVljrxckDuxyv0vxtw7CvA7N42n2ll8cJzUE9yjc8JL0vS7k1WiaEYwVQ
jzuDkjUaKLLqerOroAAKsenTtUV01uPovV+anCHka5cnngy35XBQYsiDuMM8NWu8dsj6KPlotcBH
IrBAyNFu1Psz+VqMT+SAmPPw0lMbyk8PbW5xsWWgnwIRiTPx3YFzswP/dbseDmbhKmDfe9duvq8T
fglPhHx9Q9puQgZrKBm3Oj+wx24Zz2Xd7WJNBMsS+PZY+UY6HaP/WAUJgC3CCLgw/GM1sx0ONc9l
c/loLE8XMPqwPFrAgGOIxZ3rTXEs4iUHO0a73TZdzvzZfz+T/0bhn3Lh7yCmGGGm6ollok9FANqy
8dxAp1Zj+eVepLSyJfhFpvASsMe5JbkD03sliBDWJ/0HKSNIpuQq6EaEKwbOMbl1nnFNwCMbsCOq
/XWm3cojpQOFBs9TCMSAohyRoeBHbsOBQ8EjxqEtehCH5fnb2fI8hea7IdKTvjiy92dk6aE2QBUp
U4CDXxWlKDeD67toQGhDKLpoSN6zNqsa5gYWOdthxsMbpnrON6rQTUX3CWkyMcdrpa9PHOZfpPBj
2jNnH64eJwP6GTsjYY7OimRmlD2RJDwYf2L78onghZayp2T9VjQBIwQusg9ylBzr8FoZ9O0Kq5iX
R0bSq04c2JjYnGTl/z7tSLk+CpVkuvtCBcx4w9TfHROetnSROCtln8bgKCWzOWYjkuzLW4DPrv/L
uOikzpm3KeYuAp7cpA82aURE95P364UdjPmAN3x3Ycc0IqXGIMjNpnAN7kqFNXHLBehvmHPfcqEO
q+0nEv5Q4Ser5Hc/SxH8RqRoS2gERk+ZyGCH4Gwwaa5G5QhwqsSWDBN32dMwXkwbacv0XHXk3OQ4
hSKd2xdGkA154QFvOswqDuBY7p/XnnbDmXyi49XsM4KRDS08UhDE18UercmdKithGf14mBF8t6t4
LiK8Yd65yS2bSnlJdc6QmIKaFKKaMxqCy0wRcNNUYQnrMEfcokasH/n1TUee59QmFO6S+a4to/BW
+IP9mlCEynxx3gY2BCf6Ej28F8DXtqMUXw+54EcVi3jZ0Jpz8y5ptj2dSB1nGbefMfQpz/uMg5BF
vALq+oNsoOGKq97gi2bjHADxCGis4LGZCtqSwYJO/XwARJub/uT6qG3QhIM+hi5uON0f3rrqB8Wd
VPg1q6U+qXMtWLMEzZqxK4G5FdQQqDWDlEY1PLB74QU8q37h8zHmYYK+XQI6pSMTG6ZggGhKBTID
Rr46mDgWyrXuHOAvDlw5D6bFl1BqoVXurZ9uKGxluiXR6hSz4rmQogjH9nwtOm7gipZ4EF/04nJ1
v9rcrcaOFcJ6OFD38q9b38928UK0xIfQ22MJSI/2B+t217xYFE0uoQa1qRGNHSn9PsUOl+E3j5gm
SJGHMxnf5UgJ3DU2gdY1jAFuxQ1BJqgG2uoMJUFaaMYei5q3S0tfvVl0czFujoz3C73jYWwvbMz6
aOT7Vf2Zh+4vyoS57eMnj1Ffhv6KIpqAuYHfr5m3m79obDPHrmixtRH9hbdHVzCMt17T3wrv4Dfe
/StwLH7kheNqVQRIphGEMRNdZt/gJeaK8O3V+gkEY4WtI19Z03sduDsVEPKbt/+yXksliXXXmGuw
ABxeu7VhX3nphbwIBucDZ5oLGAKo3Mu2EqA2FS1/yKbArNJ4Up1UVucEoim5IZskiXJP5cXzMyqh
9gDEulo810KiECFUkY2QmHqnbeIVHHoF76co13SB3mFqypLIWI/J9V3vNmtEV3vsF0ntniPn4/iO
SkDzP5sg+7zWw4cfiPk5NMe7m+/xlWth6qXC3E9Efym57pYk30YbIons6C9EgVh5MPymdvSsLJZp
nI5RxxNraR7HjAwXfdOSLMhdrIiO3cqQ4KavjuWeQh2Vrhw3bd063oPSp/2Geb/vAfJIerwdPo/n
+ABzIYNuA5BEtOd/inL8EnHUm9bXIweVO0t7SZHINnJ8yrN37cXDb1ahAmCExXqyrKtkVQnlojsX
M2872VWliDfVyvUU9dzGHZUdKn1l01QrnXomivU3gYlzX9cP76ME4+NHnXaU5EUmkkvTlwF+SvH1
LQ7ydHOSgkhAD02MM+61p44BymkiCweedVBfm02R5TcUD52Psgm+vyqkLBpcOU9forZW1j33Xc2i
guezw6Q9ERG1qMQGSc7d55blW/LErQAHcZQYwsRrNDFhIJBh7NLFeZDcJM2YP5t43jZuEwfMrjxy
t+ZcdVBAzGmJkdnOZqXIrr68yMsyd8sHtTRacsu++mg5C4noUcgdpY734e0bkGUQsQTi2ntPN/si
lIiVM89ciT+jQ+DvNCEbuX9eXRGhaDfPRh5pniWHruL3Cbl2bPJUCl9tZEyN6iXw2X9iO/nbPKua
xKV7KapLLBO/haYc1R6g10mkD+kfAlQnrehs7NVnBAYlcxAOm25GEimPdcYx/4glDEf42QMpEaCH
lkRavUUTM3ub+K3f0iHLbq9ywq4mTB7HTlkcy8oRbbhRJ8kFnKzFJqxva2ZhZ4BbJy6Xz0J1Wa6w
+PgLBc1EcteIv/VgQKy6CKcU9714pNVl/4iNLwoo3KpwrZwamozkqSRIfI2WiK+VOnfVFS7kSZR2
qw9cKp7K/FvPbkPlYfXWDpAKHfgGmpbb3eiqSdOavubHkg58zFhmiIKKOD3p7cMVntW6jk86uXOs
+NPY6IORAf7G1aTyioDtef9kv12/7Mj65pU7BSUGkP5GQrXXvyXJj1kwk9RHnAxzLvmP4xtXoNGw
e5EJgG8Kq6HXSSeXz0KyYtqaci30svCFlZ1+bEYNJuCStA3egh3u5U4HKenSSC9VpqAqiOA7/3SN
iSeAAPIO41tdwuOZ5ocoyOfnrE9W1uY3SU0NHqP7cRn+JK9ESWGo4cf9u9o5EyvEMGXlOgTReDuS
XCAQzjOqiMuxTq1T7a3lUcGO5kRxyjSxXGD0vk8AKUu2EhrytRWc3ql9t3j6ehhL9HeFREkYBRK3
vurUyFvrAQfBuZY5WrSU9H7pkTfIBVAUMCeMvoGM6C05Dwk2oztadDp72N4WnJV8ztO7Fdccz2dl
zwPWK6mu8Mevmr/ajnZ3a3wWNLevRYddyQev+Ldlv6+WmNicaoc/bQFJ2tEizFzFsahtcv5GtKO5
7oqj37BpYfXtcoKoS+xqEcoJcofg8eHePRlVpHktFGnBmcdDQk2Xv4vvJgwWA7BYTpqpAc8vpTF4
2cI/UomriYmSeSc1UhKSb7mRtcFGLGfAQUOHE56Ns2rnZotg1Zz5ff2DHJx2guFFh+vPidugZCzR
ZBBJYLVd/Pa0iIsts6I8cHS+qWwaotuUKMipfQpmbXiFmDHfNWPXVHWcGDn6NsIyYcYJ6BWiPNot
mmvki0EzvfDCeCzrzJCqR6gmdk/h9UR2HsekeNsHWZigl6ARbTnF8r+jDZma1vfUixzWX9Gdb2+n
god/MKL2dRyQidmh71plyPkYpLCvy7bNL+9CIoAuQGksY93gmctqtEtTjXgZuMmZH7wagqL99b9G
LdYdusthMLlxBUeQeQH3aiw0MHlGSuQoyvLM0zW3k2Q5Aipd2ojGXnEisCYJKvmkqhAygS4EUvas
O478iCJxogHin7WL39ejW40V3fKbLV+9ItZBnTJZd8TrO2DK7bYpZ6LzGwW0teolG1qSd9wrqpum
JWoVqj3YbqPZqtk4PFloZXUL6nOpQs1vGxNvx7wKQ6Jq/o64kvjYILJEfYw1bs4nm9XXukr3LM9T
uBwzF70dwntiuxvjJSE57j+IFnw2AS4ypDyw7LjUPe4RfmjMWc4CiSrRatrw6fxRhC1ZYQBCf/Uy
ywdQK7ji2iskhTf3r8LsitOJavVkDJM62nJDqIV7wwepdq21JwuXiMtl3FdK5jrAYYUfRD7AZ4/W
VcJqk65zvVXdPjHQ0wxi/eFV1je5p0G9Wcf5aLp6VUnBvILP6vvQMwWFfWItkx1YNni2nXS5D7RR
V4TjTvEM35CLotLA1sQPy0zSBXMwAJuCduKY5kids9v3voddpGYddzBGKZ27QeLkjtSTVSRsX710
3b1AKEEQ6oMLaacSGLAwN84RUZTrPfLCZ8jmpE8CvttLC4xn13HCeoEkk6DI47tQwBvxmXzJtaNO
KJ82UhIv5RpWYvzSDOdg1Mrh3UdxE55t5TNalE0i6jIBVaGKQwA82oce8W/X/kXULaX9jFVv/o57
YcOfRMWE/UaOQunn1LUoPBydQFJRWIWOv3gr6eU+vkL0+VMBseiEfdBe3ydPH7wKJup/2tf0tW5y
j0EN+coY5kLuU8uMZFotCw1HYz0dI27np+6Cbd33aqzqmer2Fi9Eb/K3N5ZEM/XlbEli1u127qhp
Ba47oZleRjMSbnzM/el/cOinq9D40rNw2zyQ5w+Z0HHWA/Jn7kOfdq2tHBDe2XylmBTqueuzQRn0
21/2qGl7IoRK440Peq4kcgSzNn19PzU9AWP75n32snD1kjO8Z//aZDTdMyKShfgu9EDLGvlgF/oT
OmrldqnNu6fsPYYh/EA3FelI70AKN+/MWFqHYqUR0M1CiMH35L5QSr30l7K3gCBawxpQqocgL1Bb
Nn7Hh4LzKXBLbXDBV78Qz8kDSU41UoMLEN8pECG1I44mxYrhfEbBysX0skOcnJppfmJTNbZeweR0
W8jKmkpnAKL8K7ljkoB4u57V34N9JEqTX7TDfFHPKaSUpjH5nJM1ik9pGnlMCJFyP2lCVH5LSJ4Y
IOIagd4RBD9Gp9mXeFHoZsbKIbc2Rq5+PVLFrC27K0/4gAQObCNL9HAhJfFU/iufehyAHWwubNqH
cFEIzm2ANonfACc+z7iyCUyU9fzEw+Ftn2y7epH0/1xB1mLtA/dkv2IOH2Mm98fF1s2yF7vgwmL5
0jMZUS187CIs/umZRj5BTAsxgzOtoDWwzhHRDPAJitbsEyDKt2VlFR63hAlVtNvfWQSOYoNGTRKI
nXxjgTqogKL9PjxOS9fOKCEPqbd0WhmDYWjCULAm/mXcvrnGO7LrhJwHGtPuug64bq6vcsxKPhyo
EADcm2AiAp4ZCVJiNOV/jfGvPMWIbzIt8HsFDiEpo/b0Nq7vxn+7L1SQkONAE8vUF5dnKrumRIMU
1Zi49t5ck8oLhk38FVaxVvu08h3uyek8wcoNViFg5meDJN8DfVMWh9naG5G7Iy/j2m8K9WTVr2Ib
JmTA7Hx261+QuW5LLLXzLj/HnqdDoMlitOIji3+N0ie7qLzCUYNll5PWfBU6cjmbBH6yT/DLBmm4
v741VolRMcEQjKZ8qsNndWwEk9mq3eMTOeUcnFxrV24miD6eC26EsfPHzGuWTbUDcfPyWDFXcqt+
+an4+LfNgg4iiQaYVZbSCPY7uxB16dyMLO+Gs/cNkRjv5OAQJA4cx8a9QyO3XoirkXhM4bHgByPD
t7Tfd38GH69mRMSqVi4XBjCSR3+jGvkBpudt5T//ZED1vJlDYr3f0a62BpWkYN6e1c1TL4bWS3RC
+iVZcDns2blENd1a49vABbAAG44uf4cwH97jNAhRgeRGPp2wa6wlZ+k1+BnV9gHYPatguA4pezgp
by4MGm27sqZBYheMJY6QHHZA7uN+VHYu3MCL8CUDiBXzXGnehKO6r8xtmW6qXNBinc4rlkUjV87Q
XxuNwf9fvqWHM8LNjfXIJIr47VEDZNEkvUzyGJG+IInsu4qVXngcDMt2ITWeJL11AQ8jc+AJD/XV
04djJnZ9Qszlhtu7RtXIfxqTkCdUDXUHtceZ5phPbxG686Lv1GaMUEAX8hTG6UIUrD3UaPKyGGa2
jB6SyOkRQnKLie+7pFkbzxZOy4xXeSL3pZpJnnUsRimXfvBCeeWFP9PXbHsU9l7TNoK5IXPWjQqV
ftsfeKKVwRozytHEndetlJIEmNui9RFbncgp0SDRgJOvmd8Vor05pYiTDrQVbFUMkRb+7ZPDT/XF
jLZw3kG3u6/XNXU/COUJmEMGgM6m/WLCh+dhnjmxTmTBDFuhcmAl7WfAFkXCdgWDJB4ULE1b8Fib
Q0774AqPjs58EudO1PZZtaBagLWguugEYwDpoHbIuApDwh4k+Ivvn3yNpqU23kbZiM90ObRytIuI
3KIAKy7LX21OyEUrsNSX2jiAfANT7/ZxYDDTaoc6tk8OaknmQpfsvxlZ7n0ho0R39uFIvGU6A54t
i3sPF36Yb1CHsyI0vxiD++RZYG6Cehzlzlxcvic0HBEF5j8x9Iy5mbj52pi1a+RJB1gd5wJzjDnt
zSP1MaId/Jx5PbalJaBvTthJMZSeCvy5jwh3kwOxQohMIggAecLSzAavWBX3YIC6dnADW9RS8k2f
qd/BeOMCEls1nTdJtH3JtIPDeVBQ0MB+zv89QOikdWeaxqALIRA2AMoyRNvqXrnL8z80ADwVS+HY
rhzq+gn9SrbvwYzeMYAph0p40/YeBDjsxo/Z/M1Bn1GgSDjUGF3/kx66NnP13UeUlFiR8x3uJ0JA
ShgD/4vPMGpyTurTZmEnKcDJKCUURM9J45ByEiJccNPHVGCt7VYSCM/lQeCpKLPUk5tfyYidsuSr
mJNq9uyp44Qy9WHtrrSOFxGmMnuWEKnEMGmEszE5oajoMv01ayPCxIN12hjMxFoUoj49bz49GzU1
ixTusQA14OsjpeBva1eKaNBm2bm/Xi7eoJ2p8Hn6rHannYN/AtAGB6kkG/Jrq1EfCcGBKCUgKSjl
eb1OV84c8ETL+z2RCIK+wyn+cs0/XqGZPpO4mvF4J3izfcB+wRfKbQ2MG/gunXTWg0IhSuaGC/Yf
xlAsCXWw33/zLAQa032JG/W5mfvgmO6l+xWQ/N+ppNlMEmveeGhsISEio7Anqn8KETf5EE6LzubA
Yn+QOexbPdB3jvjwUxolk72GPjB+UAHQ5dMAHUchnvKQpirIspJbJc8Y0xIACrdV6TElAEIxLf9I
V1F+2LivCt83B2VNXoW0ZdbuqHeuR543gyzlThHiCWJkrRm61+ven0IWPhb8Tt8bQhfZlEu9yeNh
7zqTvrMx8wSIfVtwjBVUmZrQk1rM4ZDI0cu7fcaaUYUUI5S2oXYE084FdSZghSGFX+/1SQwd6+eB
xbNI+6zSfZIvNvalwfxhk2f55c9Bdcl11kWOgvfObbHUCSu8BI/9Gbh9DVQbiTRtrSQ79GLZ//ES
CX3vqK3CBWhUlbNHs44EgLx5Py4ZAEMj2e1s7CDPM4K8kJVek9LOfP6e++xcYJh6yesFCd/CJBt2
QPdQ0SKX4ORveZqUpRcXz0e7nhAYST8WvNw1gj1+ihCYRJJLogNWNnihag5U3Fj+Vjpg/JOBSAd9
ndA/s41StKyoECw/FxKqVHmRZ8QO+ShtJYg91++Ny0QnBwQAguVYTisaKWskNWn21u/xPzZ6Viq/
hr4ZBreQurr7KYJ11CyEWFwsYNq7PgBpsVidtVUpZvo/cum2jfUG/5IC86zUJdHyBkOADiFRNkaY
TertaYqZ67KEJ6i8fGboUg+Bs6QynRkab30xehSfwjzEOQdMYEJtp4RVnqfkUQnbZhpzRM3w+7Du
apPJIJ+nkJLgBmbeYSTJSP6u8sKMmHFEGOpJuQTO2ybjTDXE2yjN6xbKNiHhZF2Go8sftE5chI5O
tXcj/c9bdcDI1h70EagpHXxyofj10sPL3MtKHsQL8ccjxOzpKWkygkDJ1b2/8BdkvraY1ShA3DDP
oBbRB0TN2Ph+wOvFvBNzTy1zCCQtSlYblzEmUSrkc3mbaV6nqW/tT/tpjaUydnzMoIvbYd+RXSQD
tlgzqTIJT2M0g0PMfGBRCeB60vB0HIUXfPUbbT7HhYUAKV0pp2Fvubh2WYx6RGcythsm9gGUSb0X
Yz9vYg2YBdVKdTUk3E9Ad9sg5Hkl+SLVpOZSjhqFcz75V1a7IUjw1k9VKlM4YVhd3eIHRXsuZpBD
5ujlcQz46p1qyb6PkQx60YMC8JY9let35rjJyscifhizj7KAI8dNFTSd5w1qQvq1Cyzyc/HZM7YL
2yu4n9S/w+1AFD7paMTUpOSWvYTYnTHRFO4MyeJ8jtXmgGldiCykH0XeetojMCru4Y+VopZZ1ZbA
nNwL0lJPAutepW7KFzBQGkmMEu3xQjRahHUV1rZAN0/Vs+WuWjDraMmJwoJNwNekrAZIdk2ZgWyi
aQqF4cw5Sls+fXmXADS8pPLavsXY/1vMNEFo6nDODHou8AhwyJspxdJpNp724Uk6V5j+RWbuPUds
exf80Y2n6Wcnjzbf/3+fxsXU2H1ulVYDM7m5TxyP6cBgTsRnWXUSExHuvOHxkAEeM8HvxbRitKp2
D4vQKjd/CLdkpwi3Gtins6nXmR5QkW3Ort2ghz9fIjnFH/sajoyvMrdqohxF+ltP0NCFRCa1EfyS
T/GzXU9ty70KwEwBPfqNHBk3ve9lwlHry4NZezjw1OUcFS1wGHC1YmU8RU85HTEAedWaPVaAW2+C
lULJ9cPFp6RrTjUGhlLTIk/Wi4xJYXkA9+SoJ5DZJHotGg/9c9f1Jmk53ifhqHmNSdMSJb22Vath
u3rXCGPw7mE1SYwvlLd6brQeLjlpufT2BhG56BAWqg0SOmUjeu7Nxihbtd7vJ3CF60Rnr1DFfyyS
LSQkY2dQDbwKV7B8VIn4BCB2Pbp69/Yx3dOhqPqNELswMrR4qH4RfTP7D/I9p8N9A351c5gAJuKO
z2+uVSsqM1vEt2S7J/sNzTJh/FXQqRKxa70yQ+TV6n/oPHlp4xMaH+hX/ouKtu9hcjvOnO3Avy2M
BWuLpxvZshzOUf4pdp/8IiTZQXdk6cVt/OWtmQFi3WeWtfTjykNNzxUErI/G+KqZPRykHttWNEFu
fGp6gkTPUYl85669jWzwV896uMG7cPoSAEkBk9NUruNXXGPMuAyUSxNci2nmBrwGxATlc5td5O5Q
Pz7cS3xPEX9QQstzTP5F5EwVNfDZPf6/8X094NSc6avv0DY4Qi55mxqa3s4yMuAgGhPxvzJOgJN6
f8yOq80VTsTYAhCAFddeJJ3IePdPRQHmXgYQi+gBXo3XP6NrzJjWgh6+LPMl5ywsksr8rTmH8EYq
jxMjH4LGNS/bqvAQpFZWxSDmQc0MRHIH/uwxVw7jofklY2NdKWrHOF19Um16Z54/PvmUBonYIPak
SOpWBjpqbuerpsjrhcR6c6QFAnvrrkKCIfFXCSX2P2gLcln7xhBrsLSxTolZfGvtzf5bb9lt4jfq
U0syMsc7uPA62lu+n1EnWr66FyFhxx0NX0vmd28aEWIfKdjG8qh63v13P9sAYAnmtUUJ90/uyuSN
Rsvc0ihBZ++y8aBpT5NBSr6HYLiylN3opd3M5UhjYN84kuCfxpGh8jzqSErRdzOadN6nvlgUu7lU
islD+pmtkpgoizfUWhshPubJg+VygCZIUSkvUfL9IN81CKLaFuGrYzKNgG17Y50h7txRilUiHNrP
lz0HxG24Wrwkw1MX9lOdK0PRAcpdq1bpxV5IVVXmDJ+7NeUxmwTIDGgSOZ68N6ugs6S2SbvbW09H
/YjJ1S4WLMlbnPe1diUsfYZCyj/Q43qLg3y+nAdmF+DmoNTLWmU180v0drgJRgim68WizDPWZu6D
8tPh+0obhesMx0VIKTj6GbkxNYM6YdQI1ezFFj4yWtOJmoeLUWXKGRQVMcBXSk6ZxdhEp1mz4RZO
MBoitGamwnx+r5QBo80RRmtt44EPb+X/7Mtt8STpbonIeIrRoQctPtUjNiMFPi1KeWuNwrKJWbOb
/CqBIauCowHlkZ+MSvygDXOwfJF2TyPlbxnzoOReO2fb+57SvHiFXPsQP7f58yMLA1n1radzGMLE
O1mKhwv1oAsGpkKHxqXKMWv5oVd3McPytGGcOZjCdXX3HFxOFMYRgdR/7DstS1oX3J1JldWWpyf3
V9AO+vnChQZ00Nyt/vA8Y5tf4/wW0Ss98vNAJ8xcVYIOHCY4JrU0w6m69kLgqWXbp1IyGwn9lUTs
U5Lh1TdixhqpU3cCcHdyB2KTaCAY6LorLzCzKyp14aLiZJ/0mN4H9EfNH2XxZtHZNpI16lJhbVRk
OCoiAVd21ZTE52SGrpSmFNmdGFtVH7WtDvkU27vyYXMiZslKXRv2dsnVSF8ssDHV1hYZA2ID+J1W
PL7+43pRh9+vLe6K40wX+Co+KSxmV30JDKN6lj8F7kGsC9ooJkE1oy6TnibzhwU7pzyoctQjPcCb
aOfStCZpywzFxRhtTJk5imDNW0kn5hNnvFvS3NEyuO0Hp44GoXNnIIz+Hjw737rRa74HsH/U2uyT
UAM+CM59ig/LO3OIESoqhFHsBuJKnj3jvAYz9f2uRxKgKbxEvpddt7aDrimkZSrKlAKmJvyHhvpu
vvpiOU7+DsHIlMT62sg1jQGBFnpC1JuCvfUdhq3fzv7d81LrQH9c0FUpSy3r3MIA+8D/0jy9wuUt
bf4peDzX2R/dfHAbu0+AusRolUTFm5OOokiMCI9IAmyWFEz+GWrMVC0ofKpi1/kJKL8q5ndUmXxb
SddsgQ/BffnI1QEKM0t3zfbKjBBbgHenk75c1hWaXbZlfxhZeUPQcxVS0sNyPrSA9DiALFE9qCjD
rq8WBNpx6c6AkgZsXG00Dj71Ng+uKX216fkEXzDtYj0n/bK6jY/6Fx2DMzsCoMyJDhsE+MD1yoMO
KXJDdkkrwe134neSGN5d6lonKauYLHKiY/6m2B+Qj+v3TmJvqv6urT6SC2qqCHpE0q9DUzN9Nx93
cwQkMFYLY5BYKX6w361PpU2axU8ueCsmT+6an2O2obsugIe3L9/zTmo6M/LIvagYov8VaXHq2pwf
0jd0ExG4umsUIAAq3T5nxfgk25cAXPz+LR9qQSv9X58wYrGzmUv2CxjcttrA2yhSSsvn6Xr3Z3+H
vmy5b1ocvg6UD+++HziGUKo4CdoTiJ7q9STdPFDRU+955iQnUsElyhDVwRuFhW3UDFQHnoEyeo9e
sg4TV10M2BDsDfkbmhOeLP8MkU1zl/cXo7QQ2GsuikfC3EWEKkGrGNUbGzlcqDoby+xE7PaD6Qm/
c4Txt2AOr9q1KZlIwkPuw8s+pbQvWIVoRYoS0c5uzwJ93CuWCezSPL8miMtXH4jVQZICvQarb84z
8omNdGh8ZlNa3FDr4lmDu+6f3GgSOxtpcXe+SsWmkpsXaBStv6q3yontfrj5eP0dTZ0fVnEbR0d3
NIaIFq7f0BX3gmEtJ5QwJHrTAyzymM0rdLuz3IScSCpBwAszSZSS2FWB9LWOiL7MfJUq9tIjTueh
DQ+/eDixGK4xzCq7+iAARgGlSfBApUT+bFRxeNY7vBNLRKwHzF20odaSJ3119CqvSjQSaDgnFYJ8
nRfzOMjh2Fey8bmdVCPro5YoqPPehuIOozCWwADzotEdEGqgWUAG2PPrbQr9eY4qG1AD6TqWinLJ
E2LyMYDasedZuJYxzEMxM13t5C6MI2DLZrGq7r4m/o7XI+7ZbfFkkEZD7x1LqAXKzdeRGOBt+xpY
Wlwcb3b07VwZ71kSeiAfJHmHfqG/akRvTGIvamPMNUqZt+kRxMUx682DqzEXQxTUzbUHxD3Pe7VY
+yQM6ZFol3p0ZKgPn7YC3zB61+o+kX7zAd23Mu4ZaUApo7brEwfLDgXjDmxNQwDXF0ribfHgf05+
iT3YCfKZEnWWYFEbT9eJ3cIjmMt1Gj0c4RcCALsIY9uxTf5R/DoL2EhSeKKni4I247X2/DNEjjDR
jWK+moWPlLc36yvoGx5/pG4Xmx5lJ733KH1CrkJ0W04f9Vz0Dpui7A142ebhDpErXuMJ7luQSuqV
4ze9F5YTH0ZCDgflhPRTOdJOfN4ndURLUH/oQL6zyykEGlqGJAQOkN7ZcEMDPCyCSectUxBh7QiR
xk7j4wjXgiUOthk4s5ZobbfRrRaL1r8pV8Ku+bt9phbV5kDE1HVlP3In9Xcz4Ta1ZLcTO3vcbRZQ
KcXKC9LbBnvNh1C1taDP9/XsyqkdG27uyC0as3nkF+lQ0Q5lF+tMwKsfOHr94xY3Juj8IQGR86v/
6eOKRzgKmUayk5YprlhWpUWsUMUCg5xX+fgrj9UXqKQpDNXyiz2Y38ejMR91aVtDwcO5rzf6HJD7
pU3FPNshNN2U8yVHrO53fg3BElXgDSygxBZxugSi8PzWsRWeDucSv6HKrYjMmaH6Iq+Hq0Re2Yj2
XKZHT37ET3xyMSkh/OPKJySpn9/r2m1ardR809afFsowad1Lp/pRUgB0/SjYcnl+HaH5pmM/UgLq
/O0qox0rS+Zzxw49dj4lQwexzwH/BgN8JLZ40+jnIyVBTWrx0JIjyUpgPJ2mfdJEuWUhBs43D3dr
VcU0R/v0hms+EVhr7M0PLDnxXfIvJPB8lnO9wcH99CLT/jSDmulpZ68s6fQA65qkt03e1S/QdeN2
glYwbwDyImxsGtsRBsi5YGc8KxbYYklCkM+wagPZ5ubCw58vaJEaxMJqhDDXFPigh2SItb5UOp5t
zjxYVBShjSoxOmYTV3O69wttaZV63NnRKd57B9B551hZl0nXkKdCKNQvkXV88d9bAsU8D1cW0d4G
GS7vxnF3B4366uO5mIiYAsZNDzs6UJ6PT42wlVUQ17IYEMWZI6YlqFzSjcWrhM3S+Qxy0oyP9Pyk
E+2fcTnA3sX0UOW1ct3Jn8UPNRx9JlGjAi0vPRyVbmSSTq9A3tIDZtW5WxMy/QicD26xtBf/Xrgv
Pu2F3QJeWb4fRlvB/yMtgT0o5qX9lHC4cHqxqyjb9nJkWoulGcLr71ArdchreExbOvEnGJYFpfPc
AkwY5x5BabYbY3+q7yzuqgfBfuo6lP8ekNbDTlM/7G4Ol7+16yOINcmD+wtT4z7ikr+kyCpwDYba
qUtSYd2tVWJcXpxAsVXcNEsiN8DgRxplkh9wF5+r7VKfz1PuxYSAno13fHw7PkdBC/rl4uL8GaUu
AfLhXjNqgqdOPPOXFXQHbG9783lh5kBdpnywV8CFWLvRkYGhjm/jnJ4a4n/JQIMEg8sUBEplwYvm
TGcIXUS82Frdd1HaaVUu9s3arvk7mzGin0bUWSE4GsAv0sT2LDj/VKPh7bl8b20LfUTq4Y4bIa77
jCyll+WBF4Yg18fLwOS5secNqQbhEwp8uFexlxqSF/Hr71PL9Uq2PIDqv4InsZ3zaPw9z9VbDd5v
Qa4sCoe9Qsy/NIIxZfIPnc78t4Z+zL+am+hzOhCU/S8q0bgRTT/GZF7WcrLk4sCBGIG6+wxYwaSN
C8IVs9yJQ6eB3uALaAI2JjQVKSXP99KYiorgUN9Wt33iYDpolGeaJTeVJW/jrB1z3iMwt4tZgr+/
qq4amHQ74Gshe4gv620BWqDNEikLFzKYIdm4uVdqbsE6bhc+eP27cGBmoLKxcEpzlT4J23NcoTSq
vk+lVSj1GCV7LImBeIIN89ETZRe6jeEWsJigZAjtQt+gkKUSKax7nSK18fDO69Jrq7CUimCnJ8N4
TD13tLtlr6X4sgFYLYi/6jKYHRAW8Yzw9xHlE7uzjWQhkToxf6bbOD2jDcFdhADdHo5x+P63s1Tp
lCWPdCzv7rI8rmb9UDyPBQ5gG4XZos9IPeIjrOXFX8bXkhyRZzUgFqaPqPWstbUCdjn7v9PH6wmN
gPw5up/GMQjJZDuf0W7L94xxjm1vgQY5WkEMXGRw4z3cWpPda5rySxsy54azDXVOSpkIR2QiJoSF
p8F08oBIQx3x2gNt7gUvlydzPNhbA6GKaTGR55VvCZv7NQllooDMM+JcgxiRIrTEFZvGQWpTokjK
ZHSeFMWenPaVmzNigZANzbGekAeSypHAmwIN+3RpUnI7KAHZN9mtubZLMRxUmnfAL3v2PUtTBrM6
SwDlYGBL8N7WT9vmqGvVaCTrGFpYGt0vyBg2GO62H14kXO5Dy+sOypGgBjh964hS8mWr6MqZXXc0
/BdoYEnFN2mO3pxn8/7Ey+I5DB1m99USltUDoFzN9UHPZLEEVGFvFop5EMKI1CywHGmfESgyGDz+
62NuBM9VWv5XfoBd4w1e0pvcKjWwmT9xJAP3iZIhqJgFOhmkOkSpF3oNrEXdZFvxcwXfKhypPtL3
iAx/ox3iAw20C9t1gDR5KKDB8xpytWXZ0Nk/j5GEWMQxkbGyMo1uotThtOS9uWDvNxd3XgAeQvfm
DVN0hx9ZyF+LIDm+fRKMAYPJYxSO37oUS5rEhY6vc0cNGHKIR8BgWAt229t01I1uj4cw4ch5DgVo
HjjMNfghkGnkIIagpbALXHrsP+cRIS6t82Pgnx3PF06NMt2NiPtJcYnikVJPNugz327MHS4fNz0Y
iJseIio4cuEoPSprWC35LDBBe75R1UlMDK4JW+VDtn7+SqQ6ntCD1RO0ILJQB7cq1knv74HMwehg
XQcoH+ihCHCUoZPZ6TmSXD6XGwHqU7/kncU0G+CCDQeVS84dJT494rEqUk80nbAmbbV3Kz7h+iPm
In56xHOklYxiR/Q+6245lz8iG5AgwrMK050vcU3nkmXJJMVldWiSAcEkapnp2mCeYuutofp71/Du
l+Kb+WZD7DxNF8ifD/u9GosWIl8u4zV8uD6/P/UbM79l8vXXDSKhKkU4GJen6DfHy/anCa6b1Ee8
eE8yg5JcTfHYcO6ygEFKrmzbV2RL7z7aGUlt75hMCRuk+z9jeuTg0/fgaadKqc+PM1jtsyIhb0M2
WT6+F13owYnj0Kwmwo0U/uhDGaKE+lTr2RsZ28TX1Znfeh2fYevUUJvdBEotCVtcHYAHldLkuHXZ
/dcWmHnqExO1+5xRKT78Rrp/pK+NxLkFVzbBTCKy+xbrIv0iNBEOGtA9TIKZ4enNMIOFql+/ygcA
xgN1HAxXs9JCdvqYu2C54RKfiKGyzaamW0TT+TkJtgWKROrEA4i9rz6OtrclE1g9l3r66eS17nUR
D3qLAXvr5bL2IG73EwWlzCvbcFejcPmHs0Yk+DKvVYAsVSECjBdxgU/sqYTbdQidhW+tCsn1fATp
+nGIUW9oEIufUZh/W9v3uXM5qyrgxqI80FS+xKDeP9GgMx+bPaI8KT2x6oNkuYC2LKU8g0qiMazE
vjO4Qh4GDhYq9EpSSmKf+CLxtZ49ypjWgK2dmNnJOTS3zaluxfBYSuMhfF8g8hoDEY6CFLmU/4S8
V6LcrYCttF0PluSTSJoeKHdWMPYCdXLoU9+ZsuQ0IeArO5E96P4+k/17HIHfKVDMXeEA1BgYsGPp
E0oupogBdAZlIazE1SRGlzBtPZWHfKtCKp70xupDGGMt7myqmvtsac+HcAxwPKeqKPc7ajwpamDT
lz3+w/i6UmxCJFfP/BQjMlrDzwRWgSqMW0OlwEeCqRsfb86kt7XZxPdpPvQZ/hf2jFUge7jiC52q
l3hpc8P9coLn8ve1rECXGpofZcM961O1Y6LbAfgpCwzaVs8ZDaL/zIjso7sNED43YeYnRwDO49Gf
A4G8rBjqyklpTyf/FnqWtjVkI4xopX51qEo4QSQfLlmqtxjA8R0SyrguTQ1j5mmCgiMekzfaVOtd
jhqkIKnnZkiGQ07LCOG6s+5EfM8fQnuC6cwghADkK402TQAvACs+DJvPN1wintmXwQZMtYKfgcqQ
dP53JwSmur3xxzUWs2jTGn4IJWs4m+H/cGRH3ygQ5LgoLnTF5Y7jMzN75LP3Yfhw3zGggFF/euJl
LCnaz9JlPLRlvpfZf/bTowRvyjlFkoeyrr6WFdCJT7+82TR/v/MU+nsdk/ViLIkerhFC1xfQSvp4
yWCyWHbc9/pujVMpDYTiTxyBIzRe1uEMUoe4l0YsMnUJhgVYvRPkWShN5OoEphoFn356sALQxhlo
pDNY+4Jv/LtpIPDuHPio+OlNAEEoj+aPIuJcx8sK/AAwzNWvXkPJeXbdlLKjysiOlQQK2ViZ1drd
lDP3TTkdIlIBrxqvkV2PjwHMBhb1yY86+wsFFnLzGCKF1K2cA8H9V1f2b8EQcSUyqHaYC6c4H9xE
rTrJ40EdNTcjSQaRSRSliZMqC1XK5rB5Ut+ALaYUy10Z8nYBrKJUB4en5jc2ItyGi7gfxxehuuhN
t7t9dFQaTjIG+Jd/6Lf7LLmcOX1EgBcASwm77JrkYTwFJSaaBo98CuTL0/hPpWDwrZqIXcHq2phw
wXOuT+vP+ayPAHBiiHq3Jwd7fJznfRa6Qn2F/XUVj69ZyML2VRNuWS9iZAsSZ6vNcTRN2kk9UNoN
lK4daiMphg0gEeZFXzMFXnUaTDiR0YmY5P5Cn3srQkWfXMefd5RdeosOVDOmy/m3HRpGV2gUbLGV
IQoAutYV+ABeovB5qNM3TEfzFoSmX6puDnnrmOeRJRjdmvMkEmipAn+cXkPZd1C8sTb69HUUf8Et
CcDJRchfoo+BEL4EYYunJAbIF/Jvm3Nyxg+fMV4NBnjaYzTHJlGJT3hWB2TKBirVa9u9ROB8Raz3
uUaa8R/y5asjdM/BjcMhVSwEVnLRcl09Nc+BKfMhhhYk5Q8mumDtYEqlFJiHgB0uvaKbEkFI33Za
rmvD+kk+XcNeA2mDQYQV0v8YnfMFLf3ikJY16NP7L7ph40lJglfDMFw1UzXiufCACN3ztW14DwNb
Qdgmoz5rh3kV1bJlGaiQBKHtMvbtcjHrDggYOEO1NVmD6vTQtFc1UsinTt+P1zjJFokCS0ejtJFb
CuQS+S6QtUNiakzCAY0bWtoS15PtUbkY+zwkXzxmw8ODWAwXSFevQ4fU6Oi8btv3vAVVv26KjEJH
D7MlEJq2inHAkOvpQABD+smh2q2Vb0eoZqyQXWz/cB1jHgJjnQmokiCemsLvaVzS8QbINDuZ9fSg
wIEDoJ+07SWRroX8q4SGbv1okfuy+KYo+kt6bErk1j1XRQZtB21GGHExoSEjsf3t/0rkXDuRVXyq
rZxMPFv6Lh6CWz4RbeG4pzZbNTewQWuJyPhIG2vHTBrapaCjm+jEUwcvKKEEGNY7rGnyYXWJIlVK
t3RcaNr3BLxvh97U8HdR2sjx0G02IxZYticyWjob/KYriK1Oc+wW3jFTLEgFyE92iPNIJrYqpD7A
X4EMybBKc/rXpGiMeL4LbRyXoQZvjRVxj3OHaBrTKhvC1yW6NMpGd8rdbIDgODv8BvFCae3rqW1J
lwh3NHzR49DT1qKioDt1spOfWAaQ88397skzJRogFyjHwJTsMoaoQYFc1DiC0XfYvD3BuOz/lLvP
yd+UWWTKYG3lXh4XI2Cx7f1XsVQ/QFPdKNdose9j03PThfJak5V/waeGA4YpV8hS8QXcGns6sBNd
+ptgkP5yjp20Y6i6vLGwWP3kdy+vuzhrKp6QiPd9A0NA/+B9dL4Igr6e1UM3qcaFJdEOPr8Vtwje
xxA81guKnUoqXVpaqUSAj6LT4CZTZllgYpr2q5TJZxA58sFC5UmK8EzWTeQUUcXFvPF4KgnuJ3PF
Lm2FpedW3Gqa5rCuIqAa++e25NC81TVzKUO6AYTdZ71xDQ8I7lVnfWm1bnIeaKySTmxxx5gdDBst
eZEmTLbvSHcuJD+CAm+23jsrQW9d3ow63GZZoP/EsLegbxKZFDVHWscoHdRNVikInhpJYdQjIzmm
Mh2+CgVRis7lCBDj0QjCsdTbaaoYFe434gjmq1WAdpAZETMi5Rp/phgMxV7NTMtaipYIxPhiXxW5
FxctJ/KjcmZdmaupe/Bo0tQ9r8wXXnwNlVucI1Dy98B5/hx8WAYZ1Ux2CatyIXkZyeOOZL8V35RV
9yXOoQ2E59/DHMBMkYKi7DB6llPod2cVmJmz26OrLMI6phvTUXvcZYo+RnTrZXyGKdNrygsiOLzL
wtMivoJ3aTxcSQl1NxrJlNzvFsxYAcqdIDRCGK7ShDzzBWQ6qzI+KtgxItsK3d4EvVI4shVFp6qN
NsYBfb2jR+k3mM20a3hauP2lV3QeXvYzl0S7C8Nb/7t0YW872VdHc+TSA06ftRdaQagnXfx1MymK
zwHQU6Op887MV0qXrkLyQcXh+0wOv/rsGm/XBmiuaXcgLoyFGFBpLJld22/ThgM98IPsBhYBkQKb
SOYafcPHSyOo0rIDBm6VcCBvCmSJ9AfGnysxh/+qxNjczkEgYesUh5A0pQGyQoptA0iUItnCzGDw
1jnV6+J70zbISo3ovExkM6fNbFwD/nXlf4tMUlXiBLDJvWWqlF5vhy2pUbomCL6aaRdm2Gl+L9ZI
GXR2JNn4kZ4Os9INBe9SEby5JHUhDTEZxqjXw4zVJfH3rztJpNWEQRrY1W2dfERzi5JTu9ebya1n
sU0f8viJbz+qzNucPpoeaRC2C3aKgnGOW1ud2EYY+PIo771OGQJ9Zo6ttsycwym0EX0FT+iuzcrr
hQY8MpfLbPhGimnTGgxOEypd4z3+lDm/gEWV3rVODajleLsPu1hp7ziv8k0SDpe3iQMoG7ShobJf
FVNx2K2hpwCSTYChQ3oKibwCKxo4UynA0K6fWnydqeYss2mlyXomApN6kpVJp+jQOF/v06XcKD4c
sUg7QjclhM1QNINdGRO+1/RPRI9JLZ9R/Wu5ljT4s7zVfFRIyiPIO4+q/Us24223cX4bm5OHHbE1
DPfSk/rCwsNKwmrWruKDIS5mEmKCq+2T8ncK8mZhzTmyVZejCfhfoAKtXTshm3EbFWoJYvLXsP8K
/w9WUX6wRT2g2uWUpZUBxntdaZwJYLbOiJJZEy7S9WAiERhvSwz9+BwhuYYUfmRRMwcYe8SCz2lE
W2JwulPtReu6N2KLFBDN/7nyE/+rDfVZanmGVkIrkEUwZjHrdq0XhXRhXDpCHvK9Ma1SLNccueOk
ruSIKHEsCQgwrNpUv2up6rKIwnbTJT2jB7917Qiuvk5hhj885JpVUODXDseni8QY88WdpnmfvC0X
cCHV3Xa91s/k5g/JcUydz9VUQLL1aAkmoyiZa68pdMF909/7y/dVzTabGiHYt4t3ZlDG71V5mRqi
zMPRZ0mJFzEfPofLaxRZdY5LwOprBoAL1l1DPkPPdXXvN1V2oR8jAxLN9fNA1uEs0qeJSMP/6HwK
aRAYnzowaN13xDfMQH1UQ93vvTRc7d+IzBSBxY7Ljd1SNgAnO0o5lESHr01Oh0sN7WCLe7TOpQmf
aa/0NUKQi9tZrlWDmMWXlU0pXBIDc867YqyZ80aOzRwscS2QBLn//9QnPl2kYmYrIqW/MLt2KP++
x9ixK/JwIQmHCfyWLIAmlBIOq3D2Bovq3SsFrvl9q8j5cM6+ONwakMH66ueos82LgzUbhWnJ9URQ
3AKQ5RQknz8psF/pe86CVYbfej0E7Dn3jIz47E66lj2pKtElrdvd4iNGbjuWo5O3jxNGwGr9yCGP
Mza8JDkj1T+jMq3FUvmqqmc0bm3WvwkD48pUUpu8S/9bQhq68kx/J6yD9NW8NsqEPSpxt1cLwQmm
SOOrowd3U3DMsB8Yw81y96QnZxkBssaPf2GzCGBTbC4s51Zlhdgj+PUp+n0Z/e9M/gcdfkDAd39N
qSSn4EFn9FSBZYOM0Xs3UkPKlJ30gsj4s6Mtzrk8RohuWt98SPkEIMxnMZpZQwYtkl5Hhn5DN+8J
3BZWqybrudlg0VEv1/I9s5VXbRMav26yAq5RrNX+ah/ENrWqE0jfnNseB+vleeNnC9fPB/Mk3r7N
6Lml+avhUj3OqUqu7ttjoEVG0+uIWQLlndpDYHSYXQZclBSl23yrQZC5YQzaJO+1lCnQ7fGkUPn4
bbS/LoV4bXx0ldxAIgWfCTchI+Mzse9X4P3J2l8ul3kw+D6aWrWu0CDkCp75fBIsHQ+y8u4RMVgm
dHinY+6O4yl2+dQOYm3s8HFD8nJ9o0y9uQQIojs8xygB/bZsvB1S4ODBHHIvvW2D6iLYdWnu668+
Z0VZPSHSNpOh/Xn8rN/FmdPj2CUDasyw3zWdcrSPxiLobz6Lifr8Bh6xdTCXCnD3fPcCeYl8pLzb
2K2Nzm1+ueI6O/r8w6f/78Vslrb37pi5mJeGzcTinieoBwm1/kFCNNYY65CFq75iFBLP1LWOzEQw
vbbyBdC8F4mXPvR2soNH2aDgPQVCH1iz6klWNDDZVYzWAD6Q2hirzjAj3NfArXWkhXP8txtvooMh
BC3hKnUm76JXnO1wsb42gfvt0/9TLPSqEHdUiDrtlEj2ZJ8iLqQZOS+b30Ou03tJgZe7YStw6Xuw
6ypBvwOQSBQ3qYA3+I5GKS2Q14I5G3k3dWqkWjdRgyC1Jcy6HrhqdXORYIr84c1nDJNb6jLYytvx
mg7qZvUlJYT28JPVMMul694aeMBVcbDw9phuOxnPol95/v6WEE+W50pbTxQUC4dOv8D8Z7jArUVI
pO/LBNZh6LX6McKuHrV+ewKX8b8UwGGqMMsEq0A8giXKtXE+SkLXWDgmAS1yQjXNQ873xLTzpfHl
Bs7w/synjOZJ5rDqVWHi+MRsQ22TN0zev1GoYubk71Y5tFjpi8A8z1GH7cBgXzY6gWu0+Z91lBnh
MbGlqx/qgw/JAGAIXkxOTBnDFxfC86RVAZEWQDA3BELZvml2R+Tbcq7v6Q3DhqfGnotUDZga/6Rf
/2YLv1V39rvSA7CbkApFXEMhYICnyruEMJr6OFP5ov9L0Ru68allL5zpZb75fDCIQsMXQ4oINBuB
HLI7TLoO+QyrHL7FICnD3qSPWEhTO+uBOKWtsLlWfa3voANg/yR/nje1XB8dENRFUWert6Bkyt5Q
vrknK7DX1DsCg8yICahW3iv098f6AitO+ZKNmCIU0vtjdiO0r2yViK+i4sALiZUC5WPCxHjPzS+U
xkbCFHiSaMgPJPXq0f0XVyBuj+1j/rkCRLjCbk02YpoptDKe3AT2nyA66sWnPAk9QYCsdF8mE4Xl
6h+QH9AE3/oBLFcdX2qtgJGz6V60EB9ZjF/xP8TrNH+RJHGdzbUmOzB/3BIpZCnlQeS77339b0ea
vE0vAau7un/W6JdH250qXBnE8cju2ayBZPAi6UeB9AmUtdxkTNX4j8SHfV98CYjx0d8w5FNtdQw/
9q4bKBozanzlANh8RQfyYcZ3iu8ofEHt/a3cU9oXknmP3YDejInQf4ybK0A0qS6/AgOMzqlANv1w
GzdY0SFOD8gf2yE6cOEDbBe25OthQz8SYio9F/4+f/WzjKIkDrt89ftmATAvLbUXMXkEpl4KNgds
aJCz3yb3Zfp1wIS59HrZDTVCNji4bsldUQEr4gn2RzaxIR14JEbT7Ke4FwCKFIXLLmlGWtbNjxID
DREQbkyGSfOlHuetj6WsJxD7M891aR1E08TqKe4GqiLr42rQepq+6FEXXxBsp1oV3tbCAt3G946S
tsl05M+mIVS6RD7Td06FRQSQ3Ak0hP19FnDY+8/rHCtygDzRiumEMXKDjbYedxu32VCqktbshSlL
g5nBY+DPxXWYKVxBfSsUr+SsEIscZZ5pXdKSslKLFffiXgfrUb2L3zKJOiFxkOXWZQCRGw1T7RjJ
mYQzlDfrJ+Hw7xdkSmFuO6w8dlwmVcpxVIaJZz2plGomb4ZZSMGVI5e0s7bV0Zt5OZRaz0po/afE
b/vpxPYwBnF2A/ao8rf9lhGd6q0MhZIgH1uxfqmvO5zxLQ9pRhIy2qKCISiC8E0ZWDBtZEL/EhvX
H4Lj0D4yiuRSL0aO9b8uurUMHZpJ9G0e6cFUPH/tOJnQltdtq0z9Sk7t+24rn7HiHBvK4pkTpRv+
u0LGhPnb5q3GFZ3B0w/+EtL9Zg3QUvKTQwINErH1L0yzSeLxNihlxj8TpGIORrnNpxo5BBQOqJWy
bDlJ2/C8ED3qq18WBYfp3qQxXW/FE/T1fAw4U6LQjQl0fOreLfHWr5W6jRS/cfAMs3I+1vqyx5+a
iJJTmQDax7Ydr5ApwgaHqK3c7W53Ud2Hq0fh2DeXx2YnLnrZ0G0l0qKsPNlHFkmO7r4JzluotkbY
pNhVLtIlGQVVIreg/wQEEafp302ZWCJFv8JGKZPRs7LT6UmPutli/WSPRNivOTDFo9+xH6jlWEVE
aAfuWCXx5TIZJyKYdepZfRLuBIMxt5Duw2LBL03hh6SNzXjjgl1iEd+oxi7O6KpIGfpj0EMCfOtS
9CUvWiko7fiXkR7WUsfBwyjGggu6034g4JsZFQnFjAcxajC1esbTYlEe33AEx+/lfn0sAP5Bc9XG
AmYMN/BPp40Iv9nzBRwnqfGWZFsU7m71gzfJw+1BlyKAd5QxSXAyvcH4UadZQVQoYKEevooUc16B
zCIw6Ps56uTLCzctYMW7WHkS4Lz0uWsmzY2761R3KQ3G8HOG+e9bIRIvcspGfW1RZaryLix9PcyF
EpBbMCK0kI0AJmGL+jSkKDPf/dd/jO9zGBDLjTZVoadbI8HW6TWvzc2IRukwPJxs7+XJHzxutmL9
xYMfEXSTrDjov6WuOdAy5/f+0z42j6Dy/ImbjUypswLmyWiL18CUhB9UO02y2xgp+aYJsppyjrcz
whFe41WfkAXfmvoH0x7/jaaAdfcSRRlOfgkOtUwzgZHwKG49d8eTZUUCEJV1UYXS+8w1VhncYOP0
UQ7Eo5I2k7Izu+Un+p9tx7zk+onbryG5xDAkommfQqnY3gqkdt7yvd/YU3DeR5eD/W59ad8+ViVo
ge5K1L8AoQpCvh4PZiO7RyWogFfgV+VKOeMOXWCKK9N7LtTkbuWWgQokbjW36BZbh1G9OpIMB1ED
hUTxLvEh5T4gWU169GTh2W+aGLXKetKkog58gHJpr4maEwxZbJml3muhyshvdC97/7iPoArS7xSa
gb8kLtwEVi/hoOwvIYUHLfE9eW+wDn+CX/wL8WDT2xgPcGd79cF46aK8uAWaPwcsIrumEDpUZLFi
m2KXziTQM83+G4kxC/88ve/MGRjZbsllhtIl6aJk1lsh7ismGE73UrYSaMXqGbz7AHAN7lgCmo0d
4JbkUzRoSLMTjTH4eWtXrmBKUsv1RN5hHQbdRZJSg5G6TS1JbHRp0lN7MPzycqtR/B3trE0jkjms
dLqa7WCZ7i6ogP26T+3NYYQYiCBjqgP0NqP8ONlPd7fOioyRG1FXVCLynYDqbmU4OYJC4nqNg/xW
QhGq3d5eOKa7zACUNhfEfzzqTh5BAuvseUFG7gFkoYbrd/NXn9liosG5OaQSDRfRhERdpKs1amyw
qWtJb0LjJ0hvLNnQAaKj2IZtZJYN/Pk/PBA2ZSCVrtAdQ+VidZB0LID3zdrQlSGoToASYltfTSqA
Sukjygzk83/tZE6s0XqadppZpqmHdWS3HtaxhPXDV2fBnlaCUWgwjEjNRCJIe4s4WSnelua7vxJp
Mo5sTsIQueYxZI548N/xdqyBGv8i2BPiygzgl26xMN3MjOejWFX6AqhcfOIfPdcds3wcHGLOca3O
3QwCniJFfZpgqdmbYVolBrYj83Nr6MJTL1pAmsj7z01Ufy2hqMq2Nm7kketHvVqjuzkeI96MSjUU
DkmOu+MqwKMD/EEBUQtp10JGPb0BbLEjtUVwyv4CgcpVjmTUc44litoykqkfn/LVrQhRdMZpqbui
bFEyxk4NNY07/sK6FNMF840im/MBmfjdaeJJBcSnDYg9Zgej5DF8p9IvJJoTMIGExS9F4b8/pgAX
GNdd/GfIfkg9nWSUiDGDyVBkEkIWw+dy+bOe3aPZUmo3mISLXp4MMrYJT0NNkH1pC71vatG/V0El
oJXBhZqkNMzOLU3AEPD0uWWCJiOBn2JeaSSgdBUWZDtY8UgTQagVmvLkv8ngB4ShhPjYNNEVeWKu
Wen4p3Y6FsSHdvP+I52XUi5HOXXCkqJt4QRVv4bKkBLCFQ5SxuIikEJD/ceFvhqSrGs/hU+Nwq6D
Df3A/WwikdZPfO7qBIjwkq3EOC2Ei5WIDeggSXoVKl7c56aGGQay6rBy6gpA/rYBKiI929m5dns6
IOv88hchn6dPBwDGObPwmd0vNFfOntIqIZi7V4p8cx0WZNV6Ef6f6Sk2DAUrglhN1IwXLx3npQhd
xMoTU4uzmdAJDAvIGMGjW+wVK3nVJfGUq2ZfWeWekr2fqPy0y85DaSwrB7RacUfxh5KTpZWHnK0Y
hisK5eZXutt7OVaQ9UwyVa1NON8C1uxzjmGXiFLvY5E2GDMCDuaTskpHJe3dwG/7KqAch+mCx5LA
Nh6NlGxLqVIiTy5NtuyTnv03hcyHMqirrzXd8we0wwyOnumikWgV09EVf3z42FPtHOTgcMn7PMuQ
lBgqF1TAGEc/BNW03p75wH+3brS/CzAaUEMCDlGW+tfSxStNcc9SQmQAmQ1ZRLJieAVucq57evVm
czh08sYxfgKvNjSLlSAw1zZvHhoSnrTHDxc/pcL6qJdiQGOvkTvIZlO38QvFXPoNaup5/XWadUlT
QsljNlFdm31c+hDmYXt9aHOnQVkqo+fDIztZjVvWvzqSDTeGA/C81NpUccMpruevOLbD5Y2Fay0l
XSEMU576w0NfbkXOITexo5UExoMyjGmA6PQaPePc+w6WFrU5m9Sl8afnEVltR3SWezUrKun2dAhI
CesMyjcZWSO5ebDDN/rQzWdr6yxFlaNLrIrAVnhLPZxfkAQF5OmIQQhmqCCowPaYRvEd7jbsBpdZ
HmEQhywObMowyk8THoDboGSv5DU3D3RSYbQkosbsxGsBz/emfxDXFYJKkgpHvORHt/d/KAtFfuNh
Kgx13oOKLwAPymFbrBOeB5plvEDZwizhK3t++x+wYKcAt1NLBWMCH0RTyY+/TmPH59BVKWy3j3X7
svAkYDFz12PVfXIoMF9CfNhQIxgbyuysdRJTd/XQfCMYHSnCWFTAph7twBZMcIQTg/Rx589PDske
btIDeCav9IUyjl3o1+DMqTAGzwyFaCtkByTAnudQB5sLKmFaJ3ehfOx+n3awZY/xLPduLvqaYHmp
UBTtVZA4Ez42akUsJPo/5zROJE3fJgkXePn8a6ANnoVFAviuSgsUXRmyreRaJw2qG7/aJttWg2ly
u1VNueMEk0wjhRIwvmvZK1LFsl2xdaZuQ+TL7S2mxMw+39aSHd18r51sRUxjNiTGXIJo3CuYapQ4
0eEPonEEPw8OMc+sF3VjUm5Ml+mKJtAra839bUe0HWU4qBNomoQWZfFkhf/8de07YqaIy7/1akTN
wJvY+U88qKURYQr9apcX0eNPbHe5pUQYLNMvfy822CvKGBFzOxbikJZZHiAJErzyO3zXeRnNKJXw
tonQTG2geXxhmDgYd6DHPkDgoHHtTJuAUixVoqzCqXvQp6Tu9UAYs1rEXARzusCB7M46Aw7LbqGo
minGY3XC7Mk7aEglY/ECxsq2sCAbnebDozd2/cFn4MAVJi6B/ZrAls3AcGBvLLKvj71M/OmkWXLm
Owh4EQ8Upe+71T70aIge5hjyyuMQhXwdC9g2RtPD9lXyNa+iEuISkq5LSWwjHEzxvhkzzFTADna2
lSxuvk8SrCokyG5MgPgm0tiQDA5shJeaVpPcngI00Jav+XCnsZbXqy+ryNcRty5ljEmWIkJSa5bN
abOJWhkR9I44KQ463k4Q3GvSax98l/JK19XWtjel8NyS6RW0CpHjWlK5wHTi2orXWhoDnFXldaJ0
BSUs1Z+Fqn54G3TVdtSZ5xAiifRv/MWGYrpFlCfjWgSzNH+zlC5YmObhQpl1tm2eGT42H0ObNEZ6
AY34kBDIcsjaLrDjH3ugmjSRbEb+DRj4f5rFyLXIqhppt0EAlLGF8gzwVlX8ZKYteQH8Ct5NFmTZ
wVXZbLq7Cy3dpfC1pJqVWGXgHuAqd/7UNmsMg+vwY598nckg5iWJ4SeIgQdr7lSRZ9tIxZt3EkoF
4xSgLb4SyUaoz4WNKSW3RM0d4pe2PVH3bT2BnCqVmojfBA0t6sKzu7sr1/llhcFGjCKUsEY2yY8S
5fJhBUQbnQOROajSvNGyV+0kBPqT5Go76jrMqcP5UHmaGbwVhqHuKv9Ucwj8L/qdkEGk1KCqJxml
H7af93zAT+jfAsN/on+oa8yRf4tvkK4wGaV3JntQYMuZfpLrRcDsiOpUYlYTAUoh94+2GNWs6UOp
f/UO5otfEmrF6n/7gVQ70Hps66Cdpq8TI+x+i9TUn6IfbRrRYnX8AAZyATRiSbY2l9xAAFs1QAVp
P6Duy/Ckp9VzDQf1VHAIEif9IOLc8boP/eBECpWSGa+XSWIdzlrE4i52K/C8cBeOD9xKmQbKsrwF
8cYzt4gsg91pZAcntYxMnYwLMvkm/XjQ+QujjIrjtdLa/d7Ns1JzznVD0nje1lNfTkLqXSw+mJyJ
Ulmit+5PxLsftgUnspACtzPp1YPessEjSBRN0YM1aAd0dm5ZXOABScJ4BxD8dEfbPhd9nhN7LwVl
SZWbnlO+m7L+wXoTxLZYww0sd5IbriTY92nLY96yRHZWSy83ioE1QUr7abdDpZxYQGQd5i0AwTjU
LRwbU5yLSzzkracbUtnhcyW3DcvEAUyxWQJcJG1WTiSpSVzidS3QTm2NvnYw/lwwrFTcJtOnbrNR
Iyeg4SFmiOVRIj7jeEBW7OEFEhY776KXLHGyWW//FoZCYi0KXxI8SElDKWoTJR0ltU4FIlbkuJhm
VJbs5uf145NQBKEdCq95p2eeX36+vacNVCl4Su2wQyhWqe1k8NbAdMRXMOuu5OvdFtBDaZMwLjl1
WU0np0imRvYgQSccAWf0GIm6mg1V9ucbpTh8f7wyawrAETPGTUsJODNYBDh3D1LoWW2cCjgvcpDg
seSfwOKv33khfJD4mtw1fF0lyZspwa1I5EK0l1Bw2MEpBKQ1ijK2qVXduTZxrG4icIwb1+yjOE6q
tktotjJ5VHHO0svOah9CJD0Cg3qtt9/jqq/D8pJ2/wlZQe077hvaN2mwrq+0pT7T5nOtuFuj4/f8
1cx5cl4yeoe//WWY+/Q3Y3kieGj3baP5PhYrxqKDa3E/NoaeiLQYTS7Z/JubD5MBZNCHJlEXPnwH
Q0LiUvGeIzAJFRTyPLtII+I8yJzZnsUdH83ffVK96gIBBCLtd/66lCwnEEv8BnIFJ4a1YoKi76Zv
O98EkyGbwJ2MdtI/H9Ok+Hnv0GdLmluDYKi4PekEKXb7b6dTYK+dZcppzMSxbdBNTKHEzCES7xCT
EWrJjx9eZfkSuaD/vNal27CX5UT+0ElKxvl87VCYahXDK9A7vcfB73dNhyErSfTj75ZJojI/kWqu
zuHaGNlXHNgMGcWkAFwyWEw7ZVpHE3aV1KeEnkSIYVBd49JUdlmc45K6kq0AQEK0fGoFGctCp5PH
fD+LMtN7MQVCOR7+dHirVQuav2H0LQ8xSCYJgMvN9/TPJbm3OJ6In0pC+tA18xxonYL+5vvSXjfL
zrsh5GbRWECLMwvhcHUHcOErH5gbVo3ydb+DHD1FqtjEFUg62Vd2ZhlvfOisDq0NYhMN4I1NGh2u
/d92gJUA8J6yZo9kEfOChhRhoBAPjKDeNnjWDhu3iuj90rGBsbv21Xv7UrFjUSXi2EuBxeXf6nLC
eDRQ/QhKGBZItrOfZGK+DsdeO28yWihTbDW6FDwSSuqy7As1pJuqdI0TN1f9UFSTPv6jXPQGDVTG
pZ5UlwUHAWbK94VPNoqBCS2fDAUaEThhGh/4aSPnhWQ7w4r8JzZSvV4HJqXIM4XY1hFeI0btouqh
RLEeBceUXaZtAKN6tMCzFXvmyRDBkr91tMZhSiU179wLX4+h0i2sFCFIcHple0g5JRhhVAkIMEtM
Qm9roTR4DuITrqFkVD860jzv8XlqDNI5fewP2Bda0t7tcVbKKS2PUROIAMz/3YeSN9n/xQw4ic4s
zy/kAv7qWpa8eDxevPXijlDxqkNkaYLiOZCl2cl9M8omibLUqj84lCjGwXUWehZp/YOd68nrfF+D
7MPxadagxPV8IIe5KGy1EoLtnsgjtGpRVsf/hHB4sUohx/OFmgbhF1IGak29jToej4iC7iZ1qCry
j5hqXKXH/lKFp9hKV3warYGYjc5aYKT5+YGwFWb+MIVd0SG/UNwK6f3F6CCx64nq2vi78fsLjH5Q
tfg3pOJe6GtlxfeCIUItsyL1W+xab816egk2ABaEh5XOjuF0NRyHthmaHdXzRK15xFMC59IffLHs
De5GNCjN1007XsAIu88g3v8T5l7NDknwU/lgPAV6JYv05HvmH8zYZLrYIxLmiM2s9YnN0/0lYMmz
8Einf4k5UXlamaSktHL7XyDiu3J4zvrANWENrh04NlFGK2W/pGIX3ETOXJMWDxE3fMBnS9aL9WQq
E3D+jrmXkjDty58cHZvJop4ndsTOco9xuhwHyiP/Uy/PWmGQiLVNVBXgFAh2gcBilJCaf1hHv1zi
x9tjn2fkau8HqNoXjIzjBFEpABNL/ZQ+KP00iU6ADXQltmgevPJNleKrW2qag3kN3MUSRhwzElrM
2CAOBox2/JewKu9xeUfiyEV/KL3XYLb0uGov7HjyMNjXPQ1xcKvJeJqRdfihZJ3O65KCLTZ7ARVT
Ivnse/4JnK5vxeQNNo9UMQdtju0AaI3fe77D2j4NT/JlS48XDDqbhdaAZ3vsnejxOnouGWeS4OiF
WOY72ZpQsjjweaNuoxwZEmRFqCMokfeu2ABU8vvASudh1TLoAftnEjEAJQM6MByT1Eo/sZWamunf
mPcSugybqIiGO8t2rPJ4OhDFL1L/YVWersySef0i5p6NJHXfACYf6QtT1Xde9p/kN++ITI8mngT/
BjtE8SwbjzD0ePW+fpI2aJFI39ZBKo0OxfLtK5hjQLUecypHSdZKihLN1dmiT/mxmR34tyO8TbFK
IMBmmysxmnFI4YAWjp8m1LsV9Ol90X8xoWy71SvvhQDnrr4VNFSnLpC+FXJiGz1xkUaP2YcUcbDX
RUWfnxO8h4dOgzN1I9nwhM3k1G0R06rsoXMSJepCquVVU+/Oo3bCCqFA1oil0NFYxywLuYHU3H6B
yu6Km25E6Ki9qqjJSfESknX1Bpzzstvlhf1arToE1DS2fTpBx38JScGk9fxtSFmMU3J0GF5c/V6r
4POX3HMaLcZ2guakSqiHrCdS3EWQLylxWwdODp0g5LskFMrWaeGX4N+G2bbzajkzOKp5d3C+ADIh
vN3DoEtnoOhSeJ71bfATEr0eEOPtbhahhHz+th567dGc5vWJ8k5i7d0y7q+rthRCeYdNK5jsC9YN
hGeRT4iOdDOlFOaQK5MBRmzloWXULbYsDB8VXYOWtCPh0nqRDjZNLhBLnIZgppj6o0h6kbUSOU04
/FysIaZhFnWjHXwTZRS858L11LO1apsvedZeblHduGiULY5JrL31ziMjdpjQsTaY+o0mEx59s3L6
SDot6u5aoQbCCX9sABfs5AMD8r6JX3TTDoa9iyP6H87LKpubG+SFkYE/lJ/44QvIvDCkxXhfKfVW
dn9J9i2ZOoVAhjfqaGVlfB9XQS6jcGb6oFo+t6vT0BItBEa6YbWA0ksH6KhFf6SJsfQ7nH+VF05w
X9AiJrD8XN/DlSzKoLuOnpD6e/KzLYGiIRHkhUjIDc5VXXae2CQfz+DaUgD42UZgJc1Yi+YIXLgC
b4C0T+cDZ/TgQlzvq/IC0gN9WKcL9s/rCmL9VdavK0OxTvj9yYGze69Zz6Z/YxBAxJhsumhMfYH9
eNZ+ljjYaCouZI5nRfc2oyoL/Qoh6WkjivV6PhwEYxqnZeNmLTDvFrV36pY2V2CfyUaa6g8oahAN
fDI75CgjOmvWVCnQfjU3sMn17ayw9CXJwuAxmKdrVLR0mQstnabcm+KlPIMsJ6kMK9C9l2ICxIZK
2+EXGsfOnHbhDrFgPiSsH4ghNOFWZ2PiVFvD0SloOQocko17cX36/9CbMaceowqfpbbuihEoX/j3
SFSdVU5tWnB/jggFcLtNgcxW+YipQsQOACJLuPjaFBTPNWtAHdWmzb7JwTNbrWbCwYpKOxEpYZZZ
Yc1gsYfUYf7kItzdZodH6lW9MrEMGx1hG5ZesOWomgErxK5UE9iqWPBDWRlb06mAFgSqKpSZGDvN
XDxc3/qqpye28KdhUgt9LVED2oRduu934pcPHnkmN753Tsq+qDvZ5AWPGhC4Tpzj5gKV6rJuNjEI
cbn70lKmIblWL+ghM8LRsP0hwtwvI2ronkbRCc8/DFgYa0aFuQVheLFcJ2PVoWfNhguQDXYA0Ldd
mMV18YTQIfJ8AK6Kf+vZWlTo7BjKlf68xsUXYjfcrDdNZaVRKUw6bgeZpM8m4vXAFCxqrJeM9epp
QWbUglcmpvgxGVbgdy5rJ98/zccm/j6qy/5BgNC6EQIzgkz3nfaB4fTLRx2AQzwhS3D6aCAWRKBo
h3rrSB1MqdVot7hBuoCnonPdWwQqeWDcr6J6mmzhAveDIETbABwHJ8wMxgP/FRCsMGa1NIRhUrol
xm7CaeO4DCtvEVeamV1o70xNxPQAY3JomUy66t3HZmsInat+OUhNwLGOUzWDaABSuDk9dlENf0kt
+GVu6M+cGeiNby9wCQFtMzJ6Gvh3pCricF2MNfwZaTOR0UQP03IWCdXWJ0oY9sGPXJpm/BoiAjYR
XN0Kt6nNDktiRiO7OS+w0nWxatRcqZg5kPlkfEJmQrobY0ajH2zENOdVZnMZIzM577QajT6gW+jb
ypWbb9SfEM8dL4DYUBNOu0XxuyXE7dBUCn+iYPXTJAOizE5dmALPF0cKJFiJ13de81/VGz7RDVVb
cj17pGyiWK8IKRl6d6yx4T6d6ZE3PfbmMqZkF0ngJo/umpODJPOKrVZ43Zv2oq/6jVWq5fh26EcA
Ve+aCOo96nMjuniKdM62uNNoQvEBC+h4+C9826dOyss1JjaEABlkz4QUelZ69E6jfCNwaoOWG/69
1n8EXltyGadoy2BFbkWJVQZ7EXScKppLloJpGFqsK/RRjRLDgcQLDLEFLgkxi7YXT42JlYKPQLg5
aljXt078N+Ora2t64rauoqsNliC/0uguICL3EWx5A3yaEjEYCc+bxaD92vu7f37ARyzVrohOddn0
bVuBltj+Q6H+sbniRfIESgzKVohF7r+hTCUv+De8W+e2pqj8BRL4mVTRQxo45tkpSb51XnCrtw3q
/m2tjI0x1H8JTYM1L2v1qIOvMXVmIbRrN3k05xd2fFMLQcnrmFcsaGIzwdz0ojzxNMmm01W+k+4L
k54WDwSUEi2WSNGsBweLVtsLqYZ2SdpJDDlg2VJHHDVJyMOlCqBqnaEORZqL0Dh8PlUOJPutATBa
kvom1D2sd/8AYR2LKKnw1j3rKiQ3iIDZo6/PiFaPrkrYCBE7y6MmRn0GABJ63IUDRbPhQ8A2/PPx
t132dG+z8uKtk5D02rbySp+m+AwSQTyybZ8DSTkQGVqurVtqsPYZ7tadI3dtvdLuQL/Y4DP6DKbb
V6c/m5AWxXr8EVm0zc3kmc2cR8sZsEonT+hWu+a9nuI/Coruv5RZH6tag0eLnaws8U/Cc+LGZthN
2AZuHKJt56xgVtLfjfKY4ImYuqUgaPmO6HASds8mXE7rgn/35cPDTADX6Ga4TPy1zc+nKZA89ABL
mddQXj+Oe1TGpyCE5aJCtK+LBhDXW3P8dHh7Ebmra73mmvTuZmo8n40tp7P4D07NTH4mdq4G3ftF
DDBCmQEnSfpZFU6ZD2tFemPxON0U29cyjy8eCUo9+omVy6iKti06CpIXquscGUjOZSVQarR/hO93
RUemaSjS0y8gMTxklMU70nzZHahxP6djB397etF0SNStCiIfV9XpYXf/SMfgoF2rtm1HO9QRjqNz
oXXs1zE3wMImGagGjku1ZMLFh30U6z2B/KUU717EOPDK5LUHJJxTCe5Jpyk/mw/6SGuoIlWvZq32
JmADFC37G+vWUjwBLvPGjD5Vnr8df7crFCkMspt349/hSHHMFNc0mmdyTlwmeUphKpmzwdct/5N9
ZUDGSTYv5tHGzkWiB06PBwcl+Z7ANxXGY0Lg9pX/fZSQNXH9DBwGHnH8IKx/PiYB6+sFAu0JJMTY
irQ3JZs5clbxd+ZtIOSmvsvJ3mzKldQl1uB/f3ZdAS6JUX9tlPeAh2yZupChGiKSHs7Wae0DPXn+
L0g/xZxf5HabAc3actLS8hxgIA/54DlPSqghgtqAgfUDb/rmh54EM925t4DFqH9Yv4+hxC6zfTOF
66nerLjOtY1jJwKVajl4ZYiH0deB14dLPmBSLUpStF9wR2IQe2PzRn8K6A5mEOm5U3XsOEAQzqyx
yU2yuKNhpi7yF2G6xz0GXBChAlBog7IY2aeqEViZ71lPrQnW5FajN5TJg40CdBgg+a/S81Gzbr/+
9sjL3SLmxqJNfXgQLSNOTbXGPIrsi0JnoWZzpb4nzb8Vjced2T1nQmvRpoDJtr1JZHgRUU9kql2l
Hul01qThTohBU59k2Jyln8xwcLHpaH0WnU+WdFUsStBukxt2yjpZFK1zANRasdyaRuj394hBzK94
TwLdBEmQ0ibU2m9zhqVtM3VyBgKdW56ZfD/tZ2hDsFFlWgxNgF82u2alkqzvlSDZ7/ZMu+1r4gqD
LS7EmusAPb/KEyZEa+WBb4LAsqo8B6B56ijaWjs8unOyenSeUKLSCWfnJKVjdPhlwPf0JsGrDUhU
Uv5BhcsiCxazfhgMzgqeGmZq3DKd+BL3hY4bIM86GLZq3+Hu4RwN+CBTUiE45oisy/BGuygpqt4k
Xqvb2YgYsgZviDmGdULAHUbck4r1Agrr8a1/HHFm4ZnjUCWbRcPMBMEPzQf5SsXaqN4pBTWn2uKF
UJerXOXMdU8HolwSEaa4t8J3w/8vx14NN815OyYiw4n+v7hdzbKSiW2ZRK+CJjXjR9m2GEbJG4aJ
GkecEpkiKJDtB4tcJ4QfSf1t9QN4Xby2QEMsboQCoOAYv7QrOHrfy/ReD61yMLOR4+rMD7fv3W0P
nh2pu507bC1gCR3/q7HeyxonF2Y/uWR7bieN4J0dXWxNWsI7ffVkbRYKr+yxz5boicQDmKLGiBG9
n4ZIbE06D/HcdzENex94L0+DYoW/FSh3dWcFD+HcE7IVDNx2/yzaiROnROWzEMNVpecNfFmLp5Yz
OPxIdtGIuJK195ugY1or/ckO//8Ac3ZU+/LqHXXtK8HBs0GyPtpgpLCPOsPbYpyIhrrGsXqOWB0c
73tZ6R1tPby24HK9pIhfyVGQMQbvD5XFk00w0YBU+pZ+FVl8Kt6RURn+jYGaXw5ukCbtYcnISJo9
jlz8rOmipbjCi+sTrTVBbrxvhtwzxRhn1T+dJpYLucgWgxRySNO/ye4suHuQRoDu1DNefx1QuLOv
JprtmNLEHPtp3uSuVKGd2heMHJuiT9gUfKDU2LRlnX0xxunJ1xFW6D0JxnDR2TUMbhnZK+UWuA0c
/1mUeOL5EaqZB4oAZNduQI7ppKq/27BhnlkMDhOEj+YLpoJ51DFWDVj+SCuwk8uEDHLyL2w3PiVr
uJn/hUvsM8eJ1Gfcrq2TymRqiG/ViEEOYoldVB/Fg0DGl2k6I9/pe0CxrabOCu3oWhNbuCBRN1UL
5n0cHo0jAFplBlX2UDNRZPBiURD2reGVIKO1s743qaxltIYwXdD8Ydkz9KhV3Z5sQ9o5KeSg3aZC
1zECcK4bcvV8KOQFo6IPWCtt43En4WdEbXlYKNp8eioVV+FpcnIhTzc5M2o8bIB8uScEMwAICqWi
UDNs+OOR60/IeG2mAI+Xeq/ogNuyqYVUIbfsKJxVqoXn3Yh8QAp0CyYyrgiGn5FwEctt8vMbkCf5
J3ZWxXpCC88gyFbBFUpm8tbpdAb+3cPwMGYZMS6Q+V5qq0PuFAWcDddk8pEUBgpZnlk49CC2UTsN
VwKYkGYiEDGyGrp3ZUuFbh99JfvAbTHACegIsAPBx9uvUpFSzZdL6DKhsYIRtVCqqWuulo36lSVR
4b1qYwOfunoR6NCuATG+LFKLH7McBzzOPvUfjqXV4tUpL7Gumwuyp5EYvWYHrEKYojPLDD0Z+4KF
E9ZoDcZz94CxRooKpWRmMVS4I78TvIUqkpmOQvkIwOIGTHPhnFpNnHaSboxFHSb2FnUgJdWc6JCH
wQErTu8SqF2YKcB+4UdrG/jZ8RBLbl1UR7t5ugUCThReN9cgE7UzaWwoHge7GpDTrBONTZ3Jg6L2
4oyIF7ClstYpbXPSdT2LYNjJonU5nO6hoxdbeYSJwVzEn/PUEfuvtSZUXE6KMFvD2BVhkj+z2lY6
ESAKG4GikhjN8e882MIo6kWxFKcqIjlCrl0IsejaatYehFYqI3KQZqcFJTS/epqwwMpBI5GsjiTU
3/61uLwrk72fGcmBB4WZkcS21+9yoQST1z4xDw6R5PZdQQvGBPSCt7Ej8KTAC8eOahUXsyRHiDmV
CUmDR04iRMxHMhZ6CZTnL+RstpnYv0N2j+Ym5CamPjbuAHwtIPPk1ki37i8COBB+Ycf7xnRvskfV
bpGHtazbpWHpWeCC3oiy6/kcMBNvB901yDcvBRXoYQNVZtV3S6YEmLm1QzilUqAj5vw2tB/rujCX
crIMl6hlNagRLhbjwHUqmV9wjhcXVvMnmLv0g4iqEB+qS9Nb8TbjV+ikf3acBaHNQidUIl+YR9FN
n28K9Bk1Ar4EjOhrL6rutcBqIiHJo4YphVgpMBErqiiCtR+HKmLtk6WB4edAP452nPaVOo3HjAKq
4M1Ph2ovCMIE8uml/GW2Avsv0QK9uTl1ons2m294AvQpbcSxp8YQDC2w3/oQUdLebA8tboKY1ek6
lLENCeYQSLHCDJSLupqJD5xKcBaXYMJYuKztNpxGz33ixgKOfuMISV/SOGtFOWmyVA++woiSqh2d
aLPspekXrntoB40xE0wDXt/DZWzh3atpishgkzYE1NGFqrOmRD8kLm9S/m5FF728sgiscPqcG8Sn
KhdoKr97GxEYyITSdZO2YZHJM68C395E9Y05+2s183B5PjMS6GgttqZZsQXjmZjf7JWAvESkJ0Pb
exhl/9naSnf8whRB+XphG+BbGmNwPH0+ljKchzwKHvW4XjA6LA9RkH9KYVhd1JzGshNZL9zF8wEp
u4EecN6q6eiy3guPqdZLYY9FAH3spL0+DbRexXHr3gNeSjGkrklDWFvLkcn37uqtwNUDgRbqG1Fv
Ri2EGoEAt55G4OvoFQaiPvgD8pNBohu4ejOVEmanuP6fAvnxiR4qZABYMIdyrsZ6r+tlg+vfpx1m
mLzDCOtLcYSVbD4T2znOjCbUMLj4tGLPU5dScS+mLbglMcRGTj0E5I2/6sLSkdtq5Ud1Ry8A6j4V
OnAFqu/ldBf3QSvT92Fte0oTx5MJyqF9H9nNByqgswotr/HhShEA6rEMYST9iI1x0F5cw2WfYnLb
7DfvTUg7vCgINSbF9WKF3m0rEoLc48Jd+Nfll67mVYINX4Xqp+q8htuIIT+85smwFpJeuh9QtNtX
IpY0QOb66i4Y/E7f9g7phWk5yRUSOE3I3DyXPz/YLkqCDqNNd1a099vff7smTrkp4Bdyphf787Cm
GUEPfngN3jDAiUGLuVMgw9RHwWILO5zPq5Rkhk8QzD36TYsMw5NRsyYLroJVuDuW53aHHXfM746P
r8Q1/M16EPwRKAPSuo/0AijajWBYm3n+JXQ6t+jAtyaoju2S5T3/8Gqm8yWNQ+sgpHtp2dzYQ88p
EcFkVNdNmwAY1FUPNyebp24LI6N0a6Lhr2EMlnGyLxrHgdiiMDbT10Wi8tvL2vmLR128khy8V5Iv
mZXYZJ+pYnPky9D8gK5yJcoZTvr2n+NnnemPtN2DvWCCmh+N685lY57rXgNXo3GF0YfHJZvTstIA
WHFbbEZftZpuoj40jtT7u+Shq2qc2m1Dj1jYZYJPjyNktZk8d3M2kaeTfxXnP32Ss64oBXGOt1ot
XHjSkwsb5ZO5xcB+aEzn4wXUZRr2Pgek+uLYt25IpNioKW7iw+EfbNQNBpgi3+jO2Sh4MioZchrW
Q0jQ+mvoNR02LZ2OCUm7qmvQ7tAyc6pc3iZjLX+B1PQUIdM/sChEPNUku0qFphRxGfDUIphwqIr0
dj5DUjR7tnFvJDp+uy97OKTaZ5pPZk02t1eqduKpctIw8FGtZebjjtgWMPzTCR8vQ7QPNVA3F+tL
Jb1z5Vuur0KCmFAia6Eb7aghbP7RriItL0qGOcxl5uDVsNAyUdBKpv9fcsYj+1gBkxVsSQnOAN0u
Di2SFBylndDRW+7AUhjRr+LslIe/Pa8GAFZ4qwAa8Md1O/6LMqW4vqfhJilu4iaoYnYRQLc0iole
2Vqnsu/zUVsDSixQ1OQ93oU7tT1qvz2CP2+OIjPPoKVkVoG+PmY6dj2mrZdNgEAB2MgMftsYwVRO
3kf5tQUj/8W4oapktZ3197uj7k8YzEkj5961wgrtUT6X1DB5fR+2zLMcO8+e7pFiw//LrvuUk6F8
FqlrMWMVG8VIfPPeqGDRc8ahE0pVvBbHmCT52I/tVWfh9YqKGlNhZhIZ3/lLceyUGHjfjrTdzuEp
I6q6qyAW9wIhuibcvzOCEthciarEnGCVs6HJIAeFkvn4dYBYvYhfdoGAb4Yy4cZdojViF0072PDB
jVhtREvD+VaOM9YFr1+1hlSuLjYoUlN9jAXAyz7RyqwW5VKUiMs6aSvHqT5A/+3HJXvFcS6AyAut
4ySBr7vudz+a2h8VwraptglBhd/9KBfkS88xDx5p7u0fAzhqGEe0ooLogZmqa+1KYTTF5l1EWjZm
TSgRChmZQHp0LKF3wJczvjv+o1PwyTwivABo9MEk+8tYe+0MMXLqTkX0zrLYIqL0E3iTf9Js9Bmh
DFlTkyNYZHXbY6sqqO4sAFGx1+prFeApDIQsti6JmyNaPesTJEAPQ8s+uAd9j0SrQae5+lJ5bvHH
MPZ9jalhemp3jPbjmUMR/n7phJUEcuJd6+BV84X5dHEFW9kTp3N6hjjT7UJdn0k8jniubNUSavNF
4Wd7Q+DGI44A7DrNkmx0oj055sqqtddcSTCqwhtXLEk4dVVtRk9TEIy/taUvPAzWosdKEQeKSFiw
73h+ry79zG8aHu/7UbZykarqV1ZTH/Wis++SqI/Z8lJPTZ5kQICcqREGLJEsxvNPin9xS5w8jPnV
cN58mwYrzyyzNZcvzFzhQ4oJowjFckOtrqOK2PN6PUxLaA1CZJZabTWXj96MmzLN2xvp0sb4E3sK
DxEj3DAzm38yJgQsxbgRlsZFEqfbtSC/N4XzhfWN9Z+k3WMJfERcaAK+R+FtVTBQI5uehuA2Gm93
PEqWh0/qLxHTiJWfxk0xPDL1eD/Mi0N7Sog3HtfIE6XY6jUCPzwcAgl4aBfXE2kTj5T6XGFrY2oh
J8wCZ2hi0xZE+MgHTl14tVBl8SNNfB4kzaJRRkRjzvo9phfEz1F3cgsF+TCnRL4kL6q9zdVwDdxy
d3b1G8TY71esdYutbADM7wGZgXADLGZu+qDkT1sN3vL/9XEQKSpW9SCQS7dYoFW+AJh/Bw7Y+ntV
ytd/sq2+d8aum8URlK7JqAduYE6IzaJ6xTh6XSn21Aa/meiGaSxStQLreVbBTWPhjCL0+1UVZXiZ
aZedNATUJLkziLNLNR2mLoitUySypADKYnZHm9w1z4d2/WCuhYOHSpwNcbT/SmhnEv/otUXn90rU
yO9O5fXDnB2YytG74cSBA/QILQ8uSHAJ8abA8xW+YuYw2Oom6z2Kf3TptZZtVh4lX/Pdw72KsU+I
eVxQMT+2OvMhci2m7ZikUwWsSlNISOOfx+OfV6Mu8zzFylrcSKITv1jAUarVpCKExMwkhqfTgD3N
mdetRm5kQFtPt/Ln6Cdy/gBJBot9Ake18QQfeYdW9vwX9E7Skmt8itrPkS163Ua/tYCaWaEMU7CQ
nqR3hAy4jW4N8qjI/QV/iBD+AQnwmmAGOcZ3t6o0uwDdOP5lz8uG++g4wLIyhrE3bVFtP6lhGVsc
EFU5qktzl8m1GX9i84V4WCk0vX3yJAV56vVb8VdgB4QHEtLatJh8aHLpDyHZNKAoopeRfix/aKR1
RCMymq4tpR4DmtSaeRPLW5n/xwAGYEu6KH1YjcHBxUEr6eIXdMuHPsMOrxDW2+hKMdKcTrgPrJJj
6oXTAfwQ9bddEEIgFSXzPSjCfeIJ7Lz20VpionXooAoj2v+bXV8p91ZffgdviT9zmVktEoeLw1Mx
kppO9mJerv63VuHvOcUYwytYNLb1JhVuXRBDWYgWHdQns5INqm2BliFhxvi8gBSl4idrXCFNg468
x5ik+CAeT2dGshI8SUC+Zhx2Cy+CFuqHtJfWO8nZdtyUf7wvmVlUuo1TYn0Udbm2JYMhngURyXH4
RAk+YEWjf4WzkW33ztFMPkerbMSATRe6lapRWB/yE/NmHaPNjglKK4PHM6KxDL1KcpY/kpYKuTi3
aVWbdPg2BpKZZONkhcu/GV51CwSTYMkPNiM1mMixRE01kXUFdzEBJVbWfgB7ZZZup6HtxWOmtlYd
3n50H9IOyBjnGFGeJXuK1mZxlWlzgSRSo/bypZ2tc/pM+jnbJJS+Z/ZzrkjdJ0/s2psHASWIsnkK
tEB2wIDsORU+8PQl1LAl9vNJHd477i7j9lABYN++b5DxwvfJyRMmum0wEczCJt9i4v576Nc8v2xQ
JRBdobdr7OznD4y61QcDLjbxuWIHZ48di+vmZChzFBoKz47/rJ4b6cIblLqpanpwOEmEY3T9AZtU
J8G0lfpds447UwFeJ/Vj+1m6exyDno0y4RW50njUPPWPY+lfMxCrF6zV3IjKGmy3FhzWy0qy1Iop
fZvvH/E8RDR5fp4SevBJ3NcxgHpzAA85U6lJkSEQSM+28yvqq9VMwL2nWusMKgp774MVU/YzaQRo
a+D5niZXOqX9su0INO1Q1ILTbEq/SYPgB4zZuew0cYHqP7jccVUl1M5mUqwcs5a9b0Kx3rY5B3RW
FCRLLS+d9A7uoZBz7YFPliKv3evbT0bUvFTzldzsZC80S78yvVBkN2brSoXljtLe/S9OoMw4H5Eg
qiGjhu9AwkLlKMkqBatBcC6CW5Rzwsm9PN7CeIQohPYrFbzAQwJ3RvlcmxvQIiZNLflUztGMj5Z/
D1ygaoHnw3vJ9DRyP2dGmQqvwKC/NaINLWA02tDqdUSYX0QaOVCKbfsFPbRIsL+pM23veMnig9AO
RuA0z7znrPDSKtTDGk5QtwRtohdJ4ApVklEVWDt8iAeZQYF/l63oVJjXxl9xElKm35hvZKIvBt8x
crgEGKyMbZ2sz99AKcOk79SLtwbxyjbBu8VVoQoGB7HS7s+6C4jxaHav9ixOA+zDq36j8Nx4JYU+
y/mf8yWdYWIiCBwKazKee/QDFVGqNA+SIJAjPxNs23sDpAJ+2od8isRAZqsap3j8yfhH7FpUDeiw
YEXcKzGQg9XAg4qCjNghJrq+Ly4/4D0P/mEiFIgRo2ExsQnIAzccQHkCPHTAg/iGyBkTs72cHJqN
EfSgCrZ235DuW6x8shnPawswA+n/tic4sdQUBL/nXkpSr69X97EYGJP9UxwOXQQqMRAZYqDhO2+i
qDZlO8hFdJ1AhSK6JHsTEMdmxtBscfgiSOq2ua6/lvNJ18U6rdUUQcQWiwIQRPW7R2N4EgQBeV8r
PKx3fAw40hd1BgKItKM4HuK5aQa7BvzWdLugqoFhYGXWmGqlLlH4A+WyJ4elfmMYsh5rD4sJ3+b7
38/ON6iF/xh7xvf5tRIhGWawwlxT/x8ingGEqZMsVL7vy69oJEZnIu+IOxl9/qg38tN/b0CevCqu
Yv2gvDA3YEyey3I+JVbsBcZr2MTStITPnN2g4K7495gt/mRSEazmZMXZNuGODDgziacGIz6gGj5h
1qGD9K6khs2RnKdrMEhFfE/C/UrHXbmjK2hwVILA4WrduCbyUYKWTBaJXz81hQ5Kez1KQMsIAOqP
4V4jZogAOf8h7dDKleq8iUThe9MWNC0AsL+gW/i7cafsbW/3eVnzF1hbntC45n6c00ftVeA9/yD7
TEd19ray2n3gDmg/5B62cL15ZRFtLBenqIH+vBOggJRrT8A4LdImeDE7vZLEiwoKRYq5Q7M/hIwF
ogVBxSF9LCYq4LNQyzNGvpMalhAvqXDL0W56olWuBSZNoYzbsBn/wUOSwrkn5o4jzoylSXSvMIGL
ob12iNFPJSpC/3igQqQy8JOti/qSz/LCHdpyKzZWCxlq/WjaWWI9v1r9dY7vcbJwSlF5xiP3edIP
CvurO5YwQcRODbHO4bg8rqy8YYVCdMYuExJqU6wFKBZWMJv+x2/bKWW75OX2wH8tKuigrYdFF87I
1vu+NJQKGYCrWlabUE8GaqF+j1cMUTbGpjjU9u/3zIsWL9miJZfsw8fpcrvgrRsE62vJBPrs3Mct
N6n2v7Mkj1fGuc6pa80ODuxaYP433O3+rwTsxBDSYbJqGpY2nBlzF0bxzy0e1JEaE7TlxbzM9Tl0
KpHu3a01YFsO4dHdOJvQWmGeHxGtDwaxViyFRHtgsukyxb+fnU4ShHakJIwYagEhk58uCYAVJwra
vKvo/zdq4ByUoC5mvBgcGwQPC2v9pSyZJqfE67bB9uDUDB7cSEtmg6MORdoqz+a9KrixySTqEEsE
BlF9HtkM1muWvevu11epW4mJDhEoan90reJEeoTxAW81NTy6TBDAwlcDTAvnW3yy6i7T5PBVdsNV
mkc6DXMhTxp3EbrWw/nWYx6DWAqT3/tTdGwvqJyFm9BfV34GZGb1wDyMyHwlE4UYWjCFhRhWRU8+
aRHoXQfQjO25ak85YxJMvybT+05aA7VRMTbWlYZ1Pds5hjszcSG+UAuycm4cZEkCbHhOrucUlTBT
1QN7fPgSYFsl6zpkzHYqt3NWyc/Yl1xF4pL/hT1DBQsR322KEOBJUB39KYavnHvm7bfNydoRIB7d
25VbalH+fiu002+lkJ5iAHk0ii7i/fwz4TWGbtebajSmMn0GyDjWAZCbRbfcr1sqdICXtIsBg9PM
YC/dftFNAsTOIV0x/3TptfNj6UaAnY6dKB0hQKcUbwBTcIINF96OrYjrL/NC3qOVWcwqsOCWbNOV
xPSwaFCcmn8nekTZl9aer1Sn0JKpj6ySNXEIOf1W6/ct+V1T53lDqLcbTvvSZSJqkLi0YOMkhNsD
RzR6XxGj2Yde/YnnXmyA1FiJ/NlopBBnaf5ZyiPq47DF/Uphzp4ovFx+a/Mt3GaTdjH5BU/2s5/7
V6BiFmUlO38CeMdHqtEp+3CwP0tCczYxVraD7kvavwyQvkmRxd/mJZzQF2cSM+iXcUGJbCHh7Jxh
/B80txISbcF9mKPeIn4s/E/mGJlzbFiVIJ/zIxP+LC/mFSn4pVLe+OocvybVfF6pwCJbaaKaMJnw
GpPJ5eOTi8+iJ9FbP7VEgCcEv05Mo2FFH/nULHMu3yKRxxRvFIBte86rVVf1qA24jZax/yri6ZRE
ThPsa1Ew6hlJhxz95giT7UdfjBxjnIlvx724qikwGXtpz9n9n+YhGb8xiNKRY6lVdD5M1MJLh69T
WPQBPhOKpdcNDfKAd3Dxbm8iBuG8O83+h9dcpVoESEgTHewQ3j1GeNnhIcmAxpy5ITFxN7obbe/b
1vJli7xOa5F65envNIxEL4mJMgU3rHMcqzZfnrnLpnsr4kl3O2dowePn/QC/Bv5LM3ZAfenZ0ZzA
meHOubasQPJnz1KBv/KKaTmU4sNqACM8fEK02tpwGnYuhG7a6e5gTcYuFaZ6chX1cBBbg0QB2D70
oud8YIMzlqEbMQBy95mKfK96SJSlXwjS9vilBfxzz3Ac+K+AxwXTp3x73X+QrOgDUxkz0rP8gN0q
RPJeOXudECVlELraQVRgCE7lBhoZC+NZZDTfgCdAh/kTfIdAybjvzngrVFiUi/QmkIrQiZgxL8Nh
8tFUsEfYrfm9WMHO390KjQ9wem0nard78xMnNEBkIDegb75o5+4BrZoZ86AORu7UHBy2fF17y5cy
L1VgiYdVHiJpx2jBV9DhuIno9U6HkMYZzpoPCiVi87/YuIu9cL8sxHmeq0h1zYSSWYE4hlSWBbdy
rYdi05uQlCKIeWlNKQPgWpAcovfjROeWn0QdHLyZrgO02gmG16tpx8Ly+r9cip2jG72Zib8bvlfT
eOn66I7j9hqhk0IxJvrAWTClGog9SJmWII0dfdTDFYYbZy2nDCxIZsWBEnA7tkhBezDoY74T4mAQ
bKNyq8flzaLmwGnTIvcdw8S79lod6H0BzuUYzugf7DdEyPWM1ZCztWXJZxjPG+vVSPDZ1bVmPQeU
KVWZrLrBEXYnqFUY2hOW6NUAOYGRLcJ9tIGFFVRBOBIku1DbgWZPLnO7S9o+6MWWdycbdkFJ1Utg
VMd+bph1lWIqltitTbn/g+dKL60sxIANIF3ttJoaskofPVJKH49crGlzvtfNlfM5MLuyqE8OqgQl
YxYjwZyQa5WTauVWr8WAQR7fIumkWFrwFj8z0sObHTrYVtFOPg1RKzIsegryOnbHRwN0QswqM5P2
pHO6YDLeK9JCJoplG4UF+5T/uoeGLJ9EL7BgINzugphv7ZUZGMwoPS+ymdynLYgaWMyjDORB/ZB4
SoCjmN5VtWTn6WnaumHAxOQRw8LyQlICFFa5JI6A3ass6KkAZqbQMZ2WobEbIczZv6+Gdc8DBP8T
Nk425CwY5j4dgFGxYsjvsgKXrA0rh9JjV99Q77NIDlIlmDj+nZqQweg4KRDNveDRHtnbCSDwFACK
xz466NyVN+aFMniQ3qmefxaNWzpfNYR3qSyHzHnWvxUgCHGiiseRWmOMxczpbzxgUBr+yybHIMxb
szjXqDaeB1snLit/2NTFh27ER6xJLjQ6mUtmFdL9uoySHS+vY0kOW0QW6iqQlPUc4uNCKu3jWl95
JSiNmrTRsbaFK0VevUpz2vkI9UFudNxHPxpPrC8ZEkB8PW0nFHlVqsrmX9uTLvyHe4SAsnqmOoz9
paW37DIPMGL59Fgib0r6kXoDX/pQLVPPQqPNh9UZrkRoS8AjxslzJdIgMoKfQp51HsprCShYCmxg
VxMerDPp/GCq84kmf0yLLLoCr1PMBc7xHoqgHSNv1wQw+VL7bnkuYkyju0dUNkAhK7f4Z7QuDpNe
U9omiWd6KJffS6UI5sqZn87q1l/vGLjHFXIrf8O+RbjbscNKdBPXRHNl9WshyMYjtHSTJj7PO+Me
QLH+U8GOXGFjivl6Vjv1C/zQq9eBtTE/BLuAPzcoqElEgGNeCfS19D/wRewGg7i5QI3R/Qae92ZV
YaYkbjaVxVb0meykJ93hPWiZvYeQ1xrqQ7yqJ+RqCgofMC5w3beJe46OPSthV1mKcAxbyavdTyy0
dArkgzYYCzKSnvEPLAkPCrh+qG3Y9gTc9uuZmbUpAPWeUYdtkcp2S+lD1EDl6hPHNYxi1NYqDmi/
wTquG3wJIC9cCy/QVzHqc7mNn+h5rWlBwOmJxfHwQ3dCQV1OL1JCleWKs1gEFYCtHGiM+pLbCFKy
wvw+JCdNxcf8P1rRD6JFr3PBaHRj7K9Kg9hSHjBn+L6z3KJCNxGeM9Qp6NTLjPxotZteYKKP0+yF
z4myaJ9zbGlydzOze5KiWWL2273zYBS5KUVKgnQDlasPdrSl+dlTl3XJ/iLiLHOsdMnihqenTTDq
giXjJZ3RbLBDWPy9j6joM/HmjkVYwqslrMOo7BHPRibYfOpLGa0rMlsoCnUteE/dKMQwvDoXK4qk
nd+2TUzQ/hbxbNlofw4aR4N3MDfFyRtVeFKvZ5q+S/UyWSBxpES6iGWmKv1qTWYiAw2tK2b4xTIr
7BhPyG7H/snn/Xg48HPPSEI75WE/K8VsHs03eFQ0mco7S91fqQyGSyKZ0fSJcrj7quDCkY4ZD4cB
F8Xrya1ZHIuCJCBbJ7lLpV5IyxCrC110s28RC52jDACEJR5LPmk9G8bNsxU+WLP7TWvi9f/T+1Et
pr/KNAwYaf+nrpX4bEtOh4rzPbl6I/kMKhfXC+fKdy5bk0DyUDVfMvdzoD5q/uqpEzelmqeZkbiQ
1rEKLyv1Jj8vF62VsU8u2Oq0YZ8Gcy0i9mQtbtRUY2I4McYctLc0JBjemPx3OKpjyRxfb7smFiPi
OcqXdkXV9pPw45BtQigjAmemCWnV0LCBNxN4EVA1kjdlr7SL3Y7+sYDa1abKmZ9Y+x7mOE3kPsvV
9WmWqi7++iCJAjxAJgTi2Zh+VlO1LTWiFU7tJLlnkcsc/zr4R391gdE0imx8P5BImOqoRN8OWc/L
VJlAytJ8ISb6FjyyzndA4XRs2rjrFRYohcZFR+9j8Nvlv3I9hBktq0WFtYAYuc915Ri8fAsuM8MU
lY1SaGkTmX+Le5mghlut9K4LzyELWqE1UuvRHxCQhLAW2Z+pOTkr6Ew1tHPjXnKx2YkKWrHiw+f1
kmktRUOTzQSFNUyuzfXrOq+YlMludiNS6U4Hz+zOcLvlmBwgJLHRSBmc1TiVrZe+vjUAZFVkw8to
An33mU+o9oA5M/60GYdynLpNpx4W9/Fvx6sOVn9jPXWafKEdD4gVF1MPxxsg+1CAll5FAeDos08P
5uKUh4exKZH9/MMFRu2D5Ibzmq3sv8wFhslRe4aKvkYas3lAOLkoMPscLaeFS00cUkpRa5cZnbgv
GewQnAq3E5NgA6CbyqLyXWijrT/Na6PScF9l8C3Npx+Wz1fPnV7KxqKHvJXjivJTRngux4IcIJQn
eF3ArBsCWqfzEU7Mw3MnYXlCZnaBTvxIXTIUQtDaaM85WxTrjv4mFQtPo7AbUq15VYo6QBsQBwYm
33zVb8FLu7EmFtJL8K6Xr36It6iCqjh/Vbu76zHFDXV5aI/zlkN0Z2CxcYSdJEFpi/FjUVuofnpb
9SCCHDIsZBl/NVWumkrDSuV2wzohiE8212ID50mOfX4ORYqDW/oHgxiAeaY7gd1RbP9sGNxl+nhH
vStsEnvIRIcONkyxFM0Av6bahvpADNw2aGFbXVY/h4yiqrx9JYpRVs6b+NDMajrMASIElvefh45z
hgUTlZsxWoJKqqUv/LVXPEZ0hb601u7QM3HnR5PQmZ0AthbIUP15EoGiEtUrvgkSMD3mOjfVQ/SU
1SQJnrNYOPh0ssM0I+ov2ZKaDbXiaboybn64bPVRRFHRBYLWjJwDSh0gzEHJmmXxwYow9C7xuwA/
k6WGLxQP1uHgK28N4kpeUSuNxRS4Zyw5EVv8tO5JZOep0BxXLV6jgJtSeF18CyrN4qqnx+l7nfAy
D1TDjQrjXlUxfUZnNtM4qkAQw+/oQjyK1FlRn9lkSyZN1B8VWYWeXcXvoIIZxOuWhhjUnuy1zN6B
pOTYVJFprMSxB7X1XU7nyKHl9/3KYyxeLkiJf/w0oNQwt98wOA7/DegMPZixtVa+NhHby1ak7OLz
PBYchP3NE9AmBlhlCvQ7o9KnJT/pdv44tWscuCM/RZSIUE7Rxlh7qTBQvlmpIhwFNNbUwRYblD/2
R4sNZ852gt83VEtug4XqCeDYrzUL5vELeiZP1Qjrmny76kTqsc3eGj+QPtjUSSuXkEO0z1Y78VLW
Vihs+2olbdnIdICqHNo3QvKDa68e5yssYpcDQ0zANK1TOhAc4KOZ7m85ckaypHA8xnka07MZOLya
+b7OpLigI9BU1ZgNSxxastwUtenvoXQ0mVgMwfCyHGkt206Rr2jmbrx9RxXCiqrIe659j4jux/Lu
5wdRZezlZQn3qu2DVi/ogXIXksASy+mPn06NYW/I3/SVYonjChygeIyVXt/QvKlhuSJzwwhA0Wsf
DC3aAtf8cIqzLlN9Fnh4cV4Lfk3HrfK2rPO5kvI3bwpbLKalpjvqO50dQY4oa9WSZMVBm6LpmXHa
869rjCpAS142xRQaFDmJGkDWGkmNW3OYv9nLMmWOPViZNM4MS7kTk4tn5HaZVvLgFtpLl4DxMXbB
1h21PInVPu6puAP1j7h56Mr+1acDFqd+UkKTZ7ZyRU8VlkjQtPKZp/PNarDUpsH9oEr/1KVK+jFr
pVi71gdtXuQ6MUySaxhN6ysPiFRyU8f/E4QbZ+xcIjpb+xLvxVj+FydzZPV97iep/Cceqimq2zd+
M0eazuBhTf38b00VDxn2Pg7OvZysFi9Ud5dBRJEYfATzGgqbuoOZFovShFfKQe6Exu47mb+hkkeQ
f/iVtAP2x4WQeV5luI/YcqKUOQB/7Y7UkS0vexkrt7/YPywOJM6eXCHwK+8YHtOVJabWGWVTCb6A
0iNXfhoTTkSI70bBGJWiB7py9sW8Yt6sCbg/QrO65sjXyoDO5OAdl2fimy/nO1huRHUnUl38z1KB
q0e2/Qkvm0KPOphCY6BMeU1STCQbazgcrBEOxzrIi0Oe6du2IbKK8k0WbSfVw7DpUGzHlcqe8TKI
1MYJCYGek+Ttd4WHs4MQLriwHxSft3Rf4Sj2saW1rgX5Xme/qwhvk7ylh2qBwHD39TtSsREajmXf
rL0sbxRxvnYjGAilucVWd1prJE9R+3zu/iRu7/mUb4GJ0Tzs0RTC3532v2I8QV0EI7/WCIjCA02I
Mm02WoUbhnlBdfqQTDC3X8Y1rN2j4hIbxRcExDkuS+hyghKAaq4VcV9861ULyPTg8i64dvfvuSnu
D6633SDxjfKJfo0rjkTKrknzXDWeOtxoaWFxecqy5hthfggSD3y3mZS7xP9rkyG7Om5WHbrQZuTh
uFpmuKlzKL9apu6YR7FhosCsLe5CraCLVq3JxGruZeb5HMgrH0nUK3KM1X6Jc9pMCgkaHm6qCOc4
1L9ybzgXorV6XMdL6xIUh2muVrCDvGMJJRsK+vJEIRfHpVMMzHRMdreBOwemMNu6eI4kMKUZvnOh
7QI4W9WfB7VqEt/3pLibNBt5vDFm14UIngsKhyxXyHsoRmg3lL53+IrlbOMbMuO5Ftid7HCkVXPN
HmqSbbic3Lq8ahslnVF0KK5U/81yivld6b1GJt6j0aUMuVWi4EcO1Oz8DoHwHzyIGrTHHsWWMiGS
ye09Nxue1RyyqL9uASkY6gM813DXFTXFdz+jHN6WkPd+niKSOIFwALeel/7toNH4DCJ5ULR4YJ/U
SXIxKAic5Aha3O2asQKK/JdXuJbfxQCLQKh/rmecDVkWGdqQWg1a6FpRTKeN2HjgAiCk0lkjGfJY
7gqNi4RzHKKgjaAPkIAhuGnbM/TIwRvDeSZktXO4FygkMoMmFjGn4U2Yi3xbtntLdAUTFQghzvL9
v3sFRxYMPujnYhRvg25kvrnVRcTKLlf2JXMivhMRKV9dFyR0eA4t+AY4ol7PNjyIw1SYTUpwjUzN
ICILEk8m+fKc3jdP3ARYcDKq7Wq1bBaoNRYa+Ke0N1AQxwlgI0pFMv4E7OUqawyTpLJX12mP/5Me
Z+cS7V1k3iRr/tPW7lapubeZXn8rBY0yrqwll4kbdLz7bPvtH9FJQ3vISm5YRNtE4xfpiSZi9Bds
H+hllT0rHcBMg9gAcq1ecRWjSnBy9sHX3WRuTyyM+3mAd5GHIGg2oIVriMVjQM+Z6bJeU6Ya4N7v
CkzlhOQlsBFqpreM6tArrarldv1EhRt/msK8uvtdfK9lprm+iVv2rPpAUX5tDxk37zy//KtSP/rt
MPTCDsywKVsb+OmG3J6604vJ/ELLPDDNKfLu6KDV5qGW9axqs6e5vhH1opuGQokEbjytPCeKwsrY
7wzVsz2VmsDof7VuKILZXGDMOliiMXN1WmHSX9wIichDNkbaA+NpB9DsuZBJilA/jr9AtE4/nQEN
5qXtyCAy7KCnBXwqceYrqwW4B0VoFibLog2qVGMt7Y2Vio0MM3uRWANJVUmNRXJ9WV0VV0GH8QCE
KgsLhzg/wIkyxqrTgRoatxT4GDBNgsV9H7P7VGbMCi9B5KjZ6LSac3iQx8ZwyYy7N/X7845cvAy4
MpETwZRQWn9xEH5hwdAL4nIBXG//BB/cMV03KZvYrouEfrgqR0TmMuMh6JkHc5LvkhOpkeZEPyhC
tMx7ZRPAsgmguIdCCqZItBkcWSdhpxwyKV894HTg/mmpKEtbrm1rn0e7728uGOhV7LoljGLX3dDp
ql1DASehtev4JXjhMD5iBEfNCdkVSlADhXgDE/BRpe2cyQzkMeDgsoetqY7wEF1KID9aHBY3O8MJ
biiMrqKcOwEKrQY7ao8CSQLRDKXhWqH1Xlq/aj5IzS7xFvNKxQzvEyrN5alCCjsJZZPgZcRf5UOm
ppAlBcHts/UXfF0g/SRD4KC9EbMvXJcqwZhDiG1FGT4LVSa48ztu5vbBsztX+zTdFC8E+PZ1YCZS
yO2xY/USRtWTEjZd18s+uRnBF0KxfWWDcERDwyLSRsp9TSyxa8cevUCXBz09YQ2K5Awy0fjRRRFS
SCnLqWx4ufcA7Z4NUIWdfRyJlZDz33DPUE7LKYjc0zCFuBG5SlXF6nViHhmAQhyDNPC+KBHZHXCY
mT+BmDi6DAtByI1bwf6Xht296tA6I7wKyvB4wpfaQc209JjcRkh72s5IBFQBNUzVPlRGPKlxRTUN
QgLLswHSe5tNBC05+dv9ij0a7wnjJ6/kRnlYtq3HWOBAxsIUkJXREAtN7nAJHBSwwMbzR8j0TOEr
EdxpV45Fa4Z/zHHjy3Rym4nbIh4NsswChhHupBGgVgRDwyN0eYWOfVrBlXAoVlQdsMkb/7frC02x
bEevnODRfOMAEsBGS50nPnrknvoaMBAdIB1dWYWz460eq9L28/l2VKE8aFqhxZ6p4MltRTABzHcO
BVXBLqQhCck3yNs5jIm6xL1+Nlbmo77IaVrjEpgABe8myAq3adWl1W4xKt2BwuxcZ7Ly7P1UAWya
4o/1UxLX+BD70ubMg/ipMTztjRF0l0GN/EF/bzxQ4tJU35lljwdwQwTEzLn3q4dAkyjciO22APSV
Mtcb3yGzkClI7BNV0Z8PFsSPOXpsFRpnQi5Su43rNqr5ipLoS8sStyqtPq+93+mIvD17l2gxBg0w
pnsQzllNEGtpuaWKlyq68pH+hmedmLeJKceusSwQx00PXR0eLaSo33iw/0geidF2BKqDpKmps3s5
obfRabs3oeLdqCZTaCfBjACZFvcmNFvSD76TKkZ86CekMmj1fpjUee4azuqP5JGd6dwj7EA6ZXYE
Q0R8rbUZyjcFlrPCCfV5Da0WKXRnpzYZHrtqOJaLMXGfQM/RBztX2jP5XHN2WdTTDX+LnW8Yuy6S
Sxzrz7dMl84PKk0EOjnboePjv1b2frxE9vqrx9HdHeYrdGtI/1MV2Zr0gcC9nnM00BeNeL9gc/EB
wWDsU3IP++go4qe2VKfm+n3S1dth9fh9J6AiEyqYH3q1lX0WOX7wESGqDdYEGOy7ZE6O1AcEgOrS
mYTkPoU3lhOnm7tQ3dqQwex+lgYUi166kTz/6aGF5Mb5zMbI5QXZJa2bMQZfRGcF4LuR94ormmdP
UKeLTJxSxjZUUwiHhq9W96e15rqMSWOjCFjG+SparlWCmfO7G/XvCSWtFlc4nkzFw+cnTAnYrbXN
lDTA1NG3N/u+twLqFglOZAWJlx3sFAsxfsZ6WC/pR2V4AcDqnxufL6deGOyENz1HrIYilFILZxEX
qED/IoX3hPbY0g2YWHjF/riCD40N3dSaeiPxMaX8RORsFVg4BkmyPU4sNsOykjzF2KWW0rSbtbHJ
lsgnQmnaSh94SZHf+oZOQo3/610fhMUwVsSZ/QiXfWStWl9sEya/JfgBGrui8kJWdDhrlWrpMCM7
8Fv/NLEHv0dpPGzBRzKsB9Yz5+tx6D+3t+y07sRgjzAaoi8s9g8rXhswhVmAMF7wdHBPx95uUaIu
yHaJkOHdMtpUB/WxLRzVcdra6iKS+w9XgNH/cD0TDYquZosGSKZL+v9eXp1shByHyV3MqliLHTNq
iRf/tNeUq7zvRJ9VLc9+KWGk+KNv5plOHdA1W/WR+031BELWN++Yn0N+w6rh1S2jZ64IfNJeGicK
MVL9fgIzNA7+FCCXJrUFLyFXtyVe0hf3uUzwrwnGRzV0ohmQm+JSL4QJTkdT36nmo73MnUCwb4Hp
eiOihzuaEdQWGBM/hooaD3z4wEDoGwrEBWDDKJSkwFeT2RUKBFVRS4oauSjgHS87q2lIT62jsHEB
T6IMV5SxOxRjGNkaoDt3TOCDW9SwmlnzhDHaQFOyR1OMYRsJUHAn6Enow1nE+1z9TTMeFF0tiW+r
il2P2Tl82m/UCL3LGg7zVAm3UFATEWVo7wISlqJ/MrLeXuimUQ5JsdjsT1doUL+edt/l+UWYzaXb
3OR7Mr68NtDRo0jpo2gBqSPRqDw0szFthhDoJxtqwuxoF/lVAFDzd1+D2zsnn+M9kNhOa0++TpRx
gSbcaRY+Em5OFBTQ28021m8U5xTg+EtSrA8rj2XVqCTLlZgwLsqB6lYVWdFzO94vl3f7oaNjoLAI
axwwATGOMagbwoyhxVFzaDat6Q7v7Tn+ywykkQxmcMG1FSK2ZKX0RhgTWh0oWoPQIBfqXHPP77Ip
PzDWC8e53DpnDRy/c6VNPNi5dOQa3dq+iTdJdENhVFFuCTnE0UdpxtypP/E2AKgGqAlr60zGnyFd
1DrguX742JKLETidS0BMaRC8C7SHjXYvl1jAI/S5MrrcYMUAhbtJoWy3MspC0aZddGn/GZ2KeRbX
O4QqkN4pAmyThmb1EMnQmx/0ODwRbwNqjModNYTOGw9zN2zFWOt+V+1d+bJ6iUS2+cypYNk1vzzk
8UFvLXRPuWgwV//KxfGop7VaHrYlx60MC0BWkzZILwVq3AlbGbxkszJgqfcmh1ReZeEkcQebb29E
npTLhiOsrU561iwAt9ydlOzMJo7Yg0hJ7cRQlOH5/ltey2NF0aRBl4jtE/nonI/4JArtwJtjU607
AJaZRZWCT9ni+cAc+iu7I9q/4iAFGbsEa83xsHQrjc1ojBJYF4fRZEZ8P3eIqKLuaUKDWU93Ommr
5/zpF8YpRSLzgjMDIesoYxpm8jN41YWjrNq7n/dkwC/aTXGmqzKk7xPMZGXTW33XfCfqDR9SKvHQ
1vKgpynE5CtgYfgSqYcuVjavmkd2uAmB4DuhByIM20m97sw59Sjv4jnbN0frefehsa8diRti+JVW
h9UnFo7TdOpDcqABIwX8zWfROUQx7bAIB0oIoCUIQRcTvf4r/JSuT0dfJncJHXjQnes+LO6aaXyC
kmUQbOLp1JZCwI+0Md8wAZoD/tIlloMRviwzBByjDNiheu6UqaW9V7MJ3mNsOJobHcT/9wCSEfV2
QzSb7oZ89xtPEec7SIio/DxAjBCcgxWD1hRFoCA/IycyG/f3AjlzztbDWNaqQn8ZERKqZILTMEYK
pMiJoydnjLcSg79+G4xF4ghkUJZ26XZYiR4XwdMxlow/TcrBx3b5TDI1wtkRdIzC+H3wSixKI85Z
kQj1O4Th77ht44uOiO/Yc1x9vlJQEJL2a0gWJzQBZPV+YjkVZ4ADbIm5eFkrdnBiBxoBwP8EGf2T
TfaqxJkn36mmU5S17b8VEq6UQcdsiPYZWFfqgS57dkNlC56GmM4pWKixIT3MffF4IUs3FJiwn3ol
ZO3aQgVRuOX3VsFYXafvMxbN1TzYQCK75Z2+kW8vB1nWeJlpDM0NXCvn/VniOvkLuB2AmHYxw3vX
qD0XY66sQwqe7LC0c+uIWslxu2VhudWSuqlPQXTj3sqzBB8tpwy4SnGTjH443KDvgOCFuOKIvEPq
Ft7y3LE+j30RF5KfghdNjD9dDzc3pjrS/G/kYHJSFN8pTQw8JXKJ1Bj2w4cms0WRfLUnbSBkHQej
jYhXwJ6X5gY6mnpQwKC98tAzaIlYRgeZ5bhpAAjx1iSpZ2/IwDDZSRDAhXx2x2Pddkpj8c50oXFD
CePptBSAQjdpFHMJ1/MA+hz1leIcqygUX92dL3pJpvG0QIaXECiGyYR9etl9LGaH0HgCs5F4oQcz
71joDK1DjVPgEojPgCUiCsGr1kRbn9/r6mip263n12sJZMFV/7Misu9qmgxagO0TD2yw/pJ6pW/4
ASsvA1KNRGUIQ/Tp0F038eT9Sca9fCQvwuEexoqXsV3uaB3LLpRosUS7Ojr3/F7tIGQMfRtV2aeP
S78Cjq28TSsMGq2kCv98+/gUk/vDmz867UtQ9Reyvz8TMTz8bRW1epntwpsieP4kq8RTmg+jJ/f/
ouXNU5exzTaGrw7WrD89iCP5wfQiptTysGTmkSs/TUa4H/ifgIFmpD1wAhIvta5u+GwyqbAzzY9K
/Bty3e43BCjhcQWcChVapb+wLQDNwXpniVGZmwghEY3ulloufuXHnrqq3eWaek3+y41T83LeZ/ec
UYL2EltkbPwRUmR2QmMMCckpR9xPTsd0cz5pbXX20eIEyEyvyJhDqM6pwhvufY5f+xUj8BKVl9M+
PLf5Npm2bX/LddSKegqKbnlP+EMKBrB/bsduP3783Q2u2LK9xEpV6JIe+LMbNpB+Ud+62cCU0PzY
8o6YfhSs04pwwS2AKsQtCBrI3EuaGpt1zjSOcTpqtKt6sL2jO0f9FZq2gOQpDQKHczcufZQzu8Tf
/YJSCUI9qeS7TKlQrIvnzUeAe883Jyv3Mg27xRv8kkSVf7PXNW01PGiCxE/COFkuYGlaPqYBV6td
9qWeoaocCWnfwH9/1ed3LOnw61elUQ+S+6LAuL9IjxE1fTFVi/CxKd3EgLN7HTyecjVNrtoKQ9Al
Dbr5WgwirrOkO2S0/LkQ2jIewFse3R9CMwvWwAyMrlx1QD9uJpQTFWp/34jtOQfBoa01MEQHIPGL
GUDhAM1sIPNEGSmAXvUb0S9xebputva1qyFMiJ7E47OKwY5WXt77mgr6JwS9WLPDmGLmq0SffTFE
mIUwF2dt3wAXAZ9O3jXHGmyBQlnnPi5IatmTdDodr7wYqKQmFfk41ubNOlmhwkqppESEZwdU/qXs
UcyY3HAqSXTdP1bP+A6/xMfgQCTgfbYZFyncJdaedsiV/ns/tF9YZnsnUdxJmuJM5C8GngMxSPIG
PLKkqGsg3cKs7UgFTvitTmtSmldHuEtoCpNtjdLLEveY1LRV5krtOI7qB6FhTwqY3URPhpldabvH
UWnoD6IAsFDaIcX5NBk8cdn8kX6zqi8XApGQwn+QB6+S3OKIMi7oNkUZP6ZflolALvlpVoK8hJqF
NWg96QiDD2ErnLLvbXXjR/8guOVhb+LC5/adUWKLThbNgqojl/s3+SV1K4rNXx4VhRXZHzpxagM0
/zsHvO7ndsM0cCaXM/eCr/gn1jnNp31XLUlaAqk6OE/41uSWnO6dq4C9Pn4gN23ZPTYIU2a2OOvl
OQiInggArSmjQiRMfGM/XV/G2b3GDeRt4mA5fcjNnn6Sy1G56KB/EdFJ29Mn0u/1S6yAlweZkg4c
VrEExc3o7476+46kcoAodySt5jTfoCCr9I2nPbKJZMYHC2Xh5833giKZN3sFNv9Uehb0DDbKq/e3
FKDyZjHPHVRJ1jjH6kaHeUVJDt3CYgCMHZGWEOK/esdMGSiyG7jL5gRycyUZMQrBEPHTrIpP1HkN
nxRtJ2u7ErPkNoXtQa3muZGUA89FyZFvVhNyZ08uKUT0xMymZNWH9sSZ/qdGjzLE9LHx3cOmi42z
2A0IgEbU99os9UVruzhmRxFbk+ehl7xmF5Dx3NAlCQv4SbYHtzW6jeFssiWB51Au/pRDo/BVmUPz
29pxr/y9a8ScoW9JTlXk6l2t/dD303zVH6KueiijHG60NdHOMNelw9yNCekJRa1Gu3AOUc2T/7bp
1FTclK8pcHZ0HglN0VKNVABd4OP+QcY4VY7Al7LO40fs/jyDFLNr5SA05MQbPt0PTqnmzErUXpdK
RYFDjuD2bxzRb7Y2iVx92ZwkzvxaxvuHJPaAI8nDkhA2dO9nL5Y5VsI8TiJ3YUylRFIQwu71nZs0
euMT25hwz2KGVsV0qd0C6NR5/SBFMaDU0gMk/MetGE12tz2/uqGiJS/ccSOe8njcomwGYdQVVR7B
FyG/zqCPZaPiqrNZs3+rCJnAaF0Rhg7qfhJM6a6n7391PokOU6ZahXH5abJVzL/uvjZqmyE7rcXS
E3P3y/1SgMn6xuZWN0wtcc7/xQhlzdThd2yzpITR3OsqxdjauY/5N8QwxZ2g7KOlxbbpBx+yPgOR
WVO7Pctleo2OOQ6Yvmy3R+sIe+9KCeNH/UdVSxSBwyzJ8g9iEiBfsviQHjKNlbrgwEXsC3CfASXW
6N23W2VufEmEvI2qUwlN9ZiffOjIBml1k3zNGkyauH3ZbVTgIrbQq8fHogJiFYPrUct2oIWqxX1a
4WeVMYJEjuwRdL390KH2LIZ0hYer7q1koGVSLdOaGpALLlhKqPWdUJl24Y7qYOB/WiZhCH5Al5ex
R2fqxEXZ1Ms3tVVGGCP5n0DjmCmSVu9BhHxZvmsvG4gnJaEotlOgGhNV44DwPXpssq35se1YR1IU
Jvm272if6CoGSy/iOkOT7EmgQMGSvlK3HIs44l2JBvyzYZAkAzYUUIqOkgN0imx2/Bx/e36nJK1c
5cANu1n02S68tbnhAppYndIgTakKhYGYNPvbK31JZgL7KSbPkBQJemAa87t1TadrP/HJJsXH8OhU
7kxqPVbvlCvJC6YEY43vTdZdCpafSgoeGAYehqbKJzNs4qcAa6J04Ok4TwKLMxGLBsrTJT7wyof4
9AhID0rXM1n6T+4yLU8p0tE6WxlKaSzb6LVFjvd58L5CNRe1wI6hRux0GmYSgKwtDO2SWuDgPpfd
zUe9wlhGyKKgtUhCObnc8joGp14pZ/ykVQRKjPcVTJt0OsY0zFEHeHIIsYbo/s0Wxd2bjtWZ+tCx
9sF4Y2SeeLtdgOKnofHefLBLDGPlZoVLQBoEWUTO9UAAa1mnE1AuQt3CrL2MOhkqSh7XMl37g6c1
7sLuz97AOFpTvWiuIu6AwcNTNSDSzTQJtx3G+69mAiVg0zsPQ8zvLaZbIcN/UvKnQASQ9hQVELqU
w2mdeQ+KJNMgh6cGQi4CE4zz7mH68FqzfE4hkKsP2cz6FZadbg/SHbErhV5VAscNSP6He0MsXhvs
mKSKaPZd0Ug2fdswE3kmTp6P0f2zPA4UopRb++eVWD+kl+AurNysFuhJf6uw9/ZlLtfPqf3mPe8E
aLu4mccBIWomufgrC4mGTPRkZtOopVuXiVKlXBGW5xeim7Moj3U5r2LJNziI70tYT13TDM986O9Q
kdpnfPnLN3uJhsW3kFgg9yjpy529x1UeLRg/stj5XdpdSbkmw9ZxEKdqjPZgfy1SQ443NYiQPINu
S0lOaA54y1X89jBCjiltxI9Xac3BWmpYSYl/7wCSowHtp/PJZs9dFbxomlf5J4Su2IFH3E/GNt18
IQDwhNx8HazpvIZxdF0JapaICAzw/Z4RV/y0o/1leMs9VP+aEjt0PbaObnPgELrky+1feG6dGct5
ndnNWCoX1RS5K98XPxFmEKInpmdiR9KiHdaSYgIAgvH/Dd3Q4NYgZ5zxBWKSoIyqgzNP/sXN45ao
BAk+/OyyNZ8Isu32tQKgzD2TVL7KGJn15aeH8JM+tmMlUI9Z6RWksGs9QfbesdpBFRtXUVLlHlgJ
6nW7EY5gz2AS8ZW/EtyLebE7hq2wSVzFE5VGrzdc54yPZ76DInAyAksI/OJ3M57MiH6Pef9QuRo2
xKmmQ6cb3xhDgsZThhq+wf/Cowh1wLd+wChYCO3S2i4M7XLB1PE1dL0O/87zZziYfL6MyAUWX335
OphXf/MaVN+dpA1NEQ89oihoTYttfU0dikZNpY/geULccOxCvdaBqoxLCRI1y+TNx1dnXP3ghLiJ
azX+WmRpFbZJ3PmL/nF0rmuLpQzGjXXOc16m69fpYa0SFSuypt5XiNUlX0Wa6xRruHVsIiANMmTl
QIg9npjqVDGUPNYVC4j0C3zJIrnO9wY5rj3M/w9juhvZVS9UNsiUFOmlJD2arBFBg1ensFvTk8i0
moX8QN8B15qpJNrbtPQg3efxcRAo5ENJbXePMVvKz/+21IP+Ra1QSFnvsCLJgdBtQ3AZ6n2kYq+F
enG/Xs3bUGLGV00sBtNe8pxgRuA3p659ALAv7KY4ekhC2Mf7q22PHcjAAwizhi94oOpd5iYyr9pT
ArQCe2ztBiGVUW3/VyREZSjD3ri+bMMlt7mtkAurUhGV/X0Ce8IMcUiTEcHnwtSsdQl/bc97c4f1
BL2hxD5IOTa3Mnz5VFcZ0Ed0/QsxUsi07RqIgk54rjqrr6bsSEiLvKcvZhHw+0Hj9gc4uB16LBrI
unmkVOA2y217uq6/znEdcy7Ac4TE/ijItpqxjv/t6VkJM3e5tX30y9kGVnjfQxBR8VZvcfh2wdBj
rR9cvCNWs0owG4qp9bo5KNgHT8e+kRl7S33hZ/aVk9A7g9S8pphaDjtioXLzY+9uhXvIDK9eOIWX
WVRL68Cm5Amk26Tt9+8XOIBRSE+v/1D/D+JI7jL5ENXSpQbdiaUcqdiXa7FqX1q4uUrN7c0REX9y
imK1Nl1LhPWBy7ylRyrwXbKtgEQXu2VXTUtKzhafe1TpA+NYVSz6hDpuvkyw1/RQq+lNnp2LVQZY
HX6L6DH8ARLJsM9ybQO21jlNnFZDLipFymSYymJ/G9ZWxaUVr8xGb0qQUcUBvm9zG5dyVQhhxheF
l2hZ4oflTGJVgku85tUsSy5Q9w8laVx4nwfulXQvMyAxH7Ka3PWp7EKaKPG6LI+4Dc9KooNRphyN
g9aZvguuJ1VsXXsuc1MEVZLxj0QZWmGfnW7WnjJ+9Lz6fQ5oBBHyOnXADiMYchRYj0U93Fmy6hhI
VSKyD+jQxFU3iXFSPrdxjZDG12fG8IRd2J4yLMHm+HeW6dZnzF6bYL7ZE2XMyv0wAZP+HUYFCTUa
frynIkekQDThP6y140OeX1uFFroa0g2Mt9khm6RKYwHBPU4TO5H72AY9SmIC/EgUDz+p5NcsTsqI
z2U2Q4rr2FqJwG1a8TUphmooL7R4ycHZOnCZIC7OmAuqNjgvSeKOmVCjeQ0DOh/RdLkx9RqUiKBJ
Am2YwFgE4Q84vIlqY+oCRjr3SafJu2LREpD/2Wuds13dFwmpIHpuxNcZP/5BjY6UtvaFN6C7WrSi
xO6+hbaR6zyobLSWLktRMXgAzHuyjwakEfGoepdYkP4gel4k6k1kvZxkCjlFod5ax7FPoqPCSxtM
v0bt2uV5DTgs8e7KLkwS6I00Ms5pQ/SoLO/TK/CMIszTIuH8O1LLLiBCQ8JMFvR1XQTp0G9gO5C0
0s1uPQfWEpVKigl/SdCQQqIPrz/XyQH/umrKI1bEU5PmZ0yUgqYM9HfFPkXCVIBQ1CX9KAiShXcl
BK7z9HAvYv8YIKeKYgaeePVy9lo0io0tOvJ0+SX6BPesnRqGfS+w3/c7gCEjlLMpYyBW+acx77Ub
CuvwA96Mygyftx5k4t9CncUN75Ws+sD6v/2MynwduErTjE3KMCBWDugYy+PJKYEX1dlEHGbrbJ3h
MXZ+T+AlqAdBjb06bW0e6OUjOivMPUHtZBgyYpehYwLHbrmH47nKMftx1OFvEieaEeDjIJZs3ONp
4dfydTz9BFIRVmoq6MZpZumYsARZufhnFHP6pp0AzeOK9XALopoICVAj5EgKm28jBBApPQynEqj7
96+z17DMJOSBzhbcU1t5DqTkqlH6sXWRMuCpyTigN2sUDa0DJhyz5N6RCO7n+oydS3SfYr4fmI2c
FENM6i3DmQL2+1z5hxMPxYY2+FDm0NkopRoRJxZhKjhhDuDJRpycrfrA0osoyR8pOHlYTbkZd/GQ
tpRN8gnPmiHWEO7CXlBLZQz6tiZBBMamBGENtlCvNtKUs5/33Nu0CAVeWoBDhTSu5CVz6hLAy1r/
KuUPrK4Yk3/v/asVtzQp0NuXJsBp4bw+97QtwPpG0bvNwdUW/rc8/d3XMfggg9IXA8vsYDF7akmg
ftSgjrbkmkzfhYJ9hud576K77R3izhiq8asxVPhleTxKDLTu5wjFxWqCWyzbCN4rXRy6UDEvcPqL
RY9SJLCcqUOekEJYDUMIuotvITsDzMRyPY5q+goMVpxEvujGxza0Q6B1QdJq8LvqEa8phKTBovPB
PLWTSPbzV0rzIfO6AobNYl7PutQx7olSWUpZRFiA1B/Lz2e3CoJn1wWbxAeeJA2RdHdSN5JWI3XU
bI7Ye+KH8HOHqgnbRmwRHvMc8/u4fxHP4AKMB0J/t8LNg2mDUVqsVlEySzNg4tJ5UX9F3asH6ve9
KBL9RuszJWY7qV2bs2mv3u+Ic0LMqSF50+eR+7wEnGUaIxustZVpXBVYOGa1nFNEErAxLnPYA6hi
qlHy5IpuMmd9mccavaiGfGWjYNPDiz6FDA+Mv7+koncKL08a2cQt0F4RAZ2Lt56+Q7QZdiExmBBV
dyD/AaY/2IElFAFJseBhGWFhYbyalDShjRwQ/zfC7k/jUK0vj8Uj21G+sEvZmtvMDuLuuSf8u0bT
3VSifptpMF4NmnjtD67bCzEpfrfoZ89GjH7WXTtkR1tTqBLdcdxqBC24Qzq6u6iURMWNshBNWl8D
snjwM6xnB2GuFuJXiUl1cIh522DYKPXH0hM+W/w1JnPQKz0qaxg5cRXTpCCD6E3Tl/OPUyInr24Z
y/G93bYjs9NPbon9FdBWxsm/JfcKe8elcwfJvrRZNtMEeG0RQgPF+0OGEtkjPVq/oMC1iLBfNrxU
9OUsLLVWR1EaudZLyNQVq0Ft1n33sfeEWl2QwaDZBIQjyYi/gzo9zNRSiZbEc2Km4KIUYq7t5SkK
6ujWTGKW8iXZ5sCkpJIqJNGDULFHHQf4Ay8z2h7IBPO9xoTdX2mL8yXA72uVyqR3ZYMEpE1dHPvE
wQ+RTLRuJxOjlmUvqqxWKGKkTiLFWcJtBS5XES6Pqt4ZHzWEsOYJD/rU9wQWTN+eZDzHoAtR+Ef5
akqAsxOnmPG7FnmCXv7szgAxen8j3IJjDDfxdq/jc2hULlXs2hGYYr9A62SlrDwa8e4P1o5CAoBw
5QCym8otmeBkdJroG1cfY32BfaSKGtXraVp9DR6NxIOKqEcULqyZtp3bFru2QtoH/EKBT/cLtgys
+OJJIBECNs6oILH5f3z38bvudtfbsXXmQ/mhpU07VZGQpnHMX8PTg/AQrGtWI7PXiLXjPzG7kwC9
GAg0VcX1fihCxkqXerhzn/tmpIfxz4ne9H8A7NGIW8RA3vJy7i52YX4NsvHt8SYrXFyn+cVOpXQk
fzKUAYa6Hc5DbcFbAEauODPCjp1Yb/IN8q7cVKbt2er3GwlQrKMxRirdAo/fdijPjp+0L6GvUJgh
nAAPLfYk7FLuBgUuQryMQ73b87TI1gayzdy6PY39Av2hLKwG/RuBhOM5xW7VqIgsIDAPlrLH8sMN
ZmtSKi6k186iKYkkVBKNXh5d0ts8Qa6ny0duVz3szzz40YB3ft8chq87Ww3hzcfaKD00HIVitAhI
+zkxJET98t42R8ktjPZS/Po9GPLp/alAhtOjGhtq2eyJw9vwB5fj5UTe2ogUf9xFo9l/sVHLpFk0
CMEC3b7GN3+Qy5bdevYNtS9rwaDhIQ2VCWmvPB/OY5RlFUfFg2gzA9we1/rosqD3a+FIaIVVf60e
Qf+7bRVV3Lmommv0e++pdVetbwWSX9hNbolh6LQdMnC92VCuF2W7E0qPjD0B7GQrdR0S11YPBLAQ
QXVmlTbGCCxipKsXEoPUdJb8rkhgFNSOMB3H9M6md5QHySCv+7hxd0b8Cg+fPQb2Ub2BAFRISB+U
qc9UxCcrRJB1mV+PDFVoObCDca+4iILGlEMct1uVECq+xJTdfOdudD4fuhRhOOSMX6wpYQGnqSAz
3qlnJYQp3wnbkfMA7I2wLHQMs+aAbeWjfF65ceJdPAYWUK8ou3ByBziSwqGnbyrZRghsDFdbywTt
faDM1+you9XcXv4LCUjAxlZtF/NYPMVceBtKdUU4wGDabJjD3ZI86GCD7fzS8ndVyDHObDkkwjiz
uFJ1cRwK6ESVxpI1y0is8grd/rGdvyOPA1ihFcsc3J7ckaDJHmdlLJZEOUjyAd1aNVIyp3LHzoXu
3ocDtZZrkbDYsm8nvcergrKWMl7agQp9oyTTA5gktui7xxrr2ZZ/B7s++ukmdssDumhBZzjLyk42
u26f2NVGEG7daEWKti5gFR8qCuqAfoq31MvIatdgUUnaBUTIiD0MgkjN5SJEjRZJWhX7C6I5V+M5
kdBvu4eNVUFlhZAjsdBxjHfxn1R69smhh3nWPKpMt1OX9FAfpr+5TNErYZX0eM5PgNHBja0y91pd
fU9VZNsNQmx4PYYQPphnmMhQH5xtdJU+mh62lML7KwPKPja/mNAl8LEHfO4JJocPjenVhHWvQFDo
6lfnzUFUsSE4IdilVX4YnYIMDnylfcMGu9cn1GNWOd2Zh55XBDlXp7yzpqgzAwhrfcLxOsXIOI00
WqjwsA5Td2HvZJgvtE+OtcJ9PlBjqQEQ3RIFqFHVRokkqLrGtqPtcXQo59FAA8eF2Q3ICJ3oIs4D
vlGI4J9bhaRNQgTr3uCs0j5wGCn1jXPcGRY0z4B5Yu2WJ+aR/Hgb6lM8fKCqX6AiaVP3vFFnBvzx
xLvsyG5RX4vGgy/TsCN9SfyhlnC8XpMkb9ClauvRBbxplPTJ5xMFPnpIngRkzquLqCFlzfQPZSgl
FW1qtF/nq4H3CHVzm/3rcjMIDfPRemOd6qpUWt3DRtWL5NEu/P19vM1h1Q8IgOKe8KQOE7EwVnU4
l32G3FtiPRBxc61OZ5qtBB2KRumfMyndz42cm7CZcjeFhlNAQeDCwWvKXJmqBn0twYH9WY9ODtlG
h2pqzTlKblqw+W/OHsQpEIdTQWtsFVXEWzyhbGKh8wYmNRsV52ejpX+qu3CKvUF+RTk1fXKbXws2
yV0YWOpff1/Xa2omC0gbUGoL6lH7Qq/yjHYjrV96nPp9C/tRcG5St9JeuG9/jGJKikUfOubZ4T+9
L75Nq1tJGMmNHdXGOSmyR9LuIQFucgB/c4OyQRsmTSbEmjVsaMuFQNJb0gzLMyOAtRW1Hdczhp4r
WuF3mJPqBRqJ2UyZ/Tx8FulsJoyBxeGUlqfn3JjHMdkpVcYhFy9LmY374YuyuUYh+Hx/s/iDbH2N
x6n+oLU8V1tHUVDc7HQ9ApzqjvYFzIVGq6BD3AkoIDqiXdabV0aqIFwUKIb9PRiouaX4O+u3WlNG
TMAid93YE2+6C1gax6rnTs0qq3cyaeN2aE2rCYqSUbvcpGq0BcBnwekMC00durcW86p++sDW7CrW
K7RdzNek90lU+LiaIF/cd4p47hOUovY+6ldsx5km+WdY9ON9alKCyPh5hKET7NXWqYcJamsCL3gO
RSvyCUZ3k1PHFFrvk/JLIIhjM2wzwURKQ/wd0xcrhYsLO5h1VREkC0NL9/kCR9jATemuc8vlBBHD
TQrIgPzT7mHgX0Q85z8xxxDVzIo0FLQ3mb9CeZ+YEALFTw9ji3B9CwFV7TCsiViBcdgK4kIcw0k+
5DdOwA4jo7ys2X2Jo3nDZ7ImcF/8nYcVFPmtfpBnQkQyWkWhYaK3jq2KtFEhGbbsqJxb/rJMxRDA
kLLfzvPWRBJ8DhlLq/iF8quqC+ZO8lBCxxvMy3Vsm6dVIxJv0NQUpkDAyY+4vIMgW+h2ipQxIUmf
Jf8/uY6nroZTRPb8kQ7qIPpUct2uJCUgc6DLPJnj1Bi0TwidsDvSymbGcYI9+TtLK9npBR5RmzMt
YH94b0DyM1t32pz5XzitEPKiZrpa8csGBMOaZC/bVDBwXQFAWg14C/3wwUSQsArS1a5asQxZTlc8
/F0e7PFv4/bE4m+c+qEFBP4lNIvuRHxVkNEj5ASzVosFrTUZXzSv1sF86h6xJcFQKVH8khqmtln4
mAfmFMscG9hbDpT5svjaPeUFrgLY/+TE55UXr9ohPiNQKopgbvqlRvzkzEjE4U4neGqXyZAYQPA+
xav/i+W3CV8I1TPZ0hszjg5NmtorrrwDG4bC+kmICHyHAr7WQM9hhtAfo/BTY+DD/NgMZRuokxvr
nRlAHSfLYoD4ClqQYwHGkIk3ljrWC0FoVvm03MoRvHm7E6mXliQTwPj2dA6mfkhSsnk1V8+ZvquJ
rv54RnVWjnB2Duz3CMt/oDl25L8FWBxOUPtwUuogiH4bYeX1U8qjLXbnEoXL/d8vEpdg6m2faooF
n7ZbQRPWGHdx93Rjp8rImpNKzUZk9kJtzayxErGF2JYxog5E04PkKxP5of6ifmJ8XAK/xhBlH44d
G9fUfvw0oLjXyJNSqR4si1duoOaE3KqsNbAIbhJ3W+x0eaOTR1Zm7TTdih7inhumEdoNOoqCgwyt
w4BLNdZr0Fynp/MEiDOUWQ6m78A3PsRbPEJCusGyVvz70H+up0lg2VJfg5u1k2GdCGZplw0rPg/v
9WDth6YYb/aRz9X/fEPZ/SzEk9tk1fGKceTtxyxs82mu1bLOGLRrcrFSUdLtVcUf1KHC2cMNYjDY
UsiW8ESRIBp+/+c04D/GUxy2D65JkESnUdR5ZKMLXoIwFPpe1Vc9Bt2ZHHyV1Jjs53f7I1TCpceV
hzRdI7ydtF9GFp3W7crBSPuVujIvFIN4AXFBl7Xet2Y+9BAIw3j5RIownlU3TDZlqqJncCzfleRX
KWdXkt04nS2ksKcPjT62jvYz5PfZFCH2mDqD/VyaPhofLlKBP+yP7VLMEhN55X1f+JAJQ+YQ1MoU
moLQOdiUiewYlaEk1DaSHoC7+BUzuXbchZEXqYh6+B3JpvSqk2HVXOjOmpjhapBejTa5EXYL+jiY
JYZfqG6dJ3OZbAHdyt5MJq5KF05fz8R/yF20nq/an+/cjrB/k5MtxxiACp3bDf6awLH55Yy2WDop
bqC//C2T5OXLRy07J/CMKkVFAEl57gjXIom9U2uMwC5aeJ2r9dvyWauloJJiVlx1leuGPyn8DChn
iYnd4TjTsRzrD5keunwCOWEV7aaZxcADL8k+sxNT7RDcPH2ZYOPwL5q3Rus2/yyFBUb2R+k5lBCi
HV0JMle+9COQp6Nrx+t2gmRy0bYuCGRzLvfC9Ors8B4BuFcm1dQ5S0tRhmv+gIm3db44iInAxyvQ
SHJ5RZUhxN+MqPVt3aomLkpVppzj//Uhqrv8dqFcLGITqv1KMiQExqGO3591bE/qOIkaj/BfyH/i
tYiefUH0rInDLy6cQatTx57u0N45wjjwsPSK/ZZTBWwWxSATa1P87bCDxKmXOVwLdPjhhahkPjnV
uhdZkQAzi4kaQcE4V5HyVB50/vCp50XsgFs5IkzbcYjTxJRA310Gg4SHczfD1RwMg2SXsxFV4aGJ
yEYr+Dg4elNf18nyjMipMXQ2YTiLir8Cj36qb0v/d6zvH5c0FRXxl3sfwfptGUOvZkqLetLjE8CT
7sw2I52zFelwNmwRyMAkNL1DvFPzd289DhB6sgE+Ek/QrifdJVUFC99q1KTi3Gcz8wrX+0pNnJ9z
jboWtruga2RxdZZKpoEQsJnVKdWatjviG1cEo55KOCNx4YTDLrBNiBXRzSDQpi792lEbBJsYZZDq
yNSM/gYAlJannqIJ/2TCgUBIaOHFDvtWnnz6a4HoaV0XTo8YKwRnxNFRLhmibb1Rwfft4VvGOsnc
7KciGsKMf+gnNN8URyhAxYHzK+vLk4qa1fDR7IK7RQ+nUkr5JvlhTebNCROa4j2MVFUn9k0m4bFE
VLH/dtHN4gr+RE4kVNTOT+Gfqltv49jNhBr4B6lCEwYp0Naujw7uI4GDoSkTV7hsp00Qf4iReYUh
nMLcbAHE4XVW63W7VwMOnxtRQcim5A26NFHUKwAUcX4MjgRYfw17INPMk/oKAuxvsh2XJnSw7UsL
+67Gj8M+Qp/emkncj8WwcD4XJt0wGykF3SteHZQ6d55r1r1D9hzTwZEwlg2mgWZFzmWNQ68T9ZhI
E3DJ4vAPPo9T2qHmlxwYmaB5HbNHXMAiM4oCzTZ1DG/kCWS7dI0HC3led1ps0luji3ekAu9wrw20
uHamug8BuiKemRLv/QpI99bW2G/6+Lf6slp/MYGzC1cDOWNhMfFNDQlo0ZDg7BTp4fStnw6+v0l8
Bm0WXmrVJ/TaSH/aeS/IX2Ylau1ZL6FqBuJN6dE5mpGQ5F3hYqKnP2WmxS1EMwbOH81r6nk1gqJU
jvowi3BAswFbTK9nUeoTstbZdixePUtlulsoXtbjuTMR2+iJdIHHR3LoVpAQcc6e/1P25Y6Whwdz
g6yfbxasUkm8UsjX8ksdPBtcMPvs2ygDRtmzxn/I+dC8JClV7/clWV9F2s8FdURxQIsMROy4PlUL
GWCqg0Cp/3P19yWXPLo8UM54m5WHn5lhEy/fDmFcd0bFyVNOkR8u8CsAScOBElH88lrSbBFnJpYz
brXpfhyS2ACeEdbVtxr/tQ0ypLW19FJayAuA+D2lLOhHd8cHTBvW0sZsvZmsvxPkY+Ub6YQSyagh
zGilPu3a/M7tTCsg1RGN2ThpJCfdmoEAuV+MaxcuY801q1GLvHCsy3/+GjR0ESu4/EPqlZrLYt3V
jhZDHkmMHuL/IuUulI1l0ujWwtl5bcN40tma2RbgcvGrnpgHeyTFOEY6lQ2jaUkkwL9/nm1I6JUE
cOijtEj0ImK3u57lTLog+vU+Ql1sl7ukRWZZVnvy4T6G5TLUEARzr2Fgb6un8l3GML0ILxvcTS46
Q+cM//6qhq3zToWYETpd5KF+TWNAYHNzoP82zn8jckrO+6aaErXuS+7SBYu8ehb9lXtjrw4FQl84
ws5E+Ovzwg9CoszjmKhYhAtljHDgM42anLzXAUjUGTigCUcQ0dESpuJ7tGdMg2gnjEBIqOYKHH6v
EFzStCh5f9l9dJ7HkPsIFMjunWyBYOqDv4mHiLlVdVPD+EdSM6bXskQ32tQeezuNgvv44BaHEJMU
faW9d/WZHunnSg9k4ioobi6mfKWZtZye5Q1ile+QPyMqSKouQr3xlt+viR86mfK31hd/zIOX4BtW
YKVKueWeWRfo4xmqx4SJmbJX/TXfGzLqfWfVxslNGnsWeLGHlCrduH3uBSJzcumN0hLtJenEUVUr
Smk0f95ZowdAMK8ExDC9ojRj2QuXG+Na9X6VG8eeQKKUH0QyCWZDLpNOeKRNqF7ywvtQwpskFp8L
4r4dplgAeNci2Af62Nmg8j7ZJ9X4ohHPQrRWdUXS2vEs2qZ+Nax7HbByt3ydZ+MWPUwyi5kAX25J
pU975mcqVdCHUytoJrVkB6Z1tezrv45+LHns4ITBN/Gar/RtZVRgUuwRFv8pExojUZOPf2QHVmk3
lHkm/vKNZELHGNHxci0F5M6A00VjEEBeQcRscHroeWmmeuxf7blU9Zg16PHVLN35zzXRvtxwyZBU
h6bhzyt3S/SG7PysiC4gkkHpK/dDVvq86ejQO3YGz2fjUld3xQpG0BW5OPYONTTMlqdpN85EO15J
444AIwTA2mQB8mambBymY4tFx7QYtqq6FnPYckyD3wBwW3Lux2DwRCAIsFv8h16mjM5jcJXH04nn
MULETzQs5TSAJy9QA92Z4qOp1WmNSZSaDaR7PJysrkrfXNxbSvDT/eYfGyMqq3sOxlpK//q7g7xT
WHjcNUoCm1uvCjXZ+YUsWRrRDS/Qlqv6iZP/0TWJR+68tTsT021ikgdfsYlBLFNEU2hkql/NVKm2
8V3eBmDEDLWZa7mLzXtjkFxoQL9Blp90qmNGV9YUeyMDe2AimllNhFtvsG8vCK+oQ8IYRIpYK2G1
K86xnWACDrzedCGgMU0g7cDqH67JyOqY8EWL4kqhxWDPmjunGXfy7dp2OZFO5BIP+WxBR51U6PTu
mR5QcjanqBJn2u5xQJIQn5GDk1XeUoNEUR0ky6KeeaeLraZnkylLsoACPZhpZj2yiVh5zA5UrY4R
fpe/lSckef1ENaU/dtT4OK5ez8tILsS0/YHBJWuyesSKk7MZ7aytd4TCwzEWAflsVVj4aSXWPxxP
Sfgxe+C3If9yk2dVwuKK5ImfN9kiJ3PYTPbGWZvYScOdTTWf7XYDZYhcvkSfpMYPgmfqTiMgpI29
aIj1zyyw+vcSwmcFIasz5DaCG1tZR3KoeSolZn0dB/EyNzxRnzjbHqItUctCmP0Amz1nXRPcXIu4
10ugZokCNhSrQl6hmqGypRB0qJZEJMajIWo1fFnDin8teHCn/v364BD0BiO7YJxZXGP0ELbjO0bV
b9Cqwf9+NnH/WRzRaHiLvEXKX1iGcj6Iac6y9v1hs12a8YTm7ngHRhNAWxnpVkS4cpfKjNL8ZZdB
Ih8j+MgLyYE+DdMfzGXl2Koa4MDOGihPIniMejuT73k3JC5KBYFC7Nq/h5FQy9J35oAtmUY+zv91
IKh1RovjtZoFOah2LVwIKF1xDfZNoM7U8NINkZONKewFQdBkHHThjSckKvi4JBqFqjgJXG4efd9d
IC7CRLGjDkirs4zRgk3Hfwupl54VlQcZKThYBhGJPMf+30iDva+/ZzTzr3T5A0UByPXCWCZJU25O
asj4zCvRpyjYwbtwciNmQEQxb+d5lia+RF9yZNoXxcfSrN6EE3rYbUoL2mF3i5CSPbIodM/bgEAd
e1JeHdwkQ7kmdiUHzGBTjK/4a0GN4roLsG7AuDNGNvuvGUVxmA78EU9pNm/oauF6yb7wPeZy/icJ
JgO/688bQnbBSUpm1HkCqrbA74zrfPQEshPKvcLVKu7P9cPlE+aoTgAnZ8u2qOT5M3C2Eyl+kYL+
pp6brWurwQfFR3SziAlyHkPjd7VJGWg+mqpC0tDy+XCf95xyBR1jaICY7C4fxHYqKPMeCSM3t3Rj
OencNC6xk1Rtc99Yb1agBfNQJJEiMWodOH0n0UgCojulfcMxbpjIFNUi41ERtnQfMf+xLc69Hi0Q
Ktdnz5zHPXrlti6KnAbIv9y0jvOodU5VBgyTapsbXpCxhvcSgdb9EixE9IdHeBr0r2eXVVKGq+gh
MubOnrnbgAF47wX+vnWUQ2bqZWGw0jx7x4EgUCPe8dmzQ+7kLwHeS3AlZeSCSr35T9ZoGJ6cmXy5
7mPKafh5YkJtegh/rIxxlVaxiNSj6QZoxq9DkqoAZz7k3jLElMAsudPrhmm+1SfU6PApY1RzziMz
mIaxHXgBCE163Q+cR/d+Y1/AKbYjZm3IDBw/NrioUgeU1UAwE/pHG/86gqRR8bVhvO/VbsV4KBQN
vJBEmUCcmrlPInzT/+CGBH6p7XvidAB+v3W4enCIBPkAMoE8Ea7+8IgvzFHLWrMsY9O8ZCRrVI8L
MJge4iMLsCjp77Oc4c2g9ysklFAOoBamaDehoRF6HVUsnzwoPJtyBf2LTKOILpkJGSCs8U7MLHMW
Hap+7z+iUd3dnUXDnaPrnK3qL/5eP0sWdoWxU/nSHpkshdsDNIi+E0+0ggINfX5D5gHlppCPR9ji
V9Uzoe50kHBTEHwETY+RJe2+QdLAxwZgSqxaqoIuyJG4qvB0Of2BfVueqiLkyERQpgstEOt+13GB
q8CsUsfzXYvVhIwFER9RyMmzc6oDaZ5DrJDWM5tYJnZcAStmXRkTKhmfjz7IQ/08xv1OeuWwceIP
CGdY+k7r5cVJorZZWuUBZWGFFouUE1XMssPEuygVnp5N+I5n71t217dR+b4PaCa9y+Gf9hjBfjAl
NgggOyTNfgX3xjdySzcdwH75YR4Uk2szBKjuNUc35lD05JksqtmEvJYWu4inLcnABJQdx25F1dBM
ldLfHBmZX8OkBIu7er+L6ZQ8vmBJTgin+n41PBKaAJZB/RTwQVhmQty0g5s1lfMZ/BTLR3UDPxDt
f96k36RoEkriFh5m+I0zpg32L7fKH/jkhLUuw0Nj5AMRQ1HxXI1kDoCOogQtVe8rPKLqSyZ30UiJ
ocVJH+oRnk7QLCidJtMa2EHft34N3L6zUDSBzO1CYXspMdGTHQRKwNEQbv0ls0rTvUdndE1vdIAM
0i10td1l+7mMThfCAQdpin6GQaiGyvqJ4atkzPppI0KSo2CRJ+FGbjjw1vlUYwpKx/G50a2dS9hC
AUCYOptV2jZBt0K1KYrMwqtwaEFzcwOdCis4oYA2OadU5to1POKMCqAC/UAoeq9+WIVrPrtQDt6T
JtUrzSDGCNlj0LQRyak1zUrR9txQPCdNR+Vvac/uGjXCBGgpOunTcosKlxN/9KNQOSo89Wu3W1ZI
C5VtQ/o6QEFa95nVhOf0koWXlyTqC8uhCJbvkiZukRRoiNNf9J81WqcU4uAk282kwHqQsc1gvdTq
/nCm2Ir6G6bbWkis3LkR/qAiWS1yTK9JW4hQsdIYXdcZNagQk1CyTg8BUUhjWLLJaGe0U/b27mhX
bQK0zyYIpxnoUiBahTlm+Fc91v9JlXx86elkUiZ3YXoE1Q/T47AilTk/SXLx9qCJg94BuIoW45XA
C+N4BwdYlyaMTun56SNuGklm2WOvdJzErhe7PpoEC0wIFlx+BWNDRLH4zpgNEIrPEf4yQxL8DUyX
ex2YHKtktK/8+Ut0dzV1w12XDZ+4k8kgI47bkcpst2rC6/4uTmaPNPnSCI3AjbS5jjhhvn+f7Quo
KqF1gy7he+f6RCL8TKJm9op5OmcUgdqcWCMnvAIRZ1TbfotdB5gPrVvc7hfi3KwnvNVaIO//A6Rm
IGD+eixAIhp7lVlB1Yup3Y71yOEdguWkaf57y6MvLzap5hKSXDK397pCbDRMrXrGmxaou9MSz5Nl
DTEzRsSJydkPwBjeSY55nJsMtO9CNTuPrbBlCkCY6CBAkyIF/WboZwYifWPlpzapo1j10vqNLIZ+
8BGlKvzjsN2HBSUj185G6ba9i5l11SisKkeFRoJ8KDn5Euh0f9oLXNTrwYAsjlhi8jCGcBH6Oymi
pXPEcprtCH0ZXAiagoRW1qn5+qE4JRaLYMzfpewakFEWLLWPglnjHphVKL4uuOz6a6pBH3IKnKzz
7tZVbV8w2hpCGMY0KdHv/RpDtE+bJf7rZfSfp1UJg/y3/e1gIo3fVNs1Rs/cNAEspEPl0nogN1Zp
bfnRzLaSD1WraHZpltP9JztFx9u05G+MdrJQ/lfimldimGUbRNrmfGFheIwSV8lOXzaodDJwz6ZF
Z0FwuWZoaA9Xxnhqx/ZTQyAdVwT/60KlMOwXArVGHIQgE4h8zq7DMExNdDPI1+/jRagtMVs5GhVu
unHNYSPlW1zWLoir9H1umx5Z6iWV06AR1cdGRQlXUa87rK0xOyqU6h/Oot1efzeEUMwFbZF0pgQn
K9Uh7lmFF6yswHpzwBOrmSrETQKc24R52v7Ks1jdbR1ggbWs+gtUwur6P7jALqQ3j2N+J8NPpr2W
Y8xjiWvQNXQrzf0r0vZp2/HSnJ54w+Ij1/XOtWXJr2XXQvPNYagLEJYmJbWvHEQA92TVYUENwqCf
ubkcu1i0DS79a/LBAWX00zYtjHPDxIoePP2K2H98IlfWpin75flF32ub/sKD5zZ3CwPfLZo+oar2
SAF+kp6qxs0pffFYwUig3lKpyhFeDVNb8g23tR2e9c+RE4pluac6hGCxciXa8BQLiejsq+82IS0g
hH9EMYa7IZNxSNdYmuU7XYoeW9tYNt4xNoD8kfKCfuTWI6nqn4U2YUboK+LtcVfO99+k54ETq8LV
0dd318YJwsCGh9ai+4u+4R9cWlbFvAnH18HJRGrvUq+WyfLKIoFu3Yf7Xr7T+pXh+8vSsIpnu7KP
NBK/wTcawd25b11um5JkETlPgwU2X7lR6d9QJTz1sdmoym05LqSN0ZBdezDQSD53P7RzWIActVa5
TXOHNIF4z1WH0gV1Ve+SPpqyi8XpIPuTqMoiScoBrW6RLn9ffmwcaVPeoRNDNTZAFwiKLKZcp/Gr
hccIbYkOJdXao0NORLZjaLAmSgYdJiqnVFWMJA0At1Tt35GJ1pVo2Jix2WKVj274ECmqHf6/B19g
pI70XuPeWd0f+oigOFreDirGOGnMPw+wWyWy4/AF6hdyGsBKWBr8lAo7n9YcwvzcKPvcxIl9W6Fk
vn7Lt+PXwcVBXWNxUbI2JBp664eDeL2A4bPu1ONSQLaytMQYP2aNlyh3YORw8p/HZMdGyXzR3Kgh
b15E0/yNoUFVAB41CzAsvWq5Xf82dx/IOnw/Hr4WEsi3XacIeNPpJ2nY8BlfXd0PzKVyA3gNECTc
05coburI3UNSpP+4ih4YgWprrWU3lwjRUG7bQFrQwUClNwEFOvuUSugjn/r0hoXYy4GrC7UUX/v0
hqSProZIO3j8TZ7h44KQgVzwK8Z0XgffzTBhGsR4K6Nsd20RtL3Ud6seXkchQfkkYR4yyLb3Ldxt
9UMIgOvmlhJpeyqWs8ho92HN4cC+iNFN0XVpKVB/VdEG3W/Hyl66lBaNyqqG2Um2bBGReYpLFHES
BJrZfozABXTTPUxMRd/W72TUrGl/083y+6Rz2qZ6UGnntEu2WPQ/Ok2E+pFFGlFKJrrVQXQrTELq
90i8x/ez3cK3Qa8J3VehwYDTVE3VsEpBlDBIfizCBlnaY0lCHOEih95sN0elEbCosItMmywmwX2L
KJRTj193Y7RiJ9NsOFJ51jrALbFaS734mJDVktPhiODM6c1x+KC/QV6qeubgXEOeYkSrmXC/L+Xn
hYQLlXBbN22DGNxlMSk9yDHKrBH5ugW3PQqH1g/GVcNfaIs2+yJLhDJxGKnhxl9W7XjX752zHETU
9mApKg7nnmDbuiwaCuc0WHjtcMYn+3L9jaXRDHEOuo5WpxX8XGB3ZhMGl60/rhqaapYbcYxRsUAr
8BfkEzBxTCri95ETSXUNcq9torQVJIAH8KWA3xMAdz1BfSQfhGO8Vr/yIUNQ0RzYOz4VMdbeBn4W
23hsVCsyivlUc0AO59W7fT37vqMItS124qVGeqMBqApaojj8Tdn6r8JS7x4SH/o+zuaOYb5sj9y+
MQvGbsbSsmi29AFGpCQecNkEuKz2IkabJ3EmZZEQjVlt08ADTB7JhtbyTJed4gPPRpPJbGJnJT5a
w/4jCFVa4xIHP6oAGbwV70t/6tLplBdNoucQQQxhwYf0T1wckG/kd2zVxcb03lZ+dD0qtW0PSuh6
9rX+NAND1SL+fgVvcBAmkFD4ueqw31kJFyv6UOceRoGaPB5fkHypI3GO+0/yP2bZUOLvGI4PqzgL
awMoWSdjnqfwTmyRefK7k2/9ofKwfyRNEV5nOvU+NgEj3dQz/ieTTJuwTl/JpOq26EKVm1JyLv1c
3CFDmfF+lVpJga7xx6Gkj6JC2oILlmAPFh+CIbyeagzYcSoja3kAez5chLaC8qUFPW8MShnyEVVL
hPazuSCxERxz2218/qYRQHcswpuEWHr7sg8L/UALvhxu8gSY/gK8kOJA7d5JVdlO3TnOFvbrApDh
yhwNnCd9D0LpRoGoDA19mulX/NMomvXHxza11kjrxQSbwTFSS35z1sFYnsfiuu2F9Po1AUB326E3
pDiZWF1nkz52P/3QXApo8VqGOLqTPkux6IQm7CNquSs5wjJiMyEPkinop8i2oD+pgt0FB4PxosjT
3BoLOeNDtcHPGAaoF6xaVBQWBksSQnvb3WlZOvHOyApW9ob+BmaKl2IW6i2wmx+6lCXMYLF7BW46
ltUD98MNnEqZX8tYCMFmqJnRwSqsRunP5XY+0vP2w20HyGYYKuVcDm9kSIyikydpUx8uXUoKD9Av
0/O5NEUOthdKT6tFBv4nPg00j5R/cggOqTFfEPZCMxNP9+RPQHe4GY5dFvgOy9KfmZAIgWAvz5VV
TTnWgWQ5oZpDnhS+VyOO/h3IF1xOGKOSM0BbmtUGl4LQX0Pd9o2wHSHnLibs7I7m7/hXYx1I6Fti
aHIq+wua3TXbt0uEVd/VYmQSanWSjfiTtTZUngdg0VBHs02HnVqHTUYoNYaYgNzyKzgSRjESGHnR
bxi90ZylmUV9qtuXLgotWTuyfDtf18C5rt7CbUauQXlhtvU9ylnvnVRNzL66QqFzG6pVRXRf0p67
YCPxmbcLYTxciIyx6Kw+Ou2VQrIorOoFtoTFORsNxV91ydrIvaCFM0cEyjvo/IYAFbJj2EaDGCn0
+ZsjajBenE/b4jUbmrNBPs231EepJpGdxfISqQNK0UQH14zTnO9bXsx1cmE7lYiT9EyFWf5/fmDR
k0nq18kbxIGdgvlpyzd+O5k/NvJKp0lTUJG9Bz1FgWOsl5UhzrZF4ml88SbmNpjQtpm1kGmyCViW
JeL09XIK+2DHs7vWSdroxeEjHbP8s+viN2C2ch0BMmUw1Ygz8tJnCjrAhDViGVUGORibH4tP3s5E
L17EI1PEtAQ+85GtzyGxJT+0OAP3pexLAj/2p6UJHrjjyAZQCz9R5T4CoppKHuzXGJ1Cjw2RNcAM
iOgGhqkQv8QbRhUbMJcEhIdMNWNO7OlZSrhF5mK6RO5Osy5l5jXNZ1XlWRU5qODLVfL8L2z/BRc5
orME4A1EkEjfcjhpghk/+JuZyfxovo1Q+aIr+H6luD2hnIOgkZVxafc+UxdQ6XzOhsdJaOViNUzo
1mgzpyq31a4vQ8ssArr0/Jizvm/dtSUNlS2VWOK/IfhNJvEkjvrMPprkKCCMjg2QmEhd4QPBnusN
Q/KTcSbIQrA3Lf0trIuznAsTrvo3hH1dT54fWJPUqvn3pEsVaiYBUTOn45duLtNPgyexa80hduH3
cxSwlkx0l2CVkwRjylXoyhfvqPn1RvmgAlIOOjHHJdfSdSqzq54rsSDgoxNw7yJilft0XOPkMLU+
KnCUyzVhnMq2uSt+QZlndV4clZvpp8arhmRuuHc3+993kfYQUQW86C8N85ryNsFL5cHadabBBe+r
UF4GejIlA7N4LA06D5T8WVzkWJlpnPXW5nyOwyXKJdfIRrgbeg9rmJt+aDqfEte57W4VjcqxlMXh
b3I+Dye+9zBwwc8gTFrj4+FhYjjrdkkq8HidI5bhDqm4P6JEdCmS3sS4+NhkPFCktUR8Y36y2CDm
hCTiUXYw2SWeZhnM5m1fYNf6uLuPbudTH5pZpm6TcbTe0nq3VlhYovZk+nGvmPoUQ98SmREqiOKB
ESHibxIvpxtQo9ZooKizCtwsdCvLBI+zuaDEhSOfVOBTmsvMch3gYW0d0jVA1m36dRgjZRyXMLi/
2gK6KusDXhKScnfGRNY4HXZi6wt7lEq9Xrsn81Sx0hYhonqUGnb8riTREph23IsxW4cc6VEGB+vd
6s5k/JqyLEJUYSILU+BU3HVJ6v3mcN7V0Za1lzvSh9/tGZrtKK5yNKFtzIKc9M+QOF8J0eoRwWoa
vyEvjY65jiHEjg2j+O+mSH42KD1qClmMtoKhGYsoZbOQClhNjO06u2dYOeZXYcYLosed+zwAuKek
OF04rI2Wz33qH1pOiXje6ULq1OEq7K6O01b6kEIHE+R5jP1uq99wCk9MYE7wcMJpHxU6FmH+n3dt
E9UzYxnhDoOaEwuu4MUq0zoO4d9Sq69Ft3OoT5pveu26TS7ODv77htEyXX9xNtselOU15+ycpFzw
JXG+0MJgO3FZbEqSZ6AAl6V+IQ4c9ANeHISQhql0UVSvhuzznoUekn9opGgEsqiON9PRW8AeRjCq
FAZ09yQDvtGx7qoiq5Rn5ptWCtLl0G95YjoWgUyxbDYEJIwXhk6RE78EpujXZTncLJ3E6uISH/Lj
LWEA1b2AMe+nTy9OPtKQluhMTD9OAYtX6l3unCIpCbc3s4L0r51VIbk3Zs18F/X5pwDPkE9v9t9m
O5YEvRD8HhZee46qyngiK9R8S03pj6bUQtHAdNaHfvxlMebILXQ3n+EY8R7WuFn0rCVjWxgBZQ2q
dYmazOisWaCwDWy36mH4oCnD3/6sf/oc139vtNCnbhwb+WLpJy8ax/DDuPdOo+U8sSWPUVVxBTEt
wSr/LnlYrm/ZhieLCwZD0I37HClGFK14aZ5w9/qLiQ1sTRJKs+1bScWGZBb1I/RcUv4FPINkFBeN
G6gXn6lKGC9Ycx8gBSQfTbR/D4foNq11eScCzEA2BPU0IwowViLDHag09vklVnYWmUA98qSyVCPB
/ENAcnhf0nqbzLkPg0N1E3AyMhEwXWNm5+L4x716rec6UXDh60LNqlisvXaALY2zUtFTQ075WGrG
ea42022qh/1/LyZwqenXz4LOhxJtZUePdas6y4o6XZCqi++z73FRJaq71Uz8y1R4SUAB19eLheXY
15OfbaI8i7RBZQlLAZk4RuMLkN3i/rSpidMhs3Yqgs+teT3OHYWqHdh1oZBrusj8LmeD+rKDrByT
i3HAjxUAh4LRkBrGT46gX/BrBoR3wbG4CxFEk8sxHHPuuDGVC1pxLDXFJawu1KfUvybZHT1YkALm
jONcLPm340fbbHMN1syrBCaz0azidoP2NBqBnQ+pnQyC5H0PINwIkJv6Lh6Nyd/vGX+x7a/2dCil
GRlOEHgWBhn7nDhScptGRioQT+fx7UKmJBMKlMq8bYOybgfJy3XUpTBNI8Md13Ip9k4eC0Nn6jTo
XPgB5LO5RM278N3AJ4HqHl3Sqp0enDygYoL3znah24V+ez4cU0FzFBbm0pEIclD5KRza0G6pU7i5
NDh9QNeBKk6xX16Ma6al3+wbBNOUkllz79h+UveRJ9cBybOa2s9xO7qcm9Yi4r6TXoCCVptxiAGR
947Ul11iU2TyWf64g/18beFDnOTyDTHHnd4tHj1ivnGSwCYtqVEE6UJNkGUNnKlAwLF462ho5EbP
9ML5W2ziw2tsdf/opt25OUC84v9YolJrja1lxXkn2kDIpdS2FMFi7GRcGkV0qdSUgccp7U25Kwgk
IhVIoyAbx7XiWxR6y8qqYBmtHl+SwTyHK6bOV6SRCbdrCMW40JdQay1bswSHOuG6rsyHaHPwrRGq
gcuicfckYPxnVS0m7uBpJE786No0NJIf3LKjKwsicwXCQC7rDKhVaWMYs7qkqmZS81pUvc83ueYB
ftHeL0Qd2gDk0hZLD57zsqVcQaze9SPYZ4c53bsrQQ8V6xE+P58peYgxNHNnu5WmdveCoeYqokhH
N7jgGwsD6h3OcS/DF6j5BpgVw5paRJgj6/ss/X5t1GGmtYEWjyqELL76jNjX6ZIXX04umMjBITuk
LSv37DOeUb8nPP0JkKoMuGzzMmQOdOLDT7aZhJL4ItLYv+Izt76b9tXBwfCNTrwjI+qmJ9zKnqbY
IT9MLuk6VBx+B7b2apBQ/exmInpvhzLXP6feNPE3qANDi1E+9vs8v5gF4o6lznD6tW2hqmf+3Ucr
6TyJ9GJ1nb15KXUf9PaXXX9ZwqJyfKQ2dNIyPtdNClZ/uMDA+8dPlio7eBtITGSurLhr5+/fJTIT
QZ5b7/KZHOGpIePtvHxHJ0qGI+Bz8iIhLo3JJfO5NHVEy6bvJHxuU3znL1J32t7tnDUWPZbdgxNZ
bnVv0kLmGjff4QxM13gsTXuhU9Hg7TIz/uWRY6SUlaxmQgTJ1ZFK7gjZIAx/jDoS4k/khD6Gf1ii
DUAXHbw5XXz5r25Wc2P/MPDFb2XcoObAajLOZWtb1jLCKwXsMQPEolZq3i8cHiqNnYqSFEmHymRc
bJeHUK0VpfSNXcbKQgEXqJPCG0h47TnkMi6ZllBExt3sKxHkqZ6FtzXGcOo2ijyL2g1Wq+eAqVqw
GQOUdyPukWLfuHdyXLY9bIMOJXSwkC15yWsN4WQAC8aBLmPju67bKsK6fJ6IudxIdN/5HHJThdVD
4yBc6uKWRetPht3VQny3a8aA1xDmxVCZosNCjrR+MaNzBvuloEJEwG+4RcVSTMd1pdmA5o681reM
BQluV3n/iF5AQvw8MU/kWqjuQPrwa83kSLe6Qs7y7QlL8mnbp74ZVmXnRHcM1NdF87SCCyFYPv8f
agxFrzjnHNYqbyMZszEFUYpEgH+jGjibSA+be/waqNE7QSolO375VbDmaNeM3Mb/lEBB98l0Wmxq
YlrkkPyRPsDSq9kB0G4RQa/SGcg1lTxZPgaKnYiwbXpf9pdIXAoPo7ExTdQfwZ2ntgUKqxUlq1DK
3l5XGvl0/7qUGfLB5L+70aQVzRLzoisSP0TzJrLZaGqKaDFn9uBJZBBYycLTACYWYENlB2pFH4DW
DynpwZSzIflAd00fPVTKolyMX7IJfiS2ldbMwN0AXP40D/O3XZ4yBIlCqGyfYKKG5MIKr04iu51o
yCoJoCRN1Yexn8UM/UEvRp3Z+RvvbO3KirKqYQEZX+Iz6CjJ9BMEKObvHz+nWq36PWgtHMgC7vPS
hXJmSB1MmoXHHi1EndpfNZSyKeVTW7pw7dPaMhsn2Ta35I+RB6q04fAb8bPrDGZfwGmnybcg3U67
zUq2CCYWpd1S5lNS6doceagnBqZE9/TzNtQzgm9lP64jPjHsYGbPQ2EMMVszruQuvSs1xaxJihxr
D5QHuAlyG9Y9dec/MNxmR2m6oCAsDWfyl9ij8xO3glFV6Wpz8W+RvnhBqsXTSrEhPl5DxTtW3ISZ
p/NX7fYcG+msvOy6KtpdJ7jlwGnS9YdsQIatamrBimhIXCwt/UUwLKtGPUZ6h7ED1M8oqv0uh1sO
sF/5pRyYROD+oGAmESLgnFlI2fApvFg5cHEF9pH9MY0Udc5vivfjRdg3pmfASLxe6q3vyhLv+C3P
BJf9hzgJfAaUcoVVRlU+6zhjnPqM/GdSA1ufiagJ7jXql0ukqTP7mj4A1JvAIxfZDgKyg7mYKWXQ
+XmMCzsvt0mppCp499F2Zut4GXhK12cx5lvcEkAi1Ul0i49UdK/Y9WcIUQ4vuHzaAjMgmWi4H5KI
mIAg+SeCIpT4bS1qdTk4dmYtAKgc34jRAczv56JCwy7/ZmglPxWYk1iHE8hnUihJICmMwKSy0Zoq
hmiOqjDSg/Etqj068dFXSlT5rZXmle6P6cJLywEzHU1VSdlWFQjrkg/kEGQJ+dJ1zLMNzuYIxZ4d
gIfmTNUKXcEKZlCasyuk7+7skQWI+POcQCKRkYOJWM0cLkBKThxmaEit/T6MYS2sBANRYa7eESw0
YAhYGTQFpoojiHL0w1FiLrwh5vzB6XeX39IsjfC/7Pb9X+unbvogX12fDT9RIby3AcxaG3ZiMJO9
o340oNMQ2soWgLRNbOJzy7UGr0MQXrMvsYF/JM70iLUzU0rbyl4vM6ZHLpWbY7oI8juHW0Dj5tMV
Y6NWP/f7NsnzqXJwwM4siarthjPCfxxTz1dTGegtcCC7YzRDBIY3u+P0Hsdo4jGgPH1dTv6kVJ3v
7Ck8EQY7pRtRVLynqatuJgVSts+RKRQ+KK7bRC15KWP2lyZiCRLzZ4uv+uDvHy903fq2I56ckCHV
j3iCEK9uBKUSUi2amD4NwETNMdlIofmjF0j+01R06aTE9XmJF2q6hkjfBvCtr8H0n18Il3Wa+9iV
dyoNPI5l5Oa0KbkpWGyAbuJYBlnDxFw/4AOTg0ND7AF+/wQlCaK/1oodmk57p3K73pL2gsrTlb+S
ScvXvtfiyGPvcve2iMXBDiA6AnCc2oUdntQ6275u20PY/Gc0kUfUK2H3bm85m+nxzMTJqhfWWEEj
alyo8Y2btDaM/FNpEvL2UKmUKiDFP2toYYC+PkgvfSogqE/8Olpc6+9Ay1UQmCHSIhQolx9opJkS
OB1iYq47SE/yRqfJaU7i3mtyx7XewMbtahj/IkIzmk6FsakbISoH9LaV7gtNgRdQeIMZdO/kOYS4
53L60JjfY/CPAPz4Tj5r3NgEF+PVdiVpBGS1R7vHZzaKaQ2PMpcITbxVyeyHEmobUFIXeKUiuEgI
8fwHnQQsm8c7fwuQnMzMfzkeu84xCrbs1266QEFzFV9S1yUVUwYh6u2OcGKt7YcwGs0sg/0MvEoI
dXysOZVa6gkvP51rVKGCDSTHsYEFK94eikjZ3+QNz7YIBcALThyVz86ODz/e9FhR5n2wHE32WnYs
PZciWx/SZ3UXeDImB8ev/fGL/Auw7Uz3MEkMl5WtKagbwhCCr7WXYlhAesnCGEZCOU/dd2AJcqHd
H6loj1v9t/pyZY0tysVFaegMlgaSO9QwyvfHeRXaCW2BY1huZz+VzsUv2L0U5alCSktRYrzvP2K1
Up0Mlz9qioavIWW9MiH0pbJP6Oergpk0tNJJJ/iOCSyDOIr+K1L1Qz7ADpJJtO38jC8/oLoOoxPK
q+C43ftQ8TgteHHvLT7aagrIhOQaS/CYjz/S1RdRYtxK1XpCJfyXhfsQIoI9znoymqr9mG/6JBCr
PrEcAPwdHPdw4mA1GYlD2pK6p2LQLdQef6/h8XwItrBv24QjU9YETkZdWisFYUt2XoaI8kAcrvxX
DIrJpeH9a197D3iKdHczGLXNf94CLnrFeeb0Q20PnHUmNyCVcdApyP4tCCFI/8U3lvAdJS8T7qkI
942PXmF3BIne2igq3fCMfrE2ZaP8XY1iP0hggm2nzSrApclJSj0/P0FR1setkRvYgjz3sL5xUQRY
AKt1X4bj4fZlGfBumOOI3/7AyRm++e9KynE62UiESIQn+wtVz+1pGX4xhHieb2aNMj0yh7rHcth4
uZh81nN5NsczWUk9gCHOJPtR4RvjLvRbHgpmI8anp6Ju164MbAhjzkpOKptOYz8tYTxuyG+YoJOB
vNidAdN0sy8JGeLJWCus/TFFBvHZXp6lrt41o031DlyMmyFVyiS/NpaG9R98uh1WpMk0XGrOCcLU
IEG3Oe4G9Viynr6H1Fql+r5HkLFna/k2RSJuz8GZgUtJAVMAXdoc5BJAP3eyX1BOie6Y4rI/hy4k
RJVstHsQ3TFUBp/oBPX9TbU5M99tdGQEfBHmtAvKQjlv1K3v3VY0TptDS1Oz6/RIwypAb3dWhBjN
Oh4y5eY47yRKYUvndW2eikX8QS2MxHeZoXl6Q5UZFZzsRoUaVAfYIR0C4ftw5U53NzawDajQmAyW
j+08Tp3ii9f7xA/S9ofEOWU+1eokW8HFLZbooJEU05gSqXJFKTRNG0/CsMhnPJNUcSu/coeWdNk4
ztCbzePL7pqeXWPRy/+q9DfH9Kzj1eonvc786JMlA0FHnUda4rktPmpdFuNCwVQZzu0pAr4ktZGa
LOtAHhUsWQyqAT7+CbM2kf/ZQBIBj0+jWPeWKSPjgGYJQj2UNWnCDkRcru+X5VKKx5X20FYXFc1W
wyCXiKC7RPD4VXhYAQMRzm2VpToeVxDgwX+QqxD0uuhwQh7M7uNJjhVeWIjULyj5QAtYhUNDTCna
ivBKg8r31cKtJkcPvVcfkagFy0UwOcwceZfLifYpiJSgCSTloD4yqShhpP8g7GpwO32DmcB1eED6
KkkkXIiez5hczRmr8P8yTPvyJUb1w2Hs25CL+cTIe3hVt2op9gXiNEqGvv0sZ9D+RegZYLbZpcAV
P6CPKiTpF0i2GRxqTaNy0KHtkOhRGfWDnL958lj6z7Rae/VFdzW/CTTOdfaqqZCaZVILd1E2fRee
SlQ2OLHnb9qCGoE18ZpUDBtsKPJWGq7m66I7DHXLQnujVUBAYPeKTBr14sTIQJeS5EqYGlbEdRHu
VRzEmFxtoPbDckH7eG9gjxvlLFtfdy4vQa55jB/SFqf/LaOsi0iQ6vtVVlQmjMCB4eU7qeyc5Fan
mZelmuv5mDH0H6YJujVw2VpqKs/JAHy2Y7vhvg3LoQFocLkErIxO1R2Mw65lVxQ9TUFP1LiWt/vh
vzMKxzkFOzBSftZdXuM5IUdAYsJptkza6SnjA5uXiTp9N2H8eOc09AgAV4mYlYOZceB93FzVhhFE
fCgV9eqV29NF/wtUcUzvXMTBszVMf1wzPAXjmSap/u49rGsd2BnJFVfEm7+lD7lW1sHCtoBvpC1+
Bd1MRaPAC2lkHVOWlCwLms4x8PCXdcFP7aNo8zWOrAHvsZNOPjRV3FNJWjgLe0OKen9FLLEKOTAM
81rx21AQ4scqisvQHX0FeLXl4dctBHl0He5FvY/BVOp8lUgCNla4UI39qgj5azRAVUqFF+Hj3svR
t3xnjxP9VtoVUF8f8FAfJm08cAvSpxssobxK0y+i0SiCoFrn2do6Rym4q5RrfX4xMRwuA0D7Bi8Z
+6bLis7/m4iggp7GChq/PE5EdlSwC8QBdOmaclJzmHiOtoft6EtKVC4R3lAAeQNbjMNzg9yoXrM6
FxqwWyCE+u1GZh8+arQKYaW+aQd2j/UaiCBmiXeDXvWXWZDDAejtGfx3PAfvuW0osiLpoFC1KFpw
72DUuUaMZehYpUAqaPP8ZO+ThtusI80FolSLf980UaOgXmdysyvQRvJDF9lIiZOrn693b3pikpgR
h22MLzPKHd4ZUIBy0m463FrIu2W8ol4w4Q1nwEWZ4+Np2A5tWsY0g0RIyH3hWhRG63rxsckizNjK
23/oUl/VbMTau4qYwPvmBb/+Gq/rSQ0Bq8G+JJsj93MtJ7A4BuyTqAz6VOjiXYtLKI3Qf6Snr+a8
1mLX9sPqEZiKx7YFfkbBTrYiVSmVmizrTZYYoC1Wx9e6PlhJnt55sZ3WEhgQX/WaU01j1mjR0Tjy
ZRb0OCmv3Jaw+9tsBNZsTaL+LMOUr5sxwKijlNxy5cUd5pplJHpP2hY/lqHmEJYAmbazVfvGjK4M
RgSGxY5CVoQB8OU2fyOsoVo38kw4cAhzNCMs0zw2/0tSTkoKHGSlmXkJyHS7viqrLwOG0dQaEgsh
2NN3z5iVsamWlqhc7BeIbPGSuO9L8Ym3jk1hTmYjedEIw1xVmR6XuVakEkYtp7b8aTtLUjjV5fEQ
bNwi4vh8DWjboV8DG/apdWjHTm3wK3JrMTjH+9gNnhDd0H/UJdBg3GYGRVz9o99j3AWfozGU/it3
r4n+d3TZzfDJNNT9/LwOHUqxiKh1ohPZlK3SffF8ZJHIaZq+2dAiTXfZLZ0yNaIeByngnQUtcSuE
coaglgWMDsjC7YOq2A1LNAD9IZW3zuAhD66VwN6Gsytw2dL3m3Awil92aQFWeMtKFPRRtYf8ahKA
1MA9XbWU1rvm71yvgPh+6VRhQIvunW0LbJKpPd3epiGtAU0MQGlhEjOB7BWGRfZSMi7xFhylaSyy
yKyO2w44xZCHKaq70ne0jB9X7XwfQn4y8FeOZmXtydUhjPNYTwLL19isys5UrTbJeeQ7okHEcnxf
QezxpYmUCetJSJX/ShTSEXCE1Z8l7eOx1NLwUNNHc96xEpYDhbmM4WcqOKl56Y4LUeUMa87+LQs/
ZidRyVTaZR6yvPrLZ/2S5ZGkb43TPu6wWWUdeGrK7HvtA+pmH4cQ2qOexBafQw3tVzWZyLuNGwaJ
xS0ly2wjv+108+ZKjUn6ulZ1T6g7c8h0vEtihE5qOz6EpXPVfDdiQa0axkc155ZMR7+mJpI1w0Sh
X8wXR42AMX7AuM2zA/EU1+ZSX3GGiGzrFyjJM4zCfdaPdIGzTEKo0aXPV+rNuP8O2R+eRee6w6aE
NHLJ1ee2Gmqrt/GwGU16Os+ycveOBhb25ZbYw8mBZCA+2xj1z/y6T5cnNqzYzFhBjhdIiB1LfnVR
A0MZ8FA1T4P9/nfWhfjfInBtpGlpxcLqRORT9rY0pARNuYlwKbFH7M5oI8P8yvfQjIzgqEd64t52
dFH8Q946j6Thexnp6VWQAPL4tNDAQlFOmE4yz2Foj3hT01HZQgy8wbY/arh8NnOFiihQMwvH7m8V
5PilSoUcz+TmnEqnEgwAV6rLTMx3NW0ujROA+lsFumSkGuKH7ppOb3gsbHd0AUMZj+Znl30IXDiY
FxELZJAsFWIBvnNqlUFIl7SOujc4VnZG51gzTJzAnOZLqMQvgj+azqoMIr96ZNEuwZJFFVQHwvl2
bfpJ9JZEzVFNUhfypbTeeo+zd+7hhlDMhHUt684zjK4lZVZMnJK0keWUJFWohl3CZI2YEqKF2SXa
xhLgm8keoOwUKvMR0KwzPfZcGzpeU95pWeUxp5dUbE2soXfrk16JOFT++ifTmWtNgO9/kw6EUH9U
PWbT97DyK0caBdfXVrkRDREL82YJ8rnpRU8xFEsbd3yB64tc0j9/2HPW3IUsc1/2z7Qh2NlbQ52L
YXf6JhdFoyjirmIhXrCEAyuBL1CTD1+4wAE5pJHrBx+Ghg42oSLoUM/IqIwwmcc4BhFVEZuSJnaN
ls09lCivoIDH1cGBP41LL16P01F9n6OKsB64GATUOwTny5CRPL1d6AOtv+gcWbICqHsrnavXb3WX
nJwaMbZDa0uaDRfhV2txQU45rDqMiTz8+dQP2FmCFDk1z5hsX7rgldnTKAxk4t9R81giwl/Hh20z
rPDfZL8+2Iyo0BTWVw0HTXAibY/YxruAKugSxC1BHDCeh9a4krLFEJtvkXEaMQAq4fuakUchstql
uFQIfGmiTTLeux3doY+4LmI536jesx3uwdUlCBSzA1YJZRP6zFrUNKV6VqRVTYXboGtz5SJ6Gvtz
p+7S4hWTnsgAivZW2QJuT0gs52bFOC245qPcpDEloif8E53sjZipF61OmPZyga0rrJ4GAfWLjY4u
GyoBi4N5nAJbN17cEMdXrBfUAkO9Kqdo18rJlFq8JTHfJ9ZT7UFQqTPjqyaRr3QpjjZCFVejPh6J
J8gtgKCfSHK8xoX7HZO1yNChg9+xfxUfFkeSmMWQNX1ByY0WDJ8oP3YwuOXOECvDosS3tRbUgbYu
smX/RtZEJxjc92M6RQJWcoR5s+Pqmvnktmi8ZgzC7MUTvpLxdJiXBUOnqKW9GjVweK0/s9Xb+AI1
d8ipcBBtYhjclARvNFv9uPfpPsKyl01InB7VRFlIX69XLPwPpOr9Euy+rp4u0vp0VolU7bJcKkja
N6+Pe2/ITFlZk7QYDdPv3waLNNaZD2smhMTePoPuroI1CWvFtEFw8KNhBdJ3IPlkj53yWsBB0TWa
tXo3P08NXo3S95XcF7ePfDqwxdfljUxFQpzrJO82iTvmBLa1og3ncwTOO/Am0ehLMpYtSbY5yJaA
Y4uTXZKfCDn/xbQRYstzZioormDARNdymHw2vjmaqQCLaZ5jY8H/ibSwFvf/S1Af/Ba+JOvLFRVS
2l4PHjMtSBCzERTPZr6R60RSjmjfvWKdrtKCeCRNqQr01Nzuo9GC/KleORBmQdQrXj/OSVnTBtd2
bB5A1aWzqayzi576R2C45WFhI0GSti9h1BZMSuEE+Z1uw8cxeOwGhU06ejLaxPFC8fyZLbVSfpXm
29OQtK9nHFn43TiAWG9ZWxx1tBt4jtAl9aQs+5BvAKCz5gkALtgU6t8QUImnF7T3vhCGzlimSMhG
Svl/xIFJOjpFNdfbJuvk1ds38eJcROl0/zun5uWIpJSTnvx3wq17PL6h4lzqVkudXb5igdOHBKjJ
Hijm82vCHf2y1Tq0HHsZqPJ2lzm7JQDfVIhD+A3JuD+Z9joPRuZBulWXTjwxQdcBtBecoT5Bszxx
NRQzWc3542OEPV2zT/9G2qVwu947z92ls3RWfU3RHCRGhPKzPHjmDXuuSvPpu7Ql4UAFnUzBONiC
kuf17YlhKWmR8X3vynFo1ilp0c5OTiDS6H7LznVkX16PHZTtbqCDG9FwOJvri2cxtG62OD7XSB2u
MuqI26+witYUfR7dW1+N6jdhEgOeY1e9KvLEMXDIulrwKWSoxb0jqWLgOnK0lbmq0j061QyzTtJd
aFCr39Q/VHj0p4M71lMNqLR5tPRyCl8E/49IkUiUkH96fU2ghWSBLL6STNLek1VTPCjRYF0yIQjl
vD1HUEBsT1keAoVbPdTUf2F6xaKvJh65g4lERQmR35gq2xBh/HcepxllZAiX1irJp9ZGXFxjgQi/
hp0yiZ7xMYmFNIIWvq3hoYsH0yijax834kS5CXX9go43uacHQslBDp9sMsdwGIkE7XLPylvfGcvP
D5gWIKIByUGjIJBqqSGuZk9crWAq9CxNdeDNMlh2NGJq21Y7kL+7jeEci6Ov3wQEVToejJ3b6lkX
E/vJ0K4kIbJFONxsR8wNV7JCOuP8hNNVZe6xrD9rzJs8glrDwd89n1+ZLVJRTKcdyoZGPcjGVa2q
2i46crKVo6xCLmNNEir+2e/qFrD3DEHRh39dcak7WAXHwujM4ckqhtU11dULj4T9Ye84JqNZNZzX
tF18TnM9hQtNi2W0b77Ql0YuJETxgkX6tJC60m0F6sl7TzlRegvSQC88ynvAcZN0vI5pJ72t3IIk
r+ekEQ+y5Bxp2tt2+gWbbpqliErOHgdlTaiym8MT4hkWQOjlOzRL1b/Wz30WVLKAKuEsw66YL4KY
85r3apIJ1ZQFuApYjwDIIDvLH4lXGaiC0jkUNH3o1IFx37qRAQQaXuQIbslKRM57LQ900tnYuU36
sMZS4puRGdMhoPe08xhqNCgL9fwidG/8mTYj9TM459cldYrT3hSz+lK+cBDDLi6tq4GfWo2xCPHu
C+mVT4zVEaztv5HQGPnF01ar8F0hsIFneFY8yS/ZMVAOx6CBfDatYyqSEtwtbNShFRVkwYbsEFwr
V+niGIypWiks5Q/hyUCu5vmll/MyVWG6dxybdhQaB+mbNwGXZFT0hyE2pUjiIU1oHzm4SUVpeQcY
Y6Tx0wpCNVcCf5klZ2vTeTzkwIag5K10BaZ/PE5O2BWGiYjIJEhG+5DmSC68Lon3lOfuhOcmlnEC
FSbTJkif79CEiwud9J9Mk0l9V1adHVfZWzKLGSuCX3ripeXYvPgPDSX57pYag7hedE5+HExg6Yy1
/pFN9jKXYfjzYLKrvWIi1yMu4Ih13etQpANIA/Ff3wU8MW4LULAEda1iMnXuvk+K4HFZ7VmKlhS8
xD8eFPJBG1MJU0RJ+myFnZOudjBjI5ci+SWcTbUVDKyV4eW16uh3m293qJ7HSCbuqNp3Y4kFj5RY
A55AOVwem68bOTHZNKNyLhi4nIidahBMloWqvml89LTsRUdJy8ErRBpvlCPVDSyO338u4Yfclq35
chFut6VcRIC+dDZe1RI5R9eq5K5GxLVgRPbz/fROCxijPHNakjtrsLeMnt+vHMNjMEYHsX/Xj22J
8F5aiOmtooJTzpFCRE7WE5oH66jRE5CwLWgWy0bUJ+O09POqRi48p+/lZLIKFLsfckKS9OpMylOK
a3FeDSqPTVaLq+hRHyMCxXhIznq2JtPZlenCwFkZHxHORv8fVP+I0Hc0uv6TQhbXYMeWuPuu5Ce/
9eLUG174rpEh2TYr/CIAQ43R47Yj90C0oS/l0eTPz1kHlZSmmzT6qUkaV5qvQ/821Q3M4+0FTzUO
1zGTqk9PSlO23oCniWV9dMfRz7QLuGBX0B8i9xeTPgwsk9jiqpTGZtOAqohYi5x9NSmqeiprz/BV
sWV74mRdcQ4WEyCILfC4qAOVzpei76WoXaW3Cmn+kwr9rEHGwCSF09yAY9oHm7cZUQVmJqHCrATp
9LmiQP/ocXQEjLDOAyH/cn1o6VmQAf+0/wjLjRhEcbonvNuk27JF6hFzOZ+lQ9xM+xEKCImdILPB
CAm2Z6qG4pAkhfmDS34+oSirR3xJifETh2FP1Qjxc24E9KvuFMkRMgJd7iXmy8hNoJjeaMcpO3R9
9YBceXOot7WCaxpTXaXpHj1aavfjWlVKsNE0OISrWMBMSfBZoe9a29UexwFNvraY7EuUKUqqYVyj
D8oPD4vN/3w6CMXiow6TnctNMYM/uYmCULroMRPYJ6fhuzBn2iSpNP66AdoL06JI+VcfpFZBc2Yf
An+ahEqseN3L3PacrHNNthK8/XrCDmY7icFBg9NLmEtf10cLSIxrS1olqwW1EkdH6foXsaUQb0ua
4ymnSyzkp1RqajsIhuS3PzEd1/DIFFdezsQBxZjzh7ebuf4AVCi7LgouYu5lHY/ZJHFfTg6LtTqq
JWUg4EtGfYTzA7EN1gSqOU/0EDrCLG1kBl/+0EfiYGeDjd9l51tQeN2zGgKMrJk5WHVPCAiJoMxi
Wm82JITcAy4BsudwQ/jNDDt9Yrk2BqrODATvtUjvRsBfeDz0jqkjiHTNjDiF4Kk7AEnCEr49Jw+y
y7eWMsnnDx//IscK8/QksL66VT4g1clfNZjMJ+ueoNc0dWDVzWXru7RpMcOGeXfZ8QsU9yBrtreC
3pxRJRwIQnN03NB4WlzYmieJYY9KqN16UpzM2exXPjAWkvnSBXumzhAr9cTgAYLUz7vOGa6JJb7B
uCoNqzKUkdFk80WSx57+9o/adGu9Mbpv3QfA71rPWJjTVhLqftWBhA8XRM/ksTFOHObPHaGvIouU
0Xsl8m+I2eHu1cD5W07kGakMzwHHj6i8g8AGBvweAOlDDgk8/37NsV7KuGsLwdYWpCYja1I+QC2X
GDre1ip2M+RoUABZ12woOpTWmPg7uZwoCoC9OUV7l35pYanh78K6mWKODCybk0vd5ZaLgxCNKIZ5
S9gA0TGeIkKKTrIFxgsrC3gf3w8HJ3cG8ZsqoP5HdalsKhB0mCYgvkdAV8uKijtEaDZDJrg18phx
JdQ9wpCFSVWRfnA6SDbBlyT2Ykj9NzNtIwhzywgPavWRxyozlpZMZuQUer95Su9+5nhH219AmDJd
ztyMALehRysVzKcPdb7AFEmPbItsqHBFZnCLaVBrgcpZ50ZTUAcaNxkM+/SwEqoODBdCHXMbODY7
C9haTREft9MnJuaKaPFOJp7PVlLBQl8Ms88EiJhS+KeUDwLUsApwp/mHuDNhfM0uY8VgCTRAHD3q
6VWo0pOauEhHWWDDHqCbilaXSOjBnCRvh4dfmqu8S2R0KBi7ofOqFs2Tv4IjhgdlNKkA7mogogVl
1VDOuC6+RYqn9tb/TWAn2ZeELgioIMVkl/TsVFUeV4zsR1nRCaH2e2ZRrunasGAwoPYbYIhk9ErO
YrOufJcHztHyoYTF1f9OQ1RP/PMs6TUMf4rQ65Ui3DLKFp3SDrOR7VkoCn07B5FUr0lu7ROW4JVZ
suqs8YeMqc87EX6FVgVzdaWRSW1zKwYHXzHwd78b7oYLM5jscD1tfIPBmiqcdBL3EO7RHLQ4mDne
AlVDwWlxJQUhZG+fxED20xprq6v0kCr37IQv7kr3/Qq7J/scCbwAduQC5R+wTxfaTFmk3A/p6oTL
nS9FpBMqyrWJ28spQLFrPGv0bnva0WyE3YvwKjiofLqJeLs5Rqze0pQNxv/cd29d58fA+sRVl0W6
cSkDPSVl9JXD5aifnTcTG7wIIIgw9xDPoHK3F8kDQwO2dyVig+5NlysFFtRijxpTLvzIZLuCzbZ5
UatwmfHEEgYTmLhZHKB6MLmDQNIm9YYqrsGObzFCPZ0WT4OJoEs2weJMD3EJuxbUS6wLnd50hlR7
qZcmlv5Z/0A1bmhQi6ZlPJJsQwekO/ci4Nq1+OTEDf8QTtc1CH6UBeLGFmn03Dd1s1CDJ+sMw+oZ
o8nM1CdI/LNl3scep883qm1R4gKzK2jJLqR3WOOXRSIYHGvk9n/DjJvZwqfxz0U5F89FPZDWaSwB
ewsZoz6dhT6PshY8ON4MXLxMr6fFwxZlaIkWC19PyN+Mnt8zTV78re4Md/FPMawJa0UfvRu6935l
GdpFhhi6jw+oNLiwvxmeMyxqt1M8U2s8SaxNuZIfLBIRVd+TyuXXcWxot7hBDtfrToJ2ho3b+8GX
6a7VfTYD/82cymCsiPJu2k4Jkf0nnAGW1N3swNEd7UfCMbdC/xYGNKt3+HAaNxNz5Bblj0E0vbEy
adxGx+ZtAo6kC2O/3ozNu5FImm3PLEG07FHwQeVIuF/mRTaEpDmOB/zQ++Amd4kGN71ytV6jDaWL
KDIZU68fCmkO8Ot2Tvygs4tgM/ZM0JOIwt6zgz4HsNM7WDvlF8Znxv47kvIgUwrkiqpdxFS2LkQZ
dvIO1QYuO24NoT2isV5ZQvXOmKsVW816DlDwBXG2EnAakcTLj5dK3g89hetrMSjXG32djiyDCVfc
B4wBEGZVtuFggWbqtuiYIYaBl/u211jiMNur7zhi/uEFo3AkBbx/CeVsZ1B1VDCVX5S9RpsLZHm7
tfivB5330cREZXcnuymtZDIHqRNEaJ5EYUP7ifQOwBY3PVZL2SV78Rzcm9hzu7P7PKV/KlPqTU1b
HlM3VY0SJfS2QqGtkvHxhl875/U6SEwYaMrhDTFo8eQhqfsWonCgEHlHbazKVdFFT+sT0+WE4x6I
YDDdMGviPYxu2ORnLx4jykccZilwGo4h6ZctOaejkOKiIN7twkUyFOGycFgfl/MlJ7THCsVW5ifv
cOhQXIZluS/wAv/IM7LztrpfMHGHKS88KRQiymrBQEjPYkVAeOAGAAHOSqotRZ0ar1YcyEsa+gYD
Zm8oOS4F8SdK56R7jsmgEGP27U8J2SXOR+kO2FrzV/EKogrqly1z8Usgdu7DhUQ0c8QV+CNmTjg8
BuWL73MaegWy85oYbFhggNI5l6WUcSoyxWL9l3h3U+w4erieSUAyxn61ppmm3IRXWPJADO8HVIIE
WprYQAnryK3CtCUQSq652Hx3Z76PPQJnSeFssmLdZbGmviyksnQa8BR5P/SeUecGC2p5+1S+GKdv
qA5NiUMziS99dRPl0kb0CTprm1iAZJCz4YNJ944hgdasPt3EvpIOwozDH6D2D7MwMDN20HDDvSZz
V1/35JrEXE1W9rl9+eEni5sKHG+2ZZHRv3By9IZXOQKQXW5i6s+FlZQpM2HszTLS7lKvNWHcHr2s
qRhaJS1OB59im5YvdDL+2osmoULI3qOAvxFM7oTqjLvBfdHrF0U/xXDX1ADknXxcNDYQJONSuEhS
vEjSoagueApJM8TOZLHeE+PKd4D7u3Mt/qK89NcY8ULP+VYkuhEeL7LpaueNCRJ0Mq33SA4AjIPk
RiRxzvziILnPNhqN1owQwa1Qo8hyv7Bo0blSDgprgrhv+fBfT5fNFFUBT3Y5vkT+/BdeNZnLcSh/
za3oPyqsAlmr/eBi0MlwzbRurgwUKQDtoRTuxgSbGPY6bGgLPRkjskUPSHGi/uqkjPjFIqRQpz9w
2O65O8aVOvVFlzR0OKuv3XUA6M0bxDznX8a3uJNr228osCm6s8VAMULVY7q9Fb7CJaIURv9CwAzI
szIg8u45ZGhqOrHidELf6xnOkdfThoiBAeHKE+kWRfs1G+3Dhr2OeyNA31e2iIILNR5QopE/5F82
HiJjxgZAecrmUoDnEv4gkCLXWH9x/lOedRMQHCqGrMhLjtMsmIEGs708+NP60Wrn997JFelrtqSr
zwLpILfv5TT48S2Utd7Smn8GSSE5kbVfq8ca7cLm6YZFxsykS/5U7iK1nemhOPorjTJcspi1qCSr
ll99ZQlxxT2q4B7+/Zm2FMrwMX9aFjHLMZMSVokpwCtGTK6m4GhdydfZiUpkcCko15WKL0Od2iOK
/vH3DOI656Rv7sciAfJXWix3pxaFg38obCK4avQHH/7tUW7PdEZVp773Z685EVP0bkoyudRNVkVm
DvhfhSfdTVFVcUPzsn0B5FslRsVk/mO3Y3tcT5AiKdOfQRvKyaI9EVUmoyL/b7LlQ4fu0t4v/2qh
N8pklcKBGwFpMQGN9eOslGl2hX/kJItWZ91dhcBLtzg+7EiB9gdMxvNtfWJQ0gVoB4ZM2NqUzJe9
qaGtfvdmXJg5eSmA+/KV/VKramoobG2nwF8gQ4lclimxQQ2KXv+rlGnO/l0fSJDhCStIXvydhpFo
Cr8/M1IO2h7eOgr8RWTa9ueilsAnBj6BGiwGMbFHjlpkxorqHu/8rWmraQ0E/AUVBTelD4qjdQhj
Q0qP7OW4inh2RZ9nxdGZR7QTSROHWmyr+UYNjaNjSFoNHIumTth8UsCDvWOXxWofehUqzNO/p0o2
ndlpIZOZ+zrbZ0TMY3niDIdLw76kmdCUKoBIKDNn1TKWwCaUtcfMcGSz7i52y9SzAjQ3SztKouIp
Fago9rcei+XTlkbwjR0jGlddFE2YCaf/KzqKhek2hHZqEl/TIqEvGXF7/AFTMR2UKsy64HtDQXHW
sR7JA2nqXtbUKgTvTWqQi0iBFATZ4KYCnZK7DlPloCTZ9bxmq4U1lNcgUI+IKsdqfwAx/XrGnXvE
pbBQNLVE4RLjUkXx32OaBjO19gmz5ICw5rU45DIbu4cwkjzk/7E94Qm17p04kMpPxyZBD3ffkV6r
Jh04aKvMbU9eRWFNT5JtP7KWVePcwXY8ZHV6om60whVYHJ+t6EbSLX8xwBJfeB2qyR9jgHfjG79C
8pPMzxC0pRCIwIeXIuiK+dIwNmd4V5q+MqC1fKrqjUSa/nQcg84Z0g6K1QbzaUZsKdhM+PnHdulP
bLb2HiFC8/NMyp6BKW0Dc8SIX4pEx9WDbhDMK5F7jLVA2NEnI1ftvbiHSv/IO1DVVUepgmPItt8D
3DhIajmjbW2VRiyEt8Jbu8n9vtLR+gjK+sPGRdDpicndVo95QWaJCl7/8fmNLdlviXviscwPV0Kz
q+lGlt0byG1WL+OyA9DmB1+21qY/pymDuntEHood+Gm69vjiSuhaO/EnyX+k6j9cDNPKCkKCmD7N
7AWcpNR6l8B65xBCg9pauRuuWxEGzGBmq7rEHT0QDPW/bdGscwtDyUu5jmkqrWOrGMfyF/Hq8rh8
R00bQy9THI8TmrZiUdpRfkNRwhG8bm56hu9DnJRxZpfgdi9WolVb2fQZs3QlAjFC1XG+hbekJ6pL
CBRR2vZJ5Bpz0k+u7cpvEM633d06eYnpZUHiXgSogJb+6+mSkDwhPhs+xwoFGYF0Uh7kC7raNugo
aOGeRe/G4IAiGN8hc1zBFSW5ng3x2z//+YeQdxrPI+AnRoNTihdVt7fdVKiGFrQvwJOFWiSWAA0I
ah3gOzHLjRKWADlmaMcvQjjtO8agMj2XkYCshBHDjvEO9ptPR0Vg+N7KnY74CE342qtaaNSc7fDG
+1ZK5+R+mNqHhCC33G4tWVn0khxmbRtpFBJY+yE47augie0CcQUQQ8XMb0bpv0zksFQ3XDpyv1IJ
0YYDpv7V+0LtCFbDFHppsVEUbHolSq+ZfDLBMmhZ4BHfUgzp2tfyDF+MpOjs6dVqxvonfd/268EF
O0zzckltE788ITHGikjYuDSSH1pjgjTtibZtQo61zWQ0rqVOh/M5o8P70A+imiXvQ8tgPS6V/DXv
gWj31zsn5LJvsQl9FmkDVwUVJznDQzwsjIHdb/MWwBnxl4K4ky1I83RcMk79nXn/lb7j+CzVPb1A
1auqXB4Bk5RoxHpVrJU9nbXpMgICUxWk/4mdA5Msv7pTanzxjFheqzqUZbG8xO42WIYG1m6BKIt/
dMbO+XEcZpMqGFVPfvy6BB0NAnR6SR1pSGWC0A5VkvPMMOgatKR76LgC6mSB9NDC82tA3vm3Yabf
4lqrQrd6VUXuui1BeL5dzHlXoFQ4faFzUENeEaw/wwnw3eOb7WBRcJ2XnJXYCSGoZTFq+moWHchw
XWHcpp75SckT7qO6dq8RK6UUoEqOMGY6ZETsTx5tS4bQ1GSzk5jVF4RXS51tonLbHgvohbgCts4M
WteU6MmBsKS9GWn+w4tFZaTBmTCZPhIuonW78CSDRrn6k9y6hUDe2ig5Q8kvIZme4je/dAS6U5uO
U/zaelU7MTc+a88GIjomA3wRIljIctyRvkM1s5B+ySXroi6UvMso7Tfg5Gv6yvbtx8cqLUc96ANn
lS3M7IMLpJE/13xWSN3JKfhgTcis0hgSExDlMkoKyCH0IPn/r2wX6K3ElUF69aZ9QSGRsFUtZdh/
tb1jtQx4yMYdLM6L1uQbCcQqt7FlvIwNiHqUFLlvd1zE9RUVlbgP9lBJ33IejwBcJnp0XkmIQZAD
C9kWPtTTV95w4GyFWDVKnRK2U+Awyu1NJIMfvFvPKFEaxGs7V6PdkUteE4QKzCxF/fwlfLin4iCi
v7mCGQA4eC9VbWhtNTJqvDe6yxUo/edDPX6qO05+eDkl6AjmKzUQQ5q9iM4xUpr3KpGK063uIJVI
Qkty8+rYeHJloOwIZe0hspxxRQWADJ/ufNM8er3bgIRa0Vc3UCwNQpmMXfY0cdx0nDKxzZGE+8rf
EgyRTNCfZVSJrgqsydq19tP7wh5BsliL/c7mRKzscVbdothF9VGpLpm//rODhhVmWY+VSqU/5xEs
/mH9eXuOoctOzHPAEZQdJZjKwt4XWj7R6RqhQBYGotti28UicfdrQVz5PZWY2QJD0GiXX1VvOhzq
j2sJeLrixSUf5Djgwq3HZQjpiYg4Zk3mJwteUfJ0aeqvzRBHs7Ly/AcqqkdwvODoHfPdhy3ULKca
2wa4LIcnY43JBnBZcJcIaxaJZDwHWrKYocdXyNITs7OJqZ9RlBzJICPrWNJtwAl6jr31KDOQTTqb
ytDX/ETGWQcw832erAIjtndumZmOaMVVCM036scFNwBdvShNb909AmsSgZWxjou0sDf1hZrPeiaP
dXYJ5cil3AAjRBNy96pSucaJH1ibIOCvA3foJxz9kg39P5qsA12W4YWZMY2SFGacUnrRFbqaq2bT
8NuDUSgVOCqW5J0FQYApbaVADfLJHfVJ69vqOwtwV7oSU8/r5g8qVFd4WpMZRvEa+ov8Jo73zdna
c3C7gTzQ6p388IpqbrbEXLYd2+bbiM+0gEHdB8B2PffNGsc5aRVNK78Y/Q80kH0dqaHLKyb8MLxI
OoY/dZCqSpebCyQpPMt5s0MYaisuaQD4c/iiYF59uVj0sNDTmbxBuuvRZR59APJMAd4mP71wl8+T
JI8Meh/29OAlJySMeVnvKs+Jqxjg3pBoGFlch3Sl0ZJt7be4cpaxSwovyItnSi+5QhfhIX8d47mn
UgKan2Ijwj0+NKIHPUrlKcU1msfgBcnOYd/a4hhb5yj/ijrnXGvFppU6XtdpI6RF9mjuA1uRtIgI
BBHMx7O67b3LR+Cy6pER3mkN4GTURGPH05Jk+TGLAhMRrBSBlt+ZJqnK+NB5FHV7pYSkaz3v/7dd
uNwzmOnq1aAbOT0TY0N98y937GZ+ExnrlDc01AUs5KrT0ERsQDhEavVUDM/EtgYr7iKSDsKFKfMZ
ih1lzD33EkvGN47uqT1CBB3XVEcx8wvdWnIe8m1AsCH/y/A3dkRG9tQLXYFH3aMxHKPGQucO1FZB
W55RFVFG/e6beFAeWN/aEt7+X5gy550s4baRkouap4sbeBaJDCQwDz8eJKgzjQEANMmaOi3caS6g
IuJljPxPGQJAxILCqhU4h64iUxuKWEAsozHvveO1/1HLGKU5LQ/SZzblBRKBBgLiVlDzqlCmltBX
hlioi6PbJTiIYWMbr4B6S6+UDWiOgNaFnscH5oD+vHYfFc2N63jMXAnc/I8im18AkWujJhUc0r6U
6MiBXSCIL3zl1u6i48DZKPAAToRTTEWyuUCzYBd9nGwE65CTRv1zitti11UW97D8bL5rYL/3ZMTv
PvVH1UIIAhPu3dORGDhUbzfll2vNYoS8GuQP35vsF/VbRCovwwsTTQo94l5M2Vsa2g414CE/TnPY
/fquX0PheRx+k+5xmrpJtg2JaSmSVb8nipL4Q+ebsVKwVv/12r3inRNUHIxhYDtTQL/VFkeGOvnO
ZOjlPOAfMA8BsaaQaTRK5EJHgSXLG3dGu31wyJtNrSZaO9NLgRQt45pqSCiuA3YLJcfI0nk8awZ1
8h2llUnYBwzmjzs0PE21fcSTVf28WhUiXj3lHpWfQixRqPkISRbMyYS6u7S1u+DFBj589aef2GWK
8Y7F2ycl17k6tI2nBrorjm81kjopdT3PGBT+IIuBGbwud1NZ8tU1e3mBoo+bzNG1OEnpqx7zh1NT
KtJBNc3JPxXnGbbHCIGxPDiAougXQy0mf1kp/HnqBSscbTkAaGFTOwOFLEtodg97aGIv2vcFYhOC
x+pgCOMXsnL3g5uZ7lWGn9/51VoqlpAYb2PHZK5pIDyFsyNcC42qdaJ/dk2NUcQRY0/AhnIKIDYX
a18hZTYEavEDKZEzU6qqvjUdefd8VULrsXtYEo29Bl0RsdKs/I4rXOa/kneZ3NvCprsd8nlI3AW8
SnZ//TBPaZB9ctsZDNRXnWTqbXf7qT4Gp9C9c+8BgcOH6DgK94iV5olZlIbuCUiO8ECPCpnpaGtr
EptXQhnBWXdaBls7YU+ToO8jaWiKpfpzyNlOvuk6f8JXtuQHaqni8rHjTy/6Quvzzv4S91eT3Kch
1tud4fG3H01pPm+V2v1tz+oG0NPdjE6kzvfz+Riz5CpHzEHpOwPHRaxUvoZIk9vmkX2wad9Af4Dq
PubsGDp7mUClxBs6OopLuCJ5rmKel6+I6p6PF/ej7b3OhMtvorhcQYhr4MAIx/32Ds+7xcUyOhPd
mKZEVEhH5UylYjWNsw/Tp8OGKKDVkFn5ZggB+4vYgB8fLMcSJIUKFZ7vwsHEZifYnVtErdbiTSc6
Wsvo9P6jAlJac0UwlCVqXC4Vt1MovPNxxbDXyjYrmOvsI/mpXWIIMdciy4MkSXdPFvQQF8CbVzFq
mcfBecTp4u9X/k/BcRaYnX+iPtAVB9NTVen3G+oTTEx+BSMf1zRebaydRVa9mf1WSxzDbkmCtKM9
Qp8+7iiR88HvQVsaPkbb7f65Ks2b1laPPPg7YFydyyYtDxtJlSy4hChEos0UwgQ3otXElS4zPulJ
YZaKTnKw5lt72lGcW4DAGVjtm+xGvK2zkiH+K8HqJSmQRdaTR48q7ary07bntyfPNDdYQpX+fiLt
sBxOIjk69aMmXZjNCrLMfNerx/P6qxjAv8Oe/NXfamA9oJt2UzFZEqAJfDyRN62OG+aJdCUI3ZFF
M2dVFq9a8NPolWjXguHAJP8oTp4BOA50F0R8uP/nrblGpCtk2GNXSA22H9jg+ylJu+pO91yCRcB1
OzWX8fhHJeuaJBbQ64/nehxHQJ4Iki1AmjJx1XzjAZLGJkPu7ZPf7YG+H+jxQbOYy/eMFKcJFeL/
X2VPxp2TuDknromGfJFaFhI367xLEKc+w0Y3WSDUoCPSR69WhTs5DIqRuB/rzGfCM1fReK4Y8lft
cTSI1yagePRN+LeZ3lXMap7DqwKkeyMKc4/CEOup/wDwAiuO0au7ijYFFST74thFsp01FOBaCQ0X
pZwSeaw4ACoIa7KDq08RmwlrfXWdeSuYdviPpIgKZdkQ7QcG14OgtCDqmV9gyWteonTyABGMEVys
bcH3sNUv+u5F5lA+vxinB1+Mi3FW+l/117D/exC0MlhRdBhV7GCkiT7Aa8SeR67iAJFD4WLOcFWB
BOlsdAxo0So8agyxZs+2ngC3x8/X+5IGHK7RDny9dlePSzPljhuVxAxne7Bf/PK3F3FRSBt4+m13
jBxqhtoTWomf0JA9ArM4NU29dky56oBa9f8kMbMSDT99bsuovMyd0UI0UdZGHNbhO81hbZ37uvdy
zP5VFf9YyjlZI3OpE9T78COGBB5+9AbLvGz64DCpVDek76p7fKA37MqSNSuV0cgVIcbcxkdY0oxw
zb57kVRl9N4aiiCSI5FHG9Btet8vaIZ5/c4JqVQF6Co4ycepBwNGMJDDkPryL0UkV3UR4TQmYquU
pENqMCZrc9hwph6SxXHa46DguDGWDF5ZJHIdtC/2/3Ur2+Vu1nyPtftZnT9lxaYC/XoLJgg2ZYyr
k1Z16OfdLeXnWhDupMdf8DY08e8IIsQZEeUDpC77kH/xICGdMmdPPK/SkJlbMuQrQUdZRSFmj0zU
P0FE/V7EuVanb53co5+mwMUFD2ITblG6Rw2lwvJajDqTwAkveQxEnAMgpEb+G8zQUePRDnn2aqZO
QkrmWSsPc/8ViuXO0Dg/DnKjNPrNrKC4p4Dz5UU7fiKQfpjjyuHved1MOZGS7t6WNiHLhHjsCo2V
qVjknzuuoK0h3Ci940k3lFla4axIervWFv1HAqz2skf9ZU1raosiqSSxnZmMjI1+LrUeuXZqfUEi
pNxrZaxIr7cGUG0dJ4kICDCGswJJFkgKl7rMKSOYIbvXl/QQc7OUo882AwK/nCS2xwHz6kMKr/3X
9Vu4oKB0qoA3rgdwLKcWWe+ZbP52BFN5PhMoMDvLrRK9A6ZTnC9B/OD+nkVojYmSZi4ENeF5q7W0
E3OX1WMnjHWw3+BW6RBBTC1ZqzLnDV9ZqvC7VoX3MH5oiD55JMOLinaQAt7L/YWNDII8W61A1Rfs
+4t9wHigZIVFlHUsYN9i+AUiwPoV3IBZEGUlkk7FLHE2p/t5VSfIveONtrOn/IX8Je+O2z1FvZZb
YV37+h2sf4ghj6Q33e5chwkLQh8XSimauWwrDaK5vkylTnVr20ZtzzTDarBM71OhCS4iwIYuDtEY
c74aFR7SIXJtCOzuaBQJYSE8jaUI1PqfCrRJh8LZI7IQCd4sIQFwBRaUguPKR6ELtTSszPM26Gae
yktMHJkiPwQCRhN8NnF66vg+dwtZD4Zl1/Tug1qupVxfqBNPGEYya8ySvIscsfpq+jUQmWJjy7NW
EMCaUb+slUCXOHXJyC0gS0yZVwpEbQi9n6BpK5uOdEbDeLnKwDF04sHPSHq6PgoIh6FGWHc9imVE
g33KTZ/HaLV7wQ6Zse5qhGMVJrKT1rGMuu/oekVOkalEgmrXtOZxFRuuBCpNmVkJBTIe2t1pO2gG
0zvv/vBJ4ZtWIh/aJxe+Nj5S/g/uLadnNftkFKCLrMUZ4ppQGc9zEd58itS9QNgoo0lrK6RzsIFa
u08q946XIG7ldAaz6QOBgVGK+enGR3ben3bzO7L4SA4mwMnZA1cc14NXUvP6q49V6WhtDBYz/RLZ
aKd7nlQjbD95g8EMWt0fxF656zPpq89gntDhLCQRqdyZhYDPhPUurJ3a36sBLdP6/fHb0MHMPTZc
CM7Vc85k9EmEmhn0I8bX8CAELloJ0uy1c6NMkygATM+ki5uEzHBGOfmQqgVCLjgqAS9IZVldOzme
o3lCLHL7WYsEfiumqyIDCnOudOFDNpbJh7flOHPZbKhqRpkceG2Gq4zsPTWke19hw+h/MhYjztQE
6C7MpkE7W36eQFPlliqWUwDQE3Qh0DeefTMwAseqjGgtA+8dxEvXN9FRDBjkMN3R80z+pv2OkNFR
jsDhFErMYNsM93aC5tn8AEzM8HWb+CGl+enwWBjmKD7qlG6h1/I2YsZbF5n2um+JUB1zXQ0wV5+R
zkiglqR4PQ1e1EJ7RxlZw2SibcVJJXZ30CXNpRRAPALnmCAQw5GpHpgLVABp4YmOycRUDF53LsfR
SSvzSqfaDFMfXQ87Iv6jNfrPXJtOYeNnM+CXN/u+sASSQq9aRlkDqcVlLpwE7gq+CPIJIDSYfek8
ulqvKNIp9V1n9u5kjQeXVzNEJfa14JfbwuQPSmCBBTPqMRbJOpCFnp11WSeYRht2vWz1r7PZ3NZD
oMqb4zu48cASPnIC5ZOlNP7HBjg+xeB4++8pPKA1Gj07mXOXBBWOIh0goXPgsY64QQ1gYNA/4LEw
S4zgMbKe1Im/wsC6ssu2TS3MtMgYXLHx5oCrBfq+g1FXNz3Fwd0/7HOApsEuLE4mbMNgv+zvjmCN
EbICOZ/9tmVcGoDkhuIAKSx8QjDTbP89/OBeYgTII3Y5pozNo6tPWDkS4cr1EFd3D+j1SlCSUxt9
pIegbYGVXCVLQRLhPUva4ZeVTOTNkXUkMdrm5PnO3W0e83oV7giHXIoF+mYuXqRj+PTmJn7IDfl2
03OZF3jVIdy27SrqwDipv3IuGuuWDS1uPFFEzBVozc2TAJuND0+CEd+ETNkibLee+dsh/fKx7pMx
texmJZTTtJh3KgkRoYmND/0L8Ohwac61bcs4MbHKBnRRmZGCX4lfacbiQQdj6rjTUPLzo306rusm
RRoMXmmhWXJToBOmsaEC66C5jdxFcU5SfKZS1BiZuUYlFSrqQrP2HOvOKDA7bn3QAVoJ5+77kvLN
4qQ0OiACil0gBNuw3+b7C09KPhodlX7CGjza5hmEEohKMPDsR8soH7VA9KaqLVQaaG5DAMwVnARH
VJu5McEey+pgjBsajRBUd4bVpgMFtqB4jVQeTsiYeek/gXYkhwAVOfSIyGJl6ZXtADy9wPUUtpI9
xS9z5gSxWrKS39M+K4qwpK2kKczj5BSGQfgNLVpidShJwL+5kDMe0NHeUFWSriTvFYfHcQPk7NvD
Dh0iG97XlUf2bjgBi5RTHao3dkTkJu6lyJhy3+70QJ80BcaF9GWdNLOOifsgBlZG/auIWqXe6u6S
MyDKviTSuKON/MNdhM1hODmW0c8GVSnH6EFGMM6TPsLwsc90jZg3ro/gZ0WU2admOGgJW3LATyWF
DE0T1y+SoirevhurQXTHk76Xu7ip590HqrKvR4IAhcvRJuahCT/HDUDYX15hgknjaBOx0pS6k2T+
KbZp054wvdYep9iQPjvAAPjZhVipRP/ZFNVRnkBHPbbQMD3oMoFEpofG6PLnC+8yDX6254zqbGCx
AHeQSV+Jr6TDeciBc/0qoU1a3ll7/uNX0smad4Zd/xD5J2zycztFbDDFBNGJjKXBuW2WDwklNJ9z
XbCN4CoYpVDA9SFNI51wbdSU6e66eSeJqiTIRMaUqktUuui43Y7pjjMT38AIbUIhx11LZuwRYNcc
PTjsOjCbEbrjhQjuGiHWzi9v7hY6xEBw+Fhwbu4I7cw4Z3A3vbV4s9VA8jz1tr0ewLhzcgA3XWgN
It8KmukUqsdpWHsv3/fZQmiAF8KKbRFh0kC3pI8/Kc8uxY4MI3beIKB5SXfJC8Bt4F+EoYT55Xea
d3j7v+wVBM7sM+JLQBjxf1pL1RnZSu+ZHcWvGZJ4eOsAYAY/aLm16lhkizx8nV3SU67qhG6Q0RoA
vALyBueoibrfB4yD2BJM38WdY7iCk2X1QcUTidtxXbhGFu3Qcypbjc2EzLAvw9nMbkd9cx2jhQmr
CaEPHqVPd3utPa1GZcteCq1K0dsLqZzPm5+Q/EcWTPYcERxUEXZxk6mO4RSmopXkEpv+7ivFICD0
DhjeB0yKRNdgB3XJfimbKgWUI7xepIp11sPcfsg2jkq4kBmxBH/Yt10w12EKivu9mKF54brr9S0Y
B9h0Eb+2xRF4OUQRmNlZj2rsR3VwZCHrpELlGSGscT/OtcbLHZSaNw6szM6RmEyeS3ROAWYGmBjo
FVy+/KEs31U5FMQstY+GGHbCeFNNm0D2nAy1iScYRkjNNGs0cyQWUnUIgVCkrGqapNOrt8UeL3jD
XUR5H6qHZA0+xfWJog3OdGhnSLmJpI1B35dtkb6kbI95w9mnZFUraeID1qpWV4/qQTuOgu8Q0BJR
ffvzOfvCnyxom94x64c1p/v8/bdl15HkvW5HqtVZ5JYEZBu80OaNiXzim8Up7O4ADt0s2Wk/jcWV
N4B0H2WrL80Tp49DB73LA4TP5/aa/exsj5ENWovd1Ya+mCwg5AmxZ4OpBRcdRDwaBavzIlt1wIPt
GmWwXWEpLF2ayq9tc4J4KCLjZgWrps2fWzY1PDHWCzLPg04Wy7+MMUvPPT6lUDD7jd7hxQrDQzHb
/lICz1ZU5sk9w4XxYISkdUYjRmDAp7a8kTO/FZ8LXHf55FDLV/PpBnDOnHltnNP50Q8KxbW+Wv99
pF2l6asd2aprFwL/s7y4Xn52eQNxVFT3xuOspnCWsJAode7771uCM2w9m8Ug0u+BvxVUlUbqUdFJ
2GEKS5n0BOQa6gLi9qiU9VNrLajrmbXDDEtWWW2k4pq/TQb0kKHX/KL2JgajUVKWb8xx9Vxjn06/
FfdrZLRZO8Rv9frdZmDMzUMeVuJP8Dt9F40igEETXSiXBQ6ikC3SprgxhjFd2aIi0iHOuMPTIqGr
hVVOME077bSRzlk4tEEqW3ITl9ZvTYAXs4NCXl6HHrO9sagGxgr8zV16D/vhwiMKRPgNukk1DAUn
90noRQX2aLTIRVxN8GvWfvXOZXa+5cqR2fcnNPE80qEZbyfK8eL4A6x9RFOLgX2MVWi2cavCByyk
AXahG8BUsy9AL3RzlBRmfcGMYUIxy93Tlcg+KgFfCBxJictP4FNLBdUA9mKEoUN0bVdEkFvWHO0f
puUiyvzH2cGZ8rZeGMXcixTV6q3q5jxYf/rCSERUXy7DE+v5o8JmC6oxFEz7gUCO5PIqDte1BXjN
RWVkGlq6PYfd7RYU53iFmIxLWvVlMGugxZ3OzNKRNFDOC/gLQxlrS5h3rMsFDfuq1N/IOCcWGNOw
EqDHuanamBoxYq1zQCB+pGZ7EABiLe2D5P0jgGLrtT06R9sREPxnjvh6A4LYJLE3Nn5lwtZwGxz3
lnCmhhIoIAevaVVB0kOl/aLSAa03KRnJVnZ9OAewzvyYKsK4hipjaVh8m/Qn0HSvuN3pdcTIYKeI
jGOfU5dppyYEHlDfICJrQYcrg+3mT7whB5BmcQOW4wKdEWJcmI7L5b6meN1kYIGscSs7ggifxOlA
u/aqhAexAqtsjuuLMvQ8X1mgaCTxirq4+ZCcQBpVd8fE6NWTsYheNrlkXqHvFUTtb1dGmDM7r+Ye
J4+HB5Fu+xZONt4KbTm54N9YsuIoNZt0+GbPRI3RLY4f65W44Y3YdjZkEx4w//sMEFu6SbASuGu2
JOaZz7Rb3SaZyfQIFlwFuqeP150K9sSLghwNqnx8S8giQTQOcfCvlV1vwiddabvYbMjl8tXyyx8W
Vnl1nKQts/XETggIxDcU61LYJhxUlALkBXwVfU5DlmehKY1kxJvzgapoYSCTK3PDJ39YgvItzVMm
1MxHls7ra/OsRzs/Kx6z1IQDmsLFLcES4GCDCTGAw/SHqlepOQZlFsuSwyTj6T7JOavh945HMRAz
56TiLt5Rhj+bY2MyPyJw+8j6Zr0OANjJ6rIR1wE7GKeMOlayKI5CO1rv+5KNpikWlcxzgvBFWDZH
C9Wmhn7QKGA5RKKPj7r/kJ726Q6dKQT8HPkkgZQaDAJoihk32fs8rQSdlCZxhOsgabjWb7mTqR0p
wFjOVN849NdIQGq/ODMuWdIiYlWOxojBUVsapMLpSz8Po9/ZFddrJnNQ1EZtTZKq1Rt8amJfP3Al
U/Rsjyi65pCc3kH/Sn+cTsbaMptW1ORmaZ+T/7QxgBzOd/y7H0olpy1DClep5sdYj8aEBZqTMWCe
8poLmQhe5DLTgE8YYfiDeOaj1Ly1FG9cy0/zwyXjIM31ORLVxWpOM64HnK8FzysUANVynynVNsll
cPwJB89nt+DxN4eXp/hTzxpVQDX0orbZzgqYHtguvinCaEXAfNv46pi211+M8rYuKfotuGM04tHJ
ufsrtaig9+MYFenZn7v3av3AmTyOBVW6VmamY91sxKaiALAZakjmZ1eQxd+hyXvsK/kV+uFvT6NA
URZDpwKjh+X7yFqjG3Nw8GRY7L0/S32m67BvVIa94xdKysl+PaTWOlncY+age/W2i/kOu/MxBQVO
uW/KWQWYKoEqbdcSt3n9KCEKug9O/XoUv8jxu/voMeBP8GJ8M6t6Ne/Jk9by3qNpRZCLRp1fHHiW
YQx8R95G7SxdWMzcIGtD64tfk2ifOXIedyRht2qQqHnewAX1FURVILQzXluAi7Xk3NcNce6ZgRf+
7QSOB3JX6gEnEAdy/L/P1zjDB55mIyMYxbow0sNSYGDfUiL6QG9lstDvvWS6xkNMgZV/Mb0owj2C
9Aws6YP+Q4x/2y5FajMC11E3iaRrnVCR5qsOPhanCSzd9btste/dIXgh55vE2pwqbONeRPu/kil1
tOAqqYqArCLritNfbvtzob8EhHJOSEh0U80rL/u8fJEM3ZW8jOUzTY7/LAcYV7chaIRWDA94HM9r
um4J58x53UIceWh7ejg2SDP84VaplnjKn8lrs99gHD4meRsvckfreU4ZD0mkKVcMu58CNqmk7Z73
2q8KilPH4OY4bT8RM85gu3Xl1FjCpIQWFIQmRHv2Dj/OX9QQoP3QxIiar6lbjl/LP6a4l+FN5Ycv
y9N1FHVER0ctSwH/Eqgd+DGvqKX7SXxy9+8q+06GyZ+uipiWR+PAxSJWjNPhnRq4M+S+XTBUqQ6W
sRpjXuO1PnegciDs4bTbq4NcNSNP2UvKv3uqTG8W8q+QfxNU/Amv30GyD4aYsyA/Lw59N1Fw5Zqv
1/0nZ40rZbfgvjVUqinigqSv1+DEeXGjlh0o2i+Wa2pE6HuaXPd1qnvEPPDdoVImvUC7UO+g/Gkr
nsJUNh46rnxFQt/TXBsjCRMiQYxl/j8SCvFPmRaxrkI76lK6BV7LakfbuA4z32N5g+7W8/h1oUCl
eaKLqW4tbHEkzq1gRGYVEqrwK5X6k+lDdsscSHKl8PphvLHcaRuJ5xvan4NfV+YzOEUbTuvpgHls
f1wQEknhTt1YExJ2uhPk1jfGYiNnHn8AzDIjYbij4ZNOURqjWIndTHTEw6QjpUk/a+97EtZ+ULR3
IO5UHIi6eSGB6CjCWVWaCDiRdUgQ9Inx0i4cbCDLK9Li9ym2VkK1WqWbh1NrB3/onxkoVJ0yfxQv
D2b97E1L47oJso/IlNvVYN4A7a2+I2C/Ef0h2ff/eR6zsEp83yfTsmIsxUENnDDyV3cQj8nrspbB
IyMD1Iys04WOIreqFGmoN/rWv72qQ06nBDkkAf0JG9yAEMigC7S2b+0TAXiz6goDDuEkNXyztB5K
oSMS5fduwUO435N1u1FNvWtwaZ3yRAmXsUq91IJuQMZYgFoL+Gnd4ZZep+IaC+kaGCbmU73j/dzi
oK177PtnBrdlSH35HxDgtRqW8hAA6/hIMdK7H8Rz7FD2Ha6xuLqOQpL8CY0tasJixAnZQNy9dbjC
yEooCFxIv5FpMkBgkmvsUjqnEx0DKfwdL6G14jmCsckrDceicyWRGUtA8A5jVsQhD4NyBF0r+0Gm
CKVsR4MiYN24pJbHPxZHwV2zmli15N+JtG8USb80tguCAJATGhfW9sj2b3614PcAg+yLk18M9Xi0
UWYRYsebAnSGb2n1dvMDaFQHkJxXcYZWIM1ULmyGTr5Ee3k63rlnRNnbh9Xz9qgBZLiIfoqiGmBX
xpczwiZU/RGd4DuFwJUtEOidn8jcXyT6bUBx9h1N5rnqn996Dus8uHzsTnTtXy/CMKOXD2SERd2v
u53IwR2IAePGRC6PVynB1vxji/2l+034JJ7r68zaa5rz35BzkGqXpNxWGiu96U3GsgnI0WJK052P
ADBMLN0e2ilm30lc2Q1UEIxsDrBktvmaaVq3DZF7nmLR6z/B2ZwPdfwx6pgF77esPlFUajFdMKZW
CVZKHNDLhLWiGq1Lkddz7EBSZEkOsh2iZUOMJ90e2gKrWr1t4lQVa5avZCq3MfYMIc2wcR3lRf/l
bXn17TO7V3mQzAbW4iRZwu8T4UBGxSiJpBbhPo7DB72Mkis09A5+LaTPiaNvbFZ91lE05MdYf3ol
3r6lA9vh442d7YVQmFa69U1opHs9T3PECfV9f6gvup+ymnDVWcEeZ70rQ/6SkI0E5D8PuR4aiyD0
4WCWKhBcELKPyVlnKQQxM63N+YSK9ljTwbnTiQswa73PqkMz64DDi7q5xV8F7t52L6gMwaLTpcij
qznSK2q4nnCVYdyRt6lTlgOKuBvVCNdktDjCiteeWF0p7lpEReZAFaVbriEGusJNSTAFNuS+DGll
j6lIrc7QZiTRkQqq0/R4mO76OYH9G9BOnRxJxYaHiG2mTD261Jybt6Fnes4FKbuES6gbZGz8HXnJ
fDeGF4rFTnz2mO5EIlIyznYkpfrKIQscQk6FdGIgq0RVmzsswZxOhsKCkyNUELFIlqre3INyR2v0
Sj+6Cu9iqOJPb1wOdv+bB6JE3Naa5JUKZB9wIXVNEJUErxObGuU98zevKDyzLfHf/YFIOZtnnyIG
2/TpFBD2X7HqrmdzdoTGBVmv112JeLlHVZlTFowDSl8YxVpYAl/B1h8zw5SXYBWMTvwQw6aFv47Y
UNN7FL49rt8yuGzCjRr0VTx1hXuaEo8Cwmd/j4bNsqKwtmO4SMJHXX1OfItSDqy/uqZH3VMxfLno
42ePOkV8UDPdzZzv77fnvr+OHS6bI+6Pwsk83wGR20HZb/T+69839biNXafOgoFFkZ36Wp5zY/Fi
x7AWrd7e7c/cfD28g3SmqNvt6ENROMrZ6KQVpucL01UzB/iuI6kp1pJ/3fTjLTwMjf5qRVYf/qua
m5t5UTttdXcVbort69qVwTwk0PEa3irBnWgzxmGSsWH0RSJJqFH0KBZ3j4ewDPDHcF7vcg0KXdSg
qBYyDoLwzcs/M81ub6w5rezKQ6d85C+FbDqaIXy8QcxyjhgLoJ6xhVP0s9gpiDinivPYAQlO+O6D
JJuty8DqJS9tIhvDhL0vix4mz7baVCZHJf/vpTXRrntZKkmsmN4nswRIe7qziF4udrpZh6tfWlAq
tWsQsQHsm2xTNOBjKhXA0cNN7IdPILOu3Vke2HAdf10jnJrRRdSNjZf7nlYWzeAIEC/4Lkg3MUr2
f7mdo1oeasKcqPU5gBPnaQsc2onRcNLF5H6dJsOIGdn48px4lIQcuFir2HcaW9AS6PeHXLDTu5MG
qBilnyY/7XHW70KFZnT2QnEjSKltdbE8qGo4YGA5aJ2DuEAbas9s6UFpzsejnh0/FiSbyl5i+KZc
wu/az7PARxbW4+XXGIt6zbyRYP3B25EfGhC0VRU8IfWwfnjeZQeqSKbL3oNKwY6JXze5lM7OhwhG
90cA4fbJWwCZxbf4Bx1H+c8GKF1LFNvTM3gHhenriJyBp/Iw5B5fPqw1XGYps97Jce56Ex5n5X2o
ZmpUfCwSYErXv5D3kbNTGmPezMTgs3cnN+5i6LL0zORsLDsdwhbVa7ngufUuspnRzkQ1M89ImdJp
gsaVV6SSAjryp6qsq5xzU31dAXd1BujGibC8y0AjoOeWEJf2oD5uSk3cFA8Z3/JeM3TtnaWEkiGj
WgQajR72id3/RnFkFFcUkp/2ESMMl0vgnDGV2JHE4FL1UpBxeDbyKyjtB4fWVOO01EAIG0B6i3tb
x0zwiiz8IrF4yDNq1hrqeoV2S/JjXroFBPbnB2vhurb+csql6WxzBTInhFoQfnWIQYWzhSrTq0Vu
3UVZ62Z50GVZ9xiW4MmVNtUn6SmjA6r2IXwSpAcqH23+MabMnFDZOeILH1v9xK5BksTR7zbMj3of
H9dzMRItZSOH/2oZWHP3fd4I5PQOVrwx+W0vY7mDN4leX+XggOeyeDkWpCSyexrqSrV/9dpfYbaH
BcwOHSM4B4uPxgqQJqi6kVwo/czibcZILH5G+0Kwrif4dghug9O+zvanhnsdLkTREQFt/4ng/9eZ
MSdJvKIxNkvctWTqz6VOQPXH2gcUpJ4quH1dV+ZzPXYj4o7A220WXbl9jG68cnwQjiwaZKFP2VZ6
Cu/tHFsDs2yMbffqoZwVclGGWKYMcvdHTV0UIxGuhlMqHTJeWX3JsjzgehCof2qrSLFmEBPNHG4E
Unv2iiYEZzBl2VYukAGg3hjfAbT0ao4DeYqjqB+A07sZ5pKiuZGpbrPsGPykjB551WNrXiLHWdC6
oFRKxYyrhT7x5Rv+dwGb6DB6HHDYV6Ed2GJdXa/cxBcj2fTCcWDdSGM0sLfMmzsJxXjikECbdGZm
x5QoLqQiCNbIgV8Rd6J0CclHesI+ZUa2on4kR4bmgdmwL6HKD3CWJF0INuAb0LavfoMdxWRe6ouZ
pFPoKMxvgfNr74MX89qJ2eL9LFWOjYpLFmFWzrgpYpfHW7QRpI06kCoJWo+Zm/kjrPA9nzG+4dXp
oqDiSgGX7+hRwcLum6h5fi+DvFJYBDwcqM9zt9q010M/oii9aBPJkLaaUpnMsMK9IoyRAJ6gPtyC
eLLPPfeZ6/XpKvkqBGxk0KAKEr5esRUgz4MNLehKM6TfRqk4+2injwfkco0JA4bSw6Aeu6fd/8cq
3qQwOwGUzX9QQ4FI0ci9+yWyFseKWC6yIGFRYoFSea39tiqbeXLdVKH9skh0QE2eFJYVPJYYmmJo
qOV2lX5mjdmQ8X5ny59BaacJo7v8q5NjZ0DvXu+YdL2Ynk31ppzK+y2my6IBjNDWnYVRQq6WY6yu
hi0FHzMf3c1O+puq4wysPOkUq9GEAWdR4BE0Ytavhoh0u1OShbFc8PcV8pTb5CQMMQEBQa6LYiCo
WPfCAVuMsK7yhQjmuJ9SRmlpfAtz+XERD12Cr3yDpi0ht9CMofqIhFcV5XiaIMVSbD+OE2c/+wFg
wH7/LdlHuopevj16sIieOQKOgNL0Bh88kir6t1sp3yl8F012Lfg5aUG8Av/KydjlPE3R+HfGbUY4
ssZJcxHlJWumI16NQ724h6P5cOs3UTH4/bnbPNGsUk3El8g8vOyt2E75IewoNSCP7QobT2AgsWRL
n4DdgIQ0jLGqoUMl+vabVipM34qHEp7n2Y1UJOrubKFAjpoQM26POxyfhXjuwX8LMDJ24hrRx3we
8KgaR25iMu5Tgfc4bb7DUqg4TYZK4cyj9Dv/kng7nzsnY8Mf2kHBr7Dpbqe9P9AaYAwZKr5yCyNY
a9WmH4ZOOvXX3xcHWK7YkAFatTrEkCABaYsXR55jih+MSsIJA90R6z10NL+bBTbh5KeTjm2PHfwF
K9GY/6a+9CPjhYGtZk87p6IK6vmGJ7nu3ZnAo8+fO6IMr0EC/DqMzXCvOWKwwS3ea/JDjK6vcCyw
NE3BZDUTYv0a8AE476g/oAnkDor5O08/k7LtpcxJgsv0AEfWJRu05uLL/uYk3Q7cUZscXXezDexA
njxziz78ntIyPJIMViWNgF8duOE0lPuy+CN9/Oshc3opS9rw68z7Rtrrv1S84JvADNEFyV1Zuw9j
GELWSf7qRfoX9a3CQAuYHenRsCPfqIvVY29C0kIXdT5zBgGCY96xrCMXmH1ipbAW6G4suwv0/74D
9+8C+fIYArXrDHAKpcdmlTueLL9Js+XdnS2aAbUptQO9PBTuo0ARz5feBPcsuFDXUAZYCVTXXo/v
Y+y+xaK9URxWTOGeyG9SCOoonmOyXk9Sk6MJ9n+WBZp+iGik6zl8oL9kBEE4y24k8U8vVitBHo5K
/popjEh7HZ2t/TRpTamfauJWqPt3Q2CHSLN+GBmDGd74umTeNOrgEIRppI0g7XFF/1ugqz7XlCVZ
nZeikln6iFRvzMUL9Yy2J2M5USKL2mgjWB77yGIfFrS+qZPPiX7AbRXBmU0p2M/iggWy9/28NQz9
O+fARIMbs6m3uvAP0RPRlkG1djH2qFHPx215X80RmAr0z0kJ25hHXJPBQe4R7OWk359BWTBTi9lW
MI7BqC1snppw1A+rJQGYpr3BCOx+6S5f2/HGLFB0cpZKyq8L9lfd0R65MLUm44cvdZKjBJzr5aap
S6pfwDnGWHGCiy1dTjEuhS5tZ2cRbxMvzAg0oPj+N2Y1C8c/DEfxUjYdWdFRhBPz6YQH0jd5jzPN
vohrjyeGEZbdeI69LBsO2e6hI/peqiBGSpoNcf+xRNm/4iBrD69bxSZ01OCtE4cUtUK11EBVXslH
eSnw+H/CmCr5Yu2YycKkELfl1FGvpRHEXylMx69TlJ1dobVBFqVj4zDtQ5KreUd4lttWnWSPm/4K
c/jywZfFP0yv5A40FOuMj092Epe07YiArdLhxPsKVwUEjsFGuf27BW05JHnNolCqs2fKfg4p04jR
cYg4YYdO44sE7yUuU7qnHdd+cJny9KAAvHqwCrArPpLzCCf+v+882An0DUGbM47PuqeGgS6sTTdf
32V1TsjwWdoXiT7Pph4J/HYHMMU4NxRAmyx2IhVLmg6uYGffiGfAC+qBh/RP41M6mVlwQ9AEPQxg
lU3cr4X8u82e2vBf3+T2qXfL/bDca28uo+hIF2+hrF67tkTqQbDq+TfBzqDSjhKSZi5m6Og7JA5U
jioYaQfAeZj03eOdDWp7cdSRFJ2L0DgVCg/XeWkBkKOhqKGrtICrKwH5YfJ+A3nQlpDQe2A20Mmk
+Uy8RFBRsXLaGz8PKTvuYzywhh/4YN0vmiiSPQlGYlNQFbmaRfhT5U4VZNDSA9mqmpR1MXfvvVia
w32jwuhCNVfVtxai390pDctadGRctlpSR0zQqbxJz0CQWw5RpVI4UPJfpHisosTqTB/fpNqDWX8P
ez/RmpCTo0wJIF6bP2pp6/00uGG/daZvWIhgREFgjaTY2AQyaxrL15PQxWz3c3KMoeXDm7ForEla
mA+w11yFEO7qHgK6+q6cGY2RpCVdRQM6Bw8solf1EdulH36FtL6WrWtSFrf7LeSftbExwGvvYVsO
gyK/jKOz8qe5IwsrbEqLYhVfm+lKKKzSXbjNuFTc2fo4w9gaS4d4t/OMkCRiROtDexoJ4bnkfICl
LaV2Wy0lpfaf1dlyJU6rjSY4XEtFg6z85HSbwiE8vsYf+ToALLhJe3RKnQbUQe/OupwVJiuvglUA
HMQZfhFryh+GvAQ7QLBIQ6ii0YXP/hhSBkhIYjS8AExBODwc7gQ00bsRLTwWiseKklfqzccz7sF2
ETIbwoFwfwwl5Noiy6cW6brJnJTwbMK/+I+c2pE+C6c5mhx4naouHij8iKv4Avvw4s1MVVtckrAd
hx4CRExH85ajGPVXaBGCdgDSkVqtk3t6FW41opgX8TGYT5Why2WdlFj0N2h6wpvk7xjRA4yiDLJW
jn3JH3RE+KKA7xbmmdJPw9AUtp5RIJJJ3p9FQY8Ue62BuBErlKqsribFdgj+aIn6MROgGwXruyGi
VY2cTdpfIMvuBDJbpJAhDWjAxnZlp1UaOL/eVN1R8k7zP5x5Ox6/eRKiPEpQoN/t/mN1iQhPBehC
CirhLg05uUI2xt7bBxuxiShb8tqaHVkkSWQHif6iqXdEVozeyuEN+0a410hWviHKPCD6tmzWonp4
IKXFQET3siDFC1TkyAkzfNl+h0nYTBhz3At8DS6Jv/CogHNj8dC1P3/egvVx5NUYth7X49Is01Fo
nVffyyb3iut3kSdBjk7DMrx3FCr284LCV/SBQGtSO73//agCspr5E8LZdvUUZmr68ztm0T7l9Jw3
HNpUQ/n6MIOlojn7md5k6U9dGfRDlMan6f+g3dbBaoaHB7vW15cYBZkIkrHaz5T8q54HJPJDB3wI
22vJp4pauEyI6acZaKYy4htmjCdzrktLHb9RFNTByVC8tGq0HroojFCGsxqm7/rZR9vWUXlTiA0O
eEZ6lnPENqleEK3+xUrBmEt/XmYA5Dd8VSfSOLSH/fHusqjLZZ2o0kgTlUY6hd+hhkS+e/Iy/8s0
8oUXv+Qacy5aUu1VIZrzyzDChkG9897uJ6+C4KSAiE9C99Mw+OFnj65O5jKf8waTZPenvLLy7y0q
hHFfgegqnhB0g2GUFha9JZu3VdPXUK97rvEU01FijIVwowTEJgzKje9c+E0R3GmBtRrIBZJ06wb2
FY2VVcVHHprmTHiSPNOYAwPrYtIOsiwqHVMfoGHPsbu41QjiefXQ18oxkIKoVPZMhF4S8oUdnujg
PyrP7tjlW+K2INXUBz4KziNz5+z8sS63Ibdu94JABP/tQwC/06dwwbls3MmlY6RF6gh1GIq6vFog
t3yGRvxCkrKTMSMwyjoD492x7UqnRglhiDos1i/d/B8P/9phWPN9k9npen6L82dT6zeQ5JjZdilL
+1SpwaoPCqUYR//yTrNRSet79ziQaZr3W/CtKVGfn7Bk0/CLTYDsW1K+RZN9jLq6fOnb0HY7N46y
/nD6Te790Ik8mD3XwG8+Vney9wwXdsIHow9xaeQIcRXsq3UjVD7kUovgasRCwTLySKotooI+yP0E
6abZHf42yPWlWYRjkb4p0/OSz7avdcZmGKAb7cmicP71Zq9ArkDJcWC+mffe0JimGL+IalznNZlx
EuqcByZeaVOv9HCvZRewYdK+VftMKaHBNTvAd9ONtl41cBakM8MCmGwUKtadYZoMfALbLOHs6I2A
grw6wuwrl/xIQdFDdY7M+IHgTpE6Ad/zcRYwRH90vUIvGhOaqn4I02DDt7NcIuHQDZSr/2tDHhm4
Kzjq5n8k3ziAlqBy3T963tsdASQLN2+f9U9ah6VBY6g2na0gk8W685mBX9VQCGYWbgDU/3DLj7C4
5AnDK9loocZ1M2c52CjNnzsOdeoxeHZjqT2+azRRwGa4hqeJ8LYrwCbIP5H5laVxMiUXcsNYACfu
kArAPeJFMt0EMRWe58dNSi7/wqT5gXHwV1nyLI2j9ZkeqiZ9suxzfs8r2MR5xthDsOLGe3M+h7VI
zDNMgK9xsKH3m7O1wcrX8dk+N3D+MEZ5M0HXSy9IhGtl15VBT0AUqprXWmCHDj9i7f/fUBDZRtFH
PIPyP/sizutIRG7IbcaaWcpyrBr3vN52hngm1iujcyIJ2B7U5+4iZlxfbO+RI2qSuaqt1bAVDkqY
TAFOVJY4RnVza//xtSAfvmkGOFXVX8BZGahrwnbLHrYGJgdtNnr3Y5rQS3qnCge6HUzZXmmGiQP/
fhkx52on9QhwvP43ZQ6DdEmq4kX1jYp8OuQuB2/CgSWlJo5olRzzOoVrf3NRguAUcYg58Dc3Uo3c
va2O2UlG5OmfGOgmkdqq+ywawnyD0dp6tg3O6uhz+ujQ79YNYHEkCO1gphN5RQwvSdYGacC20Wm1
ll/UKsQ8uAZUSSj7Z4UYIV4FX8nkP3AGX52Xg3GNlomslOn0NJsM5ONYwdIYn49CuAbiaPndfvgd
v/StFQ8HFMaDWqeoP2bTohvtlvQglBIB5gYXNMS5BXYLKys4aDiZLSljQaYpTwv0AkeKeaclR/RH
oAHGbXkp+w44Jka9MRx8T022VVPDus0Kdkl9dadeCNOXanhphCMWcR09mnQJzLZyIcFRok069nz4
ETJ5vk8gEaFnXXpmfKMQEm7SJjONagyBCUp2vL8IseYm2MksnILvbLc2IBJyODkbYgVT7G8hAgpT
27i8Oqfncja2aV4jpiHLlfdMWRGbHuLr4TgpcSTQCyHmkFrFSFaOMr3arj5uehCpgloEwGcapa2d
WKcGQqXoAd3PKA9UK8giaHjq9/USpt+0TJ3OTHDPCtAeKeqBfTlAhb+ybfIVOes/sLssZXvTjy+E
W7rtSEbtAI2dvxUY13cXp4yFSyRxXKnm8qk4fYc4z6566Zulpc2rf0z+o6N9XaZETqxCyC0+R+Oi
ocAA+9hE8pzMrBtSLNTpPpk2pwrqIfpPrTuoHFqGYxJ0PHm0a96yk3EHa3cLoLpnMdNG6lsbyqDv
R8vEJtpTw7Np5TosiLPKFszGEWs6Sil5TMbt/J09rSbJHPYG6BZF25pO444+REloOS5TjrOdkGo6
z5peFHS2JdkIygevNm4kHHLwOcVGxoHp8gC4Phky1Ej/0R9ETtuNO6pd42D+Wx6nlpf4vkd76QvA
VfGDn9XICgwmeI4fxSmN+j4PHx23D0G6KlodtitVf0Y9JK3KiCZoXNEOO221NgH9tqL8MyYm0ptc
YdhgRfLR+Prs6i1/ZOGyXv2WL6X4HWSMgazZfeqsQW8e17wJaJlKAXoG5Ja5K2LVC2QbZYb8lgDZ
JzZiljoTGLE+mNypMkzY8kJFVWi8q3f5Yh1k7aIMKN3srou3eoy3Yoh19wFqWXvWVq+WsLtJzIkm
0o1gUwmOz32CLBy1GiMgGXCz7rwSdZnf253yJFf41thqr1dM69hHXQjL91ONn16i0a2b/FQBSWTW
NH53KxfXUF707WUSabykONU9x9L16jURxPu8mBCy4MXSRcbsNF6qSA4DU5tYsLLXDI+KhgFTm16i
EFbeAz37y26I8xQDv0/U4GaRxZgZqyxrxHkZfmQFcZD78gPKpzRNDB2Ykxvim1spHrlBCbaExMYQ
8HgmZb9HlaZ+ERP8SnQ2Xlc/5v7xcrUCOI9Av6DlAnhkw1o5nJMSeTzNqgWdcS25vwYId36h3AfT
45ykFM1mEKZ1IkcqnShtxsrAtM3DXklCj7ltUM3DbIxUlVS9Dh1KxlWfbhL+6Q2TFX1utlhkfKDK
YjrIuT3wY8oIKUr/kIRQ8WUc1YREojYNXTN9jyPENfit0tMuSF4Bahm/EKSWZC3O4fBZFHUy9CHr
rDapYGdt0hgVlgIEbACn9OBQkd40yct43helL88YVaucPJJYfjTU8l7mt/SJHKpkHq13e22dIGZC
4tZqW76rchPCs5Hm+FZ4idCnY+hRvDk7hdr+vkwX1vj3lzDWpcKS19CxRi3UP5rapnRiImd5LjHL
bu7Ns3/Nh1UnHZX7mrJws9YvhBPrQ3zB8JtgTlJEgHgFDagTUxmohosTwY5QyLKpGrA4ngBFdhzr
omRl4zPOowXbr+6m0joYmdBvAkeFvCwH0ryYkiN7rF/PxVKxXOFvbBB3y3f/zvlKFPMwnPRNxMgS
A6cHx73c4tzWVr7SqreFafs7kehq3CTqg+rOKaofc9oTNXO/ErvvgZyPIsFbKlRiWxosIAMXpZ5G
lV4okSxLNkNo/ibB9DCqpZI5oTIQFjUJPCDz5HLhJMJZzvVIMjZnZmZvEWomTxUPzSVyNv/yvGBS
ZqhWybXJuR0S3C1GWZ8i5Z4nlJn6K0mnwrwZohoVQjiqJtqJWpYnrRUm0ZL56r6k66uKk74/ky54
D6iApWrgxdfPHu0DrAQOulSYmeVBbxjnfUd5mzB9k7oGkcPhJTnLyPEh0tGzb/YB2CE5cfVYPTQM
MXdmGvFPmy4d/OrM/ZSRRvr68kANlin7kMpYy+64s2REyWtAr3rYI0/2JuhJ2BQUeENaL/CeHsbv
LjBaI5nHjpk29nthKYE1wZ1VcNAKRzqtPirk8Ib9jaLEZkQj39z0R2uZlGkMax3pJ0Bq/2GDuMPs
gIXhHFzY1bIyibBAJQkTed3jGKjgP689WGennekZuC4Hfs6qNYYAXAj16NVxit/RvM6jFjc7Ybo3
GwNvsl11Ed7uQX6x0R6A7dEKiN6jH7NPagdALh4DAjAoAn5g+ySxRbsErl7pdJ9pLpiD8NqsFhCd
PrNTMguh4fo4DrcTX9iM8xjRyT1Cv4SHuxesBrCSIHd2ji4Vw/PQWOH86E4N0Gp8XSdDk82cbTzh
B3Oc8+4gBCsuCBLAa+qbutnbl0/5HTTdkF0VeUxgb+2pUsIUqEDqUZzRu7u3k2FVFofzeEmIOFZV
qA1hGg5W3ZmkzTIJgx3o4bXm7qKXWIuiy5SyMtqGAL3i9Eesn4sGMIznzDQsdf5oBY8m1ZCLksfZ
3brHiMkmKRb7cXh1lhU7ULEemLag8hsnvJcmKOfESmlun/BSmbQ7Z3ovdIObswzcN12o9c2bP+Co
okUEeq5yOSP7S97sPKYBC+2WUKN+6s0ECw4ZZgq8Fx7j4d2x/jigRPAQ/B/uK+yT+0XZiJdH44W5
qFcKeZRA0oZh0r807xjR0c3KaN0Rnm8mwn3LaBjgCxGHZ3BwnRBWM9xm0Ok09i4by7BO5TlGME8/
qmVRvUxJ+dgQpBj1IKfKctNgbDprvDNEpB8pNp9+N9SCrXNFm+Jd0qRs00Ry8GUreTmwJxc7RcF/
i47Z59B8p48U/iDqsQ3enOgPqcNd4eVJCfd4OUKr3PeG2CjPFwFaaYjVHGwvkFiXe1W/rMZXFef+
3ywlu+A10Q7WC+yEYlKi7NCO7JVflUNZMVS8UXB4fu8PJFGsZ4iJTRfRh5quUR8H4C1K3q4DcA7q
0jVBLbFN/JQMzSpNnLuouqMckZ1+6VA7YlG1jnEm7D/aBc2vsME7RMvwMaHPMzHMdIbLMk5G+4J7
GveZIQO16M9IqEKuceMIMlS3nDufOqM2oEpxXRzRCcGw6ysMByHn6CtKC6op10bB8n9MFssudRgT
a+YnEvhMsrZxVA4TSm0aDeuOkQ2jupkuPYDtf48G+N0id0OEVf5QC2TLQZhUPVghNlN1OoStHord
DoolqLjGLS2PspYq4F7ZnTEYMlFxrRgqJIS686PiDpkiGbqyTOCGaChAE/eZBkdQVCETzvOvlw0z
Cq1nIyehYsiC1rXJI/VujPkbUo+GLLSLpAh2QZbVzFKeDY8RzhLoeiN0KVmFr4H3ogd69rNN3idW
jbjcbrJLEZU9ZBYC93HOcTtUzOlMXrrrSJvkUJPE+S+ZF6iHv2J/01+ZIEFNOqiSOTxPSRZ8WXv7
YtepP8L3uDNRjXUoixzKVLz2mwm5V4Oe24CZQztM8uD2gzxnaT1ShsnZH/mylTzAdPlYe6lGk6cT
sb/hajsHGmyLrst9WTbVKSQwcpLKeFjXq64RrQPkTjuJjiGi7Lx/UJUGIEN/9My+l2XISQhiuOKp
yPmCBmBIY6HJMjtMPzLQfxRLrnAuo1hXuDcVf8IOj68e1Vs7LALcc4s59mtpFrJNWfXIUsQ8Gc3j
TZW/eJS8M8cpYlZVXgEATNgTknCAz0yKWixvsnMIaw6dlG+40K36wQKVHJZnkKjAQTEUvHZDz5Hd
6lhIOEfhmbc9lrLDd5cTlUUAKZWbTHKmQM9atHvh4SB7uLHUEKDLkZfnsspX1W4WwnfkCux97iOK
xLcAvoBwPt4Q8PqUgIf70nWVgtsVoon5qWLYYvfOIsUOstkzhjGcUZ7uioWmyLiDWi5lpgnprq2m
5Ox9/0w+HVJKBq3Glg8Hkojp8C+7dJQBSRM6R4bn8fJKzcSG0uNL463379lT+cfiU7NG/5T4Tl/2
aJ0kurM0OxEAEzH8iwoeelY+Ws1nY4TSb9t+ZuCtc6wHhwplpIM5wIXV1sbBr8+9e9gxJkJGT36j
TUa9MnIMPnCgZrHftW/hCb/SAMibQo2czanaC9jc5uNWBjvjYMMEOoZqQ2jb4nbwXkJkn4mUbCCv
Gb1cbOke47UPBc75gl713KWlt1j4USzz8J0em36HqU3frfBkQeOqvh+MRV0N6WAYGnrO4A6lsNAo
P41f470/8hrY3jKWEMj9Vx8bQOPJsLZ5B1DqYY54nZ88xj8GqaKNtBFElxmu4okZf6D7U8/hQm2C
yd/5RuFDGmz3W40oco0PmUXbY0E7PApr9peBcLPwHwipiU/MU6773Hcgm4QC7Om6YwyucrQfgve+
2tvZKCVRNXETEidUzMKaYc6HbUkaElPUIroheHXX2DY+9euUs2gbzCyFZcYO6DOH8gsp1tyiReWy
LEg2/r4IdyMOUleF9YlHE6AbiLb2Dt1N4j7kE5rg4PIvJRhIZ1uCLnA3H4pi4NskoJVTkF5Yu7gw
yyZXM5Sg67grIc+mdM7Ucpo+4tWrOwHmBrrVqFKhyQW7KX8q2QqKYMnrfm5J/1x7Gky0Apoh8xx3
MR4JU5ivV29gmXxIyx7o3GMhtJahlllOudy9ncG2esx/Rmcgb9QxryXvim0IS0dMte86IGcK972X
k+03uzSoPRGrFq6ISeamsEGhCITgde1FU/Zf5EaC8OVlbjxcQU3BfIDXxO14M2HtLTHeNlWp8SwL
/jOub0ExQjY4W4AMEbg9cVueezZKJwFIWC/RcxAxdTisJJwkRIfoXsOloBoSpdWzcCZZV0cqJebM
yd3HkEynryxvoS2Lh/DJtrKROkGKYJARr0ovkwUeSiVTdsirhhW4qFihChh2k2CfsmRoNmHCJZIy
JQ+4pam7LbKD3X4U7fy8ay8Hrn9lrCUdemJieVZ9ckIfYwoT/8IENBTPvVG8aSKRzYJ21GQVUPMg
UsmWsYpXYcc9j1EUZlWLDpj26qhEmtPSPqDg40AEpNhThbVMvPsnSgNF/VWpvQdOh0okwsx+vwIR
BL0hRwaTjMsYxh4ssZvUWIcXYMaAk+o57UsI0oUnC8sQhj1wswSJVY9LyVH74PEE6RZo+sz0z0ol
plChO+j5DY5NsKeA13KMe7EpVpdomtEs8Bs8c6+zlEcdZN/R15RFA42gHiuzfk+YYYTte5vHkFcM
rJGycvj88GfNMcGp3j9Dyt67e0o9ilsdATwwaWwnLfkAu8DUBvdpMuwpKqlEBhTulqTZuMuh43DM
3DBffBNTvM83oBePXyJqSIDAUvimI9ctYfp24LRV+ZMHY7rpAzA2/gES+TLv+Rkju22jk4SeSjab
9O+vxPWe3UW3A6HZbs/tldasSd8eHI8MQrQV2iHTFBZ0aFaxh97i4pT00YI4AN6DjiBLY/1npw9w
P4wEBA7Do21givou5UjoExOQrboLGkMOQRXTDSP5o8AwS7TkIo9m8MlCheGcTt6OJrY/SOtqknP7
/83MQzdAJ1Cs5P7Q3wg2VO/aWVoThXfawaMOmhjE9AReKXkhdLw/oMlbmaZ6BPAI7keJNyAUI/r4
j4qLqm6uaeVxGmMVdnXccNkXlWD9156SR7aH14uG73anJIhLj5U3zIlfrAqqxexfnYJ8KXyAw40D
2e2yD2mbDt7Bh7yoL9Kwek+PTxu+ZS4rAWOX5aFk3ZRiUVNIgQd6uD+ldvTHrOIoJJzII1kaM/bo
+tGWjOYumOivvSXOINvs0CIvRVSkCMaWQHVjhFfw28zf/cksCbL6rxHpVftRlAQzp20Vp7RdXhlq
Idu6gOsRbR4esB2vx5ihmEVkwPjhJrQNL7kW2ZOga3PUM7qMrEIjgVIEALA+Tyfe0DEoH1AWLezH
Ks2mV3H5X7vB68M1fYRlQ5CSvS5imtI4OAK/N3qe17khQ4DY/0uANHeG9U8DquV6qJQv3YQaEKBT
NUPMPgmQzmIZBm9iGx1Hrmnmsp9DnihlFJ/8/OxLr+uZMXjdb583ahU6evz6qEgebwn0EcmPREz4
Q61rtRpwfTS1H4NeCEIJBm09S7nCg/MS3b3PCqiwg5NjKC33Nt6O9YLcEsr1vwqoGqqCq3NA1/ss
DwMY1g7JaDwffRnjN0q6RSO2YIE02O1ZCZUwislXyPbOFERcxCX2yyYE6gsda+kmSy+UI1uBtPm/
l45VKEbsN0xpc6xQuNb7Ycq7mHNgQNFhJh7oUCVnUwLv0EDtgJTspi89oruNhkR3/AkUqDTvLd/k
HknwAx4HcRNLLi7eUcH3PMHOzouJZc8FKLpCwj7N1Z4NYZ1Nx8n0sejKBPQajTBBCoqSjjOlrZgS
5ifHo7pT9bXXjyJItX8ycqq8f/BGY8GB94ro8NlMkovaaJqy++Jenz6we3C6jKJ4Nw3wJm+0JDek
r5SQOlWguKbp+/GfqFVijIB4fShw+YxsAZwvfXtUcmD4TnmOudCTkSAanVUjdPJryWpEJWD4n+2h
za1s2ZNEroNl0rqoJoPezeVpAAGr67inLbpUWbgGKwsDlQrFIWieJfQvDzVZct+3dQvbbOBgTZr8
L5COyvJWxtdn8c0neNO080JxMSJsWFMAFDJfTRn/xOL0kr3+J5N4qOn6BvJu8X4ddJieE0sv+fFa
zu2aOw1AeBSpFahTYtRr+a5nClxihx0Hkx1Ppf5MWi92+mT2anTMSUDP2Z6tVqnqrcssNXhacw2a
bJQztxbp1XE5K+pCBE71yMKDyPmwlws1bfB07QTZmh15NuEY9pmgppENNMQGmrZZT0KAJAxSdTmO
gTuZWun/oK1o8jjQTIfl7r9kK044ZneCkTcpllChM7RzRvMGn7PIFnbYVcgOYq/tlHj2MdAa8rwM
8RSZjEYtsmK8adZ/q8K1gX8VXp/gQUjekJ1ZADLTAbC0hnZqqxxMPRSS1jpl2rni/KOCzFQMmW+h
N8Ypk30HVY+/tHXPxpur1RB4WgayZgorM+859BXOivztks5fT3zHVPJ560sTZ2GezwCUWF2XAY2J
Jx3zdxmEzinxs1cgZruu08pcFZf87TNRMcEqaAaz12UQOBTTX81L6FoHfPIzHFt2vj/dMTATTT06
bZwV9iE2NUTi0GALj3oHtbqPuzs2GzcufXzUY8JF3F7+liWaEiI3fghOIIC/KQDtZbkmIu2SRugk
fiRIq6Vh0f4CAf9/hFtWowJnB+eiOJfqzO7gez0YPPrC6nfLtsR2C/rHlLFa90ahgfTWSAkcw54n
VU7wnT5npPeQEFRWhthjRnGN19l+1A7Lcm345Ja6GrVnX1Mvkbxe8kUJyVwkTZaXLGBI+EE36g/M
Km7VvjIwuZwIUrBe9qfGQs4Vjo8tl/b8ryoA8i9R5KtuY8K8TvHv26cvQw+4nD5evtHIKdcZo+L0
56RG7rBaZ9srDc+Gj7+krDSJrVtd/rBKwXc/jenTxjNN99hpd82SGT79+Ssna1UJWMOQ+KhrHvBN
f15BTSd0K09LSZxjBZnmQOtfo3nVqSPn9J4GVqJ/LAdGXwD+UxOOFTQbmwXzIWTWCxeJtE4t0Qb3
CR6aeboIwFEQoUhO8nVJ4zuzP6j4w7BLDI0ZbuSjGcbkH72VaL+bPjQuiJIhJkLLK5F6CadHqcQr
3aM0ZYxWdO0n8/s3+QrYti5Ye5fI/Su5GvBY0aO2U+lc1CEj0kN+3ybO7QdDbPVUfNdEJ+qPxHWa
2kX/YLW6hsmkpTmIgCoUuyylguRrxhy1Wgm4qKYogxq426xsyotklwhgIlDF/h4jBtPhR8fo8HVs
4pDXM/XBBQTI/imJHFZxskPNAWOHX7zoIPwtQwPjwryxUiOSLO82kbR0C6VJOwoW7b88oQ8saMSW
HlaTngF2DtKeIXp6MPo5qkvJhMSy+Atyl74fxnC4ZYSgzyv/eZZnrokx+BwTtuoH8gDsyGz9ezai
fgF3dIoZlVQ2hWGsaz8oWosLuAoW6hlwOc9Qc87xZlXzM7MAQH38YTOTJfvvjON9Nr/X8qg05/m8
cn8fPQkWd42U/J2Qxfu0I8nlcmwlOO0awfFkRFk/6KDtDuVFcccNCBHQRrZYAtfbjhL2QLbno/vx
6PnqGlqnGFc8A2qPnWYW/1Wl25v1D6DKG8bq6SX0VieSP21FbBIS8Z3HWFXKBGOx1/6i1HardiJx
FtbWvsU9bhuPcMXVRpwtHcIz/an0wiVgjTXe+8Oy5sKeo4iqfXu24wuRHWcAH8UnV5MfLGruEzPg
pQR0UVTmwoKHsQ9rMIrbETk1c0yOQq5yxhwt/q+xLW2t1NkCQQ/uFfb/Lm4C7yVNx6Q0xO2yDv48
LUEBIFRZz8Wc/7bYP1hFLDCPxlSuA07qW/aCqhgBI9Pk41RSa8vjkt9TFPn8MyOVGbw1Ug5tfCmC
4GEWjPr+HlIaKygZ4gEhLM1sFjfWCuXJJqAGO47wvjKF4vOm9TvKxq94L9Ghxa04oMeXndlqR0QA
u8EfY1AJUvrlg1zLXreHQdS2ZAq5DcOaVnJvZZp634p+Z+V91q77HEsyXYripxRQNYWrSFClWPTi
iMiyQPKmMOfNkQ0S9s5PXWUmBrscPuz+2gZK6HPPGXjV0ctATEKiFzL2OnZ9nKLJc7+30JBKvlXb
/3vyfJhl/k+6RMbnRNJdu7D0pp17NCIUL+Mik7d6wRTqQPJOqa7QYTh8gPftVSWCX3y7qyOiyU01
YRfXhxxPzoD9kPiuBcmZ1F3MBn9QMIHeeMQhYiVYAtj8iz9MV1W11gFzUywqx3xrVFOd49vkDUTc
PQZsdMEnOFFukloNnvt9zQ1aLgAt5McsDd0UJl/0AnFfvL4gw0QGwQ1PD6QnGbLyNsKgIg+84Vl8
EXU3VZcLSw9TR2U1sv6yLOIvWVJ3YnKzKA30MKVONpcK3ErC6RXYt1odievNjJZuePffE+Bw2RTQ
Stz0n6gIb6v3ijTLRA7byY4GJCdSNRXbnUYKRjbbk0BQ0BvTwucHSbT2yzNXd5LNg0b9QgE8dUWd
E3+CdN/WQJXuIzEHgO2WzwSDy3Ncq3DJqQlDrX26MypBr6qgKy2ZozwJ6gDVRlq0RxZot3btMAYA
bZPuOnNn2eqcLER42En3ENxEoDiLTOmpFwGIcEXJY8a2Hpp1k/mRnk4Us+PNZBdMqTaUGETwmnfR
WJG9L3BZSEBD+ScFpNQnKPearR/4wxaj6uoPLs6jnNbINHPu4oMcIIOpv/7TfaG2c2reBJhAVJMj
dsEdSfK4DG+nKu0edT3c90OClzevZoIEr1IaRoaqOFfyORfb8FYFdJaro+J0ttIO5Pm/iMjmgh7T
SAkR/WPeaeH/ewbhRLSIUKtVo96I8rowq+hSq5gDGwveh/B3v461wB3dsS6CyhiC370CvawpO2Ci
ykwsvu19+VNe6sFmi0xUldmQgisjev+bFH2VDF2BxqMeBIchJON3giVoQ57Ad6/Z0PI9nMTFxJUS
HUMdvkvlsOUBOmu4g/+5q2eWDfvcfpz3lt6mU9pX1RwxDZNbErT1IGm9QqqRFC3RNtF5VdVPX+TR
/K1gbBdOwxNpDxAJ3U3CcyUZoDYlY0P3jz4agpM/VacZ44OgxJoUPwRz8Z77iHmBfa4rSBo1UEJV
h/G+cmjD8sszOQIRaYO3ibvoaa/vinV6hjY0RH7AFtzQpDisNtCWjNF+p7vl0v3S2VPrF5xjWLnf
N9ZU81NFgakkZItvwVTeNlyHnE1zXSOyS/cICrmGYpmijdW7QbCqHAEtXiqIatrmY5Kkg5gh0kCf
dJ259RqDPhfzZ/2j4yPBGUI7n37kT08QCd2a3tltXcjDW4nOjHzUQUR3MnsskTCkg6UbYRHw3ciA
Q2zfyqKOkrxUveg/z4IIQDAR4hFO+WUnK4VV+cLdrtfGc8vUESgVGc7normG6pJx+TmU/nb8jnky
a5l2ZNAwGZovCF4v0hphltycMJ1qhWqbWd/f8pvV6vEpx8V7h4xTqfzSq0Ms7WRjfvNbgymICWcm
DCIH8P3Vaivq7p3Xib3eqm/dTgtXU37dLp8C9oN4scbe0pNSKweBd5TupqHulkbWKVowcI5jcFVv
cy7xMKk/Gvhp9ZBFUAdIWJKKlicXI1aTUb5OpCAjItO97M93sUyoz7I+PWTFg8L4kSGOqd9+Z9Yi
zIInhV9W7DmNHx8GBbO9aqoBXpUtIIT+WUaN16f3rvfEJWg30+CW2Jf+kNkvTraN+7f3QBO0WhLW
zCEyIeluQMUST9XwIO39X1ZulfxQ3zUEx+GOpt538kXQDhiuYjHN8irCcz878sVEkTx8oMNJlmRM
3VckrVx7UkkV9c2mUBy+vbsVqm7XCsPkvgnrG6SXt1iuFjJwPUu0L8aWHIz/UGrgB0kgS6GNyKT7
hrtV7tujapeMgB20/gZxJ1Y55vY0qarG9k2CmB6MeBsPzuWJP/XPhkbyI6xq+QAPv3y48rPFsb7j
WY5M1AROhrZjA7+j5iv7vVQ3cPeAnEbhSbGsj+629Fz7Bg11TMRYZcBdyiSNGw/5lgORLAPW/miO
7NBYkxMzuwiujvPXcA5xEzwptNDvGTyH9oLdgWPneB9eKDNs9TNpBHWtqFljCYqjEWfTC+a4VC3X
B9EzCTZLsCcQBUP7H6W8F4U98H62pNq14Ds+G4gMhrIr5MtSKIaoVzTPZ4mRMQXtWkHieP4dldZ/
oP//4XK0uvQB9B12+AwjbCzH6cAEl22/gA+P0isNkTyS5UrBuMXPq7e8IlIpuiuDIwUinL5vjA9I
k8Of32+3Y/juRhmWQMr+/PwiTPLzumYsyHwSqxFdwwJpRv0QczhxhvYcJ3alkKGCApgNqkPNStWX
LPqxHthRRWP097CkJ/D3EUl+u1wKEznvIrInv19bL0B+2VI1LyDjOcZSyHQTltGIfMl/ezplJw2I
YkZLccGpWmDMZV73qE1DATu4PUVQKKI+6Eh5MwvbLfsIa9G3CTdt4EVEx+XfBwVU7EpfBzEs8c/E
ugpTWggnaPuCDgNOqep2IO9xoA5SmB5KIy/hG7PGMmjYLbAIzq7eFgdcVB7aXiQkdzWuH+sC2YAB
9XiJRWK0XBkB3ttWXRgZbTXYcMU9AiQIMw0fhsdD+kE16FDBCbCrGbCVyT42z7duMJXOWgiSjNyr
fTsSC6ZB/Oq5gQCq8cEbVQbwFnraL8Co04yQn8kpQ8i7pxXL9rVZHBljrz1krDZT6/jITx+DcjAG
3MgepaDKew+Q0dOxcZJCVEnDO/EGTe4P9lvKnRUozH7IBT3XqsJAlKmELWSZanfoIhNJ155X1bj1
Fca/NzUe8RotYnmZl3dWfEpfUXoaAK7nS6H/ooqofxAiZ6dXdJ7cHEhSkCtFhLbDvZdyjkTJ0dyE
27sPazPHvrlCJgSD2dHmqzpQgne9HPQwiW6NTPnASgN0x6aZ6Ot05r0U9SvgR/Zf7TjXZ74l1c1j
bYfIewKYgpk0GL2SutrzHbrafoh9o5JiIpQIJESS/Q7EOfMgdG+NEqEV2Oas0dG4h8sIJ14mqxKj
Q81tQoRm35ZLwcLJKwiSgZk9i/5ReYNBbOhu7r+bcFSEdCoMQ9e6fdIkJy1vIjTC9RdZhRox3cY1
NQp8pKCK2iFr4vsky5OtpHeEvzIJM+OYVsWX98Ltb819XPBd2kJOr+uV0Rw64Jcu3HvrIAhtU8BT
F//1eCu4tKgo0dDUGFM1nnDo0vyVkbWSZsrXPFhnHO0HFU4Rd/bApAKvzHhviKEtfw8vNRDQs6Qz
y5n/720+R3eANsHU4KTpSCboYSh8id0corj13FUA26X8F9ha+FhMz18Cp5t1mDhAUSEPAthwGsos
/W761L/u6WkliagLV7LP7rObbcZfr8M4S1mtHqBxWnGU/5bT916wZI0VWeoYYZFykx6+5gfOBa8h
ctPd/KEAPpOQRTBA0m3dNcV3fud0lrDh7WW9GyG0x0cVdviCLYwYwyZOa+781VeFWRKgqBe2iNOr
nLwdgVnoruMijMAiRVcgNYAfvUwkboT3UkXUItUbrL0ZgcaD1333tUUb7cCMVwWvOMLrcVYF0N6J
V0QeDNr4GRLwOIqJwtLtRad9Z/ulm7rjiqmFniZkMx2Z7gDlHroJuKJ/J2JMe00ouIv/PYh+tBab
7Wp57d8Kl/SAQotrTl27vHisHEQLtV3KqRBffUYPEHQ6zpXw6ie6SxnBLRt4R9xAEJKKN9FC+nuM
rtiW1GkyfGy0NrvkYNEQmn/q5qRGfPYn8LuWHPXxHxW5/YvRuT7wrPFkIgzsiwYqHlDdSXEdmXRJ
0tWsLLu9WGdTz0dyS0PW1bj+G66L+orYGJZIxc3ADe4CmUvX6Mb9Qkl1xHRFgRRJfCng8hqNw//5
DvCzdw+pOtPtdp+jCdPgJ7S1kYs+gydmga1uESFmhpcvsdHgnS5dsKryvBX7FtxXut0U54kP1bgq
4tnvCdN40tVX4QlHjYJawb9MQFvq5mefgNdnZm+09cObrlRxcSBBKF63qn/ncU3Nl2PRmad00ygm
IoDEubPT4UsaYC/ZoQu6sz0g5/3SdWReLGSgxxhQ2JqhCstmySUlDFeG3/RL2seAW7fu94hAEzGR
6rltFao+bW20bVGtcnKxuTHGXdb//ZnjlahsCuDdoZNnFAah+QXPwWIS7SkendgIIhO1ep3GdPtj
JTQZtuQQMIFq7FAbW3pNWpp1XwrV+yUIL8GQszep3883qVj6NY8XCUVVHq+dXsS5zxJsvGqI6nEp
1pfGm4jJSWEsQP0OxW3U5vtVa1jRiE+Zfsl3wpG4mjc1TZrYO5ZmiannpF1c22nbnlg3EAJ9LkKi
cC7/336p2fOffanIAaH/7CTHl/h3OIcAXyzPMRzmpHMwWhWNoa65uKQD1I42yOcJKKautoNn2cB8
JKyMIYLPxnOyR6ExguZLPLxMWi0UWY5kutA3xGXyOnSTygENh1bBDpopZz7Xk45M1Tjc3bj10MsN
1XjpPdQruIgoxdtYVP6xjxYkCWjAN7eu4teAN4X3xir3FxHVMR4jvxAhBQx0rEkQ6lFnVY39ofGq
jEooYT2tQkcIBoKsFYmA+BfOFf52R1jx9nvmzDfUYJUQ/nkSbxMRcOaJKamxJpX55gxQMV/01tHJ
ViuaOYF3gHUoFzwwoDYrMQuO/wiYDMtD0yMoRyXbmFL1et4YA7vwhGrRRga8JN278K3m2CAlLFSG
z5yjBhQVw/UAsnOJfO7SmddU7PMXmzEYknh24SDXvQNOvRAfxupedymLuu0SO+3+FqgE8usASrgy
93vnu1dwvijlz+PAaho9GTyDyft9ViH1/nWTZtVr2HYAxbhfdzczomVW2VS+GaMs/czxyWnaf0FR
kswHhWaW9O3Mqo3g4nAfw6D0lD5I8norSg+1GFp8vrV0H2c/5gp+WgO06qUYkpK9JA34QQtedAE7
ntiPchbOXKXCuBvXk9OfQPsaqxVXEuL+SbT4OyFOljXFCYn2+r4gYsniaH2hhjFXVEorBplOdVn6
f+8u+4DvjlC04Eo6UVwe9Zl0C9825Id1cfKDhhi8SppTLU/SULA6IDKpyDvLDLOIfXzzU5P4rPrL
9AY3of68DVUO8LYyU4bpefn00DbuP2Yfjbdj1SqxhnBkx91ParVm4OBGcHbqMKCNPy0ek9M7T7JR
JdUbED9Yt6i2DtELULb87taLbodk+nVmwKeTA5JHoqYVrdwX6OSple9zqd+8KEK/Cv10ANwz+p+2
YKqDdB2ORBPNxVgl5iGSJkmjZcbV0NhaUY9KArWPQO5u1fNR524o2cm/SwQE9wAUac6DcibjLGZX
ZIJPLTaxE7Uh/PqgKFipjq4HIELhxjNIhL2sUyl4j2hR9Az10/z/RWY4TsDnyIiJO+o1qSm1aEIr
StT1NxtOsYCzZPhf7G9dh1HehdOF+JReVY68YDf6EweqRqv+c7lmtp4REGYGrqlwuCI6dwe+dYZo
oPup64HZxJFMldDpBfABHT4dVyy/1Na9P53Fpp5P93ln00xJys4zJYork0vFOvrUtgC92Og6Njnj
kJ12UsudZJMGzQ79Y52dTB6PT1ZMAES/GhgpNpAEEAgUErcAuo7niR8rUMAZqV5TDgD0F5wHjQf0
9JhlaxsTbkbTkLcwNJwpLUTZ4KDJlAFfMeBwtpLgIyhe1vJBxqe46J3vSEbalzyh/jsEea9gzcUY
4yV4w+Vxaax/h5mvxqnb9S/KWUFEeDiHPP+pCxx1Ntf3hqJ/qa1WfALSxZWUhciiVpi0k9SQ0npR
ny+SFQbi2vPB838H9Itz7DjgguL+ErBXVMjvORDRwsbDdGzAFxv0xcDfRCHJeMTcyTv9Um6b/oX5
X9eZNdFTTEfiRDsTO8/0SbLNYfFVuiJQFyG3JI8SA3AJZ1LN7g7jgnIOGVbFVVlWJl7//JuxBa/D
7a1Wdn9xsAllteUazap74wDWk64AgH/GYG4DZ6XS5oNMu7SD86lTD6nqmH9Tvwc+snCaQDEDSq0N
82qBbJWxIzEXHWaG3woiLNVTgMrJkHx3E2IahlNOKl+6bzF7yTNewr2aCqbl3zxVpcLv4RmKXhgn
YPC4HImwY5tDJYSa4QO8jMnztlDMGdLlthIPl4MdUF7/v8PRQS8R6yiO2nOnBaHCkzwgxM+2M1dh
kbW8Iked2NpRdUMp0NjxdzCDthB6RLN9fFedZQVagv6qR3HKnLDZK8jPoLmwAS0QI6spKAzE0wwV
I389yoKjt0tZB3qO13xrIkF61B4Kw9Uc1mgNL2VnSi/srTeE3A3Oabur7PeH4urcZGTcIDeLGAOr
8NL3UCaq2xm021AXTersPQOYEpuYtyvJZU/U/m8tjn5PTP7dpeMwYpo/FXxhz/ECtqXufI/GaYuJ
1dJLOs6uMowHrtEd6Cwg2anBXy0xKbeVCNp4BT3UKlPLI4NvGgQp7s7Ty1gYM0wRw43xEVoaq5KD
DcaVx7qbJkKiSq4KUjlX3cRgMGER3nO0LykezZXjiUO0CUZLRkJmLSsT72ZZGAhZ2/OrwM2PKNlm
4YLsjkSbRgzZ7g3C1bsvJLimMKBIOkHvdNItIEefoU36mfvuEIY5Lgc/YVVDFabp1CU/1ePjRBDC
bfyfp32Pia3SnwCBrwxo9nxrPsbuenfhX7MX7O01RoZB7n7D5prn3X4s7ua6Pv7iuh/0QpB9iuo8
O1G2LCWQuOA4P/jddOgeENuQIZdpEiwzaenN67HA4MLdHjWfComJBS+/U3cT+3gX1XQlk9fWyg7z
e9XXoARpL32kIRTBHPreddytC7PE32ZxFjsGeQbeNfLNPgP2w/6YQfMsNdw7IPXJIszlSfVKSViC
zjzIL899eGbHBD2CKcBJmP3cQB/Scc/nyg2SFlrDduEhO/dtF0foQQ6oWnjHZzu9iYir2zIVDUQ1
NXAiiwBjYlGqOu1LMAgXzVgF1wA1CMf677XIIcguYhAnYF/OzA6ZcIaMtWk5IBITU9jgKqn+Dk1o
gmqrj3ZYoEBlGdTlwp3/xh1qiUAmlzWP97vy+6jaSsOXoi/G5L2rvEL28wD39i4+FTa2wWT5os0u
yyoJcNiRXVccJP5bjPMty9C4ikvGrcUq4QO8t1zQyYnuEX6zp3UUZE5Dh1d/tRGASnJ9UZOFflc4
QkdvEub+3ZEQNH0svVIx1a3EwkXhoxhCWfm4HJ1YOa/KpJXc6ZWMlTI/ay/pcMv2+zXX3C31or5E
tiqofsFtiQ4oP+XFJ2zNZy6qpJaozJoJCnLeL9uDsvAlWwF4Gn7FaCCaUE+1LblvuT51MDSYdJTT
RD97B6F90HYiQBOVjWuj6FvCWWPrXwDRobmKmrdLgj7jvLP6YT3cEnBqkF/8UDF0V8P0C8m2pVr3
rBC4k/EvY2/9hRGqAAX14yYN94ssLzdaN/t7C7EstA+YHpYpD6YMYOG/VaIeKK2awU/A8/aNycSE
3vTBGq6hxSZCnA9g3bKyFqZzt5aqfd2LyTaY0xcAqgYJvxZ2ATuhnkzSvxqYbGDsMQj38yV5CaPQ
pyQNFHxRydnfeaI+oeDhcZjnjOnpyTTzwN4go2K9FzNLlw4YYDyzq7WpGMf5iMmTrgu06THfhD1f
P95zj11sIcYQR4/5sx+HMbZ7MBEzBniO51SmUw16YnI6BNU+7hPvta/vt795SeNABZ+vxU9e9L2x
4FgT1/FXuj4Jy7xIUQZ3jZ7sWJ//4yr6WkxXlbKFU6rfN3Va0VHrNg4fLHog+p+bRpTR61yo6PAB
tGwuNms0Ml49JvB+oSYyYNTFdCOfqHxY5Nqm6oVJZshEkOkAwxrHmDY2dV1Cz8pzLrlAeomBYko2
pfqfHBy935mf/3MhWw4AOGruPQJVnZPj8wXGa+w4BVF7w/tZ28WS0v59dbdl3ZJ4q+MeY2GuUFp9
BLNXmL6njGeHFilq5qaY6xIuL0P1+/vJx2xpsXMfheKC7/q9tP4FrYCV99LvOGMNmCyOds7vUdRS
jVK8FYauPQ1BKMtICHK4wqLlvdC/UnBSZjRW7rOzzRm9nyP8vT5/gvpJW7T9J7R6ELQcKgrx79F2
XiHILMTM+CMaQ/PSD4XT+g3U85Is41AuNZUEoi7BUKwCezNpVKevnC+zth1Z5hF4GACK3IRYGLAf
IBF/zQ2PWIRDJz6gYonVQNwRbthOis6SlT3MysB+ScWzkG6Fd7uilPSuPCLlLRDPfr13pKJJZDKJ
ZhZbGz/CcSN6tNhH9X9hWp/FDRcp4fFqiScjlX2eYU1qxmq72lRouomNourCW56wrsxyQVPDY96d
IiMWJipelWo8aDMbycG2GHUzPZ83ulhfb3/6WHjnnRnqMI9iluReDJam9jut4CzjamqKP+Aj3E1u
T340eSTAqWOPwz0ORvL9RVCIu/2GQ9fCswiLTkmyB2+jAfanvvIMb7HadJm9a7TlJzwrXnUaY1Vu
TvcG4QHHcuFqx2KCMkCaGjWLF0hTlYVhCHMmLKFDVsCNdhwFOEcydVkMbf9hO3iQaUzepU8rU/YX
i0bsR4hCdmpIV8G+3X4E6lkPfEx230HKQ36g0hI0ZA0bhU9BcYc33lz6Y78kIGcFnIHc4sPMnBAX
reMclilIZHdIZ869twTzUvg3a0JpN/7WkBg0cBb6xIsYnO2UnT7Veek/pPY1GS2CKrmDys0JFIV3
dAg/+imLqXGvMMdbnp/i+ybO4TGqFb0fT+/GiU94Hp5IvcrrkOrpRVrZUg6yY5Phg1zLY0v0HArm
ial0FxuTe6ZMjcl0UV3oNBKMJte+o5TuJNYOORwNcqXaDFchafPPDu4ReBItgfNDY3Ufc9VuiVEH
4JodIjC1q2YCqwIZcQVeQnKVOXi7jXlhNys+75JhjJZpEn6nOGBOf81lTLSMkT+9hEJqeSbaoi/9
rgqC99EUF61iq0tngt5uPC2tNeWE3GfkvQCe3pALH/Z+CYI02n43ntGMLD6g7/nlYeomdvTpwyBj
5sF7KgvzzCAM7d9wwBjRFoGNIqizfW3NTFlU8+Y1+FQQpEOfd3oPrpcf1nqPdgYDGWjj9viE9XnU
oYDwQaXoDKYykeGPFfBxJ3Rc39oAb6LQFvC/ewOizWdAp1iRhYruqXT/oQ9t2OlDokM5UO53RSP+
Mt4+fYP83bWWIummVk4+bphbyO1WERmNQnFpfvFVP33XETF1z8gxJGEdk/VzIPOgZp3INy7tzNG1
PomQ8C1RAhJEaoVVVh4Age3EQbClzEC/Uo7R6cJC4OEl4K7sUF1z1+j4NOLkvXI6U4dw3YQdDaPg
eEvPFHl37NuOfMqd6SMacCeaDlY+KNG/zY5he4nDw4Q8A/JTOxO8xawmYsv6yiGAxPQMayCYfqbB
4QZoxEBEnjJQAvX8NNgGjCbAYKyBrsoQTFIloC2DmY860cTOTRdzp2gfvzxKlOvHwF57loVKql49
2jxB59bM5TnzCzSrNBAEG4t1nkJSegOo55JvQeQqkRGTy8DIVOrw1v8j+GGsLi/9hiG4BKapMzhp
8zNhYjj2qvCWQl9ucV+L9ix5nZ7qvj+D6ZsfWNt3kozSIfDZOHK7x1jJT7tftvQQcR4Lfljk4rLH
2YEXtx7/USFPaEzW/g1lhd8p5Tk8VpIFh4f0X3mALW4kr8xCVROVJ8cRc+GcaIIjNbcEkCGzl9Wb
DwjoJtp/Z4tqpMGMqA6+9p1aq2wnTivon5eZR9oGqgEiABXEZxnB0/KESYN93aPaPgxTzTemMiy3
XxJ4tApwEO9iFOJO+Zwo0ctyk9YAAgXzwubIL71lOuvwBbfqweLpMnqVYzAxaiFVG70Hz4UvRS0f
kB7ekrbHwP1PrEDo0fxFhEAebN80paFflP2Bl9JuKHc3rUFaoYbqj3kYJ8t0RTRLajtRKavb+RDT
kB1cVcHY0VtJ6c7M9igjcK2PfisdSJuUKCeIu2OC1Nk4XNLqi/Hg51eKZeuXi02wMVJmPGSMPm+/
y2yzdzAxSpktES3wU2pHLm6sIYG69EqhtFhLbudvq6CP0cjNgdEE0Zj3qP8RoXFUctF0dt81mO/Y
z/tXMQJxWKozoofHLEc70vxfl4z4icsYp2FoG+Fbj8dpuPRdp0ETzHetp73PptXnGgQ0nVfInBZb
stX9frrTgzJ7Bjq2jxZefmSzHvEcaTR7AViPMo0AwTce7kWRRLPmBdwXthgwUpuDfN89GLGZS7MD
7j5nUwYhX8olDvTObKUYifKawbAOc91Mmb8LAsU7nXcsglZHGhyhcyjja6lzFU0NYirV8rsfTNLl
ZkM23gouFrYbecTqefnzgrOm/LJ5Hosxxl0S//ZdwNes6Fhfn9VIMgnsBcslKKH5xqRom1ljlZ25
fGZIApBiyVJbRS1DQiDyZOGyRxidl2qaMwySKX94RRjZjN+/3Jb5RwJlI5k6KSwlRKqlQfcl6xwY
3gOtxXTXElGBS6a8aVB9luE76lfArRW+pVJN54jLBEHPRrhH86EwMaqrk3XWergYnDLovfkeEe6o
31SmXNAvsBekkUsc+dyVUR2hnRV5YC6CsyOAmaOlYtb7WN9ArqwsufYljCVMp6NqlcKTjk4BLKFW
vIMu4iwcdiNO8aPHUUYL8PJsdjaPhGUgA8tSpoN0sDASdg83H00lS8litU1pxHGdc7DJ6nHNwmYQ
PXuAoj2JqQeQM5UR8HAIpg7CvEuy62MFnKaoDnAElpShim5fuf/Sn90GWWWea7CSgHxQMmz68h2s
XpN4tqDgwF20fhe9cjW2/xbeE19gsLwJUg8P83UpMcakRtOAmvYXEAXEu5iO10ef3AUkqU35OBtR
amfGXQsiCLeWKOma0qJaX0eFhuCcmkE1rEebtar7xt6QIotOsnZJvqfJeJWOncIa9ahmR7C3keE0
jSRfkDtzu5s2thTPZFPcA5W4eD56tA31fT6bZu28KlTt7kL2ArJn1pPIfgPGSsRddCXC+db5g+1x
a4K60aL6T25TPRe/SAmw00vQ5CKXnHAu1uHUxF6UyJrK5mKDtpSjGKC9X0Bv1sOKa3mPDdlUVYVP
+b+Es3VY55Qag2oWFcqg7ZSAGzxS0BVcbE1E/ii4+NErsmz4M8XbZsGZJfpZGkRSrxxtPsw7BR5O
yLyuISG/yA0yHzGijnVWhoQFFLEodfxXcGptnKb3uchU+ML/RMvbi349RzvLEK5LSnU8+vJ2OvRo
YZTEPBddssYLh/G+OlsQXJ31BGL2ZHcXTP2VlD6cscdQtfqJQ7ttbASVN2uCzpVBXIWeK42MOU4w
Jo6uZGtN/HbxwYWt5uMZIyvY+huQh8FIcU0bxPpBa7Jusi2eow1Gs3wVY7R1scSxGUJc4Ldfs1Nx
Sd1fKBNbIOFWLg8ZHouJNTKU8kY7Aykm2x+YKFSnZ5HxCQyM/ce7WRejkNhn9GeGxPKJlP4KjnjG
h9wij/A5px8R0+2PAEUuisA07oHVHwL1xVBwIhrPKXM+2Mf/cG6C+AT04ggJv44yTkkHwDoVtFh2
etkHxmThc+iZvDRjjd3hs8kH+4OCcs5sjaIiHrGKbEli/xrN4RR2bR2QYCHPSsifm7i57xaqmGnA
wAKVrRWpMiNz4R6S0NXz/VkQGL80Gs9KnUpRTnEk2XuVf0HOMXi8+CfPg68k/8MxgatH7Bp5jkk5
mBxbI2g1ldiAzsSUALHiVCBw+fbIP+JiS3MR7Vga7TBynWlT2dCbDPwr/1Bb72BDcYZG7UYQnFwO
Ro3JbKtGOxd3axkCvtJI2YQMKBy8+zV1XAIbPwM7NP5AJwORH+wAYTGvLbNhn5Rr9/cLzv4Dt5Ms
2UU2cTElJhDsHNmWymMtt23FU1s61Uc3QoA2CvN7HAf+ZA/4qc6eZdqm/DruRGE+6pTI4ic4+ltp
0b0SMkZz9zHkGymtQESRC8WoVT3DEziP4BQZGssL1DsBg9UGuvyIZDd7NGoxeMso5CBS1Vba/vtu
duz6VisAwxk5t6LPsbSGA0uGNllmtN79Aj0BNtVO3+SvkxHHApd9aZOYhQyQiNzbCR6FJBXiVICj
OT7J7ryxl2jmYNULSBJD4aK1sorZcGhwPXn8Fl1uJEICJ07Vr+Fg3jxxKhpF0a4d9xVgpy95kEC4
SxpUXxscigxwohp/wlQCi7U3af+eIr6kPfvzgBw9gTD/6tM7LHJfmxan+qJmCm5fcmTN8daRtKXf
xzIopXwVA+/5hNqu1zC3IHkl4NrdI3faU+UC4eSbzNsvXnlGhYOHsYQajwCDe8mJzW2/aG5C8qwa
6Hvyu7UEKCTAzEfhlcuPSvg/gSDiEUrApwcRDgeplolf4vfATcrSD4FFyGrHcPP9/VNS6YmoE2T+
CUuJjRbJ/8JcTQ9dymovXLFlGndeV6mohK9mPnbkQqmxYXoeygsjeiHOvO6eZqN9Y7YGU0OFywjf
gAB0E0ptMD5i6sazFnThRxpvg7SxWYrlVhpwmeeFvKkwYJ0WXCXqvHJYhtGG3jPaXa7LkP0FMPLM
EDPCt7A4p/5M2ohaZ9UxeMtu2erAR8JVCocWEYQODmfP6RhBCzoeY9OYu45HizNKOSkxRV14BEit
l1gnzhBIYaMj6WgbkfepA0/wtUFEv9ts5SKAahLTFqmcJyWuklvuAUa02FlFdE6N91/2RadWg/j1
gPTkQ4lQxHxak8GlQRmwyY1lhruzRXfCzedQpABzu0/FpTBDJcmMxgkNUcJ0Bs756+LdARVwG8x1
FbNWC571QiK6I+A9/YgCe1x/GzhQmzi9eAr7xyWyAsK4jFmKYEAgl7JfY3137oVQ3KOfN3PCWTeo
P861F8edG1XDbhHw0q+6Ers3B+l8X68lRP8SEyKbFCtqPnH9SlLOw3Vs4zg8nqTu7wE1R9BLpIwE
5pOSTSvjvaGIrHiOVgNxV2VXVlI2vqYPyspcZvYqPFOs5LJhwx/L3Hc15ZpipLs8a7ab14aog7Ep
BL6phHQO7c1Hh6LCOVkc7MngAI7e61P15yknpdb+dhAadSh8PFMsdJB4n5+OzSZnbVch8MYyMeSX
9npVjePcyvXN2LOfNqODuQ1fakHogfWk93GWrpYmupQ/qaI0riXDQ5IWthkuNqlu8Oqh1eCOHZ9V
lWuSE2yDyKq58BnYJTJAq4UC5fkGPiDlm7eN8vesqDNGdqrumI3PNEmK4j2jByeOWl8/d5aPjgsf
xoTbRMyw1zvB3laznuqv5dPPUTgfHuf2INstcGKMQJUn+VMBZ0FKuyiCMK8tg0hmTDy/IpZAWI3r
UMBwC7KMn592BI3dh0/h35FpqMTbfe+SSVtVw0Ybf4pBCvGguShSBOGNX2ardPQ+gdfnbtidUv7f
dx4xp98yEGjRpc2BawMmw3amLQpyYQPxcSli/CTV7TDt/Sy/hmGNp+izDt/zWVEyaYNbqV8RCp76
u5YKYvEJAtlft1zU8yRl9NhzNy111xozeAoFpJV12fIQN3GHHIzyNHrI6FFMxXer3ckylgw7bBks
5VSACcpm15Mv+Et8xwWf6kNWdjCzSB3zVmAE46Vcj0dzvDqk22nWOQG+QODz5JmuEpbot0552Ssm
SBgi/BICcHkLRA7TiTWKc0l4SoVw2zGc3NKwEvzGzWzJ0pesL+Yfi3ymbEp1IAYBmEkEwPNSkMGL
SHYNyDZr461Ea4HdRg8LyTR+yRUGoLN1MeomhcFldAmkJl/7cZJ61xgQ14OX3CWfu1XZh22jMv4m
pHKaVpsCERYnrS5aEEQeOXPEDmX3XnLoHHNeynUzSAdLbr76/bkBqWQ+fof8v2kt5WkvsOgf9jRG
Gqho5ScJgZI277ZY286rYrBzIpiv9qUMCMINaIx2LxRFelFeH1UK9WJ0YEe1I4AzZM/uVvusqTsH
W51kif+9b2Meu4zimTJRJPHboxW8vvzijIxhUMBagyqhVAl8BRUtVFbyDDfmetPcCxr6kuySVCxC
Em1l6ua2mix2JTIhoQ27tIhG5x/8H6f1+qt7KMzRWX92DwciZ5Czq0OcfDuOP9wcqTmzyOj9dw/T
ZsS1xXgpPaLsz7WOlz0znM9kYmJILe5n9YwxBhxSlLfDRYsyAtKaMuTZLY0pUWpLI3YmKBIJGKoK
fr3RyCCTGxAEd/gJWM/R4mmLBDLw0gwqjn3eT1eG3WkfR5vU0IseXsbou3/DmFZxRNTrn3xEMQ4a
ncqO1Vp5cNCquE3aU8xGgIt862nd7cIT+YX+grxUk/eTPzER9xqiHRZXhY7JgBApLO8/0nFJtLr+
j5KTYZTAZU6Ki2ZWj3k6xVTK7Ivjfthn/O2wqNQVoXduWu0T9FPL79sBTr7Qby6sk31rMln30HYD
PnRQQNakaeY2DDgjewCjM0q0J14nvMZF0fxKqy7D+hA5jA1EZxr6tSdDMHzwap4yiIYJ0spu1TB7
KeIy6O6JDneY3SGX9CQ7j+i1gklP8yTQEbVzyDeVkFWDXQdv3YAneQubGIjo7foOLFKZFGf7Gpkb
yvwbUsqlq2U1tAaFsnpXIDR0+SBcP7nXWBGA/DxvWNY5DBKEGVJT0I4wZ7spqqLXZVnb4Th5ai6q
CqQC+AB+XQs8oHN7wGuTpBL19oeMrbOLHt6n5eVyL79FgXKdSc8uHBWknk5S1BKOWQINCBT1ztL9
PppF7HKRRxqYhnpjzFDM5+vxZAEOThrye9rv1/MIpKPWsLRa0q6vXIwOqWBjMdMk0abXrLsUyALD
3Vmw/nCywqIWnQK1/nrLDgd2nl+eCKaZWE3BbV2lBtbE1/WwTkKHuCy2+itzwLW0cVdHMDrdLuTV
8OqxwbQgqiNpqRncY8h+N3GmtW6ej7nl3Yh6rvuDC+N8JiUcFw/2zjSHn8hwRm2RWJ6aIm6gun6n
f1bO46aMb74RLibFE91QEQDlx5BBUBGPW1ZOVZSPijqeq9dTSMe+3DW/0h1Evfz7oSPWWOasPKXC
taKetaT3WFzfpkubpeZ06qxkO/vOpezO36MYPS+lkHr2iEDf+e92UCX6KTVu7mdl+4vytB98cYVw
noDNfJIsPYtNNqksjleL4Xbybkmq3/w+szN5eZYQab/xcar8rymVOef4Ev//3YgaKT+07rTA/OEn
gCDKJnUp0vAkNSAv4/gvB2eiv9RFgqRx1IcBimdntmDpDTD6lLvFazmIzHMsZzMYr++kIJybwxw/
D1zJWdeYBzSL1iX8p1lzb0F/1EZE3ZR4uzzm9bk5RQGNTw9vEJj9Vt4AT9uB92yISiHJnuI+GS1n
JEH7mdCe0FfVUE8VQC4ybqTCqmvxHuXRGcmPgiuCU4vGbU6ZiAfNkyNq0bmiYBXsT2vn8oTucT7+
mH3nJVM+PJMZAOoYRWnktLGpdITshQC+1vjgm8SeDJcjWR/sDLFbou1H+3uszYhCXutirLykZtcp
1xeb0WjPYFZBVpzEyGVzvJSgTloOra4M155z/4I4UkDd2y1gs/tpcmW8KenT1Yj91CLpYFD2MK5M
edsYqlw+vKUfe6W1Oad1KrRWUdYB8A1trmoxfztRCMlnzQgCC6MPmPkzUuSMlZRVsDaIONzBkTy6
WmpZn1+THDeTK4+em8FOCxB8BhlLWlkPDaq7o0zJWqlaiH8dWZB/mZUhWEuIkZcsiGcykIZoRge4
fYIB9K8Qsx/vx7vy0ca7c+4Yotw9eEMeFFDvaSGBDmZ0vop53L/sp9jeGU3L5t/EBrUV1Ge49Q3n
qy4wIr3WU21oUxWFgPDuy0bRnbFpOC/zQUtCMtUv5dBbv+7u0ORVSCLtSID7LoRxo8sWP59jQtl1
X7m1OWEPKytuVRmaVg/0lZvafeZRq9wCuCTt3XUN+Q7ZdhRETnPu0KcQYGxZnTILKvjLSqNwO2GT
yuxsdcsLXzocr5EIh0MgTRaOr/jBUzF3dYZySofSpwggz4w7Fg0DDuyImadagNv/gzLmLUWMBXfv
xQE7CEfCI1LxaTiZpmkTCLHGjo7QQuaxzFIZcPoMIrgJ+oLWvBt+UIyhIGgrBzvGZCyNaYo7DsPK
pyT4esI70w9HLHFdAdwqU1pCiZXZmYCG0YKoQDt7oHe7wpv4EVlIKkp6v1EWgsT6hZm8IG90EVTh
QO/XBn5e2iZXJr/msMlrj0BI6wy7uCPBB/4z/rOrFOs+dPnGJVVojkhQjjSxhhWzOEXSCiU/URxQ
rTcI+GJTsbZlI1fR8U7dqzOglCvdRFHgEi/Q1fbK2eMJSArLCAt5+2pfhOjYvz84lMgtmi7eSTBT
lEcEFpJPdMx0Kz8mzMdt3W4nrxUfzOYSkhYP1V/KH++D84vYL40LuN0NaqH8qvaZg1YQQMGFpBHy
CL6eWlk9Zg91sq3RxCHjPIBUQCbox3dIsyJhcw14xqBBISzmPafUkukuIIlRJ0VSzd1uAyJVcHd6
If1n1LDvcvONnPowMdS9n2pHYt5Ay4AhcPK9eDHRefVI2bR01Nw6Cf4JrDHKeYg3SRERloj5s4Ae
cMPjQgxnSAh1pShyNEbrdo0ytvn/nsOjh/o1ZyHW9yzY9w1+bLkyS6+Pw1f+9BkWdy7Jm0r6iKbg
TtTg95Or8FHcQ5x9mO0PbGNmCN0gjlNtjXSUq73/JSiEP9AGOV2xfBSWUmgXs6qXe630pDH5pLNq
GfTqEN9yXA//MpI/ON9tpCLC3VeYaKPjkBMzRGcl53sKCF1r/HGtZ/NPFdt3Cki+jTcFmgdjYIf0
Pg9k9oWutJm73o1N4qI0IDisXrJP56bKLdwdOfYkKx/gA8fvADdVtRQSvniGv8YkCg8XNnV45+gI
vMYA0IvmN2CjEWxJwPlHaLwBqVocOT7aWAJEMd0VPvn1qILfY8sn4GJdqc84ZO7EvVr6dpVQkX4/
LPIMfJhe//UfbsgS4SY+17MBMsxqmwBAF44XkyKvvj39DOka+U260TLdxR4VLhD8mwMYHwMml/KW
fDiH2DRmeaf4Vyqu7G/NNmgDNqesESXqYjvxm86gVOWdoxX0kW0HYURcSzqz+9+Fe38lzWCd5XKv
eZ+eIxmCaB4WPekQGAW/jBLyrixKEZmx2/PB0/XL+H2BDj1RhPtwITYeoPXrFeo/52JEdUTVt+SD
PSZair0L96jkdn2zC73mr+o+Pr0zX9qg8eLqFT+q/KjKnSxUI94AqeQ6LHV/7SH22U7pfdH8gZXw
qVCBQ7MGYbVhZDF3Se3l+vWsbx9qbF+tGXZGscteXN8KBS6D+nSERcgZjDSS65jHdIsrG3fzOT/S
kz4h6SGV/fBAeQfr8Wf3yXQSv7R3AMr1MlW4R+JUfr0w37bCtTVyHZz9lrzzfxONzY2xYcIk6X0O
UXAyvPPaUautF4cI7iw1wMGGQAQXdZvlWFGRLAD9vCBcWxYxSqbTGO7b49vigy60eLGYWLFNZ+Er
QKu0BG17b0r/5X9b7J4D+aBzW01awWlaXrcU4Yx7FZoterZoA7Vg1yi39JNr5B4/UWFzt5SRRHNR
a08MMoATfjrDri3OTbDcUzSK4+VVMBl5olK5PZn5J1Whc+fOq94lL4c1h+cKnzvej0wxIHRIOPna
D0BJGVLuZjTw/U8aEbYUsSQV1y2w6N0ILCdDQWJj0Nv9wQvg8aYjfumJRHbwA6hyaSmaFp9MBzxV
6ao9tW+d5ZoRnQNdIWgBXjXluaI9Mg763PV3F6gYRl8IlX8GPMnw+9S48wILw5EQzt7/Bagrjdv5
l/zRu61xpIdWlGHVU1Qg5ak6j+L0DAn4skITgXB2jYsdQZNZULMT0hSqM85uwVDRWrT3dZe4Pt1o
uLsL3J/IlNghoLrVpcUbqZthCTm+++82Wj6lP+uyrh7tVOKGlf8Gal+jNvwXWCSXjBnIxStWVEVn
FyTo5NCN77AWCLc2hrMD0JeOh6erjeb+f9q+QskMQzWt7ScT44o3x56k12ojIMjRQ7+YnDEojWj+
PygZfbZ8erHhwCH5Y/boKzFw+1s6SkGXy6e94cxPfMFfDRa3rvRB36l+Vf7O5cv5URKDXRn8nlpq
EALXOv5ik/BzXU+VgUlJM7kAi4E79PyFlYAyNNh5zt2lMOsIiGMGOjowHfyu9mK4K8ReiuCb4eRc
X+FPqjww3wDCpq8puPK2q1mdqLXicHVMCu5LmXeyowOQWAbvqxC/Tv1pkZlmBlEvP9UK4xzT2CTa
lQwtHtcIsoG2OZMDeyBgbBJDks+65eFtmvDJf12Lo3ikdzpSiT9JXQVKJBFHYUBsuPGjhCNPvV8J
p6pwDXrruZy1SkKi/4dk5qb6nlUMPYnL9btTnk+33Voq3+ODJXA86oLk5omnxALzNiVbk3EE7IW3
TBxe6mYxme9f+sjJsW2HITxpljm6yZDJxMd+hTkvBUjKaYPxmgOIbTQaqCl7SQngLPg2d/tipIHa
15xDy5hOqW7x1/+N2141v4pODN6mD0Z+UFoRrHfrOIxfTb5svhe4zvmqDYTaCyQ3SVZoIC1760cP
V7V/9WwSixC8YPjsGMTCzlyV2fR5UzUwp5FQiCY9v2KViu2otAPum2Aydm4AP86UWZ5miJWyzp7z
16arRFo+bnDZ0X1XqWJ6/SaGmBHVE5Y+sW2M141z5z2lor/HrphyoZQHI3qJwWwL4cJc6Tm4BcDx
SV5WHcZP85TqOYO2L3obxuj0XIO3iKHi94SjiWuh5UAxnkxPVsWEsXvnFywnKRPD9gljU3PnFqGX
C5P60/6iCxEtEIIdwA+wxQkXqRvXcxXdb5NQyBPtXz06/i8T6bSupRc2hwUEADwcs8CTxU3pASM+
zQ5A3mo/2nT/SyaiNnsaVPvTiqkXZA4FsMD2ur02Elu+lbQFEoldQzH4KdnAZwSZqbmsIXP0Rarn
0QYePbQw+AHRc1LFpADiRQpFzgC13MBczNRSI7gjBF4OdsoUzsYNZxUejJDzV6FJCFbphSy4lYCB
ejP7hbmN7lwKEcTG8YVGWAXibgVGjBx0pPZiqkxHWKxPgCeaQOqxYdFU1RdC0dTRv+U/9bDG78Hi
4kLL5suF48r7+jSiGJE5WgYMawJltei0IJlPfkbAFCUfI0DQDrJvgmz3rwkW8sFRRW+holpaE0Wz
M82zVj/+SyhKrwojR7Z5p6QKO5bJ67TvCVbDbF+EoYJUL2OYmc66i0hYiEvEQMV1mbwnAFJYlCR+
7s5r6fRVxxTnq0uhFparTh7MseAQy+rjYQgJukJMcvvSV5JcOl2fTMZCn0+uXWrQHXt29S8dPmXV
BcADzJjScZ6INE27jZBD+io2SPPzY2K1BLNhJj0C0A88pWtusvwZLLsMlCvGTk7uvmKO1u3itd5n
yid7g1F5cey5T+bSYvxnflHG+ArnAONJ9ZShlvdigXTrhQld8YfKC4OiZKozmifz5bUKvFwfz32y
4c5FRGpj3SFQ/OJgQA8IN8E1HFekwN+jw6ktantbRXeM8jf3KeUwUvEL1LZYFhPunl0CfDVmcdlF
IeMSZHOEvK2GfbCi8zPpcO+MhestT5VWmeQdHXAOBOUqHgvp8zGqJLWX0bBiLg4olj8guoDr/0Qy
lN/r0CiNBhWQnCm4601u1lvvN9jE/WEYaYfRwQl6EVHBA7kPivpMGpmNquhGSqWU5kloIjRgTm9C
EXnRw+IGm2CQ2hpqQzQJovSdUEZof2SY4ZTU2v6ooLogZxU6kkSMLDRiguDkSHiswrCn+kSxUMKO
pG/Zhxz26z3eNTGWN0PpKBNksQihduWrXQPMYBxWuJ4L67pDWmlbymBmCiB7Lg65kx49PbMmBwfG
pvawUPgbnacdDRmj3pK3O/UuBG8ejhz0xfOLDTSybJ2vkGnKoVn5YIbjdcJVmuE1Fgh6jabO3U83
uuWoauKemYgEX72SgnL+6x6miscgBGM37AHZTN1KixI22gR1S3FMVTXRKJLa3PNs1uqPuQTsOuCE
bvpcXofgZBRcpYvuLlEfvFDzXTKeF3oeGBJjVzLKgBsAUbMY/9wNNKQnmg+QEKBbI54SD2zAScGE
mj0B6tPI4htzoJrIKpx5eQZPQ82fm2uQhVynkWlaS8I7ViqVh5hjId2062ezhsjdeoc2mbt+0dLa
0jdrRYKRNs9eCc/O9/6uORbRaqp2/vLLlXzD1p6nXnXo+jJiFdERlmswwFN0kr2nFfoeLgkLsZT/
8FySX8ss2EURNbsfhI+eeRbZUWxiNteTxcZBmQAd3duX6FS9d8QGQfuoF94x1YKSNfzu4RXzfTEY
Bvvev2s2Izc8TYPNvjQ/c5fRcicsXy6vzmwNhi21IDQxfo9d19KaWYQ1h5/7nFR+ajtcxjcHUh4h
6aXn+U/BvsuPcmL4gOmkxYQ3InRve+NBXunnijmB1syuZ39zC4jcQ25a6pPr58Yz7t680RrAnAQS
syQzTcVS1ex+caeEjORQb/ZoUFGbol3MNlbVBYLVKsVNthS3qobPCtu6VMSfAFd049CzTxupkkkd
w1ffmr9b36fq/zorn9DwUHv8hhLfyj6RZXA34tsR/OT0Fbq+NA5LH7LFq20pJcBhrEZgNK/OVHKe
kK8r8Pria8W05MrW2yxeSeN7xiPzlqVfHSa0bgILBtTXS+pz3fKCDKe/DHvLKwARrgz0lCQ9dwLZ
4+dTK1XX1gD0C2eIpwl7kxuL8IbGVf8KeXzYNY4zGYfTMG7n/ijvtMf4ATskmntBtfAerTxXAHQ7
mqiD+ZcY1XwyXcF3gXDPM+aDpwM5rvOBxfOX2ESstX6tYBluTZkGWhmbuBSfVWEFVhZnOAa8sNuv
hRnG5ObV/Hbd6Wb1uz/6uGXerAh+iOzi6wh5pLFANdrB2uoH0vUtUqWYmXO4/NQM04JPQSL3un+h
Yn70mfUOZHIilKco+4/JC2SfYe7pmuyVTKCB44kEBY0NS7hEMaq56MrPzzy9diLwcQuN/5VTTRkB
yCZYu84j8l4yRpD2hYlZukBvNapmH54iidC5w/E72M/egXu+2GCqCfWu8ApuUrcaS6pEgkHWn5/d
Y4YNrgwvqovXfUxcByoiWwoireMFA9fEWkDCp8g9+zvVlAG+SZlVylWQ7rUpSI7c292R+6u2meUP
FAIzLxPeZgbGSNbMmb0YWoZjCavYJJoejKi9jSS2+bqulq+1Oj6VsyGiEQGrGpHv83erFequttiK
Sd9du9UBChbkPFVSZyIxyEiZ6tvmc9hh9V4HDVT6PqNlndD73GHgJQPe+D5M2NsvISRIY+9n/0ZK
14v2i0cXTcjifNMlBpzlkYyXMf7/2fjoXw3onN2szNSrQQwbgbt6A3A4LqXZBB3Wg2deN1c+OkRd
zDaUuRmPR7BEVAOFEPsFEocbAwKdIx6QZyb32Uu6yp4bd3VR1n3hfnh+W/x4P/SajCkZUL7OYsbG
njaBse6CNPSGbnfo4TupJM/D+rohL+OWHnFaQP0F/KWonP9N0mt4SBz+z/7AQhKiCBrCONj05sCc
swJGF1VNjD4Bo5Yb7Z3Pf/1pLwQExv44QvyLZxuoDPXJaIBydLSVN3hMlSQZniucRmhl68YdL1nt
Ewo93LEQLRxv1++vok865Xd4euAkKOEEdV9bDVIiMnEKpaAQvFEyn/sWwAPqLV1bfmwYkeizVfom
c8yQz8blQC+9vmrko8+w7bWtz82OLIilyLvK3TuOUqlev1uF8qWgQuJlfcUZeqdagGitRfd+auzk
MwWmgyA3XbbCz7WXE3yoGQqlf5uEPkIKutFRtJhNCrJD0qFXxQEEdEQZhq/h6izFjMMPnp0r/BJx
qDX6YdfkOe34asuvIe0takmABcYY85i6Bx1l7aN28NcrjRAYGWUmrH4IMcgL3qHD1XzPATiigUFi
wQBhv4uzSvebch392ErTgGKEOBE5RP0D3tRTyLrnK6qnTT60cSB1WIG7ZqFuYzzFMWAlU8vQq17D
OpmeaeYkVvWq2oseL7X9XJ+UbJLpEFpSQ2y0p5/i3UrLOEDklUcEPfQS1xFRvJ3Eba2yYonXdDhU
IpYdV/NIa98ZJD6XN0pvdganJCZC1bNesfx7NaeQ+nP93o4VTHb6MxSj8pagiXix4/VcBBc6CchI
hgQYbGoejcJHfgORr/y8UW7/fbsWmjUkCint8hk/4PNowWvJzKOM1V6EexB6AdSeBFxK3KAiuP/L
8imxCb65VgBrUAMID/SIIC8WbY72kvGQDiRLNzSkFCQk42/EKZ3eptrSIZgpux01XQG0Jcs3V6Gi
H/5dRj3RZaPiZ6IJojELR5SbRFi8JM1f80WlpcB4C0/A86Qj5PNKPTSBCmn3AMZqLl2N6fWNrnQl
U3zf9nNRgkBDP16PZ/EvGjyryl6F+ncJg9q8EEMy/RhIbHPVT5lDnPZNRGvcxwruEU5lbFbgSrM9
JU/VTKWSh9W9ySNcfnRkp+mqIqTCCSEvbo79aCWXigCo+RaIU1mJR8HYLSzsoJPq3gQEIYqCcM26
yxX0g74XLYNWfMX0ZyaSsXHLLeiJTvvmZYXQL9I8bbuvmJeLTmcH99mlY97GVWKO2FEdD7weswZz
8LbBx5nNAykQfB2x1scvcPVU2zvoA2FWpeFTTU4DU+Ns9XnoMta5o7mOojQ1JbIPPOeFdIBZj8mj
/OFINveeB1+JtdvPdkiJa6l6kkGvoNkm5XZiTloz9WLeRto88PnqOsPjTDX0tjwuEofOtIhT2WiR
DVwlVwQCHVmR5lKbGJV0YPeLaj8QJFD0gWR61Ns28JCd/wWDrnI8H9gvtggwa37sc1Nr+rRjZb5I
IBc4PmzZcp8FWGqxjTmnBWOxPyDvbzCmdb5XTyEPW385cBKTmLlzcYGB7RkoZYkbqZYy70dqis4j
UX93EptWSxYLYnuZxFjIM2QBUqUBVox7njYEIleGFvGw/BTUlh4EmwiTdKGWlPhpFmcWp3fKmB0t
OXi7GOTBxpYSY7iPrKad/PR0ApFlTvfZ/B5XA1gLGlNXiiLGJhFCIs2lKponyb1rrAYIMUf1rjHD
DnubuHVSdlE23QtFxW8p0F4mA1h7MPNBGMejXtIBrqBV7t+OlbNpwjUmxUt6ZK1BwHMja4wrcY9V
2DUbqz5+WxOtnAjmMF1otZcK3QpznnMeaDOixJaNUT5DptcOEfJVUK9g8SfK4i5d+ZOTZFHblOG2
qw5WAM95p3YZ4/JmTPFqqf2hwlA3WtWAfrqp6lo9/vDwKy75alL9Tmu6z3f8vf/JLmQSS4T1VknP
HWEKoJe9xbk89fkA/ZCED9LTsIr7Fg4ecaP0SWI7IiBA+gz6FysH8qn3vkolUhlLOULgyaas3eZJ
o94dyb3RRsoYs9l1c3O3ASxqqkm4amPDPDuXfD9w9Ub21svbWuvevTLKhICF4iB8gwAOFpZrxzo6
NoRhCGFlkZotjaNKkeEGAJbGYKtzvByX7RTZ9VAwq/4cNGqhEyHOFcwJTSVe+xGmeQysrJlO/hYs
D0g/+HlP3se9seu1Ydz5RYAk4Rvf5oQmBrE4dAGDe7E3v60IpX9OLUp0eH6Tek3RAf0cnrEJ/pvL
GzePMEgkXb3SX9y6Yk5Wy8yJk505i85eLYLERHJbut8QB0SIsRry2DT19wVy59Xtqt1r32ryHs5t
jZG9f0nTXac3W0nKFkAFYnyCZw1GxP+qdk9pJVdY0k3Pj51GP9DZ3Fz9lUyCvb4Kungrap2lRBbr
JUzwX4rTpYy9bfFQdlZKJTzpiFHl9JLP4wCBi9jZE6HdEydU5fWFqYCYZ/xc9/Ct5XNUjmntXj9X
vJnsHcToXA2H2/7+bHcqo4Y03xsGNpUVRLerzm66E9UfHavEA1doksG+uiyoDzK5TbLN5fkA7r8T
eCMILAUgbiZV5B93d9Bj0lnWRW8lFpt6VfDV2NfRpRBwgQAixOajNz8cL7Mb5W0o4bI62EO4wDA3
oU1JdBksxI6EL0rZCQ0Ax/y+1frm8jWhhPs8TViyZIJk+NYWMsSrlCdmLRnWDLqoHhBjirbH2Wrc
PJrU6XFgF/R6oMpZ/3OItv74RWd2kyL6CSgVC9Zq8hRTPcFHnEd9ccev7OvgGfZ0Cz9c4jhLwnMe
L7hi01I7qkkjxko/aZZcnvaKO5sNTpgji4mchuG8Wgh4RgTZVlyFZi/4lpV729/Yz0FIMnIm2ehE
IOlhh+0zPwQ58p44HdJ4iv/ukomu+/hl3HfeezpM2Nosp6W3pdhb+iioJEpvnnmtMgSoeHRF/YoF
BpZPYQh6Ep9w7hmjRAlPfc3dEuvQjYRiaHjdmb+4I3kj3w73KOQraCWPjmM8D8UxrNvO8KehlGsm
vYuc3/R6JIHdaaTYb2y90bAYcVpWjPf1JIzhrb6MsOCc24r7LpzGrEWjpU6o9AerTN1tkQC91wXi
wpseqlM37dhOjEtWYyL1Wem/WecrFKLNUz6kMAHSfBjkGpm7n3IaKZdu3xtKNm8TB9LPZUH9D2F7
6YYZ48dhSOzkj6Ts/uJA+1UREqadK+QVuM1iaLrPvl/au4IXTi9z8N9T6+SVXFKD9wLzHWl9HSUV
/ZoXY18NTvieq1X5BSmbCZf1FmA3Gee6nkFaCLcJefEMTQm/h1+5CTDHdTZihSkJXBuFZs6OBQi/
tBbhDMpvP3LNFa3EGx9dwIaIzRDo0HQBU8nAQXEMCHxo4RQsZ4REhStinHyOIj9wb9ZC/SOOO8mr
LIc3bKhTXu1oR0I1xkSlQRYGz9/u/z4qgIsQYbrUSSbLankmQwgoozntEM1xgMKzs1gYPTjAJsKx
JavmuVDbV//piL4wwemQbMLkGowE/mM4cToAtCtnxopD191cEss7LnAbOqnuhGIBsQxExBE8bQdt
SM61SOl45jYCeN78JC0e3/3UhxRzzIE6mmxiGqgisAj0Wb2oWge3JTHxiRW6vIw1djoGNB9dbjLm
OVjyk2toBe7QcBNqY0FSn9jNRH3pdn3An2wBcEJizkF4dw5x412vDimivAC2VLD6T3mB7w34Jjhb
gpaWOOlB+Rtpd4+MX/GH66EVQcKJydb8R5lcgoaE0w8TFE0HuO7M8NImFk1spBNMF/hXke3rgma6
pQHIv2z5RTjxAXwTgRtALN3Pk/sEfxF1nXOvSxKrgX7/sRQVqJxJ+6KlDwKu7mxvzsCTxjZdoBvU
rTeGB1Xee8hQvBbyhfE4uvOOvfxg2sgbj4fu73s1LhSmOkbkNiqoYSX0zvkYad7afg3tSjPDk3Cn
yvLKiCLbEM46b7ZlZW0EP0O/r/LejH4Ay2sLuU17aFwLOP4tOuj0HwJbgkcEkxCDkN3/oEmE7BT2
31nH7xZjPIS58bkjVdncDshKJMVQxdMI6jr+aGfwW0M7zglGq1xcTTkOYCk4Y9AJrY7+5lBAHsyZ
elCLMaHrYg2Cw0udh2S+cKuttOdzJ9A1vjPvbcbHUNLrARa0HIjvnyXL3fpRfElCnnr5SiKLHzMd
6+irhUEWYdbhbroPsAr0WJrjZMks0dqg+99woKhoPfhR3yi5QIjnl404EC2MHT9B+51Kon0GOl/P
5p81cs5nrFiscxWFJfpXqLcW6wNSM8rEO4GOGheuF+WovAIOWHdbaGqDXecoDOpKOADtxQr9mVmn
F4Ne4f+xrrGxo/ngosVAk5Ps8iiXIWaRoEGaT77F1hUYmACrF/mCA23ky+U7+0Zt9dxbEdcyfH7S
2Wo80PoU+0sQufXQFtsyqFWSt5IF+rLeLib+CnrZqoXx86MJkLZMuPwxHIYylA89Hr9bgAolMT//
LbWe32ScC+hi7M78fHuKQV9MAA04u01kkbIPvud8rrckCx6dhp2VYiC3igtjKOG47JK/4HLE77ss
RHoRMKK/qAOOklnc8MdiFTp3wVZ6INmAKrREL+5IM0rJ2mI4Ml0PZ0Q9dwizoPmRDFF/amIhpeld
NmlR87p+rVluQyvR6iHgb8cll5eF0Z19CYafmqqJErHV8obmrEqL+Je9XjIGQgD22tpWyc+7+CfT
9i2NPu5Pwt3HDR9XD4RSrnV5KbBakSwfI6jRVy4aXjFzcRj1HXSZe8QMDAWDZa0rVn+/4eJjp6kb
L2m6J3SboprnSQOJan/rMjweIxfEOgeOJJoW6HifCmkIGPuP8yJZkSSmswfYfLviqUYxeg4VBPWJ
adjUFsZirRWgf2gKx2C0IS31xx9OsBn/eoTUKmyrpOYBTaI2JTbgkMNLWj0SGCI8fja4M1+MSZ2x
Y6ejBYtabiEGgTC5YmAdvvOuXvGCtF5M3NHFrxTZMWkpI4v6kOKJRBSR99t2uh1AL2Fn1tKBhGYl
IlLTXzsB0xdzH5qLkdZat8brCxyzppmLhZKHNVsN4fI9rztMNlyfIhUwl5sIAzLzPJwmu3fCiLlI
mwa8eJk4hOPoeRu8cC7je13k+cLLKmfIcr/ytp8Za63ffBaSLuazqQDm7ofcWjExCxJPgvzA7QG7
vJMgxFmM//DNxxyp12KUBwLF7QnE+RtLICcYMYIG/y6C4A6Vj53ftGGXuDP4qlELMFbdKiW0wXZ6
GnCzrfwP+cdZDvMW1Mdgvl0zWaVoPSAmOh0nAh0lL8QZcKF5G0FkPNq1nhJxAYe/hH2CY8z+zPHm
lOu7D3FgvJy9xG021lywUpAsSd0HhXdqmu77jmSTYvsfeeUKW4o7bGnLaN0gatQ400/g8ykMWMta
ulLbdbE1EijvCw6++3QNqd4tMfc05hew1+nu6inY4MPemfuemurCrVakYJofhFlKEE8fS/E+LKMy
MeKBGlPSdu1oBg4fB5+6Vtu/2bLJzjoBuv5/SIg02PcqEkUizeJNiaL9dmF9QQ9vjYS5f6WN3T9p
Eczb26C9Fv7FtR8MbBQ7+TwY9yK4BSqSWMdqL0xSmaCjvSzoJeEMoSmBYuaTtr15/V7pt4Mx9I3N
mHwqBgg5NJ3Yd3fWedTPMrlr8EKHVX3QofB8xHAPpImB3FbcEVG3QZpqpUxniDKMiQBJHMPnfKQz
id0T5XDzrm6/1/SKJ9A/APkeWBVS6SHOm9REE7xzY169eib9hbCfIX/+7q9BdliSz5iDd9Xjyqlw
punuwqAqIOq4twE/Ums6KiGKLVXVa4LZwW/dp/mC8ovm6kcNsbbQhQwTrVpqDiCfQNZt9D4k1CF2
4m6r1pszVFTTKxTVhVbEoYA1C83x3xqnVnb9rvF1krBYwF3078Rxo1rLNkDtIDU1tC3bWiIRWtG3
TryEnx4NuUmhjVwuN9bL1kW0JE9bTYHOxtLVVAuvfZdJYljzJ8cb4aOeWgubwnLiYXleIkPApKXG
i/15RodLRG+J4jhNHS4V6F1Vxiu4GW405OvY79TQXqTBojL4dBxqqgFfbOicEBR8wmXMcNLfxISI
TwNqSzxQmgNaP7G6ce7/m+xidGB9uUb6nyyAZIFvdLWUCeEXlmCmNpBrhlaNiuzJy6Bow4xLIxOn
JSOcTZTyrcB+HvpG3Rv0m7iQfJgVipBpNNT1y8kw+brnJoVY+lacJti0wmHT3NeSPZW37JxNfK2K
CHHq/KPewOMSfmz3fKF1aWnsWvjFqfVPmtZEtB9cj7azzXG5EWKyOEce6EvMvxIMMKuiIii4yvfF
fWc5FQBq/bjFgzijahqtnzqtCAQt2jkSEjkrZyR0S+Ans3PxfGrxgVkOdp+4ktWKTkXR3Mb0u/oV
5r38ln6VdZoY+TBshhBVdgLvWJzoZxcjkebPucungNDHicVd8BHuwQi8UstxzDTqr1welxcXUxSf
VIfFi3V3krEpsYkOPWrlXG5whzMo3ZRFLAEnRyhQLeQTGa1UCapnq4pj2tygy1JCubsPS4JgAV46
8eeMFpQtVUG+NDWj4ajRVJhMugcyUJQgP1iujZp2qsO7egBiD7Vpphr6t6lGKkzojzyyzPXyH2Zg
lZ4GNeD3Zpr28DBpjgaSNiMYNIlwWolObizyX2QZoahRq80lKTCeZWy9aBADPRb7tB6U5buoGYTX
yYPdwW/S3Sr6jcUM6EhX4OR2X5AZOIicCzrNAq+p84mVUGFsBZ1pJe3Tp+NrOmQ2/caVSaMIyuEW
zMbBsz0mIzjiIb1mZi1GAoW3rWz5JjZ8eVUjZ/mpEd+im/VPS2k1GMJutSjmwQow5B4TO+pcbgXL
X+cO4035TdnzzjUxsnuemRSHTy9AO+euxvnJ/HcOq8bTuyTJWKQxa4sN18C5RL+Xk3O4KcArDLW5
kWS5TBawLPE8Yq5voRTGL9jY8JC/4SQyu6tX1A6KjzhM8/+j53iXen4FV2NeEzIlj+icfcwuKfD+
mvneqDDICA6uzuayQsfmtMTWwkuIA8QSSDKW0U9VN6BCps0yapuEfgtbmIbYl8A6QQ2kEEbvZ2xN
RV4mfSNCzF4UFSh9TbcTVH+Ns/oM5RubosUTQxJCceNaD9Hq4qpUG8zdAcXaVh3zVh8Dt74KVMDG
cxABfzMcmr4o4W9ii4BIY5GZajVtLaZ6A7PCBarLSWMXXIkwsURU/q6+DYq0WOEL1L+tl8tj0IM5
M7I9gG2iZOfmEacHAlDsJmxbtUYv1guvZb6zzqBnhpI1Bk7izqTNS4VFc6msR/zUdl1wqvVWHzS7
28T6w3EYeL/ELUMq+qo2VaViF9yXaGqiN6x7L5FjBsV4AHwaJNrbXm6iPpMt3mEq3NR7BHYqc5I9
VXStWbEXcWned0FS7mXVTcqjBq1zdmHHaU/lsjUID/WNeRUXUHA9qA8IpHAvFNqnuEuWkmOIlFU7
FXHLMEFgu9GY7f2Syb9PgK8QiriNjvoto8cXPsMbDmueDAjFIIsvZvQGPC4mXGwZ4jD3pmcKy3GU
nFc5PzMRpBJOmdOcAWeVefQPQCx8kUFHjhAHYnydHvy9Ve7BYwbxEhj7uWvdSaXHZDX3DGic2veg
OE3ZxUJ07Y70bcpo7gnhvW+ExVQn/MMBgD9ICxChXvYO2C4zX+4xSVEuDxmKQvwwQrfrj2kSkcfp
KuOgsDPeJSdgEZHMCaKA3T1qkHKDJjAIlchRPk102zcPimrYL8BxuRmdNbVL77BYN/v6hLpiJzC2
cwoaKyUV7lCyJiS4dzhM7DILWTRCYu6IweLvDhMfgeUUywjffLaW2XVvtRPyF71/YaRfC5nMk1x3
zLsJgR4UHNkk/ii6hrm5SwOw7FFvIv93bHg5XiXFBFRk6+/bAhNlNlDTToi/P7oaqnGFN6XUElqM
YGdr91QSOv+5056EGIdfDo+zoZ9/L4gmRSkcCMcLb9Ny6xkkwXHKxrrsNY5fuXT+D6QyIY744jUZ
hNG8Xb0Th91AXlgfDzMiTZKGHCQyw32gtT2Sb1Fv6nVqtSrpqFpXrEzASOKWQKTnkk+tyGbMRNkc
Y68e+G/vTlCb5Z3UbQWZLSxfaZqj0EdKZsv1pvFYbb6OiY1dlwncXLjn7EYNDD+3I38z74QmyDyt
LTDpzLUIExabD1NzSU/NA7AsCQ2G0fjXijxogKBeys5DvBU1Zle0OmRJy31i6pl9+hs+G3r6C/sN
OkkxChKUUyK4iKIkCVtUx96kWFN+4nZMopOBporXbydInoSV+8aCcxWk4z27pdFVXG7lv9CQ8ThS
LfpE8bVdbuePEQxtbYe5P8NTLyf1NtzCkcLtXWOLgt2PEo61bxwHcVytJE08vCvJAoH7yXBO7PEO
MqMjRk8c2xewWchLR7z8YYr5q5qZ5AEM14OUGSbKDK+Z2L44wDmL4Gx8Tdwzcram2lpqzuA06ORI
CGWhEkJUZkzmlqfj47bPfceE7paEN207KGkf/A0NO3p0ocDxxjQioGVYbFVEZ8LrnSdbaaQMWTXH
+nkogCRwzQVKKb52cJpas3kjBkuAZ4QCmUMmgrrzcp6Rw6O/aS3lD8LGw9J044JHoQM3WxuNAeze
zv3csVHdoUVqXsshfsQas3jRgt385ysKX0j6reGRr4VPOu0YTT9wgfbtxCfhYGnp9OvhBMBekPzN
QZykjErShy0PnkOiqExuDDSo1iiNY2TVr/65pJApUVGskoJQ5dp2qthzOAQTVlhRgLkwDUnRP4sj
0J4vaV2jmPbn7otk0mfWHGNH/n3O4bx93uTXeG7Ns49iFAaWMpLdEhjKD1zsy8822o1FTyzVN2EH
O4pxVATqr9kNpo2L1DqewW/nNNKkum2riG4HEbsY5FdSg1IAzn5DHfImlOVDj9WqpDSbc+h1Q2pO
Tlgt/Cztr9KKunXAJoNRrWBMmE32wEwIOPASfR2DoUS6Qsph94lF2sWq4HYCFh8HvhYT+BLqHEhD
6/G+l9xBpidML/M1CjXHJk3/8PlTvN1HcJLFs6eSNye8BtFGW76wY+TUDkHEb/FOqJYbG1nFR5ty
T5+v75M6Wx7cGMsenKPlfu7EYN46eKBr4VSvxUkBqhwzCqCMfa595e+HaZNk0pbRUJdSp7lgfkcQ
s7aUA5eLWoxkpI4AMRG0rnT/gqow6EMChlZAmx9AeAQZKeRpEFW8fEL2SMvJPqy4zVDQbGb/afWt
Mq1pLDvltqrZrTD1u8soqfj7Cr+JsJMp893HsMq88anyNCZKUieX1RREYHyA29UsxPie46sHj8cq
p8XuMrEK8oBn/XjOnMxf7daOYPeKAaRvJh/SYzO+yWHuuVAYbrrAF28XNfKIjAsem3j9SDjTy5WT
JwXickI1bgLYOQjoQ03c6gPxOor7bhGfOgy9GzH1OJbHjhjUxBvRH0CUCTkdA3rw+6jTGZxsRc/U
2nB+BBN5jh08BWwWgSuHVEuAvne75gORAT97uFjOMgAYnOvoCOx6m/00c+J5PZOyJIAjxQXY5H1t
5JpU20mxFTzcOwqXL67KVUUPCYzNL20wL4deNokre+wtoob5fEaYW05PM9LMFb28iWuHjMYFKn4S
+ly62XggwuWLyXfeXNqYARgFWXb0wJ+fU6r2aRoIdYoaAOsVM6PfHIojq20uIRJPioVu4u2+P/Is
hMJpwzwEkacdbjbsTbcDXOEX5kAMq9u3b5428LVGVp5Ys85FcPcjqlkdSo8e/CjxfIQNyhsHxZOw
JWaZ2v/rsum9zEOIA2h4FFGOC3Q/TaKxh4+h18C5GN0TygR9L2uUitNYgz68tNrolKUt9iu1q1K/
0zwd+90nKrhUTSXeLvoeIOySwz4V7mjlMv3nDkVZjZtEvm3MgD9mSdv9zGoIee7cvYNHn+4xHb0c
jh2TozaltzTsnvkYuhNiXZrtr3anMpie+13Gbm4gxXsGRgBsMOLF0FFXH6BOrwVkGgGqertr8amv
1Y2AW6Ew6kbRKLVItOqvpUB45gnNm20mqcxAC0U3Ude52v6/3Ae1tx00oAmbDSPBLx1qw9FOoCzO
d2aXyEx/A3LxI+vY/yLUnTNzb0Nq20c2nqAHY3WJUeL1qQ1x3plgMRD8tZGXauuM6GKRY/VeLHxv
FyMyp/KDDrVfh3ueMbYHkXLZ1DmfjcRRyNixckxcrclIPtVP3cifVK66/8hRXKptSGO34Oslwh38
EqPTVmwM7RjyirpRSKzQezZ0bWNhj53cTY/1yvsEt1IBKqjObVTt2dgLWjzdVB48nTZnYm6G993q
g/xUqHH6ouVYGw0d2Jwh3JCLu59dNgZAuQeagxZYRu5Z2Ll5b08WNoDdZgRlwABI6YZ61sMO9vb2
BWSFuYWkloY9yBwAuMWsiSdfKitAwYkw1Z0KNc3FBZ+J2+D0Nn2YyB8txD72kgqBJFGjwwGULMUw
X/qqGIK/qKtVSwZS4WQC1lDkR6eFOIaFYbJZZGk+5U6dqKh9cfvQqOi8FKPHc9kfXsTiWMGSo1M3
nOjVh4+YpNC2CEeN6N3CEVN+AWFCzvjCuh0Yq3Q/cL/PBJ8yur+7MB/SrFRaRp9yeMnJ2q4r/Vxz
5pufkPEF/JOJdDSUT1Iy01Dz61GSQxtzyOVmoH4xMaLd6lXftJAXgAlrqAMJO4dD3PduqK3TpTAl
ehTYbeuK2q+WNl9jhdkORR2fdOsCDN1gOhygAwiIcJYmEEG4Uo3z1/lLTDWaEsdwk4b8p44oal4j
6akbifFIB3oB03EQRrnI8rwV6yALOML160QJYXwI6rl6scSU8ehNRQxBktaDwnjpLPjeVS3t7E9E
E0hqyIQNJwBxPW0zk0o3wqNFrYEcWcoFCgzBJ5mfEvC0zozvL/GJn6M+XEWpPI1aQP0P2vMo8Ml+
8eGt0LcSqTcubS/VpsXfBPVSwFuMZw6IkqyNvR2rpoGVVpnhpHCSbP+oQqbDor3376x4rA3qANao
F340zRCD3070VvppMv682Q+0DUDMZWpJYNqQO0sI1fVPUOawqZiSMF4Hl6Wp/HfW49dtvwO1ccc7
K728FnZLfMN21RrUPFXOrgxgeOWY7J9wL21bD7prcqGQz7AOcTRqin5xCccf9C8ThvpJNRWMYqJL
c2i9AmCe/1G/40ZPAmvo5f47JFqm9cbjdQtXTEtgtL5GHJMuDJiqorKEiIwQzr/fcVVqaijOCVKn
1nW8cbemQSxIaMefexcrO5FSv3CNbdSv4ZlpgviIVSU5fH8L/Sr6jHap8OzLRXqJCeAwwSCd/E1L
p+kqsLSHgiP9J1dCXb0/xg/roJD7g/q8TK8r/W82xX9mBggldyIf/6xrjzuz1uQaBJsTCL6Ux++u
rSlmx0rJ7lPrezmf7pcAA6Axm4edCZY0k1k5XnB9Z0Uvjbq03GTeley+LNGBBtFvsEazr1NRHpfp
SBwWA+UqwFF/DMs1smolvhAe6YZY1KjlTn3mgFNKeuXQoxVzsNFxaARRW3/QGy5noeOdNKm0mP1k
gmGAHH9u7qGt3i+N14JfsQRqpgMfMFak3pf3dmupo2d15sIPQsOx+gQdgwUQfGpFnEb8iHu5+fLj
yQVcq3QW7qddqMnS9KDTsPZ7bSkfWLHs7P4pGRNK5XjDCAUhL1PvALxCMybQ6078CeipydTfHaVX
Y2YtiQVzVTYBL9bN7c+q140fDFT0T/9i6XZV/XdnniOIKimTm+/MJggJprhqbVepLuM2HtVzHq9z
u8BjzagIh2ea/gptc5XeBIGniO8d66oXY0kGlsRlcYqSD/R/u+4xSAx5xkvBz+zlbGcQwduJFZ9T
PIi2h18covm/V/08HtJXL4CEexPhzcThSvKL07EfIKUXQ7K8ztfgUZnOxgwrtD4bK9X4fxV2+iDy
hzZdMrai9YKBZ/huEMMaQJPQGPrXyHdrsm/6XKzD4YlRVaDPM1ghemY7krlrMvvFw8uyYvNI0ls3
om6R91ogCHN2odavSU4HAuNoXqLbdUARd7BCGk5BcyiN4AQE9XvCvoU9kvgh3bQBimdCrWihAuBM
sLEkN2GC/8CI8VeUqGAUq8RkYvJ/FN7CLKn8kmQ3haRF7P/zDXJK3rWPOqfZMLjNBTQGTmv6ZY9d
a4Mt9ZM+XjgnavyFDtk0eqEwOMNiiqW4Nd9R/T78gVLentsS6+4uwTdAu1IbAGTn8c/JyyIkzVfx
AYl5a4qIh+NEmd/NRgZ/twXlmBOX+PPrWCaqAJo4k5T0IOoas0RMnV/IBhT+tlAQWHHAgWlGfc2O
eGNCVQ7RV95OrqqUwf3tIptEMp24R8T+6EAjINiJhasaxCzdgEq68UgE8eIJolIysOkTVRS+5FXP
8J4IwXl0MeEEapUIBRiepm4ql3MSyQ0JH6DqiIGtbclXjjRim28tiRIL+bP+qM+kDjkgHxQUnHEr
drWa4gcP8zMkq+/OVRnEW77EXOCp0k2dYS7uTyum19U9li0CzzGHnTRvg8pfmh9Aq4aJFzTZZpmI
y7KF0DJQSiBLDZ6zFsceMd4M8L607wniMqfvtnZpz6uEms/t64dtZUCNheDkrlgxRVPWwSkRwDCw
9bT0qu4iS9xhOb7Pb86/lw01+RUdHunduse43HCLM9i7Rfl/06nTB+xXgI9glh/QCc/+g2kw3rLl
DPcjvsxAGRix++K3z2QRmE9aP5dS1Y2uXXpE5eqOQmUHtD8BSXP/EzkUWK4J+PGtCSKwagQpGiWY
SiL1y68ZqZPr1S5iGx10wbol/NaS1jjCGCDwb3I4V+285IKrgStac+EEu8Y4PhQnkabYY5iIUV9R
7dbIpcM4ul4C6empQd3q3qNVRiGZk46szJzE88BIuQOeFPSeBsODGTU9M0y9dcnyCJGrNuIDcrEB
EmeyNM2DRYGe8bs2N9wCsEwndi5V1BHPvqaxmrEnJ7cwE66W2/MyBVk5c9gJv2oVST9K543C4I50
ailJZcZnrirQU14s7ewl6e8YMrz6IDbCaGy+m+l4fPaD2CJgeWOtxh8A0XV/Nj06xBSJyO6JATKu
49Naw5/TUG/u8gblRKrQevzaNMbep6k/pDNxEsKLLfb3R/mKrIrWDFL6JHF/dSo2Klbs/zBRlCVY
6/7WLlPiiQdCGv/3XBAhDFFnnQOY+qnN3TOKPdH2KEbSktClNwCdPMq2UUMua9yd5knBT/tm4+fO
dXjwA6ArhPqz+U2bVlE6j9PxHiwnUnvhLk8LqXqCo84PEMvFui/hDhEv2cU2U7M8n8/ex4vxvHEH
tlSs4ZWyY/0iLgkcfdy052xTL7HDeh7wrcpShcKgTU840P1OFFBqOzoof+cCLYAJssuKOrAVGZcs
h0AIwaFhPx1pn6ANzFarJK1Na97HsK9OcIlKigjaNKJ99E5k8qX1Dvj+LzicG/jN+LA8RNiu45qT
ijH2MuUD2Vnjy7l05kj9ulH8LIwLQT299QnO2T6BJ/Ld7kLtjYQkEDMq3kDaomoMyJ1AiY/rlPIl
d6LaiHhHh65ITjDrwMfqnJgu0paMglHd3CqJlnxlAJrun1lVh2gglWinq5f5UjJLC1jp2y6Z3M31
8614HQAUtNlKEBIPg5rcUtenFTFk56HFw4c87nEqrCk+WzJhCyF0ezubJ0pQ1g586ghvstBsZ2H9
OPnuvM9ArK6H4Dj93XSctlO7hjIVFJaIogYBtZwecoAtgV/hn7oM89piYAbh/NqMT4fYkYIj4emk
7WooL3T7dD0ioV0Net8oaUqwAQhr23sPkw+9zyJDZoL2X4wltOeCf/JG2VT0JHmqkNuLUAzUSuMQ
RbKMgaAy3tQW+GBSjnOYgCIZJl83V4OGMDWMNhXrL2xnd1TwiLOxOz5mAgccXU/MEve3zp+3ryW/
aVzf2b2q76Hm3we1ijBIVSFOz5CH0fCgIE2X+Iz+DPk9EnB6xRNyKVKu/1ku+iMJCCQDcPdPiyLi
PQuKPWjx9FxKKxtArYK0CbQIYcWoLAx+j6HNRgR0JboUYm1eoRNQb3eCmnPjvlWG2AfHAayafukz
TIjY629+Uz/YxuS3k7Igt+UjVHgyu0JjqDkQv4EXtdRp9iJvTbnZcauqEpxg7FwE5ezN1jR7gJLT
RybFPRd1eKkNc9JyNB8ZvxfT4Ar/ZkwVtcIr2WMhlELoLPfZyF4sZlxBR2WfDnrTzloyEps928QU
bZ2dxREwYdXijf6R+0RDSwGh5HjOeyeAOL219oQYV+ba8xXlwBeslJ8BQgpK+5lc+uq/qFRg8KvP
RT7caNQTZvruxizuFQ93U3tEafsdR+eE+eliNPgAN2s4DNIYGy702TeN647ymSfXZbDBJYkcjseh
I2feiKDOoVhgwnesqwIG6EIWhH/xOCs0IsRF7IVe6fabGbfhxuj+0o8LKGXSZB3o/7/X6ijqCSa/
lYPDXee4MqEOYLh3Ga9qfsfEd+hShnCVX6yjPVuVv1dlOKW7e/3xu0EA6zZoZUvTIAB1cc0KbxHA
C8u9x+jeW3W86gpFOCct+oRAtoRTvfUv5GX7W1BE/Vr+ONMfyBXwehqizCC7fDwW5gJvH8Z1o7VT
qz8sw5TtBYMV78voiwQHNHwCzqn91fp6UIiv7+SmbrOcT2b9a0c3dEfKFyekByGSiMSv7schjEnN
8zZwA3r/BwOu5+wlknnxxrhfVTavQEI0OGlTAQH5mNHkHKxVmzjChUDWzi0lx2omY/z2uMOrK3In
I0J2NCEZdL06V+vNDJEsJo9MFAlhTRik0egBJG9NnojSUDKFNzwKWI+8CT3Vm0Xd4BuusS3nVRx1
TtJDdZdmm6XnczipB3h3kr6OLOuhILhBWsFWBYSDdz4kxYN9lIY29shuNedKib+K+ACSyJkIm8eO
nbqhUfW5fDtXQjTfFxvTgnXLhBV1tBXdlh4AdW8nACnDh2x5JAmDyCPHFrb2I57U1lPZ+EeQMyGB
0Vgy6CKs5WzXIPAKVwpliybgR9LYC9BHAfIy5JaAmjmfKiSHhRm+MhtC2c0KUco26H4LZSBnc7dk
otIxk/wEOa6iKt0qLNHslveYaXMpDELzjD/bR8bO3aDjvJiXCINS6v7B3CyggIA2fGxKNOH0W0YC
CYVs+jEi1eDp12t43qIJS8ULWs4KGK6Mx6nt2idHFyUIB2S0l4foTRbVEgYm4biubkQhvovem+QJ
8YFOSQQngxVanDlKr+hMmxuQOg22fuzPjWsFT82N6USfijUHtGozvVyOvPNFxRDSS0nHA+crWZXb
AYRXrYncAaYI6RnJdCwvGP+Cq+2f/oWGmLZGwel90bz7PENKghhbELp2rtlvnfwuULPRQjPoGNgw
+Dr6y8dLrxpZC6pUE7CmF7uNt3wpkXmpw6OY/v0zmgE/kFhZyofAORlJNWyrOo9On+dt64g8F2WB
IIfM3H+AzORwHK8rizYpT4yJZ4fUY1R3o80AUlHLKAVoy8f4qfkgBQfCshou8T2QirFhYcsWmHqD
ARwALXZbz5DidIhCNt4N/X9kpKLR+HqT0Env95xPHXMXHAzDRMKBRWfBD/2gWYQY23jllwELOxkw
RSYe4VqN0ihJX/rX6aXx8yuVqPumEv0Fm/oWXl+lug/3YfRKKRJ2v5DooF9Njcm1T3dEWkFiK4rD
2iU1mIRDVNRR15H5aWCxsOU4+g2P0ssH8lN4sifoKpnoLSwjCBMcFO8rWO701MZF1ssIpQsgOVMR
XRzZk9PXfCiH0NJSP1yZM72BirxTt6+LeE+wPgOqHzJliS0h3k5sNnjsplIw/m2ISda7JUGXdhAF
Ftembw+p85xGokkysxwZj1ueWiVkHSqEcjarCWGEyR3/59r6resYEQKSb1GnKa1eQrz8VN6oUIPF
w9zfDbMOuKvu/DKBLvuYaHhLrzbxRdNXaFr0yka8foukl4WLVw+VMeGhhcllhTPSb1wLO8eipdeb
ogbXjwpn46eWOC6WQeHoW893+1G5FhJQYoVBDwm9lFxmzHMATEaSdT+0rJgjKct1RJmrHMoqUhyf
6H6PA5kGI4UP2xUKjcyBD8lQa2YReCAVqkefdhKsfttjeg14+UYBA2iVeU8LGyqJGEUnndhSb7cQ
oXtyVZibSO4izO8YleHpdyIEc+4Xufk4Zh+XLnVuXdfzTIyP+EwA42X1gDsruK8XFJ+j/Y+tYEJl
2wXf/AM0/gMGkoAFW9oIGgbyyMHPQ6an46rhVLEnlD1K4wJXEF8mwQwzKfd6CVU/S6Fda+NLyAbG
M+iCEhM+0RY9wkCk61f4mNUL0thq2+L+Igp0YzuTzSygOz0qSXsYRfOkkSyQSPsomIUr2wOFPItZ
qiKaSNpHXWiGv+fOGmiD3RiRlukSSNzRDFWpva0GqlL3G27NmEvbF8lRMdJHrkIWNJB4HWFrS0C6
2SohWkoTSGSgm+eW3BRzart9U5LAKB7CUKVjWWI5KnEMHXzdPL6RcdKGbo/Q0gr6NJ39mLGQMeqa
mLS2KcDVfCytUfi0dZxxPBasLa8C/jCbbLw1IA+PW2Hw9gtR+vtESXd8msXpeczdd/dWVeuFF8OY
LuFxmL7pPux11qsvO3c2YvdVzQoEQ/OucrYSGau5+aqmqfOadnU1H0zAGm/aB5dxGm0IYDNbX7pO
I9ANAeN+cuDuoBNlJff4Bg6t4wJn5fCaoZiWHFbUkaNGLhF+7vGfFti6nDefnChr+nWzl+NTE2h+
JIMLdsqJXHmrSp3E0aIjX/nEY9B5M1dL37J+rP5r45vxZkhlmuFX0rUq1YFgyR6Lgon0jehfk4k3
/P/XsXIvP8+CNJEGAB2NI9qF+sO46EbrbOrnhSL7k/z9IPxQKcxjtMjzld1gXi58X0mNalONTqQ1
3Ue3mHZhulUFclLsKQh5HrI5dA/gDgfETBq6zslxTNZhr3MIVufHpYCzsoQBSB09A/BfeFM6tgEP
cmmLFUXjtJcsifdIpQOAzam3LV5InJSuU9bFjVUrEVzXUbe/YkQlXHx0Xjek3ojHMXDtYxZfWRtL
c/5+kdMJMg/3ahh2byfYrsekMVAQGraasYFWw5A+3DpSqwy/q+0OM8FT39LZX9fltcsj5D+dnLd1
lIdCN2rL4faRfboT8Q3Vz9baKHGzV9pRcqCrRq93NmJ30H3uniZfF6IQMlnfYVk8n1S7e6PXypU3
pEbRQGlDAajin5FMZgd9ssvl4F4RKJqxDwuc2aWY7Tao23yEKiNy8lMIB14T2VmwqpuFhSbRPqZs
pqap0ZWDEkFJrg9FBpzwV6yw1/U27ZWzjvwDd2AIVx6Tgh6WyOdXj6VwhNLfDV6+hfBnpeWJPFS6
JZmiXJ/Ehz/ATivU85Z+JvF4LE7Ai7Q5iDdRz43iIYGW0207vBE/4PzrE4juixzOvb52rh12eh9E
4WIcjiuz+K2Gb6HXJ8MpClCwXwoU3qFsxISmg79bM6oHlIZOaZtEx+nTaSXGPm7RedV6PNRmTi/a
AhJkPpWQftAbbBW568GVoud8XMh+P5SlIzuYxGeXrC1cfkqB//cFbupErpoXaBy516etgNcwUw0X
BpspUpQErDDj3TTSQouWnSnGroQH/NvjtsRsjsrxjht2SWMxX/iYuM8NQqr0M0fEmUHVQa84pZl7
F+h9zUfdqXo4Sg5SgSh4MykwiZNHrFuqpGOgsEwYrw2zyzq+i9CKUCx/ObiTPbr9sKPDhWNryhhp
rZFXkgD/S7ZMOcYwgXBVkDik3UZZ2ulTEqTAZX8S5VIfTBMngTxx108qlZhLgo3SUhYmnkL6obr8
g6LyZgV2XrOc7BOhVix2crSlyAshkC7CcArX9IipW6iHwbhMF40BYHjFxA8JcKhZiW165W7dEgtW
1qXUxmzh7bzOK0PapgSOJNT4agckVDRszwp5ppTsAxiwNNSwK2XpqZrY61vC6itru4QOvAGLIA22
pCG5ilVOvd880QLckTT3QHL1hHo3PWQ7RG0NvMSm/4WaA3RA72hrWx0hiwfSme1savxFAUcFDdop
mZZxQTkqKuvvlAZqj8Xjy4hbzRGJkNiFC07Gn6mw6oQ3UlnsVelCZjizclo3yDd1igqv/LNYiRxB
jmETkfLYESP8ma4fqLgc/JgIWEA1VmM16PN4MI8Q49roRWaS8vSV81RmdeEHVqn0u2/hiRVMOfoR
foxvvU1cFjDn68COgksUvfoKW/ROhpc5J4iFpdA7HeSdSnwott+fr5n0vsUCISDRq6Su9WXlKpaO
kEBhBb5Pm3dRc422eLzD6IJ+0yPuGpzXDeJpsf3CwOBKC0O6NzAh+3nc51d93zhVU7SsFmpILK0A
zyp19hXY0PGLmMYzfcM9RoFX7LtroCbB3zeKiWi72ODzbwhExs+KYZrzLLSHePoAI0TKXqLB6tlV
VSvay3Xd4TK5+Y0a3jShuH36t22BjeD/A3/CwcqC0kCYizYdVR3dnm9mrjndABc29sT9Q87H4lud
1PTNr+vMaMjtJgWMITnhHna7pHCdun+ES6nBmfCgMLsSXkR6pn2FU+mV9/Mq3Z+0kM1IY37HuVec
TKrzczItR5YXeF/suMm3KKrvu6/9BvblR8UKHZJeHVpBJu696NSUDcanbOa2U4h2PVdwkvfa252m
eCsA1ule+a6d5lht3tUDnni8+MelCtz0Ud3ARpJdLt4OU/8w13HX7rYVYYHvb7kDtfi1PFwt68nb
9Pxp6nH+WWvyY9zHjvBhX9TqpclPJ9nhgwTlELGhjDU5j9v+6MhceiMszZAzDkXS12lfFV5wh7TO
caKGju6NWhFdN7BolO2feXfWC0f3v3nzfTkOcS9g/h9RsswJB3DzmPjBRJBY7ONvyYf63VfnbROP
rQwlKojeIjdqNohMYokjHh/Asp6FEDDvKbtMxP/b+v9zTi2E1c4ZGLDr2ewNyLxM+6RM00FqAJgL
ll5i5izye70dNbKSiMGHqZ1I+r5vQob5O6BM/OVrRjEK9zWQjkn7D9C9UV9k4sRc5F/96PxcXKz7
8uGi9Fjp4s6liCpkw4kLoP+c+gRavm1ie7Ut1VSJa2lQQKzqrcSKvAvKmsN99dJxAf7aeAGzD/nX
a/o7H5kAWfA8D7AiFYIlCh+Ohcwkz4iNuHOh0NDhxrMen5iRJXyhFj/Vvos+RFeUMetP7vElIVaf
hcZ5VdcWWdhA7ejhkecFZkQ4hHJS8A4lo2lu4NxAnaxmINJs3vAdbouRRdemGLmuY7e8FNBvdsRF
j0XA3EBI8IEmxpAbEfMFzNqXs7EermKZLbkadzvR1musJGG8s8QU6cL9+CJOGXRNeUzh2/ZKUaXY
ADmbG9wAvPxvRgCipJyz5M6Qhy2qg74IV4WmjEEK2L1ajiUSJa6OuFs1flHcHJQXN5V//J4mSe8x
nhVl06varmEQXuluYf5i1iJ+ePKJ3y9VZcKZr9SrltfNnLBgk+TddbHoc+Sh5//VwYPuoW/0MmGw
Vew5D6mv2DDUX4DNNbItJiSG9ge6ARSExWtImfY6qEqWlUXrl3pgZKaFu0B/IqqGNLiuAoNXUrhc
QGohr/Exz5fRjkfdqQSGBI/0VqSfyDpEoGYIHtgAQf9XBLXON2jxz0TfquwIQSGQE9pXy1k2TGkx
+sVK34aBc4uDuaEzJAFUy53TVFIIX9qC+zzD5Osxrm3MByRTFCLyRviOELf8o5vN4O5TCk8rMgzq
7dvO4AC3d4pBhzMu11N+UK6NHPlkOeSecckKKiP2UJ/vMVzaXH8QGsuPYhMwHzHyJUt4VAh8Fxiu
dha2ncM2TWH6DzVyTdIV5gmk0ZwAsxxpuKZ9fzdTslSvHPqrQrnK9XGMLKVMpYx2k0eys/31pN4f
KKKraGX+7kVuGimJtfMJhw2X9C9WXTVtErOv8xyYJ3N3zmUye4jn1JVRQt22fExyf3fBF8gjF9vZ
CFGN+t6vq1jy/I7c6cfd08GEBgU8PPbNcaB/MRu53AOrUgrWdUBieAh8dXJqoZZS9dcSQDVosGAA
ozdGtf+xnhA9YluTbIbHHmC909qj/zHnXAFOKBE15cQ7EWXfwqZPiims9XcsGTb+vX6UekjtkfWH
Xsd6Pn0Pp8+rA+4tDU/tP6nMbEXlE+32vO3QKkNJWQbz7WeiVLXw1wcBQAcBnRtdb4QPjfKSX05j
9TwUlf5MMKszlDkWnjWT5ZtzXsxb/MmzMxqD0nppTC0ufe+Zq6XMtYXTyQKFoRlzLOcMrZv0SlYn
F2W6XN0x2i37M389uaicksPDPKdGPiqKahf0487V01vlRQXjBOzUryBi1kskgXCwzB/n95KJIQNu
nJ2qozQdSFolhqYh4S73zmAG9HrXyH6ocZaGspbMF5m7J2sXYch3Xp5B2bsmdHpvFv5IwK1ZCqy6
yj69PsoS7mInNTKzFakzdEvIVDVxSmWUEE2sOTqq6Dos7yctS9wzC1Tutkj0CTW5m5uG3unVPNlW
Hhoj/NadWrLyMWQJLAmSxxuRsud3Q5p0HT2UXJ+wqa81ssY7NoqBl0utcJAxFMiZFVmsK1CDZ5Vo
Ot3CTtnWjxAP4OldEh6ouVlJTFG6tFn+nyLd3f5KL6ozakZ2I3IUPgrKeWc/iWbWNwLuqBaHmxkP
kaeEZvT608D4tOR8kW/XEeasFWLStP/faRYRhWTBhFEWweJsPIWDwk6ChJ/ge9thCOjpl9cksV++
1vNIsHs2hY8fownR0SSdZl1nQl2QHAH8TppsI/rsKkC80C4vkurAwCLfwOB8fTtriuywf2smILFP
+81n/b2OXKtpi1NuEwrAryQ2okw9jrOOdIuIbEZzT8sqrskJmOu88qj0ygqdyfdPXc3aXOAKpQ+D
AA81VU99iSvOMVSIBwxRFGJn1hNwU/MY8M8gjbyFSK+qCyFdzLlZAd+w1uD08X1YPWC8gy6aKnaL
mk1nXODExY/oJH/zMWqXiatCZDYMGNiPOo38H8NoDHmBh36jYpaXvQZT8JwQKCWunclxDsyxekB0
QkpZlUc+4yAu0W7P70pGAvHQGA1ZP4BFmzS/c+h3cDn+AZ3YvjvMio6iMRs2dLN3sCOj1TF6CIWF
Ixltxsf562WurMi1/qExbbeyeLPiq8MWFgVJ8QQFM5vxODMdjQ86Y0pntoN6rTf6dbCF3jLmAjEo
8UChvRIdgYbGWy6XyILT1gp8v7eelpU5pMvlScTiX5XDOtj4uGC1gRZGPLwqmkP+LO8zzLHMjbUC
m6ZtNCWq6PaDgZTnja0fmjqeY2LcH4wo7hYmYcs8mVPs7DSQLrC40Mn4aCiSPP0cCO80/xBiM4TY
NVr5O17Zkkac07KhZApB/n5+aAe2+yF2CCBcYEiLg/f+yOwH7FbD4ITKgg1iRIbP0zYEM4OYlTTh
PNntQB3mnSXz/yS+pAvYieqgRfCC534YrvMFeBHKyUfR/hsoMbBdefT3DGwvZxA35NBYRvcCv/R+
dJsGmDuBAqUa8SqtAWXgfEG9afhcpHtAQ8HiyHCYJ3bg+o45XmN+L/SkqUqthPyZHbeYakFV3c6D
LDYlvLElMlQDXdIcJVMfVZYaJwKWLNLpZFO1CE75KBGaDsTyfatvo/IkcVpBcc5X3Z3HQ8Z5wgAV
yW8ENu1EFjpV6lxT7wHGN+RvoES//Kt9P/byxHAt1IU8yDUQ9XpmXZWEfvfZ3f4d5B3IQbt3yWni
7ZE/hqe6ZBC4kqCCL6TQNmCiprMAV5mpfkL9ZYiD1Twd76Ma9hqxYOY1FCtreeFg5ZuK6p+GrZwt
MtKbz8ISObMUZgR1YTTclhsu630WYnJN4J6uAqZ1GgyPOxXsyQc1vlqpscyfd+sTVz3N0MlgoG41
3Zw7Ave0A+7hYnxf9VlTzrXY3CMKWOFxcu9dv3AgcNA+xbwFW9uJSJB+tXscGm1sbT955L36o8w5
xcIxo96wbZSotd3JJ/st4p9rI81vd3oKTk7jl8sRTdewjtbywoYf4wxbU/UZphYxhCqJXvV7SYdq
1VxqlOLGd3HGSBwCbMZB6ngZMDZX+3Vx/7lhkesauLudw44buCUNZ2m3syN2+SCG8eeGH++zniS9
Vio42oLSRgfqtdtPD9SoEoBs2TbaBXtQwI5kUygTpV/P+nUGxQIoa8laxAOcbNWE02sy0O1nz7M7
07w3B16DejVl+1elN2tuVUwYwJ6zPJ3CYab6cQJQQoCU8GoDiXds1wOJhadqQdcT8pWrznGh7sWm
palh7lEoH6QQIOiDPrG04UBF3Kv9gge9TiBR3bQdWjTpnaFQJoc+xXf8CsIxORzaJ4rSg3QZRCka
IJteMYsfQmqdFT09wSklIQbGAppIg+Ga6GxCOI5hg+cqk0uToN8KO4qdRWn8q1jM0/HsXN2xx3w9
e0cV7Yt5PwIO1cwhvKYN2xGOtU0iUOk6jnuhW1Knx3I/rlZPEGgPPdZz8tzJ+OGxN8uAjSlVDIXo
3uq6PmYkttM7LMmL2gwOfXQWXWkUiWLNpHXEtvy3pf3Vtu0Yfdrb8JWOedObRCM/e4D4QVF0YoU1
VHxHF4YS80oh9rL4y2GRp2IVjNxnulTmYLvBPCYOKKNmuw5EKscCtkq3NjhS1yfw8u7BEhLexDvH
7AcrqjfMr5SGpH9iG58wvoW3oQgXepJJpMNGVqHD5LhvOgUZ8bWunSh6GQKgH/atehggoeFXm855
UJP+v+uCsdSPVxyzbYjmtFPM51nkMpXkSzzpWW7XiWzSkkWCZOv6lpyZFrhkBJRto8tWb9qOgDDy
H/W33bL+3tvvDD9RHvfJhF9M671vcRcaoUyhNMItCV/RLiJIgiroV2e3CnP6QczDaCg2zCLog8oW
dzvDpNALDSuEqnJq3f8njxPnSFeZZ/LyBxRZ1FX10IA6TiuChSohOjQYYRgT/m/HRQWVyhgz04vH
3W8XVsPYp43iTXR5482h1nK1B1XV+bkGH47Cz5Gsz+uVbEXH2Q7ApoOrdheF0lC5ugjSd4EwTzag
eMwShjtoI41Z2TwGFNKb8TcvgVPQztXHmcqgQ55WNRQSFr0dMW4xosNYZq3zslinPbbcguhCx/ej
McY1GVL0xxnYP4M7DiIckcOravcQxbWNRG2m/7BwVLWFetNMP20OKENMvsyPWauRjp5gSvh0PkJD
h/SaiI5qk2CXDnQct11EDFLcP801B8WfPy/Z6pf3q7Tjt+D8URXescEz9fMhemLx4KDf9oDgftPP
Nv/956zubUFXESVFxT6qhcQnBPPqGAO7LNA8IhStO+tHNh5cqLhtL4ghpmfqo5vu9qkUp5edjpHW
ZyzAdK6JahzBfFCRnRrg96MYWcH79oKW+dFu9HiOkk0pb8POMB2BTDh4jmpUsw7Iew1rMqq24Lbd
zAzhnTpc61AbTdCp91M1055PaSly+g2eTNowjQt9bk2xK642XRe/t7AxphjtRZGz5O0u32gzqs1p
23XZM+LYovmuMunaZjtiztTTb2m2dVN4A5/7afx8j75klkmgEy9jjuTT8N2+0rNxKXIIi9vrfGXc
Aa5PdpgfeuLCfdM21O6mxFUUOeX5G5d8kYsGF1aGXaSdYtx616hMrdtfC5IznzpN8Sltvmurr5fE
fcz1DLCGzK+JDlKOV+yd+o8Ib92eeqkOn6PHBIVSRkulgM97kIRwqru2pIOytGHQCzOw2ENCwr47
fHyzTk9TDlIRxi2ivBiP2LKmpuhU6WQdn7IO3lT3GJ/uWsJ5s9LHpfwQyHxrr8/bXxOBJFYdgXRG
SGJ7qg17Ge2xCd/gWlIhij5FKkQggQhb2ZxHt50y6Ayx6aTLnbslGHILln0UAmvAi4ssSYSECJIo
disgT+X/AmgXNkZxpJZXEPInsjXOyySqOxjwm9pohsqRps3XTtCQreXtydUKYm6zqxEFmCSQK+/Z
E0HIIPoPkvNgx82i5T+90cA1fF/8LZEq3L+XHLHx/r4v6XZ8jBTg9NeCyW9eL1t3O58SJ+zuuwWm
ziAXIc/XLl0y9M28AbpTumIqFJQ80S0ECP6byL1CDuOOvHsiFP/atZDqCqyP1NR4xcHQd7XS72JR
CmQpyv66ADBVsLRBVuXPCjROOR4eV6hQB+TiQq5kgdg6b3sPRlnDZydcyrnb1oGmx3L17M9vrGPe
T2pTZ4Bq960XC2wkOX3pICyzuKD3odFd+ajuy7OqHJfL3Kdqp1OaScHXsZMyCQKAQjfZs0UOvRNo
hkj4W6flrREXq/MBQtFkCBnjmIEDAHba9IcPSDpsMFMKgxe+8VuWBGtrZQOIYmCDLfkjL/xTkfRA
2EVzDPWrv6daKCxL5ll0d3fC4FnQQYHpZCG8BHFK/WzJvBY9LVuky1aMzpGcnjICJkS4IOYhkMvp
8YlaOrZJYJ+Elq6yF8JYOaAivPsUUL6aM7O3YJOKaa/HYW6fhCOLiiHGdAH9nCQoXqnyS3qHzrdF
ISbBJKMtYtVeU5dAiHFrJTOSxYUg3fnSSB5mq4WHvZgU0BprU2hXyLUQcCyFO0ltsv/xCfyQfS9N
Md/je2MrqBUKUzaciNJzQgg5jXqo9nu+n5wODhIj8Lk6afkzrkT2rPb3EgotvvRHz7y0ZPpsjBDG
CVE8sw+WqP1vH+L5K33W7ch3JtlHwLEOK44Jj6+hit0zSVczIH+qAkFa3B1h1/4KncnTxaM71fDi
4jPvhxQDgLdiVaD6wTscWpKzeRKesRGv+GXbX0Zk/Qu3JjI6ynG9Vr66kRNRwnOR0Th6zNv6FxrI
kULhwm5UKxhf8HO0bdmyQBfPEfq0yCWz73oYKRs7QbhIADIWWIMG8Z0/oR5xlZnApGP9kfldm/WQ
4ucNXvvM9lJDfQ3xtiZwJErgve9RHOTc56mnTAL9UsDP6BFOHtEkyhM+rbKdGyS5o58WCDuGi6SQ
vGo2/s1AGPxTqY3zD+E/hBhXvLHlBUkcPDtK+m+cRre2MzcqLnhlModVneabO7jqBrE4H7l8PD9G
+wfCBdwOgrwtNmGxgBTdYetbKPLUTqScHlbh5mj3/6COdHjnwb2MXCBsZjUI59ljFjXmXcYT6sXO
OIv+06N1OntdqLPcP/70+qdoLGs2X5Dr5FgiHzbWWjwJCW7CCOrT9NP5Vsn1Zc5QnC09t9k6kg/U
rDkIgNgll4P8JjeB3HN7hKtlDzyYg1+JKSDBeDfcXNwmc/cTI/j5hfG2x2NY/nXaXJp+rIsSaC6o
PJryatOzYoQcJC1QMvACPsgMITbFzepFS9ZPFY3gDw49TIHoMunN7HSWwjeT2NkiArM+XIPVCFGQ
gevxS0qGKklonXhHz3lapP7rqPZgXH/uuXtFOHpmrAv64QDRFU9HIfYeVovUxhdfyLux6vT7ip+A
FubTmGm4iq/UgtGp7Cn4Bkwzi5l541fxfQdb1AUbCuwXMNrLG9ZgMW9RRi9Lp+hZjOD4S+sfHSoT
HfTJi7kzXMex02XDQUe4rxTxgItySVnuH+XHfwTw57zdqIcMFnUKPT39c0+ekBpWmlGQqbcbPi1d
O4BRspzkboDXvzznSaWV5fbfyulRRWgeibzcq/aNYC9UpdyTY9JBOr2qXwBpewGnuaZpR0ixlHCQ
jjZfWw1XxeeDwx8IoB25NhO90WQypSVao9dQW0fPoVYPym1A88AAOgd0MoxiBP8D9O6Zr6qPX8f9
MWT9ZSASWAxtZUDEJm9eH206veANO+yUlpdqWcQiYdkz+n80aKoF7yXrdL1EAWQi4SV2+Xe67jJz
OxVTKvFrcW5B9ggPW+DbBorc00eNAmK4YdkOmud3dbqF/6u1EDNWg8zbtM7XNslZuhv6Tn+sfA47
IWpvrT9LMoN3EfuCK3tgKWztovvEmjcFLx9EqG9L8QIVH+FFf7SCy8Fs1qUejs/wuFDPWhjZBn4I
34l489LmaiB5/3TWqJyJyB2V7ZjQzPtpbiI026hVAY5OHNoUNnAylvu/vbuXnCA2zHS/HIqbJIJu
tv9r+5BCPpM7ZAWw2kg4q7i+pneJXuWM3FpY9YT7gDA+Bu2JBKAxHr4eYp9YTi6UNFNKqMSlkoZc
VIR2Howpd3FPtv6MqQVl7FusqBEs2wibHbIl8s1j7P29memM9iTT+fB4DAcswSgwpFcG+xsTc6mq
8DqLVwzQf9Uq0BPG8NBD7RMrEBr/f5cr+kXAkfmoJ5wg5RAalpO4jeqntPDlSk7nNf+uvwtPIq+y
jnhUPjg6pvyyx8f9COXM4pfuPnc3Vscp2Uh+9W9HaLMNB76FDSfQ0cbukpt1bQmhpxNihu9NeS9w
PMsh0RCTOLmTPn9ojg1fyJt232GqNPnjUX2Eqo/ra9YhEYtA13SEBFswtgaSVXXi+Jy1997vo7cG
szOWGyEa3CQ27q22DRsp1QO9QKp0sY+t2LiUS/+phR3OEWxXvc3Ad0Rb3qXakwNnqg7twksQAh//
bXSJnWq7NAldFMmEyti4CXrqFAifwnbDxlP7xylhx4zunvicWJXP1GJ4ssRl6eKvB1rxsybNDM/j
UrJOOfLabQG531BtafYubIu10zOOyS0QZVcsFuU/HuPKamz0FHp06nQ7LJ8G47p+zPZ54iLCWC4n
0L9ljzfTsxEBFGiQMlIkWwymTLIkExaPOhIVxdkUjPjMasbxfyJ8D28AcCYcaoXjG1BnCpuGslVf
VFW9Zu38wUxkecmDKL+wuh53hixvhFVRs74JEuhzXUBPPKyJwqXatZn2BcmKDt408W0sygb7tLwg
rGOVA4K2BCSsB8oSZVKBYoef7GE31pvSLl3jEARZOe736/ZW7rflNMA1PrDpiTh9uOyAp0a2orB4
z2yy3DR+mUch/kxiNwo3RCkCwHrfwCKklMmqr7xO5lMEJXOUjCC/j2KMqT8DHCiGzFCpnaiA/Faf
gAfidZzctGD32D7NYfH9jXCksssGroYm/u4LXEScXJaxk+XgoG5UHhR6DqBoU+fjSufxE5D2pqGK
allZnv4ztZTm1WB48XhhdaObwFbeJu9cXQ9wfl748xfzQaEU+dJSiXi/ynPDJgHZ+lVnmsAnob4O
3nIHpX7Bt/Yl7BkHWdndUJ6qzVgKAQyXZLS5INatC0aSS2DiQrZDmY0NkhdYwcKKz7c07J4YLcRZ
5rjm6j8Z4NkyJj7m7ppAuXvbyeMM1Mx3/7wq3j9SoafNuHmXw2V2S47PEXy63SmT8MojQBztbEmZ
kkaalRjFrjSymahzU9lVB7JiaqLQuiJ1zs7XS4WjQCyjuwZN/61fCh5QVPO8rcVKXxNccSNjvLiN
ZuGjkZHw/QF2mJQfZcgDgdK236Q9EPgk3GoeEFDKCxE7XY3tR5hveuAnImslEG7/AqjYgHDXA3Me
+ViXczitKw+MARGu478XyHpdx/cWsgPhXp/TeJecvggNpMJJrGbeSs/kQJhHKKhJ9r6cVeTTH1Sd
XxCBGsLk7h1Awe1Y4jpnN3MeS41lJ3dHFbAmYcYQ8VZhkSpTcqQJ1IARpN4TZIBlmPpmkTwM8rQj
pJAPKDzwa5VoBlbT1nDB4dyrqAYkfMnj0rMM3h5aetqZARHl8m2iFbJgHjy0ALRH6ANVkAyD29Wh
O5VsyY0xh4iglGs15enwe0Cs3vfb01Q7opVDxBECRqkkY/KQgxpC1ONqIR4NGBl7zH649/egNIWe
mocrdYeQ+P3a7+AOhx2e0vteOLmjy5eUf2Ur71KJKmcByBfz70YmJI5sSW+ILryZKSCZRRkAsLMS
8jDGjUmv2UzSreG6/MaRd3+U3QcAybC3ctfSwYvxgekmeA8SgpPbh9uoJWYSXMHjegP1HGweB488
lSJ+BOVekbzwDVZjFXL9AX0J0/o1MOb/X37Lgi5CcIzRnhtX9FQJrbMLIVrEQeNZQKmHDmHfYEvp
yO5WZB4N6AjvIXC99XLqIO9PXIozt5X7RFW8C1UzEe8dywgCdJU7Foe4/ZgjJPVOwmfL/k6OrX2c
y69aqCUykU1TJU/tfbr7MuXf3ThIkt0JXCOGdS/T5aJFIJBtga2J/kcBEqxyuRpHZ/3CIWPqHggl
pkA6RDgmZO/KBjy05+B1j05SoGReipQTfsa7u/6uoXeU+/mS6yIFbB7vT40nhbZndMQst+GbcAma
kB4K9LLd1hVL3RDhyg27ZrJgfAhJAqirp+gnEgH4DdjvhLUuX38yqg70X8nWaRRwcvLmKhH9OjJu
t2193ku1oaBEuRjlyiXQn3XxNb187NhwOaM6Ixxl3lJX8TRhM75SuPItsn7PkTVQKLj3Ui3u8+YN
qWPMvaHc4uqlJcc7fkRz66zbmXt17164XeYcHA480JJtRseMQhKgCPc0VDJfatPm6deLcDtKZXUs
xOiSd0x/VXtbh6BdJVJe/ST7bWlyWGcQ1bo2GfELsYok6RQSWc+v72LOjY5+AcVgYAMS+pJwu6ao
6Wo/c9J5SC94mOk7LjGCCH2hwBt1GwQ0nC8l850+aIFcjGJBBYqyGtd2UnU08f7y7A1h2HUPAuRA
lbRwIgXPksvCLnjgMjytH5rE1fA4YwUlWdh8Y1kHT+lCPLYAqTzj7O2JXKanp1Y+2BfDX/iisP/x
T3LmZXDToEQ/9ly2bH+JU0r+i939OyVQgKZNz5dqp9cKvqfW7H1rBc2tfZ4v/yIP5h/OaoYozykI
H3+obHUrPjsBQiZrwgXf77uSLWIrRGoCw3m/wy2sg9EO66bItVr96N8jgm3/ET2ceK6w+sli62p+
f2LErFCVXUORhzFrF2BX5JI9jJpPJBbBKVOltKFIrAuj0kfMc7Mdjt8oc7VmU6KMhXMKcRCfGUdM
bjMkrx2BNZXJhhLp9ASu1ZTqVmFUSkEMcQPHpe71Y/pOIDcRAIKPXqAIXR+hS9qeCOftRwH64HLG
LvOPofF91oYRL7NuJBE/Zr3ciXK9ZdcJr2t4+nj02VjNdp7Kqeevby0RYyJ3kCqgbe6cki6DzlES
gWrG9k2c8XTfCUj256SPxpsS530z5n+oX66rudAee0MeXkAGL2bSMexz48pglWuvJVNEHGojB0Ut
Qu5BwpD9eZ6v8pVSdOuvC55PEAIv5FD7L4oCyGKmWfjqfRp2MQagUwo2+Ge3SCw47tYxvJ5diiSL
RIKJcPd8h1S0FpeZgbTy22QArAgHY78gCDiLUpu4C+q/b+Xw30r6WX+YEGQuZ36Yh06CJlE1Knl3
5eNeKbnmHaugEjTAfqxNT+7cZkuURBVsRRDAw4v5wN2mIQkE4WRZ8ayUZ35kC7M8qmukPc2S3/7m
JBGS8U2xioSO28xwB+khY7i9QwYrw+QxGA8JqAaRt1DBFQUREM1scpHEN0i9GaPTk/uveYNV2KJc
F3jdgBIUtiI/bbtqF1M0te9WsksOjp3TjpJPSptqgeGn1sfRp33QQqAuVkVaYe44PzK+Ulg2N2P7
R9efrf76sgYp92Sobo7UK/1XN/e5rCxMwWf/7Rn+RVqsHg4wJFN2h1CoBL8V9mCWvEcol5wtP2KO
LOE9O171k6LgbsBuj7db2LxCSAYn2UXFG9y0/iy9q6LZYTzzjAAI4n9OzG5QzpDB1CeGtGiROfID
PTUg+u/oth9908QH67cnn7CnF8uxHgAFTgFG0DPfJqGpZe/YfswrqmHooDXoli3OjPzhKwg4FQk7
P9PgND5qnepJZXyP77jXMsc1J7f5Vo3G4awOSM1T9gSMcM1AGDRSulRBJ2nwiXGDjUQETDOrW5Du
YyDf/Ac2ZHFhHUZk3EQZptOU05ch417DyRyxO1vKNxlwZDxgcZD5TL3m+pwrkUWyHlKUV/X6EEJ7
XTgBnLAMrQHK9kwASuUyyd/M6jvOLqAXs1pRa+h3FVDoD0kPyrzKqn0EGCT5LwbPd/Se6CZOK9Yz
j5RjLuMgeBZj/t4Cu5NVSPMI918RfhW7LAZcY/gKADtEd7xU9guI9spQeYgMKH9q0qcM6cK/0mxo
AaGJB9jJ9RhZKqu2js4U43GIK1ocmT7Hli7vmrUPDGTxD1Up9BkDtiBn62IJ2/WUWPTX7FemOqXx
5TYoB0PUfNoLVmZMJO1N2Pq4eoMbcmWcliwFDciUZxy9XJL0WL1t8XkldRLkdn7e692lP5XxACUD
XwciSblpVJYZXNgyQzjP6mN+Hdi+9pUrUakrQ6f6pRwoK9r6GQO3oecMvu+pPGAPs8xV/zb3JSN7
vhjqLctVxlXTLTN1Sd7D85Gu2CIolreVDM6FzZqgeDbNW7t2cfqnILFsd0SPdNfroaTH8wQtlwvZ
XM6u8L4yViUCKcx9ScYJf4Cc6lKJ0Dpa50Q6sR5IpkTWCY01zlNZV0LH+DbVrxbk/3OaFpSvq/JX
gYwn+0+DM9xoU/BzhRHFmPixZAm5crmLROIXfpEVUAl31geBABQHWJO6Cw+aYhgCDesrGXpEqkDd
bc7XRwNcsYMN4m9Nj1Y6r0EVWwHk73VXCkcVNqqX18Rl5fsIRlGnKL5JLNu8pSkCKPTyPGBuNUTf
CL2znWI+KLwWeXIWS23Z2cEMHXwMV3++8pbqNCHl1Y9Cmv8Fpa8rXkzUG7Aw+5T+SZ5D4RFad6rB
Y8VYdI3xLJfSHxJcT1NW02wCrfryeo7NhFs6U0XbbjHTpoPt81oMTLruvs++g938+Asw3KW/TayO
gEqvtoOXj0pK6bTiCft50SwNlifRqpNNo53wAK1V1B2f0OVy2imviZqV6cMiDs9uXOyhT6q1N37S
fgfdrC0LL1bT9SxRDSBVEiVI5geQUy645CHxKFFi5ChSsKDngHhoQFui2lhNE1e7MzsC5gQ/IUov
J2NcNL9UPoBq3vo7LQIT3oBQ+CFOdqe4ydF3ku8E7DHsc+eVNLngMzUlv72qPpFjOdp6FpBZq9O2
erj44TtnLOQK7lEgAKfVc2vkrWpKARkHq1oSigkVnJxP2RMes1SeRJWJ0Qr+Z/uy9nYE6goB6+G1
7lUcYaKxZrU5VQAPXQObDhxtG2hHsOAeJxQ+8VBDbM8TW1VwBLEX4sNotD4OnJqA4HegS7mq5B/A
lP/m+1NPc1tkToiZB7J+ybfzOe5iZe9kKBRpY26/gYOXLs4xhpz3TjnhWkH6ufhEvHep1PHd5xYw
rvieG8LfbvRdruf/orqGat6Ku4xpTSNBGzYxyvMHMyihORPdVEWF+Ownp7bSRFwWVhM71twI3AyK
yflfPf1JxaZff0LLsQtlXGdl+w0a6Dkb+bbqdnfnKZy0lYPDn6Xf1auZsh+2IA6CQ9VtGioq8I4z
ohUb0tR1YUUuaPZ447edw/1AA/C0TjyGF08pgF58YIT7ZdYrFOXUcx/oIthz/+6PW6Iiw82HH2DB
e2Gr4Eb0MJ9duAlGyMB7YcWqK5S32QXkqvGs07tiylmM9tJCoYMwu+HMiEvSkY5yVPx79T7D5RPu
su0qs4CLolZrw3gPjp0otOKFdriKdhzjTtVrniPlroVip9iUVs6xixkYXV8Zu0F7xHI3Mnj+9J4V
eQ+udWHaoYbzP9GTnCXNZ2WJ5cgkby8xK8EA7nPZVV17Eh7pL0tQG/0XmPhoCe5MDchAI7wR893O
qKwRjSADLW6qbEP8wzdOm+0fQlHIvOPc2i/zg+/fjtMmFDko1O86ZUwlp0oWTQMT6y2HcYwfwdf9
ppribri2rbeMr5ZuGvxno3uJ0vWa8h5MgQnizqZwX4A4vkAYty/e1+wrO6Ux4priSG/DIGzHBFQ7
34XWofsOvpV3/M0atbaw8My5XSMvdA75fHPs/R9GaneVNJMykoz/HDjgQRqWwXCJDGga8rDt3Q9y
eU3uW33j8GAGqaxl3Er2u4qIhC33p9IKp2TkK0Ky4rQ7XbcrY279U1HLmlWd4mXDfcJ3GJBb7D5H
rQ5XJULww7CstxySWcWRTSgfnzQgHq0WZ/o21xldiKHB66niAjJuBMxLGI9c6uiHzcvb8bT5Sxl2
DRY7xTYBlJZusVEEQPAbZI3bA52W6DkcOKJgU/KX1VSJKriAPm0dfFPrumhYthrnW2ap9t6heOjt
WRKWbHBty/daZURVTMDKU3AhtZ2N2l4ntRXKF3ZqZys+NVACon1Xdsd+Kab00OxeVDSI7QOFNJWt
3qz8TaTlCLcGTUiZ4cTkOn3FyIS3bbgE7FT8v1HIwNfcjqSMW674iVf5jhf+j6c5mYKC+3zh7VjY
SZ8bYHOWXGp658GRSnb97Io3Sc/2x6NvWLpVpUIydYTznhIUOZKDtuoAOaYQwfQG1OcAXhKOGhW+
vm/9f4+A8U/b+6eFKmbEyAoirMuKrhxa/26AR48bCgvsrbJG1+k9gTWU6S29q5x9YS2xr6YNHTkW
hu8IVV5XB7Nh88mpeEDv0wSENurX+Hj6Stm2UtnIgSFM33Xzce4rdNKs+2+IJGIsLsAHzYYoT4qi
LdqlGYgAFyB5ya01Wij/lMpjnVthpWnZA+hz6j0OQZP1j+uX9sIJ9ON+n6nwGK4x3T/CswalLxsa
NMXRhSk1AwTFe5aq9HeFLteTXSmQYsedOeKorK1Sud0/z2Yf5XPiQ9BJhsYXLa7a3jdQdLSzqS8k
rw64EfuUZjfghcphRWYURvoNcISOuUi5Qrtga6VTKuFY0Ii3yHBkAwJrE/wjGgPg6YrXcBkFWQd3
5+homMKI757qrYIRe+a0Xu/rnkIYVMgxNI+foP3wYeLU5SQheRRSY5BTayCKCezxSxWwBUVpiOYr
W/rySb5/1dRDkRnQ4nLH7xgsoUJwneW0vsa2NHkMLFddABLwRwbded28brPssvJepweviB9nUlj3
VCBJSmkLwi7HhJMUlrOCJbYqbpZY7ZSSnJJcupAFmhEd0yo62Vu8DzcZMtlCkmELfAw4HCTX1NiJ
c1/7uc8ZbTr8rL6QcBmxTUHzaVOQNK8tPIqZp+pYRESKnKDM4IvsmMsd/Vf04odu78ldILMzr+m2
IFVsmXuQlKxpZG2lfo9uV1xdMJ1JI5TqoU+osyc+kfqfeWfpOBrrr4DBFPO3kPGGHIPqj6di03HC
be0RO8MjcAp3H51+PIOGkI0QTb8uskROJoVLZvrLefJzWc8iudbQW7Q2PFF6+MFBfcr1CksuT/MQ
os1/Grk5K8QTr4MzaY9uE7yUfWzbQF8W8Q27FJiBqPpDzvV5dimWpXq6qkzSTVHbC9CHEoqxjLhE
fQ3DgxJ9Y5wa0XxN+v7e++HeSEhydTWa4OmIzqPfuscsesNWJo9oZRbvc0JLW72rUNn2OPLvG44C
CsFXJTyXHxO9j/wiyoP9rh9oc+KxiwDweyYS36sfb6ckjg2IRH/939Qv9OeqBEDBTCTFaZO3tIkL
MjJ78Or5vQDnSv68K5fP+72kBrY1hfaz3ZM8gkkXWXBJEj6t0yBV4rCR/C/C9MwzJQHbjsv/6FLE
l0OVvc3gDzd/LmdWAnTWwHY87Z2riCX0KYmdZiLzMrzirw49/63uNrd6cdYSH2gfu6UmrzdQsvR/
+ySiN/757Yztu3aGLaGPxw9ZKBLBHVpd6N2UegcNKlJdAW3FXtlfgMIGwykHIJjLUsOPOR4SZnmH
nS9K8K1EJbQoLK5S0LGueYWUR11h+6vKhw12qhFIG4PPqVkJbK8pipbM7pqXUUp5YVmoHNuuBOCm
a7iDvRzKm/PPxFOuTsd9uso5zyotMbA8vKONBjJY1R9eqoIKx3lKefYXcG0BKcYwoo1YDbyI+zhb
9zPcEQI2cwPJRu61hjvTtcY80tRh/9HScpFt0tR1SuDELBOgPSZ+K0kIEmUXru0h6gCJ8WpdwCgL
vBRWnypBo4WNf6ka2AZEWwi5g0FuO9Ira4sYBDdv8xJgKIb1m+J4skiYqS54Y5dq7s5T9GzpK2DR
suA/x6CjA0gZC9xL/IyKwlYz2AV32uXKYp9gVw4oS9uHbBfrkXVCiEIfy1hcoghejjcKtkQs2sV/
KDZdglsjzsWsc+yrFoXMBlXWeBP8dtgPC5WTj4DLXBS6XPl2ix6RyUtDsTQBtzr7MwpihK+3H8Tf
0uaPgo/xB9aIb55mG1+q7m0WTYtC+SgJ/K+iei75J0ToPLgNNQqw0wOaT0pNXr9B9drVxt6en3M/
5RKJOnQEduFbpHlQJ7m+CzqheC19dHOgphomFgouPVsiTIce7XYMzB8FiyA4nzEDD2MnEkv5C+Hn
yJ+oLvSN/H/LVK4kzHmf1TDl03h1aDa1OSaDN4dfOaTrGhT8itoonrzK76NLSqa3OsxQxeOZ+9cq
SKYARjg5pm5lslOSVCfGY5wt0zP1e9OZ/AUDKchsjyeloQ5rtxajgJ2jws4DwPNaLyVRIo3iRHrE
w51vAe6z41EJ+8S/BINttNc6keT7YtAiK99WVDcS8mNFJnUT4ZzDLJY6Cc8L8Unh7+crYUBXP9z0
qjcBnuErNFG0Hu0d6ODnxfWNB5P8U8mTW0CvQ89ZI+RWB3ov9YTYTKeeuTcOGihehk2bJAzXqYsZ
Oz20S6WoCRdoWgJfAtsceblp+Kst164CY/pSk/WWsua2ApvRkKCVjBJk8le+oD/B25jQRalP+952
pKRWp7n/qQdmwnnHmmz7QsvvqlaGUjbTnEhyRs1hdE9nRPwS8N8eV8bm03Pyb9thAOFGMATLAP3C
650USoB4Gg5iAzvBDBi4hs8REi+PBkXPy026HEX8Emiv0ySiv5HPO8eubV29e98nzxC4QuW+HpZ+
KBS3wAlV6tWOM+It+g0+8sZfi1ibLwWmuMt0WH52jELni/r51RK5JaHTVYyrYtSWvRTZ8mA6PccC
xNwf5K3u6aOrQ8Tc5f+fpi7IEoEB/PPQktAlNpWGnVO8oxnYu5xRoIQmhQbmK+hEdxKL0o22NOKE
UzfRKvZkOxLzJd11MLYQfJaxAVr2EepKJ75/swnS34vOl0pX3YWk4aROYUt17vcNzXMGywOLz5e/
j3rp4BApxW4dsRDtVtiI5WHZRsJvZBYLWhkqvZwIOeEx3AWjCITNtMwwxcgZtVqiG3830ubt2Mn2
HIsG1wZBF2H2YCbPwnaAUEZncjSQ4yAT99HLLV0UewqzTCSNdIqEk5qz45L1EpR1ZDngjibHtcQR
MJ9hx3LLU+6YXsRw6H1a2Qp7tRJO8K1dZtDNRQ/OzjlMR+sUtHQTER1hZ8Es9+ht1qic8Fd3rLZ4
4eNddI2DbmFZcwF/qypu4g6hniy6crJbF9xlKXK1FdwDVmgmc6hZcP5tU/YNNiMEiUS6lGwazyff
5Rgo/bndcpOYAV1F/hJfE0qURMpVaSgHtrf4qkc8nehvtfm3pzVDG3hKD+BXfl3BK1PB3eZotFoo
0IXvaIWp56u3zLvudbz80yyq0gnb8fYe5JtggDTpb/RHwn6a438OpzAjlnWw2s4I/hablcIzGfhb
l81kE/UF6nAkQwz0wLK18/ROKsBuaWxQ4VfgNgxFiG7awpwbG5xgEu5JuYNS6aFi98G/fVMFm7g2
Bf03gSSTBG6nQHRkY6TSPIvqKN8Cl3Pk0f6MeQY4pJ24pYo2+R34CLjTk54CXkhHIVmIVMIiZcCm
sC2v65edWs/wYo4Ahq3zxfLGZalC8FtyDEH8mrmFU5FH7aIyXenWqGfVqjY4N80lyHrDSW9GElIR
XnoXG+3qtWPkOB3EETF59A7XkH0xjnQZELp7/qmo016UkXJwOgkyxoHIFMjq882Y7oTxToosutWP
SA0pYsjQTplBd+uhlzaDJA4OxqPKavc47souyy/T/5kdSLUnxGKX7m3pd7geqZVoAla5Nb3rCeuA
ekwSk+Ron+CZsWuIULtophgtigAy9d+zzARVGu4gqHkh1eDYJNK4iyimK2zfxbwRx8eiH+SUC5i9
FObTB7eRGk4Jx1EJpjeIjiPf8+YqAHmyDnK729MZodb72ca1LOwCwF83QaoW9Nx1tAJwMQGqlxxb
0FKVILhA1ocjHQeN9aHcS3BiIypAJJiu8N26CV4O6Qpb/0ztxH+Uot6C1ENN1dCILQw6UJSAqIFd
Yc0rHmrc/cZsSyKzXdLLaIjrjjbXPCp8MGmkOt8RrVWHveXvvDxpuGV+P2kVqxlV320+w5h5hII4
StLdzsX1PhSjpsp51a9+J1NMxMdp4nDLLjApTDZ/mjvuqrUH8YtudEeYeylFIr/0Az6Ck7B4ZlDZ
nDcmkove6BV032T0L3kzouVGFGTd72ST1PNiEJ9Kg2Sawo1QXxP5ftpnqxX9PJcbl/UGcZtr83ZM
lfKPFFNcZj9YiaBDz4AwQd1vK/ORnS3c7c/d6311K6+vwYXg+ZwY7KbEJV7RoOAQOicQH3tbsOKe
tIPeCgzFGS88YCpgdsxg3BhLwxaJ5cog5SN/afS+Vg98vEBn+03pOK5S7pTY0nwVgPokiXv8ulFa
ebJKVMabU03ezHtrfZAhnzDsuyOBsA0oNP4DcJlV8RiJw2WeNInoY4XeGPgyKZhMKRvNBzrT2foQ
NQe+cadfZKRYSsZc/1hhDZiLwlHkxBf9kCHst2nkbn7oBR252A61ouCDAXGa0EkeiYU3TwD0L89U
E5fBrJ3liCfEkW3966V6I81y6gos9yIKlGDs83Kx1zWKJh4favBnItPwQIkaFWfna1hYlsIBlG60
ItrPhJxs5mmdE3JF2xkMkTiqhcWUfnQCxEqQdYLHXy1Alt1dE5M97tZsuoLl3rCELPOaDm8IbVC2
NHCmf7RPCrtOa7Ked14dn3fG529QQzpwaWTnM+mmnscQ3ksBZzSs99sY8jEgRcUgQLH5n5oJYOHr
TmQW+wymG9aaORmt3sQXziyMvU+JpB7wG/Zh9QZlYRVab29NWO6eIX4iV42z8YPe579RRojUFZsQ
PjgLtXDlhlhc5qMCjejvzmD8vTHcnP9E+Cf9I0ktl/qzdD9pBkUidm7pKz/KLxvboTycGh5KTaw9
3TOzOHoR7Vm09AccmljN7elfQJOyDPuE+5vcO1Jn4b0ZWAGWAYPlpt7y1YjO933IdCLH0zgdHMXL
H30lwcb2vToPHeKy2zn5Awj5Cgxo0uPSkKoFyCKPoIb31o4EYKcalp53nNaD7NEHt6QJZ5ocZSQl
uImWQGyZkwclVnIkCdl59+TUNc3KFba1/sNybyFID3n3ctNcf9AH6heGHh55W51Kh/ue+Vm0jQ5B
suBZ7ljto+EUx25v0a7gilapokxbZ3SIlL0QVtnOAVZ9DOl+5YOh9apwK592YMJxcHfnjzSgKsqY
OuY8oab7U+VRzMfoV358vdkY3eqn5oPeXZbBoOwRDIAHm9EqD1+YW3Xt98LfJw9lFoyLDNmWM28T
EqtCh0E6VBTVS3gt+g6BMZ7jVpXWIL1fE314s2ZP/2gk+gfit+yDl77Dwb/HmookgBuy3NJkeL5X
pucrrjC3Hg9aYO47+kJV5pxVVefPdefNSr7z3Png1ryIAefGcc2Jg+YBOtJ7D7HgW3N2lGYZ5QUq
hi3OntFFr3H906pbpU8Yq6uqfaXGvS6+/YTNwNbZP0LQw2BlUXRB4oQuJGo8VKiPjKQUW9VWNrwS
gYu8IHouddc9nJc+Y4FB7sdtnEBXgl7RoTFYS9B2dbptKwPOL84E0srZeQHTTAJOa3jmwKMWFucR
Kd/lRWXdsKYKXS3hmD9ern3uVzh9bbOldHLKRT5Fv8GUfiDB0X8FWLo194vjmNtqlu1ogt9K21z2
NsYXDE6A3yJ0ryIx20Ckew6uaAcD3ToN/866PIHPqcEBPcsiACCRxd6C1spRpVlrHYNYibDbXNAv
NYvkL2b6KUEQ8M3ZqNhfZxFfNysRBSoqYYZsBWnbCh29r5dM/+UX3zdfOmBK0rZCdY/8hO+SGehD
Q13aEVRdE998Y3qYVT9YYxPgfAglpPt61zL8pEonOteSpUZkMM9fzs+4KODhHMkP/5JBBioxohlS
9AjM9hQxwGGfyUMGLk4Psde8bZaUVdeYhrv3us3Sxnc7vT7iSyGqvJmXD7eQ5CtIxsHesKxzdKnd
6RuRFO5AEOEdBXTWsdejX1kWcGwz9jFmmjzA3J3epkYTQ9WhCfA2FWp8cKiB1iGDjkQ0xfnHdTFp
icG7qMzx84UPXWOASxr6/4AuIB9nymDKb4crv0Vl59/05maHFvy2naGsXDmjekl/SfbYf99uB2RR
j7ISGzkyIsnHwFXfKa6WgRYxCcbJX9kR3yWC/Y0DehyHS2N6CwyQT3muLFJs/gNZsxv5Tkh4gYjG
8jo2cRyFj+A/trqqQtPbFOBvs1fNywKdFBYSmOC6+6vqVpoYe1bqmnrl0tSz37fKO1iODqLTkSWH
OE4aOTXeIVtTTXIaPMuP9Pz2f1jObwpaGUgGK8s+uXiUZpWvO7uuf4xy2OjX4NHzvHGBaCMM5WCI
vagZZZnrH1XLeWH4P6Tpv6lfP2yJD//HC6TBqkuLfPMZ8HkxJQoJYpPFHYF0gr2W45ljJiqkZJFZ
Rsc7i2jBILn59eXiAhyPjsY+zJppBDJZ8kEJC/VhkGyoysfORTSHWPE/bCn3WXPjCAIpxrcpTL6u
0nM4JZvlzcBNn3gIxMyGaB/tyq2UXggNVx3GSvV95DMPvW2V8FIuKo+Z93g/jBX4QlU6KSIIdmfo
vvcSG8nKTkNF1/a2hZXAv+LTmgfynUZfmni4znhbkS+/mYexEilEpaxKYyEHGyjYd2AScGjphVYZ
UNtCPovLydLHJz5HdBmwM9PLyPd+K3J4PvY2/X86e1zHUtLT37dju/unOWcsZasqQVND6tEngjKe
RKhzSBT/KnhIbVXNzb8Sp5Fieej8PmK5MfWdo0q+SAt3LRF+0wLkUDMeOnNg7lB01vPyO0+wkcW7
b39OxUuyUoQYQMq2cOHqM7vDkLLodAH6tU3zns6nID7qq/DLCF83lJOQuzm9/2Jb5+QgRgGec0ZK
04aM18K+8nLyfP06nwxMuFpVJ80DPBYctnKQP8jr4sTowlaJYV3jOcv925JowyZcZzaCMS8U3ktK
wH7EgqfOvYrinnK9Wn1S38oJCBxNhbGyqhiHZwZnkjk7Mp8WpAg9yLnNOo8/f3tiG2V75ptofddc
EWNo1rT10ppxFzqeRd+TPslhpQMh0i3Z30vGTxNFMgQA/iK2s/XLf4nv2GLfuEqi0geUfc19MnKM
IG5a8OLCI6H6oTI7xjK7Alp39CrnBziYPHHj6wOWxa8k02UV90cMSG9FTSaTNlc35pTg3cZnmsED
3b2VhJoGt4gRf3QrNmtNcRBiNQo1YtGZcLjdBs1uMaNqgGi0RJQBHoIeSHD3lWC94f3zWQI26pAv
u9n2IBF1CkE7Yo9OLeayn8mih0/n0BEMfLqujS9dkGMqBLsm7wvb7Qlm/8Uj9oruMugdccXuzsCq
oqaVcR0vmAB/nLvChatIVMJeX218u5OEqTiMHaKCiw+d32GHt7mF/X5TYlMHQ/FKArgmzdZBDbYh
XQYmIbVuc/wJ+xa9fvi0ocGKJJZrDxlj3fG/5nywkBpn7HsByDCQKbXqgN366w3Gq4zYzgsXWtQn
xcx+dSlbLftENdtNAY5SfefuuFtve03qu39CpuYMuAhLIKFWXiz5EkmHo2ReXJrRSdO9uwbq+FKA
q3SZorG+J6dlIao9b0QsdgfH7b2BEbxn+OjZ4gTB2XnPuoTtRe9bL00TvU4AA5/MTvpGhS0CZDgZ
zCS2MiwMInklINRFwtYCU3UElmyLwZYpX8cIr7I+6WKy1hZ3HWT5HBmQdx4Mf36fJCDhAtNtj7D1
qox9ve2RM0gAJZ+6NXt9qFKl9ktL/PnKryR8Q2Hcl1TsjLyK7Woi+THAgIwsBAPUekKGXn1bhX0n
5dNKw441Evwk7lQAlqp6D23sd/jPnIVvjMr8cKiKZVoYW0r0kkBwoD1qmJGbpzWPMINjAJng2ZMc
wdi4GbXTCMqv/h1EEEm0ix3vh53FhLiizhN/+5zXQPMLCFBLoTZiiqpadwbTGXSV93vZIJl9P1UX
T5ytrB1wT9SyAohfOR4xIh/m217CuccRJUiGzc2B9ScCqB+Keqoh8u3w27LUAGng0xe1t81gxu1X
6ZcP6fEEuVfiK3Yq2XMqOpLOBNQ6oRBa7Z0xR63rq0coCq5IGzlKWDgdgeYuSXuZ2u+MC4Mh0TWV
exn8UvjwOs+K+CBnoNvir/wBZp0AukURiwS2g2HS0IFTSWTGwj/a9mpUeE6b+P4mMklrtNsTXbqH
+o+jDixU4ixx9ao4hRfrWn5KHx9VkECQC/TRV7vAFoHzTUiR8jqBKv3F4pEl+dA8gLtlhw66gbEO
OoPOFLf6XfCnB/CRpAoCDFgOhq72RWiNTHMXVg3xDGy/+oNBeXP/KE/zO83niYIuzxhDI7JZ2KhE
DApe4tBI88RxVhl3PgRV86ittLzLWZ6miXZRIs3cahF74coQJRqGNlRWNCR8PtzS+gzsJkpMh6Xx
/SHQWtiUzJJSQhEI6Eu+QYWMxvj/6g1R7V0AbK1j0+zZqF6jU6ttduQ61pPQkcnGK2IVUBe9Ci6p
FoWaygBsEoULVwUSlvRsGCSC2Vjbxl9L2fGOC+5pcZR2xQGHO8O1w7nXoScSGm/y83sVr3smO5Ic
Jq2KTHiLw3UvrDUKgswavLGNHpwlVM15/Thtqqac+S9H0Sg1apn6dIwjMewvC1q15f32lZ8pLYHD
+A08BU9EBdEgEHIkrDsic9F1vQ6AF6m7LGx9QNt5sJpWCDH4VobvpUMbWODtkr8V3W7eoPxUrRO8
SaEW9LOAD0nstGwpSeMORe4AVYo8ndAve9tzhMNJG7xS7sX3A0OrjgIQ1Cw+EmtSLSEVFHvwVcwI
Te65FEq4S0JtpvwLlflFmO7pwYbFdugaaqgPF/1/VtJMrWHu2bkKDoX3dA1kVSn+Xg93ziw0tx3i
d7AOtUSHJLbFuDJjQnVxDLUv2llkk/xG9WHn0XzWTJs1X8N1sBrxP+Vd4J2Rs5npr9njuMhebSY7
xsl/DQcmLwM19+P0aL/iLjXoJZZZKdwtW8zzD5HY+j7AiMIDYs3PsKXoxPv7OyXOymouCg3ydlf6
/MSAqX+xiy44U7Gn5qUnNNdvmAtbaz1KrHrDjsd8fJ4HqgOelqzp8+kTQdYriS38YOp4DEunOSdB
/SzDKZMOdB925/lYgSgpwbndFvurmkCOMZ3tKE3ObEvyqYT6UPjjqNRa0Mf6UDXKQKOMyvvuqsrw
rtIZOszqkbfJe6QRpRoFcYCM3N1v/QhbymvoDGlXxjSESg+8yqwSFvIv/+vjoqvEZiB5+F+xGSQX
RTNz8/agsanxUHr2sxoroACyLp+e/lRRdrsNmtNL1VXj9bDpD2MPzao7Q+sGWAA8BuVo439gnpxv
ARdsn9Bs8sy+OvQIKIbBXqKipO62HstywxCLl3+8svXIICbKXvlUro8A6AzU7IWHZoVNyL4HONvI
YsZXLkhiJo68k3FLtRcKsbXeIoCnakq1+SgsLodDtWoH3p8I7si8c8B0i4zJGSuwD3bKJ0qXqRv7
iAD4DoJQtmWgB7DBvdh+SYOyambqNQ2GZUbVmj+Cuqt8VPHvjg2+cP/tdwm78UfzLXQQLGIk0Q0J
FrJePxVSXvSYzke1aiQV1kTSsLd86lQtTHJobMJ1w4knW8W+SjbEfK0IM1huha1H3WiPVC55Mbed
aQiMWPyH20JR1XrCYQ+Cvg0P9246jha2g2ef9aqXJRw9Sh1Mv2xX1oJMXb25ry7eijsxcKPnUD/1
kkLsPEx7MlmvOJEtXjs8nSgZxBCUoUmwbJxyHsn9Kt5LFlKfKin9x3GOBBJD73Wv3r8dCpNtBI1r
pFgl8MQpn/iUkCuzRIt4ZH1x9vPfZ6SDQP6XR5sGjo2W+uT2AdM4/eilFZ0Oaz5SKqBdgKl7i7x2
+WF7bcWPGsAIKrtInNaNIBPKhe7dxbphKyeahCVBqeEF6SJpVov9msMxnSaWu37eFzx1+R391tog
EUFmyf/ur/OEy2f00loy5CqB0YazLs5vl7VO6FCgugqZ2Y3SgjYZ1xwD5rcgb+L0Yh+NxuJJncO6
rWiUv6jDOZtRRuuZlpCBUtWjEtfjpEpkQ6/leL9L0ri8yS9gOK8CP8SMvHlUTchpdE/AdXY1rmeL
+1LZMQcX/wOicV7g9zYHenbJO1BJWnqB5uRl76YYeN4BwyjRBo17w1P9lB67o5YpO9TZzvmWzgVK
SjPrjXz291d+TXnzNAYuXu6Pt+xoCOSkGc6dpheNUPRqjkAHZuk4HYKjRlKKftm2mP/oZOe0xxQ9
ppt0J5ubDtAhxk3O2vTbchUcuzlj2yXV4hl+MI0hpcx4K+mWj9cxGvHN1SIxiwQb6U8439DpMT10
o+VozlCcBdg6Car5HoeNDln4Oa5AsgrGq1fBCIW2IvJRuR43vEZhJwjHX2KGUBZ5vF97Z2iFUMx9
sq+3mLwtj/KeXl8Za1CCgPilDc1yGA31EWpdqkNQgEJFc7dokr7RK6X0D737sjWaouWyBfL/wwxg
9rvL6cJozA4WqHk6bT+3DyMHJCtkE24ckIyR4DRrIrKdnkUPxj8C/o2BiZittWQi5XdnrrxgWZuc
WNGcUD7OXqF5ibk7GBcR+8JLgonnf4CXesbTC8qyKqSezU02dsRX2aJBXEs8M5PcYbUoj06F9BG+
EozeJcvXZGhMPVSBLQ2tBCNsV7FKThzBBQUNVCJs21Dhyv7tQaPNCImt3QtoNClhfhQ4fmgG4dZR
NHqRRbK2Bgi+Tl6IRkBnjOalEK2zQokG4VFkVFOyt+BIld/jxRZW1razewLgEfbQW1rZh4msfNg1
sL7fZb0m0hnsUN0dXVhHKbAOqdX/CPt6D0xC951OOc23nscEmGzHHpAAVN/4L6xCQjfsoHN20hF6
jbZeQul5wir+GcoJp0tq8eGuBqNAo0RGmNCTBKKujwg2PngVS5VkR8gd45sDV6RqkLNB1r4ppYaW
osAll+6zxdVCDArBqUtVfygcI2zsO23WnO37t5c/imAKnwER9q2fvJ7Zgz4HLjE1RNxXRvMoG13I
j0nL210K1Gf6Ex15eVvdvGGSl0OAtNge7BNYYp4kdg28Z3u2zv07Z70ixdgvQsHu5R5iML40fVI4
5xqHPG0W4V/WHeZHWo0ytcmhTuNZiq6vT0hOOy/pRE7XAt06ORe+YjCoHNqLB5gPxx4MYUnlnxNM
yF0B0tN+vZBuRqQy5fhYvYJ2EZwG/dGdvgYyiJhcye0Jd9iTXBa5KychycfNkOx5OoigvFbgmPsf
Kiv45XRBYjbcTd9CGyX4vLOzxcK1V+tuPp+VkYApS2LO/Lt2Wz92aTSnBS1HVFHZhtFm4OZhkGkz
LlvVTnFT9JAfkR6t87rMVc7Tiasp0RYLrrdGqJCUW0cByuwDuOdcAkbJ1Nn5F+15XRpAx2Y+EAYG
v9R3RxfiNXlQmWbaqGki6DheSE+T3hs91JEx7x6OiNEZzX+33GklQe6O6sOqL6vL/wMytXrWPMD0
QBCMRcfoBY+lZLro1PyzjuBTJ3Wap3MQBbuRtBJfYWn21JdvTdjSHpTJtgqMekMlNHTLmc4jgxdk
/lpgMzEaJvACYYMYnf90LYbypbBxgJc9w/2fEEs2dP+2WLC84zyPbNUVEo1TZaQcp+2+mwD9d3Qr
Rpy7n7n3AH/B2yU5pQGYqxoE17Dn4C8u3YKTOVBTph0nKfmucSbDE/BTjJflRxXbJnzDd0o23SUl
OZRcPH03sXZE6TOtgJWpv0TUREkRuy12JoCRUK1yRC/soimM1N5hJRcWHtZfVo9tHU8a2mWj5pUG
zpTnIQKc5wpt7b9je5/QEqZPZ4wpswZNvhkIVBYPcBAZ5ZVzR1Og3JmHQMN93kJYsBdRlCnahdAg
7qP2SW07xom1Utj21oUCf+RxCJ3jTP4CG4LZBskhP2U/sLBTKQX/kAXyrgpD0uRwtqqmPe+tPttX
zfBA7euX+MpqtVA+0ZGO/VBft/OQVYTL68yFCsPkqy6fBHhxuN4tnUx87U49m7OngLGv46QdarCU
f6BYjxAx91Hpox7RD/GsCzJUtWqYNjeX23S3bMCKjoiLbPnsqng8m716SKY/bwzhfgvo/YKKjlYn
6X3EvSudUsic8ofUh2MkJD2GCzACuAHNH/VG6UMDv7F6aduQrbU9QU+Zbk0+6YUZcyiVzPLTQNiZ
OCweVJL2xj2CllZJoqkzNZUaFdpTv1GNaPb8B/N3L/w1qzXJG9GmFgT18VzkyYA/EaIpF+5deGuo
twQBvVNaitiSyq76M5S0nEoRRKvIVxV188jqnAVySsbM0j4L6ckdD0nfBQwVLJFDsZ58UP9DnuI0
h3cnVKKpKymlDFahT9WVSVA2wxlAm7bezWanGg3+DbtvVlnMuXasE+K6s67jnJ5JJUfONBZ/VOzm
qkkJXAmp1/hVZnp03wp7HGiViEQkHtsfrXG6Lenp1IZR7vfKHF8wHwv8Q4lFBzIeP+ScuXo2JLFX
kKz6QzFSBx6NyME67EQGc0x/nQgqbXPLDcjBY0UQdS05E/tAAg1yPhxbWvRkYiCIllWdGzvWbUVN
1ZJFjR63ukuTIHhKid6GW7DbeVE4t5fHAf0e6sHiBQaPRr5TafqGCqh6Km/hnOOWAKzszeVLZ9P4
MFC+R0TItvVvIH78q3vWeuwPoyKTIwJz48kgaxpK4roiiQsH16HOaD3FgozpPEfwPQtziIk4wxLm
fKR9kVFcr7503OIE0mLZsKQOMmijUUh7wZmv/ZFBV8X7aOuiSLtRQzyhyw6K1h0iI09kYk4MY0t1
d/kGTwpM1j2/WUjIbb+RYBKUAb+JziDKCIhUd/CB2i3E775+pRrhsTPlWkn6aIViCfIOI41oVH/H
0e89Vh+phFiUysHFXgr99jLQZcmV2eQYL4BXj8DoFf4xjtWTTsvGoXcFuyJMZiBQhc2jGyv4lJiw
ThCupKGvPWbuWIcqrwFklQj9h430zm1TWDKCq6dpTytHp9A8WvmYdi1ymZ0TU7rDUreYPAZU+3XJ
HMQYuUgrp9mrVFkWOqg/04a1PzIyxW42osMrZtTbpxqeYhcwq8r7WGi1VXIFP1cbG4B01BPvou9G
J8qwAJsytu2V4QVkT60+xL5SggrpKu2mFDRVCm07qMOTFzbGmCNNSD0X3AMy8nu505r+Jr8hLFYr
o+nLejnuwR0V8PkXR6G4dFcVKj/2+fIV18pP4khB9qLygKLMHLCDUEbho7VF/pveDeHJ8yeBfcyT
WBSYGzmLKG3dXIlOLF3xLUnZvLE0iT0nMY+mXwOqOyV3H2TAE/8Bpi2z+K3Cra+sbXayhbNxO0VS
5I9JEw5tbAFZ5ZwHoZbLl4rwGQ9RsLtjCTBRyCBYMvHFQClMg21/Bnv+nIniH7roMRoNpsBJnuZ1
mJVx/zNCU/VICriKvysVE9fJCVedmKh45Y4uwHLgcQImqlvYuh2uEWhK9iMUjhrJWMC8mdhK4DxB
NVpy4g5f7xdRqkJt7kSbyJPT689QtrC6Upi667lpRrfS0s9eQTewbznHPzXX4Ny9vC6M1fpPQZ9f
h5ppIlq0W4c0OnmB2If3i5vYjMfSvorMXMrFSRZO5Iz4vQ5dRo9kEddmlupFlRz8tBitOQsviQiU
26l7ohE5VavnopWiWQgsnQLAOIaiP7DAPrtb0VtC/w+jdDdOMOymAsdpBIOuUYpkDgHfeGlgKv9z
ivB7xU0cEXnxydyuoxnfctd28P8mrzLoSayCmLbd8j+cb9gtqQ1YJgqIlcOoXidBVYl+wOaeaED+
DUEV0izbWzz0Mh0JW4zVTtySASk5bPTfjyTZsu7xCQTMPQUQUVwjMqku8wNQ+kj1qq6nbwxXRA3d
iJzpZE6Zs60wHQjr9s0Ow8lUM8GSMsPum6JfHB8ADCrmJ2AJKMgvbFBfALq3GhanRHxRxMG4qenT
Vu/wd81PH+W3xMF4sCiy2m96kfObbPVb8RrLjFrYNg6vQ4kTxzVRSV4Aloy86Ntwr/fFCjxbU9kp
vs45reXPOpgHkTLOsHKYCkGOv47HyDfFiHZ8Kr2fSyr2pDPdfJZubtB3Pz736/GDIB7aO+xhNhRt
a6JzWDSx7ZwEjNeG8EDfTpKXHoIRpWKb6IjmVIDgExq7XhnCao48beu18T8GmPNn32Z8SiJnTuEI
bXzTVOXjjBFftaqwqjxOwWfj+vYEZrElJdmJvzku1JcUfhkcmZ4Z7VgPVtuECxVZjC2sI1S4y8Xr
nbxifQNLUg+pS7ON7Lf7J0572uTjJ//N/N7++7X2wI1iI0BSlSnBWKsk/c6jxwbkFZRuUdmiiPWn
tc/BRlpiS7QJTd16uhPGfp/r1IJz33AO/5Qwd0i4bvXbGND4pj+OLw8ur8vQNPNN5oJX6buhSfSj
YGzxC75YjfGIh4e4/xqkD0YY/k7NB654jwxojqHM5wxz6FLaYnCr22mO9aICwz5PfxPUR6S+SopO
4pXbvGDzsg+VEfITLchWxUD4SN6GsgQExtao3hopBYQj0J2s7TqROb2s7vYPqLd5w7aJRKdFOUmP
cOtBt47y+/rE4dmcD9Y4zjWX3lL6e8pQ287YzSYrG7O2+7TS3eaNKhPt8q11M/e00sTGAO9OdFHR
hOuilBaspRvPa/XtD+MLVUAgMEDxiG7M0NGJZumJkGi7JbEXEaE657WWlqEAKcxY/dlzvUNd65xp
9pha0q0KJW76M0rPxyEyRip0LGqwnxECahpapCseystfHWYIHsq6bDpyWhFqUwcjopEQqw7WiKmv
qrisRwhg43viulux4wj7K4Ms0YuMRpoB7FA660AOp7rlCcw17auxgYBb0qOoCsp/LkdI19PLM+Ii
rzYx5IfJWfY0FX9iwEgeXDMcrL0W9JCQ9B+Eq8/j6A6ym7yg2WC60G9ZyyjpsuVHQ6n8FeXxV2xj
9dKTlZ5OMY+PoHDGFCdlLGgxL8sIx9QaV1P8ok9N2T36oe0oFDmySRPN4mN8+wQpHDfpONZqqt+v
3tVynZspQeKfXVltIrxOJHRzP+tG5nX0853pFxJzLm7LlOuA4uanwj+GZhFVscx11KLBvh5UOzpW
FK3vCodJI1w8T20rhmmSKOMSw4SAN0SID4QY+aQJwGIczZogtg1EMzvu0Kx4Tgz75NlbHyDvzr/e
iLkZnZWWMJk2C0VFwyRfk1dQ7GMmQVuXQog2DLm9mlk+84y9JmjglnHBq4ZOBtY3kx+mkXvuXwVJ
lhWLiXRtmNU6J4C4yWgWnP9IDuKGPSql8u/yN36t3OU4B9r24zbTtXqPHS5IPcmPR+yxQnUWuSW0
tD7u4NeBEIGyZucmEOOvBRNMA8FKbC05NIt45RlrC8vXW8af6ifK2HWDrneZIyJOjpw9vHFPJ/mM
QLq/B0gheYCOxNbg0v6KNdN3KzMZU1LvQrtgYhyRSeJ4HIp296g3ghYDj4/SwkWbwMsTYxAUG77z
POl/tWBALSxyQdG3uq87PF849WRpd6x6bGF2pmapwVD5Esq9oMJiV5rvYwPTx64El4qJ3Q8lMkkK
pjzMxPXZSNpn6RGj51mulMMHF0hELoJFvNXPj0w1+WaRxatel28jLfa8DyaJSnFyY0cl0ynhO5IA
sNWB4r+uPiqaxUwAW7IXl6XEWBFVpWKioFI2xLK+6cH55iGW2hDSxphEHQ4Kmgw3GwHsF7Sbqf5V
hbzAbzS8txcN0sjuFN+Z/ibTQpm+pAXakLVSo7T2z7dswGvuW/gWINAgif+laGUlx2HmE9yyM7gP
YQO573YMMx7DvFOWDsvDvss2vA+9hYd1WirmVvgmQWK/9stUy8xTSXWg3YAtRXCudb3uUhRTGYfS
4RETa5GQSAiLtRWSCsO7RWz5mca9KISB9JPF92c3XbH9ZLfDjTvlZdvivnvftmSAiXobzTzo3IDM
q4FAPMfGiLoNTD+3RnRfv/8dCX2wJ9kmfLi1GAJGDtdYtiLWQS9Q0kGRr4i1ix5h5FGieyvXttZj
AIRgFdcv9RuCJwA7osyS15kbuR6Ln4jSqbHJQXJTr63JPCwiv8PNSUm0kXq/Hg9g7VPnLvXE3RzA
7upx0IOOUVY8GQ8cXAgJiyfO8DIMjCrydYsT0aTNiP0SdsyF3WWvCCaZd23UV6/oWLfTJNScfkOy
eke0xumeybUpTiDr4gpfiCtNHVVwqOAjqJF5qtz4vMetd9tgs4q7/OyGrR5YfamX3ODd/py9BbIp
JOVzSi8G0Y78BQwN5JwdbH6lYOcJn+6Be/VsiW5NLriPz+GIr6EkkFMt7tKfctvzjksdUPUPFiXJ
rf1JQx0nhI0VwwebO3LdXBuW8VjNRORE5f0LjfWJps76LWql03Pk6WUtGAM4ZF5u0LxFEfgK8pUr
J0TZaxTc8Li7U2lX4CwdXAVS85Pu/V3CoPpvaj/4XKBKdCIu8MAWGHpsdFy/KFMdefBP/farbnNL
mAfe0rrc1AYfEcernBTb5SD6VPRWFRHvAvuXPqv6pv9EWmF/cI/6lqTL1/QtrK14WPQ4nXm0ukqM
X4pvU9AmotGRAg//ChEHpJZYJumWwtDfZjvSztesKUBCp7aHfhFsrp3DM78Ln6NzkEUCX/E+va/w
MK7oS4EKZG37+nVFPXE3kztVtzBdjPl81ee9f7ePg2q5a0ZWhTLew0O/QMoTQdhivk4AIMZ+5A2z
T10r0FkcAjiaRN2JSwSIS+LSMvj8U3Y5aXPzxytO8I002HK+2s4uRV7rXjTdPdz9ZHAlKkvTzbmV
xQFCWmmrrUJPSTWJCTEhd8C6Objj6jE4wsBEF44dxybRUe+z1sZ5sUwsrHokG+DIta5BKM2VhuxQ
kYh/m5Pb6dOmoDmYdqZ6uQ4d+O9rhXkx+zo+AfaPOdWCIY9R5+/APq7YMjj/oaYskCeZFQ2E57+3
L4Kx+X7lrokLOSoONZd1GlGuN/ykJYn+Bd7KO3FJvk924IWJ97qjZ4xXOxfdU2Z/i3ezx3mJSVU7
59M8Ic8rMzA5YhGGsU9ctNJSwQsIoEsHvyeX8WWqJsK8UIGkTt9YwCReXo0ZZXldcmCwcr/4iaXn
NOCGUrMB7ctLsuExC+W5KMz2naEDTdh4mZmdefT2ECjdeUMBfTeF2rVGQ5D5pfk7MHHjHcUAEFbH
nBwEVgmbsFB2NOy0N4hUU5pW4Xx/SDYZgYIHg33q8cFO9sULog9OulfZ9LfC/pQu21skLM1KS/GP
ylT3cZ3eaMr4pZsruCaqbnNdyCUv+rfkWJkxBW45NKcoqnWpFTaZhhOp+bY+cwjU+ujUOZtSbosC
ZjGPomxqLEa7WW3+oyiH3hIpdoQeqgH2epn1Pd4sHdPST1aoNMBFWqqmbskvrzJdEyl3Owe8TKJi
GQFCRFxNahTJ/2BF2afUgbrwqM7aTrMQCgrYBSPuem5lnulFQxufR5UCw35lObQBxuq1PnSFYu1B
MBPQIvio56Ta4pAEQNbjzRHAfT/MGvWOMvKbXxDDEmx7afCeFf4Ehu1yHYnk8nz5uCP06DGlh46n
Luvqdx9NRUjTjJtZiw6IZR50FOcri0dC99gVFnS1XEP+McmPRV9m6EGM2T75C1xPEf/GQcwzx7lN
8NWIgtjtiBIM6G5BenkUx13Rj+Nj+yCvhGxu//N7RY5t+9uob7XygrysGe0h7VFI+QjyG+7BxgS9
c7PCyMg5WpC8jzmN22PfXn/pEVBc6Mw68jHz9SiXBftkC7Om0CTvd6aJIpRG8E53Xax2KAAJ1RmB
uxMF8zp2TZeXtAoniWcEztmwnwOmacPbRO9g+BOLNhTEZ+q98H9jFftfck7uNNvgK0Bz4y1qRpiM
ytQA5MaF+XYkDyfNPrLRt/nuxB8UvRLiH3/wgz58WqX0UDLoQPR80FoOjpp8OSDxxieqDmgA99r9
ZKZqyQUqjwYweLFU1dagwFm/Pv0jvBArL5qWqgIO1nmbB579KG3WXUk2+YJt65m+Wp80tgAfJ92C
T/eaWOOg3QM6sn0FNCQ0AfXc5ec6kTQRXQ/QGkUPRPx7QDniFH5Bjd1oUWsVVPMQCP4p6bEXLf6A
Slgmn62iGO4Nl8X0QhTEWDHQBrq5czPiCuzfJDbWXJDc7d+rXMM8KnfsBn1YCiKFdsDCJtMuKSwW
jP81J9tp7QYliSVo+TTdGRwj9FTKgdUaEakp4F9IZgdzclsGDtG1mItnO3sJglvp7RtHn6H/Z+n7
oqr6MQlJCjZur7J7tV0iOyN9QMQi77wKEIIufgpAU20sEuco/djJaR/YMxyQDCJpH7UBWpDTKFol
rDimXigoegHDc3fWX6ukuv9UyzcgfPuTrQ0iTna46ktpvlmOUyW6cqfnK/luyo4tUyHYdQB2AcAA
aZy9CCw84rCIlSa8U4GN+Wz5SPm3uTt3Sy0lmrI2k5+5AXQ2J7PO/CfoY+IVI8yQN6n5/X8guOpe
0IE6X8/h5It+ZIG7UYAjgr9wGlkbfMSENYm4+pptygQYZRDggbtT0pmyfSpQbqGAN4Fr5a/QdDY4
Gf7KwZiV33sgsSKvoLHfqvQ6Gcb8ipCxx7Mser/GutLLwNhZPgSejmrbTWahzsdt23M//RD5f+74
6q6UumG5qp5npeWnPUgve0aMvposL8R+qJyyPm3K7imlfX6QtIpL2re7u6rUFvXrYXj6QVdfQBjm
OuJcJDuGH1fS4CxT5p7uo43PifCSYufNf9CGCPXxKusKg+GrvSXiX0+d0GsxGY9xCOyTx7vOsncV
ANubKAvSDGWksjlZdJo1OEq+6r911dw6PfjJJ7w43Jr3CQL0JGmX3qe4C0qhp7kZ+mPuFwLDKcUH
MkrOP11SbdJlKtQRsE1f2k5u47+qhUD1ySqpBpX35oxVht2r9uPaemBnj0sOBXA3b0XWXzsp6f5Y
E38tEtp+xNJL6+sMvuSafRN3ijioF2UysqVCOEb4OZgry4/bymiWDkwBT4YRML5lFmrRvTw8y9rV
u1bAJYwk5BkQN1+rvQBKfLkkEJbVQ0c/wQIMZ2vGlQ/qr4n3Dn9i5vxxF+ZFtzkdBknPlQGmRSV9
mgu2lfhHgEoJyRcG8xvLGCWfBUhxenwZdqPBi2QJQPVQOVYU3DkmOK/Q8R4ICHNH2EckG2ZIUKQn
J/BlaFXAhSgHdKfTNDQlPARvhSc3r+ysMaDRuWMouC7rcbkCYzDnWb9FShBMUs/E3GTAQTzAeN4w
beaOz0rrJkaPwMkYXGLwGms1krZuqFD9uyHYb8kt1VKel8h5SXJwca0ia9zepI0ngSQMA9Yjajbv
sNAgZAFvzKYoACfgvWQQhOdcYt2ebj3Q2CVTi+r9P/W3J9MDI3wtwxlQXB0cvoVBrPLNVgPF1eeb
ZHmLaqQ/dupnotIMDH+Nwrmo7Ikn9hWoUvPPIpCRQBbq/d4DgjLbc+3SUN1SbC3OWdDaU6V6dY0s
33P3Zg2ZBiQ8szZpOF4Gl0j2SoqyfIS8bzNvEusFQzItngD50GQpsw9pR98mP+NFSejdNhywpQNa
Tv7RIE9yi4i67kZjFHWWUGemsN9RXMatby1o6ZKsbaMLn/tiAk2JgOGGpLg9uzhQH+Rd+3d1X0S1
/73QTrKuLIQGGiqAslXDpFbyjOYA8uM4PNr9tMtt24neEPz6ZTKHDaLHXWp86ZmuZ19Knp0/tM+w
JzzXO2iOls3sD+R9Y94xArIZTGz3mmgPu63cTpz8k2WpLVOfHmF57ZcG9Y7lMuDToKUKPx2Ib8MH
dLe1jQ1K8gNJiYwta/22tQtpZI9wlEoN1gtls8IMl4M+vgWdJWE5E/57/El7YztgMaa+J0Sl+p7G
UkTiZeLXVPeMD+REr8RM+GY7VtAraXMzdnr2CXOl5v84TGT3XAaqB7g3BsK42y1KFtS1Sd8UjsvH
sHPrqRVonKl7ZXzdp7wuXagJ0fV6oP2S/fjTmR3P+EyFHPs4KKss4qWjb8PBJ5CeIqg015u2Hgs8
SxmLWSqp5a1BhsplUABysvF3sxtymMy9EZ3iPLvqJy4/CpQ9bO1liuHINfCL0QL+TynAkHqQ61Un
MCQ1UkWOaWiDqFqy4/TfAKJp3WTW96YNk8z1TBBuWATggsB8YN2e0o4eUJhotjuNUs3cSx0hfhxA
+sF4NawCCD4Ac4HceuZ6lS5cKUoWbpX/uGQjDOxOxhJe27U3EpFiqO/ICKjFBgwy2N53aXkiIPB3
KkUlw0fPfrtza6tk2KaIQ4b807cu0Udk/t5TTi1nAzn8WsRzwRoDKwBUI1S89xqDQ6vdXA3/ScFv
5aquqCWTLu6NIvWkCbwN2fGo/bqawEh9cJaZz7uWd2YI8pPYrdB6TiUe04tc944uoAmNExeZFq3z
fU4gIif5PUoSdoVAOcIP5V/ZN8WsLJ4IdqH4M47c0EkKL5n18Os+6j4PARMKpQgQQ+igvyZNSXwo
PEIQN8xlmG21myPWuO6Sfn7MkWVlyQGbmA+1ZHZLixuBf+R8kTEUiZF89yJ59xTQKLBI1hfeWBkl
XHIGPyU155UmdMeaP9PgzR0rIFZI2li4OrXd/vY4D9oZkbUMXWG4E8noX9nAB6qwsio+sv7F8OUD
mTFxJax2UrfLatTQvAh6SPc9QP3GB7Wg+PKHPkVE6VVPEbe78cmvfNS7h0DB8kzJ+XI9Ipv6umJX
At1mOyJzKH4P4nLSMLGACBZ2MxjJSXn1r/NaDcJdMsYCC6vR5J/BxI/IGg7TrUqHV6QBuUS3D88A
rFNNnmHBzkWpQLHncGnfWyZ1fb1UNCWBRgQgGp4ww91XRM/dAP68SGMZIoSP0CV52oUxrPrt+H2F
2GdH9xOLXr9k4pNui+ofxRe3csL2OIEGFYf+IiRNAvrrkIZUE+sYdA1HHssTrp1zsp5rbLFzggDo
uFlGjj+yI0mNn8ymDefffbMrcDn++elaoHAmk5uwMUEeSK+ZTRufZC4jQ3F5htuMeL2y+DqBnwwn
2cY/ALbW6GpXe+H/Gb+eekK1QF589jGcImqrvfH3W3/g1t4Njhfzh+UJ4CMJ3jtPEgm+6hN/G9mH
MOAZtyiX+y+ySTT2TH3sNAg8Gho8SKQ8FbiHKXbb/3H8rwT7LQblkyocaDwkMSTLmZbtsldRROLg
xMesuRyZy64UnksWAxBZzEEPLIlh/8FuUcShDMerLmiEwt/Ghb3nHX3KMZTKner10ZbgHx0OgjWa
wGyyIOMh7XcctzFTv5Yl0UxJfZebSWO3vqrUUY4j+WZ3vfLdfohPKnakQUXA+rBQTVEhURsZY987
RJfCxRLEAbaDmleJv5V8ruc/zTtMXM9DPtpzjs4ppItuTwyZS+LAqIxktWgI6E3uRh2mei3bzztR
SDARhYJlpyKFek7F8s8AHS5uzLAVb7n6GltVng0MsoIV7SOw5bnu4OTa411tqLj0zhZZ2Ttzx+ce
yb2/ghINhOMxjcvcZehRaoEIr+3zFlhJAyttgBpLX1l9hwJGVTykD2ri0rmvcq1d+NOmJorGRN6A
WKphIX0b+2wb7//QD4Rpr4mZ8JNG75bnA7XiOgQSidVpZgiHXFnEee4KWczaTnEbyPYQIUN3hMRm
5yZXeE6jjQiXJnJGtF5kObDztu0S0XM2T2O81SvWZww8ZSsGgcFddN4/oZ3qJqsnHcdCy2oKMsHe
sqNt8aVRZgGPcr9BdM6bzZ7RFYZ5W0xcGwyPDDF2A2HwYhxkq7Are375CUudLnLJS4/AiW22NIM0
fhuzxv9E8aatthG3jmw5kXH5g/tHZ61bTX2DrAa4lHNrPjUdC/Lkv/1dpflEhSt2l09tW5WBV9bu
Szt+ucUeh8qbt8WmXFK6ON+bsXvEuPG3vN2QW67j9kePGfWUn/x1OX9okZm5VGH1oLrQ6limfQXo
ePbR+PCkkB8kzPR0XlG6E7UY11F00KBNgRtRehLkLPPPNh+s/J1db33Hr1Q3WdRvgx2Eq6M/Tyuz
gkb0Pkx5/EgmmHaqo8aTNppRGPxYtlvpNgZqmjT0W0esN1r4rLbiQt9z0b5LUKL8ASDvxhU0945d
0lz3OqwGemsEy6c38mZ9QfalUuacjJ6fR57i7i+Sea9iw0IEUUIRKyte+mKr4QsvFAwIwHB98IuI
gzt5CsYO6Kid9c/VSmA8rVu4xp93EeP+/W6UdTFKFuYpwZ44bP2rHfALPVYfeWRlfz+u9jZOQz6I
9okYKelL169aTEXA+F+dCJ6s2wW9yG+ia0NkK2+6rWjIY5LRrsckqM9kI2Ne4bvQO9Jl1xQmdD29
9vI301HjdyAtOCoDL4B9KqHy4AgxvyDhM+FUIQqBwYZw9Fq52DdlFGOx4rkqLikeLFNTrL2VuisC
ikNeu2nB99h9Yt1VNpm7jO+norcPTQtGGjuSqiGKnLXK/Dhy2Volpf6oh/shXN9n39+cDMOy60K6
ZPgnkePfv024dWJ9nh86aq/x/2EFCgOg/Hl5R2/OiAgH8h0MiHztQ9kTIvtWlcQtRtMWnNjgxYn0
GsqP4UaV9YJK8RtE64eUvHpklX+u+fBRCdceWTasxsVRdgkgi7g0iU7DqKxpVM0JNIYmjz7qbP4F
1cRAscjNQ/NMJ8sD98g71dRUIcAoQ4PXMX20kecK+qUzEoZM5NSck8WYo3TyT8uzGTmlFMaeWEkZ
uCWbWzE6M+gVrb7dHZRdS5jvdDhrOMkANkc1nRjE/WwxgeWUUgbL1B8sUqJK2SDQMsIK0MHcPK5R
Dxm5cd95xFxPfDzogcKl7nPNJval+KBP1dNgubBkQ64DKbHUWVEb98jkKuYO//SXHUt9V0TQH+nz
VCpSyTgU+9l6V4pvrTcsrWRasenWRYoIaEAkZBVxlB9uTlflN2XuSqoOj6QASP+T0m6/SPlS5VWX
N46MMvTdP+NUlgePOqB6smhtFA+zSlw1pbXwVPkVxS0Hao37AqABgDBbp6bMM3VyS9//aSacQWTC
Bhc67wMjjOS3j/USVJIuHMzfM0vBRP6FaeQusVaZ3W4pCQxPY3KdQR28yqWk+5vme7N/+5+rmtft
rkB7R/j3gMZ0V0qSY6yH4WCStGjV69hGUjCvZaB+Aazs5UNvHcb/2V2FJAKeplbhd24EdSfpi8Fq
E1IvemWsqsFYrJBt2WdeonKUlDHqgK1mdt/emEFRYfupM6N7qT4Y3UxTUB4WJZ7lm1tDWi5EAlQr
Yb8SxUrJSCa9XAnLPiSgdNc/WCu7bIcZHCGw4ciN/EoeU5yqWtHHV8iOvSAz+1HpEjWi8BEmrzD4
gVNSGoxW2X3Cw/hcnMjenKAwzuOX/NQPdBDkisuHgEUZASaJHDhIoIpwjd/2Z2s1BR4f9akQDeZL
LQFZpXjkXyS6C6Ayr5w2xPwKRledu6JsQKuqPQvvafiX2P2VokicPehTLfcy5uRTncTC00UpJyHf
ek59uYDq7ajnP9m2RTuDi0e19Jg0HHomehGHpNnI1bvYxDNdotalHcoNhiGiuWgyIJyq2UX4lQ/3
GyzVBXFgz1QLKtxDUtTg4x0ZEcfS88lfpuk3poFr/o8gIUGm+/3e4rb8fFyLF7E8qd21I5IXexX9
IACwSVcZa8efsPlpgDe5n6k9+V6+I09S8lPTkG/8urncfSCOvddhbdXqHjFHwzxWMhnsmkARKhn6
AHs3ybMEOj049xq9MC7alsvLzdXtQkA8ExWZO7vN5CvUEMG/VLdzU/fRYt8D/g92OlaY1xZ82IZ+
zHsTvRbn9EEAOUynQzVKgQeRRfyg49P3mYB7isK3ykcX3E5ESb5bMsEHvJNxIe638nPej8UXKYlw
HMADUV7Zo5lSQ99CJDSxE2/ETEd37SDsr/5Mhijc+ICW9IY4q+5GkVxkTZAQNmS7mMSsnPcA2s8c
bOFkYK3F9xTjgPq87Ql735tXc9Fh5FJOBRjA+Lwm7U86kjvAjhzMpn3ETvObnmQyploDa5Ey0ma+
gh8+L+i/lmj+G0AVHTHJQUbzQO2kS0h03WA6Y58DnZ75iwyiPlVMPePeC8luCwabhEKLZVwdKvJQ
zLndIyrO2ktFQ+Ew7lMrxMGf4BL5QPxirj4d59wj116VHi/Ds4bJj3O56I/mGG7R1tg2CpyNpqxu
/jKiy4TD4szeusmltc+Cjdl6jn31O7MRYPiivDzTngeg67UjIuvidq9Dt4a8d9Kd/80e5V+HaaFu
YDE5LZtRWmmSy5hZhMkun7BQadiDHNrFeAqrxRF3rECRPEv7Fk/Cdtk3KzBhvu6aLmXJl+/wjL8B
dnqCKSOSd9XCuTmK9ANpx5OWOW53+LnNMz3Nk1FBJFum5zim3JB5dMGNqNAeTMHdfrDyqoziMudl
+abbKzZaGteRzaNoW7gc5YJrGqwEiDUIKWtdR2e8Ww03vv7k5Xri1wnV5txHEteIu3PLz3Qk3KN/
f1VeNREeaP0v5vdz5++ycaADTiasnHWmxNBnYE06PpXJSWeGkNs0DpFRz868PHD6jjipkbD5pfAa
R1nj40lyMkzZFRODE7q0Jm28V4mGLM9qrnBlAxnNfj6lk5/NruGWzJLx00TCzINJqsgSE/4sXtCo
IxFPvFY3oAEgoHZK0OH8GaB8dLQd9qu2FhQlDb7XtWZk9W+29rUIA/yzRogrWSMZc/FfEdZAOAzH
23rJ8mE1U7DcuOB5J9MYdkK4vS2/0qSgTWcZx3ELd5wrBT0FqHRQrMW62U0FtXRuNVXOF5utKe/e
48xDzwCrIYJ9RCHmGwYVOOi0cRyQ3hgZ5j0DIMxuWEwFbQ17pqD7DPg7xJDX9Mi5vdNqGVznYuMk
/GY0rAzfGonFp+hSwaiVtpdTfnVd5INl78Bc/0ye7lcqHueBjaogtrISaJ43oHG9CEGgFuDOm13I
/QJLemlkmvKECmynfcVTnlSgeM41j2e+dv00q/sw03HX2uvx6C4BEE9bzVdaDvKFajQfjco1W61s
KlO+avYGQJEzGjPkpQqErtf1BSWk9RqeUqA4Zm1QbtKocK4IGGBgemwAlnMduipaNCcmUBhm3ao1
ppXi63FgPbQuLhCNM/yGykNTS1w/joL0Uqf/HT4Nj1Tgv49Q0qOvjrp0lZ3NKUnr93fVhh5LuPZH
gNLwkbe3EpzysGfDRQkly/OYXQCJsXo3965GYBI69JF2ly+X4+b+v/xMi7Tk9Om1gKubkBiwebcF
PX/KsoYE7HK+sIVSnGQzMINh8UwNc/KJUCkuO7vKBXIjeHqgR8XDN+TC70oJzm3Y8v00A0IR7Zq8
XOONEqlJpTxKiF2biWjyeDJ2+2WXmsk3an4y1nmcDVyBhUxgbMuTxx4Hn/NhW9V4njwy0pxIZpX+
hFo0lkDxyS1uOXp9CWRrvxkJs8P41QhLqZ6qJHUTeRLrG2HjblR0IwgxZZTVrENIjq1TVu19m0cZ
kroUOhfZZFLKMhxcC6i6vvmeF58E2AONaKG3mkUBQdr9O2bcOKE8iDmRpatRGuT/h2bZezZPbpLC
RyT2KInYteCrMkO4ia6qFwEcwmo/0FNckKba+SGGDOkYM6f6LdPaNsggoBLtL2oXp7TDVyveP1DV
w8I79hFkSuDg5kpOr/riGwprqvY/nkqP8i1bTZCjBP7UeMSDhyhJYf8Pu5TP5wXtUzDJ8ZsQ6v85
4OQiVfL/vxZLEVoaS0Bw7V7NNkT/tdz6dJeQhlLJ5bCv8aQOu4eJwZFUR7qqQDvZ2gjA53edUXTE
CCmIrMUKqf0qkcmnz7aUz3kuhQQnaI9EFSTDdjJAMG9658H1rWWCzVgVDfib4ap6x+eFA1U+b7o2
NpQ8FUAXEd2cF1eHP0T6XphwCQlcMYNzohU1az6dsSpn+V2IOB8DwbbfYn2Em6N8G8Gx56yOavKV
OeRlT2LoYyIySA9YhlmLc/hoMtv1Lih8iEjsSHAGvG1MIymmSoIvFs9oxzmYrkA8jn+CUg9z6jfb
MNfcBm6uyOO8uVq4SGmfQ9CAR+v7/RWoi2EknQX6zycbcFCpgH9cMGX1vxLeyI1/cX2d41V9TY1T
o0IffdRkzE807XuVV+bGBNFQLBKG+zKAxWIu3U7W8Z6BkpFXyX3FibqD15gsAIhwizc0J0Vk1laZ
7hdG61n+GUy3BhDulwYBHasBeHO1vgYT6AUaJiJYeM2+buCAg5un8qh1HMlJGIggG7MbZo5W2m5N
yykVnJVoHXj8CAagAfyLWTzPLk5Iui7rMBo1Zw20LmE9tpkoRyW2ehqXQ+L4Jw5g5fy/iBpc1Jac
WuCX50CChsBJmFRkMlSk7Ji8g5bhPwJajr3BsvQACR/KroaCEDyXe2p2vugka/dCspZdJrttAB/g
N2iPR78l00HEL47CHESoR+8jpA/a6QucG5cd6q089bpDp35jYRCr0WOgnHy3nhM4678FZYRv9nAR
KWrlLIWlae8MlZQy2GZzBQq8vAHSsk2eeAMy+ibZvz3UDxfAocqly0QM2m64E3DQdu6Km7WXs8xk
YywZJLnUFt8Za4NrzKNj1BmnsMZLTzU0Zs5ZMPArndgyrlyqBJ/Vk9dURe5zbKYmgN8Q3fbKl4eL
KhkOcDYaHLVEfJED2PKpEg3yWa6mYd5l5IdK0ywdtEHY/AlQRkFYHHbQzwYQG+h6cl2vtERm1yCZ
+vKlB2ILFiJ2jHstTSW1IauRV5RlqpcIMMCpZU7xF1qfZaD6ppI3QW+mLZtyywUJfauAbFfbMAIE
sGoSCFlAkaodZgGtzqUZO3+n3n8uHTwEYIb6rOPISvgknyozayE+1X9jPXzwdxXH3tay/eeX3zHl
AyPtToHfY7PdJO149nAQO6qTTqmi1OWV4clzuAT3SrrCl4EI2/yD72u4sBa+gosh1WCKaAC/iT1q
kymRdQrCXdBTN44xin/fLsrU8DZvuUlwTHlhVUj4pkPsRCGdSc+sG2zPV8iCIL9Cscjx5iVWRWYD
zNKBmSoxCCacBwcF3yLvJhUJyoDhomg3iOlxKW0RlZr858kd5hUzmPN2dormjjQIdOTqTKkPwraQ
yakAE0zLQh1QLUGp9+rpq6P3QD7KF9kV91mA7JPs735hz2fV6aWJcy72dmuXX9GZh1fVUcw3N1/e
kof1NIQyG7RZSiLFrYsifs2yqyyCfMTB1gqqsN1njreGDMZ3VU2PClyvva/CyMIrGYo3lJ+flEY8
PmL51tpiM6tqzPPxSdeVXNUk4crrE6EqGigtGwlSObzmw2vNheeR+9Hzh94dVTRsZD0TIUcvWEpS
jrVbH9LKk89D0ZVfuWjdMDSXBr+Xe+bpUuaQZfPn7SRL8wfVw+1mG9HlapqK+qVMN4gr9NexGgpg
nsqxbjlKEsOsL1C4/mLPHZ4z4pzd6Ebnt9uKfco3jt9faC9tiix0yhWjmBun+ukl8QVYRoHKwHuD
UCpSNc2ttQTzKKZ5TdVr0O6jQPcGxYu2+tgPxAVxLEVBkRrNFAcCdZwL8MMwKaSrJsfSDC76Eh4O
zXnvvrjWcfnEpXR3YxG2kQrKbgMxGiXBuBM/q66hy/6wmwMv3/EPq0nngiSPFj2f9QRyZjPjx/Wt
HtziAwUll/3BXPtE9GE5wH8tG3MSfZ6q3bj5p66Vzb0Gv3OtbJlbmfU6MzXZyrO13uXqB7UZ5JLW
6LmjYbjwe/ff2Wrz5X5vvPC0O7lEc5wcDB3CtM+3BIfA4UrD38gzcFJW8pR+hxClahdJipZfKd8l
t/OGKFMV/5p+egn6b0U2UQuvURhoiwEMqlxkzXl51jPPrrzEnZIE1p7Pw3oB1orDxa2w4vellQBd
ypgHb1yi6olUem+vYUJzG0NvVBxCMTNZ0dfOb9cJzOHlIH2QRo/4eFUO0Rm/fwL26SWadnEJLg7T
qpyFNHTsOX6+O9O8p7B8SxGyPaMX2asr62lq6XlfXU+iFZXpKkayejXipoLMSn9tqibVonvUB1sG
CZUpKpeOIWbVMWwHlVhC3RP2PlXMligiyzfpMNWEjPufvFygpfmFcu/usIf05s3K04fwwuxkBh4H
OwjLLi8sd4kT3KW2mbKEc0ZxifujzoWpgjNX4hnIKzycmNCJ4M5dUqWX0VfyZdehOBnZJ9t1SB6S
uNuy6rnZBmPyB7fyqAjKrQiYI3EmPPcTV1YwJM5iNyyJ6N+7+WiF/tUFpSxiUTNwicCVPhydEi4n
UVqMjnGkpVIgRCWABBXKdylSIKvzGZ5R/REnK6dI1WLC06OqGTFH3FSNEli6q1p/GUP7oKcSnUad
38qpHdRzRbBlslL5aQvHu74vSrVfR0uFDQBjxjNbhwrD8jFjt4y3ie/yS28DKp6LLeHQ4KkcBlEN
EgBjIacn43gteZfbBDkwZwhAptzxBN22+Fkw+lg0o/VDu7cQG+OzwsIqo/7XhfAStyGFKEiFq9gF
zN92GasxKsdPRQUeuw1LrKPcKyZf52nDkfn7Xiyd5RnX3XbmvDm6fNhus+Mu5YcKm9Q77bGUr618
AMt8tqgtVfMadJ9jCVELqZWPQBVccdrcY8sJ+JA3M6iTY5+mRFpWp18fX2G+MTuilh7/5YuqKePI
OXNQHUj5sw4xD+ihXKN3QhCN/1/M5Gt8UTmTj2DwShI8o9t763LSBjEsHig+0p0kMIgoS10BOiQ9
1LpgkmSYnz4FXEUASSjGd+KQP6at1UWTYXBEsGMge9h87Owbq9cf+B/QmMfnoWJWcGZU+wC2QIxy
op4xpZuoRaI/lW2FnNc3nYmcThA2aLeVZ74J0HZ4bpS2jyrQbs8bFocNSCy+rvzsNYoTlqTv7T/b
eM8HXkxCO+2J0b3GBmgUCGSSo4yqPAULw/PijJOKwKPjhg7D/9fjFQmN8PiBc5KfEGIKj+KteWaQ
UiuyDeOjodVWMqtH/6iFA7HVy/G9vPH0VpC8OTfyqxxxK6GvFLFdJVI3K4AnajtyNVCVi8EZA1x1
YahFkAZkGUZ2TB5vtVVqPPk1J+jD3h9y/ilsi6iATvBPnaMLuehVG7Ip83DgzOWuTus86blkJWnU
gj3N2UXSaD9Eyfc7IhxSIDCp0jlEbE1ZpgtwkAViRSaDqiA7YXnRp8TB1DhwE8FI0ujYumPPoOxS
yO/0LRatH7x7cTRycNFKvXbGeDFL92uVrqhgcdtA4ZouSU4d2OG/ZoA0Vdo9cxrhcGNNCnPfQYgA
EAVNNQ9ZQMvZSQ8PuJt2DnxQ8sL5zjJ/nFtDRqBO+R80ZPba9riEB6gF3Jf2TA1ZU0+X1dmj/ZtD
zxyl3thCkJgEzMc8DDwsj6HlgpFIoC0aYs12za4g/zcAiQoZJXIkNoHQhdLiyrKTrDCmI6C8Tn4G
Z9OnxCwXf9CYtb65kPNQz4NS87x3MrNFOTxqk9cfBigQQztD8Y/WTnVclfYddn/YD2mTzGDyJCke
jXJ/I0NNk9HahQNtR0nvfL/ndadv1OmkStWyYnGSOgtLnGsCDv72k7m/uCBirc6f0oF2Xm1+ZnS6
4DI0O0wbNHAGGELP6RLWf+8bLCdjcMoFYevJaTj8UvWHWYbM1LXl4B9XL/au18QaP1vTXpF/34i2
rhMD0koFDzfJc68NnGT84vJy68boWUF81GcXq3kaOF+P3rJEc0+9ymjwkqcYDvjoDLY+oyft09IV
NjTATnLEwJUJNILM689KBn5FaLyhRuPgwMD/YtThjJPcv7ObarWc8r3x4QvD4EOysi4wb4Ag6y9y
ELI4KOUY2HWGcFvUdiG1C/Nq2rJL/p2krfrPgveCd+IEAzhlIsC5eVkKG2T03rcNeHXL21GRrqtg
RtbxA0NB8Nk4uLrNuTT1fYHwpZ6nKmIDCvF2ssL/3t82KI7JxatbIL5BbOe1lb10boWRDlpvqvUr
06t2NDaHD4M9gs6mdOVnXAi9rl78btUewfhTkyDp2H6bJQl7GANfOsSbMK3peiTolggnZ+BToX97
T5zfXoxhD/b+icUuZxSLGwTsjUg1YaNYO7C9Cbsr7o3CUs7zKcbNpBzatQMagfgsZTPlDpmuoQuq
qU4U1QZOP5PwMoHEuAoiG5uGtBiyqOSXGWH8FSQjP7nVG8TS5w/dib0OguITQT+XCdySyCRoI8YV
M+s+88MdL878sbvkQWiJxw8rxu+Avg+2CubZp0WGIR87duzZP03koVpCehEpCC+LvRaPtKu5Hc81
1KVnsS3KpZQ2VN+k4XvUgj0gRL+0A/SX0CTYrTcsYgd/W8j1HhrtenWL5/LnqJlQwjp5DEkVTtND
5K65hm0SPiNIh8l1l04uy8L/3BQrReXFZUQtv4duJH08ZGgy7t/GZ5L/nZ+brHJ5iF5bn0+vbcJX
Z765uzckAvu3kVTMQs0cqDIs2MDJq+75lHEfgcQHAlTe2ZjPSQy4ZfKaigfvN5CdkGiohU18za8i
VtiXXHboF/IaYKon53R+jT0vFFkuZCvsRh6FFt0NFQ7YIbrEKOmDwSDx+bQetm5Uq44zVT64to5v
k8Hd7UvxsH86cdMBddD2fkBQanpqRAB/CBcyPsMi81oqi4vr1UcsQZcACCGccjBIkNQQ+qzdYDB9
r68bOZMl9BpKtybRhao8BWfKfvrK7bRwA/XjBXjzihZ9IRiP9ZBOfxLkr0KeNqrvl6eY+OV0JJLP
36JP7K+51wu2fjG0LqyqoRlE8slFitOxD8QOxGZMKQDOsfIpcQKYKI9faDjFWpdJOCOVFefvW5sx
Cixx1JOdfjBLwA6tnLOzTTWKvFLuNqwlgRCiWzrcRpYipSwrXsWkFAsfwUmbo8svq4Y/IAz0tqV6
WUb+5EnjmPVp2SJWeEdPz2gfIQ6peChNBPX9ZR21eX3oSAQB54DO7x/B5WGitFCgBFuZwox+PV84
usfEi0mmgRr9wa5xXjBbPkKkyxnvTr++fxOSLI8Ob2xAZfWpEUqnZG376z0V5zWsiT7f+Im2DR6t
eifigTs8UwUkxWlnyR+/HPw9L0/zZpjCI1yXosl9VkKsoFOYv5tqMM3/Wa/Qf0hGL2yZlgFQ0QYX
NflfXOxHfrujgNXjkLdVmte9/E4TvpyUgMtddX8PxfpYusMB3Nps9RCuvLTJV/2atKY1jd3z1LEU
ELigvo7kje6thcYxmlgeCipx0Uu86LArL/bjsHYGUgy3kRe1PhrdbHUpGdJlUr4n7wbRWI2VcWbu
Ujyvxy0H67brDEfzwo1MNGLCFBwOlaehyQPq2JvSMxUeuolgg2puwRttyQJADknEMz9YfZsJEudE
BQ6onJKBwphitf7m2mGnl0QslGx7QJzCizvDfNgji2REpzsc3Ur9Al7nNVY7HGTr8bLL6zgeVMt0
WoOIRyZZ0voJYNu7p5/9ktUzY5A5qAQyYM0iF55RzwhhH55MhOTBmowVk6YJRk3vnV4G6HHDm4Th
gbMJRswQb596SNzHP1l8VNKiC60t87aca3QF++5nMMqhKeE+65fFxl8JNVa3HmPnySLbwMhpuneO
kwKaX+Qvs9kKl3j+97hv0ZvorfuDDFkDm7VQ/fahbqxkA8BvvMmatNlVu/iTI5S1VORXf6sxzO6O
FThxxX/htOS+gxGVl8o6yN/fcPmlCGQSy2dXSNlPyGtAMbKoxtJ1pktzvUq94gjqnB+h9BTO7weD
3U4NSmnIh/DCPAaCYwce2Iko26kqBJFhAmdgpusAUE5d+TYVTfrVA98wwPdPiIPTtxxGUIT9qpGU
IZNIxglHJwJHoocCTn5JhM1p9JqYqSDvI8yuh2BH/Bfnfc98AZWpc9BII4EfRGeXzKOlxhr3tlh/
+DBPmUdQoUKTm8jRf6FpYaz5Mdb8Q6a4+6yNhJ8u3y++hnvX7x2z+94yQ83DtbiLKCAw+CxVCtGt
XqyWnwUYwQ+Qn3CHahSUZg9atuxHKPTwfspoi+cFOukdgyUv2OEg7EKHAKQhQxy876XBpgMmFs4H
BXEVDjcJRVfok1lJbEtNFzWbZkdB4dtzH/vIpz+CWURMmPlVZxSlD5Xvm+Ds7bP1eR7dtH3cZtQ6
fKH0Rs9IH0fei9YPoPMq5t9ViYNFOHyH2SHSEwdu5V+jw1S2f8i8Sz14k6cecqVtZsf4s7cCaTp+
kVdrsMz0a+SczqQH0k57tnGmX3UBsA/WPF9LIUshgXKDDNUo1Lu1dduUTxpes9FfR4n58nME35Gy
xQjOWj+RCvXqjWRers80xVhrvMf0rYYreJaaoARmOgphxLP0I554YNdEFa2iTIg2DlRy6Wwzcui/
zSs83w/CE9poT+0MevRVCtlP6QpFOL5mpibRqptrzTmENGKPjoIciVNxKedF3N/GFLvlQxBgK735
DemenUX+qhy6OkxOpnOJpuzEw6jM+Xsqs/WdRdu8hrR7k4C956RhBukTZ4zHem/OxC/2xk8YO0Ih
1B8D5fyETnCfMsUZpa693rLzC43gRtDGm2gMfZ3Nyh6LjxjkdkEGlmYS+uLfnMO8Ys6qDWncPnnS
pNN9BVT9cAo1+uoyBT+4jiHyK1TURzjNvUpp0CiTA+fah/Pu5HdNb75BsaVyaCXhMuCMe4sNi2Fk
YRjKZth6yt01LE4UuCR/vhBjmGLfRxsabmJ8C5T/KgbCNBXNTOjJgp8Y4FcQOkW4ihsXInwLLwOd
/NB8VV0ZGB+qHg/o9G7ny8fRTPImKkpbNVkV3zqqvw7tU9SBTM5nH+rr39bpBznhdd911AIa9uKv
c83mHX0UO2k0p/jjHd93D8DKSxHCgMd2ssTwsnuuy4p415w0pe380BkmsjFIEYweE8ClxZYsKUGc
jQkmR0Dcqb8ZwM1SeSdt8gxk8qYFtJ5Z05lbDUkzscxV52D6KgwUY5xay2tvc5Mn+A7jpn6JljPB
V3XWSPspI/OH7sqaJmCi9G3ilzXmbb4gEQhxqpE5s97f4F+RcZJKrIVQMqSoeMWC9BhsPpN3M2x2
26um1LIB5in2ub/TW42bZQa2+fzvgzDAf1FH9UimXZIaN39NCuK+sUPIin3sYrFFJNP0Rmj9D//v
6njhpldFPVrMIpXV4bx3D/Mh/U/HsQHtqxoFyrkxnn68EnNWS1pyKgBFkokZ4k3AoM0Q1D22UapE
pICldYJ5LY7uGRtyq1V4vdevlv2LRf+KMoz9dQXpRJfO3alqvIDh5fzvPxTKT0ztwlsIWHkQQWPb
X1qZ/ZYjYGzrQrVxoGUB0oazhILIUdpocUyD1uvNzII3RuhZlr3xj6tSza9rmJPdgVg0uCAwCjp2
Svi9rcXfF0INqJi5QLTSh2W22Nw18KB0Q3eG815Zf09h52u4rhCB7yyFZVq9u6pOVGNdioo82aIQ
otExZ1TAt9pgLAK7W8W/LTs8b3B/aPCKHWKWH4cgVvIk4Z2ULfEQfVSit3p5uBXaU9veuoDe3vx4
l3j7aVLsj0QqrWt3GUhVEmp8re9AcmngEkPAReQ3io15ElGryPrps4NEJBOtY8pZMcRg0M1dRn5y
R2POR2pjL2BLky4rKsGs6x2xUc++j9L4uPDCkTYjujoaA5qqKQnLBE/cqUkUGFmNiGwm8Bi/BbR8
E20T0m3UgEXzbsHaVfq531slC1xa1DcFQsAZhfM2deBE7quXwjKXEZXgO6sCn2PQlA/hctfeTseG
T8W3SW0bJgOIM4HqrfLpOYXhlbQkJguX0xFbCMf8LP3hg+UIlWCplYif6lHWqmXLDKOx3cZNcvhJ
avhqSMxZW88gTCwdF3CJRZ1I9JmqS/MhIThw9fyy/SP3IPlJMKuYpDGiebUtKYwaqms9bwaBmdpR
ZJQng1yEXmMiwUr8NI+Jv8gjjzpEnSGok0MxSRlVW2P5nRQq5r9rASWkArNN9o4vqESGQ+k5/Prd
xea7ybTiOjlHoxC8QPT55daKm5JX2eTLkCAWitUiktvpvJ1WwZzQk3eq+l7ZJmpnt6+PjBtDOVmm
U6CH4PK5FMRkCC3bR+DfAmc7FmjJREF2VnHY544JFm7Fm7uuttaNupBU8Beld1H8RNEQu5NHIcTc
Tfmr93XoW/Oa2PIxY7jMOrgpHErDkYsM5t98ve9W7omBt4G2Mf5czlB8CIlZ9WWN7h62FSYWgMAI
VD75olzc8QgX5H1U31DGZ8r12fPjH0rLpDwHRVb7gFAZQkh2Xne8VrrUUn5hb21sS0HeBfg1naZy
+QMY6gc4HQIpYxZdmOzrdFBteFtuf0rUU/wVHmD6gGYxP7Z80Bp6lt7KPhPCH+LH1kuEiZ5lO46c
lmY5D9E5mMu/jw/JaHiwQt2peQiIatjJKwd8wGYgIRseNQg2tzTy6cdFPaiyALLggwEGuOvsYt+3
N59kAQNg6Z09x/WC+wIWpTHvjzwyAMfJqD7i2WpzpirJutHuqfyEaNiG+12vj7kJj9DTNTkKcA3d
rPJimWqLfVY51snc4B+HlBdJYlVqEb+9GGinG26k5Sm2zySSdLo3mrZyTuvWIkBv/GPTLc9G8cgF
KV+MaGrXNgfO1s+ITjWs6m1pgSlM8Dq5kfZFi62nZCZF03IeIsO0iOLv93nhl4VxwGuIxktSS4uK
NjHRe+HyepKfY36/2O8Kr7qwYyjXhvmQ3RPSZQK1EJ7ixV6Qe79H/NagXPkGZ4zHwzz3G5qdmnfP
qPUHRKcMqKKVr+GfTnvbc8/jMvoLKbaGVqbkCjFjNGu81CxDhZsleWo1rBT8c99eS0pJ+ZPPu+kj
quWFW+JahJAeeclDUxrXBbwKV+r9Za1Zd0g4LmTGH8XO9xqIowUy3SgJ2DB4ekAS+Bh3gCV3XuwC
qmH6DJ5tvVdog1VnZEY8fPdO7o4uTekiUd1uPg5OlZf550Y7YJxm2qsg2822UUGi1g52PRiT4Fu2
DEX4kQ1GlwDdz+3t3oUxxnCCm+TEK4Fn8Fz0ZYOjHHaS2VoMQ6LfyXTj7e3BbZZcH9B7lXz1vTuI
6x0+kyDbgCHJXYNCKKCFpD8W6rNvcqHiGMlQdX0PHV2lFbOilQXe1GzaH83RQwvbf2qarOk7miOX
s3MPRlaiBJXwByIQVsnTaOQaeCyJL6kneUQ/ZaDRBTB9cr1Um9fOX6AZzymOemY6kwAzFeFi7zc7
51+Lv0wkgDkDl88YZlhR33cE07/VYDLLDz4Vcuy8ZjbIaW9awaO8yxxGYebmEcIBFEV08TdyB0Zt
K6ipuE6qT0w7pK8OnCZqca6Pm/lmUXp3+s4AM29GxkTxAzOMzuYGz0r0T7aNDbtSFV812ipGKVsy
V384h+JoXsvhSz56cRZhr9wx8Hl1L3PtvDoYtLZs9E1W65lt4Di3toCUsZoNqI4LgAOHkZ/AMtDg
WEwWXpqspR6+YckzJMKu2kvW5JCJisyJ7gG8zOeVXB8Ah5SssJL12S6d1l/t7ff0Cckz82dyHI7h
wNMalk6Z4VjFW1B6ZmKLyZsHqf3oYhf8/jKZMQleJiODD1VVX7/AMB9xHTRQC5Gy0a8w5aba4g1s
eLJROYBzUFr39xDQKHmHcioPeVLXTHhbQyOpfXshhchV9vXdbAXq0Ru+J7mXxDDeBz5FR8j3k/Mb
jE59WCMkt36iHGFWSCInYWXveo53GX2duQ0E1RDDj/cB+nS94fkQQeeYrG3yHeWJ+b7HEpYiJIAb
F4MveXO+iUYVWVtBKoBCASkgN4Jx1LUIG7tuCGWNdVCP/eeoZb+9y1PT2Efry1vhNyMhN9n4x9To
wykjoFyjWy0plecumi7vSbqyNX19NNCWU2V+eaWV2KzjWbHB3OWTwqy/oX5liw6xwcpwHZxk4mdk
6FotbgLnEZVofU6NYDZrPXEHrxTLJlD+mbnG0Mlz6r7Iroe0md1ADpclTyuLSbkOA2oxxPTeJd1Y
/KLCX00YlVDVvVpL9npDRMrW6drqEuTtG0o1bix5UC1n4Joiwed6CMXwC+ge7n5COFVC24P8io1p
cleJGsX8ilproG8veVi4MTn9ip4duy6awhJeFKyWOnAvU3rT4NYhH5vuhLOLjluCc4KL7CKHIBqh
1evDpBbzROcPzFnii4/nzfeCyD38Uq+TN/2B4zBHbVj3DGp3QPBIcPCY17GjvHpbW0x82/+bVlNF
BCQYoS5wVAT+yxytHHnRb3LGZJUTfYcNp/Pl8t4aJraUgwyOEHqF8rxJenzti4ehG6VPfD/tUv9Y
KG7ebv41RjhQ5lbWPqSfdFFuIoY00r61mzl9MVrGMNrzp0rOyWF+L5yp52DHke3hVxGbFDtVvfqS
a9+YgkhfWq0QbfB5tcPFe7ZJHofMJZezgtScxavSaMfnCvErA7mAlNFI7cyr9papFleD/OEYjfiv
Mxw2XYZeAIEajMqNnYLdI3FsqqDEVUMtYWh3ET//iGvXZFhesFIsIneIWhaQtIGcZOqzZ5HLfVTy
8DLgkipgHTF7SrnWvvmnfciimWuJGrl5M+v6tPw0MEpTPRIdEj37QoEubD7xW2oQlLvQYwawyu/a
XPxG/RHs5Gt4PMiJQeC9Ovrv7xhPYQEEN6VXsL65+pcHmaZahFKKFkzGQuYoJZrF0UV1cZQqhj8h
1SIx3n0YwIalJwGahYRQLUhnefoBKhRWKDQTnKaPb00+F04TdmyM+oQn6Jfjvx/y2rSoehgaYS3c
DIES7zhpwtn0AvxY00E0AltJUJaUIB8sLxNLaK5uwDR162nSVOyAFRYEz/U+wyCndIJpSvWf3lzU
wdzCxSjeN9PUDGfw1CA25ceUEYoNjR+t1gBPGG/czUvglBpJJAiG7R6ax1aenCeVHQ8KIL9J3y88
TDqkzYcbD3Il6l8ySS2sa/gHQPEwAM4kM6NGYZHbnLmGLtF0SkEONc16ucZu0aCaZnpuwpYnrIqg
Bvvhwco9jdpWBu7nGGy4c3yfRsiFyHiusvOpslUmIJvQmgmAEMaPVP0Hjb3yd59wCRylR45FjnnQ
C4p7YWC7o/gakOg46a+7JRYDEewEDFzjOwU6kmiLphvPnVd6FlyCF1ze/iSEUOhgoGrM1YBYoHLL
7ggVbFklvQXrVJhk/tAApn7k0ujgpPhVqhFzg1Yf+jG1tt2+5zQ2KToXs2dMNBC6OsfI6pnalUgR
/hHZQ7usXt7gGa+Aid+PcKr8XLk7t5qgCt6sEqR7RrxAGfT/NbbJo/Z2Z7Mb/5R9uE5KD62LJvg9
kDNycwFUHgB8sVKWfSyqv87pFw3KBJUXeZIZFLzXlJ7NbedDIIItLCWVLDFki4lpPffUeL6KKwG8
tJoGKS9VRyXKYp/19xYr5lpma64iAqJc8XHGqQoqZz+EoHAZUNu9dhCcZRzpIUfoaWqRnAZkEZm+
w6v+0pwitgWZDdunoXJODyQ7a+zld1QiBxshWei9Tt27d0bS07jf1xwFS7uE7kMeqJs38/Puk4CJ
pbU5prrJIvNKMWa/n2nkL5Oj2LJFjIs3tuUIHQ8O/rbWU+576+BlTuGZnpy385ufkU9WlV51ZVtP
28vn7c/MUOPx2wL0E5e9ZzZYx6NaRSC7womQ6Qj+X/h2XPpLQAzuzdsz5NpZNDvUPbO29x4PWvna
bMJ2FT2fgA78mI2ml1nZ/7WsNYz6qxwv6MvATcTZZIce8OurGX6NvHu3WsnL07gS0GUyU00zWz1U
esmSQV6evGAiSLRTNKeo4DCFuX/eIv8AWUwUKTNJbCiA4nlD3f/PxsXohbg19pixFCsmqsHoVdnH
3kM/0t1qEvmRUBOQ0SxD2Vh96yVJ7YbxImHwbtqwSW6OUFbo/enBFudB9oGusG0pL5g9uCex42WB
tODrkXf2g7c68utwKh/ePfKgF+6lXF9Yot6Z6ZY2L6SRrhnYOVV1jUVAHRQJQQT/7Uj4QXbMK3zb
YnWZuPPU2cAeuA5ObpKjQDGn3KfhucuIoIu3PURIBrsSqPOJ3r3z4DHeqBzs4iOJuQvFOIJ2I/TC
woaX6PM802dJFjKde3vn0H9kEAulfRGUW+1DzKkLc6j2PsTaSSF9jZnMaT7jj/C+nr4Ad8R+e3zJ
4BXRmMGONKcEfdHgDLbD7OHzzdtxlnONXdCNSmhSqbdxKk9t/VtAJlQdfWaARB8QynBKqSqA/8vL
IwupwDcQHuXP8/d/cuC88ZuraXrNZ0s0FNjPaCJGFkA9zxrcYEUe3kLOCYJWFbOhdXQHED/Mxv5k
6QZOHCDCcAspvhB3OtKL1jKJZcs6hEOV05LLWv+/NSdudYXPgzJFurM6MrEt3yaqNv22VlPj7PIx
YFLSXO2BOrnvlfdR8ZoilRYz0Jg4FCJduEvm/tMgcPb2kBeSy+5/zgeNYS7XD1mPfg2jd39bS5Dt
hKEZDMqGOw9wGJtn4m2+OD4lM/O0q69xAEtOZxJFYsq7MokYoizzNdu0GzN7vGR0XvBZ/7Izfb+p
U3zdu77bmZWeUgWaAh99roUBgh2frsxOatb96KYtO2ycnkMMKblBY5s3m2Y51H5nvhgAOBhGArmE
kVUnyqyb2Q9RHyjk/hX23jNYBTzPtvOKCpzbT9xfSUN+ShsvnQ5JeMzJGyJNxd0fQHXYNxAAiuX2
rdyFBeZJWHFcuhO+Zs70+PPIAsdJ/c0n/IFaZRo4ckPtgDCQJL2f2n++YAwamdAFhDzsfXXtY7jT
e3ki7YI3P1D778C1evbYSOurnO8A3i+De0dxcYpkY6gi6tHEDJBtUzscrIgncbQwJam1dZa0a5b4
E/1hv9JTBIvpIM3En/k0Tz5871VxWiGsqsh8jclxSHGGswVPwARa6lyKmWm9N8j4tAPO32+yRFfm
IPH1rYPAoJgfrQiJJIDAO8my8xMuNSZ7xUqFWHJgRu+8l3wj8X6UurYYWTuFskW82iXe4atcBAng
TbOO/mBFNNdSOdKv3bB+xvRiL9OqgDBTq5EZgGEAzSB3Ch4pAjvUdC2b/d6PPKEQc1cdVdcmgjC7
nvqICxKBoNV2xnzQpxHx7dA4wFSpkn0YSBiRG01BTbElM1zmZUDcPO3qASO8Z+H/rKrAZpQaP8wk
dtDHFm7E+qG6jlhz1R2LYZsBxKhDKmg6p3N9+ttR/ZpPymMF9qMX++B+NpSsM35IvCDJ9KiIO4Gy
UDkenLtPMV/lc9en9ElpmbRMU0Fzo5OxJgK/2UveWEKu1Z3rJ19wniehcX6jjy5xMPmwbLA/6mI6
OitITaSALgKCdKhBoIKI0O+F6Gc6wzLrqlu3Ay/prOjW3szG9Yvibx38JUMLf9Z44Ihd04HWl6pp
gdKP1lKDtnBQ01cX0jvpnT/v8vlCDMoHHbtkoWifczYAPQMzG5vURlwlyzsLOl/rjqR9GAaTeMGn
bF0kk8Z75IuMc8e3aJlwZukledolIOE9UxBn+PCtUo47tc8jOlI7eZPgYJ6EJtbFMGJ+06fPaHAH
vDOL6PFFXKe4U364iq1TTYrc7hKJlQkyFbPEmKQG2InxUc39jmi/74YXWtsXdU5c1qMJjBhfZQrt
XhN+8GBk2iOQhxgEZFicI+9X40tplmNK4j3tKyhEBTgx1r7QuLPlDB+EF6gt6vb+eAoVKteJ0Yrk
RYMab3u96AXqrGCpRRfSaOGrKKVnG1/ly7fi0JUjhkivAdh5n8mqGHjy7IWnrFdyAXycsFwkULyq
YvqhO7H4m7FF5D7SX9AiGvKGr5/D9LsWZRZ7kwVESAIvSVqf0dRWzgcPAPjCti9A77+z9SOwshba
NTn4cROZ86X/Z4vRVoF07xXm2E+FLIJ+izITkovI8pSVrV6pU3iEa0L4sk2a+8pgRGG3P5OPV6xO
yT67u7/NfqscH3gOJEdDnTGZEG26rSGBxFNlMNg3kQWao8EQ8Lu58afTaJ+Kkun1KTJSByZ/Hmis
30D/Lc5vaDwjTroWFtLHVXnIFnjrK9mD2fGxUOS9616ho6D4i9M7PqrgcUw2vrUP3Z0raxztdNls
dt4r2EyWKTWzHoBzYFtszcXrFEGR67cZMQVVmVMwxMMnzFN4qAwIccEQNg/xVv29Sd2DqJmKD5nW
yUOgbup35OSFiyR2WyEMNvEZDpWzgLDd4+cDMRKpydwI1AO4Cmq5tcI2KkbSNVo7+gYK68cCg1Zy
a51IgeT+94GGf+VI/pV562unexZAx8oOqNrBkBzns/fabihh9oxTKfy9bneIM/bSWEE+UR0IlrZW
oyKvicVCiTFEXskwZt3QoMSvGiQ9BH/RVToO1tlTyz+Y5+tLLd/zHBVFEMDT9Fe+KJgI3MkX5GTF
Pp/Z/m7erPdX3zJJ2fi+OyK8zJ+XwCKHnALQ7Zax2FYNYFhbPo2sR2O3ZQDXDbmHKb1+u/UdTf9I
Su/sK06HhR7v+9HIMV5Zl6W9wFwvl0ZwToSvLDd2GrzyTeOIfHixi7rqgbnloRlBmW6gYmbpco+q
iLhxHBVMAFNM7G4y2mOfvap3s9DH4RIyyKoHjL2nji8GRAqkSP7aLQOsO6kdw5CldrP9bWB4Az77
vene25MJaqQxYMNXNDYX5JgUpD40prUangLy1LGsBtN2HnXv9+DIbhw85ION8LKGw0rySwmq6AUf
oKn+8rdTajNJUUBeQ+FqWmp433OdlDadzrBgJUZgHGH44gqLdyDgyUNtuMvgCmZ0wdgPnZAMJz/T
FcGwD1gxBL42eiEoH5IZDxIKLyMBIqZxHPNlLO51INC/m6zDJNxq/KjPqIjQprbOoFWk71PH2rAa
GI2Ag3xQ85OXVe0oaw6itMn521pr+lJJrdu8YHtBcfuRWtseyY0fYlc1WAj322dA5CA0B9LzGVg6
GliQdXL7hNgLJj2x9ELNqESGorg3z7p7Mv4emE9wQc0aOxpzh5SiHDD9QGQYL5RX6NU1IOk0e5oh
YJ9p8a2SOTesTGeA54Gz+zjER7XbegZAaGCRbxgHP/GYqsxi6vnawaMhOOSZfQxQFg6c7h92P6SO
aj+02yREJSLEhvl5yfhekI0C6HWpHw+InsqnJvku5TeDYSHffPwTUFmWkDPmPQs5Je1rq6BxhcBb
OZBbCMPHZPPRRYWHHupfYCHSpjGDfOJN4WCnrE8ITxF3t+b7x4qNaSucAO7F+iIQBfsEEgaVPD+d
ueg2XfK59/d31xJCCe0h20WHeOyFcUozHjluOpy+VVnvrSDw0dHoN/LRiEQ4ogu2377r+l4FvokC
mmWFD30+uqEj2zr+4ze8RZa8MWzRJfR8pitXhrn5ViPeYo+j2FS7hVEdl9Nxp/pg55PPWbdZ/wQ9
a8Vq1xD5nq2ZYSqEZaUPAsX/q/uJoaY8xHP+/L1LIFNhs64Fl9qOcu84+HblXSe0RlZqcTlBBkFY
pEHGlGC1RiqWRkI7Dhjs5aMT0N7plHEGcNdSeGR0f6/WlAPKzkqCUIr8zd84nfZx4WkPleoB6CbE
l8wS0Vd33DbcJxrHogX2JFhTAmI9LOGTDFMYit98BobFXWKmNMTuYVKe4IZrLCCxVTxu2B6FpOQc
DUXJP2O+deIq9V7UM0/0p9JoQgT91HITU+hWlcPLzfWk2YV3FZxyM0jcJ+mo7NNBE8TE0Fe2oXpQ
z+e18T9Na0kN87zyTeK7bUAyjrC2QFHcIDqpaKkRExZ6jMM+8y4IHC14qsaR/MqAY2OmxUHUXbD9
3709+84lGCtugENtVRVtUr5jypvZZYmn37t0qiQhJ+Py5I4BcmI+2EWTcHukWO3NHYV0SuvDFijT
BYUd7aLaOKZV7V4yLHEQQw6qpTWEJw7ps5FqLLYOnOBXPqPy58sklB3IGqg1RSuDudNS+azxEma4
zfawo3MfTS/hQpjdZy0JtOw2m/em61uTmmmnMiHSIFJsp/eWR4LWt7meASZYtB/+CFNmAVWwLgrV
KSqthrcGpChF5V9OtvcjL49Q+JePwPRlGxkET/tsJ+JizBqnQNqSFKMdobcFtUSFPLMEyzmAxeNc
JPfvlHc/zw/aACJH0rvx/LEftF/KC7rL1nVCcVhLaJtsZ1y7nxPyKTD7h/KHboYkcUZhFpFHmuIO
S73Qi3sL/ClJH249nSCGmT4rUIzyyLGw7Pz13UjIE7rBl2j/XXvSyh6c532+6nA79Eh7HF0MSi4i
aJs8gOlyQciqXHLEy/cPOPuecHEA4+9miOwIcRnRedkCiDinRH2I40cl17eHxjvN/J9hBOxYdsSm
EwvDQmJIzq3BugGpqRa9WYI4EVXHsO76KZijRzVTOaqJXctOk694w21ACZIVgaGFfRWAas2GoB6n
OkBCMkdMD9Q1oInpjp/c0mRQsuaGfHi9Tl9b6Lot8X0ChzWNy17ZjW0F8jOoccDh3r+IjnRVJk5C
Tn3nh89c66igEPN9N4v+1dwn0ihoRLQHoxiDtDe3nBCtnbF7tYsZVu+RdJLmLypRUJ6cONsmHdRX
0CZS/OaCMG8eA1KJPB6d4SahlaDrMwpXSeBT6Z/IlAHe5vc0BE0bctMmpWnbZlgnJc1NsUw4g8ax
dOLlAH3c4N7KgZjEFWdyKLhzDzb20++K94lOeosTMWlZGvXL516dGyB3m+MnhE+MRPsZEIPNGvCv
+gC9/kdHzHgyE8uOeaabSpiFQOH7CEeFnjqA204Fc142J7q8jqHZl5gEjBTyvX4w4e7Y9QJozAQF
uPIrGE+mz508+InucIi/gC6honw+l1LAWeP3cmgWBEJ2zqeKbn2XE7ANdmsMkcEiURsdlJrXovFS
qxV9TFB3zT1VZ5uBvjYdcDRxNoQbNpo3EQ0oO7+FN4sD8XQQO5KeIHEzycUZk+12zlbfvARmlpie
692d/PqxQftrCpkYZBOc06sdYF5Er2lKN9/bxnAQAtMppxY62gnaSXvQk2qkgNVOrfgz+ef85WKX
aHyM1BwnZgG0XCCSozvHtCwnZn45CS0wuUIpIojzceY3fN7DCB0zl7CLn1gE17OCoOQj2CpEQ6Zh
o8eUXml3Vr7a3tAIp5+sDE7gSt0mHKAHRnawUBNNsbp4JjPubXpqDH3DunjUTKjOe/V6zGT9TJLh
J4PasUrHRuwheEVt6fA7l/OroWcq6uBE11XvPTFCL2DlV+ABj1YhAHSxgE+a7QrqrY4AQ263FEN9
OeEfYICMttcVjh+JWAI6GTGlobUmQRWtrdcytPF+xtbnbOS487KfknBC96NNICUVgkCXw9a/9tT5
0DmR78TMMmxWqUlJhZ3GizNiK+ArzrrNnGO5ZY4ESMUchyRnFks3TBt1UVPwBOS87PDTlqDcgdBw
jadx378cSL1OsSszl1Br2KI1Rcgm5MooFDR1XFftqHqe14d+va7SEetZYx3Nr/Q5At91jY2tYjHM
WeMYJnYq/l+QCtt8gPg6focYCdwnwc10GgNbd6c2jnOW4HpRysGBU5ZX3qNHMDRezjVPEUe5VIum
eVz2ZMPVjBrrAy7vS3El2zPmg6GZ281wCSBrli4dHvu1rgLHQ6RLDaKyRqQqkpUO+iQSRw8GMGmh
ZP5G9mpoCJuFkpo6CwtcmenReLdNrjr22CJWG+bCp1RaogA6e/J0meMOchs8t79VaKFX3apwBbJV
wQakK+8LFEaJ/ZVs0NaMH66VNhVfaF0ocpK2Av1EAivpXJe80TlLohyHzkZkkPTQDJ2DFWM2zPLM
tIrbRmuaYzYrtRayskpK6suH2MYDSdO1KGbVdhcbnuFfRq0R+j5giZ3yJgGC0EBmEKzFFYCK+5Rc
aSA1I1PbuwQ4RuJ5Pok1Y8OL6JRhC97AkCqSHg288xrC8FK7nR8AGWjgArSVb18nWooCk5khkqZ7
MVwngHO0vcRqI62PrIvz5TqwSfludjvH/wXfiXIb6FQXOagm08BhqNStZUfVZ0rkBnVUY1Zv8LjX
jn1vo/JMEEwrOaz3zJd0iPQYWOCAW1HUSkMAywBNfcE7gnVIRjdpLNallqDj68cE1ro39x0obRUo
YsfBRNDobdaO73rGVVXLZt+5JsN5RGQGlK6noxRl5I90calNgxL6mbbTvIf9+YPVQ6W3NZoQuzPX
DEVbJKYdqM0pJeuFaDXyN/dfODQeZZX3Gx618b++TLo4wywjmwHe1/wkeiSWBLk/EsSoq1ZC+D1V
drzgS8LnK++qMSkGZlIyv79TxPQhhvhUm9PCO9y7Y4HaT+NP38jl290kvR2PS9L0yR0BRrKKFKbo
XeY0Zpq/oNsDtGMgXAzomuRFlUW/vR05tHHHZdcvpw1t6l035/WO/qlsxMBooKHkxgIfuRS1xUcS
8UM4MbuA2ayESEhXi1OSqLjVqp8BKoakbahWhe80GBdGGCTmn8OCSXKiP7Ec+FiRIN0woOnnOj3m
kw/yfCq8KXIOqI7VzffqBWVeo3bRTWHIWIH8W5RYiBRUJmxGBO8zqBpoPtfMwSv+pELjosVei/1H
hgquTx6p7ORXp9W1s3nrJNeHej17hdrBXjikiPX+Sd+t0fX5ahL6cPkwuwTkPL1EwLHTAOlo6ARk
7C3ek23KTEVQERBLqsv99BmhTxxx1ChuRmZoXXVvPzJzCh1IDqna0SUUUCjpveLzRPMzi4HUW2tH
J0hi08lnQxP0AWWf+5icR2MLzG0FzkA7CAxomGo7+xLuX3mChx2K6jxmAW5Z/T3tvMGW/c9zCv5I
ctavioLCCOpsslsnyUDi2guNAVL0lHTqRQnuAPrNR9ye8Pi41nGaEWRCowasQDT/+7JkrIGQG2Zi
0ZWuDu3ZvzFg5a5RymYjK4OOtYGtU8YyCZPo1tzjepznZGIN5LWJ8b6+vrPATHlZ9gxajpWoBGQd
IUxvQpXtPyuqU2NkOCsvFfvdVREZXBIeEOtJPi/xY/B7KzegG06pwZqBLluK46PdHZ6g6YCa3qUQ
c2qeWFqz52VF5o5Dz5ulbogUVAUaHkeo1tLsJ83+A4QR+W9tbbnLSlF1IV22JGMcbR49I4MMS2tK
ckQUh3exonP1l7Z1XeQjEBA+KOFRpiwpoOkrrrjBwGjoip9cQQt+fFLGqqnf94Xleh4dOaqvo1p4
3YEjqaNMQl7r9JqwNguzUYMKoaFieIwXU1SzSyPSZYBZTpr2j9j1QXeV0jFVR0lswGMsoyEWifds
wvEBMeMT0g2JmACbmGrBIVffYjReGmLipk9lCk9PfhKtA8v9mq8saCdLVzRi5PRxvXpUkKeEHdZN
f4mgQHacorse27evRGXKeETq/MOeKcTQuowEEg4P6zDNN10Uel53p7IAl0UhOUvdLRNpzsngOEtS
LdlhIDVH7qgH0f5u1LYlgYJgJkfmWBi83c+641KdZmoKxIvpY1LI0WX76a1eCRHT8feASNdrgdLp
WenILGLgguexoaJ6+ZJn4ZqKx7U2c9TRRo1s4BQgd6QYS4S+D3QwsUJXw7f/wVPVSOuevWe++xY+
DJURtTesl4dMPQs6aVKLc5f4A5AkoW+nUKw8ruKKtkLSFE3Sitkpdv4l8erlDJuUgGlJ2hw8hmpZ
4yQIzIYlEFZ0lEL78BCGXLJZURsEWsmFv8g32JwQQzVAPJrNr8ZcHX07XjPLyCyRAhmgs2ggCEgN
nNwdU2/Q1iTLV01Zdc0l6aVQK1iUJfaGAuS29E0cRayE3bnEIzjVXgrK+gFkYMxIss/rzH8oGCxI
hrpIKp8mqyL3DSDH+zI2r1X14lmqrdhd7gi9jgcJwqUO3DaBnax7IWMTDHrmVrqK5eSBhELsJqUj
yDzhYssEjtDstUW2xHY5Oe0kfNHyWDyy1bkx4Lnng+MWZoEIeL3SoeN/v+fQtlLlkpwArVF5BtFT
tlTT31j0DzMfrMyxk+tl52vSrLkyECUNiYzYvHsYfWfcD2ZtVKHlEfPpT7+dCVGq7EDpM5DA59Pb
3CL9x/tt9V73zAuPp/OKmtoVhuU5VpFoOWRA1loBZXVNE6wrvjE4g+Zb0WMkeSwc8qXy5ulN6XJj
/EjxdIytjIDUHkPDgG3x0dBZVxJ+EhV24KoFKxvtI+yyFqkFn2KA/24Txcuezzm4JJ1Nb6REYNTA
F8Ers1D+Uq/zKnJMBHJ5ytD0I9bRL0iG5URB90kvDwasKVOdTJly+p2noQDt99fEUnock/hVRowR
wQpuigufLjeBBRbgTHnOzzvWuxQkfhhFapUwstV/SGIMdrqgZhWumvtj8TQR7k1rWLGH3gIquQm0
PZO4U8kMi3GY42wWsdPIU+qWTG/t8ArMoCX4RIJUESOyb5sp/v9fQnkYuJndA+GtTX06EIUzn9xF
TwSESPdRbDNM90K7PYcd3bsUJswXENJrc53jccZewZCmeMvxrOVAgXG2A7ZQuHht5oikszVMjtAN
7/eGgARGID0ABWbDFb8ANvCosOA7rv2UspO3F1LJXGmnbnB9IjUg/IR0xC0oByoWrFwA6jt2MBs4
LP1BTqcCRpihSuOob1vZG9PtooHdW/Tcr3f0IAdyhkcTYSEBFpKfrzbqeCJgK1V7/x7/YbL5IjPe
o7q1dHGwZbdnD55CcCnqufJFI5q6cn14lQ90xecFSKJjUifXa1h/orlHpkJ5Q0QZmTzkbp69c/P0
gM/4/jk8ZhndaveZx0TShIEm4QY8rXLCoXA4ntaZr2STyhR9ZW1tbd61UDkGA4tiz7h4EsTyGmVQ
f4mDmZ7rSQ5OvckZ3eQN8sQMyCWzmxC6XCEXJv+ZT0s4YWhvYpXL9u5Jci3VBCeqDygl29ay07pA
X1cJ216uv6lIHXUHRsrLVv4OltMhWLFUzFgRZChv49ctCGmn8pvJLjPxRw6QexnIItxDxPZu9vIp
yMMFq8zVSa8PH/NT+rswaSbd0oM8cbnpIUGWB4HcJymBgB5Ihp8GR0o84Jn9lBsdLV8cD318aaCT
1xWFLJvJ82mftNkUFu2DI8VPjcH8FAPM6lJ5agZkoJK/TmxgzJbzVdciiE1ImB0sZXzwrBDVBJ5U
L+hjkRysvz7iQm3DHLe5sSZMX4gI1EmwTyIe+Toc9k5L2sh8dNbGhJsIqUQ+PjzFlyNz6ErIT/z/
ygd2ikfdu8aBz3TqUsRmSsm26KfYP8MlPqNdja5tQnV0ZTbPWtHyYnybtpetiq8h6rVQJqnk6/Ff
zgZ+8JWyvKsXKVtOxlviJ+PZ/IQR/943h0VmGHkuTNaWDyBWvKE/CQ89ZU0S4hosCC/La1VwJfb5
eMhmTAp3Y59TPjncu9/ErlOKTItqkMhDlZ/K3wcRMM+mw9834IdqF3I9KJxNE4zx5PmZptx462vt
JKASF3AkA9t917XGCIplJ5ymdw7RRmaesKwoF7umi36KzlYj4xdyIDmHiLfs0Tj34pSnM26Z9A/Q
cEJRlz7NtwnBA6Bi7oyyCUuS98d4jPDGnz1nWBKu+34PfTAg05LrPXV52mNKdxUBWes+67gO0Jho
VetvGlTNbl8LfPyqFcdB/QiBNUFlFQEgTPzwxXq/qWwYvKIlmLj8V3buyhNtT6BEKkg6qtSBIEa6
odXUIz1Xics9tBCw4vZk4J2FmDYuUwt0SNT2IEnfA4ZlTMsohy0WZkzlO/iyywEY5T8yYs0vuFnK
pWiTWJUfYEQAMI36P5pxMrVdz02BPLP8nNkIcuFa8qhWJa45djoWHD1JxLk0LTKMDW2Sr7E3DMJ4
Wh5Bz7otQtx/1iQddeDNdDL1pcZnj7op62tCsvxIwMWtOG++kHEa2cD5d0MuK9Uu1I6Y7210S3Q8
vslJemyAOV4XadEyfUo/Lbw5JHG1eL4j0YbU/3LzOCefLKlJE7C4Ky0aRAFXEvCNOmd9KjFyv2aO
GBx1FGxuCKrdu/Dif92Qu+hT33YmE9IH8xR6tnLA1QuQXsNJfFnDem1t98YWTCQdHldlYLy4UEDY
DSfsP/JyqlhzCH3eDfeALtnWA5Wv7prfogy9lqH8ZcsNyDKaDTad8mLIu1eEnaLXICl5DNIppdfK
2PDZZ3BrkzR6A6dUKcx60K0jsQ10pEXJcjBK4nuJ5DKLrqQhZuIKKCQoxow1yOdBPIaMneZyMJxv
M8CL72eD4K0O3F+CgZEt7csOyLmR+FGERnN+k/oAgRbzOn/EKEx+0hX7u8vbeahDbuIpvxnC9Q3J
FBzD3KuVEmkSwkNXP6MfpyOXPjOJ5buAneUrN/BccjitMvfc0jO+I6jUzXMhmrw3eDfCEdLE5dtg
I4iPLA0jJEF6V0FFrxeJrisG58HgAISd3FdkXLZZIlWhEIf+B/dXvbmqXvlZlbduZb0Pmni+Ec1t
pfSjxd2HOLVzPEij8oIKpGXdZcep0S9G+PAC0YpsTblNs1PDmnfh744pw0XXAHvjjW2hRrvOilUu
OdZzyYLesu5GZ7W1+nbxJqh714Y8K8G+V0ZMRVCNW+GKT20llZh7z+Z9wKLBQOqLv70x3VfNPlE4
iW3sn2mJCKSRTmvW4FlvUY0z7GBCV3RyPUeIhnEX5SPndUNahSDiR96pLw1ofM8F0U3ObBm0UwhV
xERTr2DjdbIzvWkqisyLT45iJhWb98cgDR3gn0E5fStduc8v+ww2ajP8Yc9NGR3d6Eyod3820jaq
uk3hZX2IPiTIp1FuVP27C7WZZFi5UljRXeiLwibPRB73GdHX3LtHjL4YmrO0YAq1ISKHEB3j0mzT
OgnCo8hjIobCrYK30jjsyZNQPibEINvL/gN4bX0SWAo/ecR/gT/KOTUWUY3/IlArywGMpx7t1puC
AL4T12Gc3tT9l9OevL+xBVj4Vo1unPEuW/Q6hXeJOdvbxg8bYJEdfkw1v/nnKQqbckvo97bcqyzg
DI/50M1CR0wG8lLVeI3aMEs7FujaT7ZyC+f7kNhnXstZWRlcp0286HPHEHneSV/ZT2hIGKxWNWJ2
dTbBTpABXNxxXeihYNSdHHKGH5wuPinljygo4xsd1MjKM2dZuFF/Lg7h6uItio7O1wT27xnbQPe/
pC+B5kBioHJNDRCHPlyOW8LydkYiY4rNO5/j+PBb50TuJIa+luzABYiVkAgJ9H2W5lx1quO+XFtX
NCt7YLMSJCUxHBItbRk03+VhTW6gub4BBEOAKnng8xFfSsRJDWxJsscEtXsLNvKkT2104aj9XItg
gGf0EgHvxVeu1iXD3dvvKuB2lC6U7LqToZh1TkaceBzvrMkJHQzOeRpD4sCNeFeDOF1OBDiLuLQX
w5YnAqG/uONDcTewEe/e/WFh7WnZs97bqsFwU35XZEeBu/bDti9RTEsGZh2+v6rtNnDsOXArJ1t7
iJ/x8iMPt/Itlpa/YIWVOIsL6kek59G1qGHafOF7w5R/r7TqkdKbgyn0SZrNHjtz/w4vzHS27f/O
TtAL1cVn4gvoFbwI/4ggIQETQ0eF29YAsQ8jxaNudoDtIQeEar0avYmtlLeV8ZtorHf9iO7iwVP/
rD7CUmUUnNIm1z78mYSF3QoQjj3MSbneeJi+eZVaFXijpkmmgX1z9NadCFgromnZrSnz5VnVLS4d
rmPHDvpUCGdgv3VyPFzR/6Bk6+aZG2V7vzFA0nw3ooeW66SfITojAV3OF4kXqjl9vlbif+cK9M2E
SRYf2jZS4wzuPTnGXN11EHTSQivB+4WuL6ssx43VyYX3eh87DzKi5PbEtFaJqg2gSCj1nMnXvrWa
8ChWLgMAmgpqFH0spPnRjxECHJ5sE+rC+nZ0YbZ8GvmzpKyKSAEt8PDbMTZ8fof4UHh895yFS1DB
98UgkElnUTKm/u6OJ/W8V7sabF2r2/YsrOtwlrcfKeVIdXeJ4AfgR0fw8fZ1DC4RjwK5Dhh2k0w6
Y6HJ7mYXBcFtJ6YFGgTbk+uvb+sjOmJSXvKyU8qqOL9uSy/4tlvTqfe0nEoDrdEyJUE+F9ADc9t7
to1vo1dD8W1caAMMria4NuFLokNI5wNmLv0UowDElOvIAclfHKXwc/8K8MjzPAUUqasph9yzmrVi
JuR+4uE9lp6h3Db8kZNFhXuVQC/jNSqNo6AfhxRZqIton9U4UeyQAJSQQb9L2PTdFUsgX2XeYPhg
DK4+PtaGlEUoA/NVnROaGIQ875MDfvSgp/wUSOmgGOnx20wYjLHNs4qCJgV1+F3Tor0CCdshUZ/y
RsrQ19z08oi85l6BlUiD8houYBD6YnFZRlZsb/CPcF/4DxdcGY5F+ZQ1YiNfU6xU+Uq9UN4wxJtC
AvKkMs4A7sJf/JXc7CkWqliM59DJ93kg667YfOVzk9IIeV1r2Mu/mPOMnsE6xMWeNNt8av/i5vpR
P3VELpxFQmPOSDWALWnBY8vF2TDpZILq6XeobiOEQtcFnUjtzD3StvSKpIYP0B/s63I+sabBJLM9
ApPaIn1sHjromsjMEiAI6ZWj6TsHBRmDcXiN5rLszzIxM5HFcuvcqMxeEkaYZpQj0aw5Oqk+CkGi
z6KiSG/s0wahrvrX9vH07SsSNVJO7Ts9mTQ76om5meEDMynBPc+4FNpzxISElFxPq19Eig1O0Eny
iwgg14rhj01rXrsC3aWGQDqrw1SiDG0UoFmK/UQ/4zatH0exAhLTTtLjWgDU8WIzAG4Iw17Fa3nt
boG8QF5UkvD2165iNtfKRn6rDOLquqOETHrlbOMqFLXmqszEv9p6aHzwoe2ppB+mmChrsx38v69G
eRgF6DOdaz154GiFNoo0IN05CwtKHoUve/9U8SFc1UP6qF/wpekS8s6KH+zLv+PwTz6ZBmXurBdt
2Sm2YFQ/tANcSxWRTVZ/6FiBye68xf/7iklNh4PsKfW0TIMSs/zyfTpDeyit3NUNiZycckMkIhY9
MbgV7eTb/TZyFmqBqEbQt5ioq1fZCoOtt6dxTd6IuVzyXPnu2gwI851jdiVGTtQXlG4gR/Y3XTls
rc/D8Ti6GIpHb6+6XDn1K8+ch83ximR7MBmOLaJWl7w8qzPzmtdYEFiqgpBx2pb/N8btnk2LHfyC
wuNVue0I7d0ntt+waArujeSJe/gPGfjOmpfneebBQhM/DF/igSAwug6vXNqoq4IZ6wT2GOAaaYT5
fcn7z+A2qjgLywEexc+hUJFZcB5RfyqwgoYVZa508eKQqLBzj31rEH156KEsQ02sqdJp6UNUkIOF
DP6sQhvJmiBhcwtbyC/Bjt4G5Hug5T+TjTd/fVvBC31swslPpjwmKNxh+TSf4807y/E/abkHkMO0
3bFLZLC6A9Z2Ju4XR5Xh5ez4pkcTqx+ZK3EocsD8IRa+yIc2VLtlpBobfAfyaRqJWY26EugxCiUo
3mlCRhIXmCLSIe0GWHYxaPqj5r5lspHpkWAatYj6iw4CM5RUX//6SIzZEeCTQ/9YeftuB+1xncJx
b9uFaONd2Sw3MN95PvtU84KoKj4upxrLeCNAFUFqHwmeJ1XPPvXARu3irvX8ABQ4MWPTLSInYhQn
BvYoRwoDQVDHfE+jEg95vr6YZ/VeDAY7Z/c9UiRRXcQxcUTA73XnTn2uIro19vjlyUduTFzyh+Gi
0E4TejSQF3tmMhF5zRjjssgEHRnFNFLRIwEcX9qSlv5WyBpxcXYCQtpQF+ghILf6sx1JdhP8lWxC
uOruURNaFNsNRLXZUpcSsMSjD2dkWh4/+XY7E5qShYlqdlfNAIuvvL4ZBR8tg01guGQaDQ0XxXLG
FHmUL8KHNfRXGbmkszUAaf2WeqPKVISHDn7FVtFRYHxpiTme4m+7JjK7zrVtTNcwSUrDIwnVzbRt
hTG5BRDGjtNJVhXAI7OuRi7BCOIK7Jog6FHN5G6HSqrQCkyqpAQenYyQaXcdE5DJGqUgJODcvAUf
e1qIGogIIwX7PXOUZ21CQelN5V+TGoUWdaEGgSVbqoyj2+TvcQ4JAmIP7DnqbXeXmJNIK2+2JyrP
/JX/eDtMkHe6tTvP9Mu0CIYSPGhVF+mIHj+2XML9Eb313+91r9TJLQVLht/4ViiG9ffh7Ts3z9YL
cbm3YoAjazm/axM82r2ql6KqPG7JP6HaTvu8TjzR8GAy6th31NeskjllQfSzut+fViOBnEpDCnOq
ll/Yp9/Vk14lXmiDitDaDdXkM/pt7i4c8ZBYI6eJPMe97SqaqCv6UAuOju9SV8GBALWlXUpvCHKX
lwk+aTGDE474M8QUE14aY8rqvOOJxnNzWAnO5x4A7vZ/JYjqLSznVapcTKH0wDMyI1X+D468+aqi
IuruvqJVpsmmjWdLgKTLRBl4KKlH6mUqvMFTjHsQs40ciMrsudMNkg22dtXCd0jTIqArY/xQNPHY
n5U3M7UZz+VD1arZgixQXvIQWaF6aa7vGZxcBhgd596B0bQwH98rGOORd5sDanLGCpJQnKJOSA4l
9n/gRVgrSt+IiGHwHh9H1N8ujI0cOxvDlLyaJml5NwTOR9a+Rgf8qra2WkFwbKaz6zwo7HlsH8Qu
ZdpniRposgQbaKWy8UwQzH43c9+bx42fTrnmQcKsEPAJiKT1Q8utThRpS5xb7aGQ77iYtsdY1FQb
gjGIFIhawq76hUGCrFr/0tgNjchinvn4mFzZX1EB/Qq0sO7z+ROCtW1N8FMQ9HtwWRAaR0KNow83
eLM9P2noc8ZK1rtBVluF6939EBL27zKDBY4MjI+oHS4xuHzlInR5ame4bvWp6Y8NVLIAWvU/JvWQ
8roGY9Vhek0YRkuv8ZQu/6+9yOzfEkTUxp7aCzCghWduOUE3TOnOgO5wA7zixTK5OcK2ykzx2ikM
s1AnXF+elOadK42w8D+tOguGKAiJnEMTxXA6VRJAzPf5MUDjvvUSdSZdlM5Lsg7IPERfckznW3pd
6EBnSrKH/GqCIaZraUELMZtauMaRkzxi6aimY+M14HcLY1QWl6wE1ssS0MVVic6Hrt2rwT6E7W0X
xtA/aOr2HYX1o5PLvPci4K1oFOWPVv+XB/htsPFpFjYB8bzuNqGLmAFhdGAWskUZkthJJmzh3m3+
WXQQFY9Ix+vX0gyUI1brUi6EiVXQ0kJcCQ6isxu44rXf+4QT2FjVSa7uXRhmIl1iyChGcOU+z6LW
/nRY/HX1jWglmKXPdsySmrpGzqhTikZz3xxcBnlrLX3gXBI5L+E9io5h3eRTRIYKGSYXpNVgvx9h
LX7aDa5hHX/5y7KQvSS/z7Vc3G3lVOLz7GOC3ZVDJd0dY209ql/Q3w6rKB2+2Vx12wpst8aOMQJc
oEtaLSpbKhYa2JSsDiwH8VNz2VTKzdZKQV/r2BNtuAkWCtzS/HWrN6jD7OcFaNQ5hj3NrpkE6U0F
3+BN/QbBwfDjC0K0PHEnQd9UHBu3yLJN8AT2O0JdLGrIasP74hmvOl7lP2i9TfbFTpqrWLsD5ORN
J6wIuY8hF8yymLw6M1oSGRhgtI8LLvXQQK29h7Poe0znIY0jgj8e/6TjbTQn9A2XUvpdhrOr7Rc6
eWNY/hVSredtgqjqhxihzbicqeUpKtdOfS3z0Aa9M2gS98KHR0nj2YEAi0Mkrawrh8L6iuaSnkHA
6eZmadRwUqf3UGN/tIOIYOl4JZgm4fXRQqA98MFlwh0962wznAdu4NNcv3MGmzpG+UN321leJ7e9
5Qm2/sxB1AywqhLx4hAM5xrqE5welWHe6HrMJIxURjCmzS5Hr783uVMevApG8FEQJvFDxU7sfDea
RGknDgCq2OIP+iVxtkoXnhia562rBlydYnq5s9/q3mwNVO7KIZyJ57PKWy+DmOg+z8qVTfUxfVND
XxSVcwsY7h+6iN/PtMrAaQSBeYXShf0KYWH06NTyRwTuRUMsWXmofQMQnzNYDnxwIqOn/w9wrsIr
CaoxTG1LWfQk90DYQZCoy4fW27SMaqNJgItsU0Bynd5zDclvaKpT6Cw4FYsfM1xlWh3FP2DlpF4h
mAtZI5Z1FqJT2rmz8hOlXvF6g5mzA0lRsXZMjqls/o7bM+bQPUPDx0HPUdU+KdvMVIxsvaYZHrmC
0Xs+kmzDbXSqwoqLWwq6TQXSPttymqTAu5B6x/Kwjf0GJRsd3AftWGa5OokP152MAlhHKrMeXTKE
SCOE9Upq9sDegKwr4Pv1jZjY5ToVlG1CI37JjBB0ywwAs/uvLGK+c221ck9bAd1ZPw+uXeF3NoSk
USULZa2nMlCUvWmsbvOwZjftVBoBa7T+qT8Zcwq48XBiPHt2JKsDNUne0Kuy1yWIeqKioMOS4es6
xIdshA7siEtL/UWWgw8DkRvIveJ+DdBLndI85wc+q/Lalv7W0/kIpHF2AKfg5n/kyLWo0Jm31Sr5
NGpBRa/iuQDdNmWpkbHaq4xlznnit0F4s5V7O2gditknR5BJaQCKBUKY7buj7u5F5YCOgt6m+MJH
cjvw26Z0pMn1mgeOnsR8LIL7eEzi8elmio2cMuwgrQpWGxmVhi79vj29DPu5KTTu+CUE3PPMUcph
WtsNGc1EWWLoJDwsQDQtrc2HIEE/aDiati+KLp8m/eaEaRJf+Hznvnmcffq/HxTtqVqdRhx0QP/a
/6ptlktUB4y2pxt5plL7/Qw9a63o3x6bbxl0AH+9gxReOe6BocTcZ3pASHRzvNpN9bQSdmpWdPrG
RaMizQFiTWs5uflugT0oTlX5yCfI1nVJcxn2jHfME0HW/19JzF8SBd59oiXfbHyD9MrEECLjCH+N
WO1QsbSAtVjdo/OhcyNy/vgFzsaP4OlK5SicT3Jxj7rnaamkAM5Z7WuRKZ6j8Y/9Ib//ZBu+c2Mm
vkoJ3/mRvTLqee7e3mOi0JOvfQ0h8FUDyZk9lC82n5EaIAIwmzZylD9iQRqZTtSFZKYNs0KzWPQd
0dgpVht6BLI8+O7j+13bDiogeW2bU4vV9scVtAKi74CEzG9FE0fK56+jT7O+ZodiBW978JRIoNTJ
P85jB5ZTy8PIdLmxWE95MCN9mjn4sVhEO67gRrK7w0QuHWzx6NWptaeq7sNNvcFo7BxxDG6z+LQO
XjnMxmkBR31iBsA1XOUCcgt2322bzPG3LUTf1qKgxzpN2UpLEJ8sgF09zerx1YUc0KghwIx4yx0y
U9uZ7G380u8pSmAJnLaauX5z1yeN+/7VJFqUNtPvw55vrq7rOeFvFKHtD0GbryWe98MmgqSTHJ93
9QmNzvDF8aieR+u8afg/XPcItoxde2X+KveiZTh0Z8FY7hVh4LO0OoeUWdgIAxojF3FBusGtR6ei
1lHpt362mU69crd6Dti/ID3N/YxAPnvF4AAXIkkcKITm2OqrbKpDz2BM+o+Rz+yXI5+01TS7fPXe
JezvbvMVP+scAzHK2eQTfhwO7O6Lb487oyMfjKcfDEyq1spuq1FlqDwMlH0rkAuJjWcOPkJ2weea
Wlpi8eQddprIeHpSHf0izutOghhKOkcEPe2334NJUyCG/Xm78xnvB1cpcmdHvRNh+Rceuze4lPgk
hpTFb2G99cSpfA5yI/nNT8+jYErnxpJXB+NJpBILxFuugTo1gZC0kZpKFouDCnDQ9ZNDJLKkBYJm
Ys5+q8P5u0kgtjIeci3DH7jLJJvt0Uw2o+OW65jhYwlfxBHBZ5G26s0ZWdijbMtSCeimyNnsUN1D
0EwinLYw838y2zfz7dnRTV9ELY1TQshSKM5GrbQl6LjLYelpN8LMByMpmUiTWZNfxJM30oW5ktOq
GSJWvtkMBudCR8Nz8YDHYIJ8m2eTCpf+ydjAPaxEw283CEQOFD80jou5XRn2++nHs5iJRFAPf3Ev
FSlg8ke9e9qmx2dcl3GbKdgtJ0YKmvEistvaczIbRmyg4fKpNe86qSKjXN4wbgsTiFmN2IunM0or
8dCMVylsoZbgCVE7e8oEyXGWrMuPAodOLsIX+fvFDACqg/5HoTRxTPW+m+GiIz0mYYZ26TBjPGIo
Qubl6rOt/c37duwl4F+QLnH14F0Pi8uCzYVfpB5JitjKBoMQQsmO1VQbE2HcYZ43+WlI6lPimVnD
fW19HaY2ZKpqBCJuruYlwI9BjDnZdFjONODhCLjNCsDi0ca6Q9bXKfSMVyJ1AS3OcdeumBn9UAQ7
1cbZVjj1am2unyjB6lbBedlLC2whhLIYLQD2J6LiU9O3qNUVo2Eg6tMV2XszZBqCAjqRqgKHFPln
Ncz82D3sT6t4DabsPY4zvmQgj6Dh2OzFrSqS9Abqno7ogwGyOQGtP8rnnUBXFrWsgDzsbq2kJGpV
yp6Sgdlb886uXW+X0LaGW9mXbII+EDDX6K2tniKJQrbviLT3iBZa2tFw6LpDN/7FzObxyK/qDuf+
FnvuYg7ikzXZnZ8jci31Bq4TUTYIA9MK+qZ1SEOC9byFXBdTZI0qgMKUg9sgV4hi6tyCNggRHiMs
vEmaGmCZm+c3WAzM/r2qD7sU+MTJq37hRwIaT4DrRF7lhfp/4te1TI8qBjHvgTa6obLI4/6M4Abi
0x/7dOSAv9yTBI5SpMfZlLzwqmMei+FGBs2XwmbdTaBYlFc7eSF7Bu/D1qwCErjAb8Fd4XgHXfQU
dwrtYURLGdzo9tDjjHiQPMLfyaWucZD24R2I2krF4yPGbg/rQDZXa5XExSM9a28eYjj5yK8I+8zO
27+ll/zyKnOOzyXP6dMlOvT4wy0teBeKuUrXMoL0otHNlMBP48WXo7bhu2IB8xh5hYJHb3u32qUV
81ApD8DqP7lRG0bFzV42RmhkvUVXrqp3aEthowtYFpCz4OZkKMn1o8GfaPHbTqwGavM/vccaPLoN
q8nQLJ/HcCa1EpDSEM1FpHGD4QRqEDbIjqnOSyRwlbvYem5JhAUVJYgOcBZdPbtV2E4dk7GiEfg1
kU1Qm8PP2UXU/tX3SmyWBPxkUJTiH7fFkTO+gZ8qYlm42Zh3WLRFlTFw34ZxPh1aqlxjxGLsdByi
Z79lk/csTt5OqgQQCMOJkj/AkD40yighOxuaWiaq/m+hI3UdhnG8S1vYODYwgp43M02cUedvp6Oh
+kqFMe4skkKya/rla8hM1wcIjONh0nzDnQv/PPMgz0w27D0jlp9s5azHnw5WxdHCsAzON7w9Iq6j
2bmiUcpUR6t2D+NDBjpiICnbokS0pqEGzJbM1KAZGqN5T6HPXQTZAt9eIe5XnlLrmEJbfjYgLSLt
aick+d1+1pfEzIRM6q6M52YpLbWWyZNQsYe2ZJYHqY7iK+aXfpMpB7+Px2+RFrbX9xkpI4kfiezZ
qw2GlQVyOSOh8/p6X3bLxh73wdQw0CUWzNZP8rMb/J4nyza+ekiW6PS9KNcQbRZVk273CNIS8FCS
24jhso2KRsiSUU3bna8mv0AaBrRZGhwfI4QSX2KSWOUINOq6qCNHv/KToB+c/P9fhP/Gklcfz5rU
PN7Not9mLVlqhxHbYIHp7nueLlEzS2W4B4JBxqHC6e6llamEHSC6Z6D7G6k9y9PD03Ipp2lS+uh8
n5dJRlFrofxAP1VPE+UyI6jziociIxMWl/+G3QNo3vWefkyK9fCCU2oWEqbc8xBxH6pk32V1qiGU
+orJiUKI2MluNqic76+9ZrNkQkNQzjdq7trtEm5BrlPoLE1TPs0yoGvZa5tjQXSYNYNSHg5pi4Oh
pRtAVWPqNivPJjb5XcGJLW0/4/xdn/ph+j6vPeXu5M3O2bMwAAcauvDRXtnXm/hLaMnMxIcfrqmh
Os0Bc8SWZ2peIPQrMZdA7UTNXN617IIBd/DXchuMve4Urh9hw0OF6Mv9uuxBi/xfJINSPrv9gQlD
PcDFY9VOHV53xrlizeLRTikMBRy5Ru/cXhZDcjPgf3zrlDM/kihu69RMgbifiotmn7b0cEGrg9t+
4bRx+YoKQ4t+X5UnMzCZvIMDxYuhcse7pDtXht1kcduVIZJMJa6MRuKfKBwxw3z9xYxBPz4Xdkkv
6Qve09JYfIQC8Ff3ncZAGnPgzORhrTBg/inleL4MO1nTgf88zzFYST0xHiGd1i+AH//aZSq9bsMc
XqG2Ngebr983iNSK64SFzsvpo/dvtQFSb3+ut3hbigMGGC9MzroZJNxezdJjoYe/OZItnR+NNfxH
By/A5czTT/YB6WuBo1pE9jmiiC1120gF5BN4wfVA5HuM6NNU7NrB2A3XK+qNxYroGPbQhz4Ps8hn
CTVXOXOA3JMEr+sFKBVrKW8JeBYkhinBx0rkAiQwEEMaHVdnDhJg7dG5/XFfC18om5wV5I6T80FQ
ky7GomdiomUmXWgZdf/DRcR1gKR5pF47Cb2z0taoXoXKftmkdZMOqWK4hN2tYirgGqZsta/JbUpp
vxfKzJoULfjP/YTBSI6WxzVCp19TY19i1OE5ZdmytF/cVy8AEBcZ263s9a7RoxH703uEXrO3nGjT
w56dEwT8E2BuXIE9m7JLAoEzJQ55V6ojyrJcFmPl4EdMlhgB75oATA7FpMA8VXlDikggI+5HPKSQ
f4MzlLadnqDXHWL4SpB5ZnJhMXxDFEq8RS8+AJU7DIOitJXao1ftJctYzMafnMvDo2z6fGpmJ8Fj
kOQhowbJYD1ScWNa8uZ4O1uEfsxOXFgnQrCxO1Z6JGXqdPfGsazBtVHcwfnYU4Nqvl1iMw8cawv0
+FmQFvEa2wcELw5mQAd9hL+XKh3R9rUazFEWUaTAt5o8yZY4kocFwd+xLTPpB8erB/rTIklXX4c9
F+7Kmiuj8Qa8KwYFLFHs0M9io7rK5BakS5ZvkHiEyMmHMsJRo2oZ8YCk1qTH5xM6AB/EuFCbo8IA
IEnkxmnkOO73mtO1KakEc54oCnSAkwX57phGyAPZ++e65J8mgNbjmBzvdvBMVOUp6IxTj30OQYSF
1q3QjbSCMHDMfSNha1glcDG39qatg1QcwK3uPKWMS9V8nQqLYqzgr2PwzcEeX6mbNqIedza4v1TP
zJBy34/9tDzFFhiT0J4dhMCNv29hFM+H6EC4RGTEN4d+hv4Cg4zsl2DEpnWdAkE5V0QdgrsdThBq
fTooxIYMdqyyO00kblvEddXHuCjto14uhrq+IXlRZGov/UTXh+iW4np9xjA+Ayd7KHrumIy0qlVW
hd6vN2lhO9vCKpCrh73LbGU3Q88BaoSUh8QVxpZY6QUTLtUOKOQZmPmzytr1R52ZIX+93uTo/+uF
KiCkEpQHHKPi94t0c7iDwMsoC8ziNYkYOZ3o+V1O8wX4LS6b1c4V0cD7P52S31J1MUDb960p2bBn
lEYjPONPfvcQDItM9suebIKkKKP6QWoYJgO1xyZYN2vCIOZUkR7PqjJeA1ao1Vs1uRmlYuj4mDh1
0aOSVdUML1HiHahZjkfenWFXJ+fjx9nhUTebQPYaxiuK/yeb2jYTAK65rI6WyZqrpuWFW25Ail1P
r2pzGkOUrSZ2k0CSwvw2/jj44l1SpqEjF9aDs9u223R0Mi3AYrol1XBcrqsvEJE2ZXGvUuDw8hDu
0y6sN2Dy2r/kAbV8wEqCKreFpnJgRC7ecIK6r4tyssFoBOLk32yyZfglqlnBWtmiFTLA1Tj3sZkY
rX9AVoqhgwRSqNSOKCegXq7ksMCqNjcEnyQ4QqF8IWIkfU85grr230HGdt9led3TEH6LT7Njl/YR
lhVbC241q3qdpN9bU5AsK+qhMUKIJEC4ZOquB11i8zEbCrWyhnblV1ZuYWFGAuMsT22eA/B4aBkI
GYLq1kehr/Qqt/Oh8eY7ueaxzOgz+YCXySMoBINQfotTxIdagwoniUm4spRjWQlIHe5uegJ4sf0h
kzXYe04ICTQrHs0czFJmHIw79T5zSWhHpgj1BATncXKxfxo0hwu9U5L3RZfjr7t6YIvVlbub0AhJ
sqJhwaO/34lwLBZpUNJ8xsoVmXmPiuZTIDNoaLv9FIvmyO5zlJySf+Lk8daZVrAnqJK7eMpc2FiO
7hzL7CuapGCGTSAKi7VS7P7szXWLVtbCG6F8Mivtxg4zl2aO42ybwiqfvr5FcwosBPqZc97h2/qT
9Hoh2jZd7QuneGXq/cDdob6AejlhhimRa9NfZW85fSi7yJl1EtRXBKI9b2Wixo2obfVufMcCYlHg
wOV3P9ioLKsann7VIKlNxVIyuRybPZyqslpIr01QWrpk7kEIIrIYWLlic3nOMxIUOIDFX2qS7tW2
DlhnTQnpOzBi9MLEp9gNAJW5K48R2ec3vGMqFjHI7JRxXnLnLy0sYqncTadvj35zxJbhYLKrjzms
WPe+8MTSYShz5+/Rup10a24kvmXdzIetS5JIK3zngsFp8gF54vonJguOt/+t4Q645VAMfs3zWsqg
mgauEh+GATBhqby1sReckInwzoNflufmAnRfCODacfAZarMIspc+PoeUvJEp8zRgilFrrrwMRYOG
Bxor/12W3FOpnmYrE3ttXw/W7zklQUaShl+oXaJIf9eebmNhvV4ypQNUFb4rfp2ed6PDarkqLwlh
Q8Eb9Sn7jdOG3er9tJVPEwWnif6hETn9cEWP7Cwi8bghIviGUVFIpwk1IaCqylV/V9iOu9ilftBS
jMW0Vgk0/LKbmu2nR972nm7vE8e1c2J00YjnI3cN2qLTkyRAjL7t8bZgOkAwxASzC309ruGD7xdY
CyxlCcyof04/wGBfr783hGFuDYvVnt5EpBANj9G5m5Gf+Tz8QQgFo4rCfyLvoRT+U+VQeKlOjdsz
1q6SBlT0dyeaeDK2BTesej9wEi/wD6Oefo9E6UZ5F4/bmvJtPW/iVu3DyAWM3L259AI+O55RysNi
augbq/4LZBNoD8Gem8YR1t8OQxfHe+zXbYktJXM2Xa1WP6eCwuOtbOCOll9X0n/l8Iqz+xLLenr4
P+6TlRe65MHV5w652KGIXe6Fbq0Pv/ljtBd+pPyGlcve+DlDEjrl1puCK34Rn5wwTGA7k7sShEDS
lodOqvAH+H9rkrLW+24H2yCyj68/gh2ypcJcLA37j5BF8HTmYBuprKaQAFD5xQ0+OM89wSP+zI7M
mkNVDgLePQmNZS3a/6yh6DUVCH7VIhDtmNFtwQJ+qRsE6eDHPMOwoFOlytkKDHK3tKEjuN+MNURR
A03yFz/uQKf/9rNDJGZtZhF5OhlRumbfgfCwQJyHxe+dieYPfNNwutVi8EBKzqk26+jLGssclgMs
Qer0D/OKCSqHx3Dwv+XIyRYZqfO4fBMKd64nn2Skfl5YznNzOz4evAUEjbmGKwceDgji7U1IV3Iu
MSv2O/BNxpO5Q+pV7FB8SYPeriW+Y+f/RNUFx/hVTv/DT/6U6JnKGFtCu00Tq7u5dIZbtEAXHObX
/THB/NY5Q4IIUF87/VXTrzz2k9a11FBu/fyrs1BX6dxNKictVbTqS0tZ7/opZ5h6YUlbebZEr9Yf
T0TOgBmh7n9W/CXF37Ih0PAjkwVv6DsPBKyZnTDOpJrv81v8lNOWtN2wwP9ncIgfXmJ3u7+lIQ7z
MScXPs6FYLGXSmPa5sNj8jo2P0caEpO3EZ/wEfuLqeqspIk4GEylLGFfW6y3EhgnnRgqgK7l0Wt3
4cQq1j7EMViLjpNCeQLULsgQR4z3Yg3mVGhkK+Abs+9KjXlZnn5j6Beb8U3z+0d6Pr5+LEnJvo7c
sW/mu1oVmytYFq4nyZEqabqpxe+PdxvwfvLeHIIHUHiiMhNdVtoJw7lnlsoC8BoKfljVxv3HbrVZ
1yK4FY5roRl3Rtr8Oj+JJUH2QgJOIlfpocc507UMs8Aa6d94r5tM+Z1t630uyrAZEwF11z5RElBP
LkIoURlK+utPp+VsXHuGPDL4sg6WhO/bKs6x9M9jZCBevc32cWO9RU48Q4a+5jmqhE8xXlfPkpX1
F58CDYrMaJmkzxyTLsH1WE6+A9DUfqv2lvBR/OSjHOkfaZJOVNxCoogYzFQJsmruleZzUaxxFTLT
PqfTSZCmazVnkqZkdPe55ib95MJ/R59Z9NkFn07BZaCCYyxAD7tNcSzy+NebWGF6e0E/PzJUt5bN
hdZ0PNjEjRr2ngAr1JPMs+Enj1JTYF8Czp/QhASuqafoURaNXRoez8URE64pgoE10SD2FzOEHAkj
jdEKKQlAyKBpJ14SGZUGv0gpnceLEDuP6sdqTGfsb8rgLA04j1S7jUeh444ImWBDqtUsYG0Nbvj+
JZaFYdF+x2UOKv1iQN+CQJwPrSJyhMCaXIRxLOzMj9vvMENMm1b12A/NCbz1SUIO4VnAnOPJZRII
cX/URlLh0/5TLbcENNhj2OSUlE3/SsOGMU4eXJzCoH/7hy7aFTLKdmkH9Cw8CfsGYQf8bWA40C/6
SyhoEKZs1XtyA9oy1bWMmU3P4X3Nfe2uD0QlbieQ3UvAoiM+WxcJbGZPvq+yASffcTxTF84kYJye
NJ5LHIC31LeqyoPEqUJgj478UO3Nme5IywaghqNuvDyYcnLRTj6o0xV6y8tD97ClM/QoPUen64OF
TtI3K4Q5cx5OK8Icmk+1lHrwtTyVjTkTzI7IfyXMK8/W1rQsoEANbH+kDN2hwDSDvecvFmDRn8mk
O4oC2pTuJ8l5+03/sKsp4Gk2LChHnD52IaWor2FQ0MCkhy14wNRyvRziWeaRH5LsnVxp5AqnN/HM
WqDI2fyn7CJ1tDIGppPSLvAcSnKY/1Wyh9okSCu+HUaddxBIrC/dtqCj4rUbzyDoYx3cJ8M6FBAI
i5s31jY8a+/AMPhc8RGyIRX26yrSH52iuhJY4jlDURVGFHuqSAKdcPRv+jBnwe16lncmQcVkP/JQ
Ld8d6C+Wlld/L1K376gW8mFtayWd9l/pNAWwNbqpC+25pX+R3qWWY8FYBt4YHirfnHGsZlc6fyJo
XYv62X9WJjvq3hC618/iF1mNv9JX/DDIa6mFAz1gZdOFYmj5pf6Y16ffafRTXYQcFaekt28ODlZD
vBN56m9XTAy3stvlnN0uErbN4UYtecQbUUjCjAXkABz4JVsYwOibCnRfH60/MKdKHbj5AIognV+0
+O4GsDYnwFOQCFOrB4Vr98IN0DX3TVuH3BNJV8NMdQQATg73SCkunuPuHCFJo4nGgw5w4jFQweni
aIC4JRDdXzjg6297hO3hn8NybHRQL63M4qhaLMa5JTsjHQaDF57wTOsbvcpeXd3+bduXttD1bWXv
lgqjF/MdMeRSZxGtqxXzLqaNHNNoz1CCXfnqjvo5ZeJ0UMjNApr01u4lopaIpR677SkDn3OfkHVC
+DqOJwPePyU4HCqmel3UU8rWwGY9RfM1/+IHa8O2pVTSM53QFwvhQ6hfaDsrbv5c78VJqwDk4o0I
OCRmVhJQPeZ5ZD64waX7DQ6CIqA1fF0alE4EjG+uW37Wv0jDHRTPA66nf9ZFTUvXVNTTdLmY1B0T
vu3kfWl0lYUgvnhd3nQHvauvB0ZsOLB3cAmfJ3ELwkoXGS8ZPpXwexhoB4OGKu1N8/UmWmobeLUn
Au3o0dALhVhU5dqT9SoEKjSWqnjcONH9Uae+wwSaHUkloWXDXG4iT3pLnvkk52yIo941rAY3dSo+
KNB85mPPX+1ZxIT2dGcRkNUIOfIrercgn45XB8T0zDEQZDk3o5ibaAMirK4EiClpb0+sF1o0PCNN
aMQhqBt4nVrEzuyxwsK5xD/l+RyYSMQ7gL1mkZHhwntzimENOuEWbiUlt+0WddBQfES11E/2MqNo
qKFvQxkwSnNss7x1GZmph81kpYiSFpmslJs2IpQx+UrOCJ4UC7qOjuLQaJ7Blq7Q6ESBEgghpnZI
Ka0NIUwjV/sIINi/IhSuxHsRTNeu+0nokEg+IKy347a8yCS87WLr4hD6NV0lFAE4A5F6W52xbQDJ
hZFj4pt5s5x16n+PTbHf33omX1ngNxTxWIz4ryxfWuP0nmdUbAKRAoxq7FOehV7RiUvo3TZa/DRb
Vf0y4+/1M/XhauNrAonBZV3NQmSUjxhuPZIQQBQpVBbndGSCeHIxxJSQniSUKfvF6DSs5ExXnNck
1Ikk8kmPGlibn8pOnf0yHTQ3uO5pV+57b4xfAivSTFR6LrmF8A2wvhs/fn6tLbPB2StFFcrUYa+Y
OsSTEsMKp9BJawC3f7WynMc8SQhOyeCntXZrJ2MpdQW4hVY2gLiE3DgOKtsfEVq7GrJkExpDqZEo
azJz5tvU1dfRnFTTeHX87pjEyf5sFykUpgQ+jQJF0B807DaUtPz3aukYqAVfMpL3pE2sw5LOPoPY
YgBsi7bsEHRTLBcm8ibfrFQiNTi65dimKNqLebWxUi9nIctau/65OyCA7wdX00jDM9CaM2f5Mr/D
zGhLBsxbmQb8F/X1A7qHI668CFKXIUMg+B8yid0IbVfWh3dwsmbZgmJi5iIjfThO9K+KOG/LsPKn
6K8tQ2P7arRLo2S37WcCyGl+8sGn1zc1F2YQX3zMiJcS+679Xx4/8yaTellpZ8A6KnFk1QVW/ORM
vD6j/VRmBT0OVKjweINx7Exsf2tbjwH8za7Y7zC5+3D38ZomHMSkc9z7DfFMncoqX9Nf/hZNkoaB
T7+JNMrHDyBOCfS7uaTdoa1rHaetVZbn6cbJRwYMcXm2O3yKNcsFshCEn+uicxW6GQHM5w4+qum7
qzJ0wpniSPEvUHLwY+ggn9qA7tCBkq+cpLcMgthZ6P28DEAlB3d7G+FsHH65PhYf48/55/2y3gjw
guibgjDWZ0mc+mvvbmTqpqzJj/JNx0u/JGeB6yv2oY4U+n2L+4CZROuR3k6Xh7M++253X3XAjess
6JulQsAp4sR6oY1xtM33zlbohQTfUMLdSLhwwo3sFB7EZDC8+WqYrX3AIrNpl2gQlq9ukzq3g7MI
xuWJfFHOS3SOFNykd0hnYROpIMPZfeebqzC1UM8+DXPSuMe6QmlOFxXbZXDeJQ/Y0lcFYdals0ZL
QMToirhejv5WnV9u8qZ8IOKW6ERttKSTRcOaA5cVv3uIwfUYGLX+17QEGR+8x80XMhr8DNibMnsp
TIGae1EDFOqu35qrsItBw1RYu+LrEevhW285gFhLr3fBMeH0g4kCpi3S7k0VCrGZoAel2d4sZUx/
FO7qJmEXCVW5SJ/9aab+Td6b1SKSgEfCTayAjpDf0B/vJdUZI8tbgPdz5dvjgI3P4CxRnwEPWKg1
9PdZ7QNtWRMkVv6Tdb/YV7cXRqWhhz4/GgTG/qHHjT96uZQG8zHqxLFBatfhRdKOhXoFZKVux7u0
6S6FZCaRaOkMjTM2UyWqRF7lC9XPHev2kmQJuHBxGLTK8BSET1deXckvJTx3xFxwBMyJYjCNluF0
RUoCQvjUJVUtU56Ux3oDqZkSqGW5OqRxVoH9mLcLzAWUb8w64DVFoE5UJVZDMLkUqyqrJ1SfH8xw
26U+A/g1ZEXbMRlm1YZ/9klqI6KMzfE+vu9fameAUNlWT/e6HMsGMf4KhYYYWfs8h+dhoRUIh/Xd
dEpDNNJm0WFk1TlYTbcXpF+D4Q3Jg9hQnQ03M49Axe4pMukHTPLzOkUL0bqPlonrZJ/LJ9ZeWpbx
Nl23B+kUp/uZ/6g+Mo7oDJhgHu2Ioj6wLfc0Igkt+6086gBnUb/l4Uqkd2IupfEPTAETiT+VT8Pj
0yIiCpYI3ELww4bm1eLmY90Gk0gvv3XNqP33qiq0U26TGxII5kJZcSt3V2GO5sqQ7d1x+TPwarCo
E5zUqgyarpll+k/VtCS0Ns2upaOnwJvX3UK3ShLtHmOqGOOIBLxo/Zu2ICnTIJUuoW2Kisc4Muc4
5vteVg/b4o9IoF9zDjNwMiSkquLf2TPyv8We6Oq4NUmP64zyvAhRqJy7kkeHcDTnZ3/0ecVnYzvJ
yIoT93VllYcT8O35wn9rT1AiEtSm7P+mX8CNOCpNW9FNZg3pw1GQSmwHNc7NnD4mrMgM+Zn5iCcR
180FJRAbPYnPGOpF/7lDz8i7YJeWozYGVrmGcLECBAziZoUMlYZwzT0Ok9h8OdzBZKNMQkjCHLxW
Kz36oToyz7hV5XNGApNx1czQs5nqXnVeREu8Ziw+1pHQcpsLQ8KLZmah38EjgMUVLUwdqAd0PKGT
CYSSkX6yRGBHCWLjg9YrPBHQvDid+Qj8qg/StXdqQuYSXJPcrkx+AB89oc33vc/Y29objFDC0NEj
lld2Dbl6Tb+1V8B9+38NJ5HBAVqG/rL/q3TRO/RXOo1EoEmhCzV9Y/kdHbBJUvddaQtHSOQtqYXR
XL4MOvmYcF+Mt6EgEJV9KigNGGo2+AXVYPq3CwR6BnU9qHzGEB3h98SsRt8r+rXyu1ZRlyuS1IdQ
kkLM1mfnGBxVIYatRKpTfR7RUqulb791KOpixsF65wEGLRfpjj7OF3/rgxxM0uL8JvLBlvuB+kJp
ctjatEQBU8i0gvClBYRFPUEbcyvAPr61OVRhTpjVUNkSoVPk/ZIxt2DpsyL4tpGj5BTH5Dz0CSKD
UHe3XvmUUf3KFYoFdO4chga7EGJxuIP17igK3teXjHPuGzCQ2iwZMdEDmAyIhs2U2SBBuU5K+0KV
UXcUVMAmuyTsgeKdWAk7gZoTjT0hWTA6NpYGH86NpjBy13YitCX21mriGANUCYofyLah699VdGnO
w/+bPO41QT8I/9fA1aeuPXAuV/Ppvqi/ezbkxDap46ie8vyGiYyUIKgQKNZq5iF0C7Z5Nw6YLM7N
Yx8H/SZoRu1J1RHWTOo5Zea9NIPWbaNGMBeJKo9OdKLiFvC+iLyOg1vUYuiC38S4Xj6qKR0oYrFj
n18A51NkQ82TlMbbAL0gB8sU5TCoT/poC0BHpZwkOjti/1oa7q4NpOP4aEj2TTuMdhgu9h3cLp7u
EFkypf3UA73ELDdJn3Jdked+H2Rtim0VJ1HsnIviLAzhgn7mL/EIkayFxjtgUzZRlxBsdIRRClEa
xTju6CEHvD504OfVhlmC5dfppW/WntQyapZMSLudAFXYztYcs7f+AJEvFkMeCwTSLMXyKEvwuWko
Rsu9UufDCRqIpScVbwbnE9m6KYAmTL5bBYSeOwuxHOHyBjgkYCf0VC05w0lE3w0oTg+5sHiQlRMT
Uft1yV1YE1EjcT/VBFFyTJfWfERfKVAdmhSz+nWcg5FFKm6ScvSS7jXK0p/jICVgL/VIb+4Qtms8
WCKb1lCx8UqosI36rbOLMchsJE4lmTWHOTP3aXWFBgQZVnvjMiy6drT2LyMwZHG7MWDap1302Bbf
RgpxxBghZNdM1kJeOxQjcf4J71u6EvkdXyasN/nspy22ZIF75LxBY3Ebsoi7leAfzex+K36yobmy
i8VMwQX7PDj6QvlVLzXA35zYR6bMV+QL/ohW23qQnTHhK7lR+6A7L9HPwb4QqUCzmET6VFf6B/Cx
KgqRrgG3eW7cwiXh2QMJFirisbkA5r3JgwGz67YEyD4N2PxnI1cbglGTqsG8dBuohWw4fC5JvDK9
fqARymX/C0qca58AjniQj4oyFDUAWmQk45nDNcxh3L3eprOqlPf96dR4/gDLcZ3XnglytfKTwggK
gWS6sxgAxNO3u0mJqahXPLvUmZCvpkGaMrPB/Ic6gkU0QmAyG4jte6RH6GzeTX+Ua9CT2U5ZkV6s
8DGV0PJlGaP5RKkTTPA4DvUxkeijf/pPtF+7cXxx0zMmAoShG5Gxdo5h4XjmIhJmUVpulWsmfWKs
evUHYLp7g9UgQ9oPxYBzSeRJ3+QtZT1vCC++eqAVDVO7fzKZCZFgBVd8LSeiE540GNdG077Djw5I
MO4oqwrQKxhohRc8H4FtX3RLGcqMtMDzPhVQHpaHjDkoyiZZjP01dcrgDuLa4wnjiSylR+VKvk8P
zyDAyHDKfmsCM6LV9Z1oSgG9Lfqq3J22++0e+4PLIUSuSrD9RsdoLKE2hhnPx5VcBLZT/hsYzPoz
HHR+7QeV7W30MtYG5xsfEUond0VlaSwhYtT6qtVcBLAw6Y6iMxQpZA5aTP+YfaukdbvD2ufDD4bK
B4u/bitNFv8r8rklHzyuk8HkGhbL1cgOgpZ9+e8S8ApdVJPi4Tpljq/6ZxNAcaOHi42jmigi5qoj
KMWy9j7FVddfR6IwDiSZWW0NQFN9J2J8lYoznNg54eiydeXHhazgyJchCHpb52Dcox/Qc6DWiddH
NBs7giOMoUPclktYxDIZy4SJf5nhdS+FWbwLeoYWjMsMb1uu0OVlcPGCxQMJa8oUVsbxwhRgZi10
ngNv7IRec8JbbwPBP7UDb6AONPu7Jf9NkH3qFtQQ03Hdt93YNaY7+ogrx5HY4RKtDemLbj2iz+fb
iSRAuf8KKbDBKTXsoV77OU1rsTyqWu70Y+hL1ij//g7+36ZJxVixG3XzIgnwE8aQO9PQvYP4JeEZ
Lk6xjNwYheSKtUjCMzXogR/rbbPBoUfGsJP1C3g9Evowxbm0WnXtCfQdsnI4S7doKbENQTFYgHBy
yNufnc1E62HA8CRTFIyo8YcZ4FpnJhpkF+kIzClKuKR6uOfes4+g1PV0RAJwIlYWVKPxuNosYcfS
XP4h1GVs+CduztUaxc//X59UgDgWoO5W6dKWJoWHrqJFX2+WiMhyMGGyxghAhmVnBaruUvTQ8fqZ
x5VMvgF3/zh63OZbqFCrtO6vQLegX2Ympx5kPS0bNgNXJNkukv9I9+Ugi3NAV7OALL3gLwkZqxia
7EDIVB4m5QSBy3Ke7YCT7I4fDwEXKdtPlH2BiJimrPQZMwmobH98JqQkZlf23xkecPJn775o4tEM
yTdK2NucGtip9TJ+AMZtNnQ+pUwBxuMHcb62+byUcLV3z6cJSD8q71jcjrBFxc39VcJUT5PKtLL6
AbLoNwBK/D7OKB1MoOrXousgamwk6wb9rzV9zkHfWt8vBK+jC+HdAX82BNFB8WkNt4AOjFCefwrB
MP4ARECQC0U35jWT/pTnaBN9C3rvL639oq/3fB+k+CpbbqpqQuFtrNhJ9ULaF1GQmyW/CefZ2AWP
FPQhTsMf4D4LA7iNgk20c4VmshrB+hyzaD2kbKKyBLFIIjLNfVcex/BpMbu9XCJsgKjqPzgkW20g
foZIx50Q0frGybWsczzVTtvUQUFaon+jwemYDE5NfNLa2J0VT0nSlDv7y7ts0VyA2hlqLAJoczSS
Un5+W7Gp67h1rXY3RCJ7HHw3RjdqZ8SOLCZTSnyC04sYi2FnsyKZ3Hz8XTT7TedmTSqPWtO5rfUU
MTu0mV3LANOpttojsxLAM8bEO5aG441yiQo5ukXhDDbXYacFtmpFLoCtmNfw3gJotWHlwT86cmrk
ZUiXbcwRbKexqjW8kFxENYQZO7PqTXn4YH3RGfGzPhbQKvWetJzV8SvIM4x7IrxTzkxBtCBx5i+P
mFJvTRncbhV6HzwNlN0DX6vhk2OPmeWZ4KJ6pQNAb/oLWwSQj6RdHa3udlUljhlmDEFvF3BL1rh+
cxnpS7pCyzRZL36OrqPYtZl2JT1aPvELm8w9N0jp6e2s+JHmVVflARbz/itY9KPwOgzDQgygt/Qy
AUBWl8Qqo/hVMKoUoi1v2RFd9Nq9cUnlyPKF1kRob8MyI302ADVoszgZUIOGtIy4B5a51Kbf6kES
tCLGghDuYY4lCGHDRqXgRXx0iLniejCQwvZ6cpX1qwvmeHxJ+52GZWGRVwjIjLi71s7ktLXs5ESH
BKmHK3Pz/9N2dp9z2bRpp61UdgOGiz9xl9MdIefxpN/mxxHxlZnpqBtQw8DNfWXOlgVgWWghbzEc
pRAb6HlVcjbO4lKb3qkHLz5trRT95pYKq1L6hoNAvDviMkoLn995vAeOYXGgtz2W2dgIr5aAF6c/
RPGO/CcHJDuBnM4xqaaZZSyrGKn7zszXNfahbXfac3zxKZrriVS+wbCp6BpedKrIvgyHNzkY4bLp
MFcTizzCA+WQmnPNiqV25FHNoqail3JpaUhezl54Imf2S97+1p6EQjng4JK+FIB5NnfvTU70qXIu
jCh2yB0pYA0BpxGnQf0YmZB+DLNmGALZxMNz1LanIT6sx4q4AHgBQyr3ir6YV7Ym3L/gGK37nkpR
OgKVf7C44P7f/ZioqvYXdPuoxlcgAwtyyAioEgYDLDAEh5hW0ezJw2oaHJBLAmUlPo+Hpn1q67h6
F2xcqQXUHPKEQItu4lW8alThjdZu8tAjv9fZ4didrDtmTwl3hNTj1oao6k0jzqchAJLf+zwjAlt3
PVG9NoHCUK70qeyVQzhyeaYCLM7fVVvCAlR49ac7wBIQoZAEZdP5gDe+mkfDGovAwIPF4MOOZxAO
7K6fuZY5eAkx9pJW+snkPkm+H3YaM9WrmpnQaeBmcLEXplwEmGntcR+vLtlobUQWAjBbgxRvr7Gr
FbQc2M8Y/wvI1+fE8m1ZTpE6O6SZzJVNc+qfNtfpx0ZBlqEAVkHTPMl+WEIGWrOUJjnNboYZ1vsN
1f9LYqeeAu+yohVySjvlYh9qH3ruTKnsPt1IBjEYKsneM4MYC6BK1L+BWIsdOOZ8TXaMPJuU7UVt
IOSihR0NcFA0wmkmMsuryBqH12yGRG2krLxKhrt9wmFnzlMiZ8VwKWz0ztADxM1GD9FLpyQGd1bo
vSAF3JDcGyIuBf37VEE1g7lwayQVnM/2q8nubbYhob8eLjeIjO2U3Ya+/iz4430je4RKeDukzuiD
bqIyYYamMnOOzGJj0iyk+HXtG7atPt3qCyFgaXI6tTIa2H5JqDQoKCYjgUKxFyXkEC2irWrf+f1/
JSqhOlKDt8QcOOsKoCvjwVabVNV3uT2dXbhBOaXGaFWDdoKIQvkBerQ3m+zA1SOeia/qJB1x3FiR
ubc4kaBMCsg+++roh5oyuw7JZl8vYSmPXQkN09Ktjbux9qqqMWX8EQUA79C0ktoUrhsK84pmfZ3V
OZtCRpVj0rLk1/79BLW8ZHOTOscgSwtFhfZb7qFq94HncbrKEA7dHLmgbXOjtYreVOGQ88Esb0kV
/9ku+UG7bH96rjdTXbESgkUT5VQr+uQAj7ibc7L/x0VKNzk4FItTnHbmtMXg/Y+N8YEpgA/ocC5K
bJuva5wERkWK13ZLV0yeN3oVuaWLrWIjBAk0/7CD82jrUP1Y+1Tj1dW5mCESHiW+26AYQACUjgKi
8VfhRWp9YLtmlMt3xa7BmjOv6yGUxsPMHxwFNLiIO+za9Gkh2PGaewHGT7nBGCqHzNOI6HwKzQji
Jk4tYkU8PdXrZh5Re4Bfoq4D8noEhUil7Yc5pFvMizZXIYXubGmz6+NJwElP5Wo0+V4yh1Q4Ehrq
aAmcmT/Fl8srj3nUGqTb5P/NG2je6uW5EIz/LaZKsehi1mHVVjh8V0X0Wf+3zVQzPvLaJRJRNhil
VU8nOE6EYJrdEVoDRKVsdIj5IFTOeEbUZXp+xR9IOJMYVxino0MBPfWcaVlXiXGDHqDPzeOUylt7
3opsk7anIBXaJzpugL0dC+BSpzuQvTeeY78okNJh5dgNtTlF8RgOdgAeDNgipB1R/zarfX7luR0g
xtzKPxSJIvCZ/8IpWwwL6tHCJCC5+9LrIMFkp/3Omn7EP8kaA8d4TRcup5QG7vXXwg+SzWJ2DswH
5mVAWg2RZbg+J9IypRB2+GIcNnAcKMLvakeW0HxAEgbMbTlpOnk8wiWX2gvpOaw0xVziF2puZlFg
957xw2mEhw5hYSTESLP/EKLjbZ4CUi2unEgf1tVySQ19GExAKhshMXUW611jPEsEkFNoowJuBNAX
mfYiJo3qAYTOeVhsfyS2lVyQCxCgSIZseBJOK2vB1VjmI8hMQSS+BvyL4GbZQNaLL4aWLwb7L9dH
26n4o1J5slps2h7JpvbE+q66d8tWQ2iGYNiJHEjCAEfiHPXJjnmzsP2lIngVaHXSfTw1Xp1r2kgq
/D7CeehHpTKDmYDt8B9Q4gZw/9Zb4X9Q/F32LEpBXn1Pm5juSI1ye/ePrI5mI5C07EVZzVvEgQL5
7uRpwxfn0vKN7k7C0cgQofxT/+wttNNVZSRsmGMWI7y/zBehHdsIhjCyAYwtfyKRMnwplP0+ZG2t
KaHMbNRk3OHmtOiQkEbrzx/bquXz/aEYTQmu0JuG5GD0d05uxMlzQlPmpl2TmvbLejVPvvElAXhd
Ea+ejPBsFETXBp0tpjmfwDO7l0Gd242s7OQgY1amCtOxjE4/19SzUxG/0kz8j1FhokYBSttJwZbq
55Xd8YYZsrOuSeJV4sD/W1nYJm8unmL7TNELbJ7mt92Oe4xVtupvZTy90TWUci29U6+k8cj+dhR3
mje1LVc9LVpJoHFTZaKC0YSewC1uhLu+mTbdOR78GJa0YvWSn0YX1UHuzO9qcW/d3Xie7NlSVwAf
G2O3KD3t4Md8k0xXvnSilZb3c1gTgNO3WpwfA1VDR8q5540CT12wubUdD7Cotrfg3XUA3gsKq5hg
pDmVNn7ojbGEi1g/6uQZBpCDD3BuxFKKjM0a4SEmjZGGz81G+U7buIxlbWgZBQYInDcTLkedmEcU
4XOevYiAqvCEpau2sj0VzUPfnZqup1mBxanT6QycLGAE44Cw5zqLcvQmUBGs7Jcnio2AVc0TBQ1L
mImmzeIclihUh3fIjcx5EeRi1ERldrkRutQZo9sA5Z41nVqW5T9B4Aq2wua98UeoJmxAOpX3Murh
3oBZdzBUZXPX7oZ8yErWXaHkzFuxvoDfVwJax8OR6FsxYZ1hThDB6sl0hxJHkl3O+/0QAA+9I0Pf
oxq9BjyjZ79+k2HErOlwRmEZR9sGjnIX+7ZaBFJy9pQ7H0g4uy1TXBExZk9lhULdfK0Xmr3O9jCm
A1j1bo6BjnvPUhmhgr/cDJsdaYMnqZuI+gkb/VkmTahR0BGLA6tE6OsCt8skHXTk7PX+1B3uB1TK
56MIqc7RrdGLS5M6pIgKYlB2XxP4nlo1QLP1lzwap7vUIUTTqMse/qP16NMp+0rugE+ceqthizQg
cezPL3hUP934f3VXkFhcZCMUYrZ4m/3wG1FCnFbGcGlITtL5uDgTMjexploQ5L358zR5hEHfRg5J
Nj19OD6n+RubaIGI4APTkjcrwKdSddwPg8riEuo8ZU51X/JqEt9EK+pSIA2IXdx3DJ7XY05GUjK7
UNnvcJTbuwAr32PIJAX0+WFF9JeJM5qsSGtBW87qdCH+0ayk3iiXW/CO8xgfoiR8+cfSdTD/2wq6
hBYnDxRlcKlcmQXYuKeXRmSSLP8Y/Yp1pF4WqfEYYa1V0ehXk8cfVUoo0Wj5l+G8TEG639r/oab+
tuXJrxm4ja1mnTNkfBhbL+2ngo+sFwt6dXp+mdXW8DHWekDklyOWF5HDCsClTa0Y6/7O8Y+g7heH
sfhO7RyBlOCHwUablbc9MvU801iD/NElb+mx/3XS9GJJKRePS4duEVd1CPUSw0EtPMFFU9zmwMO6
XPsDenXXJkDSjmGgJPQ/z19gfI6iSWTrsvdIrPQCIwAiKd8uJxDkkMknO8Nd0lz3m/khRd2sTo9z
Bv9xecgi2qk9PqLY+rIMqPafaGMdCUE0C8YP/Th3INMbQU2vvllW/SRvUE6qKSUuxrnbSE9QzhFC
/Nx8gqrkNpUJFBGjJaWUNumCUc5wrIYj+jjkkVMzIvNA/u3kmIE2fjd5kCsVj7KT9GmfWdJqNpHT
rPdvP13s650eZHMhkB8ApR8Da520ksjnv4wGdIsuQa/3mU0YgrvWFIPdkzft/bqajiKrmgUivA6x
6I6PeYCAmSNMnU7SBJhDGQEGjJM5iwrB6d2RqyfEPY7XHAwVkVCfbUM1ob9Vg4okMTdquykl5k80
bt83ykHnUSEMgE+iIZweA5uPfSreBs5jUWqT2l0aUPT8s6deCbITi64TlQgQKz5Nd2kLxTOnhkCb
nCb3zkWmWh7Z7l/ykK24P0flClW0nNVJjUj3XCbj64zmT9HqcO03MnESgXjZIRWYAUgWnPaAwVQs
awtXShQLfYnMosiLQ44gLCtqaudi7b3b7vyo0sHEISTja6PS3rhqhGwlg8mi4zE3XVgJGCZE9n3F
p7WBqZHMhtr9+YLi7+qVL7pomAT7osWlqBMxuzZCzQGPMxi9GVCOJW1vFhQL+WtHfU8V7/4CLJ8W
4ki2q5BfKgJKDZ2l2YmzNFUP8yKrD4u4eQoHI3wTdT+CK66LW1h3JzhG5wxAaYYljbbjyTD1OC6+
pSdT1wBxc7oqpo5vYTE1NxeVl0rXMykruZr1Rb7612sEuRHMtW2n5P/EaFNzsLn88Fuxf7x9iGf3
/R39PNPCEwKuBBwzMqd839DruswUMxilXx7j7FYCyrM5MB45KmNNsoSw2DKz/Qv3Bg7kPGdkZ3AE
wQCVPm9imNIo7ov4rV/XyytQHeqBehG5OYUP2zAi2cHP3oeup/BRnHqlhD8cW4WpVdlDcJMdZKrS
kG4RTLeNDyHBvz/M7sCr3IQG/bGMtTC6FqmmwYKSw9VebTnhOrfdmsSuWNZv6yksfT/RgU+ehflw
LMrB6QhwaXlddLRgA3daEmsgIK1ajsutYJ5Igri2rLrSX4g64idzLjlMcgJLb70nG6y53bkptvcW
qUIoKhDdzR1EK9bXplrAhcx+4PCxUZsPU137V94GwVlCihPUQkA0dJBpa675YVz/AUOY189F6chz
jzJwryOPYqiUOBqubPrN9qziPAcu4eYj2wL7vFAR9zMM3eecZmT1xbZL3N2F+R2ukCl71XQofoCP
hMMZYxOybtZqnKr2ZSIG1HtWtLtZRW6RNWFGpxcTjMU/EPZNZvWPuHHZ3FJtM4IgX3PqqqUQeyco
ZUi66oCHwMfBAHHJ9dTTTaP5zR8Rj0lR5Q2ceIFhI2GIR4kDTkdAeZNPxxbVBseE0LlVNp0N/7uD
whlkouJSliN90pFUnJ6S0HylAsIBeZH3iRhEMfcA3sdhtzBA404Fe36tXCZWubay+1929YAnz9+Z
7f6rj+cWiR4M9AbBvjxzFy8SBO0tjB/3UzaNKCL04RKKeUvbYwHACRYAsxkC+LXdMAxz3dztq7Jd
++9V6TtMy93SjcUCBRowLwdLK632rNV18fXATIqy55jAH06TVLWM8Byk25A2LoQr61HlJoYVysoK
aPY23UCF8X+/knvaqngZPX4Z7iL9Ey1OuRE0L80NAj89F/8VYP5SIGiQ6Ehx8bbaoRCLmC6X4e1+
sOu1h21abi1Qkk+Q+vd2seJdz+XjoLN94ZRKRvuopIaw5whdZI+J7Urnnz/KhB0pXDV9d/c8rFlB
oF2z4Flsb6Cug1xl8rYRIIHViKSZRkVKf7H8AYKbPckhsaRDUYjRGDwKV3Ub/Yn2lUoLX6T3BS+e
omp8vMilR0H5tDAG+vcywP0G6j8D4ApX9U+UUwwUvHz81XlQQD3ah6JehOspOauhN9elQcTF+iRk
AHNClI+JkXKkudaA17nmbE6yRV16PASjzeSHI+MYV8Mxsw+SuqfEeqCW2YCfzk6nfaoxN3Mrg9OP
cGWq8tMeVfK4yDDhB154C1Z3y/1Byai8nxwr4GstOb94pL0iZxJjj+qBK4QFZa1Ku9zBVQ9capgw
XLI8yRo6edBBPqRkeH5PBof+NFryysiJyQ1kDy/v4m2RuQwQ2XXrxw+dHWqbFwMgTqg+cCHHOgm7
L8tNkxDaTWfLGl8oaZoHZ9j80dbGaaLdSBSsXGD4Mtb2lQsXXVeaRVX1DxW0czjnT5cKUWQK5XFF
8niOuztTQcw7fQNgCtkAASUeFb2vJTRSfb1QQ+a+2zyztZK05DPuDzDuvDZSv5LMfyqMRBgXjuiB
Ke0pYk9cYjYagoicZ1ZXtqE77eENBdtFwh8mRTaJC63h7896VvKXZXGil2e6QoXqf9FRt5vFYVvU
SG9ZVUX/97UNtZYChey/LSM317QRcxFN92pvGPSE89oDXSftmtccSdVvIiEjc7XuN0iHxG9XcOFW
xcXW+73LAQIYgmMRJ08m+19qxhf91Tovw9AQrRNmE9VYWfCmurFLRfmhBUh4mKMtd8t+cLqA4pwP
x3D9NiV21T2LApxGx9gx6b4cQwGSV2uFdfPy+Ez58Hq2HwuClVG49h031mIqPEKjCoquBlY5120T
pINdETwgAvIQ+E5jFi1UYIn5G5uh5vSkSDFcUsQdh/vM804XrTb3Per54+IncJ8gDYSD/E8awAYd
6OFGfneccwnj36pCvVasNdiLYCFfJTUL/pVxVgke1T/L2NjUS4lmkVWshTlBJkslX1fx3S3POdv0
DZkPsUurhrUmyRxbG9vPwKHeXf9wpe54fQszh6hoLFufwljIe7G58lqvKjAVWxtAwT++ObUW+1jg
IayxTwDgBKX5ForedSagnH1jN80HoX9ucZgHanH+ptxlQXUkWRUwb5lETUDhvNfmoz56u1XECuVm
1AKA0iQ351O3gWwJ6pp0Npcqm/RMBuVqR4LjSBCUPHGipaExHtRwElpQwtQy0hqv5DBTFtJzOk2E
yGmIgvKMh1Xq6voFfo3q1cJKGjsJu4of06gaiU6Gu63zm90tPi+0C88xzS+iHzSOGj73R4tZINAM
INIoTLh1+nKNcU2pO1Lw/d/NnPY9ARLe9FqL3dmwql2VwE+TxsK+kn5HIPjhOdiAq3l32wvLid0M
G/kRl7p11QxAzYMGKhCAZ0NC0gXLu2SIzbaFOUJLpDJCAo8oqZVNKMWMeE25uK0aw4FO8Q4uiWUg
a/rq/jZ1QVvFlBbQkCMwtlY1jxsmNZf5Itm1jPVxddZz/WbpLkI9pi5EWrcJnj3h8saCG1ZdsuEF
wPoHQGfyQPcPaG03EVow3Dt8EcXnjo2pD81cDH3D2yvP1PINMX82IkvOelO5vNOiYcJjkHOhz6+z
STEqqXv7DkRvGzGlGv5QCnziTXJIK8ONBkZD3Y73p+9AA1zfnb40qy1XkswpL7QX46ZgRIY5/z+L
1pGDgF4bqUGadKQ4wKtF5Zm20CEPKyBr5oI03LuDZWkt1Krr3P7xJoIBlKPSI8HcHTszETFlbVDh
N1qe/0P3YJOHRrskxcCwtLsexS1ogsRhV6sAE+OXXxRERVRGMBBN/P4IgA1NAGYa3mkOHK3GcxmM
Kqm49zInhbq495WzlBjS2F4kanab1rzZOgzBE+DDpaoCEFXqVTuWIl8bVx0Zayajep5nebXznbkw
SCgOro9HvrW7X7GIc37uFkXHtcC8r8Mg+I5b2R82hgTNBpaqgLdhBfHDyhsMr+OFl/LiQYitn53m
pzpL/gN/k7H/FT1bfPieyVfUuJJRFqJhd58Um+i4QLBjpwlZyyoK5/Pwe0YB8r/Cm/Ebn8cuydpX
66WVZzg8MqZ9DxBMQWBzRqX52OXDycqH0dzL2z0iShzkuqJqo6tUK/F00dFVJblmEuhD2i3Bymyr
RkJE/74ZccW2YrFuhxZpBEi3TulWmkfxBw57nItjufcqJhkEtS/T8f21T3VDTQnvEaIVZIgBIi/b
FD15YuL42vaC8F18wqrPzHS4z+IfOzfu7UPF7jdnfvcgjiqaVA9G9yZxaSr9NsrJFUA38b6na1Ym
/Ef3hD0a3hikbR3A2aS5XJ2ScVg2FTiz0OUNIulGphycCr+9YZNoSA6Ze4qeoLBrz9adqW4myTz9
GuxAoAU4IOOt3+FPHKwnSZCR089OHrTgz0RDOLiV2wMfdYgnX2yweYMlQQX1Brstcn8EZjTB6GPC
db2FqtwwmHl8fHpg7fL3CL3vAf7tSB7fNglmUMsoeLMZ9FZHfHFkVXsVlO/AFFpfIUnDm3iqawQ0
nYHvWpKNAQQLt22iyNz52HBnhOcZUSfSZvF91wreMuPPlWdkGDQCTRUySva2Y9aD42UTLC3GfGaZ
vBLtyfeB/DY852hzICJpYHM677wOo/Bs4cfzwq+YKgFilpf43Ptm4bBtPWrq1G1TlzsUzMwWv5xr
70BtBwHWc1EgxmW5L7Ohicta5il5b5rbKlEn5mTw3KwHCYj2Z+M72EtC9v6n3wyOv7/nviFTcvMT
2sbRn1f7Ztg/Ib6TJshANFW8jTUyKLazzSgquUfNTwMsGE3ogrJ0vR2VJQxEoJB5rgO2pxQnWKmE
V+6/bjlB8EQ33qXL6s5dL8XBwUh1BldNiXecsgJAKg6suT19/QQjd1eZqclR/89VHf/BeVFh+imH
vKc/+FogbD4Nq5VlxFv0dCKSy5hf6MNU8nxS96tB1MRUzwMim/SMo1hwXsmz0nFS3aoGKBLMf/oS
eRWPT68vjoDhHavH7pZcPem1Y/EpcM1yk2+ZpllfGb5NNOGPH3x88+Od/zIrllBTf4Kcdbe2noEc
Ve1MtDbsCxiKYTUSoLXGab+JOl4tApRona5G9xgky40WIOrvR8Gca49DfEGOZ/RGK6xbDHc8kJ23
b6p4ZBUFGOvxLi+IsCNAo07NMFflWSuH9+AxaanqThseEWVFWr8wu0OxyoOo+wLaaYfnYifm94j7
LykXewCAt2v4D3xuJ9HsFoiSpTkTeUfMC8ZQppOb2ttXAO/AG5/LWbs/Xr9QH5+Huecugc3IHdg6
MOVQLsXH3Q2wzJGiAGoceWdy4pw/grybiQuWayWlTmtZblgzSEWjvBE0dCqI7E4z62koNjlHahP0
BnHyNmD/Hank6hlX27DtGxSEdn76O33py4JDVg5ic4WxlJTt43KL/vpTchY46FSHc9/Plh/OnjaE
cCZizPmUDWglicPjka9XfeOqAf9E7phQua9TMXSCYUXp64ojli73wyskVirNjPW2/9XgODs6fz0r
Q0nIwrJK1bzZ+NxXyEvMRT9HKW3bIod/PJmqudmjV5rG1MN8AaW/0jRTQNvL8EJ6mQYPcV3c5mHG
0htPvshP5xtnrUMXDBJmHaOYEMmu9sp4xZ42HcSUs8lUYyX98gyyv226mwiS4vdr4FDX7tu9JAwV
5PUcZlPudT5asYBGnnH7XOVKyCzCUUnNAjE2Cg9CHkLQVjymRc0XkXtNcjBrh0x1WPtJ0JgbXBHp
RKHUZ1EsxCymOTWRjXJtaVIxzn6U25s0TDMI0V1ZSYxO4lxle0emmXO1bPkxZloC1kJICke1s6De
eEEuBlOqTUmQwfBUhFGpt6Y4RwYHeFCAYSMKDZ6wV3qW4pt3JKKU5GLhH+MBJ4zmWXtcknAe8xGH
5hc5fRexz6cY04NVYx9Abx95aB2wnX19qfimgD/jLvqeOwYut9z/l1s0cVI9zO27TZiqMIUcznqg
i1hDr8QoUgttrqeGbxRxn2Karzv3RJwY8GMiVTMfqy62tOa1H/0CkT1TUPmSzt7hPQgmy6KG4TIL
6ypLT96A9qVDwpe4YSSUWaMwZZR9ww8oKq81YC607MvjjffLrtTsZbh0wSyVfGNE8rkWdl4ypupF
u8d25MIgGQ/tqbIIM/N1Y/jXklNML5oCx7DOdEgWgv+veZbOn5miY2rMprKm+JKFPtHH/qjpAEMz
/rgAfzm5cK3xkBUXXGbKk8KLKThs5ItApu2tgmjakdaBqEuZfO1SW4/eMYAv3DO2/jPs+H/penHx
pRAMNnGOkEi+MyNDewq0eMUc5O7uSJcxwbcx4aBF/Y1doYsDa0tasHAl+Mp4f31+M3OjEAdDjIHp
qBkyYvIi7pGEHF7vRxIbKKu/7BrFdL5Qhru0g11eHa2/jJVKse9j/8XJh0nb8Gr5j09T1he879Na
+RGb4EmUoWSo4VhwvTqhz4qJ1kIF0EWU8vXdPoqv7AGgARzWLoZt54BAIHneUkhkBnvW6CpAutd1
3HtvdbiPaItaxl4TiybUkZbskEaw+6Nl3+wVOoowk0sDqz7d/XI0dYz3kd4digNvQipykLKaVs4d
rL/8bI4ivxfEVMOJuLMnDoLu3fwtxtAT766OMxiB3AOzK6gRV6SK/aTEYTNfS/Nazp+jVH6v5ViL
83Xd6HRE2H7GCH5N63gTEqCy1yr+iV02mdcWvqk9kLM48qlwW/E/0TDqT1FfI35o6nA5HRAXmPJ9
TpPdedXJXWEXHKnxR9Yt6XqyqPkCzHlfVOWz+Pas4fSkHjzIedD4M9BnOL+03E0XCfXGa6jW05US
EbW1d2ktYVL13NsHMVpKqUxL+aCne4xoVcD+WLhpu0Pkj5PxSmbs13Fi6xQuqWdL7ZDmh2kTegmg
78Nn63uk0L9rah0iVWBbwUF+tUpP5PwPNWy2W8LTmvKzkDkePwiqqu7uvMNVSOfAfkfUxo6nGSxM
E7T2SuZzizmrlzDvyr7BaWIsS1zlq57KghXz1oJJe5xD4EMP6a0sXYPJ0nCzcteB9bw6IZb17xog
XZS9221FtU4bS70ynl2GX/EIQtxUuTFWqHjbLAqEcsAtYG1UR2ghpz/122tjGqJz+3fDnkH8i+ey
9JzWN3NHmbobCvykE8iBwuSUIghQ8t24FPVhY2bPoFMoLAwVsZ51t3JnadHHs51DjWMzqRni6jJu
29MPkW0X8QT+FBLsYJYHXmkPB7dkE7JHCVTsx7g7dYtCG8ScWJSKJ4gwfmTdULkg/UbujmWVY8Le
HwkMscvgo/w67mY2Kz4k/RNWzJpRegAmLiTMA7xqHerEth3CIEeZWGWJEF7B7pq1hOhmg5a8BT3G
UUcP8A4r/Dc08VihoYaPrIoBCI433zYG1H8z+aDvII8X8vsoAV88rm0qfBItJAsWnnrLYu0ltO7R
XFyUORdgAMJonykcCvBRbh0FcodA3bUAJ2ewnMP5q+LiF1TgjosKJ0fJNHCUUpMjN02hlYiQfO3y
rv7qDYNS5NcordF4imtdE9pYvfzzJ0hh1QmmxwV3oj+p8QUehAaSBhGuZAH7YZuFuYJW2ZQpgNcg
5s5QjKhDt2ZyIDW5qfnDUC0mJhhzGWa6a7h/cBygq4ecYkeIoAP/T3GMosBlfevzU5qPEEs6elgy
MEZiIZ0f2BhK4jjsLGzomNi2sPodMuj+5z5HRJ4xjGi+GJsgBqfLef4abLv4eeSKS8yq4oJhwLnf
my/7n3EiTSlzDqNwFVCjn41S+EuvPN1Fmi0CXrAYEGdC8GRBLSEcpALhP4L/ou1hEgqGlKpywMJ7
AofhplSwZ3NgbtpOE1bZyH5wxgS8llVmLTMU8IeL/69Hcwl/DPeP4bk4BboR5lv7t3lKaWKilMuE
PfDDPtje50GuR9qNGKVwEq0sXThtHrEUcT37WVsfCBDNm0v6Dqa4YDR0ZIp8108/qq2eAFfkIvns
z8xZ/O3FlrgayfQhxg11WsHfK2NrilSEH/sRmQVLB9uQbKR5ITTjpOIo1iG/x4R8fW6mkcaKpThC
21MnCuAHW8gHIx1EYRvpSoTkhTKYm7mJJmz4FBPGdcgFo9/3xXtTBn0ybTjK+NwfUEZBpbpbwzYt
Wu1U/3wxjX229Ag3U6EUZMa32f7vajN9vJIIuUL+tsfaKTsDPUKIv/++KneC8Z3LgUOYfV/RuaC1
KlceZisNRPX+eDKWQUwpR7/w9U3ZItniz6EYklTLVfYroWhclJATDklX18Y4sKNC8y9Xnj7OAACm
HfUhoFFFESmHgbTxsZNnEvBhwJrh7mYpz3wlBkxUs0wQIa1vZFPdxF5uaFqSWGrvhYhLEi4aEppf
Y7tDdiPYJvda0e+H+GloneVnDWPkgV92MadWotE1Wn7LQdFX2jWn152gpFa8VAz0uGxUwX0zN/FH
OyHjQCCq2yAeh7SIzQWbSDDkhqXjSG1cIO/ETGLnOUuP+FNIimQruKe+KhhubcG+Ulq8nK7D8eL1
HPkTuBxvbmZj1AP55nohAL03uHEwU1DAt5NT1INvICU6A/+LQP4M6DE3Qgovs4si+3u0xwLIRhT9
m0mAqdvy9G9Yujvw8yeqDXFNtkNGoCTpPeClEJ2wz0nH+yciUwB1l5VYvA73tZ31EL5J+sFR0YN4
0imVSTFwrN7CkL5jjbnF3Lf1r7cx1PaU6NgGYPleugWb/QSs+4kab1WdQcJ4pznNiln0hpKvQ7S7
kZHzzyFDCWL6bo/ZL7nT21HAzW3x0VjACuOJp9zyD/eFNLGf6eSSMjCzw0HizX103p+buYLp8EJe
bGNp2jn7NV39TWkGBt8hLW8X9D6M+x8bTGj6Ak2kdcBaIxe8Y1STy2ASURPygW1Y6eoKmCA9oFO5
exU40T9ZiMXA/SFazQdsfZ1MIZ1rDGEJZFODe1728UpeMBxkbFFRpASB3PiwdxJkmd2F3TO/7EO8
tqU2aQpAmHKTng05HdtPBeI/ezMv6ElDU1LtWFlHTwchdUXOf6dE1SD6felk+SFiwWbSb0B4iJ5S
XchMcdlczB5rpFqSOdEXtqzn984hMG+cTRy0DIr5Dp8z9+iraonBPsYwZ0u168uXckyHMbqLhr26
f3tgDaNp7lOQrTRTop5vUuyFB8Y3OFU7xdhjuqQM2zSLRZhDNziuFwaCkQtQgX6DkrH/B7HW4amw
2CpyFtFtaf/JM9FpVbTgCTSyMUdZMRupf88cJ+0fIt+MdOzcJTffgcnGlQYW0uFAe+BYTQNITSeH
qyEN+8to3Nu3zBwgwTvTlSksSQ+S+cmCfvhdVJPdyPxhX1K9IRUKKU0PxO69AceMb52LH8QMR3/3
/jhsi20Y3FRFNX1L09sucOasBLz7aN9joAdfzTooJ4EJ0KGkwfOz6qgGSnPZpJTifboHPIwdlJ4d
0URc4JzHGXYGdvlX/8fh9fUc+pY3wDq4EuiyfdQsdJ851BpJkLXl6sfRiDgY5AEwUCOwmSJtJnuh
wIRedSFc9EwAM490zFoVQCW1aYDEKSMYy/SpFq+ZrhhzfLDeIxV0mjaZSnmRXtBkf5EmGkoymBWI
Io6lRIkk4opntBEctK1rp2QxwtYR0lYcyh5dM/5QDwMfn2xuqoYtGVd2+CgDUUz+c63L4UC/23P9
zR0dFEVnUB+Ieui2UxtAY2cEjNTXjbRn6CtGUQeKVxlyfr2unWcRD3PYDqZqz1gwQf0K8ZtCAsZq
EWXYwFesVXA8Ck3WwuKDHyP59hQb3sD8dHFamQ+m+FqxjEPXOXdmUugfKkmlkzWU26YzQq5RJVXO
qXOtEvMPaGd+F5g+TKPIbmAzuz8YpY+NR0GpKcVoHk9p4nYQMtkWaXIHPAyU7wNzRh8lcW4/rNUm
l2+t2zJk9k1/VIp8PFAuwc5KCSFgUtwlQVdOlJ5zU87sFsPtSaWYcLU68QYSw8zYAgPLHW9U9YLH
ZocQF+cMD3N0DD7H0eYEAiNiZpepRNdy1B8SGdwSEiaVT34dV5jUo7w74z4igU4h34JX8iBuy111
gfiIHD2siSes9vM11u+Q7aoiZEpOpbnb+hFucm+8KkvXN6IZH69ugUSs1trTHRlVLFYTttjuXHC9
Byc8J4h2PO/CHg3T0MvM4VnjUULKGtYFsvRROILMd5igzuDePh+gCD6IYinGmbImxOHtqEGC+k9e
zVu/78N0HrGKg0T5sdjGhJJDNZu5pG3E/l5P5oYnxQiRPbeMIqskimP6EIyTPBg+e1nsOELkz6WF
ynkThazdn9C10j5W4wLUW8AJQK2yfbxX7qFUkmAMOvwNHBeGf55DY6HbbCJOOWadFX8zWz03LLZ7
BZnHC0AoTFjNsPqsMsPybfO6y5r8djI7D9uOF5af7pZVBHZK61y0yyi/W6yBqMn53q/obRFL2Ghe
pGD6hX7JswqmCywwSlU5GsXp4tcLQvkvHV21y2asR6yCCm0BoQmxUV6ZzS1/YrOItU8lj9DPbv2U
H0HcrC3cDocA6PESzfBZLW+UtvgdF48aKfH7pSwx5EZGNVrfoGJOE8K/ekMnEsgPzOMPvIIb9+pd
SuI3yU1EVYUtmc5FgNSR01XJGndX51RitpXiN7bjMFeaiwJDSOShQmHhBe19NdjkR/pcYbh1S02L
YSKAFe45nr10cH8en/r27a5nVk3uXyHqmAPMKcrEkHMQEgm1I80ylnHIZsF+RuMYTSOoun2yHPpr
N+0dTrjzZRicLxIa41ReC9vK7x0FkFAD6eYyyeRv6A8U1M9A8iyVW/GW36jwHg2yWJ3h4n03qZdr
TlBXiiyWEJFpuLV3MQmixWfIH6w9u/PN31A48Yc4PnAYaFjyrC49RDC4YSkAbu+jEPgt4XFiCDR1
W/M37xLtu1Ji9ItUfae5VBKmKv2cWb5B++YKTxoxXUuKFFNrIXBiX1OYZr7n63e/pPmRgsoVTkGC
MewGGZUugFqrRnqgvynmFYG67g/1egO4Vs1NBlrr9PZLKNXt0TKQIWknQfhmQkAwR/jclqgSd3BH
9BEadz0jm8s3v+2FhijasTAyrTFVJY79BxXSLfwLKz21f+7TJcIGGMpo8QbqIuDmxtrBqcxywsD/
y1iGNmNqZbLAGciSS0xiCux/763Rgsy3zKsc3mjJG7GNuA61hW8WhnyCUdT/0UT/XgB9fuO6JMd7
v1y/WLcJFTaFUOkWbcGAsbo9GxQJoAj6N/K8g5Bzfi2GNO0gxtSwvY6aTFzklNOQEBlbA8qPGtV4
zMUtCjBBn6LqDiEYwCev9AYRwYHpmteanp4v15WKnc9kB8RGRMURB3myOuwv+imTBW+AOSSyOddK
8s4LgCs5BHyV5D7H+RPLJe6lWR+CTun2BiQXeCppzFEJb7vNvD/FUNsGeAWkk1Spq19WG5IAJMbW
EI8YSVHGC8RY8vW5DF1UKzOG1uUO5fG4UKE93u2mf3/XLbSH5Fgfb+l52IypGzfPPb+9MhCss+Hr
mTZ/e4ypaEMHMnt22MN76jSDEP9BDvhqQbjIymrJNSm16/767bsMVuyE7S1g1JinfH67elWqA1br
2RtvaUtWVdBbAZHcQO/T4PbxuuyFKvd7H0P6UqcNjwViSvc35sLXCBfiYFlW3U/8GkGgCN9xI7u7
3uaROyVFKTFvF22zfvpGM34te8bXEc1NRdvhSnM8bLs7WbiwrjmoMPu9aRs3sLiwSbXMGrx1gsai
XpAQbQpOgsFhFynszjvXqtZ1qj7vw3mTKHC8PFHBPefbHJPgTaUIhq//yM3/seh6l3u7SBVNhleI
Dt7XELtX+SlmGmcR5/czzqr4Mmo6SGaHv2Xl9uIAowOB5kjb2U1ZjQvc3886+MljWc36BCMfw2ci
UkXMu4Uy3idBi0DlNtgWXp7cPF/2NEuBw32vSHmZuMk0MGiuqXASZtRujr4TozeUMXKdYh7mP464
ZcctuCtnWW9PA9ksDD3iL4Kv2OIkDSXdc8xLAZs2CTQuwkdVSL2tiFOwWcCF+92qSqogfShgyO2M
251I4V0ft0CKMp76z9LPZJBOyZcXnkJRYovMGHf+cqMzP/1HgCz7vTxpRIt5x0EBDi44qBoXnV6a
otxUQOp5lFUdjGcYbvQocMLyEKj9TLsQ2i+lZ/boMRUkaytjcN0q4STsGOw+0T5VmyTUxxDNa2nU
gpj341ODtCMzn+/zds4OANZsuV2kiM1g1pLiYXXlox/HWQXDkD61fw67/dB08cm48zVNwlm8o+db
iSwllMSGcBSB2O5t302XXnUzUhkHG1tfe7Hqdd/T6WBhemfDngsY7VSkWkzz9OY5vSAi9OzMrx+7
m4RL8syDXxk+o3+n12E6sCXTuogFv/+k+Szc9H/KZwuA/CepdrXW+opGsU9ReM0gKl58TII6iwrP
1wISO+Vut206fTPkfi1JO5zQydLnYqeLfzn1lw6lXbb2hAhMNy6AyRS1DOtDiBbBSRnEpCfbFYTW
NyLFoUK5U7xn/RiSUAdocNxWWWxWR1XMl7x1zc91FkMGPm8GwhMNZJ7P9aw5uOkyQg0q8TLK0ZAA
3pM7aswBcUGwQzLL2dcpPIKOqPos0hrY0Y1D1dTu/UBViDogul2D2WewJuG44Yyhwow1NELwfePz
/nCWc0qmo5ppPyPStYw+NM5stoJ1mPdgJZ9sTDiWix5n5GcFrwgvsMmHKr+HGh6Pp2lih/XZ1MA0
lUirOcUDR1Y1GT/R819R680bGMKrXhm9Nr696ZEB5A3X1R/G5PDGbwr16Tm9pkjFB0bLkTBe4qa+
CZTadeZVAgMQHRGFbcmcpIgbQsDJ5pLcexy7703h4wEO+p2qSsEEyPDTz3WRbjCD0ql8ystqSCMH
2L4Ehrm6OuxhID0BCa8iMYsQUx0BDodKbGQ4iMXG0pvLL3MSV7puTZiobmZBNEPtQsCzuW9M0kO8
T8UpFXiBNTWAj5LxkaSw2f9WSNpC3+Y65uEs3GXKC97JtmtX9R09uCHhf+3S1cj/4RXeFkG+ZqGY
ug1tWuysGYZoHbSElLzBkTyNjH1n/wG0pqR77XWh0wxLBIKT5ImjNMy+846qUqANEL1RO+GDqDVP
Z5epg+YFricnJhjtZY8UC2+gMSYQo2A3biCgACnfeMYCNr+NX8474H8Mk2M7m6IDjSYtz3o6MzDi
kReenlW0zUY6gOoBx0Id8pE0yEUBjrOhPr0hX53W1J54HYKIR+9JcBUheU7BGn/IMDvi+gIjCcZz
G+PUAzHo7nKd8BpYWfBtI/93gCgWm063s71E88wWFJLtZGQSDv1qP071oScL1FvMxgf0eUiHej9N
J16AEe4njyxrqr6Bj+qoXKM9DKrYuf9aeOd1jL0bPoyZY7gCz15NPwOWxq7NZs3v+SnUiGhazibD
fw8xctjD6D31Lo2Wbn6a1HBvo98FWXTun1uzqnc0uXghyjdrbCNa/8QrKZDwYm7SNfh0oceewZ6n
HZsXXWVGQHPahy08/mk6T1ni6rNyPt7R+h1RYwsX5RuGl6PLWfTaHFs1SLT+KkB2vX35JA5aErKf
r4IKXntJPA+2tORhbr3WC2VEhP/STidKJlu9Ujw7ZRAq9JmdzLqTHueFwnQmVgB2ca9e252gZk5H
uuPW3o3PNBxSf2pFtF38tQ0TFv3weGzfwUV+D8BqGs5VS89L0HNcvf34Ttp72w1eb4GmURKlM822
dOr65UvRTOvz2fQBAaS7GQxaTr0VBjgJZlMIvhGs68/t0aErQ99LAQKD/oQSASjUdVpjVIgA6uf5
6c3fWe1UdkXdrIHtiDZyjdC4mqnHQnCc3iLrqrGFzLtE1WDmGPmk/ST3Cikkk483XeMiSoEfel8K
aBmT1PmK+sK/yGDn2W5fv75SCxOO8AorF/fdZ5ZK2kq1Q1i48ibVRIY8rPH7E3gzeMf+wuM0iaj4
ggWZvMEMGlDkse0x1GNBw/+Nsj1FDIzzvBGlCh1JbKQwSMD95Gee2ihWe76P7DHGnK+BdKQPywZ9
sNl3Op4CoLbcX+Nia5jPGyyO+v1WIeX7GlO5cTg88Y0bdqDesJoCOfBV8FBSqWLsAaBKb9QyKObv
0rU2pou6zaKXNEKFl4DCVGREPGbPtCmmCOsMmAb2IkL29SXNxrykFFunrqmNvrZrWgHAdViD9nGy
+hsbxGOVbg2odTMJ1m8OEm8ELnYioes2CRwzHLZ/nQCw+ikkiu1Rt5ISgEdissKqGnbXBoCmn0Ay
SRojzdO03DajeeVPxIOFPf0fvM6Cpg13Ks/06P6st2Y+3sUKR2Zt6b3q8YLfQedUXE2dDpw4O+De
+MH2u7N7D9DRq+iwBSmKdfQ3bczUNz5rU1Qj/Ir+UQyQMmiPigCyIAZBgTLZLVBroMqiYPJra/Ry
WqEsDL1ugXAjFpDjB2WDBVZtPa8VT+gODR1Or4h2Q3Er09KdTyx2SdRxrR3gTCwVYcQHDsqovNsY
XjlmvZzO7FHvpqTp16vgkzMvahSIjYfYceuksZpw4hTytr3ee8IUsFOQSb9auCa7H+f5DHDTWD38
ISUfdERaaXy8yEbhREQ0bxX0oKRDgwFYRlGXH0A46fkFQborzKtuheY2PG0SdbhsXPJ3SYso0UlI
RAiIU/iGzHSBdBbfAaHB62TXo6Vi5yyklFfw5lLxULm4RoZLayW410fPaBmFwoEOXME+MzHEnjxu
3oFabGzBcbKcleU7SHLVo67DmBu2g5/wJYD9NKxVwkRERkLekxpOxEyscA8Q87+QJ4kIp20iV0lG
0yKSPmQ32TgEPSDsjf6yFKbVh8DcEtrsJngawnnlfYGIbh2TBhOu8YsSl2rlFcE422BAez/lasUc
dbjei9dITGg0bgQaSqU8t0KwQkFmJxCkvWZHTeuWHrRButaIIrVmpLYXo4u9R3t2wJjQi5jYQVFr
Ofj4/uZPizJRqR9Il35IASCWxVvakk+URsUlRjsK3DgO6Ppr7f9K4EKNQmEE7PkH8dPG8slMH+kT
yjX6uR77f+3BvI4OBXVWfp72EwrjH3Q/UtE/5EDX+oV6FiPtdZ5sBDGY4KxZKWrSuEJRaOIcgu6L
1K8JiLNT6CUaNsP9HkIehONMTxBWrV/bNnNJEGZ/aeWk1AOusLqRj+3BiJjORlgecS9gix26Be56
cDD0jb3nU9eK7Wj61yDk6M1r3ZqsckSX8cDet5BXrLU6aGrDuwSmbiCcfx/dPubLItvOyifj83O4
IDr5RHHHqD79ZxK48rjoZdNVHepXiKuRAgDTlCejjNxe/+CqWhXHhHv3CIzeULTikW5lpV/pxt5n
2tOfYWHwrzT2ku+F2zbvJRz8jeoPCicMTlBgMU74tHnE6XtHdrKCN2PLmEd1tyZDUJ1aAyXFZKlJ
sjH6T5L6w+C33HKcg/lzclpAlAFVS/IWDR1SS4pTp32nF6kgFwHhJhPOPctvDAf/DA5zqN8zt5DB
RARc13GI7JqCxwP0QvYleVzkod7RzywZwhXZYWnycorIQtWophXGKzF6d4L+7Ty8ThxFGE/F457L
0xpbyVPdNp1xdllGHz740CEGqid2a+lns1AT6FOIKi3ToJFYQPs3cLlBARDbgV5zebYLrmwqyhr8
7eQDzXJ7r2X4+Pv6xYTKk/cyLjpp5nR2lKf6hQAO67XZnHqvuNEDMewQ0tjTNM5iOcqCYTYTUVTC
b66gxP350WhQMFQON4oQc8rx9mpnlW08ib1cLHCRthtIPHFOx8s/218it7PNuS/kPV+S8jqXQVk+
27R0bzdA4BTBFGjnxegw5jqoOKfSxGFXjqzYrPrrSxK1obqPBCkX60a9mtsFVnwq6LZ64eVf0kTn
yhQICAf7KH72a44PKyuvSA1811o/YPA6ECZ8rll+TRxHmMZK6P3Qxwugw/vhcjXl38bXB7WMsidE
JFGT8t7dfKb4UyMdhSQBXqQsvu095REnY7Za7LDS9AsgCsmV4aAgSvsHwyfAuJoSDYaYfdX6ALU6
3ZvnSQ3v0G/Dih4yEEt0S80LrdRPiLOXiM2EQC6yONSPSh+ruK/K0AXW8FL/m7jg+yDc6tnrtRRI
lFQIIqXfRRrodbyI/NwYS4sCDGU+GbnNE+7rAwiuSmTCr95iAgERDHD5cti/D56EP6yXjvoAGlP6
Qz0eCArn9+C5xchD7wCerhSb223W4TAWpKbDmNmkqsGRER/q7wlOp+VcnLvEIqUNk18cfSmXt149
HCWH7j+5Y2G9vPavMK1prHOE8g6T5u+ukXvto+vhJ6cXIx+09vfPpMeXyEJ/a/eq6STkNZiFErUJ
8bVSbRAg93hAs9I3zJZduiY9HB/+Hs3Cc0cYPxV5uowMyAkJec7h4b/K1t8EZ+OZgW4JoeC93lXt
B2NJ2NQA0zl9+WAD3c/M/HNyLHR08MkhLt/9S0AiOXa1m+XQX1q8kym5Dt0FASAgDyRfXqSJP+Mx
8bwsx7j5f7Jvvp6U38Wgi+tnt9QHgy3wIJR1hyD3nbMirH/avzYZWAvzHTk84Hu1SjSiVzctjBPJ
fPQDzp1BejfBmaKV0zc7lW0+EEqEVcCC/q3l4Q7f7d/iNc94X0wqNRYW5Vqn20Q0tuWvqxH5Ryp8
pMAMGTBMEbc16wIGXXoueZlPDaUxASi//lL4Kf9iy4J+nyLf95GI4mYqZ6ONdxEdhSY6xaLaTZE+
9MDCe64Vt4riYg1UDvUIeA5e+6aKsw8fNSowHaFzs3/fA6es0xv3ZiHiCT6hFqIgYAT0mRFpTdAp
OVvXzToHDJKbWUsLY91w7bhr/swZxanyzkFqvLrHdBqfVPv8jPYrC1M8ScUnnidSFifunfgnK4w+
rsR889cziKWp9sx/B1OAuFyBM1qeg/plzT0H4fWHHOvjos0qpuJDSmZH7XOu2XRZK9RM13WB7Tb9
0Inp+mrVlVyotXr4QXghthVy5GrvYb2oCUzyR46WKu3ocCeEp5Jcw7Oa17NFyRi5Y9dFu2Oj6+Mv
7//irPEDgRg6PXImvI/etfg4RdufEhXJ3j1ybzyZMKSpA2ffaXeN1+6wckgaEHahauUIMrnHuzvW
+SF8IHqTEcO717Y8BX8KfVGD91iYU4NRrAW5QTdUUtnqnsAUcaSNeeJWqiWF72MRnq9t5YXvutbo
n1hf1FRCK8XUEODUfaTfJcudggdH8BXH/bIecqCv63eRYOPy5Paq7h/esaBhynI2MkFFt326DImJ
u67w6DIPI3kPMPlwl9LXuzyaa2X2mIxu0wH5s++b0+uOXHOZlnxfyni6STmPDvYvVwPVQuZwei6/
BHixD9oUlmI+YRH8KyVHkg3sctc71+FNApjuRbJex6+/oU52g3/WfGrnMW9NfI1v9sEVRbPBEbUo
we3lGTWeofYvXlz/Y+oYieYxZpMrVducvHBrXnvXGFKOhNT3KWrz6AFtIlGFZ8Pa4W4hp4+JG7ME
LNMVVcySYnLEVmFC776byyjmkiLrIS6mmG9GrgUgqFTtygW9zsTAvvtrRvlHmyulHMfuf9LBEAiR
0YMQA5fbFq4YiQvQTByHqcjivj4cCoExINi/sO0Ci9OqjbwacHFoAFmhWzkV4Tvcb3nUTcQ28hha
S7SpNXErhKF2Dmp2EbEGkf25kDsLFfkrBeqDXZOv618QndW8C4MebniyTqE7weh1UirFusb+CYdz
l2l/G9jCGn0O8EDy0YTEBeLVeVBKGmLLzkO4HxCiM9+AEgWzwblddLMpkVlEn4vHhHCUaGaiaffT
Gaqxdri2lmXJpGcywfgyA/xOnrsZCBh4dVQtDkLFDs+ZUpbekMg390mQfotJ2BupnWxk4XieGPcK
MZCKty7JvfCYLOy9SnELKUOh7hch7GRV3frtFcAutdL+d8J50V9oM3mNP6lb4gtsVmqVj/44jhVg
4KBEiz6YwlnbnY972WWEKRK8ozNzRLZYYTbRCaVf0lSylVa+dKdTPgrWawhtlW+qz2+ztch3edgk
Ox0IY3vLPFQfPARy+KjjhyKIOgHXyi3Hon+Ep9X8QnOSe3XvVHvJV4TPGznsaxeCCugBNo/CVbFk
ftSGgpj8yt8eCQMDYlsdqwIgNDq0UpGJhXMBaIz269QQ/TZiIAP9uDfkDamGsUpABMIwLW3dikve
+QUM2i/+RD/qYlB9pi78VA603KcVIUl4JA1Twz0e6begvd7XVcoB+uFDcVulCZ/aSsYxaWR1oDf/
FLCS7BBQfwKOWenEHwQPDebYyZrACWT5nIfRpBlLgm+8qwPJrYYtScrefqZbZ31Dvhj2+6iYjPDv
Wv9aorhInUxSnhLfO+ohVGSINbl/m1jtse5n/XKO+YYu4s9rsisVJJjo1bUIm9ajA4w7zo2Jw6k/
vKQo5gTZEnTwMOg98WVhUndIuE41JVhsc6UXlxl4BTR3k8GcyXNoOvPgSuisqDw6quh7+1g7D23l
sq0i/K3vdc/8T18QrxWMZu/CeejSu2XTeVpUr0q4gEHhBwGqclGwqvXhJZxH5YPRrNRIYzWODkbr
e39htznz2LFKbKQFh5f4YZ8oj2oUvvfwDuxmxinxpmplyoEUKMotd0lCRkiFr7xdBYuPC4QQwMgG
/axZVvi0Yo+1wml+bTPDCErqjlnaJ7DroCg5JkgqRfgY4IqjvkP6FlheamZrPGq5B3FWaeAvdR73
Y2wh6XkukSNmJVHD/T5wdrv4sxSp7TvrKYETjoe5CMWDIn/hIt6r+ES8l0BDlX0aNtbwH3jhJUjL
OJUIcQuria4FZFavq+vI9Vy/zlK2lcIOK5X7w8qWLgOxsmlPmYvYDQsO7NLxnADoZPYVd7A+4/JG
6gT1MD3qIH7ROACQejgnQ9z3Qm/BNSt6em18b99id/QzXneeTwcxUByTfq70mHQx1M9Qyu3twSxJ
KQyKP2h+lEtRvD/VpLzVjghnxPTEIgwAebDy4DnSJrXXzEkfphzoML2Xwq+24hBIScft8rxk0Eg3
EKPA0wl2kE0mFfmamAl4z3OrFueg8vHE7QJSupaiQOg7glEF5JGMMmXdIwYKjDLNEHMDj0vOGCHI
xWzGJdjFZdDNdBjS52O56BcrlX1i3TooXDFdBMm5QAn72ohxKAgGdGpy2tpptiYKy8tKiq60XfTK
ht1fjncxrThMK2qoVu4ViCvroAEHc0Xlnop1mz/IHMMf/iEV5cSYOxAahj/EbJbHT07RXAZ6A10i
GMMefJlHBUuezmEylayecqu6d+14tYUGCt/kIktSAR1kkaU5Cu5HMaFXbQCmc7VcuEd8tULfNIhp
g+vf6UD4bBU4WJ2TKt0ajuryApGrD6fRKvq5YJMJrMf4ePpAepxeFdzEF/Nt5Mf5FraVjqqx33Oq
UPXlnJSh0dHy63He1pULfl4lyYjvnKdhQi+3FcmVTxCWbQrRRtMdO0ROSavXTowGqlN6F7ZpWWvJ
FzNcADIacwEmThM7kWILDHiv4S+7HgccSd7jEicZ7kSsPFLdkvgT0WSKD2JWbRE0YWUoDheeOwb3
Zf2m4fT8FF7blCy3r9fICUSoydGYdtLITp6lIAiXxYvRmymt+mK4trYtTW1diijFc+Vi/yi8BUdL
IBzVwVyYmEo5lo1nNujcOjanGcneiGnsvaUjADgeOIrjGRbh3pqi/qeAFTGVEhICeEMXnqfX6MgB
oNgXN2y9QohYMdH3kcoiwIPh/dWUUI60FFazWSVx+I/4XB0Oen4dY3vVorjTEzktsmptzQG4bIfo
mIakBMk2ao1gyOoZDD3fevIGG+N0+aUSgCD9ZEpkbYSGwhEPWEWCJnHvkaurns33VLeDvTg5+Ohe
SxPLgh3/ZnFCkUWP4D39wWUUTcV916LTZnTqs5sMG3XoY611SvPpMQR/BNx2N7cuLiM54ObX+97S
xH3pQuQAf4fJnHV8WOghkyjWQt0VwFNfUXTY8/lHXszhNV3yHi+3ygmCtq1tRGoqmAvlNtlWWyDs
fp1A5Y86zJIZKTY4RaAttKfEb1COTyXec8VZKfV94T0QK//p/gDcsD6cq0DfyiXnOXel++jNS2L9
NXR5pigXYBxug2LMrauPGgwrkrql/y0lhqqsDTgdBpuwlub54dCmvw2WkwIh54TXmgecvd22vKM3
JacRCQtM0NThazeNJzO1kiXKCFAZKerqp8sGK5ktZf3vJSTKCY6+AmMl97wS8Hv5bzin4RbUhQwq
FWxv/miIi1334zBMsTnkCbdx7HS7M6GlzFrpQP3vQlbEk9EvdmZqCESgbfzv1jTuH80odIwD5Qe/
D9wWupI2PjOrvQ+nHo763h9wSoBex7ZB00dSlnfbn2ZYujfDtdTAb+bGJbMsdewxpGZB2mtsvmIR
xb1VkTpNbVrHPL9p7igJKzzacPoRLegSQD9nNXhjudr6M3TGToqiNA8y4scV/S+RwvMqOh+V0/iL
/04tmJRsfyNLJNfb3BzPkPM4tyjmJSyvkA72LZGn52/SMsvdPpFow2LZoWQ66QNIUalxmRhxBWTQ
YcWZWknjJDet4d1WTx9oNAx78hL8c25mIYEuoqOZHIDg9rtVIJmnapy/A8k5WsE5H2tFLHuhCzYC
CVi/KcBPIZdMxluS7C2ez797onJKUo0hfYZEl8imfxdgXyqsZfiC7+HsaAGmWBnKFKoHUr06RU5N
I5dB7ZMne3SHlgwXGsFelNXmAoIOyOY8AikPh//e+Kllx/PoLSlxwduuvBqNcGtjTiJuthe1/1V9
tAiOQqebU4OFzISta9I8AdTYiVLdnNFhbsWNSVHG+bPWJxaA8ThmLQnpyWtMAGsAqL8uaVNl95vu
aGBJHY4PGhIl5MMdJMoawLYKvYzex8CZC3hbpnu7HFaQFXTyeiiJ7XvQj+tnEaU/auRfRYLMbAkF
pzYcpKgs3hwzxgPMr9Gx76nkaofHmLIo1Hdz6Bv6qKVAnY5e3c52an77B2ELu//g1Z0ooZsDGWeo
MZKdHdTY8slGd7IVjbTDmCc9hsNOYFZmNVzCapyKZFhXHl3PmMwbsCosebokMsC+PagBM+DImC8r
ZthEOqUg7XDhYmBrowzvhcvWzq0AMlmH7c9RsY7uQmDH31onEULCHNqaRdAPjIypMwjhJTJFVl9n
RWYxsmHRs6mW+U8gbmPy3GpS2Fpfnf1DSOvRaKjJ0fGEX6vu0R8Pnp8iklvIoEJrbhR6W6/xP8U/
kWA7gKiJ7wGioV/CBeDJO2sEsdJzd+//0XkG6lbe9m8FNxxJJ6hNyTZs+yXD748Go6h7Ze4sx525
cnHYmk5wpyDZXPS4W/GDCBMXqjNlyN2zletAfPreU+c5qLD56SyEMlC38R5XWRzdEuA7HcMM0rjf
U+vYU9Jp1644fMkPCYIgFZdJHhFDTeQVQQMGaQvkBbgEKnyvZa+OvENYGwvRtKVF47/pppYSUgsg
ifrl3XamDhpnkbiu0YqIMcZyyrCI+AWXtWBiIQ1QNMf6cqpEXjmJqsmB3DOmSQI8CdD0mU7gI/+/
Apg7b4cEZwnxG+kGqYEf7s8z9fqipml3GT0Z+hJabdCS5jc/RJK2linq/M4H4BnR+H2qiMjJ2ILE
7Z7Eb5E8wlkKvgsQS6uErRzujaBqgi16kzJ1PONlfTCFiLt1e62z+JgxkpMV5HuX2a8wC7oRYk8t
a7KEmSIIX+KRbasQQ4/gKC6JiH08k/q2DrLxl2nHsHiVDNF8K323iv1Cshm0CeBUUzZM0aQkb4rO
YYAfV9kbg3slI35qBtO+W7zD15aR6sYpjcrsauFDjrBruhtRpxsk+mI5Y83GKgdLinReZoGynJKK
XGEVlnpcDXBmvXhN8roqR9CL6AwIXV0bmASEX85jbGGCyLpG2hRy8b3Faxmrpc4V2Lrx1HhEpIeS
dlUjBQJMZVtH4pr9bKHC+VHkohhZjD5cUiBO9PwgEkKNSFOjoLeO0sdWrkSOngi4cqZ3eVVhOoG6
M8dRJqtuV8F+g944HQt++6bWyekv78mz1W17LOghj/LjJWxTq+3T+MrquAv4x/i+uVmTfmHyEjYt
TEEmd2MgbB0F1ZxI7MeetrDzQXTn23/a56MhzJS3CLqox41WU5X1Bi3ytxqwZxbSsBO1YHFZ3+5a
846X3FuJiYsRNni/9ea7CQIM/8ouol4NKo2hq8pZJR0PBu3N627eORgCWI1eAlxSe9nH+I2kIkyN
+fCrktYS8iZaRWHadBC4sI7ToPz7NSsTA/W8v/8hPrGQ218ODRE40U+FrTs0tugqjGzG26qZBx6W
/e7RRndEaP4nTY3jVydGNuXaDWkecLkR1sxKdbrDCNQW4mbIx33/lCncoUedNm3Q68mtLLVGo4jJ
eji7LfHBBib8z/nu/WzZzuOXcdP/2mIOHQiE7NeVIZzsBpzZ2fl9IWtMv7jgt4l9qvwwKf+nmCqx
9CgxcGtLtJcVu+GqKG9mSRCHdVNEKuz/Y44uo6TLQRjFf46PocB2llk6TOHpmWhuzSbApkIL90IX
V71a5m9QZlf2bBzXBZGQMQb3oHZOuDB56G5fSz3CnEJf4ilT8Zx0DonNO3D054utLi7xUWJN6RfC
CPV2QYxIHi8rA2qxvWs/mVYbcY/Ga9nayw7/0RCro3cLxnbu2X4Z/iwCZKG6qqdqGUDSflWchnph
CjlN959BdEBXq7klLImnYYhZupkAPRnwf4fXLxodq+CoHiHGHKKxpva+dUD0+bC8efiSXyWHv/hj
SkcBOrhuT7PmitlTRvXxyP7fegaWmr0PStMWAH+3tTt7wCH3pRW+DH1gK4mZh0d+GRrQaoRXF/e2
Ho3yHMmGQT3MK+wwmV5W2suWt0rLmp5OoygO6IuFApvdhFPn3V2Ork/8QgvbvBCrtZC2yIbZbTK8
LWvBNnSIUWUDt1glDp9nGG4I8hdBcuMRg5O0HYELHVJegnWWf75PRo33NjaUJ8jAEJMyhxfftJDq
KPpTfpNy6FjLVLCGsSg9wxi1/E1v/3Sdvc8kx7plJPfStRu8Z+YrNgD+BhTDjdwEg7t7mTFzNbn5
nIbXfVtPOnkOHBQQeDMpzzYE8ggNOgdhiU2RykkLiUSCV6cwrAl2txuThIBr9cCW7SunyVQN86jF
SEeVs37q4MnZZsEQuUTqRGp9c6n1uJ1RcLkHm5kh6Q9Rav9PqlUi2pGKp8e41JCMxkiFZYfUPMPg
bAgrHOYAcKgVVcWug7qyfEWJhRsKyI+KJY94aVTtZVU2ZjWYAuotVcc3cxPHPuYxi5bN0HTDnoBm
/FepuJb3b5lrqGCn9eRE/L5+Gk+qAj2SfLzSGB6QI8Zxg6cOkX3FVoIH/ELUM3AdoRf4PcZMO5MN
85pqU+ZJ+sItcWV/oD05ct7WK+O/GHm/mL3p+XC4SstCB37U4QtPLpMHX4KvfBndnqgUbOq/wH/T
2qKjRKmmDfKhu3zKjWwUWhL94E/rJzi+a4/eDiMWeo7pAgL9QnQvtHC1E20EYwaAD2SYWo5o/+VD
ZgerBfXCGOQdcmgRNK8GHo7RZbrVLVpHptPUkarMk5h/YNywZWQQ5riGSZwDztkTO6BL0FZcpJ0f
4M3+Fv8cnaNSmHttdjcQ5FFNTl4duQXhkcoLIxVJXchMpbt1Q3d5cZxwejwvkzRWsLTU+QMqAcIN
WS5MDw40lIcuAxr8cpqyqh4k1U/i2zMRNhqept0L9s8+NQHEp6/RA4DbkxBJAmYGWr0cFn1rdxP6
fuPzMbOWM5VU4BorOFPbzmGgbdWrSJmySqbNVDtW9Adnw7V7PH+cca10PGLXKpzishqV75L39oLX
7Funm4FINcNDr99Q05JvIY6g9dassVIlQuzDpDTniO3ALxLOPDJP2LQ7sU99uwx7oByKaTGh1XFp
/a/eV4c7KhV29ETK8k+yi/sX1FFPGGKPfacBgWR0HKu+P6FZW3OCrMX4JZZOR9DQLJDyQEj93FI4
7xWY/9hagjFz8Ky0aEtXcMg9HvseXWtD4yWHXv8mq6hP7MU5GfzdcgeNXQo2Hoka2sNDmOV0T3ty
wrPXnMJ8vwVp0S7Sv/gNbywQmF2GvR7Kejjd565C+bq+kkXAAAzgoqnIKiOKl0oHViWxRh0StWul
o47gkuW4J4vDO0LYzxcAL5Q8VI97/P44yLdnGksE2lISlB4DUEfy0sPjN6CQc45nTz9PJ/Gd6ikt
I2BLgKGIUMUNlNgGBct+lmyqVm/GlO0c93YzQot+sqYQDWUUyY9f37LvR70ACf++X2wupvPtoo+Z
xHj/FlAtLTR5qbZWZ0+oBATDNwi09SdRhMpW1LMXYM21e/pUTyr4tdpQsTu3JYKZT5bobB/ujTq6
OBU8w8oqmTPvVRXVxryuCcWpzBQo9cJgA4yQg4zH40FNvCDzbZO/a28Cs4TR1qv0vTl9OH3tiMJv
HNj7RIbEYXgDAMfwOtgWfl9a8IaKrmSGEJUocOqjQzY45uz6MkeRHPLL/v3RnayAWzTCcUnEb4Dy
vgj8nFxVIx5nuUJ9Px4U2zeGhFHVvgeNi1uF95K7jFZEHjLYDrp9BgnbUhp9bnjibWCHcNBSNarA
4f/7TkoTcnywc+n6tP6JATObUkePmWbohA7XhGpi4B4UYPpzEC49v1bgolCDl+mWl54kkLiFU0qP
zN6Lm7nhkwosKylUBdx54vr7zFkc1rxaROWPcQtUk+B4DIuuw7fQ48xUBLSPb2T5CO56fa6F0j9o
WYDi13S0MF1l2mGZx2EPe6LRaaMIhi2OGlb+UX/URXhZYuwA4264y7cG1LToYUKD+OVanGbIOSOE
fONtPfGEWCfA+R936SCFMhzcK+RSLA3N1eqdZavRsN0YhfSVxTAarqBOc+Iou7NbUktB9mb6MJVp
avg5roB2BGUeGW89l44MPkmVL/LVe3mIpqM0RqyKj/kxHttH6Q8Y2StMw63BJsmbjxCiR8z5BI6B
nGMc+qYpm78CF4ZYDcbQ5LGbBlHAkjsz4QeBk2/E7co3GSMbxLzNgDIvIi5AfGMst6uWqf1y/Ynr
1w5ZlDP0tb3BfJmGhJasCsy15zKowCdhqkPD4qYZkXlWptfp4rqDU21wl0GHktd5krYxRMTGeCWS
uduNGgAa+vLIaiA9uf7i0ALf61VPHQQqggSvZo+OHL36LvE485FaFyaWH4AcyMjfDTNoBsR2sJMG
aRmJN1HoyW99+qXP7NGiHcH3pK/p3Xfa1zM6ZzD3kPFhpoYyLDBq8rZyfGfqaGb0k4Rp+Engge6y
Aqj5pIaT0WDm1WO9P7yZsnHBYdUZ6UZEA1AhhSwAdf++KAkn2TkX51kNbsrJ/aSfqLYLACKqGM7V
mur8Tf4tzngGrqgU76cgny/fyVQVepAX1zKtAU+1x8qTvIlRps8+pIy/OS3Fh1mcWczWJhx0FxNo
HJ9hxNnOrna71QU9L/GXauW/w5DL5YpIXXUa11tnY3NJ9uLi6y5KIMVrMINmphiZNP/WrvAuKUJv
mKp4VFazcE4FE098mXAzIbVrHVlLvH8Sp5T4k9dMKEGPOW5kVxC9olZnIrO9Z4hZ39PYnrzQDoJ4
005tebPTw1P+Qnz5hR5xU2id8qaONLIUX4bW+cvCJ6TvGqK/1UVumVjb95nv/tDKDL3uo5FRnP/p
16O7fvlca3FKFBA1qxX0ccYkx4FkZRdP0klfWiDuOQWeldLsXDftHIffGzHumtbQLDoAErySgvU9
mPTiadEgPSbwkP+PSf4Gj1DOgIpFqayRDsrh7XjVrdveZFvlwLg5VWfwR6jvKxPOGqPu4yjj5DWO
ZhhKvwFdwXU9Q1Ef5tvFRS6RZDtdu4soVHhqn2nfgILiHU+v7/cLoGm2OFBfkeyos/ZkMyD2axpm
RCB/Bm5+SNU9OZbGjncFUTxChMUKZ3H0TBKYj2Tw2Vb3LdpmHw6AW3WHCiukLKcCuP8vUoiyEXYt
r5CMJTrZQcIRTluPy2tREnTEn4uosU3PU+51pMiqdZp+EyJDyGUGysDc/xaIjEb0NLl29KxiIdyM
H3869wRA/mg3AfdFrWhpOc0JMWGFYx7CAz/4bTzbFIWvGUCz/09/8jezEAQ5yx7/skNtZNH8JFin
lXFBrKFlsMPQlhC/DLN+SBMtCl2KEJudMEyDGPH3Oqu8GCX9iXWjMd5dOTzOAMzbmOWgzOtU8q7k
nLsPVI18vTpizp3CSZQ1L9ZqIV8zb1yGMOQgqInO9vmI9vWqmDVSbGqj85RgJRlYuq35iN7Vvy3Z
VnwWy9SH3nc51cmZNl4LaGcGV9O1L3KsPWAgqaYyWc9sq2XLczRNYnpdcXE02uMdbU5XnK8SGg/b
/El1GrSsyniXJUPbJYGixcKVywct14/xn2lzL5QIPLV1SoMUK9FhWqvQoZPA/muROTpEMxh8H2Cu
CwH4tsgCanMCW0aA0DqCFOEjLj38d4/GY6LSPXCl4ZC/DgKufoXcBbnlp2ZjOG+xFosjIJCssIxP
kwBYraaiKBBXjlYdLqvNR5Wv4IOGQ1++rbv9EN4gNzVafAv9LuHyOdktfNNJS/6B5n+3vga/8qnN
PE2xFHB1A9rDDcSGzKNnSYhlD8aOZdV1VMWHpaCHp+Y8m+Y2yV1wbXwJj7QlZ90CRtju0aU4Q86p
88qHWFuLVdxNFkYDMn5bQS+tTQTdgbMf9mRoqKkKjwGe7UyA2GVzR9MNBJcIcXFcfbduYkfN/OmU
0KfXeSKkhqgG1EHFD4xpIpkNu0bg0kEPto18TgVvidDl+6C6k1lFteqBjJnGtOV4diK3gkMgNyXy
6mtklC+CCQqArLF1fjwdtb0XWA2nSqwL2mWeQ08/v/kAWNhg2vbVlAIAK5J9NsYckzSEYtf5hSow
5KCrdWD3G5WvVsiIBjWKPz96lUsbzU2f/2sDnpIk9VpF2FZd2pxyn1DVYMYDok48n55/gx2Sni8T
UID8zkqXY2pHselOSwjsbwHjq6AkAg+637Ve4hRZcfHpiIe4fmjVvakz75mlloNUp2Rjlblk/YNZ
lUer68X/8NJs2UjbIzLHJArPNqy4xG0j4c9MQ03Hak5gUDkSPeQTOJo2YQue4wFVvTOPrndh5vLD
L4NfuTxbeO8iHw3FC3XjTbc5tKNUA1qK5ifwlfQoYR4gDyMTgxSnbxXmqddJG4BVDZa4yfp1RCqj
4XLLL9NMOp7ClHYLRESPhb2ac8Dtr804cPMYt96Ev+3Bi4SyNQaKG8EQ57/SRVwLEHeALcHEA1no
uAoDaSv0FQrYXrDmEThCbrE1rkoizA+OzsUU81jVaBqV3SMS5RJ0Sxzor3puPvWo4qr2bYW9il8C
psVqsuTVP1ofvQBLPYpY5v2fMFWlm5AOllKARpYZX3VhOXkpCx34PrLFMuxL/POeyaXyyfPv/Fwo
/P6CgKsrQYX0/BsjStLtVgYh+7zUjbgJjlHJivjJHGlzgNVNuTlm1J7vHeMtNdpPYvH2MlaDOlE9
ycdb8H8sOLafaKwUVysNWwazR/Vhvg/t7MAgnJTkaG2//D7dQTedlSDn9kRLTLuh6YJVTaotLcaC
tXaXMjqB/c9Wa2j2Hw4ZCboVr5mkk9+1cfwO0K9o85oRS96yXxmS2lRHWXSpqRq0XkvGpbyOpUKj
AiQ8rB1mPNUqHJSllFl+YVwy0CAd9VZjKmUzT0seaU7gEatCeJEzAjoTadDPeKYfju+J8GGfTpFl
10yhcdAiwUX8/g596CILBDPGRuj2NTMWEf4nfGLd/PSh5mdVI5JhT5aMO8gUwcmdRmPutfTTu1HJ
+ZwRMvV07TDSVI8Cw6e0sxlnhcl1gSeUfZh8siufovbCORs6AkFViJqMyCecm9tEjOKEybnptleF
VvNB0LPWJziu9twszzpdtRnQWEeQyWa79jWo2D48PoIPoPYnCUECN4irSNkUepo9FJXYvf9k6y4d
P71gXXK3OG0cWN+ygqz1fpVwYUagIm8X4JjgmZRhthhMcLWc3Z2Z2PV09tcw3WLmKIMyUZLLjvOP
1E20VmVdwvfamE+hMqNC0Ts+EcueWE9z4/5fGb0xaRn/X7WPEGeWhMhyDH0BQtqCpgpP2565A2Ix
XND5I6LnIZLZlpMB+2kngo1YlO6YAEDW65DQKCNc4aVaqnqrn5iq+g/pzv7RoznNq0Q5oG+NJTG9
hVkQuzlP0/dQDUEP/XEj5V58cL8f0FMDgNcVYf92fsuNZuLwQXqwCjK8wK9t1mM+pkXs0h4wCITv
TeGMCu2jeIO9tQcC0Rgt/JkvY9oDezsEG5eMz3O9Eii7XPf5iOv2WB+dnG7VQ8NV3URIzASsyRkk
3GQririTlZYmUyWnAkfhzWobJFl/mq13QQ56s2+OIwTrzpaIWexYYwgATzR2HsWRYGrMt3XHiZzP
RD8HT7JRuosF4viYrBYIIdfvTgVzz6+c/MAm+lMZndemTUQpLHKseCvpMmJjqwXvSjhcURHpKacC
t10467QAO+aYOPVldSyi8AlPg3H/H1DOMvABVLwO3OUe5E6y/uE2gWZr1qSUKrMWF69M3VY0wsFn
s6Lcs3lGfsi4EfbqsiGVIAhrLmkshFsip78CpRnxCMr6KSVoFU9cibq+fnFvIB0OrdJVtpbd8/M/
j+FNwcNQ2uUhFwgx7PcD7TD3dIcl01C0Sl/QjFBGwyIldCWG3vdPnV6M03T2hxAxbD6r136/Nvnt
cXI+aSk7sQsmSUsKpD0EHukZl83GXUD5oBVYRhubEyuVVZct9qb4tTAqa1b7n2EI4+87c2vW9yjU
0c7EC3KPiL5pkJ/D4KMwcEajwJWo+NwZ5eO1eyVbOzmXvfB8zasPhN1u/nEICtWgLKJf0ePwqM7a
xoRvYTOJR/GT4fnflXR9QquXhFpxQb2ozf1gb1Lc7Z47IeHCHmTmN/zN5ow37sK/qyLxQsBlWUjj
BnkgTTQ+AP3ESj3A5AANxWwXmz2im59Qdiz7Fm51KY6/bagu4j/1Y7Vofoake6keU2BYutaZtHJD
WE4uiNVGtjBbCFLkLmG1eUVqNs4ccjbYfLvVp1jY9dlLzs6edrM77BZE6vYTpumwR/n14jll0aWy
kCG1rPYATxDvbuaiXFeFfd3bsfcKZNhtwkP6qOx76jkdtOwxFzQ6K5e6yl1E3yrEbV39JkciJPPs
cSU3RBWU0LD5h68Q2WuHXmt8580VeMtjRfnzW6hydpyX9w8vfKz1Sp9MdirQ2tLAowFWPV6d0oh3
plK3ineCEx1j+iu53PMmG+Zl1u0+L7DDuSAqY1b0oY7HAWRy5XK58NE9sSOIIMTIizq5blWW6zYg
4yGEtvrj8xkrwmhon05m9GnWU7mw3ay6zu/a9hwYoAGsAxFGKlTg8YxNpS1rWfUh6rVlLymPcypy
NR0UTVLCxONxdPdN4iLTp2Vxfrf4ReKF60z66F73cYyneLahdmvX2c70+9hsxMMB3tp5a2gFiPej
sAskp7/pXughI9K/R9l8FuwyED00L3qAa+eowkBTD24509jDqjNl1feyz8zzE5Wm6NL0X2XsX+Xj
ZEM03sAcPNTmn5bz6kvTdH1Kw5r+UPAiD4YW+XJ71rtrEunCqao7q91BTfZSt2tBl3LLwG0Zvedw
0183mnd1ZyNKrN5jSGhsXZR71WL2rG5kU4rM7peF1kISusa7MmTDES2/LqkgYp5mnVo8IrZrPLyz
9bPOOuXWRXAsg7qerMv475HaubyRGGTcMgrUMVHfPSPRfrfUY1frHw+ujfvn5I6JDfM8mHFMAkE+
7WRngP3EBVaTWb914KupCZZGWUOXgXve0M+o+aL0GkvgWpy2bij2OF3X75S/BmcTzAiZJYzBGIcV
tJnrKjlhRDYHjsn45rO9YpbEDn2jDq+Wy8auND2i/mvVk9X6lM3nnDYFJ4qF7cxuQ7+LT7rmxKbN
641bXpuxQoC58+BRIuQwPCbaZ+Y/+ioO33NXCyikpi9Zd0G8oz1OJ3eqVSUtVDQCtHQO1F6OWYwR
OhpnpvxJ8+koUBTi0012qcrmu0S71QISoCrvFXOnK34PkqfYgeH1z9FSU6vqbb8ND9Kyvjg0AlhB
FFHKI1vHPrHJ8/AiMCcVwdE3E0y61JjyKQePba2imAm4O2Sfh7g18or4eW3NZZxJC4Z0ki89FayU
m74DssBOJ54Z1s4ejfIJZssZB6YGid03cF60flb60ggPsm73cSAZwx7o0GR3IdLTEAScywAQkU/s
l/isrnn1+JLJd3BJg+B1VxdHhEv91zfJoohCvX8Y4lZvi21KxBjXn2zN4S/o+I0iyebWsRDlbWeQ
bE9Jul9Ac7nk0W3Z0gMPoJ74NiWqNdfE53ZVDIpqeCZiVKYTI3NQrZEdwhxlAgTKsBcg+xd+nqZo
2FLPgfw8MtAYvxnb5BtASwjdX2ivwncWj7lERNoyMZK/bEQjabGd7dQ3LBilY043p746vka1+SYB
twfyH0PTCO0SrgS9GsPY8pXKYkEQf2VjyT2bYoL8sT5xVDrNcu73QyTz0sUpTDyzQgqI+gVm6jfA
zSv4iBG1Xwuk8UCdr0sRz0JhEuIYFSvdQsPkEueav0lOXCG3Q44dItF2MR4ozBA7hQoia+piCnaT
HH6jWmCDpCbLmK2Gq7SYa0Q6J8A3qYdRHB8pIEdlHuWI+ewTYDQYSPZAQBVNPY8bw1tgxBe1l7i2
24dvQTkIDezvPSjJ3iNdpYmLgyclDf1dVi2HcgZ51f6x25eyPikHz/Ap272euWY22lyejzuIY04Q
XtwnmqhrQDDIttXSytU0Fh1pBJ9C9EoMElJ7ZC9EbvyMLmSlA+1ThkoW05R/mMAOoacd6g6jo0Zp
buTHEqj6TS2EfQOHYmX8CZbA3wtwCIC7Qa4oO9qQI3RsHpeSBW6WC7pKDb0yq8Ih3ijtfDnwqqFr
AV9sVna24fRY8wnEsc5c0SQFu72Se/i91jtCsYsNyBD13ueMRfDoNxvh563iYAnRuN/0CEHRxV3T
FTcq8T/ZXNmomypGIDLBvqAMuNhaQhs8aL9LdqBc5JK9VkiSUS/iGnF/qfP2XCMBVK1bh/MDCbjR
qacCfmb+xbgCwc34UghQPG4CS+8eL31lz43fhEUyVdiXN/Y/qTmEpOspny8xF8T2cbdVty4XJaYT
Jmabn3EbUNvMNhONVk65ndqvYCdok0P5wPhOPYR6ONhVVn2Jlam6k11Hu2+oh/YzT35iEhmmlN6B
pzSm/HKm91puKMBTamiYQriAecnbaPZZH42pEluRl8VNAkSyzONc6mBAVQnEh8EzJO+KkFXHwMGD
9D5ruSFrp94fUCjzrcUX0+le41styUt/FWcNYbVHajWI2C/OCKQIiKtl6UH+0+7PtdDfep1/mPDc
xZ7p3d7hEFW2H/cafifuCcLYE78zAT77s0gq48UkfiQcBZ9lTe0Ahu9+b0lEtc9Kz7igPRsaCOf1
ieTNO5XQLl8XjnO6v1L5C80AvOl5MzZ7hbeYr/pIa2o9mduHYM6KoYVIsGnJN4VDteldJwUuZjzP
L8sWE4EX7xVVbM1wcJ6IN2ZY2CoJvt+PwWsjidfW+a8BF8fHV0dYIgBPAnm3KdlIB7y7Kr11e8/E
xp7A7xN+Mz9ohD3qonb4CxQbZh6Xi4VrFH3TKT/jHigOoiQMY6y1/9u2e8FfDuQdjFYCaZjSSPMg
yFlS8HBbd46R/V/uZ1EKNKZlNbbR8BOeuPx6an9CJ4ZHLCIEX/EmWVMV5GChAFw+mMIc0x0chrok
LasYaPvsV4kwkmIj6yohrkjTqqf2KSMDi5jLReeee4+ngcXbrRpngMo8tGAEYFX2efpENB/yM1G7
EpkWqpvsLPK7DiPIc0JSjbZUmA/D+4mHB1duSQkrA76epRoVFiT0ZUpwn704+FJDKvypUnGIIQTU
Q4++JkNvuvpIYbRlhRBmBYXHirwAbN54vfUx6EobGcNJVTODNtjGkMcq2/gcs2IdfqHDV29povTj
7kAmtS8tGzHJxGISuUWi2FiRCoyaCIQnU+fz/3fjJgtLeO9qYzf2KY3dTxYMT3T5g8mSIi2LtXwj
cf5pBXVZ9nUcYfVHYW7oW9oD7AmRbkPzCUCWqWHdFeeIlClNQZbqlVaz18yEuJkhyNzJGm3ethqP
GDhUIkzz2/yW7VSq98j1nVwtO88D12m9nVTiw1/wzRMwgotJl6mGNJr4j++ZDPa//p0+ka0JXcUw
tNAwsxylynLWhnLdTEqFzAjADBOtewZkADUCeOKAtEvHGMPpmG662ShKsGFgZXODjwT/GQAkFsR3
oyUPVdfwrIapucBy9Aejc2oxohborLrmCDT7ffpYGZSemkJpXkGGiey9gl5GBTQxjGxk7VY38Bxt
xRuMv9skIl/rmnw0Unn+aUljebGoLG1jRVab7j+nalj3utoqTP9eA4I1+hG6/5HaB72d7mIc8oiR
kCgTKOsQKfg0fxqmq9qkMlXAZI9rlzruUlOrRCrlM5BvBYlFJu85yw5op3goa2QRDdIvsXM5az7n
fe0GCWHjSrp2e++GjlfsH1BCG7tgY2u7ECI5owVaTyU/r7ZZt/nWOHZLJG1O+kvCvdnmXGFDBDaJ
C/Z24TAIvOffLN+CmJ7lWBGsNB3lUm8FWEuQaLYf3YXsvsi02t5QlUWBkDSGnu61opA1rqkK335T
Hfzup+Ot7fKeKNul/a/HnQBlWKumPxD2yYDY/ELqVDHWt3NVGO7bgly4zetlxkzUudZSGETy85nR
DBGg8oCNuc8p8nr4dqD+PfyQIXhK5r2dgL9MZkjopQsQsB24BpYVG0uwyNdESZcvp6bqsGOvV0OD
q/2v7gt69JiihLmjFL4ZsErqvD22YABB4U/LLl/cNdknr+41Vq8jIzgRyyY/i6VXJxH7yFyJRvaS
St9gM7CZXnadTBMtAXLMA+IQVD8TAvSQWBX04sdUxh8PNQn8rLWdULHPQPQu/nLfwI8RoohLtGuD
igBoaRcoybmionb5affFbGiVdIbHYjpM7uH/eIHRwVu5VcdKp2DF9LEJAGOCpc0TawXKwchWYEVL
ReAuZ+K4ZRniZKiv/MWj6tvXaslKLlmz4Eg1+CmvFMIiA9UAndS0ur59+AeAKshc0L6i3hMK4dea
mctWDd0456zkOFhB2GR7mB5NX1nO35yxrsfUelOdTpYJsSVds/RLqyZIAszQJl+vXZhkz03/TXiu
rcbnRDMGzHAyREC9tgc0RZRVPwnkG3wFLqiG9lqKMOzBYCa5qzdw/h6PAJC7ZGFtjKS4/XYmIPv0
C9QTZJarsNhERJt2/yOmSQHp8bixj713Iae0Ybq2FMlYIu6RqgdC/cgPwzAHvfqsYmQu2Oe45eay
VZVmzlBYFFMDf9pOby/9nCpuQ9jDR74z60C1eQF0E6sSaacY8TRbWT1YNsnObvg/JVybB3hxUnEA
N0/asRpyZdUPl0jww/CgdBps1sV2AVsU3/0qSNAxW3ymB9knlLAXm3SM2wCG+4qE9my/eu/hJqTv
mpyg4cYqtRPtkFSNwS6eX4nwXHY704lcp6wZ3Zr1fCKYM7WOf1vOSbp2v1fD+iZB7Njuq0vkxkc7
6fUO0itCw4l+F37/jlK53N+Bswjf0fdVG00LCNqu5nNb9hGeZP42Wl9mUI7ZOsfMbKTF/0HQ2b4Y
V0bLHRWLDrrWpqYEywvRz+6jb9X1cB463QAsAJv00AQQZ3vBC2MdU/SO3yOOT/zV2QZgmRGu5cdA
EnX1RyIapM/rZN+qsbf65CMnxVg9ckrZ9W70N6/e+eOXLkqPcfVVJ8l+VObIMmMEpuU/JmI8C1WR
b7A+SkVo8cck+hQVaDj3gNfg4zXekRtzdIltT3Y1FB2CVefGY3OhhC+Y9mvhsPgJpENZJLpRuki0
H/aunhD4OoXGzeJR2KZpj4qzyq3hmxPMJhb2KL5iDtv6OJOKbV/Qu7AZG5tOEJMYumGcBOEjUpAW
X1CyEaO1963AyzCZzPx6Ko/bCbzjV/PJkWNr3C8T/0ilwK/InZ0dXGS/wYhwouKfSU0j6dbC8fTx
BADGP+pTd/AAyg3sw4HNJFTmnnGlaNSqrjlMtIk8eWeZYHLiKW0PNp1BNipIfffdSb7vz9ZkGi1S
1xnU+b4Fd5X1blNN6PJ5SQcFq32nJuOaVTmarnEH7E3MalJ5vtktiG6SAsjgbGpc1oWa/ZYiXGc1
Ze3EtKU4howfA17PW3ibu/PWqgOeFIdUNbQPEIXcVHWx1hUi3nsCwOuyB6KcQ93KafuyAB+Wa1Eh
/tVsaWVVKYpgqvtFCAv0wctzpzmHXbYcoeXGMco6lGRgyxmtKJH946dIUMnhxMCoWAStzi2XP/sh
klq9cCTGd5I5LarD9Paz4XCfcAZas0MAE+exjasbdbWbPjg1n8jlElhms+WHijkG0fHGNLSsukps
qbbJZor1lJccy22orww1D6q7IURYDxDQHc1QsF8k8DbAT4JJnOOnGhCW2LD0Z2WwNzMuJy7lE/GV
iOVSVb1P2bm8CI+aPsq0uA/IxuACHCNgV3dvxZ98x1bqCQUQlkl7BOaf16KtLJRsgBHHYlHuNS55
wETI7l3FBgApgTgu4C1MbiVY5Np7ZJhGo0u6OBQ7TYkhvkIURqVdOcEiyFqTdgSsj2OOWHLAF5FC
gNsnYnnCjjh2uJxYkERIMQAes9A/L38bgD7G6o1vQ5P3gMUbR/NaLw4BK+Say0qPZezryUHV/Qxy
dkC7RNOUldpSQBanQKejzlbquAHmcdkYQedcNgG27D+mwJ8ftVbplJDxKD6lPlHmHhVfY1yDkA9V
ARHr4bq3zGnduE9R5D7BJwrfReAayAQGn3hj5Amiv7Xoj3mrKNhxUKs759mlvdYy/WDgVqGiDxb2
q+vWuyi9zbmAVHJ1piE5neyQbVomWYlEszU/21XfIexuSsuIelue6xac76uxawC2Bi7t8Wpy6hYl
T6Ls93Nvs8ooD9hOfoKglw2uQKSic2sF3U7AE/eLVtEUOLlP8TBl8m8Ywa8t/BpFgk1Uan2Igns/
jjouBtmNa5WRJtIDQVs/NlNkNeVT7vaexAPA36jPnLoV44+dieBpsAeRkZmqMDYszmsFiHa5A+NT
FgB65mUd8H9I7+QQoU5ktYs9WLM7o3aFcOUzU7t95m+pHzL6mABt15Zc9KZV/sKclT1ECcFBP/vz
eNsjFop84/vulhT5nik3bpHYBOjtLb1E5HDthH64jXAJMDptun7R1dtvpli9f3FI5sXgTItfxZ+6
355SRCaRNNA9NydqBf4EsqCRT36kZDpFQOUxDf9uVspKuSDELSObNXnfADV4ty9p+APXDOHaD3WX
gEh9cJxxf891WQ0HvFs1Tt/FxcRQz+pUZEA0Fa4PDveHHgeqyy9ZD7ZZyx8v/TBqpfkqqy47wrdt
jENazBx9E+iOAzUpKJEjseLSoUvqM0KoSuD5ntpmNtEhQMZa5G5f1GczICSwSR2qyPxG0qafEzPW
+10uWH1FvXPSEAfP7dqTN/+pjoKlvq+jVnd0AsX+8+DW/TmcZrj3TFhhwUc3AookvMi99ZSLvF4a
ONyv+qqFtqj0rn6E+OYYpQv+TzxT2Zx78SJ03h131M6eq1DLufgZGJ5X7N0ENYaFMms+Bh9Lip5t
z7YSD8VFUPLd8JCeP+4TQh3YjLRoM881AhUYXpPvJLAJasb3sSQ1+4kDdtoQk9mYbTI61DviaCoa
L0biHu6pzXBSjh9e2kDtANItqRwDsO5yG+ZyaGfgel6p3wMjI/b5QDuMBOb7UTSGiHmZCmDPtG+0
XwbvIopgWmG5XpnqFLQq+U9ZE+xaolOTKspZPniP7NMUhGn3g8vllwwpJLsu+L4blmPScPfLdHm/
VMwbRHid935EivZ+QBGNLb7YjoJuVS/LdVQ4rEbRmrlWRtrrjrzf7yaEWig9nmnAa0JJWLrCgVsY
B0yQ055WzB/HzzI1HxES/LciBpy79pVYV3H2OFHIjcKrjIZRCx8CYV8RZx8B7+YGotOUc2YmZC5D
1Hk77qyIMD99rPQtCjfQw+ZYanDoUgqhYJ3ZhcqahwGQUXIMJvRk0xw2+Ovv3QukjOstcRMml5nS
VA716azgh0aNJK7flf57uM9TPaR66Sv7VZwO+SWzbjRpR65pap+DD5iq371jqevSKvjCby4BPsRD
TlPkjGqfROK81zBcBWyd4IB4JBMlmhBJe8Hw/Q0+lRc/TCz+g9WhTXp+goWNdvbgoBbwYI0k5TeZ
HmYKEgPUttjtfZ2jYpapAJC431deuHj5swZg78MJRsRMm9J2NYuq/SUeAYccSvfiBRRnwkVK8aSI
tCCtMX+7OlWhRb3sROIbEBCe3GGhkUzQFK7r3ji9oX30LC5fStBVgXpIG5vAfqXsmH4ufN7RQ26D
XrTQVY+IGyyn0qV01k0sAASV0utmozwjrFY1ZPNWTZghf/6pwI9c4lRG83uVMuWaKjE1emMwH5eq
0PAmd6GLPxus7YmfG298NVgwxRAzKtHQLUP8S2S2onlhQORWfIMJmKv7gRIB3pnXCD1KHUXRQoVV
Ml2lexTNCShNGxldeOVhWhgSDUx77dvezi1rup746QzA1ab2fAe3/V2xQoCeWtcD5CPg1+5c4IdU
qk89f4vApNhdD4j8dZYH2m7sDf4MHJAl34+4EtSoxiu95FpqG7/CcMKEC1KOP3M+rvH6KHQgGRhz
8B5t5AoadOPr3KHeUSFe+bBA4bF79b0iZFpN48lt/RCZfGsMiD1J5DmiQin9+hcY0HG1YUYDTYxt
2SPXOJMhgc1oVPh/Tx6vw4esadC/MdV039tm9wWxUPrZBq8BMeEA6V78JiEy0CIYpdpAVZak0qGv
lpd2ZCQj9SdtPHM/9IXJTRbeszg4nx2oGCRU2f4kkdyg5Ln2z2bVPwqXrTrJZRfRoz/dLfFSB4bp
CbbwhkhXUEzhp0E2S9oglLxW7NhqOGPNEGd290dGc4VBj/TFEaRKzSLuVFQ10cvVR0bZnp3WMLvu
6R/47IsbRnJkX4jq5RRN6X6t02y29H/kOLkuoDDZ3amyh2y/0jlF02yhfBEChwU/UFfJsbUeCnJn
+ThCjElcwdhWLAzUAemxYcMKqsPIUqNExM7bTPz+5/U2nI5wwquG+a07B/+N78zBAYjMwgMvNQH7
ccAbKsTvOdxx0P50BtdzQDkQokI+p3m9QbHw4IhXMu0BA0J1uPwmR528sdGguh0n2zCA66oYEZDJ
WHWrMTglm46sfdCKC1Ipc0Lkkj0MZkwHyWlQfqu7cTEab2FimEstc4wqSBreJ2jDkIgMgvY5Bcgk
rUaiMBY9SlSdCYGIjFPkaCTYnbwXWfsazjzzUGiMJG42a7MnhoWYU+N8DcMGTjU6chGPb3BttNI4
5/eKvBT/1c5QLd9kZ8LpcBJJIkjbN8FOFCWTW9VQf0lVJIiLTKH9N1yZQsF4ViRb8XHXqGnSnLWO
IdyrdbrssgMEHIDKtMDLK3I2Yb2jumTwYcZefT0bTtI63OOe7mIUzk+23gL6yOc283/eJr/jF90/
PtMIXxBrAG3nkTDYOo2IzM8jMh4xxEFKjl9WhlUPfZtngmmwIoTMcYhftNmigvX91GEcqx0Nv978
zmCctWsVn1Y5U6ktBGsx0Rk0K72ll4XxE47OY3RiOXFugoTON++Qh5XmM6EtWq311/f8TZGwCkk2
Ju/06Ob6Eiyrs2jC/ITbURTC2CGmH2yMHnHfogwMzD6AHLeHCu+VUeGMDVvcbR0WEECZqqdfevU2
19p2kzDafIfKFcK4BEeMzpejnhRtJkXPN/Qtn/ScG+dlNTDCz4OPjKXqXvvvo701weTSgx7YK6o0
xn2+FD3Es7KdyrMLI1QMUzP6+pxXH/rM3N2i8oehYZtjekdfr1x5KMsJcM02vjD16KVnWn9Eyn0O
PJohIlBWaHBS7Rk6Gi3ren11IpjrQuJWxAm8ee9ZDJ7W8va/ogghZ594CQh6UF1ZFY9XUKRgizY9
rjHvKJACe9xu1yH+2cFRcx8M6Mc/2W3Tky8+tjNdq/azJt1nKBZpZiQa+a/FZsJlwSv/bikApDeL
IPXMQLlcv32z2LdDiaaTeYLpiQQLtcZRO5pw7/75ikA9TL7nrXixbEL9GCs0pAqMPSJ6gmdTLeWl
NxA/tLQkDEEbOImVCqvXTZ27WIqO0z5GUcgzvgA+m2bfa2YAB4EZ2NKQ560vuxEbYA/eS6h/NBMC
d0Dy8nF1s35Z9pdBV9Qf3tX93FYpADC7DmoGGK0oiSlrBUy60/O8dVIqezr2d/VIE1eoy2sgQEOd
GAswE35Qle6V2yom0FSzDJ1M0l9sWsa60OcBbvONHs0f4bHegrKKDuC6tZJaQO1lm1C/BX0v0JY8
9Sv/kfBdkERfo945GuyXjX4PH5Dk1QVUTTjAHYHE/x6RGCXbmY+g41VXvduvJmy8TpRF5JhdXFcV
Y5Up/HIx2WX89It6fgcnQaOV/I0GQA3kfOVW22AhYQMO/7lv15jzOleQ4pOxeYt2pu6QzWYAhHSe
o741cvW3PEWx7Tk45JRRbXXPJ8IbKglFqpTBzkUOS6ofi3tnHpaaW8qOIG+YrZaOs3GHCT3sgl6U
5JByRzAIlpAXkjS13ZF0ysQC+xIgbrIj9L3xlt+jjn/lIcWDdhqlMSDgOzLBLXrNCCHeGBcTpl/J
vAfj3rY2FqUD0RlqMLaiO7ud38pF1raj76INsgJ0li9pjYA+ReoQchs1PBo+R9GaXNQoTwYltuFi
An8uCSIerVS37dlCB2piTXfIX/BAPYQrmqQ7cCK3LA50VvPo9A3g3lK+eNMBKik1hVtr7F7C5ECP
uyti3njzKTlc+Afx8g+SuEfZhEYZX9Y7JGzVknWxrRPyRBdL2q/83ROu3AKwKdzN2vfPkMqFAzBF
ac8sx/RgdrwaBt8lolEJ4NJYbkdLN7LhFac4e5VR72aEC9kpHvWPYekcXMkn8cL5tsF30i5+xI5k
TYctU0wI2kdR0HEESMSU/pRBllzWSVoMdEWiTsE9qbsysoSsCxL8YzlxHvEfn1OTKSGu+3Nh8Q8j
IscjzCBPuJUMZDlasb62pCeVxhJJw1NRQKYkymjG4u2rebh8b/T2vtmuhwKzkzuE15g2F+vvW5jH
W571zpoi3bGBy76+6HpS7GqLOlMs7J1J+wVgSyxINWQgYUJ7EWQf+9ZeG5ICZyukbCnWAmd90HDS
8SWIOEJJAeCGvHYhYaPf6OGRjhM53VgNgnqvcZBh1oYEnrf6atfXyy5P5F2xxoXkuTLZnrMJIYFW
fL0pa2itUYQcLXoQML2gnVelxk/9NicSiQoC8LzKCsgsglD3th3KSzJLTXEI7YqUWCtHA4/1ze2h
dta2YXknMdJMvKfRHKU1+GI9eacoi5pFbicjBhpBfd+k7+5UwgFu4KXP4Zyk6+Tjq3fjPxAYQeQV
v3124Y9NDwnh6mfuFPgeffJzJgjlY7GRmP7XuVF1Ut/W+xvrCIt3h4511c0JgkJbyLN+Pckyz35C
aYEdhi78C1ri2utKGbgui1w6cPlMCWUjENBeWaeWO3goyNmFSGvJKoVFIg/4xJ4DUtuYUIG8+nzj
RGNnUfhRhnUPmcZeytVJ+erbg+L1cFaA/5qovLbJbScVJ5eO3IvAkiMY/iCZA4lJUFQ51+PTYHkW
K/XgXIBpOetYduP+4lRMlchDtVl1Cacc0tZjAnPbwGQ6FWTcbG6g5uRkgSgm/Z0Gc4Iby7A+D/Qp
J9y6EVv0L90n007OUi40PMZL3RgHz+EGdm1fDAZQBsSQqMKKBoYEPA6ZDrREDuN7GxgDBnn3rBkX
jC7hbKMBSoKVEN810cv56FaIiIpqcFFwBMs6ApE1yDpiNrPRtpKutyq97ETQem0xktdc1d6Q6RBs
7QNRQ8/1hkiFshp+TnDaLtGEX/8cOIJxSNSXWfkbVKNqolZWkraByk2nfueFa7Oz4/hXpBWs0bIG
PYhSGNvGemd0sZFypnwctF+1PbSJ5EljQBfRjiC8q7WMpaLCHF8n9hZi+OIK9vzN/ruW/ftm71S/
k5dblKPKpK+d5SKBOpfrwEWU4tUweExtJ4Dzm8f9nYD0xdDrV2/jXAc/gPqXkCSvWbGOkPgwsLHG
CHFPkZ8l/rHGMFTL+Wt9ZfNTEkJ7BePnFHLd73QpEkNfuCBlMdXOceo6UftpCYk/DuJxVqt+lgxP
ohkwSZJTAOMFFgXyZzLr/W74zDq6MG4ntubCT/a86fhF1sc+xoWk/oXmPFgYMDpL/MeI6ZBmu4rT
z+yt282V8yGuIO8YXCf0173GVk9lj1stDRrTWzKM9fwsdRtaAxgE7D5Bwq3JAP7wAPd/P54VU98P
R3aFXULbeLKXKBsUxwhRx56I02ac2QaGUngVEyCMyf9sa0ykNAFabdNS3GLUvWYb+WwmwCNKtIUP
5uR1mRaL8rBWxRxAErW3wIGY8zK03Kut5MdwfVkWBXPvv90lsO2OuRcYBa+93qynpI8DuQocM13l
iwHRUFEQl2FS2XI2Aol3CJCxl7YuqgdrMtHs6TK/0kcaqxZA8mEMnRfXFzD1kPE8Ft6lYHBYhPC8
7blRSfCD7eoD5Qc7KIEYkEox4PJGKoUesLenqF6kzZ96UBFN6Ea/qwhwAhmbcIiFZrz9a3bc0PKj
t8eWs7zKIsANV3hg4qy4VbZY+emkhc4tOLXBmAeJaQzaV71BQvfGs5tu3+2P6522IlIN9RymkF4u
/rkGqnGTC0py43todfunyP+0cpAeP4JvWEjZkhAzHp0bXeS8mfhJS/HNFapkqn1Rq/CHfGr9rO3i
ezYDFssCyaI55OiZdsV6XIa+y2fg07CzRg8+AzSngzQ2TzVSEfAb//E8RFYEg/YyneSEqbUaOgkU
Xt3aHwIvneD1BVRUYH9g6awC5LLGUFNrA1hcTGw8k4IGTVUq/olgi5jBvTWFObNJjvvzRJibWGes
wVTo/K1fwjTbiZ5hwWBmiqAMHPCR2bwlb98yGjuCGTsDwrDzFe4gGCFFd8o4mS2bpd/CwT38z0tZ
unSJlDPhFKhxC7D46A6ni29oumsDET3/Q3bNUp1rHnzojNozX8wzs+ZwOCCVwmoJUq5XGc/k0LPy
1x1cu8xFjjHieyTEdjrkGTpw6KJXdY3iJqm2JItNIbnwmnAdTAUxk4UnzUWI2kbIIXHr5uYoc3JT
go70WfJ00kTvj+bq2UiA6ex19wlFRaxSbl9/UdkeVFjYI7kD15Ku7E7KHYmYxtdevI4x8D9sSOeN
INXEDA3zusBJvUAReNP9eof679B5zt4gozaLWM1mb6lH8VXpmZ+3WvJP/VzcMvlPnRVMm/RCD9Or
Mo29UiHqyTYJBLXxIAIeYJ60oPtRvSg3dfCc9q3UC+4+xqOiFVFwAL72YgLlPCy6y5morrx2yub9
eNA7KodlvbccdHoInQcxfAPdx41nCstMRA0vdKBKrTGz+kADn7qfRutPV6KF3AReKAY9EhH0IykP
sqrDmHeM9ju9Y8q0OrPoY63Aunf33nL0rMvKuL2VVZnzClo1eetzpFzZCXwH6I0I71mG6X+F1Yxt
BoGOCbjFbSWiqawT38aRQMMY7Yl67AHH1RjyDxaNseziNrjIkIwllm2bEtiT5oKxiIwO5R6EHUnG
xXRCjoqLtt31zO9TVgv4JaDx0yGIboHJW49Ru6F/jqUJziOZhvMlrkmoa3hwktAx/+1fz3SCG5su
2J+ckkXp+DF7f+drcym8upN+NpVwcgaeFOjI6TtdGh/5YgZORBn+n1WVR/uyowYSqGAKgYR54Yeb
9oTHzlWVitHOgX3jvRxsvi/wHI9UOtoDONd3GNDp/ohgrpEtAPjaYiaXxiT4l6wE6KAjUIPpHckd
YOyg2OAx39dXaTDvos4lNnZV4dHp+odfAap0/Vo+LrZQuy9kSfNT2TyT6lQdzngbI2QfWuXVKy1/
F+5tg0K27CO6Kw7Cqf/Yk6MizIotpNOZRdQC7ZN3MQr5ClY1dy0FSSgGvqt9OeC+HwJvVFnljSt/
BXkt8KdZetk7/S3wj84osg6+ciX3dudTeQQAWqcfcnjDUI6TEg2q5Cr7U8p1UWcCCwD6pPUbf627
Q1etAYEak51TwHdLwVktayuYsIfcAXtazDARTwc9YyRtPtHruUQ9kCKg9pmXU+gLpcdYTF0vKz4C
qx/wornURLYXni7dReyMq+7LDGYRNMlkArBJvPUwIKVAU9loA5yKksZVUQgVFv4tTFzcU8baHJh/
/VJ9oijruCL3oLvYt5NUaky06uN0onZeFJ4EYlskq9xXS+oUfEASn0vUHJQITDl908oCDktA4ev5
ZltwMhUd3lqWTWtI1iGHoMmQUgXFDiQu1ImR4Ik53VMWsq94jM4VxvzSZD6MlsQLw2XtA60y55XF
2NfAmbZcBpfsVeDLUcdnsLI4kKVDh/kClWmb+CAEgUdjcVmQa5RIgEPPpdznndudTLamyWzRZDm0
cWuN0enxwOGY4kaW50RnVANYsXsNy9SHmMdChA0gd7Uo1eZCHYf5brDburxlBW5OgnNHbN6L8rgP
m1wsgNUWlk9nIu7Z2XOzq76DTS/unamlqKkS+Wyvf/RoXJmMdyicuJmFeFdwYvsbIX38zm//jgGq
FvOAjIKUUWF24l/v3glCEusktL7+Y86DIyTDsejMFaSNIKqH0Wd2bl7yZ//1ucM+8GuCc7RzjK29
K4Z1Op2V8WEjSSskQQh9NM5a2s8Dmr/RDAtQPs8QpNaWsIXvwSHoWhyHwBZyVSIdFuCSlgHYgmg6
E9hbhvFqc6K3IYQ4GZIVdG0+2kCCtPy4NBuG/aRpLYPVhftDWRJylOnT8t0NKZW8j+HfZGixM3Uh
iw+YOpttvfGNViBoJXtXxKdUEzMUVX7mtRuhrqLGAf9bOm5zMeuxaqlpvO7jZIFw1Arei68mLhFh
fynmLASQ4rpQyB8gRwcWkC0GxAZ/wPcX7rIDCJN7pWxaQlDkS/Rul1SFR/axD7VGk6CtWb7aSISB
bnI9PXrAbaFrQrcy/mxny8sh7pk64k/Rjazic9hJdCxWiNZwWbBVdiewDBAt2DM+car76umhO+Dv
J+tna/gzyX2p3MFR1zB43KlUA/N1j/nIdOXUuGd1v+mOA3DPZjUL+IKz64slTAphJl1erO4nkeMh
GUMBsAAQ7rWvb/TZRTvMturXVhVr8Epp7rW/iMR4i+V2yqNi7ZcYPiejhLOKsPWE7OpPsBGe6uNi
WpvsgBEaI9BLWf7ypcIYJy8ZGWLZClRsiR9cs/YGlsGWNSU5hMzC9PigQ0W+D5HX986RxITsAHoN
y6gTxSDLX7TCd98Wuo141ptT2+mtZRISVd1eRHaB1aFX3uX26wWKGFpBxdKBjqO2Dz2WxQIiNdSM
MQUUGpPrIxohf8Uq/sJ4yOeSpFrWjFrOz/ARDVniqZkgbKgVSmCbwbOz5uyPfef7EDjF+fDS6+Y9
QV0HzY7hxNQl1l8rXacmtlcyoRqAaJfuIc6JUBAu80mA1xXlJPn/uicBGSAgUt5j+lMPXjDsuMKv
7rtCsUlhYBI8j2nKDiwFb8HYB0GSEuPvmoQWWS4LYdYBP4Ei1ZgzZir+g1tvVMZZFlffV3q0+tbc
+aztIRDC2E+I+iOeYfiKqRjjbHnOBqfN6YYZa3PbHNAD7ebe1PrpEI68DmwWAJ54N5ErzCqRLojj
G60L72tiwdryUV29X2WOX5djcLvDkIw3bIY4EU7tx5vym2PU79LKpBgE42BYo1X+o3L70KV8T7Ql
FuVtzOM8Dh7GETAFSExgDY7tYB3PHuOyoLhtoPYyNhAsGTyvjWZsa5aJX5sqK1Z5bO25CXAUJPbX
qnr4m7UDUahl6x+azXlUwReM6580MT832yLe3t0wO47kO6uz5QZte2yrEoU96k4wplEmJV6r7ep7
j5G0a0/2KS9U4wmaYEJDAZeAX3Jm3JET/+P/lDUGRCFSPFw4frOGECMJl0vPE2Dh71KXipMZr9Qj
7gHWD39f4L4Raacia7TP4o5xXcAQWLVM7tg612p98k9wKXOW4VCA4Fl/sLsm9BT5AAvU8bksOrdM
iLage1vGAWtGc9Gb0fX/L7ifjYuHlxmYGtgVZUrtMda5vGd93fNNSHiApOfAyIjfXHfAylg2/OkQ
459QOL6pU/S+NiRJ95HnXiFvc5E4YBbnDMYjguCR+vGWL0sXC6xnNJ7IOluhn8jJIwDz2TQSQvA6
2CYqDiF9McK5Dwj4htx6VwBdbcWIyndvFkZT5tZzF7cqlUMEgg7iZMizDZ4V/+fEvuAo0zQ/w8E3
6XPju9W2m6cvubDm8VhLNfpjrqicaIswRLysTPP7+oPj/LFuyL9MV16ETXH627OfVUeh0606T0C8
nh5DBElGeu9M+yOcATJpGUKO5Kr1P4D0g3f6NYdknPvAuKECOFpZ4oDuAi1U7WyZ2IG9K5JEBz3w
jH2d2K7TkMcttwIttXab3aFz5od0vnAUcZ00nhbRyeVApFWDqYKuBjSf3VxQiWVTpTlSyE8c+zXB
j3e4evWS7KWbycfVKZQ532O9vd8My1//spCkeibgwFAlRoipP+mQy5NIbfpJEGpd6aZykIOEWcjd
EX3rU/Qq4ltZXyDyGPooZcaPTl4AMvv6Wm2Vvb4YtbM6aj2OVEhz78ecVJA4rOgtMHb17ciNQy/y
OZcx82f6utoKriz0PO4UlKi8XuuzuJvhsQQEOitK4ZCOYjI8RlfyB+3TxdfRBqxwUhkRF4cjduBj
h3iviOXH6QcgJmddUwFqx6vBUyySYlENdWYgotkP4Ol8ZqLpyk70EsaHwl1Dt3Bh875NRUmKApOa
EL3fS+pJRea2mFpoOD/FqsspNDAiPRm4t5AkY4kGcgfOrjYDCPhrlx/yYqpg9i7NKjDJG+x5xsLc
ZSg25+Do7KFvamhUWHS/qWRaoouL3cqh1nqnnnzGihzixKTeeYSZa4H2gdBqpCj83GodBvPPddo5
xfCLM5kzRkPKdK4wBxZtm+m+gfeHZjXrWJxX+FxwQ8pHGvkY+AW7gV3NZCWI7l8mo2ytOJkHykxV
9Z5zEP0HXolsDTBqKVI38PQ4NROrXqwAJemoGBha/VRYiA0D/8ma9Zi1RSGqNLK2rKVvW/KIqrT9
qxqxs+Cg44G3ww3U2dLaZHsgEgJbeE6ca/mgr4NTeVoj/raPrv+IdK7tOyXafRuZD4A4A3OvQO1p
zR3b5BT+PrBQyGV2ALsUd1jZIqGUoqD5srcTDxWwzFxg5Ae4JKcdgSLC0xqgfcHvq1/7YlQ9ZwnA
ErcHViL0i+B0a5GmxHm04IjB3LxxUDtvw3x27Q9VyP1+GEnqtlbdDWP3X9skpuGs05rNq6/3YGFZ
uwRjmOMdhc4aZSTM02m/B+27rFaJSeA0bmref4qeXjKqrAuqJS59+REo/syFNjtNQ127IId8NyBv
xuNTD10n+fcEa3/+xLveRk0H6oNT1/fnqnyB87rBS24PHT9wsEYRkuJGi8j2qqAUwHy9zcHIRyEF
zR/rYQt02zo7G7TNeXv7dq45rw9w58xHloGzh7LEavMDgUw8/KwRsE3FawCfxBXftptaPVQ4RaG8
IWlMqJ2egjHMT6TDEuEiKsHfsHZq+XyVMX0+p8rAsEfxj8DsDJY2OUcKoy5fsXGM90Tm99F4iv2+
2g0f7ksnTN7Xcf5HItJ/SHH/jMs3PFSGv5B/kUQympYnv/NcD5Vm7J0qATcKZX+3rp6jMRh3z9Bk
+QRR1kRTLI45VLTI+SrcXktZ+C4KIUbfyqHYjPHNaYQB/yXhYv8J6kANYDe5+ZXycWKDb3L1NCnS
1deEfLnDcAomjSrKndzt3cQxxOZyPuR3o6+bVzAI+OHWR1pv78dcWLiji33UHrq19bEQ2jhkraZS
deM1ev/pRxzyjvJqsWx+unN5CxcBTO09CUgZp7v+OLCosR9iLOOsveo0VFu0U4xyQL5s7FGx2+na
rThAL4Jrk9l8rYR6wVm1kA1QpgUsvq/jHNyT1K2ps2SBNsrDtg9TvyNVNhuBaSeW9IQA3lkHFqkp
Atd4DkdJ7zKDbcj3aLD15OeOCmrciH3lwWJ/HGHwsFnpz3gOGoXI5S5trfLOUYUoXSno44b69/8M
VbDK/aeCWxlHdZGoxZVwv6VnwZgwn4YNykmcwSTRlm7Z0s29e8+tPflgW0SC39XAbLGsgXbwBsWi
6nCbW646PgYowFNq5rUGvfysXO9th0zPrWQXrB5DH2ZPjBASa2XcCUWlG9bGFuM2uQHp/O/wbrv0
YS5fd4O+ghOybUnbVqOClwEhDWSyMVtnCbyZwv6Wrk2Z88JUe4buMq5JVyJzoriabsjiT89M89a2
CK+5i5/Tit0J1dgiAfExojlNUTF32UzCPIWM7EBWoFYOcBM+8NwP3e5AVPACaAQA91g5byzYd9Vn
B/bSyhyFb13BPtkPfQb/Fyqp5t2Hn4dwgoCeBOYymmiaUzK46A8d/LnFN6RgGZPV9yT2YvinZhZO
PFxA8mDTtOs/Br8EkiXjQ/fLuTovNidfXC6MBno4/8Q5veq16Z0pJyEow51JjgJIyPFLVEI/pyUR
W1CzstlYHT/wUUp5ynMNYu8kWO+dkgF1oB33w40564BzBPx32Mqk6Kf85tcOZXqnAtvI+iw9B9td
6j7uK3AXw7IxE9HSgEHd4VKZfX++Jz28qxHJairsaUHz47B/7IoRaPcJoaMT+l0kx0dUE2TmdPFw
NDpAO1vpj71ThKeZ9btbvYbZCOeHUa7/o7RE9C2NQXzLXAh78UZ7lsIhhR0PFDR8JdH9jC/EfOfD
cxai8rxVs1gX9hzNk4gWTj0kW91tdd6ihSEhNZro8rbRRsVofTWN3nGq2J61+HNA00VpBG/Ix5f9
HWBwP7+k86dm8iNeJvZJU+QWYjXtDyM+HQHSFC1N7Zxm5gw7WyWkV73eECGy6Wco/vqji66Zq2Md
Gg+qBpoF3rj7O9frs8Uqcb+FTy5YIveeJ8d3RQh2HZruRZJi2SF7kyNmboMac/dGxd5vwO57IEtW
76CWhUStsiGN7zO2asALbP/ajwXHFhOwqzeQ63Bi1oYlRFdAN9VfTUl/eQ4b+XI8aWjv5WTIPlPO
ACcFYBCj5OqqCfhE0WuYlF4hQcsMLQTOgoILwZNwfoDVt5EOIv3/eFBUlyhJMBxOW5f3ZZzDbl7A
96htD+pbLsoJt6LW7uiG66i2HUTvG194umGB0sg2HY5FWHKYacWQzmHbhNQAMTXe4DvSTyKEusFQ
kkBsCE+6tLeKZ5Op1br51zRbrtr97vfSpTtt5Cgrmak2H+pHiFPYyVXnKRvn7fpFjGUm/Q8okjJI
srMnQ4a0azHvMg0skeqzxcI/La+zK78zwc4SRg1eMj5scgmF15bboiuMJiai3telPWLeMRdmcuEa
QjiADaCgczN7bgV36oHMT/IihkK1sQYKGOc97Zbm7wtTHcRb5UJ+kZr6NFpg8R3skA5w3kUHpyBy
VkiJ90tGcmRyn8L7mPDdtSUi2E7XNMPChYeYsoK+RIA5RuQgVZdf/BNhJc8lB3YJhx8NJt0lL6cn
VgAhv8Jra9d9O2Ih9dSjkOITWj5qdMQVZeVPdZRKZp/0O1ibfRERxBCOcclYtbXh1FCkkLqzmoXV
cRJahxz/0m/GH3rxgV56mzhuAUDnFpXmN1/b2y4L9mynqCbz5zePLWOlzRRDnZw9L+gHp91zmXUj
tPsqrAkPa5LLlFaiefopArqulP8azYxlQ+1g83sAl0t0f+DvvdUhWCNhCDtPM162PWq5cz/JlWGj
z7zjsrYHFdPX4ZgxNTmIJp/MzWfE7sGnN3wv87N4JfGjn6cXfHVwszsmwJPfPkOCV1inwfg/soHs
CJS/f5R5pbiP2iL5pTM8v+A9pmjOIl0sTQgqwLLhaRlXqVQj2/rhZ1Sapf48uI3cWcXtGwk+St61
pl16LuRIL5W0cOQBeuHQCef3i70ZN8n9to5FK+aoh9m4+CjlHCKODVk6ueaCdv4kwYvcfOfV0GYE
ZOkMvKkqlufSBQXzyIpI0/vW8sMGvraHqaJFm0W0y49FZa2dNnWEILJhisrRyUP9CSi8JBIEFz7O
GX/uirWPheCmq8++VBFifxpDovLaNSLmXzMiT+8jMDxrB5Krc6ODdgx33z+alsdxNCwlMNzksV2j
a5c+BDAYGEalWQrfN3LnDMMYcXjum3k1rQy/0ZZMpbeeNqZPN8sMBwV1R101iWDW5zQKOlN4MHay
/YTjW8FGOgpGvkUrHjAiecskOn74G/FTDosSc7gdTSCQljJJDTmjXQiedRmEQzz4HZAB+7yPubio
ezjCftVk26uuIplOnrHJbl6IzJiY37p5XIB+L/5dW0shsFWSR/MBxXkta0czLUGST578MC/FdGYK
I5q9a72EzPaSjeN4PGV2fNnow2xN7DV0V1kQax/A6W0PwxKzNeuB6Xf1PXqQNZhclRSwrHYFMabh
lN1P2awCsOBMW+Pv6fkzwcuVzsopPHAinqwMLATE6mvUCLHhkcKXN6/YF7Imxft+m/y42J9cWplU
8QMG3KGcbiEna80mVvnOeYXe7jZLL9uYI5R4IZQhB3c0SEFvpBjHi4v+Ch2E0mZRNOY0LEypE4YX
9WHSwowkVZBYL8SgOPIr16fmwLyhcLnxeRzW4YmsNANuYxvLJxYbHwKy+tPzRFyp9YckFd3p+DNr
PHF+GIRfsYjt3f6LExj+F7z5MPT8Hho6NTmw1nKFb5ds+R2ztD6ne5ajSuLsu1O9JCoYrjEIr7SE
Y7EuriT+Dvf70RvaCG4ELTUxxd3PRInFmI0GnRPwqUyy1TwpWF01b9GhOcGy4/ehmRMMti9UuPud
yWq2gELi4qT6TM/ib4wET3UczVRlP9OueBLPe7NG3ZY4SG4LLzTbva4UiM4EwDDZoev1z0X8qu+z
B7/IFeGGV+jDuXWh9wLWNCS1djwCg+vRoW4/8/SqMPihWnWnYxW5Nd4JHruLz5L65aUUX1SaKpGG
p5owI4UnFlJ7b6NLCl1L9G1avl3NberV+FPvCVil083ffdbB0aWcox8f9moWmJ7sNlNNxH9J1X7g
UnOHMmxw0KLnfA5y5xXyRZy/ppCW7KFHUJ02F89v6rQ5HCihPAFhG128+88qHJEjMuXWKcMAyQwi
g6iuj5eZFB0QM/cnF300cgQKJFZ+9OKkzNqIFY6pf+I2lJdVZfaB9i3xoNgjtngFD5zQwEcMhVfw
0cJTuILYp7+hqBbcp67mT9LWoz88PY4suB62ybH6KRd9BW9vpe26f0nn7cQdSEwJAkHM1FtwGl/l
yUoo/ewwDDh8pt+6Sb8iLQLRiLf8nmB+DnS+hbSUMtiGvvKCo8Zq0quskgVqp9huKOnM04/Qj15+
LXq+2Y+7Cb5ENvn+uft4kJlftKEBEvr5fsavvl4aPGPpWX4nF736CKmYziDccExZbv/G1mjUbPLf
IeKR7mYFrZhAxG54u2HsFrvwFWwfiUGv5SoyMcaqJKQMshhJEev51w+mrwAtqJn3EO3M8L15Z7En
P/vh3ITfO89sR2OznIBxU/NpjHS4wNvzu1iF+TEAEJV9n/aeRe12jwnkDV07d5fuZu/IcakCoOMf
YJxprL75HHlEDtxF2FuCXyiMSw6ViBUlljWImLN65aGcGnQ1nDJjqlDzDROwELMtyjDVM78w3KUF
+7JFDlMzta+p3iK86BdNbzrhci/RRz8rDrHQd804C08LDQxLh89Mv2sd9WWRvpHjM1raReh4qY9S
bRc+rn4ZrU5P3qYskGC1WQ5tfUZYysCAA2lOnlBZCVbFPDKKILLOhdJ9hrk7fEP7isbjlZ81fUbo
A76H9Z2ftvKI+l9oPq7+LM7yd0jcOwlVqsclROtAxFB+rck2tHS5ZXk6eOllqMSgAIv9aakrdly6
rA9w+XgjPNrtnZ1P8RjdEZVLHUlPlg+KTTyn/r8ifC1YfpoumvRNQOkE0TEzEvs9lw14270QDuuA
BNk8zzPOHDZakAvR6RZxhqbwmJgPgAJ3fm2LMyc0xa0EPQNIuvrN5ToEkeRfW0+fXM4y4jJxe+96
XXLfw5y+I8mv1BpLRKCm0HBIjYcM5akZ+ylFTq87uI9OQS0if9XHIWWLwMzYR0RjN51TFJFFnMS+
suFdSSHIRbHdQMVbjAZR2E0nsfNDo83bImDxmZbqyb/iFHhYmB6O5kpCUqXPmBMxNlEFtY8lqRXv
IJoKYRrZMjylKdXROg/+cg1bBzRuaYDWL09wXPzJ7TGxX8j5leAMd+vkowvgs5hlh5qtgy319sy/
ng7MVXoaWeScUYO7Cwc/88Aw1VlwPzZTQWI8n72Up95Mk1Aimj/2ECLpwuct4Qt7BSaDBjf9YdVC
wpFrZxR6662YBf6G2KM6uluNg+k2DG0NH0skclaBLn7wKSTocwcnnyehI15h9RaBF5bCvlJtBVeu
V+vVmsUCp8D0BGtCFz/Re10VPKqNPXzWAPRbzRAWhYEuuoS27/nHphT+KffcEunixE8FNSxsAset
8CpG23k1+F2CHjBm/rUkBS0Zc+EupD63GL7uAYVFKHKytwT537m96sIs7adUIT/jXudATYHYof3w
1KfnK1lTdyZnFUCSgvHxkl1FI59ABkl29hY7gYvDnsaPxpItQR2ctnoGbL+Jt+frQ2kKGSPBF5Wr
UxYNwzvl1ZFyp1cYqXWEfNTcjnBI14uOqFYkWTeT+oySjDt/LhVZtatX3+LGP3wNUYwCA2heT0IF
szlh7FxfVgyEBRdw7uipRH8ZuF35HbrBE82dlYQPZvMJnHdIGG335VmzBz4SkU4i5KCIJg1xDDLU
GlV1CbpLwP4NUyXqrbXWzSAVN0E0qEW8tnJlyn2dX+FDvzUn4FXizxA7b3S67FcMtgA3Rr5n/e/f
Ez/EFUHDBppCpWiXlrBMS2Ms0qlECgQQrrWObLtiF/Xl1FKC952PGk3tHx9iciEdoHGcpGfm+mFC
z9+LiJLfUyT2dUtc29yNMUb/Y5UlhQ/LjOClqHSRCGGZxAF27y5VAzFEsHJZV6SBgYqtLO3QiLoM
dSIlwaxAlPUYL6YnfeeAc9xgo5pXWaX7R0rOeBVyRDM/TxkMA5Sx/8+3GPzKoX/sBBAyPHvw/6bl
b9fG585ZO4lY5+RmW9CDQB6byM2KvgSTG+R+vfFsxeao/o88/grS7TKRzb3HBE3YOmGReTKHy0Ts
ivJIFgevRm80CqrTW0HWsWZY4Ty9rRAI53hkJhpMsSn8oJrIzYDCVdIzwk3xZkVtuK5rB9TuedPC
dkFRcOZJhWzhP6UF9+n8xPoksKtpUf4nnWrhmPNQfn3ywNg/5r+FqwF03uU+PjjdQRTxGBL5bBQR
aqVr+Guw7m6u2uxvrekxu1WDtz9WRXVch3J9Y6cJ2NyvkODdoThY+GKnK2vAfkrI4l4UBidtmpJU
oHLMHhf7pFzdY/ZfjpjidZbaGq8Acpzwm7P2/3BU7aQfQ7HBKtSNru3gD9dP331JROHbzThy1hIu
jYE57eWfDKGRsbgn0xE+hGIYC9mavytfQuhIjKabS06xZ2CJFJmGCI0G2CrYOXXChlS92MgKAmvE
WVVSro1HIQ4jjS7s1RiGqnkYPY+Y8QZ9eO2vlXL/FSUNMrfRxnG7hihqGC2q7L1m4mDMVKA4Fj5F
gzB/4zjH5RFxJiS81qvu/6sWPoEF9izBDwF7Vfd5iLKRvyCsp1yMO9hxD4Z7Y3RJ4wVocJNTJmNq
IQ6HD1ba78UeF3NuX/jqy7eGrBb6mKG9Xg9Zl5kCwGXWUwX622WjSU6RaXgQPwHS19fKxvZqdL0G
AOP+H/ANyk4FgBfDWTb7hVektw4KD/TMTLte5uyV0hMwCJ9JatqVnruePFColxNRsrmYDqrvSdpn
GXom9SdOEwZ/NuklXhRuc+yWnSsZIf/l7KY/Db6DEo/Bs5gKekN44Np/FBp2sM3lMHjhHjwRhDIx
tv0IkV+MkSnMShaxI05EX3ZfWl2vH+CgzcbbDxk8jD7nqEwZVv0k6vErcGIo8oR0imtoEdN6vFRs
UtZQRgqsQoOXSK9KhfbOgyirJY1OE4k4LltdFbo6iLjtFSkmJgLHIrouOz2CAH7vaWGACqEOooLw
S9XNYNTX8lXH0Z7kck5OC4Mlp6g6mN7Ql+MxJTRn8LiJpHQPnVvnR9nkBqOWwRrWyyvNRgUP2d9E
TzWWLU5Dlmc/WaDZdMZg7ENkm/yFCRP+cpBk4CBstCoB6b/nr+vGcmES4+VuZDrQdKrTKcy+PIRu
xgUND/KrXLEoPjIHWjQn66Eas5FAekCyu76AYrHzBmJAf+sZ0H2gRy7ogG0rxBLx740MYkyrinUy
rRa7wrwWX1oS9dPZEpD+DcpzYDaClpg64DFZcJu0V9h1FVv5fg9AqtkJQ/DsNPBOCMLJhD/UyHSv
EOL1E3g70lYW05w8qrCLZUxhwUBRiojhZLN1PXyPmlum2K1iMNvkfhbrGtociUv0+lIvt0e2RL76
G4N+FjTpvcp2YuhXljeHzm1R85LtNmDjM42WVYYc9AjuTpcribxDztgfQKnasZfxyYChL3vWdNPs
9FlfIFsbgy59SNxzsIn//rjyIZGo2pVEmCcj+tNFrv5gXcTwBix/FvjPJA/CQCItJcqI2uaYlWhE
7DdwxIbhmFBsPsLvcr1EQhwAeImDCJlf0eIBXvB52USsn8I24FpBOjzPrzuRc1GqHJaQTV4SYcfB
0/SrBhzcCRbkXAN5PSw/wo77K1dIoUx/2PrAinQvVtwoQn5LenjjqrwA4j18bQYpN0HJqbXtcaSM
xENrTti9tvrxSMLM1snJn1sscHaY3ppcrzABFxmkQTXX/lk1qPN7FbbzaShQ5q1TYpkSTf5VLlA4
IOrjQ23viZ/AzVJwbzpkFZENQcIhnSXQsdz0pIluTyF/4dDWrmk+lcFICFqLTHxBQR7pFJzZzHAj
LZhukpKaKJjmus1WnbuC5TpCcHlDS/gAd/uZYzr4hpo5qkzKEFJaFhRM0I77QJ9LYjADLMtGClxE
P1kaaWcZCYAOrg743A2R7o1o0SMhmC2mwgv6uqM3oLTOwwSK/Ru5duke3+8+zWpNnbLRdGambPV7
BWPVNNk9mD4+LFBq9OQ7syi9Hw0IO9WNEntOQbw3U7Exwn2hr/h+C7AcPwiS/7tKMA6pBjELtN6B
lHAbY4rc45f5w6A001XjfjJVlC7gLmrdErbx+MjQK8GdZ0XAwJLxjghGW8LnN3IJRvb7nXC0zTFu
opR/J8I6FfAkEXOvadhnTrzgiwFHnnXtwOQ9RqTkj49HZrqpGPu31GEHHGPvBfK2YK8FjR9Q5WV4
rVB7CtTF4lHN3MBPN0k5ehKqLeYnkgfbGBq7+JklyKPaV5N7srYx2Q4NiJep2hvIgjYihKJdtFNr
tfz6/19sshsJvpksnBekH0xVipatRSnUAMlPKNDr4aFfBsSlQ6M0lxVEoCW6Jh6qax0aVZRcHUkC
Tb0TOwwpRkAec9Fr7auFCQgVMBgLzx2+EcVA0keXayl30x5oipH8lr0xhg0GmHhrWSFyb6cxtykU
+oo+m61Qh8nLH6I7UjhnuBR4K/FvnyYZr1aIyizCLM+NgUcv3z+0+CwVhvt0JlOZ8Tfz8yudavdN
g5MHuZlSpAkFPwsDKh2n0YSDkST6yqoEQi/c+YVCpOoXQEdfVJkU1l/xiq3qLSwu8zW+ubDC3XIi
PkWLa3VsPR9cmxIG9TT0VqDCwrvT0uPhF/kr6oM1cpB0Gj8zYHqITTGfZEWIIivIrHoNO2t05n4d
45KTCiTtDaoTbpyOr6UCTejOTWJ2n5/SrKTdwIjnxatHVo2/qoO9Yzgzs2xD2UTsdPjzl9WTrLrg
1HnJKeXlpnp0X5vaiwJ2FO0HDBU734ADGnGJhbhBZ3HJ8zwg+n1EgwrFc11fAVELctmhXurUcGYf
TFOr8dRFDzbY9KMD8Dp+Ezvmpf2OvXh1rTzipt2SLtRt+Cc0+MVjB7DMNNznhtxQsKvTxMrpNtlK
xsPwz7pyhZtDtiAf+htFjPZ/dc/VA78ysY72t/bIrujIEaluT0X59dATdLWauttxssfrrYqckbjd
kORM9H/nq/N5Mrsg1uk5+xhErldepA0qEJpOv10sGzTUy3/yYWASaHtEYF0YwsFMwVf7Svbj9tpb
UJl96BYwsKFEJJZN/atNgPe0GD/Z62SXNR4jtgv4Xz263hEyToTzBTrU3tvmLDjmWwuLmRURKhg6
a0lmHFB7o5Jkkp0cPfjLWANejQPZ7TpZNCNJyHWf+OtgdWk80gOMPek26QT2yrVahoxV/tpkTWR5
XKGrBMMmpddx4vcWedrWob5ouP6eEhbzS/FSVx7l45wqjmuGZqtjo7ltpBurT+hbhQK9Fu7h/8Br
uziWwBJJ8D/Nudcto26TinmCcRORsghX4B9dMC6FhCdygpTu6iUKmWAPEVySoHs5yoTPsBKurAfl
1t0ZRA3MvgjKGbqm2IsnXps8l7Ya8Gho+2DAspmXKTMUD7XMHLbwVPH1gLqnUZlpKSfwYTUEfw3a
h7nH6WMYj86bKM/GwvFxbodABmvtzSl8DAKSvsxDUWLUGG3mA8wom6enIViTC/ICF8OoqcSLDCPz
HtrTXbHxXCEUgC4PbqGnI4a9aQg4PkwuFf1tklxg+ethvD5Vyq4SWVbx6Y53Wb/qA18TVG90V+jc
v7GdYe3iARRpANltXoGqbw2Q3Aws0aFzWTpp1H3TfA7KjgsHpZrw+vbJHVEBuVBuRXg3NL6iywH+
HY2NYjPT1Je++uvQjKlvavG2pdZV8qdmQL94K3ACICfo/v/yMGc1EyJ/c8HMNBXjYZ66qxnLMiXv
d8SUqtTuC54vTUpA9hLkZTxvpm2UqcAZsnJ2yeKlWCpOsRyevuvSJNWRbyNjveknrO8tsy9bCWEH
JU+vfwUfQ/105O1EZa5PkZMA7ON4/K7Q9Ud4Fr/dubnV6cfIkej0r0Jvr7+G1VjeiXWL7R65usM2
4FDlq6SIUIlgoLj1+il8wvej8laY1ErziPclHCqkpbnAnHEhCNjUapFmNHAXKN4raJok31EKTo4E
0oWj4cOEosXTyQOHkd3Eur6lafPHCaEDFaoTrAvzJGPMpkAWYKVLA9mPTUSQSy/WHWvHQQqV/inj
IZhWnUix6SHBhV/U/sGUlK0z9wFcPyApfhk3wSvTCr0SMIycQ4MtC9vC5XPtjF4nRvrpgoqw0/oT
NBnF8VlI+3zngjj4Jif7uZM03wz3YauU5c23dwYm0/2zsHAtodst88jlgpQocRyZkHN3qVTH6QLw
0pBy7xBj0DoYONRdgUfLsyWTlYtKbp4+L+5elcuNl67sTO0B5K2rPcrn802r9HVxzotvo7/R+hCQ
mnTcWdEYHQAXK+5pl2vqo12dzrW3XFoAa7/sobWd0BmzTzrt34t5Bs/lfsSYs47dqNL1et0EvLwE
joEx7VAzS7pFgbDo9k696v0n+kvHalu/mfohKLmoqX+hHpTPFljPCYWDwQ96gp1yEmr+bo5eWUN8
2O9TOMpWkCOM5W9loWU8wTz22kmc3+hGRb0BMdWEe7crAsKHWWJlb8HHLy/1hb2K5YOsUoL0QXJl
1VdWeK072ZxI9Bmk4+xkDYK5+b6mDRAgQsS3h/CR+QfD84pCFCVeW8BG7Icvmm5YcXQUI58ha3jv
GBfto5G3eJz9iz4hup7ihUrg0QD4br5Vhst3nqttG3cHzyOnpES8wMEizkAElS4T56alqxbqns1p
WyhBlbJklpcEpYpHLtB+lTtRHacYvt4rglC9DucWvDIMmjj1YFEbMUfXGA37Kg7Cfehhv6QH9uBu
3PAGwo4GPKSZP5w6pu5er6m2W1fhfTpmIHyzPZulDqERqm2A7fiWYLrRetppXUMwLb6n/1C9vcrk
BgdnEeq5JEhuXem1KFGgHCb0ApWzFZaOUNrgv5L8rdRldLsGlTGvUrfRAtd4Iu2scjpCUr/njm9U
aonut96Oi3dpC0SlzaWroOHfd7vHS4QUrUWEVBDxmt4zZc/9a+vUi1UkDy1s00utfOceUkMNyONY
jhp8NNJs9ct0Xaqoci/vrLy0B4WbZ1STco5Hc+Yn4nJrBhc8c5zYtv2TmcQUQrNt/JM+LTBbJw8z
K2hJLDFCoIt+jLHCDdUhuEqLJbK2wXJdgH2xIxqTiq7zp2kd2JojGv58RO5flFPPzdgIBwM0C8mM
/CVY+7ws21jFBACPiG1nEkeZi0VL9diPTMWgMUjA1gjfw4qwFvpRnJbHI5Dl18SPYep5WgGNpHKK
IGFRf8cKBAmvG7Mpsd8MRiSdNqeoR1khAkI/RDx3plyKtQuwb8dHDbVRW2CLA6dB4hRMebOn6geu
LwCftAopY9vGI+E0JW0vBwcO4yC1OGT10VdnC5ItPowYzhd6uUHCJb6743xCTewaBNldrU2L2zO4
nYfPE3nfBudYzvtWD/jnTAQ/d3c+cnzKHkJzPT0vShnaUVidNNM0wZis+zvkNvAnPH7fMiTWD6tJ
ojTya2rFrLA0CCXXn1e2MfJ3JEZLRub/yU9pwa+qKZYX0VkGZcnmbMxcn1D7w8xbcgcj/0S01jJd
F8z/tCW+6afpBraTTy2B/gIdRbrLjyicFCRXkChRmHYDBPAOe9dF+tsUTRoiAGQm3OyRFChloJTJ
l2f+LcylNvXFUgvvnSMt5GydRr6V2ommP3h9Z2uzAe4LMcRDwnbXV/9TzTZNlAcZiVesfLYITHn+
SsNn6fA6KJ5TWmfwFSY3rMijBrFXCdAL1P/QYRre6NgJyO5K26gO4ieTDLzhcC6exG3P/NR8y2J7
YS1UgTuvu4TEQ7XcDF9zPAg60dxIqaa3a408pk8Bs9MqtYiINUsSITfUgBRL49ZrKoom1fuR8ELV
mz/BtiBdPrpTOyy/iaU9H5BlMZqJXhDdXVTyaY9VGno4133MYSCK8ddajAwLCvhnhtqWiUYMLXKQ
2RUGfowfESz6seUKF20Qy/hYRzl8jXQ3uHdjlOEtMG39z14oq3roBb2XCM9vBT3p7m2hMpi72eog
g3Gdj/AO45u24v0EXJ74ZQtLM9KiXpaYocUYPxugdMn150qt1ZMhkw01H2HAVYpq8gPI/ONkyrTU
YncCXzxcEyrGHkKNY9bMC7MR7VB+TJ1akYWZUws1JHLRcZNYZ2ezrwRTlkqMDc2JT15iW4AW8obv
5Jq27LCXF8WLABOLvt8ZJrzPITX3Rri+SsWZ4NhsOxdRFC+Xd/WNrv4kg1HZ1kFRW35Uhlmq6jhe
dabsMC2P8Bc/oLbmInOTspRIQcAnmpMA4tc0d9CBJMtVmZ3omxvTWe/acK75yY474D7KMLo1dT4o
vQPiPZq/JY78PHs/z8qHUaeysGi0CXsLosuAa+OvMEcZFeigje8P9ozrELbuFI+24kvnXc6mwAeN
l947CR04fb2waGvgfcYRvvReEAfHU7KFu9lwbjVdNEtkoNx5EzEfI2dDxtrY/H2YLqOcSIHrb3W6
Z05inX0I3JG4yYyfAMZKH1qkpbTGImcGjUnBAwyEXO9DSVB7aVXphB5jAlVtnVl/hTTT3VMhFbh5
ZEYl3OOtWVmRN+/5c1d3ne8cyVX23AXZGIZKE+KlYVat8KTZslzVjHLN7JkVh88xv16uxquqCXP5
Fh54VzQnwmjUf1Yy+zqVwcfG15rpHO9/6R4kD5oXIMnyE3ZboCcB4ihEGoF5iucE2n+WK8sIdfZI
1MnrtOSEEv/9GwmF+9OeNKcWim3CGs8r7fc7BTJzeWrveAgOBnCwJmGCxv6a5e3JbYUK1oiR325M
+k74Kv6TK23h8ynfJpMI4LZYQXW3Ic1llLkHOkZ//bADNWufYM2///exoVj0d3FU1iyHPiolUWTB
hu/3he9h6tW/BuqNh49AFSufja927F6u526J3xhByeC69VR5z4Ee6i6efA3ScjappcJ8zDC5Z/Br
jweXR8q6avG9sRGp4asBSRnnsxqCu1zfQFPjqofHV31kSi97KZvlOLOxVRvvudxrqFvUAxT2so8L
1Y+Uwcn72MzDnCKHVDd0zEtU4olLhh47iNSLsKwfrTBjr+jsj/Z4i34/6JuE7SvOEaE00bHyeCnj
ilvcvr0kDrS2S/lFQ3XO2j9YWOnC6Zqs+UG8siFoyxaSVACTncnvdB8LsIfvqH35DsRst3VyV65V
Ki/HeA10xm9sEuu44meCTdH124x7+MUlw0dN7syLYGMtQ29kwkGmBuLmE/qiCiOxqWWVtb6bbs4Q
f0KzLBUsjOnVKeErQIMKIg/+HXE4I0vN7h+JuNIvRvZl0f9j1WAHtEQSHd+tp+q/vEX/106/rJVi
YgPtC2/4y1/v0OcwB8YdLZUkA1L0+A+SYdAQdXJpIpoYMRxT0C4sD45bn4+8XYSJeoiOwCy5MkgZ
x/UlCKDMQbQl5LiTJ8FoABLz1y2vfkeCPbiDWKDME6EHUnkZYUmNwbhrT7NVFtoupGtwz/GosqZf
2+5A0iShJrSTJaaqCyaR4/zWg9hT3yXmx3edbavhiH5fN4z1XL03Srnlx9Z1h+eCOmR8flBhqjXs
BJwRADET/YRfn9QCRu+/jqplxCz5ciOXgQvtpNwVMJBul63WTmBQEUx3X0uRy136uay8C9tFue2R
jd8a7hYemKvvgMdgK5m23qRztELspZfd8GP2FrI5qVSfdYoRFLxk+s9A1KTOX8NBdFLMWh4PrBFS
nR8RazSk2/96gK3Lntjto4CXxsDiK1d+LL2KtxilzvKWd8JOHvRhdpij3IkWtZR+UwdXiGCPQDZu
ZW3piyu6Se3jyXJCkqKgJPHoJp0uY/uXJYy6/KUkIj5Jl2cE8s9v5wFVmF3W5eEtoJ7NOMmmwuTv
gLi2/BoFIe4ay7GIxEBNeXDrzZzgSIAxaGh43dO2fb1kJEVMF93rvfMNuiwuN4SmM+KieMFOyYxC
0emLluHXPoXMyOYM7PQEp4BuyGemk0x1y2BWocnGgEi8Yhne3btqC9npkAHOzp8opbUdtMZIIa0x
SEdPiPW3QKSAxFqD4YzSWQ1mn01qFKvERQq6HqtNJiSVE1v+4XJewv4USs1EvwsUEcLbjMNU0gOc
ABj/ENgVM+1Wl+kOeuwxr6Y9ZJI7OZwFq/K17o0aUr2Yv0UfF66E5RtGw4AdmuX4oVwSG0Zpgf2Y
k1fu9VaI4sMmEY+vUAtDsR8Yz/0h4+d/fX9UCECMyPQBOobxtflSCOPmM+JdZxJzL1ECen61UVl6
koV2ItEogSKkfv73yFSUnIsBChjbrF3FJEMTL36v2VE4CBUjHKg2J4do0opP4CgQ0NOuvsUTfikr
d+znEMJtIm/hDPaMg3W4Rdt4s0YioVT3x4yf2fD4crf0u5aboc76skiH3G3dpBPgYG+Vv2gPf/I+
BnRXxGwm4+IYTcUYarZUU5N4xlHH3QOrhCFSKNlh7EnOiaTZQ628aU1Mz6ra/AQh+OqQKZo0kdL+
dFTAblSYvMjli9be200naQjpMEdiVOhIkoCgg62eHx9Edb31r6VhTGvN7XuW9w10kFOGiA/NGyTJ
UAPLpZfeTazY9ssjpXe4Ude+8udAn2WyuOCzJnBQCPDj3PWgaOamY7cxLqySeSXsJt9X9NUWyzwB
uIOLR9bs0Z60U5m9ysihGzJrfrFH5hWBQ+qelTcJngRG/djSZ0ZBK33ldUkiJuRx1mli0WolMYJ7
GE/70FUXEAPmrPtsT8r3uEap2GdFm5CKQ9jH8fs4AYGRV8B5wO7mjcSf5GCcayUiB8A7CU8nCHU8
rHSADf6ewWYurSNwuCacpM5FnN1xRf7rJixt/cYrkn4faDJkGA0prWZ0XZrwA/oLbuC+35DE0sCP
qLBwOQhv2vRrvW+6D/YN4GPyiolGwlTK0gbl9TyVwbtRwdywoem2KP3XxMBU4awhVe9F6wvQOEVi
pQaEF0nzsL46eBREsjKGowQkAtSjSDzcb8LqLOAh5AXP238PZ6G7lAizrHyD1BxL1Oa/N3oG33uN
S4r6dN/KjQ0/XO3hR9drAjM4bMbqNA0EfEizJuzA6t3VKIyAVO9hrBgO5z034e0OoiKBIQEVNZju
UYmR2G142HO0xcIrymhs1H2g02S3FeWklA9+aV8T2O6z49RKpODm3r+LjWfXfxQ0V7oVW3sDDdBp
vRN03Xd80eGyJ2WMNXyW3k7bWd1cf6vgIJgrA7LzH2h1hvlEnhF12nzdcO6aqq+rc71MpH/ne6Lg
pdIHl1wRFzM1rk7u/tXKfL/Xb6rGmwXYRjyIWNZK5XRhBtXEq+72MxnkJqadnEBsprfW5L4VTmkM
jiYCQ0M16zcb6g3YkkbDv59tAnBK0w5ZLvvbjMRnzAf4BdrIUfheKz0wjj829yabmloV+/fzg/eF
HDrHiSNTdMy9CAj3TVDPz3ReXVbVY6Tn1D8wL/BhbtqTtZCXX7bo6JYEEzVqa0GFiMhNqZp4c08u
IGPcTXnlBJcotPZrd852i2eyGztZAOBrDn+E1Apnox0wCRxh0DV3Nn4v6KtF0m86p7AnDsmaPWm2
wboP8ZcnD/1UZWJ/518boDlh0DOsPqwpvGFlyT8qkwKbsypv1uNvOVdPomNz5wWva5KS1SFJ7yog
T7B5d3zNq/FPBaruUCCmX339bTiXtQnUDOaxjQJGxWGdGCVbSmspYLtuZQSLM1KEUG08XRZWdmw5
v5bkVtRYA43x9Muk59vU5cE2rKrWhUrl6n790BoKu8ADLqwZDj8NYmV9pslbLceBfKw31ZYlYdT0
JHCJsmRObZt7DNXwZDA5dwfc7lAlCrb+B8ORPnrSxh0Iteb7kxufoU3341X5PXyHGT9Ozn7KHz8h
jvBGjZfiKi9g0RmDKpfOnnDlOeSwOyXgRRyULpk39ktHfq5JTjsJmy8ZBcWpu1++FoHtUhmcf41L
X2uPLhTGOX9bPxqiluKNjwMYfh236j+6tEer+i61uZ0z9zy6uaNwXVtRXuUK/nTeF64jS0R2Jgvu
gFz9Pf05h/a2HEarXafpvkAXlMSoHpKvJOOxWRdJSjpYp0JU8SJGS9YJhz+rsZHVARhB5whGWCOE
5O9rU2TyWCNiXPEFUkkNMebsMuEWnlhccN+vZwViw2SmUsV1SCErHUGyLzCx7beNvOxAlfvd71Mg
Hw/UXfagJjkz72r/gL3sYG9u4vi8NWWF3xrrbv4cW6QbtOBDcKLj7i2gRE7+I0DHuxlaUwalrB5v
x4TQk9i7o33BmV6ozCwVr+d29/SdMNtvgKJX+R7PeaBnH8mIKyEc1hc3KwJtXwUzHDv2zKmEpEpp
x5n6BxZUXDh6ZvhwZa7MGlZAnmUu+8BHtjdhbdyquBpPHhamqiZe9cfXcqwCOxAb+9+trg0QzFhM
XSDSYmUZ4g+lwodd+ONEuoRGFgWXYOVd05+coZtF0gzgNBINyQhcPc9UbIEtDr+7II92uwVuGjZw
M2FyYqRwKozsRyBmpFcQ9ah3u2qVjswfVaPtryZYeWdC0DjuvTchOeF4RsUnUOn2MrhUJ7IU7sdB
6UhXFZ0frUuBKvMY/ScptAB/NxGgjafHQXoLLCCjkbj5IyCfqsHE7DwZSio2VG3sBmgJrteLHktU
7g9UlIl3rRpyowm1Ec6x0hTZUjeLxWzUt25wU9GHgcSM6GkLiUF0tTiDqPn/G79JX6JO3orMG4ls
IAu2JgV9mT5GbjeEJTkRI586yZVEiyUPgLGHEXpkf2tO6W4E8dT5p39p5Vq+bJu24MyctxMQWowp
muy7qwBAQGk9cwY1sqjmOYVU8GsSKm+l+O3Li4OiStx1P9BoZzi141rdoJURFfxBdVGk0fHrREhI
yKczbY2Gulk4SliUPbVSNtAEyg6mMJiiGZ7rNT/oO7pBgFAFF057sU07apUNlIV12L0yiTBYHfoo
wNnBWPHBsPTj58j0lWyzOIaPWXrX/kzjgSe0wsCto6dxsTYz6EKwtQwSMGwWBS1OU1gpso9Zo2yz
gaHeFxsZ40AyvoJ1ncbcJ7MZfwJCNAc0/sXUDjnvOj1UQQWuzKKDQIG8m+hLLqnmCV47nu6lVH+H
AWWNbLYFe97CR5dM1bYhAy8RMDUWNVL6FywAHTmSC74ohF0vP9PtukAQZPSqQDYwvK4afd15ev0B
9GCBJlb0BgC3haVIABeUYXUgXmb14Fw3kUGfTJ9x53Alk23ocKNwKJpSb4C7C8CwYyNwDYNKhyFU
hD6t53vr3NCLwGSSi+ZWnaRv79mIn3Qt7ewQQVXEe3QZlNM604EYhMmCzz0bwUw3fA7q/fe+O2IM
NOhIbkf8QihY6+0IUDjhfl3sR7x1cFk4sqfP2II2X0Z8/36bvxgwj4Bf1gn0URxJvcDSVm0MDl9S
sXh93WiM4dU/ZarjWAhWbypqJOJZhNE1AR65oxw5cL2t/oQLmoAfSVKpiuujM8fsVYgqWEowHgAr
HD6RXAvXmiEga6RmbVABcTCJvE5rS3GWom84NBNVvD4ZrSZpr3maOGZHXI+BoQJ+gXVR5AWg5QLv
xqdV8TMP8Rd6OiJ4AwAMmKABpEAuxzeNzv5wit/MoadN0feyrk8E0dPyK/8eMkJSn8ZLNvmwpP2u
ObkVeAD938+MNHwMX2XjeVfntR4qcG8atgp8g0s4WthT+35GHEl3jKrV2MaNl9nL0Y6d4nqXp/9p
yFAQYYCkPXKZvnKMxMtpIYRaH6KyrRACPeGYkbDltTMRKuy3LSq8oo6y437g6Sr8bbUJTgAM6XVo
7x1wiaWaATb0VCUed07CaPZxK8qyEt19Iq/joqkbBmZ0a4QapaHxyTaDWLqQfNSvyMpo5JQaI/oY
BXXTCnWpzD1nrwiz6+p9XxP/3+XIDkkZRbyHLM6cRsKUmnKjDIzoeoH11Y4e6lwiifuprOKrAT16
qnZ6vffO9WDGXipvF1n8cZSCrfY6Qvfm4o9pSe21Ncx+X1uGN4TErcGgaXT0EuTGbxuNc7H1q0rT
rc2nFaHUWpehMyh3znigPnw+K93HV3peTG1PmvIYCqIM64HSkV5PhkiWDJ1C8zH7pDdpItRJBY7P
3HHQeIZip7PuDY9KZf46oX4LZVXqRpOuSff3NnpIUUSavqmzJ3D/4WPkdw8VbGwNr5HEClWZWIQV
YctLyojSORZixWgGIgESYPTyPLOF+RyAZIyt6kGt1DGQ8mvbQQJJEAKlwc8Nt61/rgrdrq3Pr1Rx
NCjXqrK6FgNpfwQgZ/Ey0DTEFnUOiPgYHg1yPISFwY6Iu9rUw21kO6dbsvmbUAF2hCxjhYzIEqjS
K6MQFLraTRb4LOCiI6jTYsJm5eTFCvbOu/JnAsYb3etBjewOrXNId6GM36mFpFNA/JFkIvdjwokI
Ff27Q8bmnLcxe9/VJ844AdwkJFnBxeUcWLTeqsIjtxHgua2IZRWOMubeuWTefFFMR7rGrWl1IRnl
2b5HOWpVNUHRhvss5GBMYUHui+/fuEYCrWzP36KGrN8RIRcJQz+sLGr+HspIZOv96u6DBTfZK+F3
/ijAEPQpQyz16+xlHnmMgsIXTaeXOnX9I1jLIW5v4yp57q94q8Rx6Ck/bBvnlg1BR6XVDZyE4qm1
2b6NyiP7SRVixJ0453ZnE8Jrq0C05ocL/LPfHa30678I18LT2oP18IWLOKThcPLoO3ziO1K9gEu0
bMwxrVP04OLl8/4fc8AP6KbwXrSIJSUK1VAJSvnbbT8IbWWDIRwp38jDnCLZ5Pzt527z+CY4xTUY
qITnotRAqTIfhydyfNrFEOMObmkvPCwQtwmsLd5uMpz6ltkcb0vWauLD4EL9Jp7fhz9fgcinsOxR
XJL9r1Uu8nPVFS4vJNyTW591Ffip8p/iarDE2NoKaf9e5sMOxssVuJPwPmitNLBmXyWfBv8INRSv
nVFH2dOhlHAYNSeRj4/a8gsJDouBYvKwgH4XHw+JHfp9iV+7f84e4XyPBMh2EoJNYL4unVVtGPvW
6ZqF1DkAakb/Cl1fymVngnm0aCNOiBCCk4K/e1qg7uNd8efhl9AV6SlMCAYveqxptbV4K5rNP9Hs
YVXOg+OUpMxXcS22ZDzzDJMCjCWhLkRdfI7agbbmmHVmXMexZ+jF88/FasXUZWo1jlDwaSKdnKMb
oQRqEUhzp61dDtexVZgfR1rTw1UT6+N2keZ9YS1NqIwmWO0dvp8msAo3p+ibnuhmu6KQChKNnaTk
PmVSZf6yzLqqqdclF0NB5h7r6E6gkUy1yZPT69Sx0gA32kEcyJVg0iwILxGzBmoQJV1UFAF3kF/f
ylI/Cu+tCcKKNgB+PPD7AABhz2NQw+u+So5eCC1+jeDfRyd564KlJgLTnGF/7bcvFpUAZZ5yGv58
ckFjsmy+mNKgo6g0jdig1iWrZMCXtFdM6nm5rigEszCZs5UnJwt1maYMSfozVTXDcbydFKX9uM7d
IveJWFMQchqviS4eMHYEfljiGEOqnJGNvAvMA2NgIP/H2HdMfjiQOkVeLIZV6+3SN5ZNL0fo0lW0
UqA5dIe4ZptKC0M+yyhbBV65K70rUn6joDtwbq/79bytr3XXIhS/+ZCk5ta3uqn4wJK9dmepHDM+
/QEzvzH0hinDK3ftaJtvfeSKUC/qvbuSQIw+YcBvsKYKT/55C7ZB9NRl5jiSTQnYYUI02Wf9+H1N
+uIYcY1MefkMdclp4apHiryrfajFRSs6D0hArThT6A5iEv8HDYOOAjlYPp9SBwviN4pozTAUeaH4
4WBgBBA/fQGR2QOGlm8WoA6LqBg1HkPSJry8ZG13ZhWOPLS9lH2AgZPJtRtOOOKZQ5rs8VX5Weur
aVyTxziRAYkbsM/V69l4dlQRYszXWkhD6eVXnLCj3A0B45J0ki7KOFtzhdQJtBE1ujTFJbGF/B4s
1G5aM5AX8oPHh96YRvMX2Wung9/KLRoiirXkwSZVKyuFP84j2jn8C7kQNPjzVKE3BxOOI+2rrzY0
44bJdUjxcGdbNFvEFWkGw76YOr1ZJcbuGzPz7YoUBJYLn69fO1cJxUSn1drPOKVJjgbG8B3uB2SG
zJuTR4VjtPWb0oEalxkDM6EwaXBRrZF/LBFbb32cfIVLvKEMdcHpNqBJAgcCoQ8Dyco0YW/rwYPc
1cHb5XBl1aUN0qpcAgWzsYUCdQ6M2erZDWDPaKXu4ZDTIxT/Pfv8RkxCsMgw6kH5aTSTcFmSNrQK
6DOuOA7PMoOA2PYSY4JJPBLPSesAFb5g5vzKOUTYMaeg4vb8GqykNpVrQORVfdxllMtRM6twmDNX
LOxCBTPecxReYq3WdaMoihPMoJIlSkVK0SFLNlmN+ghpjwxKJnPTh6WKIM6kAdhu60Xdy/e7qp55
+eAxuQVpXOLMhndLLnxLxyBie50akpaGuSDPDtLURNgCrIT+eLqEJT/r0LB5O81szuFnlgkQ7PcJ
Sm8SBVg5XOtnq9sIapqjKW/wO5zlH8Z8Fe1QTXgdhTWTG/YRFVzi0gL7h5UwDwydOGq9N+ym4c8i
Lf3h3rI82ZcOSx6ceWRH0xlji0V+mt9vFiDzEDEojU99ZITtVA5JKZZFex10rjfknuW5q+u1zOWU
nE7kphIUGOTxt+CeN2605sHnyWF1Cf1HoJoRCyPWg8lpzoX1jNKgL6zks3I6IrK49jAOlUHP4Qmm
SBF5OPv6lsoX3tfpgqivGn3ezUZBRFTVeRBhmmS2tz7GQtLAV0AwxUZo8m172BMzG5IAUVFW7HFg
u3rpxCa+OlGc8ZkrBHEfbd8TjK1LJZ1DS0sEcdKN/A8nhkZ8W57TpbtAvIo1ie7RdC2IZD8RuVMv
ea66nWuRef0Xv69pwBIDd3xM54HHUxzJWgsRvGsuRKhgZmMxDqPrGGjmdIeMJWXk4DS76bDtDGpo
1dsLhjatTrt0gkSqm2viTKh7Pq9EHrqxWb27pLMfTgZ159jKEyFPUI+seUgj8ZAxM6O9PSRZ/ueo
gNYmP6Uva9rr/kYb77Qo7W+OaGVd4r87xULuNVz37lM4xIJulafGso3uEt5WFHaZbesV9QCSm4OY
3WcHIQveoS/POItEHMPQyutD6QxnmCMN2Sydau5Zys7yitjKvH03e6DrOO5pa4vs/0iNgToIQ5LJ
4pqP29UrpNlHRkPEezAvZPuGGQAhfzHxtC8tGZy03ck70ppBApOH0szEP9VeIq6+g/4kt9LkWuoB
ffUlfOifzdn1ywU+rfAHv8BcGhVGLn1lvYCSSibx8NgMQAK7aPVAhpH5UR3vlCSmlFZM7KRJGdqR
4ULLolebOHXXDncOehETOpkZcvah/7O9xiTBrofhOMoNcaahdL5P+aH1uYkCP3IK62yXnNEEBXvq
xmuUW6D0u7qoG6xhkM3KruXti0fRXU51Biu4TWCJu9oQ/nrdpz+/Llg5pqHLNejWzVHjXZoSAb+s
x54NmjUY7n25I4ccp4zM3VpU3ftCS+zgfwiHeCqgpNR2vbhyrHlxQ3bSp/ZShAIK/yUq09C4u20U
mCgbhBITgraqIo0LbMim1xlyWdbRdaXfdke4RBdU1g+BJPvT15oN45B6kDeTbZ3mqV11VsJHh71e
eY6mbUWB+WqnqjQL82cZGWbrV3GA/givcAF/E/QWxID2rwgUdu62mYb51BveLrnG4ZtBRbd7ct01
m7vCzeTJN1NZX8tDzQCDkCXjL/o+E69UEa34iVMgL6uNjYPvae0DnzhSC/Ig3+7UXjiOSW7hJMnR
ZWhK+G/0R4PIQJwpPCgfxgHfbyUqWqnA0+Uy8dbHNMniAqYDCEjRv4CIpoCwsGUfelpZp6ySWij+
+mRR2wWx3b2HHDHRhJYB/x60yq2DdhxBvEi1NpzZv9tT7VCzLF4ZXCJWLJ/V0iYH7YMb4nZ4cSfM
Q73g+PUQula3b20+cEKqYRPiU2SKRC2rar+BquGJF0x924cAzvL3bKCSXZ+cW6pa+6ldvBEFZTx3
rS8ldvKV0wdqnq3IGC/PjqeHUHp57o6tKIPfeN8e5IbQBNyx5Db6t3MXxQEbjZRiJVqElcI9eFoL
gHyJ+IWiApaXywXAvMvzu+zaiRv7DggRgQHsHsq1MPVg428zOo8ZcM+vl1zE1MWNWM8yqG7zTSCe
apINmTJmIgkT9zMHXjUyEKkpd95RzBCWCOo7UNbzyiiWzehkuEAQtsJFALFfPU02VVvjT9QRu/3X
lCSVw2h1Zyq4XT+7Cu5KUKFEvJVQ9xT6mb3nc9sbNJyKtObzZu711zdkTlzcOjkxi4K3p+D56x2e
oNPf/Od3NwWkFVT5MMSZV/+Zsq/iAyy5IJu6EvNhyrVauyaGcovYaVdPIQHYu9sd9lymEgG57MAV
g+ajyQmwPkBBcYELV/I2XiZUkaiBT/Nrzv1J5fWFjcGhhjk2wRVsVUPwG3+c29kug3RT/f5d5OLD
LhwViEzxClGPVb6rx8vA5XLW5h840aomqCq/27+C7flM35PSoOEBqiBIzBXzzjgrRq4mVh2m9gQr
/NuB6Bduwxr4ASOgKSfi0All5BxO2HOps1YTzzDzURbP3iSmqWQ6WBCegW1Clj8q4DhCimDSlSMg
wibfFWgwrNnAbJss8uo9eAwPL1IdRyLARP4tsDdAG+V8XwRYsY7jDhqQIx0k3paBTIZBUlYfH42o
w5axSZFwGqLcOmAUPnQWbiF2aYr6Fm7kdvUFixPYjEn1c9fUpXXBa4FH6Y2q7l0to1MVAY6kF4sj
dp24ZhuZsGQY0PSJ41EFy8rzH6qbyM3lQASjNZBB7zwN6cLQtO5w3p6Ki7cJDRfXSgMnL7B2jpQA
Z2f0FNkTu625Ej0/bquTS33dikQJphJM16H9YHH2N3jAdhUtnG1sgDUslgtwWvk5ZJEnjjzbkxxS
n1L5vbW256MKILPiPs27V1KFrLfyg3LLk+hD59IhApHooM2MPdZGHeSAUqS6/7FMGXRBCGRNQ6MC
emr9Hih03VSVOfHGGGS6SujnNHP4dU0gpU094Hx9s3N6cDM3Ua4fk2qddMTf9oEFS/EGe3DX8xA6
VUSDHHr9kV55g/cw3d01N5TMaCBbgj00sdTtbCg4urBl8VZhhFNcK3IYZMjrWCotcOabgARVIXqe
T+n34ntU40qiSZbyRWxBDLGrMdx6UpO2D7EesM7qw5cuwWKItB3RSyICiClkTiv16k3FUb3yVwOK
+L/161lPoQVQOopYYj1zNjELj3XfWLqCqkcsR1DCeFeJr4FiRVFPyDSn6oN0zxyBIrbvvjp6mlt1
TPGx5Ht7omCteHOInYmpvB02P6rVsSQsLZ12aqPKU/YBdSa/5s1jYqV7EoeUTPolU4QtzHOSkTOi
uwxxWpzcoa30DXXDaZQKo4GvJ8V0l3s4CQScjuYP+MNvnyOF+BCv4Kj+OX5NSMEFlKEKOZC9jT9b
3DgmMLPh8oiGDOkNpYGLLaQIhayqRZFeA4Nvuhn9aw1fTYbgFujBKWYMrRSWxiJnRfPYNllp9qxJ
U72YKyLbmZ5BEys7O+nrD8Qy7pyfXPgOqBbeNvmZw8oa6BgkG291vWouMePLz2gwxQnRX60ielmg
F6oEPeqQFmFnZzFI8bpuLZGUvT45dayWCNv+rM8D1kB90AkerHNeADV259U1mF+b+idlQvmnUmjN
jimqrU6Ei1jxNLSQJPtog50mwUDGUyom2/U1Y/mFyhoDHshmRcsi0hSTAaWKnJ43AKsGxWV3PSwi
b0347CiDdfbTtDTI1SpovWaLIzPGtaxfSIvKFW3PLKAtAr3SLcl9FmBPUqGIXNsJf/ZjcWvPQIXp
2MoWN41qBCQ6jfHmhBXIbeCkgAbSmhF7MsuKiIo43gWxw+SIJN9EpgUG/I3vlAMfT1SDuxE5CENr
tJWfyqaYM4Qel+2qGtMq+xIty7JYU+6NGWgWVJ7t7nCnaof5shJckV6jiHS2VeGQdqTl4hjkz1Ao
3I+DEFd2NFJxgC+mhZwc3Bz0Fpb7eqfXwqNo+DSMfE8fV0tMvQmLomOzgvMJ96nMa27KryobPlh6
qzOjiA8uxpGDQhDHRE2RtJ5tRI2TwKJVKM3V3N5jhMcW6Q8wZdhkMaH7ZeOFYeiB2bgiwHgFHXUz
PT5P+0fQBGWiYJufvORtvuzHj7PoPg2geKFjX3a6dCX3Lks4YftQ5preNDFDCuKsBS1RFX9xbEau
nZ3otqBMAm7VC2Bk1T1gxv0czVaC32Uaz5JLPh2+vuscpN5MQzYxbg94d9xEs8JfGTBP4Rvne5PS
xBImMCD0z44fX22flQf7ihLid4IyWNvy2SD5hrPuFkPBFgvlYiEbLTixuKiaVbwRw1HqqzQzn8O6
fIs4ESL3rXKiNdiaJErpKWfw7PiRVMpf4BCTpYAofuvcgDGrQXpaz36lZO/h9YOjueJJb35k8L7x
Cl0NzA/5goIGHhokf3HAVpVr2gyiVFgIfrQE7J+nEGTwhnn82yGDG9dkqpW2DhHlE0ovsOxkmH/N
UgUJ6BjlN/qVhiqOBkLQFO8PtMID8TINTAU3lgXMGlCl/Y8M7V5HzGA/zFm5QvqP8+FGripEK2zQ
OHcaeHWMjJHJCZUFcdeoTnTZEBjd1IoVSCCyWCssqZXcehXiwLXttx+FMaDiunNc4wPbPuLR4IOb
MIFNISjqA82cQasI+x78lgx59DvlT5tVQ3gzLNZ4AO9O8M3JJAsBFuLZLgC96FjbusdSSx/fzCva
hUdj3lsDlPm/kwuxaNvydeBNAD84nEHE9zpYBXiMUpQ5VuwZMF0okxQZnB0s9tID7DXZw4bsGa+o
D8Dj12YcqqOOYabqsXn7JkcBAvnQK8Cp//qnINAV9jfB/tTeUqgvn8zLSRBxR+DauqmAWo4PUzAA
DbUyDkEj4ezQzICwZQEePTTXbTsiunDFVlBefaGPsFa6qGBt0/hwQJU04iHcTaVSYQJ3njQb999K
dZPMdT39SEfeZ0JXfPn7wxwHKNCPRbDQtku0CIHVW2cwvX7hGXxoaf0vDDKj2DSxTnv5C9Upzxz2
A7Ia9SmFE9LIlt9Q4EOQ+06/cF6g6NN5jROnSLCj1OoFVfrEyRHBGYKY3bhM5ERlsggn5Y54solo
RCr2zZNvyJSrmR4RKgji/CFBRmwrQko/WtP9836dYpWN6gN5TAPhmWACdL6jEOwDIkFscISMdtYa
ltzmOOaXO8LjVGJI+xVLX4u/4fBXmLhm45tFJdVst6c70Y0bDQo3jImtWlZoKbb4AD0v1baI35gN
htcTKMqEpLcE/K+kcZ8mkePYMGGukVMJ3hNYAX54GO/6ZNRiGNwf879M2PhiVC5RFp94DFl3bU7P
s5oGSPp/qZFhkD22ooicvhXzUN3GTDgYrhzsQB0wLoJ1NtMyQlvWUG0qn9pjl5LOglVZpUMS5Mje
emsrRTffRiNYehSfD8MtX8ab0BKqgo4FQ+le6ZpK4AO4muOwo19iF3YsQQcaMz/eceVE7WKydrnA
M8MQxdtUpENq7w9jZY/vRcqU6ft11eEcy2a3NfWmeqtfopygRl3UvLX53ybI0OjvMEeeKj/6SleE
UiIJ81jGByeeg02YKHRVXCohrRz5bgfHSB9og4ndsZtkYoTUWgMNaOIQ33iNrR/FKlZTazlIpGqF
5nylqoxiWZS9XJUK1mU69nru9PCE7kCTKEZkiRPwD0nJoJt8muc9lkxtyr5KxLKPhgNFBule1omb
iaselvjWBoOGU5pqM7CxaAcQas6RAzdJQwTt1Dz6lwA60v/qrQaWDdWwwjw6Lrz1xVrgZ4IKeM5d
uor1cs8iKUf9dgFymO0yPXdF5WbvAyMNN3PgMdP4qP1NgyJuz0bzzVL7PdqYsYdyfd+IQWbB5IWO
cGjZAdanm9/A0Q2MzuBETBynZHeIk3ZJnSkWTSDhT/OQAh4bcisNZ7B4qdUAQMa1x/RsnfbTlNlK
KX3ZEDUEzF8dgF4SjL9p9WzFYTW66yItAOcqoRHwxd9MFBGnCGkpFl2ybz/uHL31Q/vBJjWx0Un2
HoM5nOw1zT6srGGSuTPp9U3pV2WRV7cKTiNdX5YqQXP2vcKdOEjOzFNMMCHoLVYol8oh48nMLv/j
CwwMpmlzuS4htNVtU+S1KBtZNqfQYW49bQQfU4mgOYPBmTFEHTXCE6XZvgJjTy25ZsL1cwobvKji
d9az5+V1a/fehv+FgZ0arqyPQOJAgDURbR65uKiUj762mAZ1fsiuVDV1UAdfYs4JiucAuPfrWbSD
0EuSBFckTHJD1KMgkGwIE5k6KH8rDaws6TQLfDn5pAmXbXdyhQQU+P0aywymA2LTV03MQO+RFxLy
feI92DwW1hSkul3NH6I+iGGDxUjMTYbzMzk+RNFunBPC+IrzAvRWAfgtoq6o7BKgjTvJaazvnY6u
1IHeeFZhnW+PXZpQW9r2e6v7shF2UTaNTEmSiP8OJ+n4/OJyxRKCMRIQUJPhCQkVC6BVQA+tRQma
WQqWUl6XYTERUi6J5ACbaDWURn7RS2nyIyJGErI+ZnYmZvxQvscHPSU5YhqAesAmNTVHD8nOCPyk
sMpYSOTsLIS2Yq5TUcGyT6Q+TRbBvrsDv2WOEdUMBCCAlLoGcZdb5ywv4zPWeiV6X0APLAf05rZ5
8NmvlVp3nmz+ypamP5AuCCvDJD3dYPJ2uRlkUa7YczSrQBRAXtpXrqX+Qm65MEo1B8NvTUkRGS7b
jIwSUP7BEFr/y6uQHB5iSfUajmXhCjNcM4KZXh9YWWgOVThyxmCJnJA39sm2Qh/RZG3FNht6KjPp
QroVYOtvHDySSIEV8oEOKhGW3+lAXiFDexlfSK2xKPsWNocUeRq/MXqHEEFBCoVfMUwyJFOU+KLA
DVYDn84SyD7jJARoYAtlCTCW7nTLbl8K0sC0ekCHyczBk1yDKhRQfj/ZYYKEWIe3dCBbmeHNZp5o
+bAJ9Yvix6MkeUgieJyMGZAxmjPXqu1b7RhL3b3yV3A8wdnVOzBGc2BIfVFt8uqiC816C1aQshJJ
c6laReL/oVznNOIcyBDwCQjkxumeYrXYZXt0dOc1ibC4ghKdmN6rFbkUmNKMT+cBkK32dyXH9AiT
z7U0vVyjgtmBpekG/y8kJXSFY3SUhx+8xeUyl8l+ior8e0e7KOqCUuTCbgK6YVgPcJB5c96rzpX0
L18pXWz8PJIFRhsOMnEitzTv9yOuIv7aoU9SVM+CEpjqHYvn54sZXmxtbG2w8PY4l3YtNP98xu1H
V8F79eBBXD3CL/ebhdbZsfsNgzbMQRsaCSs3P7V8XUP+cWyb1ywcROxuAD9C3H5fo+9G1A9ymzC/
1AORHCbSl4LyLpKmd4q1XZxsEOjzEVWG24uQXq/E+1SZOkwHHsgzCDc6puk4V6Qs7vBq7ToFxwIV
ibePn93veGm7m/wag2TaiIr/l5g0LMgvrW8EBszLuX0FKZNaUVIDzxEA1fIXYjc6twkN+xwqe9PO
96glYIfMsCsRQvDoMTt1bmZpFeSWnZCJ9atjfswAGY2eVOoTqwEzgyuNt15dP1mSaRIjG3rDHlPS
k7vI77VtYjq2CzxDERSN6TN4qm39jVPhaY9McvKMKSovSMhzTnL/oLhEj0aZj8GdZeJEb3F6SMpG
H3U3b9BrgNrSS0CiynwyQQGAldCKEZMjlhHe0sPTq8y7u9ODAaRETa31ffIKafXJzYYiGIdop6ZK
ZhCJu24ZJr84V9lTVrw4WLO3LHvmDWb/QWmNrB8n9BjTTz8M9p4b6QVl9GcUeen+kdD7I1ZL3ao8
n1ffS6P7EWqdOrMssWUFQsmFSHx6MlO96wzh4W1gYIuQtsuFZKI2K/eK7pI2LW+PUxGl7ANrEO28
DdJGhFJ7d69ULW3VJh3Ia5VMMGBvW9+anQqfRnpSe9amPXfqY53FrY+Rv4UvM6iEoq8sb8HkmqAU
MWooYGZ6zzrLnULqcDaVqi0yoUEyAXcig8Uj9GC3hxaw8wpr7bpZpS+X7X8e8y4fkHWmJrVE0Pw3
SwrOIoHhN2VC5/LUJ2OYRZ5BMTOnKKgcKRDvcamgJkMcJOerNGOpK5ZQZojJo5O8kQZ4gN9LsoPE
cwxoUYbXdMNKWBDb64w5VYI+kEw8+D84JWueK74QT9COJapYucqKBkZn69FPqiH+4iAGye+MNSU+
UBlH0dyGu7Jm5QTwTPv+UK1XaEtgtmskgt7NLg1Gu6PUE8IFY3/RqAxcuY0jb/IRyzsVuzUsIKgf
Btk5kT3RYVQ0ze8bJQ5kMDFqnzLo9AVJd/RC83auGZkSp2DO00+qCbrGtvuehBAwBNuhzt+z1Umf
ZIcu5yi/1nFNyAdPMNxnIn75+F5SoszBDI370fjS3ByUQbpQtRe6dQgNwkIa93aNt2wRtEJTu9Eh
dhAayR+rkY6tNoQNaj19ySiJ4f+XymiwbZgTES73p7qWW8AH8UTQLi9Kvu3eFk2BbLok0XqsFP5J
wcfcpIbYDKgU88wHO3u0kQvs1vdZDpkmrwommelUPvCRYNIWX1lEBryYwejA8KJ14twxMjM5Oy80
y4+YFcAmG6yWgqSYVerZnbXJtA0iuVZ0sUzDJP5gGEkHoeQ+ZHFKI/eIhedDybxs/MQw/I1X7ATm
YfY+5VU5J15/M/dK6usgY2rjFtYcn82w4KInPR1UfJMOcHf2u9rIbd3J326pB2/K41gV27783LR4
l26y8o0OcZ8ATPSxv6dd2s66IGrVj7jz9SIYrWdiV4Bjcn82usBeunbu/7bwxH7vN1RpUz/w7TXI
cSX0wu11XvuOi+VougTp/3hOjRkmTGDLfMMu70Z6xj0QOvkbIUfZwWy0d5H/aqqihQZ24MXA4hxr
YMcM37iL9ONLIJ7aL/RUUXkfAEgOX+ldSvnLVEC4T2iw43NT9A9RMyQx6HU/UzgNq69i+YTa/h7f
9dOsCxE2TMLVoQdMGoL303iAN5aZpEC4OXLqhQSXv5r1aYhRlUCM3I21HatQLiVA/mx9TmHcgyj0
46NRnP62MYpu/nvPTFsFwE4VumC4Ymkr/oH/TsDzyCuaWxhgW1GeSnhT8KRJN24lbAN7W+r/RrtO
YtfSk36A/AXBnytpT/tmdJOroQGbqd+ZKEQquOgTDeODN0N+m9Y1MsQryTSMbyuyMnLKnAjbUNAI
kO+YHKHvXW9fb03ekWzB3r1crxpHgLqRKdPwGfHfAKSm5CdxpBmgRNCJ7ytodMi/b1BwuEPaLut2
tTe9ZmSs8aerXJr4YLBNAWrNMLPOb23bEd35KgDjwvx4FHeE76I8dkNuHK3FlvRSQ+WdtetfHZEx
v35LOBO3NIj5lLXMH5RmHkrjU/2251rOM9uY+r/z8gTergFJd+ohsJf5rz5lqZPmcDMjStpTxyBK
S1LJQt60LahW4vcKkIPVDx1+UJRjytVv8m4lhEApz12hIHJq4WIBSyjBw6Cp9hMb86zQ7v3s7BXr
zixjTGT8O2utDlIoEySMfekA6VqI7SktKuP34wrJAWgQCYhHw+HKHVMJTb/nJOyVQ0UguVdssanM
7NfzZE5mHkyQYVpWOoM5pRuUJ3YkQ1rUM0RFZiKVZM1y+wT7lEtPJH61pM5FCMxfdudirSv+zQ06
cHtCLCggejjSafQ9Jhg9vEKJrppK0EAcVctGw0Ko0c/Js8YzifrbhQkb6HUliJQdCP4EM1Vk5spX
8cdINIln4vzCCHdZ1HaN4qFNE5Ez3eiYwkTdHIenriSLNGllscQdfC6ytuJmnus7OwcdKq95NZel
4BH0H+nJBIRrXDGn+ZjqBYnGb049DNTOsGOJABl6i2TWeqshoeoFvnD1kWAu3oxnIds1xW2h6V4K
+gqcwZs6+JIV1ay1fq60G9aS/1LcUqfP1np9fvSKBM60qVOjqOpaJSE3V4kSBVYxcaQ5ku8IgX0/
c2meQCkkq/l6cKBk8LbFBFFPb7daSnoz+ToFsBvDWWEvXwqDEGYew6h/3tPlLtISZFDB5HjWvrRc
hKHViGMNXCXK+FhqAjf8LuF1cJvZRQYgGFQxcNwSHVCqPRw7/jXp7/9xcTSqw01oXwIRZBfEefF/
qOvJJN1/94yAu2fEJ6QIHarrjojxvvURh/WFxxCulb+9sDi9beed2oeunwMGYW+KCfWwf9aQPKyP
laY5lKCAQohuPfGs44b88oEHBCZrJXFv8AQvLftzaCTnSJcFCKb4/o6ZurH5/0kOpwCDljN370EC
dP0vMAtBijX6Au1ecE4vxyGo81dPVCz1Hxr4uTxtHIUfqdSe0HIP6LbD7UPsFXnnHi6LmbIoCx+T
HeqPL0GAllEgq9Gw3uPQ6dAuGlGl8Dw0ZeRX80TIm07Uij3hb02IhAIhBwiSMErawAFITtCsVzH6
H8/3JpWCbVmFi8MHtc8p4o2kCqtQLGokyDTMlKUyQBVuaqs1XgEwXV4RpgB7oOIvdEHpp1W8/MB0
oFdhmoskZQy3JYWnhEY+CQUXrIv3+NRU2rJVQISFhO6kEMRkzByzg123SL3gqBonzwqh76zfa/GE
vTn3oZNqWW5QX2g5IDis0Cse/yNb1cwyTtT+bUobCiZqBwC5eOXlFKH91zx/+rMHSEsXzgiEecen
DJOxwjXGPqyuWB46eW3WKfZFtBZdad+iMbO2b+v4G8JW+4c9UpCZvK7HMVF7EoJT6BrGAHYWvmoQ
LNFo7EsqKFeKqPEBMElxRfzMxTS0RwAKcxx9k3BKrZP3/kUWvHBZxEABQdkHfYdKATdaXf4PNVKL
ZVWI9rkzaULgOQakZ7RKN+J9cpCXZryXqKvPJ1yGjXsP+RI5KLOoW3hmyonM0m/mNjR0qV5JWA6B
bqcjqJxszCO4A4kushLl7jTr15NfvpgRr8KHIO36cMSDvrs8Qj9VF6OanD1huIcaDLiz4+xSw0Mx
GrtwFolTv+Ftr+nPWDb6DbISZq1htdG/cYJQZIikGf5MQH+PmnKa23uQTEGOUKbpgSoG5NchxVEW
/SMkg7t3FUZs6pDGLgDiZThnBbZkfoPYvzpcrsHuGxqu+/5q8QrH51g4FMPvpWVcgDrfcfWkqzmz
CqunvNI4v+lWiakRptVaus7P3tCi8WWqWrSciGO2Uy3FNyf5NxA0hebftKOGm9WRVvN0t8BPO1Qk
81VzO6rlnTSmqefXlaWYs+BM3EBESpj3g+44uHGr9Wvmo+UMEowExqcfyeU+ywHG6pNDEHrTJwzj
JoX3jQoakNst37eUW+VsxLXwvClVl+LluKb6R4JuW9TEUQ2axEXyVPEr4ps7VLo1QQf+9zPinQuU
J7icrHU46waJqrGRF8jorSTxuv3lgD4hhKpbiWAWnJrF8xDTCn/AAWgzEQhkIVTjVAzUSjvv7LfT
NxzG7Gm+MFCelE+FJXXe/McF8Un1GhlENaSywTrw5SuU7Kx9x14txngrX+spglIATr4pvCGABAR1
nOCxSv72DfXAXRf35GkzQfV/LUgt9Y/dWbPFRhEUaImoaEee0TqDFLlBR3PHMWF+s0qFNn3Yv5HM
tUMh55chlD5E5u373n95M7c6oNAmGPAt1jgAXKei2s5/eUOFOcfBS6v+0pACcFLehZ3/oeD1ss7W
mQsHUR70+BMTtoxspvG1ZeU1JGG9c9skuctZqhb+BdJD7AqG52jAaTy4gSKb2gQQkXvZ5mWrr9vn
IYVt3XOEWv/zbuGtx4ePFT9TSWwBz13/jhW5BJmlfJeVJWwJHW5ExczvaXnmsiqfp0agNW2tVJVS
nDbMoMK/2vFweL3cjm9tuuGhqcfd8wBHIghqQRCJ3vtdqjAzAWqggxI1jFzLtr76fDQkfo9b+5Ax
ssqjE8rxzmt47sUJN8yh8xU2sxjB+dkvMJdCcNXO0gRE2DQMnXu6hqBBxq2AmK5PVvH4HYEe7CwZ
07LL8otWav+CmkD6++h0PLn5oRXyJ3bvMT+16Bav2ktQ4h/+ovIur460wvCFL0h+F0rYrpH+xmuH
WrFX2rN7Vhw2JTlbm7dgetNEaGmWuuv/+nIRFhXid29Bb68hYFrR+bmKsgG8m/ExgCbvzQU4s3tV
utzljNpi9z7man2KhX/3u4WmCuzXUujvLlYLEtHi+AG8gsQZPSI2b+oxQlXxGrRF5y6RcnhmdGRU
KiRrEYV8x9Ipy4nvcUz3DTJOcKtLxgd62y5GDcwqiRlFERjpe9DfZdiyb2xUUbhEoj8w1jJqFSTA
oqLncLxGQCO0SbXjsgNxAuZb8TJ7jXWRnLh8/5iy5onj8rE+6aj0Jk6/36lEeO5veEbPjeRCdytz
Usk3F+2WaOfzb6pCSLbNH7vx+Qk9qaXPWr61kYEYrDSuow5m6PUWlbGVaX07nOr6GcwBV/50S/77
SE2U+9YOjhxE08shUvLrErCUGyoygxsAyVFJrWJiixy5dzQkWEes0wwXqUQzzi7xuNHaDC4vXzaa
ODjoufmYzA62COF/Rts5/wi0hVcqNPaLWQOXb2flqU5vWL5GjSQ98Uxf4D6Ln/0QKJWgx6CmyEAZ
IL0UXay1VqORP++TZRwwPp4gwOVNPd7BRvbBeYjSCFb2JLldqtBDp6xw0WEYi74UxbNz4dNWL4Hm
9RQrkEApleX//fG7y2QnsUjmfDfo7JUTrxsQOveQprl3vmUhDPRN7gYTayBxiCN9RANquRTUMg/g
MZmjaohSzEdAQ3HQGuHw7NkOA4efcasctEGCryp1g3m+Ke09np6TogKUV6HSIr28+SRVx+tjBPBM
kvWR+A4EjxJU3/3CmLGFeCXmRqk/n9BRSlZ99N7f2BN7jxnuDJilL3HoaZhcrcxq56bH9jHH7nOn
MJ0eGL74/m9A85T9Dz6HZUXm7E5j+RAx8MX/GHNSHn43N+Xp0Zp8E3MvnZHqKGeiQNMgiEBasj9J
pCTcoISeB9j6lg4brdp0ivd8VmLfJJdhMyglVfA6Xa3vFIweu9QXl4uNEfbt93imxzipWFYXRvYq
Vk0UW8+u21JE4+tvw3QAysJqAL6mnwXdv7abLKAI4ELt+yJKxmLRefthBB/jQ59JUQfo1Unku6xH
/WuQ7gMfUn58EaZCbPj9nJHXeYA73CzQlyddBlWnyoDHroZcLe7ALTgRxqiBh7wU6xXoABILSBsb
EyuTBfDFGwzfwltXV9NNeKtbDngEEtOIYmWBaqXiw/sVXXU6puD8L4S4t3zo00M5yf/HNcEG3ohz
Klr+cvhphRRlI/JJh/6XqX84Fjink+Eyjd12ugnu09BE8SAJck1ZAq47oAaGVUQ34QK1RvlBSmfy
Nyl6GzOERlTUbY6JIRpZD2yKdbcSjTR2tIy4jHPRsVzzEKtSlgbWnwXIro4FIVrnjJqIGxyxpzpp
BE4L5yow3sd7vAIJ7DjOa2ns+3g+wy54bHhO/rnF/0ehm1CwsR4D57QOvnAbNtmV090Zroq7+NZW
n+KczczqmuNL6qf+b1HgSDruRaAYNsPp1pZa7psBlSIbF+u3oglb993I8pn+c/SsGwSeRCmv1cRF
4z+cyG4DkS/WNASvqbP+b7F4Iqx7BNTV1/S93w/Rf3HopkAdFOSsKvxFVctLzCm8/QxuuVXjhD9j
DBLX8NnrL0aEBDk3DeJiaWZYrXZizPCTTY+17A805Jeyc4A9n+28ERz8w5JG7Opvl+u5xxqavJyg
J7pVF5e8H04IWQQwppoGMOsMs09ivgZfn2Edv//q0vLtHE9f2W33UUdAJRGXuLGhlI1jPXeslTtV
XpGGq/rM5+30T7Sa4WMaSSfmO38SdxyqxaIeQdjq9KvnlPiMh8ruXNF67pMc9VhR7tXsuqxj6bpN
6B7T+IHWQfVNREb6KfU+z5VpfqfBgl7LanSr3LM3MGRev8Vn+2gg1Pvq+osz9PjMWQvuhnMuEwAQ
xSJgAU9mC05Z5BUqY/CvXpQ/hcBgVA7K5WSbwv3POF6cXYUX9veNY+cDpb47qWXq48e6jhznrlcM
Y/2ec6VOXlOm3ZhkiFmuwXJnriSqiq9Vm+qEkOktyzHvcOFSR7w5fA57KuYGObnkr4Sn/XJtkMt9
zY8TnU10ApBTUdqIXeAKH43XR/QQqOoTGBHOTbBFij6FXeoeO9Ko0IEAO2Kl6dHmbmAaR0emVDCP
E5Bh681i2zzQnZ2kPb2n8SxRpxK58fuDXYfGADpojmJlr9sFdHc1SndldgtlKZunT8xrjgZbzhbk
sEsxVJXKVugYEhlQS99g6cU+rn8MVT3Qq2qa4I5gpYNsQ15AqDNOedJTL5aNFR1+Ke6+HaNfc8aE
sqt7rxwNvJ2dEh/OGhgCPkWe2P+0B4vXr/kqmvun/zg1Ql7Ja37W38m4mF7HOMrX5IDv53/XnLDI
/5Athe2BJdgXIMikrrnaJwT4XSOfBNVMPpks0POIU9L0irJVWL9lqRg+//uZMPPQkD2FGwY/0PA4
htzY1mK2h6XUbhc2r/9dMSEicbRKwqvK3kM0iuQdg5gIOUfwbD+Jr+Qr+JI0CYJQTBOroGItAzwZ
ek7SoPMR7oHeZiicymm9Xuz+kfbcYOqGTCcipLqo9k0E0cU2CrEKp00tXdJy75InxaLMDQ5RyQKO
R5sCjpjzVBoB9eoyzFsYArcQSw+4d06eKdNAhjuUcIdVlAHmCw7LRxLJGUZyEnJvS6GllHXCVC/d
34bssc4oE3jmt7yTk/Zia7b2cbzg1hm3VatJ/OGlsPlHTGqCGmbB6/ukVOAomF0Z+Plxwjde7xwr
fJZs4wg11Va0cugStpSvgqWw69FOJCCNJsLRGCEopZLw9xJBNQ3AgWf651S0W+JVLDB/4tRXazzi
sUJSAxzMWEKDxV8v6l3HMXvX59fVJ7l/g36YcVeHAEY8vqtIHRTDzJfqe4LXY5DZrmKruLq7/LSM
Yu3TvUxQ9navIw7sNFBssJ9x2+z+YjR4sDQD5YViQrLUQVOazRPIMHpCn6IPWKBglVmRiUQNdoa7
z+iBQb17ne6kwKOWF4KMF8t6E0ZrTP01BSMSrnry6I/IFeRuIBWBQ4XwvDJAl6k5YdqlTUQ5buv4
HhWFo+8Pu2QXqMO/mh310NAwZVvGDv4EJ/t7DSoy3XuY5VUa3PlsrzD9szMM43K5/TX2e7vSgm9d
9dDW3ZcOPBDtpqHnlQU4iBoYBon45AVl4EpGeEe9G42bK08OjzyN4zRIjKO4sanHmawNEC3wKSbh
yH8uCsqHc0kI4YhSxDQEV+1z3LysDqkCsDQaG2bFXHMpl/l63pTxslx2PIpbTBb7Td9Gr5A1thXW
bfJfoDk+2Kqgx0cEhtZNOH1AWYW838f/4y+abI1mOFPP9MgQR+NMmkN5xCpgYbGERcuXBAVIonLx
HWck1jVfSGrnbowtSr4gOGTcJW3cK56jXGEhPF9ZxOypDgpkyK5E5s+3Bbfdr+tNhhhgc+h4C4bY
v/T+uUHIwAzP+DfvE8A9W7Gf21VXO776RPGdHFwtDIcsVwznX5e6cQYIXV9f1niTal03v3PSECz/
i4zla5GSqDGrso04YVvWfOr8MzA0K/YIjr34PtmkOs0vS7su3aM0+lSbClOFNjsh+xKJ9JPdHXBt
yRE3c9Iwesj5A+qT+4gfj+ASLUKMBbYKC1S9Vtsa36gi8+yFc+IcsR+P0smCdDCaDQuBcRMMelaR
B+kSpynxWnZLnvHVDVnItFt1bPE2siSQgnuyQYH+6xwght0IjEjEkeykIOP2nZgXWO5oTE+xT/20
n9AMR0lcLWyCXAWMQd7KrQIKjxUNvSa/Kwm7LRsURrmkXe7WWZPMveBazIkvg0JYh58Y5OyDUbiA
7IYmadW+agenpWz+bhrlM6EZbwXfj7lxiomNUpoG61HVTLSm0DfIkgxOCS4hs7GLjnXQVtMILTmE
QZkxoJpK2sBZeJdEuW0SIAh06fgTI5BtvG+ZTuxwkfUHkd+vvD+jcsGjaWmQFZ84IupAtGArFpw6
42/q0fR4yRwLXQrzZ2EPN5aUdAnOOO5PObPWTvsEI/IzFJ6uH/fqbAQNiv+IopyC71niuf5KIlwG
iw+vc5DfSKGiTktl0WVogvFiZU2Yw55PzOgoJnRNkTRfFF8rSIAogFp2ogkETuOb69TbNj0WjPEN
UZHXEoPqgm9aLnE0BwXwd8pYK6lnHvGxqlEY3DSLw9DjIwvkBPq0KyVO8mjxY5z741N+o1tRWcNZ
JiRvB7t++AXvNEag/OV+Xs3bG/ObBe1irRuNJWFuhwiXx9nLZqxwhc0suTC4yiHfYfp7jStW92ea
gSBTxLjrj3N/t+ltz9nG1kvljigMwxFJQunTB0T9E2BdZneJUo66XYRXbl8I1/sQNWRH4ouDevau
kjlf39AftGZra+f2EiIAqDs/NSfMApbw6UhtysomDqeOZnV+VkpSELSXIE+IhXwbGwlLvuvH01Wn
7LF2dirO4MVASHrynpy71S6reiJaz1f6oZbo608D/DD/XUDVMLjItfX3zYAAyqTiG4/vhu2fd/3F
akbkz0tb1Y0U9jcTCgew6BP45c9SENVeU04Wk4EhWHCdsgOjQJwDKaYVnviTBe9CeEbW94GPNdos
dsfjMK+/h1JnUdIadsJsjlHb+G89UyMistcKT56dgK6rEzhhunFJCgm3+ystdEAfVt6Zf9MxA+Mf
gcq09kNBrXphgF+l8+V9ogawpOMuuqJ4E0/1v7i463rGTEOrB7a6Mys2KEEwzUMoOh8bsaFjygmA
rPZbSGTTAxNr0vh+SxXQcoEEXFMfpn/vwiTMxVMqqvOKTT+KqS9a1o5i1OzP7tGkwfleswRtXtsu
Kr8clKa/FIY+0CiZAW3ZH80r+yAR8wAl9f/lS4ckPRUicMS37lbHGLEH50sBY+bWvlWLw60FZOuM
ybxvzSdtG/CejH7TsEb0AHR39la2TEAuHGqIgpmRa+/Y417iJgv2C+gVvof2OgA1tg94sb0yhDzC
UWPUxD/ULLbDq+Gv1tmWMbgAGQggD7nULOtxGMebtTWncNUlh0Zp7XN+ETlRdTMbx0941oJU0u+w
1rmu+GNwdcRDC1wUdOKGld25EMKYJ33DMad5YFHFY6sK19Eeq1G7uXX02bji7MILDTRG2jhoKMja
+HjAtl51d+y9gG5hfqlB6H7XMTQJjRN5wnr2jZyrExDUXAFpMq9FgX7gPbigmMcEAchzosMe69dZ
JNy05Xwp+t2xNQeSQ60TqMfzcZBs7pMJoRX4j/kA+nB6Bd6dVSaVJxcLfvrQT6ASsRFYtp39lVEf
9sR6mMDBmoPJcsZD3preM1BsdEwPTHJBWrq5SSy92AhYxD6C2BiLbSrkl8stmlY9yD1Xr/tgiAEG
dCsOGB4z1hufCZt4WHSvCd72fFOHxpyqQfRE0Ni26XTDn9duQJjAMnNHCk3CMwNawfHY4srn9U0c
XSwpNDEWBc7zqRxyuBRs41Q6nTka9MadtAxOkuYRt2YtuyPDKhlXeuR8tptICaFGzVUMrs9nw+hp
uSiKc3PEz5bXw/H0xR9SWiV5QTLkXHmz38fAtOPa/uyiuopbBVEPgVv/WGhynTOcQmMH6zp6Xoz5
bwCTzN13jSk3FWCpWbQcsMpDXferVwDmpO2IzG2GBRdHeY3o1vhNkUNVfQgS5KrGR4wINRUXzFTO
c2qCPFbMI30KavdavN9YpTdtMMPLeOD/zgCU8e9kl4idLk8YWFT3lmhb+JXfTyswGniyCxi3QTJL
VKzXhAAh4Zvnl/FA+mA6lZ3OUdRWEUMOXYRpjqaR3hWa13zZHO6Z7eIs1dihOaWpvJYamX6YyI5P
H0sMsjrnPAaysZ3q02Oos59DLlMcbj+OdqzuQl5E2jlUj77OV/sJgRl+RotQKIK4n4n2c7GKSE0+
8xl/GiqREgvJukf2Pnzdh8VuZk88HOwDOfCPc/nokZsBXCvlzLd8Vnt0bo6S6MEGoAMLKYN4Lz/4
FMmkRrpD7IJnLCtCx+33l2ZBMg4nnHojHwQWzsIfgY2LAEfhgMbTeE92gt9ekQUxP/agsOUc8CGQ
/Mr+8wsKkKFHK2J3YBKy0zdLmCsuAx4L0bc3RvZ59XiHUIJrsq394yQunPrLcjFnIJoG8t8hyRyE
/hgyc3z6zeI/vf1MzdeBf7o7LVvLyY/YoQz8qrFYqNrOULPzh5JNgEQjYyMWyFHoS58v+4oLCvwI
rW5UQc4DCNO/2ZdEo+FCFUzFjvJNb+rWb2erQXpO/qOQoEnYq4rmE3310GP/tqWy7rEfNn+A9H3D
4ULRrbX0BbOpAZlmSaZBJgp2q+8ZLoQZa2GSeGzgexEN0pXXF61Vm4XQSqaZANvq2T4IrP3+JjgP
D8ON6a9TMpZgYKUun52UChGafrja+dXMtaQLofzkP52FEpKwG/FGkz3zMuubnlRKPwxFn2gAUYwa
uysRH8Dx/ewtZHjpMZIWRuBmTUxST5Gj8yka4HnqI69sH/Rr6MKPDWC/2CbkT+ZiUPZN39fNCFQ4
V2dZNypsD3e3TabY3IKc8te1myM7kRK4Zfy+YaFXqjN8A2lkC8+GcL94DwOIF6y61o7FhSvMYAUw
Cam2hV0wWzMQyCVfxKnrXV/For6FCxOOfzYjRzIMRfe51A4fiit58QLBOUCq8lOura1irV3iEM5Y
xmERG2aVlC2WeHwjkQeZsEVFhSTzxKlXAHg9G1OkH0v5VXALwDGf6H2tWgIGFz1s8RwI2SQ7Olov
iWOgOrHZO8omPAEqI7hLHqcZjA4FyYCB8ryQa6jeiVVrVJGAhRGCCvZUmkmG07sfaDlPoQ2gvkQa
FqGCg93wuLc+vYvKNTsSiGIoJ4sYxH2Up/OLwtFr4M0qDTdZl9kN6FYdofGnX/Z6acX9OoQf+Mnj
OMacgl0kWR0gi43TbjcZ1a4lYKpPlXJyzEMSA8IVR5i2Weokv/3J0i+5OswLbsfli3mZsw3+m5hG
8SwrUzxWL3QJ4HYj1AYHpqQdPriIYcrmIcuwMlkCXjAsGRpAL1D6MYeBEDMfThUvzKl8aYaK6PMT
gsTB5oGgx1+I4n4fUYAqdJrkFuko6R2sXR6gSs3XE7IgygsImRf1cROPR4j6KlLEJIcsK8WvOQr2
B55H/wax1htZPBygwF683ktpYZ1kx5TGQMm6Xqx9Tu3xFLirPgq3Wtbe4UkR/pS3jhR2BrAEi/qT
izeJU7Wh+UJm/QOHcQaWpJJJoNATsFJqX8iDKWMHMzuGa92jCMJiI812V8OSZvGKAwOGNEkaFlrm
gImJHqSs4QGjqpfN/4V0yEult61Ap2P30lsbOjxUIVIUPgEJHphMnwoJf0agaMgfghEz5BGhNNqS
pyRq+XabrxYnuT1uTMjyrtyhAZ5ICRsYDkxtZmCy1OZG/7mO9NK/d1G64pmJxqWLzfjFns76SNJV
ashcUK3dYMUbx7SZctSy/kixrIAzOlRi++Bg9M6oF2XLglbY2qgdk1O9FZxx5X7SRMHmwS0rhb/t
vzeqhK1a59/PYv1uMJoIYAHzt5OZnv5xF1U00C3sfxk5Cz7cNYTXurLQwfYjnCJCIJUXwM8x2US0
JpJkt/LNJhMqGSqzFHrGrkFpmiPwB7YB9LA+xtfCK/qdhmWmBCebRfe9mIvxX5iHWec8iC4QxdRg
2/HOfte3ls/rM+eyikAZ9sE5lSF5kTaSZbxrD+2CDr7+Lfs4/M7hE133WlcN/NgYgdFVyCA7R4ji
o/hj2yrNyIlM/P8o8g7VD3ZjhPrUBmtLJSNQoICuEaKF9LNYhxQgz1Ft1TMcHJPF3ITp97Q5R9VW
CORXULs4jJAyKUnHun+0rNuNIos/PwGuC1nNZ2r/XZCeO1K/k/qJsWTDNAfI53FsiYNlTndQs02s
oBrjdCRevAs2KqPSI46+QXd0m1HegHlSJWrs7A+tQG+j8tEXBJeDR46uknKNk+IgU3Eb0i3stzTl
T6nVi/3NeLR30HUFkpkJ82DVRaT9F/wI4bLwp3Ydzun/+6+ipwB2fNKq5Y6cGjCNJVoK9gHmVjzF
UDE2XM37WrhnXer1Lp11+B8f0sFNOIklXAx9TJUAScmW3NfgobA9pNcMenfRhCddp1T36yxvsMia
nhr8duW99abtl8TuHQ15yjHcQe19O6DHazHlSXMidrqxTJxqWvqEt9wZGL4FXESgiODDwvBr4yxi
UEt/RQwJwIPfHMN/uqMrnGMswegvAtNvdQaqUFzwSl4dm67GXYtbxuM7jRQgUkm2jdDYWgy0vXdI
Kbh2OJ+EbpPC6h25n7ZiO3GNs4adg4t+KQAH0sc69y8K0x9p1jo8BiL7/2qDYGN83+kiQGjHoh4T
vFfndeOQIs/64Sl/+/kPMIHXWkNwHeeURzVtM561B9hmxmXiUzkpL6zw4/ChSJ4wb5NVCPGKtZhI
KyH6yh8I+qRn3TaYtZMUcevWxX/rp7Q2a9+V/6a1O3yrsLWNXtkz8k3xfLkzrfgyccTA88g6wTza
mSiV7irh3AnSg2Nzh+wYgSQ5GbyuabLk/ushwDCIyzR4+hDW8VPEy2fknnxcTpzs0NN35r2EuZrP
5c8Gw4skicqcP3AysGXInjNqyJ+oDRUQ1klqcALmqRUipI3bfI8+X1/qlAPGRHJVEo1zf2lBwBqE
a27I/hP19ZNQbPRXiYkUI7jyA7GoI/3ZHOwVHhC5RrXnjFd2o66HPcppKAMWD0WHll8Ryu01yG0F
Q91kuxf+0Rveu30AG8I75bTOB/nnjTqZjcqvGAsnZsaLOOFJiHWN8ZHmweMmjGTc7Vghypjd9yED
Z9SYvdnPnIps686Bc3oKwBF18s2zeawjWk5a6EbUx4YFNMd5Cu4OSY00J4yj4z6ZPepR81jBD0oS
fXHcYmBQJMIX+CjFFayIQ5q90J/OkXeDsuPo8hTuyj0MUVbVDaWr9nO7CROzW9eQFvh4sJAbDHn0
EMQs1UM1xBEi/dCm8nfGBvYCvW8pUODqkz0l1Ne1TaXWNH8EOJyqalVoU27kaZJYEEB5jlvzuIiY
QlyH3HJtrwYyYlkNN4wmhKK4RXyZmjnZJAAxNU/bWUsRUd1mfoV9BFou/I38BL96HHWVSYMTu52v
W092IZHNt1lqoQ24d/M+kOdLiP7voxghLn/xSr/4Q9UAHAy4hc3V+qHTgfgwjk+9/JLy+seQADko
JHjV9wYnNUQ8e5N/+2p2twDwwwPrBKBGsfqAjcWYMXfrwMq4s5NPYi9meplfmodKkZG56MChuH+N
VHaIoZrGQsWk/AhEb4bVcHUMbg8NX027FuWP5vnvIk9siqRS1BNAzEboHNCyibDfQfb/diIlKzBI
aa4Fl8BxFidvVtstRChblmd4KijIcDrSA4ZOZ+BQ1xYV1bcfUFxA5CO5OzQDL97pnmdUeRpXvFkD
d1H8CiHFwDbp/2UICK/Jd1XFsrsZkeAxv7lwmM43yV9dAlDO2yTLOj8D+IIdOd3v0BPfsPVNE/B0
6Lhx0NTiw7XggMNDXH1VYzm7vZo1x4FdslDyqtM1fVncrXfiGG3cf58oe39xUTISRBTSlXoCMIik
cQk9lFA2ofCSTEqRoRRqeSFTF7CXEsCAwGsY02Mzo35BsvAnFzWd3T97cUJahldK0LYjXm4yJJ+I
MP0v1074ycRtauQr+zx/gvBBxwp/vsj3BU45aOL3B0dO+4jkVWR0qS2pSjlOCGh5HvG7xG4ib0TX
Eh/DTBDMcFc0g5hwW64QcGsxp46U0OmCBXrdEmz0Qeq8GnbmoIIOoCoHj6JojRIS5ODwfWhUDfKm
jbP0Fqo9EJygA1izKMhbfsvaWH10d2OZ3WIGRAMaUSXVp3j9I4dhq3eDaHpXeQ9bR0mNffm5E33p
UZasd02Q2IGO+sdTxAnuDYjUY9iqdwJfx0HluCELSokEStSatonAMAWTUOpMpHq7xxpY7xzZOlB8
eY09ogBqAmk9QqjbatJGAcT+d7mlqlJ9+abn4/njNGW8GM75eAI5sHyM5bKqXhKktco5V+6kkGFz
8V9xSBmuoDp4Q+uxwu8djnpgxZinxebxO5Lq9DXOMjakJAvVEp6aQtnsr9wyZ7iLom/mydABNW+q
HtQWvIX2/GDsXto5LXMM+LHIPG761eq+a+bnA0y+Jt5/4uey6A5Fug7eMmH2ejip857npRD0SJEg
w+/Mf8pLMAcxlV8mS2HmMyN8ijgLqQSqx+bLR2v38MqLiVSmhm+XA93q0fzGvdNNWL0HfqtGlH2F
x1GJx7cSL7/13Rtl6Eti0e6J/2KWIbwFyvQ7urH9Vlb6kcFEwuTip9luSIH/SUkN+XTfo7MPUhB7
8m3YA1B0x0u7RHYL/xbCz3qRfbJMH3W0Tl1meIJb5/WkrwnbnI6ideI/cbNci+raIwGBb3unjkiL
rkin1S9dE8CAMo5hoDje6MtIlzAfD4IcfhQP7DCkPDuaWu0OIL9C0OMvJtx5I49bwAP6HhSPxuVt
Ht/Ht2Jmr2gM/20oPuCYNZqmJhN/oFg+atIO+CojHUGg40LVeSVX9sLdI9fcCq/gGDWFM3bMfSHC
Xh/yen+8fShQzDhcVKpEBdQpFbpAExO7/sBrv9N1pZvm/anEJ1XQF3ERmPIhKOTGEBjgJEMLD8SI
4fHMmlJ1m13vvRdoyYvkYBH4eDV8As4u6mQA0aMcrweqY1ams7UM8+v0BFV0FVjViIe6y6VC62he
Q63syZCK4nIX0zBfY/2cNUQnJADeAWJzKNS4ppXt6le9M/koCEA1D5QV6IJ7l1Q2/79pho+7dFC9
CczxGM+gCu2vcBLTVAio0LVIQwbBCB2NYtvuPZ4mlSfZhKjGBKyrqFn40vz89O9riNXUGokRnkyJ
qBgb4NO9Uq1IT5KwkeBjCtQNESDNDz8ylfL0Y8prXQ7y3ePG/dV0pWq0b2TQksonGbfiG8H9tpDP
nsQb/nbfyo6mNSASD6Z6rg5rayzN991c/49pXS1KtXK6KLeJovosCtaE3zXD/OH8a7PB1uBGnTjU
obSZgJ1zaWnD3WFWOn6jwcKIqfiZ7aLLKxsF0skThIXtfQFbwOC9SVPCRgg5ASrR44wzftg2ltOm
P9bf4WGG5dYs9wrPkFvMOxpNFp3PjsuaKVsVYW/QEHf2t/gCcaMisYIsmd1qeNf8C4mvuJl1JXje
pvGNeUCCgMknQIguOM3BmoaPuGW4/ChSbkLTVceiddwS/yc5x/Usg5tj1UdM0+amzPDLuQN/KSGL
X9v1jJOFODbLxhd10apF2Nj+N2MqxkCiAAy4L13Go1/MJhBsr2bFawEDgn6/H1GM0Zm5CUP2qf76
Resuhcqk7QbgYXxJcn09U/EHVo06S4LGp0ALIFVaApHDg6a15q2BuRynSbY/j+KsQFntot35qkeB
yMMutPrHJakz6+BACEWF6fxp6rdaMptfROlfFhUF/mYNNe7tsz1MUcShfBoQfmaSlz317MaucFom
qPsZh0UvQ+J12UnaJwV+E0haf6FZVVjcCDJvV6dzhxqeYBNiju9ndwlH9DVB49/XyqYis7rEYyql
slWVepw6NeBCyss/zty2yhZmVJ8A9j8PPbtuWtTIgK424E2/pOI2JI0qlDPFGotBBB4e4vnyUVsL
y0QbWERzGnHkSqg4DnYkRdFJ3nqsBqNRh8tgvqFhG5fJ4zpRo3B6W+fe5S6UJ31jCSICiujS1sSL
lFCqmMiTKo+nqHImVex6cjqlfaBch0eb6zVL2piSSdzs09vNYEh6euZ8QQK9pnGRHx1ntNzIe2S7
JOUFKDMmFGFOOwgHnkSqVDLx2OOE78F4IRz8bQILqQwWViIom1zlQJ/VotFHfZhTz1Cjl94zXdeM
IYSghekh7IFUYM6ykRiJbJcgmO2pxmW8yvyolJaUgjP+J/aL7QaZSf+7mH+rea/blxCtTLlXq6Fg
IHIO8oYSb6jyVBg3QCLMieBXvO+99nDj2bfl5IwcNkJTmnzsDuo0uNUhfwAyBg0Vk1x5c4UPES+z
I28N/QcNfcvLM20uJwiIM2ElNONJZRWRPHWJ2NDQRt4Cb3RBFyJZsPFUDvNMEr6T87RiqJMgn1XE
C0NhFw1hcKtVJn5sR8+oculIJedftqx1yRFQvc+xSWdNdpKeuPIjavb/nskA+SufjzWEYBNLXw9l
4rcFOtMrrvDaxHqYpDzzkRgKpiMZtHel3XHsDMP6/G6QZIZ9MAldamjAtDdwpRnAq3Rq0ROcgXwc
RPYFZ5CGa4HR22GSyWhLmzhiD6AViiVoGbO/5LyR8AYHT9CDrcwcWG0bg6+4NsxNeDv3pCpe/C4r
+n1I53J59yehJ+jute/0Y1KReyOZvlYDmuKlNVHX1l0mAVeUoQyA0xvOAZVKMN6audX6BC6W2mHn
jQhGVSENWz0cvEYnSIGsz0gPXl9qc6bdyoz2kLtrJc5FFmxN3Ky480okwPrSMBDRMQ1I7XnpTWfM
UHeCFX8A4/SbDo48+74RMr3x3CDauMz+M3prWY6SOoNwuixMdFcPzAkydlmUy3s5ITdI4COeVVyN
1HfQa188qOlWEnAgHcyLXoznfkUxnpvOdN+SkgOlRk1wfKxZum/WVUX4qaJ8YiohU8/qKDSkvHCD
tbJPdNpPXW1mz4fU+VV6vZMqg4kOj139neaplVNKsqesllFW2y1t5QIY5gyTAvTEr622ldoIA3zQ
9BNRnD023IEf2U+N0pW9WMxYcILeN5IN1/As9epglsxkW3BfZEcZG+DTVKT9Pzi8y+zhpr1PUycM
BHrnQLixfkL16o+vNElCoB58xht7WQiRXzf2m5/QRWSRJuXHLEw78WiligXxd+uMrTwy6Ohd+ZIF
CkSqL8+U2fzSmzOAiqHZYEJSLTgtoNbPOuBA4jzXElWtzqRcRDsrnN3GufIWsqUOV+5oWPK7IdZ+
phjHQeaBczWHMV97kJxbioik61VwL4qyrMShADNYNkXfdME6M5oHawdEV2S+U8B+Feru1yJ/UtNT
ksWPOepn0MzmMXGzrAzwenHrHJFnK1HGjMYLkqm5VVQPC+B7Jf8sKkPQbRg28eY79mCqTExMKjDH
itYVm3QoqzYEf2qKO/O6vtvR3ohLKdfwk3gr4VsMlhiSKrcsykIrXIYWgvvdMIC59IwKZtSNMVvY
30iU6YIGxEYMrvP7YkoVLGnZctTz1JrSSYcqaqXZU3BRLsjGvRJcZPCgx0pBsp1ZperAXPffanzq
tpL8HQIriSaPbNIj2sp+0Z6bdFh9kW+b2MU/iFcj91qZhTcphVqpxdGuURCsaJrCLSuyqZ6I6hEB
aP+c/SDNhxZlqpV7XlN73G1os28ltOl+10Q3GTEfQk9Hrq1ozulFfw6az7pNpfO8iEhjbQnoqCXa
Ni/OoLhX4+vPWt1kqPp3ekGL5yS/GrBrfIYW0sqekDTgHYzKxbCP/fmL99GGMtt82TYC22JkLe7K
KYKAijcj9FjRXlFQ//amWKknWE5CIT5vZ1K6+RNYnIniFK4Mub7VjmzEQiCRL10JQL0saZ4o7XEx
TYYBHZ7zLU8rIK5ULAeqlGxwqTp1X+j1OAJ28eA9O6ac086ow09aumOxc/cErmheK23a3x6FrPRZ
HF2hCrUScYlEqN/toblZLAcY92xw2OzrYRINqeHrBGk54yRuHagEzGhnVAJoLd3OwXbfndK/2+yG
y8DaBuLUHBIgRVnS1E8bo64lcIxk1xjMnSTl2onU2WYUomZao/UDQdmu5+5iWrC5eFXr04CTX1u9
hbtbdjSWBu+VR/ThThZWPvCpQpgVV+i2kmOrV60T58hlgPKfABFX5EI9pKGhkZV7hcqav2Z2yxo/
y6hKdkDl3XRzobhxM6ienJ8uiGMgtYqutXLb+8SzZEqwac+QORIE/cCEMuIet1TN3Y2ETSwh0hGh
54sZUqQLOPFHpBfGPKkuV/QHJTqEt55QYJyzFbG/xHx0xgcCiXTcj4SL/T18TS7Ccirwt1XoDW5N
/T6FrYCo7CSogzesA5PjPPhBD/wEflNtDWmeH8oGjOlA6Ha3Ak7s2BXFGCNpVeZP2vVCuSHS7mPl
m3Lz5qhHEsSFwv3cTYBAkrl3D2lOoTCUcuLNH2VsUjYT1ryGK2RusHzPPmH6AC4oiYRHwBQqQszT
iuQ/t0HflC/4i9CGZd5w1rWYkgHxfbt3DmxFvQXhUomtmp9NwxhjkAJX+QwVQJjDoW2qpIUy0FPT
5jQWlrpcZbGqPUYHCmHC/8587gKL5ZpDW05LHHUelP0IBnAw50lBlzQ7huDnjRoKhOonri11a8sz
w29bVRWvcgQ0W1qGe5aIkKvWthNMqUKtwQA44GtCe/uvHH+VSY1R0ga2iLrxeseMzA805aQasgFc
mayiZv9q3J+384jhtzA82GjG7018z4gQ196YNozvwK6CGXSwLQ7fZwwESQ43YMAiV4n7FHQBcaAF
sgRugv+G0ozj8bkETYMoRcXI5W2OHpdk08s/47KNMi1Oz65/qxAMdEjL7RMErwB781NPG5WTjH9R
DgpZ2TYPo92F2nRteTNNPmoT4eesMgAwjkVgRTflw/xqrXlb3vc2hyV057+cSVcjp1HkghZkGbzO
8tBddsWVaObdq6mGTeSazmCE32waSU0gdl1/9JiCyMWn7zoc5ayYKZdLdZFi69Yf6Zbu4Zizx54y
9CDy8mO5YyHYK0ZSncD1UKkJv/DacRYbFcv5uFCJCaQDOrPAMLNitOxPJFI3lp1FOKfzLbx3boKP
z2teEMhJuBKynsm2EK/VQ+VL3LODpi4MYF1TIIig368QvJKJwXEe7fG0NGDGsTwIwjUL45eJQzc0
khcQ/XhZxs0JNcMINklGEb7W07pi5EccTPNpWMeIhuH6fTdZXaUUBfnTffklUcTDbLCxC461fUJC
7Chw34EuG7Z9ZHrs1oKQ3ma84zY+nXvNPMovkpS2v9xLsIHGHr7BY/zyHLMZpIOCL4XFFpnuxDra
XOGQwPme0UN5hgJVZ3lS/H7RdfMLOY6/2+rkCYa6i7+nmm/8+bKkJPqdhN1mIhqXJVCyakeHqQN3
Wb3nCsAo+nDM9Cenm9YFbUa4s+zt8D7DrZbYe3JlNasrXKyVC3QQOGs3AjgFkiVRh0zYgVimn7us
v4F1+KcL48mQyjBPmVXQDH+9xHbJwDU36Lmd/dw0jKftHzrUcto4mtj9HBnyoKWf3Jbwc6iDZvhy
zMNjeszvr/XS1ceZkf6H+MBiUmgkr8Wes0XA2EB9ye9vc9uGb0hSLA+tPkRaaIBusY48HiT6FdpP
6w5QDu6gz+FE32/HXFKjy/bVhcMp7pstfQPDTH1zr2RV4t6lMcb3VI7qsQvEYk9v/itlbho8fzs/
Vx+xl4nVujjmc5BRXleFHmsmtQSMGU6uAno1XyhqV3fNsCNNniopofMgo2kd69p9Y06TUSzQc2Yp
JW4ypQWQcXwrmh2Dngli3V8LaExr6hD0qdYr+4PCN7ieD4XhGoSfstGJLLQ0Hz6WxmsdjQ42lkWK
RXYGMNPWqwZ48eH07DDz+Zl8d5hU2kmVyhmXasVrrL5JVaD3ZBdlBjIc7N6xuNIcJln2gKc2W1+V
G4yJnSo+Dpjhrn0Q+5i58g1Ov6/DWVMRGCRLNJZ/SFC2vefBoEOqSYT2fIRW2STnzpfQL9mV/wz4
tg41ilkTfSis076qHXsz5xD+hBX1jYVw/UzlBvrD3mRxC4GMji6l1kN+z3dsNQZpJYkHSYVoe76Y
XurOZkRZKh46OYe8D4t0uZHis3JThEOsblBKdL2DNf9SvWaN8IRm0M3x7SJFt4xUlnzFlD4lRbSD
LHOmMrihwneghU/FQKamxhQUaW15L83j1JZjJ4wVrOtfrBEVZ9wf9UnLW+WPXGnXXvRLHPQS34+e
8wvDzwQmC9gGZ1Q2ZDmNbjI4DYKzC8WM5df+274YXsveXhvCwSmulLAku++9D4a13EV2ImBKqCjp
vauNU2cWZrTNTKIQZdD3UfsYLUmn+C9aTiiA4iQ0F5dbIoxXkfZ31WreWiFqBbWbVGE89LV3jnaZ
Ty7jgsNaKPy2SXTkSE2mxJMANHFIg0mp9AkUw0ch2ljmyl2EXsuuelxSMlNR7iiCTRMIxcgVqtgt
kmFOB/a8uytl5rrwhN8PiM55Po1kNLEpEZgmbuRLOfTb0oSTRR8wtTqoZGKXq2KUpwaaeS63gB1x
xxsRyTQxCKQH/3NOgkppRpjZ5pSiJZK3HGW+ylwUpc8MyqoJ3tJn2mrhRcp9qDQwKqdyJlG8/AlJ
vio4iRuWQCwqFA/CyxraH4aUp+i+0PVQMajqI0kS0D1ue3ttr2bwTiWqgk8LWDXYveW+Fo68wj5J
Dc+1N4WC5tfJZ92LFQCOR9Txf0XnkQfMriXxyQn38tTFFz8EWiQBNEZMY9EmsHV3EK9PuXqlIFyN
cck8jmuphWKlHqOv46581rRARiB3WNqyiSS6m1Ezvk91Olo3fK/iZMudSpt8rzaKpQeUzEDAxDii
ogmGrfq3QfT1SLQuvBksD6jT7r3gYjEv/5EnXp9m380UEyobOVw1AjI2xBQS74rjyikMsuulOBzU
Jn7SEmxzHxXm89Jmz98nuKvI2tUzZn0LizIwFAF/nGGYClHOl3RBtB1X+zlD0/S+qNXcwQCaT3+F
AJ5dZMvhSGb3dgQrZqqDfARZDpwZkWjwj+PdqOI7QgC+4Q9iF1rAiL4a2ron1TBxgLGA1vZyrvAi
wN9v9QZVJEpQOnlfeK/xyjF+NXxRiBv760HGMVx9xvCSOSZ5YrR+NdIDJOT4Zov2rQk+rC772rnQ
va1yj5rqvFyMHpeWUEEfETnhB2v/c8sjc+jvv4EGqV94rOX7tG/I2kFou2cit8q16hWmCYWOz/1m
K3guzo0LRlpDbjlUDzRULEqtoiNPDts0fP9g8TkgCV8lffuVDaMERaFXNevUVGjLuEJOAs03N3vZ
fxa/GqbRLewvdKjfKOT6ZbHEwNUp4rd8qGHTQ/0TUbuo1QQ5DwzRINvInOAR+ddgyl09xLyP/Fgl
YaRCTIyia3Wmaaeg8jGRcCtnWZfd15q0885GArud3XjUBGp6IY6eyHxAm+I47Zmb3+BJ9lMXNnDw
0cQrt1juw9/u2Pv0VnlikeJ9n//zCM9iPOCK5K9i71yJHE72gTLV9/KQ6ric4aXdLd9meuax5d0g
dS1wyfGnkLO1rHQObLlo0EmPF0RJWdbAq4SDG2zT4Lfd2iRhz8mH50GRbuY9YNruIopEwD+wGqJ5
Ix/dax/kwRE/MC6TNusREWAEIjPYlEyoasdSr6FeIxCew1Rz3BYLV2UR+5wxU9UBadBw7t6tGvOG
BLa6yIF7YPH7DYz865wL5BAxEljLdxuj/P18XvnAx3Qo/NWI7ColudSLCi+0bKZTj1ykzJGQDIf3
HRmHwcPXVwTKmE0ZTxdCfCXdG7Q8hCwMh6mY73zUbVuKYrflcxfq/EpWTMliL22m5Mu9wBCfdeG1
/5Y8rscqNgMZMXdfyiD66MZ98DyvH3shTXkZt/oYLxrbyBO1umEdo0ZYkvHkL/OQWSmyUTh3zu2g
naWIBIEpaiUe+rZZu3I4MswZRUtaI/pGReDPl5MfBWMuwKMrqw8gUkb99YjHQH3SNuj1HteBLinQ
0NJgRDOvxacV3kQNk9VKjaEkBRLzuyIzCg033491NUfmVK1IotCB+9fYSyzssbZwQpDZYxU9OjA4
u1x90TR/cC7smlGPGz56aNeZnAdA15QwoSSCjFs5osXyFeSE98xJUPRlDqor3Z3lBjyc8LEYzYkj
aWTDXqJUaLWCHf7ByuUsNjNiOV9AC6G9qInPz87kBiLLVjScpQrTmYoutrEskyX/6CcEGOU2E27Z
g0IePaKxVLO9wxsEqHDRXqGx+Ao5L3h0ZZP+d3fC0Wf3OYigtUbUHPb0Ewhm4Pm7d1tXxn5D3Ss8
MT/yYU0/pe7L1x468Jz9akSm3bXyGfzV4vk6tXvPdkw0VPFJeT5sLMRZ+175dBx/HlmJv4VqaP8v
zjLkO+ZRrqfAkg9vo/+Nu+30C/OZgedhNQP4narcU20UItZ4y7VBJic1Xy1RPwEEYBPa2Ph1b15t
/4x8KgloZN1Tz8kvwCFd5u4Gv09/fek2qZYKUkz6/fAHQ2xJ2zmDNigVdo9gUJ1aKzES13ieHgf4
fnOYYJOWtVTuZEUrZVPmQ+bD8KUFDAqyzYEzHNkO4Xn1BDeQPLHs5PHsWs8PWK/U+tde+gWBTZKh
+q3mk73USYgdqZyu+xovbIn5kovP80PUKXXL3GjfrgSMz+Yc3Eldb7ZwoFCEXz7U5ZbV5a5l/tXd
UcTdLF9qcxasU+Ilg+oYLHwJDKRlNSMX1jr1i9l8IUINsXGDAGGRTGmuAqJ9pCS6tzu+0Djd6Uh9
67mSibyuyMiEvzc+wlBNRXZlUMtEB1ZioOKCj0wepbVRebK7ORUl49+vMF0ejfSvprMW7dLJPC/C
7vz5b8AvV9N6VA53Ba3ORzmEij9J3Rlzhl7zycEPIFG6wB4mubFLA+pMC3O71JrauRQf1FGWGCYt
fxow00DHiyZs7s9lXTAaEZmvg9fijYSIE/2Fi7wLrB6OnIsEbc9aiXJZY7WOMEUpDz2kuo80uo/c
olZJrNpmop80XSPgc1/pUf4M4wtwAtBZ2XbybhFRV9TuXkQt9zVc/OmOAfxc7H0z1g1Aw+U3wZW1
4BR8h2lYsPzpCQMCIXZLlH9aL2+X9zPQwI8AZk6fDs2iz4TJATcUATRl/OrCKWoyXgVt16boo1eM
R9f5XHKP3YqJvium6/hogPTfXhkHmnjsKmElK9nRFCsNjST074DjFxRM5haRLnXsurWdAk/RywFe
70+U3/ZPjNt+KcSZYaob6j89/LWMcAsjgsHwzLDw6rmy6NnEKUtGTCy/JaHY/y8EHPghQ48NGWui
GoJcXKD3bvc882ofncQ+IMaPa7GlsveAyAAg2e15BDniS2RRIZK63zLf0UfRlPyLmGGFhG597IkR
nShQ6NNRH6vb9B1hKJzbRMfk+lOoHGNEGRbKpQ9WhpPeEd+Vo45iV63QTcvCbt5RF2JGOez1Whph
rtBwQ7BuRoiiPQaNwk0+MQT6zzJ/IHM6huqnEb9r4nzLiFU77pXSt0gJfKS8bQy9Gg4uH61fERF5
uw9fjt7hLCGSKDGzo/6xPVlLChdKmK6n+0YZ5M1qSDYtK9+lete/wKIWAU/l163U8JGOr22sSnrU
UOUbkNHigciV9+21l/43U1DhoTN9wGXhKiOy2LtZV+IYEShHR9Kb76U9jKx0HvYjsLo1csllHFc3
lekS+4P/lSc95zHnwDuGMTSwSm/ko3UWx9ceYbPZWg/RuEQUvlvM58maQaXLnMpEIomJwNUmWjQl
+Z0g3xf9YHk2jMOFJOpypS1/Tc772uFpSKP/AaHXr9hiFBfpNtjx9RJMmbbGPiws3FrG766zFWMi
879xkjCd+m0yQrusEeqQ93G9R/kAK0DEA3IiNwlWeGQX7Tw3f3+WLMYIQGvUXxBYUV+N2aiu+vHd
1ySwTrp/PMhFM1vREEuXfBwym+x98K4/ajU1Z0a/m7ZXcj3GWIlY2dvfXfudx26KN40OH49oRx3W
x7mC6iTVo6RXFtZyR0ebKRFleTdyV4yNS/0jOurxXFIUHHbB6Y0mBE74xElFZQtCTaPEp3fLFak0
dd65ySPt25a7Yj2oWkF+b2/3A7Do29dz4c65S2sd6zu3TMN6K01eBD7/JDrKUtGiQstkB6upoekk
8H2d7dMvGdU3OLdmGeXadHJXEhwsuQO4FFgxfvgGqdNWhS9x1VC03KUuRI3WL7vW+/AgXT+iY9cg
G4tyHMHNhjBoB3XW9ma8emBNWPj7VWIipWZbnvT/bIa6l8pkolzLcedgA8sJJ1BC3xUDUofaP90L
R4ciK0IfXRQMGLH+3XcVPbgMeyeRWQtsfT46/7rTc4MnbYqVmE9rzNzYI/PLYXQcGUvAP3yRWW0R
7eTQx0qxiqSUZx2V9TzeRBApytA9lIviJku/oXqgxqyr/SRrXd+vfwUt34kzHFWwIN41nPFI59Nh
0eAa41Xr9iFubE/9Vte7OMEgpRbM6TIvjVoCEaKmEl2ubXnpLnrL+VTc8LvHomEQ3CkzeH9gyUJK
B0C9yaoshnQ187cfGL1EiPKBdcsBJmXscs/mg0OdZ9uS6Y8ybyfht99SvTQ53d6evz+jRxx41Idt
iaAU6HyFNPMsyzxcgarE5eg5wLCCKtuK7QXfwyAT+oxP7BeRkJPq9ro995TItPE8zAYGrwn2ZjVC
IfaDGerahcaq2BIdSTQtB9lp0JlgawKzpnFo/+XlZo6JX7YfmmaQ9cmLT3fKlimD6itLfM8fskLR
pXc1/m5FXVymGhgjywYaiwwym/fRaAIHDlVxDM9SR3JpfWBLrcmKmahreVfuWPCP9ZwvWvIbOr2l
vKNflMiGG5/3vd+kP2d/xjDjfb20buHTOJm2p/lV+7wBpyRevPIxyxxk36yd+T1I2y8e7FWf71Br
dBV9lWb7xWcMh3iMJetfDCcRL4PTsOZ8ZmfCcVyB40WDfeBvJuT6BCl/wKlHTz3Gqm25WDxCIYKo
f3s3jo4E8VFdnQ9IrJiOVU13eJgBlzSL9n4fBJrgvxN0fUmb3Y/UPqpzItPXnneQG6uRUQz6jnvz
vu40ft4RjWhBDT9XyBd7Tt5jdW6ybrc8ZQYi3sfxo/touGiA7tF1aJ6tgVkvreYy0vAvLv4siFc0
m16/dNrK6Pp7u2HklLOruEEUfbAbtUNt9CeY3hXl0X/1/ff2ZV9wMyutq5Dhrx7Gc9SflDHQ22/W
INXimgKeitDsV++iuvSQ405BFbA7i3gPV05Yt41QcfS4Y9t2bJ2qfv8x+GooekA4/6yzXG7Dzkvl
pDKvCmqicgcyVLSy7bAuMl2s7Njyzkvo2F0OpKNGmiXB8mqL1VdgKme64S7eJFSlRTvhKx6f2qt/
DLoefv+H1SSP1BVhP/vT3ldHOowTG3h0rKl2OxpfRJN7YxlIa9n1gAM9+gP/lW5FQ58/5gKJ/NUp
xkgl9sxSKRq9cKS6ixalEJqcYNkWNThhD4yUgS4XqI+nD66cDyTJLiImgKybj5NqMIkdjbDMvBWg
G79TOvRReb+Wa+JsZgQiK7I0u3Xggi9DUQdq+jArRlbffEuFQroPFvzkBIJD1i2YIaKla+LwjJBv
lsOYzH9BqLn9pLz1lqSjY/cgtPOPjDeFYj/pjxzfpU5gs48oDVfxGozyyAPnMj8gSmgq39oE978X
XinW2EnbB8aQflwz5/e44ZHql49fIj9+KCLrCrdzD3qsEWmMGeAde5rVUKkh4xrzgLEhcLoPzSVz
RkWYxqHkmJbGmyJFG4SaS95+JYLFGH8p6KaD4QEl1+woHSJZIfSr7zvvqr0FJOwHQZoXXKvf5aSL
W5hjKgLolXximNq5Qh6izaIKAo5G3zlXdnx5BGa9tY/0unOGUfCcByDiDBF/J4L9G2DyALNBggHc
yGyoygTb5MvNXKoBeuQ+VOy/s3ZNaXzCCAXkcVnY4ZQX8MITptW9UiVLFZDEbyBGge77z4CnkFle
reP+TD57Uw80KwPXwxQ4UDlbpq16vNNmE2UgvO9grUaGnBURhFY+yTzN5/DAhAUN6xTxq0TcQ1zZ
UEXUtEkoZHixsv8beRd1QzrIaYBz8oW/idgkYJFRr4e43gPhB3iwxDKR8SkecJXlFD4cjPLXl0kz
OoKnisOHvcn/+cVwp376p0O2YtP2iH/GZNUNRm/Y9DKDtTmso8LFiNaHwHkNn2JCYosnpsKgHzfG
Zb0Z4aRz7/OmXskU5HweujsxdMVk0cdY2VyVGa7wn/49icVNa6AAaX9imSkoNn1Xeb+FXDruCaG/
Jtm48ENVX5IQJLVIu8nyNPEbCHSlAx4tXTcJcsjYLuTXLFlLL/f2P2EGB+CO91BwKSGPA9BgJevh
D4NQs/hV+iuIs/pCk50odfFuoX82tZ1o/KP8sPdL9GsX0GksN/abEeuGykCAxJ0sm5unDglouDQ9
Sw/SU/As+8ojM5DAORiiXFDFRtIU35f1bgyVtQI80RYyM+y5NHi0wKP1aYUvNrLIVqegXZP/lZ+p
/Bi36ZD/4hnDWW4M70u7Q1wSJCpPpSQ0J+mP3qSdFgwcpublFt9dXqpcnO0NrPWgfUWJT1uZBgNv
gQywWcuS/0pPZZlXS3H9WffiUxUxfgvxvCbbSGGiz4fKuLFTI9wUZmfT7VuZgljSwnrFA8JkAhsO
VKuSbsz3SXhm+rIb0JLASmg0GtQmcDjTzJhhm2tOQFPBbdu3DXU0iUv8voPXsGdznwzhtmqTreI9
DVaiPvUbSR3vl4n/qA1S/Y/x4fruVhG3FSW8T3vLPMhKLS5hOTOiwaFjAfa7r8HaI9iDu6g1DmLs
9xV3OH7X8d22y0LtiH45YueXluxq2BbHipOjLtslOc2QhpFn2MoOOu+LFZMTNWYJIyxLhc/4xDH9
uq7UECDKdi75pvzGpoTdbYlsCOqmVh/xn3O+AJwwrjBojw5f4KY72QdhVurC/XFAs/0Typ8zx62T
y080t9sSjNRCuW9lhhjo3Ene8xQ0Elv3n3tOVeCFiRHYhjj02XSiygGDUJZ0iJbqLQjyGTb+7FlY
KnmRHtAG/B8cHeoVyWesF0x8+x5dHr09egsWLLvZBCPx3LX0u1ryoSdycTuT2nQEc4V5SY/uOe6G
empie2McUEq3t3AHVjjTnVGNCNWD38Domc15oHy+ulpRoN+z/gUj/v7GpfYiRppCSciqshPjhrbS
BNg8QFZnzGMEu8pUL6BSFYvBp1jCvnfm8DPF/YR6KniWuMc5sVuoiu0PVk6BE0ObCRY7eQRyft6D
G4HFEV3RPB1ocK7Sj11g2+y3K6yw6l8EBIjRLHH0x8uMCFojz1mvy2hndWNzdUAPRWncdohqR3g3
80lCTojpRgIaSEGXH0nmq/7/VyP5sETaT30wNqQBsBbMrHHd6hvBDrm8xPdiAHu/sBRT155NbDqx
ikMSgV1LH4iqq3nDwaoMtaBw4uKCNT8YKMP2e3IKxQ+aI+OGzHuR+WcpVFqAgjTogEUC1osUBK2F
ptYZ1VlNpldUNiHbNg+SWmDOV/3XmEUGpAUV41p95/efM5AdD4lmpRdql9/KRpbgacZb7K3Kslvg
LonSwVg0xJlqMpyuO1kabxPRrKUp5Hzanfhk0bBZiE1RJ0pQlvzZg8abFr97RpUEQrpgqLAulLfu
sRQV08/zwCZ4vtu9IY57V7KsgrEUbLO/Db0RLDFVVPPZtZjkH0Hh9O3RPevjB23pqt6xENkoGOxZ
UcqPLaPAHQjDYJEpgol6i7UqjCgrrRisTGxfH69t57XqguJQR8v3QWLH402GOvV/tkWebQ66U3L0
/sVTxHjSKBVwHTUTX0iyUHYjtWhywQVARd9UCgVIdLF7hNY/PRwpadCb26U8vFeGarLCC55EmzWs
Ll/n5+/X5buxvJiMkP2C65pBJLJfVK4XDwzS5agK6Vq6kPJYVZ9+SIHOBxzI1DLRGyY7gllXB3Nf
GRABT9bocLCRT0cEzEhkfH9kt6iK8796v5HqbkR6TOTy4EqGcc3WmL2aJcT83ky5UR3JECOlmfHB
ohE2H3rsl5WJSsx9h54vo8Pw8JpdBvrZFctgwRrop7B8iABeWvjEFUvLWQO4ymoFoSSx3aqyaE3O
UpMNjzLGHwY7tKAqMV32bCsqOZLKSbCQ9uflaRGApoI3giDEKuEZ+Q2iH8f2ByTFyygSIk2DGbtL
1UbVANIXnFapKreoHC/TEcCMP23CEFJ5t2RIj1Jwc2jAkU+SQxnzoOE5/FrPlTg07naAn9C57Ul4
hXJlkOjzyw7EPuISKc7dD6LfWpQKnV5sXH4FhUrku0spvP6VznAeCP6Q7T3wEpKpHfciRAKRAncF
AovSGc0QCv0VxuqSBzBCS/0W5Ul3XVhBDJtUT/31oJCHVWiKReJaLb5ktrDhP+VhQiUCNGR//wRP
rq/wbVaDXmYn81o6FsqqTdzU1O3Ka1cb7GTQ5ZPq1R7iCilQ8PfrZpjgAkxRFOx4xtZhYTax9vpn
voO7s6wfB0W0M7KMk3cXb+hle6irhA9QyZrXJTDVVgZjAtg1XNe1maX+athOzMhAUUQuJo9CLw4s
64J+ow2hfF0m7X2diIto8KoPRe6ZGnuDdQUSfswApWriVLe2D0EhDyUCgZNLvk9TBZ80lW/AZmgk
yPBNEvDXrWJjK7c0Oj3yb+A/l+IRMjaNsTSStRi27PM0wZ/6Z9sRx1vNidkXDNaBH0+rdyv2+63h
qXOat5McSe64la9O41mXtagch1Gckgkfh3g8HtkO/9mfFvdcNmp2h/D2lRG/6iCBY6yB/n0VtKyH
67VUnde97DATjztUzG8xNMnwlBM0L15pg/x2nJvR+CKQ3M7C/12kWx9bzGOkRMeYklL0sNw+UFnW
qY8hsPD7QdPoeyPILLLmUAaeRGE7T5CQXhJQkcV8uYrqb9N+sAOEmPzsiVgjDx0g46ZQSuUKirxK
jXg7ojxRG3++4ncJ3ZdjGcBhVsXN010J5pSCV4CXFKKCSc1NrTax2UYlp1Xw0xSjFyoK3Yo08TFu
HjXUttrXDgz6oHSuG0n1AAuL1RiVVdNhHqUdDH6B8Xo0HIzDECg0ckpRBdraHhdCpaC5g5UvtH8Y
iPY8yWwH94O7+mC1BoFuHUQ3VQ9sfS/dF074EfoF35LZe60rHGLM4OhuPQOq1HapX8HozI+kouj6
qmWx62ZLZcc5mZgEOs6R+teEi/XQM1zDPjlsXjUT9VE8zCtSrlU6RCWbEcod+HCsGwW0WVrOpe+P
ZjWjqF9wADzoohfB+gCSQ5AoCsySDLR9o5p6FBqQf2nscIk7laCmCOkpoI4MDNN+Hj972a7PGWY/
wVIU7/n7QJA3+pxoB+c3T771ZjrjaDuTj7UjOa7Ra6R9850vTaYiy8AdVAWkpnvFoj5KEGkfpxFR
SZVo2eSY/y3uUPDpvlXRc31ZoGTYfO+nUjf1m89FBpkoVxuH3oIMDVHHH+qKmL2oH0nhNhu8s033
e68S/l/M8kVLF0W07J3eembO7enKEmYkn2yu8yrnzvDDe742e3Bv6C5eu0rIDD6xwyBY8dsA1CvO
TqDRmt33yntChJ0oLXOP3ws4JZVIgkeFmptLYa2I8o/vwAF9mPBxynPWCEBQS4WJgcOT4Z2EzuLX
uDAV93cPxVM/6Y2w4bFtHVxLte1XoFgPzw37AOpT1zapnwaZnZ/H6Lc4uDJk0024FaLX29fTjuUj
egmNdWc72cwV+VuK4A6PgYZQa0DCrDEwCqwKqRrppfKZLI/V7bGg2YYcV20hsKBFNK7Yf9uNvjP8
0lecJKBdlUqoBT77fgNLAki3n70YMwpUAJgVwfWZBpkNgdO0dMygAxKpetOPmzxb6mWKJS2NimNX
rA/oM1MgwrOcAaNC5B97JCNxpuN8XoPGFi23iiuJvrAegufwwy/9BBexGyf0mQSZVr62/LFA/gKo
stie3nQasUjovrt01JvVKDcwo1Hf8WIrOauA/LN7NSd4OPHXhS4cx5w52ST6TBI2fAkt4HJzbzol
SzjyAhtelTZsBA7WUY0fi2fS9/AQu2Cslqlr138ligJvNazStiujqV+6tLsibVYLJXJqPzC3MIR5
2Q8z6lxWkfUqUg0/oil5yJOUtxyfA18LLbgHx3/LKkYqE+BLPRqQuSU/TVOfX/TTypcy8i+tK4fp
EpwHU5ct3hPMBDlzFns4fcxADXqKRMy3q9dMgs1/grXAH0DC63FAlgpZck4VEwbYIC2RFxIjfMs3
hgcrnyCDrkA/rCkdyzKMN6izWnwKky20EDwFuRou4lMDLshYo6DqBp3XRgWL7u98E/4hxJo7sySr
S3cS/jukiZuRqxaMJIfB/RsiOu05skxPyewyKDX7C11yuRQv7n4mevz5XE/eABvNs3IMYV8wKCp4
qq2tYhf8E5baOBCtVzMdtjuFNh9u3mv38s//ec5Foj/bA3Qm6G0KINI/xq+KnTHhDYJljkXPbL0j
ZVCTV6w0+hLl0w2g7yhCdwY4GnllVUoJM3A4IWIpW11PV4A8deczTqtcJ6KlTAkk99454IVQiqbD
7X5rX77EZY48o/t3hv0l8Dp202UtQxn/PBGH7qCuJV3MsRulKcYo1s7DdiwLJ8znBEmQ747HPgrX
U+7/0wMOCe22iNCI+I0KAiXGImv1MvotecQen5pQM7I3nZWi56eWktI2tjdXbbPce6L6R2BRAtQI
WumCR8gyAES7eMd6dHQF1iVhpj3Icp8bMaNWCrXeTfZfcsVTIWjKm7ZSgiWI3xKM5g5L6zP/fxwW
WcGWDy3797PyYsCLeuu1oIyXhCyYBvljoMAWhl9TaQPa2pdZwYApxWbhtwB7xIh0uCuX+skB0r0s
+9T6c4wbZqMwieFxHuIkTrYog1zF6FgVXqpRPkhWwSLSwvqOk+4N65WYE4ncX7ywe8+esfQv3jq9
+jC3mzCGL+GTuVkgCgVcG5aq2aUtxiQ0QWzCYsOs/z2wfnw+bUwKRbpzsuTYJ0vjTiDHTi4h/qLS
O+YwdMWaw4wAv6eqX4OoBATzbzzRWSWp9u5SRGq97q9D6Vu3yhIJp7EQKN1OWwgry37bm+tpoN99
DK2hPGNcKK8DYdj3dS1FA9ONHrKBSvPnD1sf9bXYem16sUSzDQUp6Ru+giJzR8J31Qfgs1eHpyLn
ACFgprAGkEMpxFRr9K5S598ov658gRqgkRznvbps+gzDrA51uBf60F8cNp49G2om/VGqHoiQESf7
gUA91gmrgIIK7HDiTghwTa75i4p8wi9/RVLr/w2oHKZ1AdnuauX5CmO+Q8mR4So3LrtgXbhZ69RT
W6QV2ETt2sfqhQ2lkZk9vf93Kmj6oZ7JLflxdZpNUKxPCSh+V9a+wOUwGw5SPCS0XRf6DfzKqk5x
rvoYeZCjJXMzvdkrnnRGQFPL0bWvhw/wUOY35PtTP/IFZn2RPozgiFPdvX8YQuS6qV1LRFp+APRL
2YpialQGSg9fTWXfxdQWAlsevv96WB0fB/R05nmXtmFm3+pRqXrRpDymOnKy2N+2OD10DjNXafRk
rym01FKrTaHZiV23DpLYtRu42oklcZvVzTCaV3xN3ojyfCsOrojtAHkiTjDO/SeIpP7GgF/lzyNx
oYGRCK2fOHtNAz9YdrfnHXo4A9XmC0cur3KDAyqqKlru+RfaG5OG4fZ+7Ip3r4yGBNI0w9ZLx6Cw
NSNE3aOGKMsHcZ7AZ34Lk9avZm3I8Qvwr0lVxC1DEp8ikBfndml/TzSH/Vkk6AWg3vMkerGitiZY
SwpddPHj1ezpBCD1oAOoKkhqq2+QAyWC+uFA+0ZlPjSIsdjDWK2Ev+sLBH3RSIn7dmSyTB7ot3hW
f22XGon8cflB0Na3E2+mXSdNF1ptyAHfTOgEZBLa3O637obWB3mlZA7cpeHjLQgsZyvfySdyjrjP
SL/unyTOaq5c7qUjpb1PVN+jq3byuQcpchqdqLNgXgMf8goGYb8L2Tx5hX8jlOQfEo0zzQgtk57x
c/pqr9ck9UpJZxWvBhIKzXAAMLdajoIQzpzzL0ewUvE9xpObc5/z1rRpEp1MBpaAXW++EApCqNTG
KqkskHeL9tKvbq6sxoKejEdJQF79BXe6wIM7I0Z+F8yb6agXeM+lgoaDwdtiYD0kOZnyHONJT8jf
YP+GO2blquTiA7oH9Fzn3G2IG5VnUI7PQR1DUjF3eP+FdsxLTkNfW/7UMrdDCv28i9RD1a/39o97
ojF/0c+LxfD89WKwqYo/rCnLyipyTJ2/qKXtPiS3Q7OpbQzaYADROIUGSIWvPIULej32ErQpc3sO
UBDmpWkc/Tbt6WLkQGm5Suh5+0lDQ3T3IklQmBLZ7CA60FRNfgeJ9cCi1VfL4SXcBDzl4tQV7pcS
of3Qz5tZvmwGWTSrSS14Tx6Rp92aGmmNr3y3bVq8pHgsQ2QJHyyEuBrnqFusbe63V1JOEeYr67OD
kcrAnZ7QmDJxxkZZN/hI2ghCDzco9/2DqmVYQ6G1M0qZNbgENYX/4Jycyu7AVtq5muYNKo6/q+x/
DchBxoB8aT0jCBTP4SS6XduF2BaESbHAHkhsos1h62CB60ru7XZEES1bc1COwzdKsgmIJc/ETn6/
apaE9FpaLRpO9gTXZo7V9RJa5yI0neuq6JYGFdYq33jF5kjb7eDYMDaUQUaW40a0eVmvi5C2HK+z
a0HAovw+Iq422fhNGsww6RDNNRbA5ZGHh4X2RkRTlIISLOkiuuGSFFKZV7+VWMeRiO3xDTsnp5zD
3SkLk8R6Mi/DmZ2zNwBs4hKVq0AvWj+b2v7XoQs1sQryMC2dR15qSVGmL54cV0qSOq63YAp/fDSE
8TPOz0JYyI0gLJ1UEXawxgMVMrSLJEMKY6O42x5duk5YhV5iOUx8u+VlhGvnXHnr8EEZCOugIt9L
kxU0neZqKxZV3bJ+EFRWtJhIxF8s0P3HaYtbhuSbIglovnb5Np53QkdIXvXGHCpAhvO7Ob1XT7D7
cHGqJRm22WFPaqqH7AWnn6ESGZpWkN7JE+Kr/EDgrthgpC+SsKdj8fcMPr87iRjCkpR5OCj7FlwR
m5YnWRdmT4jr0Uh96NOLw8Dw1gq9I709Zc32ZeUIBvJ76cj4Iy5e7/jfa5c1luRCtxkfyNTlF6xz
0U7txePcEZzjiGflaViX1qKKbw4a0rCC/mi+kbN8xc0lFsFoqtE64lSRdSHJ2cXmflnrrOfkFhDU
MP6lOfWkLUbE4VUS6CQmQQGtd8LtCcvPix96C7zlpcm9pxQ64h0ygdQjdsVPOgOt+WdSxOqyI7Y5
tTp8GW+Jmd4ME8l/pw63SRks/+kg/4YBYqfeqZLbYCMrbL/XBEN0ImXDJKSSXXa7OBd/qQlrm3ym
kJE6ctJzkjJzzQto6jJG5sfaY+2CzSLRGt8Ff0T77HfVrmiVpda96wBj3fq32MiINTxZVXuyScRM
JICMhO9kzDiXRLkXCbrc481Zt9Rgc/gz9jXWgL/uo/Qz703dKhS3bmybBRX1ZVYenhvkHlGBoe+/
zavJ+sPqhVJ4R4pI1+V9gfN8zOBfzj8ONrosyPGwMFJ3VvKK1btgaJzUGCW9jvG3Tm6o73xo087z
TQBecuq+piMbLJUvslgGTXCDtJSVIQw9Bi03uC45ejGUA2+e8hacGVP3uqAgDPECI/0jSQHQooXW
n9QZoCyL9eoPA2ME5MFt2y3xl9dfweJTl6LYF6UAQtezTUaKYpehGkaXKBwsGfJUAWj6fVCqWG7t
D4N+i0IeT5LCPRVKXi2hRzawUS7ThWftR1osASI1C4YBf0f3o8yiDcNrh3wsdSnJ9VDteG+Kz+Pd
y87D3KAv2VlAivdFJdgBsdMJKIVN2phRKFKnbdhcPsZd3qx+ZymRtHAgbK9X9hHqp7dUB26t28Ue
Gzv43f+1zk89gXVz+GoPko995Cqzj/qdYivKexKWcrbSAlEiv/u8TlL9m2C8eVTemD3LPc2i74lJ
o0MPpZpstlvLLE14NL/bucIBcJKxRIOEsnLfE7X7AxUydBivAglQlo4j6esOQg7QKPjMX65wj2de
P4Mw2BTwdS/OOUosb1Bt0zK9jwgkO8UVN9CJ+yQo91gz/2tGsrVggGnTmkI8wFf3Y47rRxzed0MX
E2FGgLHDVjQjTRnf69H5oi27AI60OuXthPMkDPsFzk/Qj4ys5MmyPXSJjq67fOOqnW55df9hEUCI
4FDAKXIFr6vWjWiwibx7LQ5gk9EwBoWo/RexmcWkYeR73N/w0RT4Cm39RFM1E+Xhjb+ONn8Bs9wi
QJVFGTp9jhLnIXBOWNofugCbC+4wBKoKDZf4L1n2hiwqpwKUn5Jc1jJGVYGnWLSD6c/RHW7IAzJj
yxeJefwiBjFIFbBauuz/2lZ6hQb4jBnm13Is3NynbRBAITTbOivd0tt+1IeMVhGMOhJpYHTxBFcI
gLp3ugoofLvsyxl1lBAOW3fMMlCHOoDhVwzr/YQJVXlIpu9JJcdzHzRyEudohtOdpnqBg/8HUo7w
ZI4bWFHNZhtSJ7bosy42m7V1SK1isU5UD/G2mgxFW1VWbFhsebxYO7ofHqfQlASPV3y9yByTGD5I
gpIfT4Yyri0Gg3cHWjutLJi4gKuezgjDyKyiLVlYgU4+CqAR2+bHDDVJJGOBm68swT9MerZcIqLM
ioR6lX+ooN9AIVDHMT1hqM3KxLUstoeDpZ/bzMHvOt2kyzEEgDo0aA12pahk4tE56FQESq2TG1Ya
MJfirXeihjFbo2/CCC0INrl8MwzVtULYn/M1WSJakALiU65VF6MdTrqIPAB48We8B3JEr9+GMiMW
rUq3rE721BTf9kAzpVCYbIazQLHVrZxGshY5qK9NJSGQjzBYtY+xN7m0t1YIJARIIdqiNMwwHWph
3X72fxnapO+6FQ/S72pXz5at07jAfpGgQFIClo9PaR4pGx4TbQzAS3F1XQF8n6bCA7Vp35VViMSo
0vzEepb1wlqqlkW4HD3qboFxHhx6WSBx3lH/ajpS6+CAtHitxhCPI+ZqsLTLyuzSGiqgoxNQzsMb
BdpTINc58StrhHDcbpmHfnjYkD4V+wlel2e/uom6vc5jy1l6vBXYcnOhZF5JOfM7DyTXZW0Ibi1V
MShlmFToUFlwtLEqPWptdU6w27adMh7fGkmMKGcvLQIbFFgklCbm87hSJyfseXhj6IJHc4B1LHUd
/RfUDNRGkR6fLV0iP3YcXmIqJCmkFARThRx8WibeBvG2YV8JdDeKsG+QiqcTyX61pzB3T+GTOxzO
qoS68Wh/s65OI3fTSQQLSSMqU7VCNu5bnS9w74heSctflVmhZvFfiBr8XCGp1PmfyYlFAkh3r7+A
vgIZtEpeTlWvfHCRR9fUCK8HElxRUvRfXFa62oW0VnererfnzBb0vCq/tthttwUmoPVC4SrYTmgU
HCtjkPe5UekiH8APCFj0SO7C2A6wgU5TqBolNjPFBqWi+mX6Io0VK+TRA043DzRS6uvyiD/CsMl7
/DxhLntBCcyl+fmY8pfDqtDum49BDySUTZDkhBepwC4805zqbyAaa/vkP1QJVSFfHSE6hyNHk1Gx
51xpOeIWgmGVyenboUAAy6eZHwi9dmRPHP5SHEfAU3+MpmNGEhgWpf7ImivGrZCMsM/CDdfynP2O
0d4Kc8Z/6fUWphSS+Fo9Qrqara77GyqAuLmGaSQ/Mgp24GlPVk34KkOd95cb937CU+Uu1a3YSHrY
oNGsh/MoeSdBFiBBkJ0JhiuIreihsLYIdCttSNIoYufD4cVI8aQNvPcQOGgzS1USzHy5pe+fxXVD
dFG0kS9+2FE1S7LO9siVEXxpNDvmPDxC/SiCwEge382qc+Y91nbUyl30B+9Cq5NDAStw0RYjrKjr
GncYxiV6pSjqIRlG9eYbBIF1KzZtHVWX5sE8PSaBNehDY8oK34/wec4XAC86gef0QyVVMIDJRP04
+5iLFG9VXCjp4GAiZtgiwpLMeBwlUjgxi+UpfT8Pk0Zc8XxoBewmKey3QBFTmpbIqmKqrm5g/ynR
VI50M3FUIAJPfFFq9iK2dMaaGs5NNO/OP6+fKjH6ZWYoCpmlZnpuXPrSrOiI08NzCFJPTTssTYMy
wX26rpipidSVKELLKV3z4vlM6Ne2Mu8H4h+j+ZmXcrqak/p2Kf3/1SRPRL0ImG6Y0Gy7coN789lB
qzn0N/b9RHh7t7mPsGT+9yl0sdN59+bPaLKjyD5skc7GnuesgH4fQkdoDAYg6mgvaTACfNV6LcQj
fs5eiKoQsURfYSXHMqCzyadWTkuDRhRZrVWDU4MeU+ziGFdA0hpSZp/Gn7kc4l405e/DsTSXd8ro
Z0ilDkjjPTmRSQGKN3ILCrVVZW9rYNG8k2ubIPdaT42ZGTjqvZsIYaOWQm1izmnl4I18Yj/jb0c/
kDOSyKy1wJhjarVc9KXGa1scqT9VPqPi/TDhwsjjociYPNrLRK+Ui0e8NW2lfgkS9mBX0LZPSbad
OlPHQwc+HdKyOrjft7dBYK/Ey+tZvSXR2d4EaYsuOKt0SYPiUrsPtu1TbnH4Za8RzdUAAMVOnJD1
Z/GeBr2rj57Xj2dZmdxogCn+1ELKMMjHdGNxiJwaz9QxJMxfKo0NsfyB/jKURiKWDtb/kK03flvy
mgRqh+0T5df7NB3T7Q/5E5AWPyiF9nn8JQyE6Z7E90BZRfaZgOj2MCYRIB/9rr7GKq3wNVovHzOD
OJMCK8HLjF1XIjrXvdpcfEdF3LIKwH89vW2nBpoxSqXRITec6Le/MILnP/nr+QiWQaHzKnvy/1vs
da/a2qxrV9jqvOkBx+Lz3J+O3xIEWjf+y52yV6tokOeuSctKbSt9Gys+8TTIJJh3ALjBGOtEE6dB
QcEv01/w5yLxXZwK+YsxpeVsYex6aDJCTV7M8dGJpinTodq27bi02GlDLn3WEXTstzxqc2C9RAX2
2sx6Psv0/bFcvSd6KTjE+8XglHe0cFhC79aLqZtY33m2jJZz02ZYsPtt/QW3oehaH3h3kzw50do8
S4fr9UA2U1Zn7znX5uDu/LcuFmKpwqvTSCsKoZon+/PJpnBGO54tGW0ioZlFEBzE/9maBVh0/Sax
9CY6+z4BqOIZN9nA+mEcpdm+64LhtqewOT6fuYcsym2b08METjEFvx016d9KSwKE6hAtxg5L6OhJ
ToqsZ3yp4RTYFwIV4IpJmdwT5taiWURDXZ48LVrEJMXyxXtZSH68eXD2k+dcGNd2eUqYOZP1v5JT
p+Vhv+pvgub77WIAsItseR5RXchLJ0ubWEksfScO5pJ8EznCHbsVfR8K+5gWwHhS5x4ntSWpSwS/
4BMgyJsJFgFYpYl+bkYEI7jGGRxSk7kLkPD3llnsLaakL/67FCZyL1K0foTZ1AE5NqrezfkcQ0Xd
0oaRiBLXbyyhlS6kqzXvfzz20fudqdH6JS5V6RdE+fcvxQx/Fz8+lEyzHKGEgeF3+HYVe8vWCpfY
VPXz6avatZ9amPyn+tlnUps66DaGotK4MDR+L2Wg4tikJS62UB68Ys2EyJOcRuY3Wem2lswQXA0q
uoJjhjqsZ3SR5AgMVbemJiIjSw5TcpkoLTA5F6Wt4cVgODjK5rixVeqZS4Exhg5I60cTwFp7kYCM
bMfVpCPbae1cs8eVq0RUyhHOfK3XIRWrCBX96aDZzV6zey1cpzuHLlU8UDtUI+SR7CY2ISEuxDec
SiGcNvBdQz05ioc/eRHDUjyIH58Q5OjcGyTfGJfBfw0KzjPepCXunMz8hdeDQQmH8q/nOBk4PF9G
RI6cqKecyRR1OHC8Jrnxodbmu3UcE32OU2TjQz+AOmNB05MpzVpDLyYeSXHyD8kegHtNXf4gby1l
Q1P7iB4UoJGA3Io8FHU4iJVJ+jRTQy+P0HLYGbm1kYLGr8Pp5JGDh1w9yhXA6i+fv53sX7vbUBS0
QsQAYbZzekiogto9i6EWkP5tRbZMgGMS47YgRxNyNBrG7lEnaIDdsBNsltNCQDyzp8gH6vGESRfB
78U3cg2uNU/EERGt9PQZGzKdewq7s3Y/80mrfxGrOkHWTq/A8WgGfpZwHzv/aEHZm8SWRE7GXPg4
+ufDkBPoORNO2JZe/uKEbf5FIqTnPKy+gOGNXi6BNlOzuiXpuw3MNWuLuLAm0B4t1URm9CvgdjWy
LbAqdy5XsRX6DZZ/0CaLlPPLgX9R+4G8GkmTN+4vS7+zxNReYP5TNSdYuyjtzVjLT49KOl4sKoyx
cmuxvzuFSBdXOuHZ8Nt1xG9ImNxX1r/iKbip56MBTA3V7j9RWJDzIdOT8P+DZSov7YmuJOoblS65
AtOaXq2/8BREMD43J4TSr69OFIQ6hWrXzln4mnezmQ2rTzWgXj3G6AbFBVBfHb54IzzFy6IVlDE/
KJABXk/bRddrwg4WJLpUeP6YE8xdPdsUSk2z8zLbEouqW0qgBFkocLnobJphb9HkgkP5+aiT9jty
zg15t3ktc9kcMj57rWLzIAgLNWlO1uWBNVNWsEONnZlnchn2f9fSrWi823SmmTOrS71rhXzqPWjW
e1WRpw0W5IHpUJW5RhWtYQdfLQxCUOIu/OV+neqa7+mrC0p928gQYyZ1KBdLCofi+mMqBxYtnGSV
tTLxW3AGalr7l32TKM+jlAf8KeqhKb0xoUJA/wPTdV2m8WLgGaljaPiTrHZBsrxKugvzDrhj9w3b
vI4bKwC4zhpbTsaJOWAZhPRYZvVXtK5A4ZAq3nj/wHBaenqEXmUGDh3p4Jq7yum9lECXmN2/hC4d
JYxT07I+R1Aes/OE2C+D5h9BdqLIgw7UGxSjDMXaJfJuWYDTbibPMiy2tLV6pmzBM6yT6E5eCrRI
Lsy3X6d8+l2Hox/Ijvgq2kyTp0to0m4Os52SlZag2dc5wRMDUxmbM5fmOkNb01oXTcLdXvdWA/kf
MBYpAO/ZFZGdRCbWNU7HjK3K/zDNmlpfiH9DWSjjb8TKnKOOy3P7Sxnp+JD81tKGDTAhnZlB1Vgg
5Qpb/MSuw8bpIaVulDynMtPEw0/eMwVqEsFm2NlnDNfVAGnA+HA+TJqQhXBaB2g2Z/dvspblCrWp
Mq6JpswdY7OABx5g343Gd8ZQfoXZFINkd617CAru5mzqwg6W9hjbVN1m9aE5qKqU5mLIHnwcnKUQ
ZDT06EWz7ksF/o9ochl+8bILbWc69j3rzgJNdjvWlBQHdshgpWyOyLDulsvfvvx0c7dnPpI2pwvB
/ud5qE97h1eglcKfKyDsQSP6pKzxXfoOkeAhkpHV0quHMlnSkqL1v1r8LpUSTB9slhGcJFhCP2i8
S8P9AJHnZ19A/ZXUNfRulCFILRSLdvQCdhsx0GNUMDqIzoqrsJSZF1lAinoTVCjRhGS2DXfOWdYn
ic8Q0RomSM1z2weQvJLqdAlyV04UyFUzWpazB3UHOU0AK1M62jnosH7ul0YTG9OI8HDY5FCIEZOB
7cLCqUwQ48Jlo1VznrBcEwGBJjN3tUPxRFZh5vEDvRY42NtdubOLJLLI99xLD4DA+kUUGslxYwXp
tF3EOdzBcWsc1d9NbT+7wgQ1gtsgrW8t572Pz3+htvH3s1MutdK3v5XKTa7oiGRCPspZB+/YIKDc
rJkriqNyXMQ95BaFHvKW0QHnCx+Beb30oHkek1RRqdB1GHb5ZA+n8hX+Rm6cJPt3kPCtCOObb0IL
VemICFXkrIxbqz6I1m4KBCPcGQEJUMfGu7ZHUKA2ZRIrcodjg6dsSVA/5CuE2ECoLcIPg8+6Qp+J
VPWzYiGXkwCiB/Cj2Le42YlczXBJ8KeO2LtTvYdJT+4aSIfWuPt6yG3MuKcLUHiAh3EY3WTiGl/K
PZvRx4qQRmV1irvmdCpB/XUDBJzTHEtcOmd4ImX8vl4/9ydcJxAsKvtFgsNOGvws5n2Hd5kFl+Tu
+1JrzD+1qYMFZMpTedAzmtOZ1y7wPXAKSostoDEy2sNpjDMLXFV54hbbq4AP/rIe+WtAv80Fz7Kw
NKePx6YLRnv7hlz135MlWJXYs62VVQUyWcWrUrMTsVP5PHC7APM4W+dAO0DXkhqUHfup5GUbKw/6
FRKRUu7dY0yPUsu390mwnAB/weEX9FEIXPUnIJeg0o+nGMMm3hfMaMxrdWG5AF7piBDTPVn3NvR3
1DESYjaG9q69KG88IDz2pozwk8xGJphtgWSaTPGkzLxThYCrZzM4Gd5OIAvaBjAZKQfChTrWec85
BCJXvXeE78H1IhB8eqMSzXGTIa1sDSAFnldgBjf0qigrgmJ+n+rHzcHme7qRZdswcMNEg9kshtvC
Zrp15buo7DZDx70zPnjAP4Az1SUn6OJ+/wq+wQlMfG7ZEzoTONPDeqNA+twM5g78Hmju6Q4jy0bz
x+BIkUXYzu439UnkRdJFc3WbmL1eaojyWJum7WRfLzkqhEn/o1TbcNMOMe9uDpy/f5itbfLw+3Sr
xQNiwnMAK9SEyh0/ZYndvP5EWuzxm4jgTbtH3rdvofNGQeuz22TZoicyzlLF7ZtVnNlHqk5PyXqJ
8RCH5N+4ySzDP0Um97dvs+kRVS8Ow5zvSYIEKbKSh9HXoKEyW8JnCwcSQab99jdGinHmzJwLlEIW
t2NwvgKkbQpGeGG8QUu637ZdwVJK4fCSefFdfi4i6w3yQDw5kI76ucxvnhclmQYH3P3175yFJyI2
BdeVhQ98fqKoBkHZBdSq5L5v2HR1zHAvyRLhXIinLKz1vxHUb/U4rF4Uw7qN0a96IBFAsb9ThA31
iRxqoeSBc25oOQ6ViQjLk1KZXT4SCwArjr8umeG9TDNPW1TDtcWLq5gvIuPD8eHQFOiCA2VHqPt/
NW0u/GcHxtQAxejlOsBeBiMR1TGyp3jGMnFbHuQACg0h/l++kIqL2beooft0vI6jROmoOnX01Ade
4uSQBWonhubJFnVRtn1NmGIzuQNnaEIoGO4MDh7cJf0U8E9/fP+JLBaSoNmtpxDynK1zcixj6cI0
YdTg1kuyyEPkb2obCyEH+Hq7Xio8e1J0NPcPwZHuyXwOZtpq28pSzYuRBaD7jC+vAWtA8PzQFdQW
b/L80KZTbWD1BT53pXT+XWlsLd/W78x3AewvQ7nAJJ6Of9GnLXPbR5G9dbAETrJXKJg1ViP5cfNO
lILCXfOWBPhPP77rlKzje9d1BrYIXx0IfoCy0wp2+bLCINqKoBOMc6AqGOimYXoPnUSRZVBPvwJb
/szggI27O+A0IL+RWC/edO86/2vCExui1jgfJ+gPNj+7g0LtPIaY8GZ/61frb2XDMeQXtlygkkKW
NDZ07KYxEPitQgKIH65lFC4+9cOfZCErD7lt9mYWn62CwD2SccnJ1kl7qCOL5iGxijLfW/fsEbSI
P3QntfXPrAt5QKtKMzw/SOn5quLZsjxY6x185c15eeg7IyTL5KuFhmPNw5yac5rC9XJJTM9cmHgi
F5Kg+JvpZi1NnHdrF3RFXImZCr2mfkm0jBO+40GVJ09TES+o203EJWdFk16nL4kbiwLr/ThwCxss
6RCJDf9S1W70waQeOdRfeKsrqjKZs1OZioZR+lDdje01+ruNLTaGbMfKPpqoZuugUK96keY74xe1
FktnfQhA4qx5CoyE+WOAynlPyxL74tQC5f4IJvCSOIZsShO3dcVuFWg8KCypXJADDsqsjyxZboYd
Id7+tjdc9/JOtgL4dpjEjU35lb84xIirpkgRVyTNNSnjbJkN4ecnMXGV7lO0l229vcJWw22i9GAu
Xb+sL9yacCHp5sYdBQKxs0Mhg8cblBIHfV4IutAgvNM82CxLKkcKwPhaPt+CQpB9SAPgBvNy5H0Z
0GfCI+30F0UbM9vSpHhl5xcZBLBv7QCmUrwjH9b5YXUdAsUuhx3DvTf1UB+NJL/ZZk9eJZ9Q1SCw
/a0QzJ2CKWa/JFIJpDAXugCBmL+sg70OuiZVf39EkFLPn0V4sqOUvRUOwuhnmQ2YEo+/l87hGJer
Un7DI8ui5tSYfI4TklVOENrG5Wp+eC+xuZ+UUgVmGEiY9sxNgqnGDDNCTEO5IeLMHdkOtosDTI4l
Mb3nz6B+bm8N2UgHf9GQ8sFmlk5gXkRq1lYX7GkKs7mOxyPwvlZRTwZVCddbnsCOjVrWKIsv7mZB
5mB4AijGhTDRFohxM3pGjHqQYhyLYbUfbsfHBWi0cRxlhj5PKQdUD3qUnonuDrYBPylaN3q74z/k
LwiAp+nDSvsUBf04MTz2YWdZLK8V/fcbuadk3L/PUnDt41OR9sG1NEVu+jkvcTJZVBK8Fc8D6O1X
H9e0Qx5hZEe/doCXznOI1A5SQqI2avPlj9IDmWizgjdZiVq/mEa81dCAlbpJOvrS5qmmFVvTkMWK
JE9EKgJ/pE2lFrOaDAFG+RrgfYKG1BDe7T/EzN2l1k7A41JINLGwQ+h/wa4gT7MnlJVk+6xettNM
22T0kTRUPgl0gIzRWKLLW0QAQ1f8PUDueldlVfT/LJ62IM8dVZ7Y1tmE7vU6XSPAVg9cqZ1G6L7O
vGFvW2888f81XpA57tc4nBN0GhdlQ2B2ZlVPtKGl+LdU0yFeeIDKVY90Jr5IaI5Y7k9970IKCrQG
kmm1EsT/iagfjylElMKji5gII64uEqvFPETJR9YUtYkUIdbC2WaaqsYM90Esrjqo7rsWEw5/SgVr
XHTi5sE9uGmG67TpfkdR3KwBI856sUu9Wo84+IfRuPOXzdFdxhgM8p8aJhbfCFc2bhL7lMuj+p1L
tpaYliYBAnfHFvo8uOK7o13+JUBwxQv6PNsuvvQ/b21hxVkPnhr6Q14bBtmycNRiTNMNHOtwX/vB
2Zs9n+Nb9hdHn4KhAloph7hzovf8cTqAbNPnTzXCd4AByCsHAqZSqyXUtjW1LTQJPOI495SwZvgj
QM/U3qlfGVM6v81Jzi5QYehiXpXchEGyOX/Kv0wOsackZ4e/mCSXQBrxOFktk7r1I7zaT6lbJq/V
/lzsCw/tyGaVx/HJZxFZsi+Wio0hO5qMEUGRD38ERzdfh6Zcz6zVU3/fn6lv5UAYWkbg32OUtlRL
uhr6ehvQMp+OfkQmlayQMzFm37ce0cSoIolRJCGjBXzg0W96pIfknPthQxEpjkelwBAduNZoBa5z
wpKNb5pCwGjUe3dNxSXvqq7JYNXQYfdEAM66rh05Sq+Oq8bXMhpCR52l1jraM7J8pCsPMBLopgDp
juis2AtqM7UcSYuNRcIohzlsKDzYXSQQe+KGgNwB6GOTicPUnYuZ6E9Q47lN2QTIBi6fpkpZVSgO
jExMi1/jcjCDy48IT6zPzinC3Hh5kk864/afKvJfV7TKt5VJi2LloJCfE89SYfke/l2MAGh/zkd1
izB1Z2AnRayq6UZUWwFqweBB0SkEMogvwoFe1W4Q34VbXsFrDay0yZ6NiNbz2Mf0RUajW53HFlM4
eU9GKWv3JeqkmmhM62WqVZsBrrUyKmKLUAM8txSd0uuZX11Y1DFQgxiBiZXp3+52ipFikgQZcOeb
Cse7oZt0hifrU+lOUTSTyAUurx7hsZThuJidvyiPcCqw0GR35AE59VvXrA7lardErC5bq12xVps7
oNqpBA+LLGWfkKL0thzBbd3wGfOjwzJ2uDj3OOYIdyumHPjOxIsWR92K/kUnoGqhU7OWDlQnAwLv
OqAYjON2cSFx3oWz9k9NbFFR7jbUT4GOzoOWIv5oqTKuL39Jk0FrgFIPQeQSXO9XoNdWPEk1hGDy
+lczTdBN6hI8NTGftIKUI09cr/IdkSV5Ap6PBqUGHRDMdtuQbedgKJXn6RBSX8qS6qzBRmufQVR9
+SFs4/B6QW+2Wc2xH3HFyX9p03okcXMvpwuZnN86fi4DzIzrF83b1E+vH2ALhbjQXM4i9hY64j71
LUDoVlNrp0M0R73f4RpuTpZ2afyHjDrtlBsE6KS5h7fgA0YJCg1sBIOHluJOPoM+hYb0wdaRiw67
2CmVaEwIEShwd/2u/NyfBhfctoIkKMtpChPX7k5j+psjoWvaTKHXp9iNH1CRkuOvT4MqT0J14QGo
cweZJ2Po5gKrr3gUS24/fO7kKq70F9jvlnDRrjiw5mkx6Y8/3fmAsrKdSlqyKFP7ov660GiB/SDh
IQiYVnULPngyLsJLqAaFm+4x8apBVYxP5pXQYfcFVSAXiG3R9K74cj5S07rPWbGW/FiAgZ7d2yWx
dWN9DhqGfyqopz8tZ9CVPR5xWw5IUj6AbgEghfW+Kx6SYa5JcYUL+s9URskTKQZmi98Rc8UnyioC
xOO54zszr/yW2KpHuI4k2DsR/VuUlItXXHf+02vyJiNCAtDfbyen+TQzogB/3no/jpn4dJ3rV20m
8sSiMyqqtKnZ/OnwNnxqj0VGt2vvOrtmPbis6yjA3aeG04ED6fSn7CMrDDGaNZTfBVV3k7fs6pap
8EJsEkssCuuRBDx4HoXmRqRQvGa5Vp+L6KsBM+GqAYqjBKQMqzyau3vJrb59VxvWlw7PlHQa8Qxn
ayIM/tsToyQl2Gcd3NcUuc2FkcuvqHZk2qLj3uuehYUZ7X2/CGn44cmWI46DHHqYdHGjy3UlCFSm
bK7IRfScPvZlvFwZF72xVMk2gVC1ZxE+shnU9E3MjXekPh71s+8KSBqnucmKhWNOQvz75VYfFjke
qerQwaDaEuOxJgqnVFX9GK6yTH7fdzfEl1fjlacT09DhpcTYr6jhXOc+RYCZs6F/tr6gs+WcO3o5
z799fZpnKc8HsRg5luYv74YbnhdOIam83417gwP0bGQDXxZwA8foHBe5qcPGkheTZzlMMdJZjZqG
wW7+bOK2BHv/rC0WIcT1zGOuy5YuDGIhtdDEM8+M+cYskCxp/xvybJjMwGzXefSF50oRzxtZyBOo
tLxHWEfvADOWH4jCCdWtCEZ1tdkdRYRvSkPn3uT25AfyrXivrdGx/J2ERCcKF1RKba1xWm050lKP
vWPHDk8fnn5WrRiUkTnhh5HXr2OD6KV/weU6qlqCtE6l2isNoOrEWsHmnQfMA2Vmyg+Q+M9WYTEo
5h0t5CVpMkmR1nTJBl1vLXwdWWmVqdDql6M3AaOVntR1ZCt8FMDh3576yOfioqqvKFDOOgiswMG5
rmKny1M1m/W9PDhgf+vio1VCcSykN7vJeu/N9DMm935teQAtfo8+TFkqeeu19LY+xqjVEDtqyCbQ
qMQP7MmBk8ijY7I1a3TjySjUSgnAwXxSyBuQQGhfOGLwALboC0cgZD09fwgnbaFKo80FblNEcgyX
Jyh5vkY+bYwtlq/mvLxx53allqyCLTTyMP7e7xwPKWNVtZoSvkTr7Nr11aEXOzBUXVh09BwyGNib
MrEE4znM7J1PoJrL2DepRbrSwwg1ZG9nAKNLqOsbXW3PcA6xrNt8iwwwTYhaZPV3YBF/5rH80eH1
2+hFVu2/atqI8nM2wVrA+Fwc1piapRfOmJFhb7z2A69N3+sddYhqdHnqyQLdzSLyxh6/NK3gP1wG
lbmJXLYREp4Flcn25po+eiL4muAk4q8n17UE0l1MtGmN77UlkmddF9hechumLQP6teCt77+2K3RE
z1FVft5EYRddrmPCluPOrUUUexpk/617AxhqmM3ZdqfXM5ZFkwch8QhNZRh5UVI0LiNUHC8Iwg5e
qeDU2JsLARIz/pbTrzzBCaoq+MwY1VzGQrQaKMnkoaACtJZmQGwALu7gOd0s7btarGBN+YFrrLWg
PEK+2MRJpWpuz3Qx8RcppZKUfBpy4qnw2aVGunbbAKu9PY4A9bWXbJ44CCQlBFhHQhegv2djPP0V
N31v8UIDpUG0hVFgQgiu5DOIc35fpW3XsgeN6bzORY/xPs43c0xVWXoX8G95mUE9eq4KuZOKHKAW
aUeEzFC6nwCCwaZOEeUnsBN1JHiVQWONg4xA5IYO0+O/W7vzVAeDOkhWQf30V1Ch33rEdYV9tHot
OHhfwfPu8xreueIE6iK4jsr6P5WM6MOcm4Idz5sRKlpgnjuztqu6knJF8mU+V5iEEs8vIJusxcI4
Mglc15b8o/4hdGRIxUy4FCnVnaAR3E3RMN3U9nYaqHQSlHukgt17HJb2W3MJw3anE9TRO12Q+Y22
9RS501a64Iz784k+k9iNQGfb4VFV9dqBroCAYkBhoXfGbR+esrWMDI7r8+FHgkGUqRRTw0jAgb5Q
mP+I0C+7u8PPfjb2qx8xM5ebwHFyiWlWzDSNN3lkjzdIEE+uzDqnUBh09DBq5IqAuwyzWrL1Jctm
l++Cbq5Yzf9xO53E5I2QQJ84RhZ8aN7h1rZI15Mpko/4YjOl40ePS+PcrUSbD7bMuVyS4gmpMHOs
4r4uBeb9lAiN/n3u6PI/b/i2spsVkPpjQwW6bCCsOeXekFtdewr1l3zmIx23ZQuTicpJjBgQCPHp
fIfhh6TNvk551yAGyCBWSwDCFZ+ykqtqCE59ZJq5UWh/efoF0CWzQcpa0imYVpN+rFAKen1QWapN
FB1+ZDCOn2RSJo+bBFHUKOu1/JyQFPo3EHKJ0JyioG7l5gGVfDeF7C5TAEwt2xEuOOFVZ/JWRCIH
8AxtqHoZPLcpY6qTezMtMKQ7hhjlZmkzalG0i2V7tIND9+qgutfjJisaeFr1wB0Z0diCQ4eYgHgb
XYPXHteVVHqT3EaHveCK7RZ3qYOknOunrKt9SnVLGaBYQQzAwm4dXhGpSRfhH3hmGCcTiLW3Acq8
f4zyyLX9eUAy1JNYvJqDH7UwPCKXQjs85+yLukU23TzdnCVyRziN0t5J3sa2wjoU/NOnZGtACD37
/IiCfOrL+2TQzsI1+WLWkPfSY9rAgEhdJ/1f+tw7ZB9foGbWhVX21raZHZROfEEe4CtB675NLgzA
kbzJ2JYUMTcDmr5wwsCl5+7bs5Bw6jtXDoERvrmMD9jYXJzP2NtMN+z8+mn5Xr1dspyDWUAq5P+O
L7ldHo9Kh93W0MNKRIdZwk8ONlT7rd/JsZZnghr6tdFzvycO+GiWKx/v5FsRmOwQ6jfjBhkFGZ6k
2adB8lAAkvuc4zOfyRvJcu9jiCGRF6i6AsxZF9aZ8ohKqN8MSegfEuu8Hi7iGFcwJzTW1A5v1fEG
LXzd2JXMPcA/Ra7O+RQR39OfPRLR9Z/ZI8zYkX5TkHU9Q0GzoK3mfolqNgyEb2p9qwDfgL2R0HJl
jBhANtDbDpx5y0zBkJUGcpiltSLUjZIbHLM/w4XzX9RWo+g2k4/QJWVqe86sFaSVM3WYvlf/UQDv
JL1TvpXz2YpzIb3MpMEqTbZ18F8xIAn1eOK8iZYOxzT/qpgLLORtDxF3bxmqVgpOpQg2irirKlXF
JTerhmeA8/pde/L3cJzOBGf2q9ED+Bq+23tfDx9T8fiTpDj1Vnanee6eFcTPSwsQXj5m82iELecv
raNts7O6JeyopsUaZofiMp1o0QqbhXetWeVk88U8VVtW9mF7tGmSBzJtUMXTP1lCuTw6hLE+HSr2
PmSlOVl8/qUWJdjRpykGeNDfRXRLrm35foSpAphh6x4xBnrAR3SWOPQON2kynxk0cyj7BtyPVYhd
4W4dKv9l0hE6PCaQ4Hdd6gr3rCu9JcdJK4Oh5RLckAHOx8VdZQPJoQO2ex9xQ1lBG6USvHx/VtFi
6T6eS02KgYedcIP9MwikDI2d1+se3Ea/YKWe2hB7vW/HItXTn9+F0aO2GRtj8Ga1X2GyMh1x7vrF
/MKNZvNyryGrFpSTeZCJ75mZUp6pRKrYEDu/2Z6scLlLRhX+0r2i6/aBARTN94Xe//U4s6Y9G4D6
X2t+0bixIW4fWVc8D/f0ZyCIwv9KENXnCjZhtfRCENewJhk6yrgXxmJEHS4kH3f6vbbhunE/MOwL
oRPi1fwgrU2Mn5HIkunf+pj4CQriCWpCAEe6lFUAvbCi8yKIPNqGTZjG3j73/XySxzr0uBs/eE82
NSEJQrT6AQ9IGoA4oneaZCQBB9sLwOXKLRFJEnJ8WpHeS3xrj4EZDw058/5XEkO0EgyqoxKicCJ5
zFVTCYL+SO4izNqsysisJiKbMrypkdW01HbiRnxCv1ubxFv/Joq3Yo54v2ZCOe/mKbe8xapcVa7R
HawTsu/vD3PhdI5qrYo4qA5ZehFlDXLEwuM83lsv4IB9FcDrz+zgath/eZII1XtH4fW4Idftn3L4
wf+QWC9wLYod/q5PewMHtCujOaR7yQWmtv3FjaWipEGTRdY6FqLVaz6PkYEB5p5iDxnWAdMY7jiU
ezVAFbKsjCexIHyQRchcAxXXYgkLbtITd6ClLC2exkIK61d0D3BTUHK5N8jJ0Fr35iPP/xxV9VFo
cTta0F8KEcaWrjicKLUE/w9/OdyWmtudW/g6O4mlAPoSiBf5S/cmnCRxSOu1TxJ/BCcgm8CJVZQB
zxlQTWBh7IAVRBjUMMKOV/VwUYmEQt0+g9qSrO0fkMGxZ5ZB6E8aWtetd2Nv4Hul/yRFFNN3SaT7
m0EdUGLs3s0eLwjjPZrHkdHR7kkLKb1ge9TQ3q9K7D0Vp3iYoOAUzfDIi08Jm04tkEukbvbPOMTb
HNfNFC5/20FpAFo654q008Bn8t1y4Xf7GiomZhSDcig7K6fMBxDInzEtP37J9d7aMTmNUpJ2//jx
PjZ796b60eveM0x+6pNKDeZ9VaOfUBRO1mvsrMgnFq/AsYKMZ4/wLwVrOVo58AiwUu+WRVrA+pGt
CyQiHdnjx3EE8/KGsHhwv79nID/oankH1DxLc7wOze2XJQiBPcsC4RGYyHGTqFzW6T5r6XYGlCmX
PgRIHIv9+vkHZ65Jx4fQx/K5Nx1jruZTABEkb8sCXuANMK0N3FdtoqOdwSey44IZW+XWGh7p3m6q
z8+uFag0/15m1GnIld8xl2buOnxESESO26Py6EFiwvXWs2DqcABfLgM9pkurPbKQjfB12N/aywEg
6PyT5hkvxiEKs1Ju3599uq8nAXm+p+tTlDf7dnlZzCCWYr5TF1xKZBeBn0ZtC8Q97K7vy0m9OBIg
1g0WfRJY3ZfjNppK6D4ZW+X/Q9RV+/XbYPFB63zoWkY3WRBVO+angeYKCMJ0MPx1oyp81WVR13iX
pmy80A5dfOElBcBd5SqkzC9wqEqkBj+hKIzorlhll+8SutpMEt4euR8mQ7/NinND8dJbcS28Q1oM
fn5bTMgmytLCLjygUJjCMY/ESRbvJ97LLDqeWV0Xdw0DaWBzsol6bSPYOgB1f7NjKuthVcnZg/p+
hHcsvuXNfVFq/wUcWPb55H1UNDJhacyTJ9JeSqMYrE0RYlwXOTuhM1dXVVyomPnkFl2S2vaN4wEN
/QvW8AmCp/q7F59yS8QTVovWQExrWiROsfZMqQr2JAfqkuxo8WNCasbmyLIyyxIyi0SV41LBHOGl
S6jH+5jbynU1N9BmDoyxwaETB5ZA7aAChCIsaRj26oGGCwq6+ALMwiziLHZklVHs58/hC4LciirC
JEiRjy6/F3oiRzcKilvIIi8AT+inmi85ajns0n5vWZFh2aET9S6oXiXG7ETPAiXmQHcstHjMjmK7
tbg6UUCV8qk8HrZJdkP2TqW9LEv2/xeECZJTEtWvHl58xYVnvxdowHiqHejqmIGplh6GaFzq1mnZ
DhCMjr4LidFttO5tDbww6MGQC9AyRX7kRRdp64zKnX6HZqoG/82J5X//LOnwTjirvQGjc/qUajhh
b5ojmZ7ZYlXVuZGrJEORMYSV4jivlVczpG9u09wDWtkBma8ZAaAOVjot0nfidYK+yOnjtJEcJQXI
HIbQUgt7ixFfJqLmKhMrU3NPKxw7FfXD7PruM0m+eTAAn0OtVuf0+M+BOBH7kWBPne+SnqcL2BuV
bl1pG8Se0Ckz5K0/aFx4Latu82JXqK4mLvqwzXPGOIVJGTIChq/x48kz4/zAAu6s2AniDvoaXZEK
/3dKlHFFxeo79F00ffJ9op/b1GiyFkwXamKvsHv507cdVHMpg1VB8c3C10htE8LNBeGIUg/ZFlBx
9yykru8JRh3kCtdl18oy38KgHfEV0Uf4ofHF382y/GLPKrG8yXN/NMBrBWOkaG+dADNRM52vi6JP
6nYVvfmIKmejaCZyEEeVTKJVRGzW+DwfQwxfgjCG4T9m/STbwA8kaglYdn/+K5Y7Hx6ouqhgXitu
jnwQa+fle5k3CaRSU1/HVRnhyqMvWvmS2lQcF17s/izRHP+Fx8kbV9R7Rcm95yJUUHBRrTaFRa8h
FxEZTKOL5AnwjsvFQ5DvkED7PqfpDxr2K15MlmeGwjk9n4dbDsO0tZ8YF92jK/GPh02iTBdSXYLI
zTnjtlL9j7wNPR527XMFy9ij6JPnMv/XGs+EIjJwr59IjYvwR8hiKa8ISjL1N9SsrgUa8wTWvXbI
MLBKP2r8rqV0rdyEptskBxU/Q3w+XsFw5nlZsZcKBwhiyMhSYKkIB10Q8k2T2bSoz+VGZyYHMEGI
+deytT5DnEFKFlaCGUtNxGRykTcFkZuuHb5j/VMT6pbB0/QID7XeU1UAackPZkwnGpz/44Kdcx93
aB33PzNKUlKGgAwC6DDq8Qtumc4eyBFghK/+b4AspK8Nh9FOaYFP868lUarF2JPw6W2ve2jYqxPk
yhQERTHYFfWPfYoSyhKfniYiVNZILQw+RoUlbOfQ4ifTMfbhoR2lyqXb2ex6fK0v3RCyzJRdHvhr
jypmhH03b7eDvDXHptlknLQWuEn/n5Sb/9JIt07d3evC/IuGWR4t7vu0pXc0ON1yOI9EXVjQXy6O
X3PtFoJf9AU2a4ZBVPty8nSXSgGFDmLmgIFHXzufJwB/XZHleg8NN5R+3JCZB8taz9novE05ZYgn
DQT6dsIBEtxvrUGsal6WfKi5mKGnXl3+jmo/DtUV9r2mI31tMrt9mlVo6/ZcrnEflQO+XXIOAiEe
wn0SEBF1awgGwPi78qzXEF/NYxb7RZ1mpoCvioUdDCKi4x0aqISpCGjB0xoozwKVEh5DbGHz48O/
88vdvfIOqPvLYFOZmR8u6m3lqUTcUFxg4TntaP1lGeSbbTFikBjiFsQq7T0EdOxhgGIBS/TU8R3z
Pc97RjI+TWGLEeOplkJDktcQxJPVt4lENHI1XX2NRRep4AdeNzp9SRzvX38CWGOJmNahKfKE3ijw
h/XZKLskWBlcEx5lH3Eyf0tdnmqy1tMvfif56nlpBBONfVBzq3pSfHSGaBoM/oK7KgumTDbqSkYK
s99WmvVsnnyIDYEfcJeOxM32OVUIpDoqptN0eosGDjkjHaHgDSS171QtDFpMH0SVfESpHFZnNbz/
R9E8GARSXuIK8RIQR6AGqP+knF3z/m7bA5MFhG6CsIeisck7f0M0FTNmuNSl5rY+6BjZPF+kJ2lf
ploLVjYXaWDZ23bP5UNvm6rTRsDNwE0cCuYZey1dIv4/CTMaIcRGU7vVHk1u8NhFE/jmlRiP+XEh
HHN42CBgtkK303ZjfaZLKED8mp0izGjeNEJXi77lcUF5tDvTXS6N5ZIZGNFdRQPUR1aEtFaJ9kUG
FC5GAmlwKFMzMjPQgZiwUoBVwLGghuNM+r7XaO8nL8XTqpfLC4qZdbbXmkwGuP04hfx3w6+bHfVI
m2i0THUtBZ6i21nYQo7snT0B9mjUoC/iYIc+xZn2IUP8cuxpCJfa92QJ1uZipfw2n1PJ+SSdtCF8
ukHxW6jN0uG38FNsK8Ft9QHlE6wWqAfKkX9ufzrhFAnsJIBAJqNuKZ3NZN7YBMp/tybPvgtnJuFm
MNvGdMmBsbnujKgUGS/8d8rdnR5EMTNbVHkZMNUGW8mRQIyNuZ9++JZUHt1kLqL0mT4nTQhkp0wV
j5/DIbF1bst/4+6oBG82AHxv661grwjXyOwWjZadW5fqHpsY4ECLRhglNWm9T92cxvnEpQIHgjcx
abGar4B6MyHOBK5pqaDiPFYqmwrGumzESBjKaJFzFJPFep0BR+x4m6oaMkAkMOrdzd0vBQZaMel5
zS+Xgxdh3rhO6aaYm2xWfz6jT8q9r/xxSDlQw6tZDo3Dz/qodAhO0vYfjnlVyJcmQmvRbGbl6URb
fcI+uIr2C00sb7/6Nknfg15HaNU1prohHT2x0ks83ECnnDV185apiOwnL9EUqbBe35p2hw1llTUk
cF20laeJqszzpYzxBJiZ6RvbbfyanvNAJoL2PPtG8QQ0JAdzqrIGH+GBDu0q/An+sTVcnvjblH1F
lpojfliaat7icmVE1cSW8jSfIqbPDJq2rqTYnlLluLHH3vs7b5o4A/hUtv1bpJR7sOZi5kgtBZLZ
kuqePaIIpB0bTeWCZiLV2xujET9JBvyueRolgt7pi4Hc+x3qbAsT1swqcdq/EKv8hfEqPnaHIEOR
PQTi+aKYKpveRyQ6O8nKIdYr0blVlSpfprrfCqioHxnBNlk4rL4p+e6EfLAXtCnfkAPwy9BgQHUP
6Ukaph0g5ps2w0ERYgsuEVloFLBWZgJYr2dupzhH5RnsCgwIoLAKZkwq+A6cKMaXX/T4mhU++FCn
0svIoZECZxXgy5YNXsAM/eRYvtprSSfocsENREh0OTHpfGa1ciLg8akyyATsQtdk1K/dHFblwUsX
SBDwplhbFRB75zNIgD61blFPMtTubSohtpqvm/g/GY8NJqS/QFg3XQXRQkMKIxlQxWpglWpYxX+m
DKFSczx5sf16XG3y7zh6e9NKZvso73OTYTdhbaluHEm7654vY68jWnk3FXD8dC0TgAQtgqU+Ye/S
ouXxLgjBFV/1X89wqA2P+itJc0U7fj39vVn1abYPC5UXymmrp45kaasOTrbmlN2PiH0F9Lp/IbSe
Q0OBGwPR2qCeCqMJgpKiaNR8lg8/Golf96ScqTo6HLHtIpG8VZHnWKW4+//0BPg5uRqemXlPaYPb
RYiJPR2GGAdfwVPCsVPlJpuHTetr1s8kmAJ8m0BPKw/FIKEoSeMHIevXIRxQRA2NeBkIyu8XCf6v
NPOsmssoFkrXOah0pmOVeMQbv+gmuWYurg76zRcoGvTbKZ6ThmMXZb+7IHUc4LQslliSQIifSs2p
Zo9yTVglCV4zm79B5ptWZyGT76S3XOWFbuZhhrGi90EASLKZ6HgBa4WeT81qeRcr7AtH/174vPPi
qETs+Cpl1IAZFrHPWH5IDsXKkXrmoiNZZzSyE6B+xc6qjvcI9ZLmMoMvPSe9ZB3koGoJW432n3Kb
49p7EAz3gSS2Hn4XBSNu7BNYArbNN8XVzj+1QHz3TGgyszAgBX99p1r0edWb8CJYbkCbE9PuqTWC
WG7yhrAiUZgNPvXKx1FetV+rTd5aS2p7vQREQPKBUaveYZSaBJys74/mKG/mQ+no9iAJOVGpf7x/
EYCtrLZoU7ps1O5tt5g1XoD0DK5/WsDiXE02HzB460ZQ1GVOO63wwpV+kw8qV4/frr8cwE/oRyNq
8jT5l7Qq2W7x7flyP9h+3ni/0/jezkDtVmtyFnVnsumP+0TQD9NUBgLcrvX75zQb0zBVeIW89MXY
tEj8SteAq2DdZiDGMXMeMOmnleCB4t1lC80jmnMn5nDkt4ne5voexr3/9l0HzA4QhmfJiYf+2Cr4
vzVttMfG6SxrsIqxwE5Xc0qnUtPd68bW8f5auSAymy/cGIEMI6y2q1lByrksNONIPD25OxF8ou+u
iQZYqW+FsovCZl9y+UH1r4oL/C9/fieP6zA1JbG4k8iF9zLxLQlqSlEIiUwlriGmGsxtVcu7OfjN
HQDURE0MzqX/V6ugIWZPxlS7CseZB0KMCxrDoWjc7uTXMyv8PVnQ1H0rHBcu/RdddvH04TzEmeRK
mzwlpA9sB2EZVdVpx1MhZuWpkd74Ngr84jhQQ8XA3V0IMY3pFXUqzSZVu1+IrsI+mAMtA25jY/r0
Z4Y1+8nIPBW4K1RRJiHcACVgJGVU4dJ9dClaVRAzBOdDsvw1QEPb8BJujWdzi4Ua+tkS5lu0s5By
1h4EHoIhbDFYhajxlSZOoxTGDLA8Lz0AhDffg4N65Rir8GHmtE3+hgvChN5sM2X090/7AmL2YH6u
Q7Bk6J61XOYPy+Rt2y95mdY/AgXA2qs3MpoPvp4bHosXmI3Ukr5Ppa7SsIc+P9x38HEJ1wRqdPj3
GJPb6+AT98cF7wwcIwhjWPBtOdBZYS8KztbFA452hLdI5QrTJHpHf9f3hJ+Kjp5m5YD3g0VznQfA
RE9wZr8sKM9ubEd27LNHKYel5wL+ycZKvEdL/KFw8f4pSNHmsYqYaeg7BrdqvQ1/FQ2fs+pkoe16
ufsUc64RkV/eQ6+8Jwm1na0dNOo8jXyuBswLMgj6+UnRM8QzSjWKu8QHSwaAloYjh8PRSDf0C4Yu
cQuHNnwP0SiFH7/XgJPz+g34ehm5QrBHYQPUMWU1+6V5HG078oh7UkbZvQs/GL4I48UZ1eQtUTdw
toAlUGXgBpBKWy/YDn632fxqMlfsO6GxWEdg4a2HCD9Oud8NdRDRoKyLBCFXKxVa2YRWVQM6ncQz
r/REDU5xfqJeLiFwhVDWuH+gRVH80ydfR7YVvgzpwPpAcapDI4ajHorMRjGolfVo8yrO2jhEtSBb
l2Y+cIucftitUfjOINGJ2XX+6RuFmDYPLZJKnOarIugInfNPAK4VgEz+QUAOPEmJrZF8OgiIri3c
1UM20Su/mjTLQv1OMgPDvBJ5rMUB0shluQVcp8k5iicf5WStdpSF847xYKvYiBgA6XL7+SZBz3/z
ZxeA0GdPnV3OA0G/OQokeLJNd57Rksz2LBnn/Qzi6umiOvFCfe3iimO7k/9vy+nwEBAcgM+FAy04
fDbJtz+bvJX5tOi6YxI3nkA8coV/gra6l2RNA0df4jsq7mXvzLh2/F9xYEfS1zqXNB1QFfF//O7K
5tRmuYh3mf4vfwX9Mcym4ohdfs8shP6zlc5dMjzu2uWGuEhdmjDrTV8tNagCNXwbobtB1qp5S3Pe
Tm9biXMhnEe/67umScb5BmdNDZ/yeE65Q2CDYULu0bg2Clp5Uq5rWuzYOZoVQJHe0UVur6zVQqFC
uCF2HYD75vFD3HnxzI0PXQkaqeWv1JCRuoAcLvtH/vbSPRbGN2+CPqHG+z7/t3Ehd1PGhyQVEtWV
Hieoo94yvWIYJCHY5640wJSeQywRoQtQ3C5SdQAX02AaU4rNHcR68dXe+2WMyJLlUnIrAgvbXDh0
XlIuFEpvoEG96i7LQBT7j7QD2/ZLs3aWk8pfdFQfWIAYwfT3xXKs6gpOW2R+MH8vaTOvL5RusYZx
3dKCPli2xQjr4Tz7Qm6U6poY2ii3TWo8if3HSTpLvYXv+xl1IFqa7fE3GAkLUo+qVvx+gzcrPG1Z
PTBKXnfo9lKHq4cywsQ6mpyOvAQkaoHhuIQGyxRrGlLFPZyImgERkHRgBwP8tqR8aAaNxZShPeUx
K8T63lxeVtiPdtgkjUWzO5w9KTp7LZIK98ZI0kBnTOaiCuLitxMaxy5wSa7gDWDPKXLhXmcPY4bj
oritbRnIK8+EY1sdQW6QcVbXaT3XoXnhmm4Ho7fusxAeR3AkjpnifwSK2WhIwtfCvej+02e6Ih75
2p2GzYH8XDhGymLjqU9FUzAlPw8O4A7CO6FQuM/CDT2D13zZDUOBMMQ7i8KPQ7gZPl2KR2Joh2zu
2EfrClXTHL6z6Mtu+ICVDb19jFlTARCf659y/SI/1hwvwI/vkNPzVlqqa1t7yBlBtmJJ4BKyJ2H5
ObDsSz1zPwi8BONDOHeYVNy8NUEvOTQEiIyR41P6LmWVMkrc94Lpg0jTtxpx4TFjzFDBxYO7mdCf
MP+y/3ExCaGATNApWscSqEhWaTx4GmqmRDmNDMHelUlOrl26sqeckfVH1+gbGDzEaRPzjK9l4rlq
0cVghYTvvNaKC08jcHvMXR7TEq5ltOcb3NFA6hE+ZmzyGHXD6bnXl5rwA85mHUzJV08L7cLJnwa3
lmwZlpOGALZNA4Dpl/2b4xSC0oApN13Ge22EjNQD8WU1Bf1s8mZFGodKlIK7KM7wEl6i7zEtx26C
BgpbLRVVHKkI+5BoZHq6+dItwhxG7VfzHip/s4ixIS91mGIrMPvVCg5NRNDi26/X3va/FWtBnej9
+ho+iHmjK7oGTfrzVcMNmbGhwpAXg5crZFmlkrN6tUA3CIKvFB15Hu9lfJ2vRN1rkzMTWHEm4ue7
aMGIMyV7fNoEwIjpXQyGQqcS6fF7EpYfYdymGN+g0hs0ChS9fsHdVni2Ipe0kRxJNeHZ05k/n3eR
s92Z9ue6MJZAKu9TWKR1fWp/WSLoLwmQuyuu6fZo5fPCGIRjGZgsbx9hLG4gbXTHzETRf81fThdd
iK1NZSp8eKuFVTkZe2vY3c6DyPPIiLSpusGTaaj5m82tt/ogDoxHS7ppWC61jGpm/xSVJmHMhXJm
4X5QRKdUjpANRiNoYPKblFVdQ7W9gsWrUVCV1tBmQwaCknLB9/hneVWciWzdAK0AG9Q2D6Mk6/IL
dpLEuqeglaUuvMsK9+SUNGhFxteMpVQ8HT/yXeBkdSdWlXNpZfUT0TBUvsoE0l0khIL1BN306ZBc
vsAWGUdfJ6Mnyg6VOYB+piKaAfzOUlmIw3By4MaEG9OX4BMfqUubHPah7tRt98f9vy0RKCf2FkpF
1AIhzVsX1LD+TcenXJQPvLLQ0H7ERBVvH2Jc34SQzkypuazRKZcemGYuUaU/WFxAVnxQTZRnxCXa
2ZAsKvlpuDojgDz/YoFFcMHDQENpp/U3gdBRXcBG5exvfLLMtLPbYB/TjDiKpePgqEbtPJ+tP7ov
53wyJzZLHI3C5G95uvK3aSCxKOhZ/Aou9foH9kmVOHU2FIYAtVhI/2/kY9U0D6MaICbVjxV+rDc9
ym6/mwrMzW00kjwXNLf9n83IkHDpMQglMBzXQfDyeARo8L8tXiJkZfWGOFGGyh9hxPiO4Y1lj57C
rcX9gD7KKo54edkj8XOW+WG5KgTFC1/c6S/trCBetbgAney7mlAQkQQOOfTacXdhiYLsGIqIXSX2
rBvOLgyaJ0z87bgzs6fnvM70QpMxt8dTyimwG2NuBm4L9U2OLdRCCbXCqZjIXrDxj/Hos9QgUE2j
XB/GKuRz+fvRLotq3tPPmi+WYbXLoLJfRQIBjDxureCTFxgR5Xc95CEJNBfnJybEcPalrG+UeyA+
8eTSdhqL0RDfjxk0gPT1ajIpqYLwWaR/W07plmfAqHnrWUE96xlYDChnw85asiUBMGCsckaqHd3a
zmVej40z07mQr0z0dKCLWxfS6VBT//5oZFj4G9Pgk8+O5OkIhlHm2GqDv0WjpBHMTEDtcbKeSa7n
OH4UOLUgHvTfO/ukDn+pz+rpwh9Tiwj/YH58jli6EgG6y7LpQWm5x2vKp2HVUM+GNp6PrM0BbYpy
CoWQ37Bl7gqVPcDry2dEitQCMQErReDqVd8V+7sTUKFtlK35dOP1aLZdi5ubpA+z/kD5lvljdgHM
VY+hVz5zDyGcfT1T6zWxdRLZuqKf7vRJFTEM/U00IjqXDwzMbZzITKMTCQj11JZO5LHFYn6tyxeu
Vlb2St/hsLhrwFB7SbJe5CVaVIudjG89TUiK72oEpel53Zssx3flErivAmchBASdUWxYP830p4Et
U3TBhI9lThkpBJP4l2ni/ff52hvQZuYkkWD24HLCPzPabA1XPaMAnNJTQjb0DylirFQ2ycXriQv1
Wp0wkOZ7U8zEpoMFegAlbZx/8vFa44nj2ow7TC/ThOHzgyA9LsawQzKOlPXXUbGu86Mk3KFjOuS3
0OkvePtxlDD983z8nZgazxVq345GpAe/G7P0GQAwxZPFh/xZ2b8LVko/3ylCFyPmzrj9qOR3uw5G
oItHqP377Rkbc20kNiOojl+AqvjiIaj38wKM7noXko0TDYW7C+vnVarDn73JFDvSWXlmPd1GTxFR
da4mAmFx73iD5SRWm8gxYzQRStkDoHyabwUzsCLzqZiJwL8pLKaXkCAVMYPeEmmnKFQq4n8nOlXD
9TSWmYOwQHfNF58jqwMqL5mtHULo7Mv8MYO5axRhLZEvdj5MHrUS/R9WPCyk+L8Fa+AsNsA9uvdj
26T7k8yOGfSK24uST8ZSZfTUtrpZR/4EpbBjkGuwB6zpSGOtewDHTeVVB+CIuY2ohdQABFS+OGsD
qVD8Cvlisd0o04dQB+rA4QBMIsfG7cI2MJZC/jsy7FeO7RaxDDC3ngZoRUC5jTGSAd/N10Lov5h6
tcF3u4i6MDiDngc3qGxFlg5K5smOXT8v1O84SuWrfH56PfWo5y+2Am4UNOh6vB7urSAXcopAPRGP
RP1PwcT17JETItv5G4JFDDPf6uepni5/VCHvN6md3tplXlZdMUtWPRQzai1DDK/S8TnDr43sx1iL
mt1ssZDhG7dXJ1sHs3F2H5zVqlC4nqNmA623DFiGmzWlhvCHrCZoz3ck7vJpLG2jBAmpYD+/CnmC
JQaOH+/j1UcRh+tpMZH54jMKnYv9+MQVoSaU/MbI7A68tQKS883oVil7sJgBpzyud68DPGKSc1LG
4iEjIPA8jRHQrrozbTJTUS+Gnq6wJo2w1cHL5ONdkc0tVuBK4yhT9uptm2c7vqrwzhsbP6RFzehQ
goVkNXXuancQcCb6iYJAtfX3c1md8BRowXbNaOKYjLVrEQpo58ZR2yCBqatAC/iuvr9F8TpT29a0
4emvu1NuJx++qICHiwv7EeCW+h2gvGR+qlPbZlap+lX1wKUaAgSh9qIOX0ZuRo8NmloIf1gYp+Zr
emgok8TyCePyViQKtVMLQfw0alWwtGKEEnev5i88NB2yLs7DFExuiBTKwykrQnhnn9eWeCeKMC3w
S778SsBpdCjev9cSjjhhqZR79Sm8gg6SPgyYB7wT/DNQRRRRTE2FPG0CRcRnSIn4nXmoCcusvCIo
+2lhVDubrNQ8nNwzZYv26lFgQGfV/wA/uHJJq3vccw4e2Rg4R3sfEOcKueIRdzTCuBcb6X/6jYsp
/KdKnYwE+tj/X4kLkLClCJqr/MU9VXFZ2V8J7rLs95dAZY9oji7TArFuHu5FMJt4RfGF0wEv8qw6
94neQ2MXSPYC157xdFzAiQwPuGh0i06bry1iXBt8se/P6NiKNbR3AqQ2FykF+KFQ1wymzlccCwuv
MNO9JHef+vog8+wPPcqwB7YDiTlu3ZdTlyad0g15zQN69LLhyMgNTEZC1fCPMc+IRUssliZ90cv1
XvkWMQ4cYNU+BDTkJLuj7A61qgkbomA1B1KG5SGqxqAdCanT3KqfsEgsi/NqLEF/Ah0Bop7Vr6il
vbApOZ8t3uM9C34LmlWq4UhV6pjndyTVvbUenDtSkuPHwL+B26GQpM0i063YHw0Lc2GdqEn80o4b
sKqWJEnzLzUygriKLweyrTMaX/dZZFOWOeygqxQd9g8IY7m2u3g991X+mGw7n4KLcG7bUERgdYQQ
kZjItGCXrz2idScBkbD3zKZKGJJj01Zd38MbiH/27HDZKFtJ8vkQlZ3AuTKDlM8YnzFl5P95+ZO/
FmCTc1p2slT19HIDfXAG98N/wfhhu1y7RHfRrm1n2C307wCsZPjiQ5GhwYNRpOx30kNAPrANX2CJ
Hk1iN+wt9SHFELTEFQlbkhohbet7/fMdOMle1KPjGDRCtA1dYZVKtbU7HQ1xO9LWkVWi4dpiqNiQ
N6oqQU2z1TyoLDN7Vcsf31FsxmM/DcfNG+o/ymIRJSo7gAensLuGq0khOxTVd4IIK8MHGRQiU8Qi
cIOuwMm6LXd/RwCa7kZPq8eiJmUeQhjUvFJQ3et25+EOrVYzSiBZ64PBoqf7GPCiMjd+ISddif5C
oX1MNswcngwIa7k6RsZ/oflNJQabp4fSwH1Ymmsvq/LszzZUagVrPRuSfZ618ywILTSBLxpaYiOe
TkbZW8Q+sCo0LI74DlF3MJVThyr3c3CjS/gQHS0U1mWffo05ikjk4y64nmN52cqKgFil0k/YciG2
GT17hQggsAetb4r0OfQBQcpEhzGT25XhdJ7hKZeDh/n9FSyA346Evai7jOuyEybZazQDhFvV2KN7
OwhXIO6Aanv5lMTc3au6zbqdw79hmja+dY6jDJtJAC3/nN+EYqaCrGCdM1uacSAo5PWxCJ3DMYwd
frquEPpdry+khKcE/2mQaVv304T8lBqIBLnfUuWL9YDiY7gMusYdAfSALEJz4vCKHNFawCi0k7u8
QBygllk+lyNiqXM8bxSCKO7Uf6ateAKVrxcGJS/o+Jsho/jlpPbSWz6pnGnItri8EY23e+ax9OZh
0x1a9qPqGJRKhfzBMEMX1ui0A741TzB6Op3EHVbql7WVMYiW0PbHulYL8d0a88/WORH85GrbhTg1
YVRrRfX8SHabc/vcUOv5s0tpbjol/LO722TIP3rJ1cFiH1HVqr0h7j2kjxCEAw0F1AfgyVkSOVQH
sDgi8DRJmtgOaq4YIV9KgoByf8q4i22jR36mRAYGAHfx7yahtK5SYt43LwTqnbdcVNEB4mmR81MN
QFJu44VDTNXRG3mhPELTP3a85gSCayHhoC374M7EQX9cxv+UMt3100u+Pj3yW7YXbgeyFQcRN+RX
EZiAv3qmyXpGc3lrqwpFEr/vQjjjdEQTaFw5WAOgQCvKmwzN36/mrKEoWi+/8ESxIrsbjWnxHMeW
jgL6ZQvDymHDRabrwQ3tbuSw4T/Vi4nWL2rpo+c2dh70CN3Lfo+QNpReGEcK/3d4amQGBm/AAJ5R
JtCg8KCQoXJue2KFdnAjHWtyxuSLHKHIy3h8yl5XuNXVOjyvmR4gHw99YNFuHpMGlwWRVShK3Qvc
Gu15TSQJzjy2Gw3fIAQ9UynZBuwnn+GF/kaAmzoAAt005UGv+mq+b8E/xKeV1EI3F+kjjTjEONUA
3QdXR+101NH9uIal43b3s/Q5sHKN3O/7J3vWleTH6qaUXT68wtBQE5L8Aek0Ughpq+Lq2pQfxh9Z
/fkh0Bz5SOmyNkyaDFcuM9L3EE5UWy6PHx6RARHZxBplMW7x04T7vFX+6fD6GBiW+1VohXPVk6Qy
tOV07+5ufJ1DUKSJV3l6B4auvZq8K85sSFGUy85G4Q3DD57odUtj2nD3oWOApND6nv16y8JzRkWb
gjgM4/mKyASKS+Yxu1k5d/45L7r8sdB6qRbKp8L1mCjpKtLjlutgloXpbvLuZ0MZK3IpeiiHlIJ1
+uzW6RDr2a3v3fWBSWFZg4G6EFXp5wQ8R554G36qBtHWCmQtDSf8+48Ug2YU6iQuSL8rkMiU6H4u
xQ1AeE7d2UFxbqvEaOM+UymAfNUE/Ro5ddKndpGaaVcJlF4czIEnxUFErLSflfclqAFB8++JOYZE
2QxIUFAO82/NI5mpY4aEVKN0lMDYSP+1S0xNiOn2IyKWmZFezvINihzykZw6Mv8/KlxjxTIqzXYP
pUWhMCh/oKpXEMZTJDTrziiq5xlrWx5M0qFAl26bF34Pg6x8nDjVxin8x+i0jek6qnq8djfVkdcU
/3MkQteXp7Zb3z4CvKmRHMF5ksqR2OG0Q2VXnJCeBlXi+YmLeA9sORlL+55yBBTgALrCdUiczcok
ig9x+RH65Q3Ox4AJR8L97a8RD41UcMyUSkOcOdtHR3Hoc8DD706i5SemWiAMUPpJvg4qMyLoNC0F
px0nwvb7XaNFmk7KT7klkJsTiMet9cPfvZ5kBoOYWxgozaKPW4jkR4zssKKT6rqgSdXpaBUCzFeb
CMl/t6WZPQjDNdexX7ccel+1oQk45KlrBr/uFj2deXJSzFnUw6gZOduC4zg0m+PquCag6vznXumC
FsFQt76GnzQacZQ+/EUNp+/sw/pcy8vUf+wByqYbY69YCMCVFlR+KGJfJ9LbdUPozTKdjeSh7DN4
dI84wdFqobqnGiKK8ChNAZpHJzaihOeTfNJuRxy8DcpfsGcxHhF/IGaJMLhaNf5YXA9/SVklc9+r
8H/bUgbRF7C8b3TYoj0tniBKpbzYkqDO2eR2Ei7f8Tizd59iRCQfbjeGsrRuB0mxPTXMcegApn3m
bz+1QI2R3OGSytSXfia5CnPSgHkX5UZ2aNtBWXlFw/fqRevyI0H8KsFlArfegstunhIBKU8DTOsW
zgs47Zw2Sio/Hweuokxxcj8f0hHINeoV6g357gnla7zODspI3kzepz0kEkhGOD4kyLhoTjUPOr4a
bQC9kV2IGPA2JeqfirVR3eM7dImJxafawOi4+RUCHyUgaQgbZm3JCkQ6wDpPJelm1i1DbBQTwkrS
Lk+1b7R5nQTPZ8CmBAUTjHDWgqBGhRAzjNwAhSr3WFCCfO+r794t8YpGJJ7JAzS8Saz47ApfcaEt
W2f1M9G5IAwp9jo7wyg5lQDdR7FihU2xl83l/nada075gKJ53bfPbOwu7sbyWKgtKuhYGyYACPda
ZaLgXDkcIfYQEJ+N27o8HbIwqOrl31n01A3SBK7C2C71HBOPlNbSwMqlO6X3FM6PT51/EJUa+0JI
UwXgpHGa/y32ufdvQ7tr1ty2zkAJ0aAMsKiTBcczy6HoS7RLMko1F2D4qX2OY6b6/ZPo3yw9reUA
UV915IeMUr5uRkEonj3a5L7i3TuR+iIM1gqg+iHd9uoxqhr9ohiJP1+ogeGK+q/A6ZCcqPMGHuwm
0EPks1+jcjuGM0gNsSLER2TqJduhOn909JH+89qhQZ4t/9sMy+7hMascmq0spqV95vF1gGe58LzJ
JblP1lLgXg0PIIEIonvGCRuq7wIoXxZD/xTsmZ1TsNN8/Ej4TiKHFs5MWmBmbP5v6yOrCc220juR
AKDw3WWZXzbTKbogMkbEA5PeSlMrCqlya4ISqM8A93+Ho8kmFJiOKPAvI6yNtaEybBLGXN+XLiGX
MrzRzWW5TSpn7ElgabdwdBw0RyXqTloeICMuNa6L0lKkqGUNgh500z6lZQddNoGKtxC0CltkJT1M
OeBnQJgNjYz+9rMaP5debV1ApkSsvgjjjfHueuR5YntsJfn19Z84rTITGH//juOw64UPtv9dUqvm
hLzuVUp601jAxyNC3R49coAmOrDh7CDjYntJGmnjG2fxfvWDSuEkfnxk5xNOGKdK8a+m3adorVjv
bu5+tcyKZ436ti/FvRwExVf488lcGPS4VdWz1lbFbfYejNSBUsHUckwJTsZjHYgzVYQ30+mInmUU
vOwyV2kb0GPGwvTcd9QujlwNKKpj75F3iUlB+XV+DL09V8fc+PyQD6g5w+4DL6IxvW7I23flHqU7
ZHu+2FV25uU8N81ZtceNnbcFxpvX9b3oCeWg79FdhqLW3X/ZxmjchHgRkpS1LtLmBO/FFkDX4W5K
OuhpxXpkD+vJbeRzBGv3qLpQOh93q3gsPUOTTxB+70PubySntuscR/8ajEyO327XyQ6184N+VM8T
Zlnsvbfr2Gj05qR7XZ8AoifAYl0laa/ITjdT17O/KLICgtSzOfxHzgho2uVU90WnLE7T9NVS1BH7
09fMc/+zne4tQfi2rYB9esOLtM6X827ztIxCdcy2gdeaCU5GOArTr7Qej4CqS6MjS80uzS3W5jc1
SsR8kOyOfl/KKupc9LDw+lvDWHS13hcEcgcVeSpA7qVv34I4uvsQAk0QHE+Tx8ew438QQNaxLfvz
gRtL02XKvPQBhfyOtNNQ5EXn6wpiW95ZbCg6hnz1Jn6FvK/tkNzoFNnymGOlnUc+RAMAjQ7ZIfAt
7vQH1XtQrQuZgzHVB8NrucD05boohgnl7RVNa8fITo0RC/J/uGFffsfrGTzUKZRq8DFX2uPp/Bnx
YgzRRKSLdo8FYF0z7wnnOXSrDQFa6vmW0RFidqZkh0lMN0jj1gCiNe9/3UxozVmiprbpnsBRJw0k
C2Fw8ZsxJRDB8Mn1edNpqHiZQPOhywyOOh4f5b2a0Oavt+ewN8EevYwJD7gJrfZAVRLEbDU3YT9m
R6J1vw+y0nUS+EhVLLRbwY9i6sUBhZj8byKCt3DHlVTeQAiG4IoXig6HRnSFv79zubHCuKU6CPHz
UbF9sfUy5qEtvoVlcRaa5fGlAfUCMQkUQFZPGbQtvw1DbryMDzSpxYVg013LhFLwU5XdHPkgeCys
UTUr71EJrBb1/23Q1mA2p5iNsH0CZwxq7O2uEM6veVv1SwsYIqMsIfDg/OZifLEF0BrtT7hUCCRn
carcjnHYSQQLGO8Qvi1E+3r8N0/KQICKLiwe/qNK1oB0gFAnRb6ENWX/Un67v5qaMfiWgme+US2d
j+i79fQqWY4cOU2IBr3oL2PG/8DESkmf2th9vAu5MCZByaPMxYfYQSbzKeaEPoK8jQKICcVwNLZx
sz4+1p+O3ENDi4fgG7pD9Le77QDwm4RS7lfbZmuTptl+x+CHpl/Hgsg+3Ss0kVVR78BdR5UHp5hv
V4nmHpWqlSiBcfEiJzrKQlGtOUG4VtXll4wW4F5Pzdg0lzvQXMN99Hn4djy2N9eneBu5YeNbQ6D2
MlxMZuHjJcsK6MU+hUYo7shktHv/Iy4skltaO1vmVZL2HMYDhHrVeH1YsMaDHSflIBGctY8t1/8b
n7SIPpWgD5t3IviB1okVY8o/zHYcAGMNvhFzv+8ZSeCWGuudtxwVZV1ezuyrsTX6Gh7+ybV4kIh3
ZmOywrruXpm/vQm8aqOJbYX2v1mlu078JdYUBs5OBGhjzx+B8IpoodvwtbYD0oqMi2pEI5vuwYvj
O7kHBlVhOdzfU9V6QYGaSUmEfN+Ctbfyx1fremQ3H/8hd+Z6zwbAjFABbcZyMIBmXxJaHeRgtGz8
oGwXlKs1PL2ypi/R6RHK7KSTFJYtV1ysQU3zcWmaju8865Df6CszlTIMniUx9ZIg6FjEUukgbTIu
bhAiQc9eCqBaJy6P27/KQ2PKh0pnIwc7CjjvylX8nn2lvPfz91bkrMScQi7y0Aihn0/BUiTuZeGR
6ZfXed7RTObBk1AOygpTS5iuq5cIqbY67XVdCgFjJrj/qdIEUpN3+aB7pubRXO8nHzKpVqNiwr4F
YPlKK8d0iRR/9h3UUY+bIjP+nCefaLsFxMaIoDhWU6Tat+To2uAh8El89K/rNIK1u1+nLyb7FHum
DS336A43sUC6wmdiU2lGLTrj8p7y5075ys1Kf3d1CBQYgfiZixt8uBtcRJ6ZYnslvgmlKq8/kF9J
om5BdofvtG71so2F7ltr8gDe0g8RkU7doQZEB/lQtyUt5EPBbiwgTjEsPbzMwomOy7RsQmphSfuC
3krOwFi1BBNO1FoZQGfxXk+tW4jE2FYUY47JsC0BgrZN33V9GO66rzOxZIBCfYqjYOuZKP6vYTTL
vT2iDEsLGp7ZvLl0tObE1Csfz9rVUmwsT0hmbz4yKDjiRFZ2O9JkiHgkhR3BJbiV00SQtn6oVhwP
IHRyBg2BJDXSbwfzi0B3818LQQPPoE2n2uicOaQ4tBIGIMj6rt/yjyjE9XYMoh3x3Ahq+IQtitYP
uZ31ujIAqXX69qseeXmYDRMtUcalPml7SDFCeeHLJHQzHtuVuCAtI4/uxgxrGPrVL7KpsGT9asqa
bsRR9yeHbsHPPZC62/O4NhhnxCHCr4Ul40GqL48WgZO7mvK201gbohnvXnyxOcbcN6XPIEws8gCd
0N/9y73tnPONHmLlV63NOjTPw6TO9ONLX+9jQNOiDiH01A2AfgJmXpNLtbv0HlkPvOIREmTEpqFb
RfOrn4e9/0NSdWw7k8HpocsLgsuCITIhbcqH2bzAjU7ECyqYiDLi2hN2haNbMtTuUD8KUS/bNCMm
l6AFfpeuqhkCIU99/GSByEG1sWHGrH9y5rWvK6y0d/Er9rOz9D38hNQoL2lC4ru9FAgnvSYpbLjK
mV6IOmwEODfg40WJCUe9+xePS67MQs692UCp1PCP+IJ5CgcQxyO/jGtNaAr4jeZCMGnL7kH72MUm
TDs+QxZSbg5TCKq/O7LE//GIa3SABxtk+QSh2mg0WwzLu02R5KcqjK6oK0Wr9qRQxKrDDDqgnBGF
TGSThMfVunC5oc29QN5IL7PfYpYhseNzSW+Wo31Wlboptep6gAZMgdxL8poeN5W0PxXeeurxJm6C
jZ/D/h5XdEnzWi5pOop5XpXbK3laS5SKXjZjkOBSbRWGE6YwcQvlQVc5bK8sliSH+XEReSPn4JXs
pGPWTRfJs+TxB6qdTMqOo7g9GYGPMQVl47dcomW7+ZcJ7G0Y83CxFAiogqE0k6WrYyoBL+pPzQpT
aHAgFiWA7mp99eqUkNSViMkAdYmu+cR7oxElL0tSkFdWerKBpJqvTrBSR5yyQTaT3qSETFeQateo
FWuqKdtPkJbzx/k0Q7TGDyCiZmysno+0RtCsd95K0Kv5emdQAlpZLv3oPlklsb0no1d/CXZEyLHt
7Yqq8ZXeGSRxIW1w6Ik2Zyz6vcez/rUZ4WKmzQCAxnbhCJ7A4Nf6fyl4cCTcMovVuy8EE5RcJNEt
OHRsOitJWJ3jOLIcdd0c6NVr64gNRe15HpMfUMp6CokUIKkKhGyUGs3LaXBuyBw3HFfVVNyMOoOu
WTn+/oX0dmuMq1FsMJc0eh6adQ4X70CNhHzrs20fYejD3jWFJFviA98iKG5kXYbjNiGt4cUKPYqt
miKtdK50pd5luFeFaXMk7WNXfPwt02PYC2ThKDm5w4qubwWD62P2UHnRtM7ZRTAp4S/UwzPgqPsg
4RHREP+T4YtDM19SpVGagrg4Ck1W+IuvxdRWwcdZQaVSRF13UsCzlHLoo+ZkySRdpFKqThLw9l0E
wh5fqfyJFkHdPWlqmSll5OYMSmQ3oeFaGMdBwcawsK/gCQ1a/J6g2fXeTGWcP5kuJ9Mjjd71BJkv
mZbO8/lLy+HuvnivNUMpvl9UX3xu1BjhYmPMLUL+7DdKRaWOO8mLaOXtpSBLVAK0psqdJ/68Epa6
GaER9IqUfxWBVOG3oAUYXGPOr8MifcWvo/gFJ0i0nfZNbLvabvp8x7gXEaMwpXSrcRSFW144rA28
H9QVbCKTc1DV7y77r3toKntHCWSwDa9nRD/d/Q+SqZXvabtLqpSqQk/JJVncRfFXAR95T6BTSMRK
+dYNU+ayUaWOVDeDrArEtNsnvKb9OJg0SZ/tSAWIBUAYI6CDxiogvBPgZLEcnFCNQBhaovdJpsTM
HdHbAF85CLcY9yhNSykcuxCkqNZcNAbtDRnEBLs5vvDMYUo6Il7Ej7ry2x5I41V9B9LEeCqK6t6g
yI4FHg+pqiz/tGOtV5kIdlhdI1CSGkUy86WsyJJn+XJHcfmmiBReKX2hQXsZR6aQTaBoGJWbbGrT
5UkMndUmNfGXHbZooDcBmf60o+ldgmSBcd8T3rW+9kaS/psxx3Dnb/XKlQpB64EdYPhIyG6eLZ3/
9R+D03TV27Dhw/+GKPGfPHK3S+0nzSTLcbK+zHmbyG9dvB3j1O3bTPXPR6Kbc1QWI674x0lRso6a
/2exg/0S0qpt1Np1ETBdpVW2LeIEa63t73truIZArsTHGCFOWzCtn6LtNjybdAto9jFl6DBVgYvk
rw+8nyRUWgZvN56QjvDKCarBtVmic0hm4T9/QkbVTPR6qGrC8LDrYmx4qIHv2psZm8O6heZ8bWuc
PV57Yop93S4WJ/ATADJss69pUcajPO7X7fQMQdWykKNFwLo1K53DoShN8soBriBg/hzct9FRSF2I
fUwdsoMKz5MgxrNTIE7gGsHmvl0yRIdrGPO6up/AqT3dzRUWvl+zV4wmS0EGyDAEXEdT0aPaGnW0
JmxWSIzn/GUcSEhYLxPK/S26hONv4P4FYrbWH6v8sDeKAzvqMUuVfr8jmBDLiTvjj+JN0vWuG8Ck
PXgXlulyMbXkR3Nw7cw2GndWlRwQc5YAbAue1+8YcYeP0C6HFIj+j8kQU37ZL4YEm3VoCqKzC/kL
aYjY7qYqqm9gMDUWhylc/DqrGYV+qjalZki6M1J/5Obe7LzqJF0sbkv6vzub2jlESRaCqjOB2MUz
3xNGsoHOmX6sdOFroqHh/iDXKwwVQfhH+aTuJPzdcut0pq2KuMWlzklD5jb1N0UHQrKkFGUgOq0i
dQrWLkXUuMIfGiQwmfMKxcahoGiwJiHjbE66MOu/DDehmXjWjgM9X8cM9UmzVyh/ZAZsT/kM+Ewl
n+c/Ajf47evwC5UyQoRtIEN6A2nxINKimHRmq/rrLPTfP51epzR6Sq9mGhjQVHI7tu/IXzB+hxY9
emx/3Yp5hIkplvOShsNFaD3VYrfwuMyE+E2Z/YcHnFaam5vAG1QV06OqSjVAOMFESwVqXNGWKdXl
uRwBPRT6erLx8QLJxkkEysn9p9jlR7HySe+sM7G9DFBy0AFvAVRELTjOeEo2jyZllVdYFAzDkAVN
ombhedJSB/SOV8IPTSyMUswz/BCvlGA+8apL/4WEPcAsgHB00fuowJ8dcuCTNnpvWl2r6rFEDSYE
UzpWdu2xn6/9SN8Vp1h8HvIOkq1vhIEvQMkMlTJK5Sdiuwr+U5c4CiURaTETiICeDBCLFeR+zEzq
HnidpNYDpeclHeb6oYtLo+WyhvCS2CFT6MSe6yYMXI5WmPusR2Rzvj67mcjvBtlK1+lAFlOE+8vc
mEU/l5iKtLZFg0taR6eDnMmUH01zTjrbIRKp0JX4VWUku61J7hkuQW6lOvHAdgNjygjYLRfD16iM
pivRyq+4CimNCBGvv4JS/Zcr21h7hUP9ZC6+t1ZanJ5g0BKmi1AwconZnpij4zEH6dvt0jR4P4Qw
h/3YsW3l+BmqsmRe8SOB6JZIZ3vPTws/3prVE4gHqEqP/r00xOBzlrDHN37xv6vNTjFglxFExuKE
vich8BB1nEZ35mFpTIoBut8XsbVJmIEAL+KFi8AJInAsmRShxdtyX7INzLyT9620iHYmiqrJ7Ij1
66f9ikkRmIOYUxYOmys+nI0fBpgnxF9spdO9g+jLDrnMLwC0tGcORALOIllZX0gILGqUmsud0xa9
uSUJfb1dfG7tFFOM8sRhAagGu9BgijJTbGVDX4o7B0JBcIyoESdY5DgMISSt/pyGVlgwgVJPWBFA
4nF1IklKJw6m1P8+Z41zM3Hsl3te8QXKWx048+Skms2PoosRjMUUZx7Dmx3iXWcT3SpcwavxKguw
HyBnghtGF3p8mHh+8GrxXu2R3c87bUi1ZHZaLNwEgbSCtbOuUyKRRbMWOa0nOzflb3dKAjeTM20I
aaKgURg4Y9rVLOr0l9T84Y0T/iYd3Usvq1pginI7/7YMmBpanegKlMj/K81iT1dnookzPVhcn3dO
Ow6KpvIBNVpl2z5cF4V91wBfMiRhjFQY33iPrZPzzIA4ZNZm4OgsXk5vOTScD2dDaIQqAu1o5Q6v
iczgs+Nq3D/MjH/lKvu+O8Kap+pUNdZW753lHroduXiC8hZL4wHrzYUI4m6lI7N1GA0whLswI417
QcQVCvyE/PIvJbwowy1F3i58zuodk9Kts0LFYAvl++6lquYMCxjfOFUi3fOx6jNJB0ORC1BEt4Mq
AZ068L6HnUZCz/IUr2iZz4KvspI/bxEPDVZGaLRKlEOeTM2Cjz1KOJA8s6hdbFtd0KZpodg8Vm6P
HQ7yONbyC4nrqduFHx2huIIJCt+deS9N/LKupl3nZN1PwL/lKJx/FGCqDYrrZbXQjX414ndAlw/9
r5Fbt4quVjDiOqKH7sxA+XCIcxh2M7mlIsQlm5scLgkqlIxNKVfB7HCqXP+1E0keEly6boersChD
EzZdYuc7yECX2ns+Oh7V8Hygz2yUe/pMdIM10JQNVYQtCSfAjPg73t6r6lMMwtHBtM4bRyAHqnbA
2D8kDPQzU4DAtI+5tC3hL+kuRqrx+3D8GbUhvIYoVsznYMzCaULMSd4FoOP2AwNkJISV1vugdwzv
8gJnbpgU+pqiS4o/W/R0XooNBschxpp5/e2wEdIozo/onf4f2ddYbgC6nBhkRNfpTN4ABZoeaoKr
ykF25PD/cAmRbL2WsDAWtNFDQLPfefYsJQZ0wQv4FIPKf1y1vdscjmOqX8IAfdBphG//2BsGLDaI
No+s1ncWLE6FwfEt3DBdu9Yw8VCzCzpanC+N7q2KvzWzChzbkh/qNbv/XjyiDL9k9tz9Uae1mUeS
H1FP/FLA12QmKllpzQ1TM1geJlbGDA/byjPqUTpTFiE/3dsHXOIjbtq5DyTKlho3lnAIGYmWbDc+
Hg0lqAyWCgBSRNXgo2IR6Akmp1bBU5GWWt07uOyASHp3r3nNeUE3u3MaDWwlJABUhDWiXWCh5+An
vNSbIq2UvKowWfBq6BBGr/rRbgJe/CCECLfWGqLwigwLTl7m0CWPM5c01Mm9CO5q7hJvIwB50Xlr
gBkNgyT6thwts35F7nm1eXBMrbb8ExJLoLvjIWOWnFgt7bnDtsrg4oktORmJWXWS8aNYn82qFj0r
Uo+T+DJfwTagrlzGm1dywpSyZXPVf5syGqe2a56+SDnIKWcCvhGHqMMp11v0qZ24Xw/mDssNCYU8
rZiLT+/ihSsdIkSjgfWReCp00UfPGSnXXd0Lqkf5QakZoPV6a7mfCmksHavx5nVP8sNQeecBtMtK
CR2LiYJ8mqDCP8sJA6Q6bGpAdwl923ciU3+JDn2oUGyXZKQR5qgCNyAYcv6kQoyTlFEo+f4NODMb
oC1ikDSt62pc7ti8sagryr2j1N5iiRYMluFOMBAzoX374vIVQDkesnpmRJWavABnDQIZTZYVKo2m
zV0aYUxKli7zUkEL9qd419dvuHm/Tbb0qiNAhOKhBKI+d7So9paLGdKOvfVr9uBWElcHnSahizNh
TDljQPxB/LPGazIw2yZe4fo+NnnG+PJCmSTFegCSJ0XotQPKQUBotsrQFUyzUnTHOKQg/qBGnEoR
BX3Bz+CZVdSda32nu3Y67RqhVcyO7foPdPSEZsFoZ/m2MftPqIbY8IHyBU6ztON9xikfIVe8LSHx
A+Ce6COmU6Km7yGP/dE0AjCvQBZDiQ0FuQMvgdRjsPIOuZ9oMvCZyyuDrOXUeX84V/FTbGsFj2Lq
IiYbNWnynU7KcXJfWFXIdW7ChX6xXwLc+3HK0uQHOCxRHynSya35vBUIHal+utrm4+yrnQ6m3OSj
8EvVoGRFev69iP8Lh0WwmsSGXA7YPBsCDgy2ZiLoORWOZTzrqctYew7wNeDwQImRD78H0QBaC6t2
qGLWSianqKsbGXqJ9wVQ1U4Obmj3y/GE9oI6zaDFVHFssiElauBJMNuZ9AWMU2JYKLEddYpNu1a/
59+ZV0VOPbdi6fcNl4L9Zqhu32TPJ4GYv1dFNfNd+9Gx3KOHxMe/fa+fggXH86fnSso5D9WdPp5y
Sz1YAxRO7NtlubJGdMbDQ8wxrYQ7mNr+pPCGTbhQNwlgtEkDHlLl9IiCwndsDrJ+7G0yE9nCilor
qZCodJIt59b8N+RDSe2MGEaV3E5ET8KPU6HeEfJ+FbMh0Q+gRLfS++LANSgKBV0gGEU3IqlE99lE
ux/bJtI4BBp7eVbOR4g1RynJYFexYbfUvAi6BCduTdM+odRQmKWKZBlpCxf+9PmOR2d+pNh0bSHd
vSucIePqy5Y/abvQ9YKIoMjJltERryExxIdsHgkJC7ovusFxUPL9ERwiqPONQcSlDYqSekqxlKzJ
n9xtsdsao0jWb1pVA8kLDJ9kkj7L2TOZnXlgEATtv1YH+iursWYx4vFll2xJZmz/iZ0ZgFV7K9lP
1tFB38u7HgZuSFOaFQ4z8P1T0OAbTDZ6aN1wcm3kMWV8ya8Cl1rhQl6/OKTdcuWcYW4baUrphg/m
ltWFF/bIWWclujmB81MRjfd1+P6H1w7zI1UJvGDrgDV7TOAo2It6FTjocDeZmbcMoErRr/8LidZO
JG3e427ih+0fn+XlD6e2NnTYyF5D/xTpE4065jSZsKRcUG34/1NNia5VdYnYVslnsZm0XU4Av9gj
RgOlDmiEAJncCpkgibL+0ogdrvIFA/+2lqMcMoz7eyCp2K+S0zYh1aWyDMMkYkfBs67ns3TKglgc
OHShFBDFu49gFArCsu/T9w+4ABE+bJvWm+4tOqMM5PxkCCjvlvT2liT6CxG9808c89jYefkGIPb/
Tj0yaH7259q4r96r2ftVTejVB6lKXqxJO3CUlCUVJFnzVA9pQtnRqmBdNPDLXX4BPCSTgHs8NO90
et42O5k04o/mUJKFSqRjxTtBeBSV7XHYv/EGf1V/3y7jBB2m/G/y+b4ZAyHXD8EGBMGv30otz3kE
K49xd/enwXSXyo30xTByDEqvshdw130vUNBTMdZYgKaHOEt0f+pkopoJHfaB7lJshvv5Qn/WfBKG
X+1T8N+SuBbH73esQsQ4EIwPQIIcsgSC1ZoNGjBuFS878eVwVoQBiO4E4leK6qDYi2jrso1uaLLW
N/3QEpD7bMSI1GheeSUtZIy2qYLaxwzdu9bbvDnwWYhNlDrkoWfuMuMchjG0E4H+C2RdnCEDaBnI
aW5f5PvBR1j2fph5bypsOtYXNHfnmdJi1pQoAxcIsGvptVvfzsixKK7HF0cXzgf7ihJlwLdJ/3Q1
ZLcHsIxOTVVh0hAVt/RfOrNOGxVsfpjXtAFP45c4pGlKnuW32fDUnnEdldcW4QsHkti7xYE+T83Y
Gjvp8ZHPkvip0sp4mY222r54jEqfYePqKCF/9YXRD0HtYworpRBO2HxRvyFM9A2MdNnpXa38h5x7
aQbY8KvjiaMCSVHTRCANCoSISv5H7B2mvpA8FWwiel/bjhs45qnEMxbBXhliIXryG/JNN8huyIXZ
gRJP5nIOoe9VluPshJP/3ec6T0bM5mGvCPM7Be49PJdxLTSceZ7lXMfr6LBK1VLZRorRuGLxqJuV
lomLqWBkMcG53JKqhdCKXThV48zNY3woQaerE3t0DDCBaX8ZgfN+sn2+QYmbQtVYQKOnYMTuE/Jy
5n5U/UpS6ErHrxGu+6SY1fyKrEMc9G2DTRVJnyrK6/8vmtYarQ51S9NIDvQu54M1bHiwZI7kaSeH
i3e1aKZORspvQpCd0tDkbHwNx/nk6PmCjL0uG3Dbmke123IeDZTNiPLeLVcHAkvkFxVxga8GcZ4R
RF0EeOhqKrsl+49UQCv2b3elgUw9lIU88NzcvkFr4iNubaQ4ZI43+uuggluPoFQvORyHFKKwGuL7
p+Ro5Y+3yM+Fwr3k2lJVPf0+2+uDazTKCxdGPM9fyR9yF8uT3fpCD1+hDkRJNKC8zngCoGFRsqXi
wUVrgF/En1tZo+MFyETEM3yTv5O+l7Pe/ezmLX/ShOnDpwWvUG+L+9KN2PLcYRMCL5xjpjhNj5Oy
jFa3geLuMKEKwGVXeRnM5Jsk+c+xlpQpdO7t8B32G6T2p199kNWZXJ3foBVRxOF5DR2PguencLzL
l7BYOI6CzS9erwruV6Ky4ndvfg9VKK4azwZpEdWMJNGbeewJCQfOV0buXgyEh5aMioh+pp8zzbJl
zo3xYL+K/na9Z9cBrg7TCVJ4Lrn2QhzxpXdaqEmE4+iO3hB8Tqr2M4njVWL8T7AFpT0GF374APlj
RLabP6H6r7fhJtPQ2psLNFf+ZqzJutOyx6D5pCi3ssrXxGygjUrv1SFwGpaD7EgMdHcuB5qrb3mP
DPVPpY79hEfYHnTxQbUxlhylmCniSW03KvHVu0y250fYBJssNSXbwObNhQ8CTQm6lH3rMYfx5a0y
TYdiOLTNu4Py5/HgzU5aGGR/WVHeBDBADA5wbfOX5QlYbmA/5YmIp7rr+/KVoeFryPJ2hge9Agu6
UqAv2ig+dqO2VvpyyDd6jEg4iSZYx4RnsJgndOFZLLMcgYc6hj/1uV/LEhifBc2/6JsPwzl/vG5K
F4/+PPZQGn1PJPVE/J9OMfvCz56GM76gI0za1FP4CQyc4osjI250GZoavW7mg7DiNvudYa1EO3o5
xlItHW+VRy3Bhr3TGUtw2N0A3jGOLxgb0Nm7jVmwd3M7g7JHyXQw/PVn0VvtmloSOdd6kHQkgMkv
hxwXM6B2xxm0fGTBFPVUGraCaT+Rfwgr37dOneZDOjPv6E9YECrgBhP2JbPi/GRuOr08/FFkEmqb
NHdErDpKS0c6qZvY3s/VTTj8/vJrYFFUdt7Rcc0q6oqFljPrK9EExethvvnyuRO5mBS/cg61/QYK
Jy0Rd5bp+tQO1eznfmkXdvtmyPfPH1ssGRyGstGAV2bkKXFeYRXUoxn37IGZkFprj3rkA3dpstXy
5Ao/zXZ5oaymAR7hZhyy5a0WFHE94ySeK/Y92A4NEIGN4zAkBLFwOvMzLI30E8K4aL6jyjMYDZdU
ih6GEW458gWQ4u3d+naoewQN81JSPY3hcZsRnJSPZxqc7T+M7K6dqlTbwEzebcgPvO6/D1+WW4e/
Wjiquow1hvjRc0f7qYg2HgB1BRI2xs9sLhveD3vwytuG0Irl8NZB+9pgfeiykNiIWibZz9+17PYg
S14ciw68LGfpOsuJl2G5arYX2tyzXSC0zfywnaVU2VYHP6UiS2BjqEVXrACXgk1eBunXMUp7EEX+
vcxkkqe/S78JY0O5Ys3LJmEZXB06xreHFlvLdLipAlBGRhmHFovFVbafRT0BcXEbcPkwG/0tk1nq
Arx0F1O28G8ZWUbgiV2fcAdx8Sr83DEoIaFqeiGEQirZteQ0dOLrodOcm6r8roB6ohOYtkA9OvLc
MqO8icVwULJxLvYRFq6aXRlkbJJ371QRXBI6yAhAKr1IpVz6KcRNNoQGyuYGo3jLZo9V4IU0UgBV
jV6i0DyUyKPyiy71cUrF/K/nSEf3AtXWgk8iLcm8cSCW1k6CZHoV03zvV1kty0UQGeoiSYZ7Ledz
0q3KQyI0ejtmjEzYS9oYbtS+zG3XcaugZA18JX7izJOj+XbSCNdqWMb+ce1/vh0W9Ia/eJkQLpeu
mw/SxhJdXFU2pf0h7Mb+ZyV7rd9nsQhS0p2c5aIShTGdrvLcqxVXbVtL9gq4hzdSIzpjxZv86FrO
7lfGt/r+nncBAQUuLW4T3Gyp8fnqGnPW8Tz/EUACYI1vJg84sA+73jjU/tDDgm9JH2XzwuISHi5w
uh3E2rr7f1fh8dXR4tjolTtWvuVb0GxneoAxUjhSzwl66a7njrefdgE1iwRbPoBMMYGHglo4mtNh
OWMsl/mrBgXOFBo0HTbyCfS1uD448Tk2stv0ivjcnuL2KGP7OFv9WK8Og7FrOFZ14sDXhklQmoIp
YNMyukux94JzelPqNL7yfEET2hNbYRtGkTHc48dWh2vNKWZTuIaO7vJMdjZfIpC1H2aPm6CbcjEy
Vqvt5/b8fBQM036s7SduiXRiAZlYVBukQKs04fwb5h71aF0nOuzIp8WyDzrR37wgW0hHX/zBBSXs
6KjGV4Os7jJqJEfSxY2gLJCiYq8iJwjFL2UV/HHffhHrpi0uhtr+8ify2u3tTrmlS74++xm9gA6d
SttQlgOWlehm9SQdC/XwljqHRtiJI3ugxhHurIlmjUShR6Morhmb+zEVgT8Ae796pRF+Mk6kDwmD
J6I4pSqgnO3ylMMPrNs1w1F0m1Su1tMlDxtyLm6TryO07Vh2SPFLfekUETWnQ7M/3f1uZF4c0k0Z
2T2AHEoeTYwhyZ55XMrpd3UdImHuNGhqiVaGXbNmbnHyhUTdPzFqPx26mJudkKi8FVJ5kjaXv0W1
UcW9XEH2D5wjLP+mEYz9w+WRwNx+c5gTDm2wxqAHSfOjTi7b4rObU+MzTUEUs0Ponn9P9YlQAj1J
bGRFp39xghlOlBwmsePMv2xFGb1GM2RuEDC1++aOlZJyHeb97sAwsfJLoOAEpIQrUHODJNMLbMTp
Z0kA6MfspiAbAuVODIii3D41OglncXZtd/dHps7jjP+8Dp1o1DFC/sQmG9XHHAJj+NuFA7TgqF+w
kDMdqaQFpao6gll1xeQw5UJ8T/6Rn5GrKXLQVpITiEZ431a0eYlttZc1THvp9PlnWfxO27NXHcFR
n+jH+OGe7dCAvLz8r8FLHMxAvCVo6rtAWKBXuC4evfaAZ+OBLi/9dfmoxU7vaOR/EZyQgCC5j5yM
15Qz+Kf3ICvp++QZouJUXkT9K4rCwblZUUuvBhrTWmnEWsxW1wAnEc0hg2j80/z5VmPREZwy1QWE
SsOtMGqcQtOqR3fAW6Iw/iatqp7xbFyINQMqsfJLRFwBHawzRhTzukBTvFj+zu5nJpq/C79fOg5q
dXIf3C/D7Nfkk1DaMownAoIryothdTs6B8sHiZplSF5EdwTciltrVM2N6f0z/9X+QkiZBNWKSrZ4
JMTFsInJDfLxCFrd9G1JGFgYiXCqF3Q3WjdFskfuWiGA8UMgArISguOlAe2ica/rmzReFB3ycQsY
BOotGoq1wy0/UCj7ucxM7Wu8z/aQJT29+JrsUtg6iyuNayHHBMOcV5lFosvgY5zxNyAgwLXovSgB
9k41WWvGe+ryYDa/C+zEgm2jQIs3p/AtACAlerPqh/rDejgyjCKQzfUgC+2h1ow/pkUCBt21uSMd
9oVU4oZnvE/HTyl5sQvVIS9ufcp9bQkuGdcWzSVeDJRu/fFWSOjMiwG8R5F7dz3JNYlEjdEuO0w2
XvBpaa5foj7whMsF1j4v3k3U2RrjpscZL73nY/YHFEWx1nIYp1/GsHtQ8FliqcHb/AJxa3sTag+5
RKrRH1iwOubSoVmlS8yeulTuaZp1KPoy7oNC/EPXeDptHcXiJCCI29fBbKAPwpn9gKF5tn96wwBS
07MHwfeQ+n5/K6K4tEltvjbbQqNG78HoVCFdP6xggD0H8Br6WdaBSwlVi4Eis8CwtJHfNzteFYpJ
vIcIbtxTsQdPBQtInhrVPxb0ql1aYZRDJ4N7PcFUtDesXjtoJusdnfW8Z9PRFIOyVqPxPVjLa9aw
kf9DfgY+5DNJmSnxn2ns7Dz4AMfM/G7S++UlhC1NTvElfhKc34n2MuLUaaYYpMrYgmF2UB23pB51
NA/b+Uf5naWy+XUuXMjjDJBCL3cjz2X0pd4E925DlxCCcgX/uUQs0QXLfbNn23wvEX77pBj1oLWm
6bkb0GZAjcxZOLqS5b9nK4i/1EsrzVbAdJvTYvtKBOwCZAR+uT8p7N940NEksCdNNFi2COSYK7I4
mebu0nsLy9KRaqrEle1/mFgJy6/a4wk/Iqkmq20rxPzMYwq7yO/wnhBx2D7+qeeygjns3hRzVHlY
CWdGTo1KsBzox06KPU7hZb0Lc06WaEE6vdrUNHIuTdZkSuCPo0F7Zk+H9jdcxLv/HuEtr/5NvEfg
Hv2Gwb4CsNrlWFJEEftfmTEKQ7kchXRQTI2fpSCmyUbHyfBdOr/pfrCsqyHPICXGgbykao+f50ak
niteY2fLMoA5z5T0YP2hQmQ4Eg0Oml0yrd3bWFS7MAs9wg/kdZIA2BJcQNGpHOx1GOs/k+5Y3wJQ
Vj1vPACSm9TmDJT2NOxY82IU7m+4WXsGqsA3BcaMvTBFjzHXm3ebcLOSwGScknLr15BDh2ein2Zn
yTktGyuw3HZTEXJL4ZESC2umDAFHzAeyO9QU7MXMzsJ2c8M/tHOoT2ymYhKrmCkPIwLwRwzkNtI5
wv17l9BRxgaOgCphmjRx3VAn08HqSpmV4qPRQo0E5yTxLYQkiIx9358o/xlOCyLTE6FRjKVzEG8B
l8XJvfRIxB1aTouV1DdQyqZafRWQwrxebDvpOmt22tADsjG/2zoRNZoEKnX/H2tKYRV6JkukE57i
UYBfWll4CVdedZz9qllB7ii/QBhLoj/keRiqgJitNY0bxHGTNADOfQpbLsAvgF0tLo1qNgvmEjzp
eg/sUZ/gA8avrAah+J5jj80dfbQzSKVe9b4Tc6xVFgcpW9DaGepd9RtqRa6wCn8zc3rKdEuGjX3j
s5jEBm9IZhxsPLHWF/PdFW2URpWi9VkwYNOFkQRkeSc08YgghN9fabQchK41LZNJ14u7juZVlVw2
IKl6BWAIOGkobn1MwRm6m1XJZwzuFuOZUGq5yhq/EdEQirGDNUuxYGdDEN4p+G3CEt5BwqccYFDp
Yh8Hh8i0uTVFBELyFlvPMXkl9c1vcJdSd51L0XolGe1XJx+Z8spUTes8BjMivhqrnwONpq2sV7yU
XCyI5FVxrMqogDvPKnYx5c/TzOzzxj7MuRaE81BSaDvtco6Ae2O4baeutlMf5hFi0Ml8dpABpZXi
nmyduwLKclf4jXgcemMvU3DsYTjbU7rmydeOSEJXUt59EaGlb8YZvfsL5fgVfGN8eWyoQQtE61Mi
XuR+j/3KSHt7/mtsbE5nnG20JbBzfAa0AVBgJn0FJr1b8KsGGdzuNtATlejQGXca6Wj/w39lH180
+gLzJI+0iy9CRs7OMg1xFwSjWU9mdctxwguleEpdDQzdh8MBlAClmwS67bssvQzrq7uJYvz7vLgU
pGyD6l5BxwKLcjzWKpDFgjvsGpeJo/9aRCl4NkZQhVXMjMywqf1SYDT2c402ek+S30+WzmZ18ETs
0d6+2iMPOYkgCoCq5xr/Zi00vZ1iEUqaSMBUDUCiJJb3N0wydZWXZzftqLzc1+dXN1tC/GL9hOwE
/dYVSjRYREKRWT6R2GuL8CEf4fADryTXks88SZk7G54tvgov3FjHHb4VruyVyfEIyoG+yBcy4CIh
+MMzcIoW2nsy1rauUw2N1msr3T+Qk44at1BIYltrzK5sPu2u66vcb+KAAQQv9e0x9GdyA+rn1qWW
B97pU4zUMq5lWogldRYDOLdkpwtAJQeJL/NqUCWs07f1Bd5trjj0HZztCG/7MVOx8CRWx2ckxCbd
PlrLa1meyehIOtxAvqyrKFHNiRzaBxfZHyWNLQLM1N7ddB4z8U2Gar4JnLWdbcJd7lF2vmIEV/4c
jJHUkP8PZwyBn7UJzfY76BWFSsRHB8wDfpF36BfhzHVTEEU2UNs6uXmJE1SikE0R75rv9BlIQHvs
Bbh+aKgAwTmzDA8S+4jnBEIAV96i8+XeJ607VJtXWtTEdioblT+Xbbtr63QnKNF7tladd4teMLQt
SdlI3EWYlui6e9syfMttHVwoSM0CkfnnMKSBwu9Buy2dZ/P0s5Gi1qhdbY48C489w7xUUBGamGOW
Llza4WXOqOTJTT8u1Nfql/1gGD3UFnCGdw9fNyj5jlpNi/3e8m8ejSI/L3hxVUe47CS0RqQEwyIg
AQt9wdgGmEXd5lFrzMlkL6R1KcHT0AAkM5Jhr8zq3WFbqts/a9vXPV6ZIy/S28U0kTUgLUsuikx9
MNzjfDJRq/QajDvnh1Qp+dMzvNsIHAXvJjLUbdUMYeV9YutqSR9D58MGBLjzdwLlvtXeEWitKDKK
onR4Dn1LNsoV9t/J6cQOGCRWll1xttjJKsNVMa67syIuTC+d772LrHgchIjuY1teVvra8meFbUdV
52l5uxyBQdGQbVCI3gPNwcREN3ugWo2APfXvssW36IPh1pyCybW7ra823Xxl2NOwhNOlFypu4DtU
wzFekoR0VOXxDKwCqOyh9kZAWpjsiXW4ZM5g7nzUogH0DCz1ls1qJpJVD4bSIKnMSkeVQ8opPdlA
i1ffm/j8gxZ3PT9VZTN10H0yq00AkvfYNimsYPiJ8rATWNV+aQ12y7VKmR3UdinenOxoOseCNpTi
K6r1EDVZt1QSOhOOWjt0Pajt9JD0boIsKMy5Lj8fxCgwIpB10Fz/p+AXAuarWXT6PstW/KtlyVA5
egR5qt/1kx2k5cAgnA3TOysS4OtUEfpDu/qJYkMMv1GmzqF/CwY9zvIa3qMbWpYnAESfNm0ZUjLh
Bud0bl21cwiY9vgkT/e1V7nDdyxgqJ5pySl6rNXC/RtTufmTH58iUHLKwfTI/NbLob1OjfbhQfdP
4J9hTsgPo6zpFNI0yvT8eAoEVL5vn67Ki0CkW4bp3Cuq2dGNpyqq/689Pj0cT+VkrS0XTXUaWGln
EZY3h5FZQpIX+OHDbtdNiUkN9+prwYnQNAcm8KZ8zRzOPkAhiE8DG433XpTh2S/c4Z2fvH9GqzSD
xkeY5PLCbhvkF/PSbzrLWpaVPmyUJB6K+vkoBv2f+vsZEzeX7qkys/lI5lsob37VkzaqsBBc4jyg
SiAXVGEwjSw9BES13BdnNc3qYYZyVvKq3/adqvVJ6k/DQn0GyFmK5JhVI74SGKGUHFpBg09tDhdc
GLRe3KyMx2VU9Ez9ktP+vz9VJeQtpxqn3YhQl9tgoCpT3892ogKSDAXASfQXeS+HcIfO8BueH7aO
Mt02GXPzHW3/Wq9k2+WQciZJbLmAaXMXkYV1QsfM7ZoYFq1CTLnpT9pECHKWHfiuq7UgrhH7+T76
HUO2sE1kIIdbBm0vvZJn3XDZKCgEMQ8JLoSyxI8TML8+Tj8MeHFSNE7CLWBlmax5Z+v774ByeJNf
J55eAN+wmGQsTgZmUXZ5qPwuDpdhmBDGHAqhrrg374Ju+m8PSHWWuE1CPi/xgFeVKgTEUXPhOW+b
5/ArIZI3bbw7f9tVqvtKX60oIAgUCu5+0EwnhwAghU9eHjYSj04WE5s8Eg/lKnBPMa2isGIm5Nsl
v1he66K8VTDualWMKDoLcbC095MDqNM8P8T9TJjW3ZaElLanpjDitgfWX9m4Uk8o81Rg9DuK0bVk
hZDwmCirb17IerHoWiwTtWR7QmGJwX/Vur659Qp1rxak6MTj3uoowMP7hw3NRtndrbq+u/oQxrtY
1Z97H7g95P8clJFuhOtQrfWSo6OBlD9hZ2CCb3EBZhyH87z05n1KKwZ8ED6bI8sidub/46CDqzaN
5ms+RGf9yXAWGaenpF+u1piksMmlaYLJI0PKSJxobkRyzsdRFxI5qiVkFn8kV32YNttVMLzZa9Eh
Q0rTt9uc8aAVEbgwZ+42cY/tsBHXQIedstjkW1YHoCTSHA4qe2nC9Jbs4wU9miSNEjSkzvfGQ840
DBP6fTU6A9jcl8cBzVB+kWozcBV+i8qrBRDy6TNNfslt4wXvVqbob/fZ3GeVbpWC/3FCHCCTiTWW
C6ixZ82EUSLh/OnP1eiCxvDhJc5AH/fTqpQKR+wXkilyRUGdBN+zTsXiZ+qu8Pa735SH6peG+n1f
X1pJqIQXZD95zUMV3Q89KfEnx5OA3kVmJxT4xT+5Za+ryIRB/2mxTiqCkuZY1dBpg/75TWupyzPm
6HFmXVI565oxUtRxjY4aAfD2V2iDwLZ0w3Pmw0a9UPx7uKAI/Km7NFI+NU8sQPgj6rndgfsIkllN
NkXOCEtvBRgXK5Ki0zRYbTZhJdr6Hk2GxrXSyOnK1xGTzOqFMzslkTc19qEFgQZkjuSn9UFYkwWN
Rngmz8pD006bf6y2pBnp2IKU7gwOh3M+U4u0Yff39kbiDMMn8BwZzY1gWg2jculhGDqumQKZ+P6Y
Atx+Emptos2nP/gnKrcnJuXwro5IUiG5yHu4rR6F3MsfEZ18Q9WSHdIyB6fvKMTdbkC91l4X6Dub
7bQe6i+8IG2jX+VIodBBaA3zRswY5vPAXlcFzfefX2xS6cMO2FSVSHIYkPGxowk1PfUfKlmkfMuJ
pf1X6/bXmyjp1DPjzTTptrOv8yD5chz0ilo67XIm1JUuZ21sqxgGGh/x7yCIkf7lJsGD9rb027wc
BPEVOecsGQL2mtNjAHf2LZ2M6woBd+W0QEhHvH8GRHtj+V1IJCQVkKPaNWR2kkbYM5pgLPhGiePi
W0DxusNSwGxm4XCi8hbD2QbDPKtMaCSdQcqJC4Nf9jKCGGlShhjBjKRgQ2aUlJtCqmzQkzIWVU1C
qOcpUCfxrf6Uv/r/N1VtRWOgWxFDlagRZb7QLvEWUpahoDNnmzkDyP6stQ4RAW9AvtJmVAn3hRqi
oMsxg8rLpSc1zoBRpYJ7G4Z0oubcqJM/hM2wh7E0ZPTd+qkzaFP6rP51hCsYz7iG7XjOw9RwCOI8
WrbzfDdLMAw2+IOOLK3rcGzDlf5Hihb/XrYKO/ecgbECZP91f4fLPY6T/IHzN5SCPulSEzpZk19o
5crfIpwnP26L0/4GdatKiYyc61bTbA67WlNFWZrgl7RF+dKozDfju6lahhNdB55V9BETV8J471P0
MWlIkdrhD6/0867OTlmqb2AI7v5N0KefUF6g/vuzfaMDj4iYQgZAIhbTXPktEFlXgX9gUomycm+T
tNLUHB0onFLUAeT2sGRXpv7AGoXADDQ6k+eu3qKvxOUyrKs5aBiAmwXC8pxMEMxPpP/3EzlBaYAd
AzuOcQqH0lB4VS4p99FtVKsKLS1CmQHwCeNx35El3tV9aWoqtDerhCFRznQV57UBcbtySA+TpJk0
Uz2OhKc2Q5BiljR2fI+cOAmReizCJ/Q0VooGu6R2Iu84mEdb0ffHPRwrNHsk3qWp8yhlGCNkpmAW
+WFZHySRhxKf0Y+56XMvGD3UVpoeENdhl0KLr9xZnRnt6MFGOe35GOZFzs3Fne1EATLztJm/+ngT
t5ClNqdx7RE2xJmFhRH05COHHdWCpU+UWJytbXErSpQ/lQBk57eiL3bqQlSOLABDwQzsxoGoZ47C
mDXewLd0BPMAEbM3IaGQcog1df1koCEJ6S1MxOfjICRLy3RVGdM/o8XUQujZo8StRUWOTO/925U+
CriXuFXvbJhNqpbq8F3nst2jQ4iZOtZahpc5s/PDRu7yEKH/TkTkphe/jlBwn9lxi8yBhB8iKs9C
Z2Dt7CR5Qtq/pe9npMRwB1lEwwGzg3MB4fqsCZDje8acGGbDu2G5CytIRr3414/qtL15GR+SpDZc
6REiCHGbBdmJ/TDfbvzVO+zlAp183Y9KUGURaqvML3ACwxHG7G1twr33xBYsX9Oo+iOZ0Nh4ldxm
0nMPKoV/D6wD0Jf98Z3DN9EsJkhXkSIT86nY2/lyg8B8/hojL8Ey2IQLlptyudi1JZTcHfr/M+VS
Sg9j4B9XJtnJ29rBi8jpKw2Lud24FYGHw4hr8IyepFeZC+stB07LPUOqe39hy2FFkrhdSjc0C/xb
tH/ns2sFPgr5p73mloiEFVJ4K19E/sP0XB6zD4u8o1Xymq5qvNMw6ld8aHqshPuL2OBLqvaO0eFE
1NRfT6cyYSNZiXUf25AXVDRcG8PAbU06vwHqR9Id0OaDn4VGkm9VrNExQTj/EThmo6HAUbRtYl1T
oxF8guJAKz8B+N8aHEZYfbPQY/UT1jcYBJwZSQLKFVDAMHkd7rKokx7CJxjPUsXbhVTs3jkvrLVf
wAdPaKSJ1czTiWvX0pNDsXj737NqDJq/1yQPEPkoqfbIPZ//OJpRQn0m58XhectlkXcnp0Qu9Oaj
d7e9bzm+SwYVVo1Qp+8OtNxLLKlH87k7R1el0nJcMEGyaDys4gZS+570VGWhsP2NZu9HNDMwVtof
Ta5Tzd3CqgNtfKmyAGJI1bB8+ntB4D5U1IMyHp+D79ecGMrl4kNYL3+UE1XCT4Le/k7OCymghK++
ggp4g1NdiwB9pXufNi7gXBLvqBv+yMgJl6Gyo0do3DiFWKZoI/1Zpq0hb4tklDsY0q2W756H+GJJ
S9VFkmBTjmkXgIgoORbv8WeaxL3UM0xcIgaCjmYHW0y8uuALj6t2zJmArggi4j3hbm2f40nvKA+B
7xpR9OMKrDTvbATDaxogxQ/NHZo6E7TR5saVa+hi7WPKJH6UUTPJXEWEtehiPDPoy4ggDtrvZBNp
eIpqC7ZVtePgzr+Ys6l8YBeTkPAjphLCHcix2heMGn3Fr5Kknzc8jFVsjXE1MdtPQOG/kXoNF+u+
RCorfO1W2oqVEV3nYiFJe5bxq9U5el6v3krxvXRtOggYJLhd2sueq+7PMTKlG5x/6+jLIFhje35D
S1QGyG2V2JFUn5WYHavMbKr3vjauhzn8x6qRW0uvqvQw6+CLo5cwOXCm7F/h7mGm/56TBlE3UeBl
SuWozo5imyHlpRVuuiodX0eeX8b2WMOz38hGRzibWfRUp9sBaB4OOJnko8P9vbeiNJJFxEUIUrGy
LfVWtzRf3R8Ve6bzWT6JE0xZTZ2h8d17xSjW8a3sqOZdxr3oWfKwmRJjtWhYzv/mIN6lM263lJp6
3lHM2+zKmVtNkfGd2VeHEzwrxn+xELIAV7s3Vsvdoi9/HSVH9j0RE9iSu4lssKUpt6KvkwhZJEiH
LY4bBrDbc8yZ/sP46+2zXfuG5TkxiTiXgaSiTDa4LuZXJEFCJSR252gElqTXOYzxpp9+mhdHC7u3
bvBoMx2cIyD9UHNVmowRgH1SOWAl++acixyoUEubUOP3UseulolcFgkVwK8e/+6k4nTQGyXeHl5h
iT9pwzN7jbNKJ8VRajDbLNJ875SnRt8e/hNx/j5IYht36eLDNJmN1AVzK3TVTK25nn3lD7CBPNck
GUS6KX7Z1csdPafo+JfBWrlDMANSH1eL45w9+gkUn/UKhkTmC7dRr/Zax7EvUTTXaNmBmFgLDJMD
jxdLj9CK3YVHWSHHeWmsEUX7FjZtt9hY90rv8VdY6X3tQmOAEYjm/3LLawPjtOv3/shTjI/pTSJo
51+WVwNc8UpVr1ANpYeMybA/WvVQGV2np6TQHIQg70RhPxvpFpqBHv64rt/kwECaRZaRHsA9jdQV
q74qn7yU4ejdAT7uh+WaQ6r1xo+qkxbwsNOAB3wOUztqrcyCOu01CgLeC/4T+XtJJjfwqKdPL7Fq
eOOL8vLd3ry158J04yqpHEn3iee65AEY0HXglHerVjpfQzpCm3k4aP7zffTsJXFIsZOCwzgA2Xo8
Jz7EbBE08+CKGqOk0R0pHc1y0s+o3NeMeiUiWuqln95vonRc4H8ESSUxCdpxqkrtY4pi/Vg+nwF3
FMtSYYyV872hQUlx79c7pbWCA4Iou3zQvh0catX0C7IDbktPwSRIDUTWZx9EtCGNPzS+Yb7pksfV
zB+X6KsGEnuw3UHNOPzNokGphbTC8zOd+dXGpdvUO46KebFQ6xypMwUVGIauc7NFINm+MtaksLma
2WZSU5JGBr4ft81AtmZhv22GaDT4qvmddvFqd609/w/EApJplULBqvfJnuBWeHuvGXwOF4GgXTDS
E8YOnD4pAblxPOAyBBH35mhq1vpqIndroFQobOv17TO5qgNg/oo5oKuiGQXyr8uAjW1JjofDVlie
npvd5r6LCDgt6/7NT099+dkirXWycKR4yShsLO4EqVTWlHVFQ6qE6Wlg+IkwWvhc3xJRiX9hJrXd
BP4vyvQULbnKMdUm8RA7iO+dBNWo174+mBpjLoMljZFSZpnPFDmFEA93tcgjY1ckENvFkkrnpACb
H6iwTy0Cusd9AhokC/RQiYbx81J2mB/7WIM67Si1u2gSawyzw3Km3nGACTnZMt6YBXgATZARKc8p
t2TwY3hMLCtCbn98AVx+KDCMjViWyNK1W0vwl4VcfR8UjFcZZwREFfL0NFixy0sTwKNgFmrKaOc1
9ngJ76S7vhHhlx+W41khgnz9kYOhBmLK/s5HePlZyyFPXn2QvStCTojKVx19y90taMXWLGx4ZuH7
BlHXMSH7KWbKhDGJJ2hdMDjqVQcXSaDmFcvqD9ni2a/D3qc44PSagHkQqvo1amfhiJPpsorWnmWx
fuvb9L1UicEbwokjf7Tw5L+uqaYbOkiFpGWl/J/jE2+nPwsl0QDEud1K6eQlljE3HmrL0YY/pKaP
SMNero8NldVphzq8ozMz76mVwZgHuGxDLDLSUfBmEiIWweWuP5EL7Q/5+49s/ZtflkkgWKQ40O6M
3OQeO3tigUUYKzFkAPgtfAJWju+PThbaDEYzXn+tLulO+iFCgTtbsHzScSavJnQExSdpCiKhFu2E
WMa3gzzKyhYtMRGwiLzq4SM6RmQbBnu9arDvat8o1AJ4iUcPbe2cG3vZNi6ZZqdoCyYHZwXer3m5
k3RO3NUinOQ5G8wGWbmcPZYEtEzdipIvf1vLkhjsfFAMcUfPs3va0+RdHZLr6v8qYfRGL41VIOtg
yC/KMvW4F69Pgbprlas7vXsgaWSVLE/yMOx8aZM0KODC28SCWv8bUrkAO7kHEcWqCSBHaVonSvPP
clEpvb5o18z1XzrDETehrCw5l94NrkLpXf2qZCasWaRF+OhTMuUCf7HwH+yfF7EXWWAb8t80msbt
fsExrNtIAKBABSbn/GkwtjzkTPeMwZCLt1AFGubfx2CDC8h3I6UXdpp3gY8QDcaNFKRSYjbYdEOO
tqysm9aZy9gBZO/UJNdX5aqrylAonH3+oL9hTv1gwxniQzVdfsxTD/muM/KeYFDjDYTU7wh+O3Qg
7NLgMV3tFhs18bUtJaPyuQqr5CFTGAfjgZPmx6UHRlH3XqK45GyLo7Ydx1f1swmdZsHdBczpKZxg
JkzFuHSoj69LfoW5is4dATV7XfpL5fyz3t139klQQSBL+3CnFBG9hCqouoUCIBDu1ZGkjdUpWAQa
kQptmJHcrv21UjP9xvubpHtP6LtNHWBqhhRs6YSP6+ZRpy1uPi7kQqbF9yaYV6hQjzvACF4kyBo3
gaSCanyvImxyz3xGECk3ApAJO/gkmL8p3bRFCRJ3AkcjD9ekF7X8R0STipsgSIE7wxxBCSyxvFsX
NUa7heO0TZ3+yQ9SL+fLtg4TveR595oIHyCnd1erxMH0GNCFnXPTLEYPSd0IaZfzEmYO1fJb/mAm
RJUC3nSJZ6safdWXKoIeYmFfUKgWYxplRfCZc0TacDrMuhVdsNGGX1QF5vt3EO5Jx5A3tOfIqUwz
SPZtmn3fM4NUwY2L2Vx9QiU6rOViyKAXhjSR0ioQpLwqCKcLziD+leWnNokM/m9vvRs4hFhaO8+g
3mQExP0Ho3MUcDO8LEwXITHrK90B77geK8QOxR5+sbKiPz4N4iBZEEcra5kwrz99pebRgChfTE3K
lZjN3J7umvvctMQhMpzX/lCJrcruXMkCrFnLp6TonWNLNSFDn4ADNv1B53OxMg/Zg7bZyLCDutaZ
b9d1s4z1K89db8vnoIGORVc2i9Qi8BQ8Y7VSxEZ6NTEBil67kUC2d0B0btDN5mXpBhnQjltjCh+p
rhrT894MDC1JsJA9Wm+iLwGh0qTi+1zTuzPN9ilVpyL80LEGwKVLFb8IBL4m0epG/ujSzyqyugGc
CAB063PJ5/FXl687hl4/yuELRVUdps1F2UxDXfoRxfqPR8l08lt2BY09mviBr3fRqBFwuyzhvhR4
b1Wy8N6emUSWps6RgSOw3Y20OMDdxIsL8I5vjOBGrjxioiTs4db1CFARe95s7TbVACIslUhpztWf
jQH8UYNn1Z0s6iRTETodxQ+qjiC1YAlaMDl1Sh50nueBxgqvu5Y/fL+OkXa99CLJDzD39uQagts6
nmufoTGboGZKvtyH8p/1cUHi3CRxtYDFBEr8lGG9Hpr1Qdf9MQYU+L2a6cPiA3932idE6O6lEpUl
jcG22LlmY6xUOZsqxpUlyMqZb6ztOXNrhZ7CfQQczGh6mwRFI9sT088MkZBRj4Zf0l9b6O59ouHu
i1JFbuRi8D+CIdh38rppdO6m0uw5lrXBmhGLUggZGrSMUv4ZnlqSlEJDkrCDdlg0FAC3WFBPs/4s
kYwtYemPs+TZnJsAqEMK5GnWbaa8dLzt7ksyzVAT0sJ6lUXFE9Jh/tmYq3k9L+oRHC7TqAWBG2iy
TFqF/rFDCK3Ijk8MffNdBUkS90TFmrFzonI5Bviorn+Ut7MhgcX9yG2066MdWTwbv77ZYyK8liwY
FtRtRMlvbnphOgiccXU8i7d7DK6nKc9PTSpYf5ZzhGkFkdo/dxIXTIIdJva1K7jmrYlLMF2mXM+D
ortId/0B5QyhaMdzQEFrU6qCbtyjpk8U4JURa1kjVAb0JnolHCzRsc/WYVRaFTvW8Kn4/NK0M+AO
aBp5UhuDkGeguXJd8aLhX6cUU99Cd/Pr03A9+EouClJC362fnI0TRljI61NZzzNf9DyWKcYOeTp7
4lRIqtT4SD/bkPnNyzd9dQ+pHWIwYodZ1K978msj9eRx+BdwKulhhJV+Kd4unCw8gsUBcMtXYCw3
yItoABtV4vi2DuOwWiZNaH+Xr8n3XpAmOuWK2gvOtR1YWwUyR50fFyuScnoqvAVERP83FiV2eT/A
9EDHxJz8jr6vFzUVlO0l9fICrdL1XwJqX18/IpFSR/SX4MWs+o1p8aRYFt/m8cUvGZuqBZsI3DIt
vkk1vCR/JVemso51K4rpwyKN9dwE4UtIYTR6viwlsZ6Svh4ahb1/yzLihL/LVCEnHsPSB1vw1lyY
kIP5NcTytyv/8o2ClyOatrUe8Pewfq/hXZyuiFYZQxNqaqn4G4EmG9xjAu0nMDjEr+GrXyFhS18+
apZq48F17uFSX0HGP4HpzKcrzu2S2X7Rlm9NcxHYxK+VWATJoEqKfvHv4sis6IURAg/8+Ntf2biH
snCyWFu20XVuNOqEGYzXa27419BfEhuy8WiPLwHhGGRAlkXxZghAazu2odR97qI32gIw7Z3jqYlK
oph/wdyMLKcyEVaFbZaTCuhefNbdLmQeAQDFVTHGeMLVKK0mNIv7jYKTmKYfclojLIeQX2lLDtpL
uWRxaEQrRoMnEZbPXO8O2HfYYjKhBJWq0rVkJnGOUSmiGWsRBS9z4wkx4fg1t4NBsx/Si90KwuIA
wc+5O/IJEby7Q23lqx1R5cASUP9QgC2KBHzLbdQuta6+4EgxXJYnxfBsaDmtiKR5aWjiFw5gu9lI
rCaPKJedf3b4PsCFNm2R8KbFTGt3kZHS1xv8pOCBZU6gDWAwTVSXrQwtXxvbLBFXoDW8A1ODrhF5
N+KkEk1f4n3XztRMGHz1DkBWX0v1l1sTnOUId/337U6rmKkK+i09SHYgmSxnWKoP+g1S0g80UObc
kAxjMZijPyKn6CfBw2olQlUkSnqaD7ZET9mvixmDzeOY7px6zGTbd17G4UN/n7Qob76pG3LWSi4T
fQ0BLZZeg5+oenOkIHgy0eda/me+/JmcN7cWxXvBIvEb334URhrd+vZ8kFu0oIrbFmnsWHfpOLKr
So0/7ALUIf8SpvDHEhYF4JcF7dxVfcoB6ry0lSy9Ad57r+6cZmbVc3eyyGnj+4gL+v/4rZZWBXQW
TeZlGMv7Ilo9DFzn5fBkgbYFvh03kJjxamjCNvmLGiqfQVEiaiYT4lLzZIqizamIBJ5Y5EJlfgMn
i0lrfx1WucD29srwVN6B4lTaajY7euspq2VuMURQ79D/4TaXzX/sWVopoI/s7sMyNLmnlwy6LKfA
X1hj1Ly6KSHrtP47tWYF7WC9IlFQJEFPUsOcAch4x+fCKpp6kIWiRRfbRjEK7VTQTvxWPstzBGjq
0Aj67vxGy0dmkz0xGDncZX9+qkQDB4JJ3XNVZl4nrYKuQnjN/8UjTm0XQMC7foR+NURs21vTyvxq
B0tuoCBlobWu2Mutle8ju5Ax/tpK2i0EDhxrln1NjpboXNLdZOLGCCqnHCkN9tDyup0PoohBO9FG
WnHy7ER9P75EPGvNLAmedMuX4yY8OZELlpCrCzXt6VYEpinaGuW+3qooqa67FpzR2N46q2kHH1RG
WioALy6tcyGhZE2r6CJ2FuL43V62coZrP5MS5OGbDvR1eDfNZOd/cX9teuyMqcYhaKUkUaJAS7bF
K5M07LT/xzo5AyAFUIHe935cgm3/AYmYoomYz1MhmpkX5aiBQZEOooTD0rwEQZIGbgjbXRXbObGu
mERQ7oEbMRDcWFVFKyocafTCsgkl7N6OXqAkFfEI8cYHOD9ugcyolnJJnGcNizuD/RoFZVm5WQOf
XYi0VEnLXIRAm3i6vkiSWXR+zk/alXfT5IHvcbFlmWcCBUIvZlQbLLZ9NVq2opmab16vkk2PUWIQ
7iqbItLgc+X2M2350esr8OFim9G1AxvmLlgmYzIqZFMowVmG0QpyevWiaL5hh848KnI9cNJzgklz
+rcErU5jz3nRYWSL98BnVIijVWmXvJ0nG2LZNPtO6ApipkvOrsIAelHOuOUfrFfEhc0FmbyKl2tb
ck9jlUvrK7HeG/grc8wNeMPsPPN7mEFl7vEWu7JYHuXa2+dwSASvO/m4EPgezZp0mI49DK5im+sg
nwOrRY6XC4+AOSJMpm8an/7niESJeQy66I/iDAj0ptNnR8iIsIEKZ19Vplt9I4t/dtbPwLD7hPO6
vZQK5l3aQt2iaqAsuEoEjZJkqx5PHYWR9GOIQkkWXx5msZT4Rc71+R1o8588b6axGU2aq8g1MBNU
13c9VWwe3A+K9cdzJRu92eGYJfj4mOWLL0SYPZfP4fsR6ET0xTWlavZxugoKuaI+2Zu6bG/krE3b
ltSkv+yo7azmWmAXACOpusnp5baVwGSybaW2V7Gc3Blm72I48ZuOTGRUcSaads4AbwU8lWpkbBQr
4qty6oVSfzZtjaI/a0a1rEt4y7TEs2vjUAvHeRBNzPaEt70Mc9n5V8mRk6rHzh1GYSLd4xcJ4UeO
Jj1Q1uSgKAqJI1ng4VwQIehFUHpESPzQnxjkmKqB4Dtvdnk6kY3zvoR6SuJ5grb5D/2gUoxU1W/e
EV0AnPr5jVQvYRAUb23U2JSssV1Vei7VZTK5C4vmUG2Ta9JOe0CbOihlzEg8Lovsd+wOCdXx3JUu
4dOVNLLq82oe1R+V0jeSj8QIjk0TziiwovIkOhwXIdgaiKbce9Ae7RV8LMvr14BLovqPlVTEnEn9
Q0LYz4cBXn9+DEJJbdqiRJYkh4Uf018LnNOXe609Z5mO2WcD/oWiT6k3CpjnO97QBUX/i7YviG5U
gRso5/n3A1/AdZ4c6p2K2Zq+A78i618fiqH1cWbxRGKGmFq2B6pJ2Z/gOrrFRQXSLD0c36iwJIas
6UWWnZoAbu+kTYHWas5RG5tIR4lQXKX3yfkeCiQ7PoXc24zdcvOG3gPktTdE93tpLww6iI3uXrQM
Tq85RQzHR9vGYitcj6IJrohgMfV2VsMTijZk8Zon6Rqo79yFpl6hD8j/oVkaQsu2DQqF3TDiNypK
TeEA0xHk1AIPBJAdo4FVFx+hkPLjn7mFen0avBaJurSKHDHjWXpKDJcL9HIeC+wzq4EBkvNMlF7s
zRogUoyeiSZ18rxO0y6BwjVYOkbbzMhXQHkhgw5MG23fcv/mdOobzMMD7nohE+vCAitOgO29YoXl
EEHmH5qK9lXVdMr5+eETbsXHGOaG+GPVeIlV+nY0SoQfwPxdubOXwxoVDUbHMhJb+n5TJpz+h8v4
qUUYIheMrpfmfRvB4SJjdHmN1Y43O5/W1VRXL5CFYNuu0Jn6pJWFg7JvdecQ4rLUmfH501oyhmMe
8KBDdry7TBmPzbkL/6z6ZRDNk4w+Vyj8QNL/N/7B/jJ1CiFIwGlmw1hzUcmMI3iPUv+21RmPYmTj
DvXAD1f6kz1J+zRBbZ8+ikSHYXTsTDjWt0FuHhJf8jcF9l4hZi6dBKHsAd7PQVJF9btsKV3qJn40
1jNK6IXdZbkPQwFN9a74i1gU5CIAexoL1vI4xaK+bElaGBEuC8ULsOb/OvbSPIYrUFUZEpCaY/iI
1BSh/xsAJjLL5l1/+/IKWKqs3hQJyGYRuSoZNmaWHvqzHbgJvZX/iaexEZX2N7md2PraxLImFfV3
vfhVIevwkx2vLilnQ1E+2xL0zQVuUOjgBhnxKVl8oB8/tmSSlmbziD1D7ikvcic09Ew8CONdB6iS
DZeQZxFKY2CwQapXZvBEH1ExfqOCRNOW+L/OXqtduXxvVCLw62NkL55ZusWnCqIkeK1ULU0dY7cq
vBp3V47kVQvJLw1OqRLYu7+NuE/zh4dfko65ogjwy8U72VUVbxGgHlGOJvvbEch1miy1sUcLiQWx
olDDGnaj6nbHX0aH9rNIG1guQ5wxAgsrsdkwiF9CCyikX0iP+PSWqWnB6brSC8wIBNaZgOj7k+DT
XMfjI0DAtXDZSqkLtmWfEe0liNzApHCYZJJcvH99v2JLW0vEheR0LgGLM3uWyJgPL1RWUsrNMd1M
zjuf6J2EppZhMR9VvjIeL/WOABV20Zux2szdAgL6n+qauABgNMY2Nn14z3p/GfLbD+OqLotMZXrU
og3GVfINpu2T3mVEgiaK3eybYrYfFXuUGW6emStA0XFUyRPCg/pewlN/EsquSzSXtkldP70kPAgJ
USsr+MxfKtcG0COpW3T5oRXzJylkJzFXU0C3+DD4EnWudsKlHFUV30zedQFgDZaFfEE+5ofCgDOc
tjryj9bGMeEWFPXe0lhAhbGeLmKzH93LZVhGpmEb1EZX9mcDKaq54bIUoCzK1sR6tKIh/uijacLm
eo3X27y60KCye1PSGOeGOFZK+H7Aqz2rjemDzGGUnhLkCakGrPcvAIsWpQ+6Y3MHD6gW65vWxGwI
T8lAKu7wyNs+SZyv+s/kF9Nhc1iK7O8XAfn7L3JPPsp8yl/H1SpNezMktQWvm9uTk8++9VmkmUiO
LhSRRY/Ont/eH6G34EU4SETX4fR8TxdLouPEUUcOBt539U9Q5LargfsLvt9LEcwGOUuu/yhU2sSc
yXCPKImh2b7oAET1lq6lOicPRCIp/1Yek9C2xbW/8bWlTZHZ7JeuhfbiyxucwQLvLORJigCIrkfu
17HraRpCdy5SDqDOQjgyddM+x5dEjpuQfx64mhZphcax/rgKmn18JkAom4vy0vAbTWRuvjgzF7Zv
DZxBykR5WMs9QdZHLfnproiTZywG21m6YQvdudmtc+GB3mLuXskH2P+Zx+8b+6WaxKCrFLr/+g7n
kMn7FMae5kh0B9rBLh7mBGQwVAVqpV0bMhL3h0rQ+TduNA5PldlqxYmKnnE7lHsxN8MF0ldxuNXy
mGygGA3j3BjuyYqxpO/SOkX4T6UWvNm+pLgXlDMQ7YlR1FlVRw0FkWnnBrauCR12QO+JWWPizBTX
nnmbX6aE0fQDbG6vsszH54Kd6Qd0kyDFzAJ7CVEHh8Mny2c3vS6WylWQX385wASgBKt/MzeQW2S7
d5HBjqEBa56E7sL2uAiwM8I4d1MBbAtUqkpyJxTtSNKCXlAmT/cLvNa4g3a2KqZnjJ4y/0l9+qme
HlBUvhJerXn1mDCvWFJWGfHifmMG6saimN2SsUoI/FguItyCFfb+jy9uQCah/a/yOnfTENix5cfm
4hvtZsJ/YAa2Huzcp5dggiA25Qg+nmroMo/e/IdRjDAFLacBx7qcbuamqs/H61t6TdqBQdGt9o4b
8whoqQWYoWkDToSR4P7PvKQjDF2E7d4zNW7LYliYqZF7QmpppUaiQ2lcGh79aGDqb2yzBcnfy7PU
AkKDONP5H8P0sW9hmvyZDWSfXPfd52+zkteazxUy44B9WS2d9RDlLI9dZ62IIMlA2qpuO8WsVgLK
EhHxPtD8CA6l/iK1Cc2dPmAqERiucBvsRgIqW/FkMlebMlxR4n9b1e32nDDMIWcxS9uE/8Re3Cdm
kubX2VibbQWKv6fV9QRcGTBgF2k+f8oFiZiX+abCiaVmday5uu2o8NO4W5xVevf2fYDHEJFuC90U
KZ6ofqCu6CpFBnMrVy0hEO5rvN/ciHwRo+smPqMDx6/RK1nTx75ZwgT2zzoC5/4O6FuNPsiIPsi2
QLxgkAhl5Y2+vv0K3MbGmGQPgLvp9woAsa/7aDpejQjDVEovhrwTWyHDT5q++YynVopHA+xEM/gv
jmxbV4kPJglA0U5pGC9telM2DUxAEjfErPF/8q2DeGnbp/UxOETLfDLYlckztqvy8PWOU9KNKC0d
Na4CBux70LNanY5Lw7uUcx1wWBi4ci218ky/zos8VWUYySNGgnMOz8A7xiZ7oopIo34dBwlROoSq
yDpatczcj+LdWIqSK2D04TV3AiKHL23p9ydmdIA3/TyiklBHdjDjuKIPqq5CQNuOXsRY8/h6bzOC
CO8jYnr/VS0uD/r7QBAKvAl+KUw0kq2Ce247p5DY6feVBNkXXnlY9k9PSoGX1xRZLI6xKNNYpNwU
VEBKnqEEJRSOzwQL3hD4FhHppyKchV1kVGhgdL1L+lk5FZcGIILOp1UmKE+AErwDEjNGypjsJXyi
/iefbsk4eejn0ASs9tn3FvPOjuolQ0mM9ZOtS58T9/vCTH6E3oYVthLDqrw4DT4jGCujQxkyopsd
0SMbxl8qH6eUFejjbhyJ4lTQg8oYakPkKKictPRCotjfjBJwqLOwwUUPjVJw8/9RxVvMGjSUi4RY
xoeNABsk+x6mngBQuJKyP6WYaBTGzfLUPMVH1n91FAbSKmv/qAkhLSeZNuXO10Y6FPQS5JSybo6j
AmuuwAs/4WjrMO2lTg/sM/A6pJAizfuEqRGd/FWrpjjha1G3yGf1KTeW2Zzt3bIYQ4oM1+eGO6hR
LlpuZWXxwcl6gDvs1W8xuby9yZr/ryVvavkoYdOIfXLnXdW18iGY/ZLfiFCCwW1hTSAPyqLuHywN
ZqPUcngyxqjzbA3acde6YVvczlythTBR/Yu5xO9mN5vi6lcRAIIipXh+9IYw8O5OQvE+7F/j6XqP
8CRvyKvUYAnx7yNtq3i4hyNVHbtAcHrrXK+fdInOGVzCtAiGYUSg/tuD2vRTT5KGvCqHu5HtCz6J
nV1l8e96vSzZ/bm6DV8ni+mSM1lVQvalihWk8p5dS9e3h2WN00mtEdnvDWmwINfH5XV6rcN2c0pg
KNSa+S568FvfBkF9vDmxbmNiLRJZKsiDuNaQVxvoGkKm3AoeFRwSLkr6E1xa9KtXkQ9tUfvUK/yK
/8LyU7rHrcpjpJ3r9t0ZthhXcc7n1Bly1jzEIFxH3xAnDVeMvSD6GlMGza9XC15AYdXFwVhxWFO3
IanccU7s1Fp5EFtrOGHuo3PnkwpRTp50Xw9n60fqOxjj1CoQ2FrJXM6E9Shs5jy7XHn8x9y6oSqD
EVoRlOqEzUA4erKyZ2OyzDZhU7qKu8WLYK5rtrnbpvQwbBDfh2DagcgYn1/Zgr+RGBvedsKshuTq
RfKZhAQKCnrHGh3OyXHwdxznUOWQ0N2aDW28jyfqp+/YcuHyolW6D2PL+/HoPiFYx08QqqmXvMKl
dDG1aUFIpq6pHWQXitfL1q+adjv4Gm+69Yv01JrR+EgcZr43PvJGmGPMNg/X0+cc0ODQlh7wJDv6
IRfH08k1eVnAgEW7wFAKNoljp9BIBJw74IsjsAVJXeQTwfWi5J6tGhYnXgiBVYJiP7iDrfoBTNwS
Ieu3wxI1Jqg8JPAqc+pTh3IM80Lwc3sPruE2F6XGyLodY6mygJOytUs3hyzaUsiBvJTilUtWxYWp
7LVtKKfnQcRCFTgEATq3tqj0ZPJ1xuCRjsPvbOemDFGowTfPu+BQNd8may/ah5R+G/Pr+fV7e0Gw
12hr+AFXt08cdizA8iv2yIq3oiLTnWkYN+GYIYDnEv5nzdnn2iZfO972xfGqvUspdwFntA9s0xgf
DTvLzrRstfO5/80lJa8H78lmPsE2sM8mLy3GEBmfgxciv9RytIvFS+bYlngNe/tJ9abACJoI6PBV
S402M/ebACTIJNKuPk4spbH2RuLS13qoAS/vW0NU231nKK8bkLcXuX31wkxlqi+H4SRj2iREJcVf
vCnY+0FbGL0p+Wmduj3RATI1CBQOjzKHHlrS72Vp9JWuVYlakY9dYH3hMzTx4TB3Db2d2pG7Gbbr
viTyhRmaR1VlFi6/fj0iZt3L30BOHcBpKs6WGU0QGoP5mEW/ZXvjKSwHZQvNF7w+Z2LKH6alVw1y
xjbidB5CvnPrtv2lBQHgmPawnA8L2wmN2JOXGnpoaXrZlUbqDpsGRexH7vLsr2UEb74I2Lnk89wA
OLjPHJgH4XPZ0it4H5FcEPEzczYF/y5wf1D/+Fong1frB79yZSXNOXA6gLSkKMt6s15fYOjsQ4ic
wVh+ZKG+1cILHzk9FZJN1TZ9mPCBYC2w7rFX2g0Judb5jLewuV0sLFlLAjHmz8iW0r1ZNO9Ec6ql
zsp87kH3ZVsYsEPfjG2wTl5sr6sW5WMyZPU8t9pO6g+Al6gTMiVjTnOopinRgdffnq80Dkzv9T9o
R5vIbYvwY7bBWxg0H1Rc4pTt/PJFsGN6m6+UW2D7FMvq/UE+xd1eb3ZDhPJY+ah66UqNjE3+/vEP
yfjlqlVYE4kcT7QzPvmK/avWRXKmhJVMcPjnmzTuGiLMlb1EwSO64e+920p59Ij20qoGSDUss7rF
Cx4c7V1l4ACx1Lcw29tQPVuyzciCjfUvh99wyOwsemhN4GoGI0+DBiC726Am28bvpfWmtrPytw98
FKHRXSX2kqXr9/xEDxordB2hoIjHn3hrhmpjMI2MhuIblN5nHA1HXDYdHoTaKThqgdXzVF0dVnld
jg7UkYEowNlKXgx7ftUjpw/5SOrC3lH/kLaz7ZBRrn8cUMHarlquiRH1vcboY1Wn6YfLk66hdy2d
MgFFOmnrYOi37Tyt1LWGQKhGgdrLJE22TAb7wA+rDMEKQmDhmr02MI/tX4pDLx21UA8V2Cl1TLr5
xej51Fr9jWjN56sE3Co+bZluXka5jpxbvcugXqWykSC2M7CvKnkWiTZzoVV1AqNyXeSfYx8zVJYO
wGPD4tfPcZ/7DOsd5QY6Ajm9iXBY+B+qzkRvKzN4znSk5g8ml7Q5XBmWAyUy4YECnJNHBMeV2mVJ
h8kWk3WOtEsBQnzAv5OcwCMopCT0NgrNQBWegKLEgqnPK5pwWNi7PGy68sa1yo/5nTmghfMzDK3s
XdvuXsxwzIp8O2Gtg1eu/F6CXfuWP5NZOashYv69vGgIQhqjXXp0NMDvPm+A4TiiNajPfF6x4vca
CnkmsK1stptRbz6xV3s+c3C5V+28fjRIQnHwRk/fh9fap1W3MuZ+tRVCG5ZTmDzYFhZTxhF7VkB3
DADv9UK5SAYkuKfjle4HRtN3+hFAPrPuTqSod7eZMWG68J+YHI43kx2BYGBwz+84Ej+O5890KRH0
Ow29c0Hd9A6VMoKABfZmVkNHwQi6A36W0GZZ32Xck+9kMkyGNWMosMOSSw6HmpSMfv2MsH8oD4I1
52ZGGBBNuI2eZkqqfI1Yx3lLiqm8mRHsMVvH4zZ2xv6iAsndTxctB9cn+E0xgRTgPFrmtbhCDSk0
Qc26tMswXQJAJX1foGzZhBQF+MaY/4sEWH/jECQcYkvEKFuArXbiFvltVYKvmXtg1eapFfGPcRd5
LIcQ5Xkw2iamiUHL2GjHstFt8hIE8WZ2CxuHU5HUwxuFpKglQOjdw7JBzTAucP9LPYUIszbBxzt0
FoA54KQrNWSvhzPQaujzvi+M5SA14Lbq8Ioos5g753l1Cx+7Uq6Yqiu5lAs0MsruCQrxblN48bq4
r/9UUOfnHl7b6QgCmCs3tBv5ygjJWLo37+X52aA9Q5VQ2NDMjJwY14Mza1/CXN4xNZBaSY+uKlD7
NRIm5Wi1mudmWqvtZjha9zfSzjZCFPYHn928vA3B8RWHUh4CSK0XhcNY6NyRlZC3GeWiYH5Pycgp
ODVOPj9ipmISRr5jm7RTP2ab2h/cxfftsTNaP3crPVOEfSByvKL6zjA1JJoFox1oOoCP0ruHfGBL
crki0jxuNBMin2Q9owEHPq9uPEq2NNEC5ULKaN/Ci3jU9fhN63IsIm5T0wR8+AtlpjctwwcgknA8
xWH0ImJaBQcM1gfiCzsQ3Z26HoHyISjwnCTJlpCRKQnth5Ug/8yxIBwqYkggbSFszeKWkDRF9bL3
nnIbk9Fr04MObfBsZaVn2GC3j9BikfnV/T2CC7KLAlzaUQ7GpIYer7cqvaCwOse6UXOUjl0uJmZq
7FfSuFDGScq3SrXLFuIo1mJ1sAfPGZs4xFJPjb6k+ikbzYUp3VaRcmSIvuS4Z3p/pJybjXcJkc6O
ZeB+sM2voducApQuuQAelRTU8kc1r1mFIo5GFo3DKYLZ+bUwQv07wIQoJmGrvBmL/WalDIs/9cQz
XxbJipBiStyBJih1/G8EzYthVt+o364R/ekhMneH9py3wJTAN75/68TlMdj52q4mJsglzvprSmqh
t9yUue+581dnjwOL7Mpbbx7jmnQGhRgCzNp4gwGI+jntCkY/IDPIJPqg5yKtuaUT6xFa7uWelvF+
k9xv0W/BS/c/PpZgPq8AGgCUPrrBwZ/mYgljjpx0OtsXDX6HIonV5OS6rYY/ZcuI96tYpb46g3xn
CBkwNxGZ0D2YyFu7phz+Gb9lJtwZsteYMee1cdm0+umj6d0V3HK/8FpRg+CnIcVjj7DsKgnhDa9m
twnHhYf+/XSy5FLWBRE8bfPnceBqekcldgnlZHOqceF+gSPb/gaz3IyQsoSGgt9yNZTZPWoDnEhL
l3o2zTXBVjxq6VkSWJhIlCaD553jwQ8ROXw2dVZRwQTzNq2aJWPJeauLn5ZFjdPV7/IdZIlAlnUt
T7SDuy5juJtpnQL7+QRUpNObY7tC4SVBzmyboz2NVng4hOQk9F3NLSjKn3L3ZPiosC7Dej3un0r0
s7LIiJ3pdOXCHmqQMfz2RWu5l3mVLTDgPD8AimpQa5l90dLTXqbGzzkr3zO3yKw4SVfXG+pi+sIR
E7QtW8aCORk9k+RCFGGtrjXPG9wFuHwjMLYv1y/Dgn0ekIn7whmb1dQZNSxjxCdpfCl2kiGqB90P
I3XZJ8maBlzi3m83jKfijLUSSjMBL7ZO36NrV9fE6YCW52wkgkt340I2l0lYm4YF4IGzv5qmJXge
bEyvEBeHeMFM88v8ErG4wqiZOKZsUw7wYnRuaBBK4rxtKZi6Hfp3FRlzuBW5SLbFp4qY/iYI7JpF
6/4k1sQpmSeIP+AqnLC6cSuxnPZr9m/g3NdDv0QpSl9qMn8/Tf+zrjvB2YJlvb3a11O4pzOBqjvt
F+V6GcWDpMIsVrYxep6JyLaTF3hU+3DT7HfxtsPnkkkbq7G10yTCSxAoi59IaE+vjgVY2rGeI2Tn
YftA1EAV5hibTMNYOf9YaQuEuO4jkPDn3rd/tJNX2wNN3Gb7hu/OxahAsdQKiy7IZ6S75HRTPpWE
5ZteV2J23Pxs4PM3CxJJP5jj0KCtCQBpY1qy0o6BCQpOmdiDTS7HQQ0VNl8TikcIptJkJ9RJzPcj
XOQOVgG5TIZtrLrDkgfItjlJqumWKfTH/fG8nul10+LJIZZiraklOz+eH1XKWuKJHNUXCFV9a6za
lQZSUP/WUaEnf52RK5zs+juiHa/VFg2L3TgbndU5c4gDt3m6yBlY+UAbIDHmP1jbWyX9EfZM9T2d
SHRvixR/P+w1QJtse6wqLrVNTSwtEWLvFjQnQKdaYyU2AzK7tCtRUWS2S9KJdzzcgrFYC+AGE+T6
foQOKJx9panjv73alD+lA3sgiBsMUbFBOEtO0AOqCjeruM/9wqxHq4TcM24ZSzi3XMMnEwQ/hFyH
SUe34TtL61L+OLfHWk/V5l80ShWhOsJBuoKUA+VqeKw61OvwH9CODVe4v4IeUo2I0Qfcw4b2Yk46
fTDwFuU3EJAp8YIRSpf4IF4XZOo0X6oCmX4LZaGK83X63xyPoPDFq9KH+T7f4ADK3UJWAHeSwiWG
5hICtgiktUCnVeuQmQr76Acm1gyHTOxqr/ugox+3u48aQZZ+CK6XF6GKFdik63N8YOA/a6bD6omE
TbCkjM4zbKIwlFCGt6vwV3W8Jn5OzQ4QjeX2jYOmFC3W8Y35RsWVva8kXPxRuTBpQcad9n7kcV1Q
b7DRERIDtlaPsdcfdMHyPr4er190Udu3qqY7BXaec+kQnrlSOZEC4trlSMgWE6fTEKAO3K6Sf/ac
33kDgnKByG+TlxlsX/dAgmf6exZQRVJHuqpZ/1zjXAS4P8f6lJ4ZJCqyDPp0ip2v96pf93bGocUK
y9ciMEjbln24fz7/4stEouyCwevq77/IGIlT753ZTfZIDMXeV0edW0XkNTUr8wpIuGz00LgaEeO1
a2ih7fT4EQcQVmCNmiP0a289w2obrZ3FJkMQdFqMeZLMbuQEeWXWqQVMPonM0/uObQj6YLwIosqA
MKurcnYBRVovjfPX++PvvF7YdKEoR3ZC0WzRQoX6nyhYCHUuOIylQG+LZnE9whvfg3HRsyCuQWqi
Oq0JOhmgVwxKgQ9VtaBb6QXgBgys83ntI89FmG07eW4MrSY3pRFvriKLgYHNjd3IHkNuaSmO6M/B
ax/Pq+noWkJuzcwKbgwts7uiJ8VicV6Hg/enCUvPJz3FmVF6Cr/Hf3sxL+sHjYeXKQYKXVqIZAfO
luKL7S/V4R0416jOcVRk2fpsqvhvxS8r3nLoI30HgARSIGWXpekJ3vRHJGQKzueYEhljzmCJCgsw
48XHFzsNFDxPyW67ohqOkleGRndlJogqNACbTZ2j7uMzuvqy4eYsxFpIe0trQ/uzXiUIU/net2an
eJf4fpLrRxBgO7Hu1BkoJidV/V4AOCdtUmXQML/O1UnOY1QhtcK83kLsbcgpKPPwz/t010mxSOGZ
HPDRbnIVu4YDP1dnsVXxnnUTNd54zZDsFP007UsCit4Lv6Jb1etFGK5e4g7RAjiBjaPD1qf6qIt0
8t1s9ZrYva5LkNxANln7ib4btIcPGIodAMYUXjK+TASqgZxy26GO7PxoZThGj3dsB8g31r5BMn+o
ejIxzb41sPD0Io8mt3THgpakUttJuL2x7xYF2R0bxEILD8uXx8b7cd0Eaf/76qLDoGktPDbFKjPm
XRMGlPqQZy8lOV0Ra7xU6UvWSXFyX5WklzHhiTFTjvLDhsEZmgrIiAQq1vzUypiTQWWSvtEQUcRr
3I6KGAibFNn+iLJQKOSwK/3VlCN/+ViarTyfC26XvZFTbmApWtj+CvMcsh7/kXdlJhYLXwpy5u/Y
N9dnc8Jj57pOy4hQtryMgBPqezGNJh68LIaqlzew8wwCjMgQtCpA0VC4v2BvjkoNVJCyVzfKL+xI
jVvnvlFNAsH7s3KUDADdGRuFOvIuTX7I440gUa3iunhZlvbQIkA9eEd0sh9F/WFY0B0begfbZ4Sa
vVnrho8zxBqmCfoq5ayhcURrv57rPj30g3MgYS5Hgt1dAWww0oR/y/piBxgRja1zKbc9X6BXFn6e
sTvXh9tpbPdXULkxICtxvtDPKbZ7M2Dz4+X99UdUfkZil1KJe7cDtYTGEsKUvm/Nl2xtsOXgMD2o
Fj9KBpKrSLpMQyYYZw2l5p5yvq8RDwUCT/H90nhPyMmZTicAYO+nfjp6eiETaKIzTxJ9qNIypj59
P1q1QFPxtDyrUGC3uBWr6zAgvBrG9RkJjQHK7lr7yIyBofsmVhnQZqxeL7lReCP10KoTfReYUsaZ
sTd1a1Z7m5N/ZViXSjHcx0+9cenV1xxYU4wWfK4gAPAkDfAYBLde+ULoDVJhqDW3zVE5cnryfC7O
UkzsBgmhDnVbw841nyN0/nw8AkWOnTdD94f78JYw9nzDdo1m7EUXcLfQRBtlWC20MTPVwnBmw/gk
VNbgLzwW8M7r0mY4dw/GQbUpFDj5RygM9bMPcdDCaUUEnxfge7GtOc3EG5jLMH+FB/4hSTAEFMhh
gBGeT1oPThe38CDl1f+2vJmSAYxncafETioHWZl4yy7wVtMXGirkPKiG3VvcWeapDoBzOjr4KbBE
Dvzl3vqxOA4lFj+SJMoAdnWkbmev0Yd/RupphSfjT2VdGRq9nihJV++mCxJ1oyTswcUNAb69m758
qoj0WafLGcLLrmtrRbfqPrP6taGTq4pRlGWwtL6BcJTKkcPSJwfUUyRBSZgxNdrA0Yx0V/d6tEnr
NfDhQLKOFYEbFr5MLZ0Dpj+xzdDR+teuanweXZGtdgX0sorLTlcoCLTBT22XiePpBkczUvlWjixR
RvkvFwy9F1L2mIBS5oCTbubLCcHO/WfS/PSJhXne6fwjJDQrnghQ/JTAXwusTBupYHpqMGkYnDzy
zWWrq1fYf3ZWF9xAdD3m1FdShKcd5/QOG7NjpVE0N9VCdbXaO0yA9wMkmciAO1JmsSuIPlFSE8tP
3i+IfdazwAA+KlKOKqGc43KS3JeYRqHnIrrp9r1Ss3oNJ279dJF2NzJtUwCCRaoBp4Rg2Avo1saM
7gI7APaa9eYc9tcZAb0KoEALp6dWzBJYKI5rOcH1mtNi8/+gHRtUC5SBfSCGLfWddS+sn0eHBefn
BUokYE203bWh7o4uVFgTTyort6diK/PW7XP7HNu73vlyoFkmT8g0A6VFQfXqhM32crrLpS05+tu0
R5Yykz4esHPu9+voan3MHFeSUyvw4WhQI092lx8DU+4ufA9k90D1B0Nqx1U/qn4pNz77LVhmO70D
++LW+k7BvQ7kGlYXg6Dqj7pHjlq3PT4KE/GLbt2wnAGCne6+ZfGvm3+J0So80ZHV8DXNs6MHBwUw
wdsFAhp20pjbLW/PGJ55fzVCFsScHjYVwXeuXHilAQWtiUeqYh++U0z+P1D6q7ddKLPJWsLi04sm
epVNyUyeO3PFkHqsdPINfIAmfAqM1Ul9r6gjTGu0Rs3K1MD0qdmXbYi3mL9i/9loHvZaA9P8cAfD
oXw/r639vb283Ab5uV6E17Ytq5USy4MTcD1b+YjI1oFIQZ+zePTEVEiyKqKgd5SIH9ZUzsUCHsRR
PAmO/C35/d1IeOyctvHZKq/VYie6D9bhp11uhzclD46cdUYqzFqK/VtUVO+GgqQiKxtPbp5dbFdR
cYx0SuGIHtA+EdNllzHQv9ekweN605Zj3Z8lHvqnhzh6IHxgM0fguKrI0J/+2MqfLGnewanZ3Rcr
rFr3ehlVcK9ocZP36h2YjPAB+FFLzxAnvYEJOp11GasEBW+5yCjTL308WKXhkqog0yT5QqOSJkBn
MVLdvxRDUXvCqslzZxUA8mQ6Y7gPF4A0CvqfdfNLr690B4vQRGeScTUWG5FeAzojGmVwwnY6Wblz
CwUURKg7mXqW0F3xc/t5eFy/dNw4/aydi6hGx4Nb3bX06DpdW5UqFq8UQ5ymqm7U52IyC7E8nKVY
55G0KMdT3IC2A9adOzy76JCk786dbO7gKm+Usxx+4Z/MH6xMwc5BaQZADcwT4X+Sdj67ZIPJw4HJ
Bosg2r8vyXNiMRreW9BmpZnQiWt5GOPPl9R4Vr+TkuKAUPGG+PAJlnF66r84PadwOS4Kj3XquP/d
VFaUdOx8nktI4h2qyW+KVthCpkISOjN4YLTLbH7CTDV+hg4OElh6MVFe/PAJAr26atX69oYDErGZ
vk8sdT88ln/LsiQrQI+Bh8XxnGWZ/2bCa8PebQhWZNZlHrhAb1fjA4ZqxlnZS9LHR8jLDVC//o/8
tKYcJqLFgWKea7xCqzbicWCBguEimLOzcnNniiQ4VZrIVQ0kWKoa7UnZwGtLbKnQw0fYKyWq5XHZ
zTlDh3kbKcm300Je/L96j83L5CCVZiJ/FM9TskBbIZR1o9xbrmG6AJ7GibATkyv0znxHIucvNLQy
DZNyPaPT8aZjYXMtbYn8M+5b0JoO3XVUispRsXQGJYztwkEoZFeimhO2ul97xaejf42TTIOelKvx
BRDjwG5ztk+a2ewePZq8vA9jfPKQemvaR2dwVM5srzXEu+oyqRQPMt9Gg/13eHohOtqZ2G527wHG
+1vPXtDqDRx4IzYnFTH5Fr3uHm9DkydHz900e/ieLuieMbA7M8uzYuBcq6BVQPYPhsTp0DnIXki+
+cU7ZfwaZmQD1c7J94ENJYnK5Zo9gzQCVWq9WgP0A6tu506oWi73zTVnQOZUcBRifzhJJiVcgGP9
+cDDHA6orGlPGUekN7Gjp6gZT3nxIWFJ0Klb0UUQ+O3JxTWApqP7ew65WWY/Th4RRhZVRLbObyQl
Tz+nwCi4GX1JOwBriXs+A9TsyOOwrmWTPLRpizQxCO0LxyfQdq3GbdKY15tjyBs9UzV+c2YNfQg3
goQsAZN58XBakWDoUThrk+tbH2/UO16GatLjj/Zb/b8KxqsHts97ihDzYUBjfynW9vFehvWq6M8B
Bd17zfM91MAXN4CR43wTgeWzSTUiWR1qyBcInpcNEF7hUtGC93f5Eh64B/FrmHm1QRI8gLTsf0Lu
+5fE/rYhKK4S70dSOjyRxPpsuPfTtOCZx+YSAoS7L16jPMafLP6/GX+Pfz+VT3cIejcobz8tTFi7
fkGtRWZeDxdmsQNqmWiXEzCHbesXgeAEoMYwDR4kPOLju1+Lo4DO4qQIKUzqyur1EUL1725vLhFf
itW0mQtVD0x1M0xBRWosy2BGnltJBNOpkUisvrhoI2rdSZkmdlPDEBk49jh04ngwBC6l+W33I3Aq
ad3ZfLumZVKhZiSwL8LUhCbaOsmvwkgPzIfJHx9u/bAKOlgltxJAvSbb2hwE8Jzh2Gi49DXnbvoq
x++uSCZCPuwxXjJBC8/CP4qEzOhms6UzrGRaZRJTRBGrlXazoSov279eFsOgi1+E95NH1b+iw1SP
IugVNFaUjLDJHOIet+FP2Mtmy+1sK6oF24LXrZimDhg/JjPgB7D6qf5CQKsy4ha2n9M8P7OX2mIS
QqE2NPPPBm8yvrYa0AQ0hG0GG/xMvUbjWKXyqPk60GJQ9SjI2KA/at1T/xvfSmUfwy7HRJtYcuPG
I5CJPTQDyMSb0j/skANNRdAPLuvJl8jz0agcRfbyekSDcachpDpr6YToWHxrXp+9/QDO87psCYn6
b/eTrzV6R9zD8AY38o9GR/wzqFC9SRxwabe7+TYsW7TI28vND/ZNmrLLk17nM3nGs64tfNegzfo2
rN+81x8H6crt64dTC3IMa3kamk1/HYFDvB+WOZWKTBdnKsu7o5TYREvMrQOnLaCp6XO6nzdE0loz
IdmbQgN+wN3F1k+1Kubmsq1vhzLLUDjLbqkOmrzb00e7MHtFcn0+OTHboilO+XgMP5PvoQHm1an+
5nql6CNr+BoLbXmmZXyiRrpOsJOi14dxRfdl76Oj5u6LxWXXUhaIFuwhsKdFbcb0bay1QCneCqJ3
GtQjv2JwKdVA2JIaTxvU+qJqucsycIV6ePVx4oTjF6l8Ly4dR3E48pkChOerlDHEcmXDGadK9ajK
lKAKYCaApWJVmBmbxIR56t34wknHQ48diB5Xwbd+ugE+vyoZ73jKoXuVgmG3TjKfD+xkx171ghC3
c2DSenhO+e6YkWDKNfwQlX+sf7Y6lVKZGfH/MAksS4y5Tgjw1yy569eBeg7K0USdCywNpD1hF2hU
jNqzDguEoK+A7MH20MQuD0D8Raxr+RSPVMqNj9/xEdCtxF+GmvCR0bovemNm8kG95v2ST1fmg8r0
R6Sn99GzuDRbs+jOjiuskDdpigaehMs+WjZfOTwOBnduU0tk3Fb74DE9VZTXOs8GltZBHM7EnoHz
iEkIQL4bLIU95KWqieaHsxPzhYX5I+szIHAg/NRuY05SRRUSnrQk7EwvfxRLVthj5KWAcuvup1jC
mo99uk0bk5IyXE/MLocGQJvj4v/jABRA+b4izaWsV2soO6tV+gr2htaTFnUYHhHC49IfowAPp4Ad
TO5XQ5pH5E7f/YchTcJ12FSFSNYpqEhZQfejWvXpNgi05TYp/SQP762rFQ7PKlovMb8uWqTLTpZw
OJjW+hYKNHCxuboCmwuiI/PPjqCKDNdbum33bskl22HH97QnNmpiCcxEiCj5pG9uB1uB9PR69/Kh
lLETE0/Gmrf3vBWTyk8IwgeTgBTwllSpSCypSVUdpmHCmpCSZbUQHpR6LqX2hpL7tUB6KC5aW4jX
5K2nDysIXty4q4MXeHKoF8Vo+Y6k6dwi8fbm6G9OHQQUSnQTad5czzavSql6SpLQGwFjFFYs56BO
/g2DcWWlXbTTPfZT1EjnlJ7z8DJZnQuoNEw4gQHW1AtgYEc8N+W0x7YNax6App9XNebWjd3WBh03
c1Wvp/RMWddPKFcWHdQCOLtAZ0z1PBLPSGFe532QGO5rkqqPKP5EsJXJRJDLuux3jV+sc/CV2C9y
R3FzB9Vh5R/S8mfiwxP/SdfT/n5i9jBOuoF1x+VYoqPTmxuP7e4QeBQ6qhMSPXkdqwUOGLBBPyjI
XiH/lxh5JvLqHq5+MqVwPCqCK3lNSYgIRL2kGTpXNY7SUes7/VEp+xkemJntdT1++4FIR8JQhQnI
9thZ0pTZLKdIWaUj+EIak6yiWowPo4tEnCuZgCKCfgRoQd/5XXf1Ol1qhnrWP7KSyTIBwMGn4wJj
a9B9vCvtV/Td+l1v9t9VMF/seyLoN+dCAk/JZVUFe7eMnsfMp1sJkCZ3LAchNSCs539po0xfeCkK
HkM6z6Mt7XToMTA/gt+8oFbZensqfw5xoPe/zWy40aJlg2dRKHE3TTv3rDniXRMpgRlmM/UKIDyr
3eh6t1lb6uVk16/dRixnd5JFrUQ+Yd0ihoUX3TtoDpJkjv3GLVfySvc8vz9gtbNiu5oSqINzPP34
FoMd1pQiSN44zR6To9jpDmPnrts5cjnJVz9hieH9jy2EyL+Wzvjtdc1iziYgiUFlRkOeP3MHGoys
R9ggYNA/UolvasWbjno59c6ThjcFPX8vehZOAsqogJeqZy38PgJLYLzpWRIrdG2vzhBIep2/AtFs
ssaRDe3Nw2kt5vj/K7/gteCrZyV7yTjrlQLMc2seWkOFcG00+RBITUnIiN0/JVYvpgF9jQMRfxJy
FYnr9M+Ys3ncfJBOmoTRjpqpM0GFOIYigbf1W8hDXSkZw+qYrDQxY77lyqSWmr1L4arHiO9kZl62
Ud8/NweB3a+6FjOvE9psNryxHfEmyMkRLKhkUE4Qc5qMzrFqvYa9DzZYDUthpNScJPOHn/wd8hlu
cxVYBXodMy1mfbgu0gbXh+1MTgmpEGdrAxhYQVjrpkdwOHpo9Jpjuen0W/zZY6aDhdR/zrtjP6Vv
i85PupdRcvfz8Vc7H+1qiln5Wx7xqD5xHEN7a5yNEyfJKxXccHdlCbh5dyCjWedm+lI+eg2x/VDS
4ff2RsWcFVC4rUZJVJyPl3wRWeA0hAKhKryp1pLa+z7HBuYOm9F9+wbMfIoR4PL1Cv/UaghXyidD
TRMw/inbRW89GckWoK4pojERIphr6ez63bq85k1s0KSBL4dUvCAC2WgWc5FDla6Ct4gOAg93mQnq
ewPYCwjofBcYYcRPWQyMFcNsODakY0G0OFYeGeA3NqbXfOFgQzVWC8fSHVEa6YTuMjp5J3CXfgG6
b+uSORDhzvDBLeRxjxYmVYZYuMCqRpFrC7kg0vsIc4aQ11oxWaY8ErdjQCI3rYLFksB9qZJvgN+y
LQLW9IyYvDBeHmKMOcvqoPlvjHHiEUZ4iiJ6zDOresb4ctMCH0G+VU9tt1G7HVGPI1UDECjZCAow
h/Nu6n49N6F+Go0jMPREvOgHFA12D8J+QgnrdKuJigNR613DZaYYWEe9WUdJ1cY+7AbrOJQIRMMD
P++N1G04hAu3cu29MC6J3pvZuqx6GewaDuTb+a/fKLqkZ2/zKsHm+KH/t+wQrZkXvyziyHkUXCKC
8cDyVb1mJazQ9MDKywHJSsakYNVtdZdqqr1ORRrwZVbQetKuUw99RNfI0DE+u/asSZxPYlaKVVLB
lEkfDTZV3yRfZM/SKvgJZthAIQzPBRBmnpadMlMIWzLNgQ0IqkteaPTB0LrsBuWcX40XS77MHDnq
BBHtnbbDRqBM9/VvRKz4ex/2QureJOfyW6lIDQNKjLqxpSGs4i8I23M5F/4cr1rl+7Yansvq9YNy
FNWXcsCFcE6JPW7MEGG/M1Zz0wrT2HsijOKsS7S5MOndW6JDkB0S7MSNNMDYMqhtJV4Saq6BJb96
LJN/MOKxEiMtXJjl2/VTPyr2WQt5VY1XXoct/xX+N1jlTkPzRT/UhoRcvus0WPgs1ZD5InNfdEgT
I8+gQGZFW0pJnHUos3WXS6hqeBfuF+fN9EEJ8n8rnFvHk+T0yKJogJcaAgrTtrsVN/17bgjaLedp
+RmucgBnwtSnIzQXwJogPQkajZ3PXyo9xtb+Xqy87HWKTeSCeeV4HfJXFx4pjM7K5EjAkiROE+/g
GGz0XuDn/2iwyDsm92PlW6IuzsfFu7q/SvRejyZbOsIn3M8FGVCFhgT10j9+eWNroXiw7oY5/wQ3
Y1pBFWhYt5wIVcSUBTbG0gyR7yy0TFUecg3do2paTQoaXNoDw0tRiRjaM7QldowFLzCq2uHlUIBJ
wRbKr3piu3Q/hvsEomW7lj12mkZJKFBLKlYrdpcB5E2RiZxXdL3KfcZYClvZQ3vipVSWrPUqL06L
4yvxUqkMhzadzV4sB3d3xnirs8QFIc1yr7e8BfUIKC/kVx5MqcqekcgrJtC/NTHZXLUYF2uxzwIa
9uF3etQ6xGB4OeGRUD+thI0xwOrl/fDuvMI8AibLLvndvTzLKvfPpqerRV4jK2SU+wKzCzlEPRwj
j+lwzUY70CyQU3HblCv9Kf3Mx/Kz3dqTFeQuH0GYwIwfoJOoUxFkEdI3lUrZBpNzeE8eaqLAkgNp
y1IR865Rr2oZS1x23LM33dw22wMqvLKMkqupA1QUaTnLqHGpzBFsDb5sGLzuhn9I51vPzcbQZV2j
8dCo9s3IqBhPyKE1uTu7iZIvHMyU08ZcF7eH2ayor34HUZvzFJX0lmSYCX0taScgzQybTfxoZE5J
Q7HNqzcTpy0bMc7mh1yDCmCrHWR7bKS+ujy0RaeTD22E6adT50PMG9p6nKCfKVWb/INqrLr4amf2
K0adixd1QKw2RWE8Sw6xjcm5YeOxKLppA0Op+kpQ3fKmmV8JHXf+0oFGeTpAeGhMLRlWkpvYZIBf
EU7LZtM2bODzjGw0+YMI5ydwEW5yBiR8DXo1aEBrk5FMViD2odguzU379dMvG4FRayEosq+9HpUF
qqMDURaEox+FPJ7C/LBIuJuplS+J1mq2gvFxrH/VTzyezLc9Yn9dz4+3zQmy+n5WEszujVHmex44
ue74YobZpSvK/A/HyQlJxmxzjmNfto4QmiODkqmujj7nXg0TefCt2AoVElxnK0mezDM2TjrH65HV
V2Qyu3zlU8DcV+POvhqBvF3rry6qXSZdNeGp+JWAbB8vJUNjU3TFwe5oJQm9twlDIT9qakuHYQqK
7NjMn5PcfqTYJ7wGCqU/6Hcsi/VEKnQeT7aqBis/9nKTaS6KvciVj5s9JZinpig+XwQnkiZhQ97C
xJWktCwfIoRN065E7aZ5d8jRacms83AC3PXUnM+qcB1xvOwQChVE9jtMz3TqlvwRR0O/3AOK2wRV
SSMzViMufr+0t+o+awbWvBArPEbU4ArocSDGaJ3kD5wNzqyBxkCIdzWVdpzKqhsi7BYiE1sHK0az
EEYrxwComZRfVHyx38EO6CDeJ8yF+Z6H11aWyXIxm6gTofiRMmqzKtIRmohFH4LpEqHbU9/05md+
d6OyIemr3TttzXNhPJ5JhwHw1YhCTXDpyTpLq85lW/WDFf9AhM6VcMHMTlhvVp39XxEuteN3PmU4
JTSKluOAuY3n5GkqKH2JL7Did8DZwOeZLwUeWkqHtRetyP/gLAzN8O1YyaVX5lrQOlEOwd70+VvL
K7q88F5ClTeKL/fx8ACJpxnNzvYQXKclSHdJxuterDXQJVUFSD7wfBCvYBGF78JxpHFQDKwzLBQW
ze0+LIBkEqAh46wMR+pGc/TQH4Hgm/0Dq2sKdinMt+lGJ3YqzEPSyUymmztVV4QxKWZUC9ruCdH/
v3A2KBRSzg5SVIYwe8yCUtrjhA6wINtyEj2W1MVePhxAksGpWlV9d8CgkN2natnsoG68VHwRVG0r
b7jKQneTmMD8Oq5zuY2A+bQhXkMzZ+L+STn2x2U5DJON2iAOBbgi0nNBR0+Kxzr2V1skJtN+L63M
6Y1Q8qwU/4YPdl/w1vg3p8gPh8dwDOULeyrWotPJ4+EwHYKdZihfNPqXeZ7o8PKctwtHkMJiIHHD
ECCSjtgY1GRWnQoY+JXtcwpNy4KYYLApkGYFfvEVH75TLm6/cZ5MGQUk674i+m2hvm7nqRJmDkiT
lJD+dikJSbIbbRLOlZXmGFYZXP4k2cN+QOiV9qs7FBRixPk2nbXAlhgp/H13iJovPNpEuKGdJKVc
JyGh9hNKm9f2lJu+TFw9KhemhBFx5ppuIPSDTBMgR76/nZ2GqL/L5Sxc9ZL8kMYHjn4qwqiU5I9K
9gyuOl23LvjFZ4Bm+/7VQkDgl2VgEPNezvjwPmyTeVJFcgbJaSBYKJ8zhf01dxFVYAYfmiPsK4Gz
kcSUO3QWLlWbo1VIP49fBjQc5GWkqLRsjBBgVk78Ls/gRUnD6HvycuXPIY585WIS0NqAuBMQHLMI
zZ45h75KlkzB8t+Z1TQLuZiollNAvXWwqo3yoj/AP9ZUMl0Sivekqd6626zyEgwxj16tX0yd+NRZ
MK1kBVHHyto+h/wA24bYMymDJLcyobenPeVU85MwkLthNUNece/VgscGejYlTs8swVK18HBu8NDH
WdYVJiurRwBdf1pTef/Ua5u0X5AmY9Wj8NRWWuJzikSfBqKeodb9WnSwdQUms3xPmwYw7bsYi4xR
BjyGdQnAWyOc/JQzcIr2XMV23Z39M85De7vH1u+73nYeHnhFfsBJldfvwFHHlI1Ni4itCeplvQCT
w0xrLyKgJdr60MwqRscSx41gy8QSQK18qsJCdULmsVLEhOsCswV04O/H9BwbzjXdttRE659D0MPD
3pnzoOXGfGmi3kVjd8PKz06RfEc0eMFgE7hhCnMHVHXZp7RwBA6IM8aIf6oKaVxkZrTBKzXNp5sF
eCYzj9+egb/QRO5dNBY+cgT8ivCEZmpyyGzeS7Diwwq4IqSmYvIFOBRgW0uEJunEWhUlsOBCPXON
xbo+R1nUP/+Yg1wvmdYkQFUcp0P4VJKk7WFzdbnBdiBBClXNafP6s9bt4f89fP+Nd9bSUhK8iI3Q
C1dSIXXlnbTw2oXIOytw616Uw2VTW88soRKFolgSUOZJYXYl40Wlz7rKrFwXjIkL8tQMZv4qbgmO
yFuxgjRX03bWVqocCWy7B295qyK0sk50kvO9Nd0YUvpvVDKzGa02/eWOkWoakNJ/jCogdhrcvU0m
dpTLOtBb5x1cCGL+8VBEMzAxDKxbXpLliDW8H1yTQSu52h9SpIJlApVR6cU//lGf3YEGjAgBomVS
PL+/OBTWiY783I+7ELPrjDFN0DgqYXtlHTIktcUvGcWUWdUvjzJnv1cMZe2DEr+HXCh2rURZHXPD
EWbufuVJUtTioRgO/tFehf449UgL55AFBSApspruoQ810759MzkzGvgBWDrSkPIqpnsJ+P1PGC6l
46NS821KBzIundzlh08r+BwtXvNpHlF8weQWUIMYSMb8Em4o308FK2xyyJVDu+AGMJC2CRjV8Nco
V5fKvJrjLhhdpo+53kGbvVLa92M4CI/Y6HYE9vbDXp3PhWJtJQ6h+nOG9iMNh5Bul7VpRuf9Ps3L
+JhHkhaP5ZJkmzETaBcNIs2PA3ud6zrC+2gCWSp0qLwm7pAplZq4aahUkop+Pt6L0ndaXKwfywmH
wqzjCRx4MqfvZEKDh+wrN0/oj9e9HJxCY6fuc2N6e5fhiMeDzW7GsX56AZgDBhbaVYkyzFPfj2yI
JL1+4dOBCAAeYA+KO0Is375GcOuzOjwlqLKpnCT0sOvVt3DOkciiGr8pDqjvWv5D733Qf/qiZPA0
Gv1jzKm2moQEXKn/4O99TEkhZkBB1Q315klLqBmvlxgEedUWAk0Ph1lnod8RwvBLpstKfdCjLaff
s2VWz5yyI55cQ6A3HSBBZL53d+K7/IioQ4qWoyo/8qr7tPXJS4DS8N4OcPi40UEpQ6aQKlc/YFX5
qG02KS+/qfGY+C4W6WCygq+PxFL6uY4mct5YeBwi1nZswfzZTeZWNy/maADJq132u+dVr01rKcWI
RHtM7GKDjKzyWcW/x0qkPddNwlEBFItvlPsBiJ7UtDwpHf19XFEkOReJCyHrhdDH3sJOyQ8FB2Q/
TjKP2rR28HkeOqOOBlBsyGzuNfIb6CCgv6uRvk4KU6ImLlP8FKPW7qtOFFHRCSfIVGXxfXEDMr8d
0RuHX9YMgRHqq+p722jfF6IJtp8VaTpi8JSHvPjnKHvtTJJCF4WahU3Qk2RBtnscNnxbqHqJyXil
HuCzubTsqVe8kmFSbBPeWFjNqDpppSaAvV72jrM3Jvm9t4id37m+ofBo75PO5Ls8zSzp53diszMT
nz4c2SWoeqUTrRVQRvHBkLb6CkXufjixcWmn4CwssNBQe/g8+T2ok1eQM5jKv5DLU862oG+W0ntA
5qGbRFYvdhU2RNz7t568XhzkqSFngbZazWhUZeT+aeKMzvdhaDcC3f0iBUN9N1pZ4oPwiyr7F+kR
NS5H7Z4+ATapTYhApBZ5e/iSwL8WBiCTqw8N488MgZimkKUIYDvA8STCTpa+zKOHO1m13SWUp0BE
eGowGEiZQIBUogw2U3op+XQV2siYq/jaxoXbWWDm+4Z6YoWSpsPZwmF6GnC6BatOh4UfEIU2QChH
iUI9IgtWpK58Hn1azTwu7myTjXvQ0M3oc1ApBC3R16KGw6odyX9XjxHFY82QOPOYH7HlXuWujkAu
mKwpFRUbPSdBW92xkHEpeRx0pcb27z9DAyWtA7YtshddmdOyCDJ8YfHLkicBP8VGySFIUUeSZpO0
5TUHY+/UXyjbVUqrOYrcEMUuQ/M1GzL/wGAZloAunUTxbQSK2mDNF25QL0piWGQ3xB5atuSSNzoj
+al9vDVAvogidKAw0EA6+LYy55NPQtWSKusgrtdPrbCOe1ka24Bkd5109CjoHCXOmlgK7FcIpbNj
uXSBTWv+VO+1+QO2khsveYQTv3dpdXSdrXkExszoaOzBIeYnpn+2bTLBZB3aWS/f8Bc07X3AqnqH
JP28MQp03hXyhg214ywDr3L17dXxAjkrgDL/6UEtQW+s4y+PBPC2k24EzZm5IVKGPAmpTYsMsAFI
xRMWNHec9TYZT3IyKNxC4OsGhNySKtep2usdyqNUIRUp7a4CH575GghzS2Lh2rUDJlwa1fdZ7pro
QZF/35hQViXgQ01Zb7et0vsMTbGLOxzwkqx3yD9kqnR4kAP/htLw/wTKP4RfpcS3XiFGSUBdIpv4
7iOTiOo0CS77HNQhrVfF0Y43h0kJDJF15Zjd4lejZGbXSbt5QH/GCWk7rKb03M/rFyBfCTL3+p4f
INVqyO3GFOwhrM1VsnW2woUvu3k5D8a+ivJ3OYwA2ezE/qJ5YtcqodCAWalBG40pJ5Fq+ZvIv5Dn
DrB9t858pkgp7//efGCdYh2/5Sdg+dOqRp48EXkxA0s8VgBPIYCQ5xCEgKuuaOizYZ5CAG5hmrYf
GyLiwZvJkqSHr8yHo3nhDpWdI+EUIoA/ucI387MOa6ApbrRe8u1DUxbAsU1+OGQn1xKlPuWryasY
DDQo80PllBFiFwFnYPUf4DNnej5aC2ZrJyudeOUdb2yW28WY+++AMXCZOFqLpGWuONMZ9+UmK5K1
u47XfqAzaNaLDVGvtne1IZtJZUQaE6N1vmHLazovrW8wspWrxLFuBtIBcCwLiDu/FNfVDlLwsWyn
y7fjLWPljr0M7N/EK0AwLNv+4UQfJWFvmTRdg04SRhf3vQosL2h17wH+Z2Y3gZsmDvJ7XuQQr0Ty
whwd3ii0hiaqSDc+LGnPii6kmzDhZHHF/2l2qwO8Y8J3Gx2EIRRItQSOUUUGNINGfFwi0CskYd6A
VBQTSAjT52Ir17nZVoiDTbbijOgMIe6ydZ3J//MkzjEXLB6DKOo00DZqqy7SAKjHryMp8rhklBp6
FdNkzFPSBxzAf1MEv73+zKLBLfliDwm8blG6wWClNTcGeWVhp4WHhDvBBfMiomoyMue9awqAXcEV
vegYTe7YBtR4Od3hfl4+rnQ85CIjEO5Nr5z15N8M2+N68zLtuaAxAmw+jwiDku6k09TSrFsrr0QA
idCOXs18Ige9c2eySYcObHWkPOrLgPS51dT/jP1uqDrCSzCYN2Hihl3d0yQ1ovU5wahXhpVNKkAG
rNaMz9CeCP+LtVhL3xtuzfAdBW8aOoyynGRGdwWiJcKfPBTUJmHhAQXzMs/Ux+oVGvRTo5Dwn1eW
J/imQFX3Nk2OfMclEJGlOxj7s2EZawZqo6M3XTBepQmfjqeXTqP3zVuQjDRtw+VX/VNRBk+hwMRW
3cKDcjO7QhEj99v3NAtXwdEh+bbqHS+ADVSq4JBsBeRqvgL2KnjeguqiA/bs2XeNdzCz10yLUmNH
PlYwZuyiHiQPgpOrw2cDl1nl2zHdioy7Mgqu0WhAHogg2Ivw02xfV1ZO2u1fIU8ObZsLs54lIWVi
YDfVUJhBujanc+dEaJLCr67sqCXxMEPoDB0zkZ/8kZmNi0J7x8Czh7Lt/xfY83te8kj85wWhCbba
8mjMJvrwgttV7gKVxFdCMk5pagO5sVcdoQGv4vr5TVEO6k6KDHnu6BxLKGZf6Uqu8NEACNK2pZmp
DYIcJ7usojyvK1QrrhCQfyOJi4HqrIxkSgfW/Yb/uJL1wX+8V2hrRJ3b3TeqQalZERR2imKK4WNf
Dj92WLM2gtSM7YmXXnc3654x5ni4/sPle4cWS6U3z678MZnPYqriRIYxRujoFWiIWsO8+HRysl9V
rQcuBxERc8076EhZ6my3YzOypyYRUR20cUv9n0e9MvWxJ1d7USXPX9SL6o0uOiIqSPoUiunUg6bI
sDCAvez7jf6yyjvMNkglQ6/e0m9gvFaW063xckJXndek/tayeIqKf/1yfTticZtcP8KYGVaI9ZlB
aK53o17a+eR0vhjDi3nQStFFPZ0+onK8apC6avV9hFYWNYxkDFpeWze2N4SnfGDBvn5Uf3/wi4DR
20IBrGxFFCc4NRp9Rf1QtPE6xkGHsdx4lK9YvMtSR0pD9k0yIQiPXFp9Z92UuAqw0tKhOnySnqPv
rCKnBanSsFoQwv9SE6JrgtTXnSL/elH1IHp3kXE2JW3Nt6PsNpBT7+pSSU/JauYE3fE+Qt2qEzOV
f0r0RV4jsRXJRGbZOVxwq0cuWF7IgC9U4k3B5xYLbSyz43Om7gnbIVrXYstTqu1n54fNUv+GFAJ6
rDEmgGenXuIApt+Dq273cgdg09YCEfKDEOmJHfStp9s1e0k2SxXH6o+MYlPElsf8kfdLBBYpXsz0
2qC0UQzlUJejLO9nk7pVvd/O9MnKcrfQ0prQpFQ42dV/R0Mb1QrDUc31JSPCbJ05IvQ/wq4QWxty
ZHH/08ZT3IYFX9yi/DV0FvuHaF0D5CKhFCO8g/ibXB6HRq8VN8JvqfUQH4bD+dRYaGJRSSg/B5cZ
YrFKeUifwRhAuCu0XjwS6njdPU4oH6nbALF7L4vrbF6bTLjp5+fxAy2W0QO8IzLv5I/x3e+ljjcS
vcyVik32Z/yeU4fv2lo9MAydU76tir2ZlPe3na6MDo0cxmGpklmT6uemBy4XEguUD0OjylWjyHOl
J/FHCQyHdsUuslNUIPwfcHvp/I8s6cvd487r8Jh1IdJrtDEHbYpFwgEsPGApy2QdNpUUedtTVX4W
3ZLPyjp7MDg5jNetlhZ6gymUHET1qlwR/ntbb/znJ/a055W5aDdMjUl60TwKaoHzrpU0bXyJjVDg
SkKo7cI3qlX6qHbOpaWnimOb7iZlLLxgo8YueHdOyputM3Dw2gLO0vPCY2UQ8a0CtnkIWdpMj8Wz
f5ojtLdAXp0I3i/ICVMretVNAsBzFUSWEiOf6F1OtqjzIvAW/a2Bbt1UM7I8QNLXic4aUK/1qgHd
6SAbi/E9WVxMLi2kWfVnpKQKOaPhTyUMrTrWGgeHvrHBjrYm3/D3JwXGgakOOD0MVoJYlVPE3nX7
s3nFFjacvjtWEkCWEK0fPFHT12XKywrbzrqypTKSJMr7K0xIRDJUDSE+KkTrnK7j47tx0ZXcrRIg
e8M4gNhVmWzhd9Jyjvot5fdXmS5Ze7XKduCQu/9xNvsnigvAmTOFD16C8Z/BT/m/6f4oDpBZF0Pa
MWUHtQqWk51KEEzSQfeYa6Pvc0dymoZB+6fdzS8Q7QAy3ETdIbON+ix1cfV6hThti7itZaHDng5P
mIIcwUOCMCO0CEtwDfB40+JhpRky4nZEBlWTVkUcFGvVqwe4JNQGdXpWNCpsroVIIW5+0W0x34Hy
xzaI6SCIfyhySzwg5MPTxeJgIDf8aoIpsOFN+S+rjl67EqHjXwzLMTjkEEfNtbPiiNK9g+RN4zgo
hfmnqw8nbq3jmDhmC0HQENyKobPrdaz9QXNTk3vrC8I05LSEQSIhgGQ3Nl8y5M+E9dP6UyG0eFT3
Y8mgljAIqLXerI9EomjBmDjwyNEyoD+YpuLa4U4PL5MFMX8osi3EiJul5+I0l/HCeZ50Dq9585Vq
dRxu2O2H3Z0PCoZ1ml2iF/+iEZFMvCo3bf+sgsuYSg78nwiTMp3uZkDt9VpNrNDcn7RJ7Q/UclP+
PChBYaXXpNrocRZBCwY6s7TKR9mbunRrt40kWkuYu2RaIaqxXDWPvrJ/ctFj+RBLYCFBqC61wjvx
D1y7i//uRq/hTOfTefpp2bty+72J0aOYLHiA2B8R+A+XugtTNyUagFDmVbaL4NH+1NKlTzCQI/YW
dS1rYOKw3fTlitFM+xdyMcvMwiQqDir/MroKkbrQvSTBLWFDuvYFvVfyDkdgljbnGRd2lu4iXftq
bNsp21atTuwGCYNSFNUkIggyx/3SRpFEOQdVZtWrpL0VR2Fx3sLsAR5Yh4iu59p/lGuSjlgMWNFn
lq0FAv/RLzVmOQnDLb4PzLhOBmKrVJs+4TnW63lukqJwwVKzbPeASRxem+WVUOIA6GWFVJVdGP0L
ThRmkYehP/LVZXTmfzWgIc8QUDF1610EmOV5yRbTWy0mi/i2PrKCrETxPLbj4w2JX8KMS5enJNj0
4sriZHlcmO4Zd9BU/5ai3hh1FqlsvwetRjX0sXA9JwUFqoHK9t334BpfHx5myXh4afsWbXkfFhTc
XcloFO+pYKfLDnQRZIy6QXNY+EOmq7YZ8rFMvDdtES/AkheA9SSY+O4fQfvEgqD7dr7yU0qC9lSN
kpnYdIaWLllmlXXZyq2bthgcXAHXydJ4tV6d+fK4f1MLHDGb1Ca5GqhildAkOqc9eCofXDM706kX
DHSvjZPFcNtnPv+U7Dh7mND0YX9ARaq5vcSEJubvV3UiSe5PK9ryscStlrcLqzLnK6v8MzqYi6B8
uBiVNwDqAhwBv4ps0HLSqrZqwkOK3PUxIuaiGY4P3hal5wjMMgohQaRF8EsP0t5LGl4eAClAEJ8b
7Oh4j91/u8GeSM00zp/xJ+5WRBhJDb0utlXDi1bov3JsxfJ7PZcbPsu965bRh++xHZ0lw5W7qF1R
A2OkVZISDvkRq/9sgI7MJ2rqx57yjaTN3XYJ4uktAkeNnLWllszgdzxpzkBPLs1MUnW3gq2IkgCD
XvXJE4QWIq7x8FuHUf/BOtqcKZ+oNmbjzeDZFS/XoskT8vPrefLlAEaPqO2mHx4K56yNzkf8bEwN
0J5Q1/HI4xSmSvTfav6/gRqhP68wW0Mji0seI5UGvuuSo4r6mWvQIDeoIm7l8BZoZJrkRIObBbN4
xLyyI/SEngqW1zRDa5qtUDBZczoQPXJ9z4fqnAOzOa+896xvdzD4NF50sgC7I6C6dcm32NS2hEJv
RdI77dVv1oyxH28thwgYVnnGX4w3r15TBCvFU8h/Zd9tZUMoAWFIW102u6Uor5EyxiwhKE7hQ0yD
wd5Nz0C9LJWr8zjmpoVFsIf4lGEAtyKGZusynY/uvbYPqq1r7CkZw9Sq6tNvkktEGI/MM3tvrn42
k2qzOw3LmcAJ9xE43FguJp4Avr0hKIaTxiSvUMnuDN8sFKNVqECjbZofH0V3DU3XxbxSmJG/Ubhl
5OG/gf0wjYCNrhsAFfT4XLEPeJx4VJUw6ra03DBcJ5fbq4T7boQjCyueRXCVSE9MucoDPM30DktC
TdStJ+GwkGn2gBpXhwsD00mOSRtLjMgnzYNhQm91VsPiJSDPcYeeePXgrREK9oD4K7Skzlpw4lah
K3+cPQaefkMfjFylMiIRDGfHbCJyAoAFa9lmpgL0OhRgN9/BQIDldct3Ouh8x/Cq77xA4p0ZHTFj
uYz002DBmpwEOfTO0uzehmwcHE8jIMZz2wpPZVBN5tKES0wfdyGGAm3gytIDHh3wWmLfkXSNeVg9
mXsb1f+GLpioPhXel69T5/gyyAZDXofze1jCb+2BHx1avsOIyMvgWr7GpSvP9fyV5VX/xKPzjKsc
LLPRjY/Zq6JU4g/EbJh80jJf4IxN8hPqSvTar/2LG2AY/kySkOmzmmjX1U1NX8cJe6GBAfPiyHSv
tAHMOgjP30TUb+i3zUu6/lZWLpeL0VF+XkT4GFFgRhjf47hg0XDnCPsY0ieSfgW+6T7JZL3VTB71
lopyvuRMkWdu+n1yJhZmIXP4KmkZs2O+uHlDIYs2SNCM+q09GpRGrAekT2JBHnnjxpZlD6UDEwf4
Up1pVz1qT4i24Ertuw1uLRd+2Zbn0o5DcwngEmsUItDNl9MdrfbZ6tW7Qq5ZXFGp8oX3NYP7EreU
zKiKF3wA86K7VlEGbpdCsg8kQ8UvLzRLWtsl/bpXjTQ46KtPReglfodCxew5hDwL5SBhTzvmpolY
lxcwoS8u8pnfaPkzVnMowe0GRjHsJXQ5cUUBVDwPDKk0mByaMRq0mDwxB5/j/0AV8mhKHL0Wa+kD
lzUGGnyM62qlukdptlCBqnGlfnX2C37cr+Wrr/4CxaBkq4fRJNIVA+91qPhNRGEFkBUfrB7+PIsA
+fI2aTxrGrQHbZqG6LoMvq5DxpG6U7dMxI5hz0fjUT0muYhwasv+wBXghULp88tWHf5bKnbp7NDg
g73OA7wH6Xt0I2iQkIj94UUzf4gkfsO9b+mIK4BI6i5j2Fu1H3McXyMLlSryyrTNFSLQccpFkWTw
7iyMra7msNYkyIsjV7q3WFXWs7phzcT3tcDwHca7+FjJpWPqqMEKryb0b1gy1DHdgvDeToeKc0I3
hHn3c5u+nsKxLFFJGPohJHUDE5SQ8ELe2F3Msv///j0ItiCGI2oK1VY61JrGFkJonpyIIDjeP04l
g/m/CUbnSm9RHcD4qPyDMaicZLYCPZpsq6ImUzanEik2KBm4wKBWUMuwN4lG5itjEXiTrT8jTZ15
Hqvlw3bBnNSlhp9zwGokcSLEM/rrHQC6JHMXXGXwcdGDc87TwXXJjimgKXFlhpb6qpoY+QbZtMrq
+Pr7HFJ7Kk5xOVDWLJVNMFa0ooRjvgRVbnDBeFe41JLdaeKIVxWzmrY22SgHdw+kQaLhbCCx+urs
zRO1tufgIj9ENQYAMPV9O3IPqk0obxICHxZsx7sNVRUE3XcjAEOlVO2CsGCCDWr3riImtQZjIM8N
PHNgth1mK7Uxwr88soInC6xaZhKPKae5C1/sOHX3Kdwc1eowfFG2UAG4PB1Y7002AHqqDvC4Lmb8
eXfjk4kEuhEKJ3qp6TPJbvfb4VRVSv5JfsuFSVr5LlGsUvR7nYIWK75oEgUh0mYSAZg83wnmgiK3
jc4kSp9h9SezGYnpoLY2kkiu+blQVVGArz+QhjEjyOpfFkkRb9J64qEmTmjoB8hR7HNVB5skp1DS
X3uItT3u/YPxhfe8Vpaquc2FrsvW3chFBEjQfu5cBbprt3BQxLiIgOjcQh/J1C8OJ/8JWsL/yRjA
Fje94qmMB35Z3ye+J3PtS110lC9K0TBZpajq3b9FYygXos6Ekort3PjHZuIG4d6ppvqBEGUH2dEO
sLHAby+JumOKIkgV/hCy22xJ3N2M55nVYQ6y3XtzXpV3PPNB2vXYTtaC3/VhDoMU4Ctua4DVgQVj
2K+pS2l9vXYa/lhrHAew0i9f2CZ4LqAJx+nz3AVlu8MDzaMFVcWYmsVsz1so5F/xMP2K/J52Mrt+
b9vjvl4H+iCaqu60w1Fda254ZSarXRwwn75qEEOCLWqPE3Q3W//vogNjLYzquqd3bJlRd9S0L9Qp
UOWWr9qZ7l9MZiAMk6srMhhJWkDqtpC3q3XYE1TLqhhZZaMwhcZPd6lgybcTCkYOWJJ4vBgxG1h+
7sro1yU7wSJrGI6/C9l7LgiCSCme9yzJTPrRcC1lxZLAuhiqZL2GJdKfirzNwt1Tu2WjKx/2WUxY
hF+VETU7+PjQ16lBJvSsAvSq2WThfpkw0UYCTPOn7q7I+/tbcOV/Z1TBPJxbqhwvHEfBPg5nX1U+
ynHQ/5M3fIXnch1VTxN3SCb64DQ7Bu+LF2vZhce9BKnO7lJjRJDjVtMOo9r3/QYVTUVefSRFpOp8
Y5L8lWzW0xILpF8J0m+I3qlMZAjDlrpO2ka6ArnwpjKa9SToeLxXQqWg+br5X2N1v9OkVmkn17nJ
OcE6HgqmaOMkzl4OB/vXVEbWGJFUsP5co/S2ZixXSs99m6sZFb5TQPoG//5pXZ55a3W7meZQYCOy
zQ5Aga8dsztFqRwJmw/v83iEfw1mZB1esWA5yAN0Fu+/sFwzM0QbPAJnPsMXVrMVqXPIRrUk7XJu
d5zUeqSBL9Z5DA6UY+1T60vF99hTCNa4RHClsCHiSO5mVKEoZJj4gHe+M7MMYGUzFhF2b+UFsHbg
PgBp4r1CFRXM6VkfnUBgLuuGVoKSNl1N3XRIVU6RRB6kkyQBRfuMHcEJWXNuRW/5RVxslCuguQwq
m3JKTqMnO+T5/MXOoXlzLcGYIQ3CVI60NlXQtEp+UAUET5sDA11XVDGwcaLgAe6eiQDsWm7hHgOn
kV3fgxPmvIUjnerfKnV1HXz/XCj8XheoQF3PmhSeNbRCjekPSjapZhBk+eORZDDJZe2sw5Asiy3n
e0RWJENZRD67dDbHxXIW+Ww8Z4VvrlKYWdRZ6vamcSSply8GGs5mlYCFRUHRzInXIig6cG4wNHBL
kPiPyTmo2DbZ4jrPH5ytjiwVzHOYpU3inxyT/e8NWg==
`pragma protect end_protected

// 
