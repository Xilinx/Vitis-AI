`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKheddr0WV7P2kxeqgiADYgV1YkXFGC3Pu48MKz38M4/PUTETzzD24v8Vuy
NiVyTPjeen8yjXdf8xepEQs2PzGiblTj3PQNiWW+sgDLOJNB7S0YM3nPNY6Ja5LTHHBmhbdChehP
OnGU8jzGLbiOgc16EAA4ObxwrPXDF9navpHS+/P2FZih8JOx/B7VeOcvAQoeE/Plm6NYwk/KPf4j
LQGC9hg64rpJ05luW2fijTuwbPkUzChIgFKXKR2v5BBpoBGibBvKyysUJbFI0qCqrnn68EuVbTgI
4bsMYTNEhp2MgSRTXr3zCWWZtKWAGXjSWSwmiHaJiefEqCWiNuV5mMDxnLPthwVjwnqLnSujFInz
q5SbOzpjlrU+iTetzfqJCbWJv5C71DTD9MDq9E7xUjzpIlOUk0lbFggca7ROAnoJxmlXyPj5T/9U
yzvYfpspMRINllHpnAAzDwpXIdWucAY5lg9wCrl5ZLO/rVW7W3wPd+BHD9TD4smx04a1xX/5owwV
wzEf04v2iVO2WyOjceBfkx4gCaBn+DNIMcnEqiKqiNpSm/TzcQpSC9xDTxImu4ijaX9g7so6gGPq
ZqzoxDVXZvGFxIsXqnerC/bglzp8SIHbnxvMHsA20xwgAgfphN15EdGeg/nBs19XSvPGe1gKd3qT
J4d41jSfq+D77vVCJByOHwdTX5vX1w79o5577HFmxAr17P5aO/w8yCTRGrQ1QTiiLIj63y4Vh4o9
zKfxXwDAJUhkHSahSFw6GJlj2M5avnXk5sEit8yJ8dOt9cyhPXkP4MqplB776HmPqt2KPUBJFrI2
1ujXtlbS6dBrfwc0q/PdRxlkVZG7/GZzs74vj9IGv0HiILsYdD85qPBQgtef5qgalh7opZsvxC/5
ZMHxPDQY1SLHX56uHGLtO6h4QSA4w4djRr3YkvgnOhkdXCCijiVEBt1erHMZoQjNBUviZFC+EZnG
6bUmL774eIZ1+dBZ7ZQzUDX9WPcgsyVuDwGSgHz2Tk4AOwAyIy6cEeP+auoMDc6lcwdEoeyZWET7
axMOCUETjx72WW9tLW9h52K31XpGzCAMFRDvc8mHcvhZxTRcdmmwd4cg8i2vWZ6IaMUMie7/e5Qz
gaCo6s4eDtWeAJRMwYqDx2IEjpJGzJfac9pDPCxshOsqJIa93jWAx6bwfF6gpp0jduZZMQwH1vss
It6sEJIrdQdfiGuA9NFGM6+kKZEoNeCHJeAjMa6TEbSCxvvQv9BAP2xzkbHLp/0oBVlJ9DI19Yq2
kTN2o9xyLKdxbWhUpgeZ2Wbv8h8ZMZrpjpumGCDHZw6JtesSBHzJyabjiDateb+8yX/J+940D80r
CgbW5w2rTuGCU4iwQHuaHgNWh1BxwVfaq70KS3DjR0YYdC5NRGUcbdqLwNonnhhPOOFYxqHPmXa1
vY+TL7dxYrsItp/LBdx1qRs0xofZv2rX+b+haHUiYLXP/CXMKwU/MkZv0eIxHQ9MAAXZgzzi3/t5
8EMJb/kth5G1jQj8FhRfcdC9+Pj5pzxYjuGJKwFiWBHhNQJKA9kvdE0XzrXlALCUYos6UxeNvzno
M34x/23Dpk7VlNbk22dOUOFv2HFPZMO0v4duXWTnsNr2LQsvq0iQOi3Wu11sZKSHHzHT6U56kz9s
lAEspcRXzjvtNgees0cyCEkapR8SkS8liuL33AHcCZ2OMQUXLoAaTyW6ujUUam977/PJkDpklr5P
7bDlX9pdjASdvt/vCw2BminFGyD8pq5cSIko4RmtPDOojxfdZCHDq05rhiH1xQMPZGTK3tywHbXo
mqb30bOmNPg60yS0YqiUjL+OgApxD/pTRVeHleXhnnDBMKswqTAz7Oh18GhO49j/rhEO1DkMTPSt
m+KytVk9UM3KcUTz4pplzwRrTD6cCDP/NVUWVD1vUnURUbMx+Ful0n0LatEyYO9+n1I3j+4ei+BR
QlicuhoOFPdf/a1CuFJAX1fsmDeNwNRCp19XUqvIOpg/aqXWKbID/ZzgXfCIILtXl3fzVPc8dWUu
Fzx0x3gsnaXmG9cMCShpi5tvebky7Bl8WNtxHfXf2/VNQpj0MAZULXtxP/fPSo493XEWZ3lHwqX0
warWfMsNRvaqbYL6jTqA2wLn7qQbTVpZrh9yZ4yBlHvrlUMIMxlxsVu7Wil4LltvG+SPkvPMvIOi
/8Mzpk+FYhsONVjbNiZsHEpoqtNlouulfE3MaL6rU4SXEC/1bJpB01GihPdTb+aHCxiM/zDVvswB
huXuQ7Qi6Vn37CensCOSr0nlOi7bEQ+u5EyAXMOr8MOv1psZQCvoO1I9xr1QWi7lB88O8jySIYYc
2/Pw1/BNbkLx2Szh/rRa+U5w0lOHAWJiZ9EX9gHKb31KdPYrzt+Z3tSLJ8sJm5saIsE54pFxe33U
7uPksLHq4nXcNHT0XWIGgVvXmMkz4CgGqnDecJLqLTJWrgdf5vLoRWl/AUaCe9eIV+mao4i0tYFu
k6G9ZiF4yo1WnLwf1rm7JAn3J89gF6CI24wcdYGKQTQ35dU+FgDbED5YW3eDKXznOFrlWWgbk/q0
Jqcuwm3Zcgi/RqoFqNVgvOxctyMbxZTXge2N5mdDO6qh/oyM+Z1ug+3v3okeIP0ZPASL59haCs9V
vXzZRBsjnpj1cevx/AP44Pb8zevWZkESsMghcQUWm/A328FrcKXkInN1p0f7ptxizpNrdGvmJr2S
lMw+V0AnMBff332NokqXhLZ+gZASLsLlY2t6vOLeu2Xg8U4HF0sn5P+UI0Cpvkl0HJUW+dPlBY5V
FZArl7UPlvtFU/zfKiwt7ISKUBjTfjtAirN+6PJc3wz/NBHYmjCJYF0fk284DnVEmqXlgbdWpq6L
7W5UJRThOsaioa+CNLa+hZnreoomEQNCSomPvBNnQf0YgqeIsHUkzwm31Vg3oZ6A/MMy+U8ILA9x
dKviQSoAxhAjWNVXFoB1pOK8+MGVDaN327kwsYJbRSEx2yQRaxi66knG2IgeRItLy4uY2/Fm27va
zp5XzKYlX9V87AzefIoI+NutAKNQ7yLbF2o3uP4UVby1yZp+3M/LWLv2bMsv02eYLL5qbTe8doeH
A1Xoeaggs/RUftq2dxRB5WcfJQ70TdWa8deZhPrDUNtEXNVGFDQfBBnMRl+cwV2t5J9Yq/+hiOaX
2Fws3i4DzYgRx5mGbRauO04s+y0TfLCiIYryj7d7bDrGSffiuskfyAiS5rAn7g61jH1ERJkc4kiL
QMhuwkull03F+GEZwHK0MTR8pd0Xb89nU3PPwvX/J3wt9N7a4g7fS1P/uZKAyf1V0anqewKklVD/
2zzXR1mwPHO9EcNWCT6/9tjLUm1zRV7GpFaz6X8jRqrFh5oevrTESfZErA4OD3/JNDWhJoJGZsU8
71HtmWQZ/BPczFVQ9c+0vgVC6CdJzEUW5K80motV1qnxce8Zb0GB07zTGkYBR+RxcHiYhvAm87Hj
NgCooxuuUPCf/q3XJeTCWH3cB+OLKVk7TbmGaeou8QiFcyOcTMTWGcpHKiy/Vu/7S/LNDhRlGyoS
53s6KOri+d7pscSbfR6qHspKn3vX5Uo3um4WVoQc2VLEclc9il9a2lkGvqLzpj0aljwHRIUcv/h1
yAhReq9Weff1zqfvjF/S0j0Fedhn/3/NnC4qxIeaBJBNq/0a8dkq3CW6EkGtegw88s8guBWh5RHd
0vq6c+kLbWPQN0gAtMs1VIl1h9pEZcbxgbCcKI0AIPwuWsBFUOMrohviRjZvU1UmCrN8OKPwsl+w
6onFzZbpM6PPCY/tmMS2ys5F92ZvW5Vy6H0qu3H5gdcbxqa4vxhD7t+hUBZUHTC7E3VmRuU+Vngd
So/G+LFjE1jI5bsL/EhSRh2YZHWSXMx///dJTcoHrRZLaXCCderHlFlZWFSty92L6kTo3XP6vy8U
xrbq6qkCKHVqfaU2MilStIAdVguXzbeQbJZuEazib4Y0FKdXJdFsS4iwSxlW4ALrOuQ149nepL62
zX0wT2tKeNIFsMh/z4aVbg9e/1AatrqWFc0ZDbvXOemgjNhnHBQ0xbPiNphelYEY7eduNsF4bQ3m
e4Emia9DOi1qV03SXcOdamb42kb5fBxfslDYLhoKfxCQMuy5RMG9A5oAPo0hZHhPiFotSAbRUSD4
UAY3kw0n5+N+HaGtC6wwzjnmyXB6KTKceNaYzHUS98GbLqFBo5yrQD07NbHIlNFLkpUebaltaVTC
sCBugTbNC4u8f3GYeFNqJOZN9ZqFfiG4lnDSOy5co/TWeY0CkTd86rosszN57m7bzi6nKgoancD9
deLZBQL7isBepPgDjpSRHRK3kl3x+KL6TPvHiSvVPJTGS9sypKVEMewIvjK3IwHuN5kl5BG9fPJZ
ey2Nawl8sOKxPqAvqGm+5JyGozu3O1gKYkp8Ke7ZA9jzGP2avKo5hR67lM2yezvjNs9p1K/yd16S
zDT6myj45Mj+p3NEzNKQygPxHugsD/ybNFblhjupO4Ns9PYk9fdIt5cDg/MZ9NOHLJH68kZsZ7XE
R5VPQHT0ZIQKyWwlkWHqGv+4C10Mu9jpsGXfNJYQogxP4UsNRqCV2SJIvA/H64bt9iSf1S8aPEfc
AkJQBBDHM3mN/Fpks16SBXracXqbjdPkogCGzU5vEdaZyydUF7PGM1nbQQDdCaI7OSyQNWG1xPGK
vqlGRqmUgx4L3xGX7Pm0VFu5HWfmDNEogK3UK8v2UMxtW4Eq4ZDtjaLsCucudropF/A+08DZxi/x
0aOcyp7MtXBAei5EW9HAxjs/AO92STDlHZ9S6mXCY/Rp/SCGqh0IKBhVFUiBbEWEybovBj7ljpFa
+mjpKAFFcOgMU2vbSDyYc9qw1bEGAXMuSDhfBkRUC2JWYbWFaqkxzeIWngvQg8faX5ctccnS+qtW
G66+e5yKLqouvTK169GGvMQh2SanOfBiHOLoc+6alu7sjhbi4ZZ6QnQP5ZMuO6CrrU6r9xUbZ8Us
XcN6iSMp5B7QNXrW3M80vRGJMjsAUMecGgQBJMuBgOaDFZfgKOltXaTUZNLKKdK31HPgEGLM9RBf
EUDZhchFHmQ37d3o1If2CNKzgnCmDeCLqYrclnEFM9JtgOoRKm+2dcZb0iAlREmRiivyyW0hhOYF
WEbZVbOde2qUVwNCZxhx0ih3WZQH7OgDp/apWFH0rCkqGQuuLVo8YPAbPUlkVcUxwV0V/CPa3CoA
S8PuKbe8E930altl6zR7pB2G4BTYR/bv/CYLcg7n9LH6+hzlOV0bS9reDXGaAeyQZopJwjWpGYMB
yexFpepeVT0iXEQSEDc8f9yj8phiMVoEpLj3MeN7cvoglo9QchC+r/F5/PKXhO21qlZHZQiGKFbZ
EAFGdRUNbuogNVWjl/o6Hc8fgjQ2/JcuIEAoPNJb/ki3jUpIzuJn3MsDWQ7dvDYSZf3e+CUUyocJ
30PNKboFb7h738QgoY1D3uemKCLc66eR6off19gD2sQbHOR8/RedNon1yPYCw+2Vrn1hdphJwHem
mt8SWV3hPrGhqvhwr8OMw9G7ajXPFNG2/pGoYAhD4hLx/IpkrBulIyFyPH5ZKwnWAFx3rMT5Kk7a
9BzmNR/nqGQ9jngz70eeADYQTlPixY3++fHphLY/0HzQMU6DqmqBmFodJPKkB9Srk0hxBQOz+IOJ
GuvZQIkyHY5iCGxi0ckDAylbODhzm5Ma1rSVCuUc3/nCxctJKnsNyZwPFQeY4I56BwfHckKO8Kjt
fiv2oVYdiY12WBtBCH6YD6OUR8ImuNpnFhebl5jo8IJo4BspfKxPPNrQrsDmTjMBjlc4vL8BL5k2
oEdHzjViUTBpmzxaWcY7RHTyEUj6y2a0IvxWvhw3C3GDdXptYlj8TY5Rgpa13jd1HAQYQbhmT3Xi
vNI+k5RCYtcgarxfYSGZXtJctHXhJGgX/+OtZkZ7p2xLisLp7p/StFGjABZfhVNB7tCWilMOdqOP
KwvzzpazHBmQde0KOJadf3MatI7TuQwOjzJnL8/WoXsWAzmgDX8t256xnisroOIYY8qBHuRqetHf
5XJsR2UbuzbMgrquvEHSWt9yEwq3+OKDDajDlNCChhvqqnrRyTx1NqCE6UoPGSUcEf5kw4Nau0TJ
WoNnHcNCVd7Ksd1dN2+vGlI8+hSe6UKrNpTMJvf3koRyo0wS7l7WYObvoSGtjlseX1tLoamzCKy8
GdJfk6pVg5S4u7giZY1t8t9iJsioT8HCrj7d9BgaewquDpXn6Y8FF1YqEqobouYI5nZvLi/OUu9S
ODamoG2t8bf8Gus4+NGMksG+MqBQp9PkopujcT2Y84Og1/uiQ7iJZ1knVWT0ptkdmaXZKuYqN+Gb
V17Rao3cO1rCWj8TWPFrgmgqceuwZ5j5GgMOgHSQYQ++5PQrBTeuTpMW1sXyZkcna59L2zoOLzsQ
d8tzSY6nppH0UUBGifyAIbuyjVCaM8v+yib6YxOE1JUY1Ab4e5IxylVIWB6ckznD4OAijP6MmVyj
8U9pREVerWCfETSDOr1RDbeSch6+KYhelegYJUxfHoGOxLJqzgylbKXdN0sgPeblR9jZ6OBcZ7UX
akyi9u5lkaj5qjYTFugnjAkQA/RIR2jgxxTe9aR4hqwTwPn/Erd3I/qywEkBe1Lq3z8ewIut2m8x
GaFQcx7sK3cJyj6p8DknmOxvSyXHgzsQcbjBDv36hjX4KvhXDTop2YuemLRPneL6cWA+l7cnexco
+VDvFFZLbvCfdXBKmoHJoHm7/Olc3lR5yQ0BwtD9zKjNicNDeWTAxsLEPamYW+SV01bw88Qlk8gv
yKBedtUm7ftImqOKJXpMB5kwnb1LnhJOwHycK6X+hKj7y3NB2ibWuvutCf0/eQJf3DoSuz6fL+RX
0Z4JEAF3faF6eMrbM0bxxmi9hDwF5//fxz7ky4ac8RRhacCSJZTURU3TEeBr7sJr2ga0W0lXbRpZ
SaptggzhybeKx2YeSsAkO8r39BL6KgE6F7cug+t2lRfghCq2EX7IhJpzbLS/TD6ZekqGCXwr2PKz
1QTZuZwpxajZofubHVYVSpR8IvN0PQXHUag00+ieQrX0nkK10xfJJd+WM6c6hlHMzuaD/36lMJiJ
CcbHHd//HM23ig26IRXUu9cwdfUVFfHKtjabOo13sJmPMgOQinjsm2vTZTogtNVfnyXY7T0/AJdf
Ul0LA8C8M02DHU+oFOMXIQBHo5OQlUtbidpnVM2Crp3ihFT2T+BzK03vstCJl6ZOnHnB3VUPU9Ji
czF2fXY++gXJMjYlUBPljLRrRwdPFcGd9WkoDMEbUy/7w+5WeqglKdFQWdBC4ib/+u+7SPjmhDlX
po5ifo6u9qnZUORfsLG2bqg28KdnPg+o9XvczPFQQeuTShkOSBq9D21bpClSO0aj+GsWaWLKsAZ2
pnvnLlhBkMz0mSmLuuEr5LaG7wGqrC/wZjFasyJo/l0Q4VjSxb6aVLwWZb1ZYh+hge4jpdQqlOC/
NpFcEKU=
`pragma protect end_protected
