/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2944)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAEqs/9I6SBGHpv++TEeHS/dhExIjL/29mq5EnZlN57b7du4NZJ/ROZSJ
C5W1BvgK+S1ObXIvOhPa1pzA2mUHOhXWxrU60bwfnmjaPXIlkwG4NSMrq6c35zfg8BBOa/LKQpCi
0UBOTb6Lo2Zs/JiCht0M5TcAK/SBcCWK4qxQkaJwPOTRXcQ4E2psfFAw32qkqBSJ3+ly0k3CM9iW
joZkUAAu8pml+mq6aBPL7MBl33Cj9KCCc7sL3NqLfuDWbeiYHlRcWQaRp9C1FM7iBfBE37BvltQR
hIpK9lmi+mSsVV10COA4XhhFKz7KsbkiBRoNcui20cC/qrrWmKAe3sT9YDQWx2wPy1x0iXLpBAJi
y4nB7bggkL/BNQZJavyNUi+mBO7nA6ErMi4aof6R6Q4ZmeeCoIt4JJxI0p4nfc6t7QZ8vEawGcCI
3I8JA3GI2lLpn+9l8xPmnAKvu0ZYyqyi8ZOFicuUZAtUXOrdJH2YRPO7Xzm0lHNP2T19zAnnG7SI
+YTecu36yl4JkGgsk2sZE2vFDMqCwCARy+vVC0RMDbR0V4gSsbKl5LJuqSUaBmimsKOKRF8sSeN/
TKd9pf1Fib157jnV+vBfO1PpUgmh5itEcfsQA7xhlK5pZ4hx5fxLj295xG/tRqP0jIR+TXtkNJY4
oZKAniowXQpxiRgZwZZ3RC2q8C4s5M0sl2VJaRi2Ac7p29POAYsf/a6tg6TecImfpDecQg5AExR2
75D/1KCOyJeGWdTcVMSouEALgMVOOujO+la4zX0Nihz3x8AM8+bHtRBshwnOHUll3Ra1e/bZCTnR
OTDjQ3kDXoXniTbTaiGIZ3uGdO0V+GRmnK67Kcemrf5359BTGhwnS5zM8jLgBoYvJkUi4O774Pg6
CotF4JIearQblPVxAK3Ii5o77yxNjPyxMfb/SOB3pzxa5wsmwC2IyqX8s15ezfm7fE5qM7mUViDb
HRTWTfE5nkPuNjMILX/3gcvQsEI6rxxJ5Ltg4ya4QD74Nz5wdu68JkjKLfkwQUdl2K+2d+iMz+jY
Nyg6uHhXoq5WQHHwh3EIVqMMqkOqsSS7btTGkZXJzYXXsqFee7RFG/3ccZCdfUkmsHeBahonOUwr
Hv4a+WOQnDud5x+urNhkJntvSx2LIUHVP5PLQb9/zLzQqwUYMwEjriIbsS9oFTDMn4Txu0tdgxNG
9SBPaWQkCPlHVafPEyD/29T+7tljJca+9PBNZ3XEALTmkpaPzdVdzP3dryeCVc4jJA050YKQzaG6
ffHLtCa6D593NBzdtG053KmAaYDmlZGVjEw7MLpQfvz8xTmVFvEdHpUcMMZtle2KYYx4Zo0mN9XE
BLWQ/VDjDLdesJ9txsCy0XjZDMQUbI6vR+osU7ZnzHRFFZguhsqhfS5LuoLSCQ03bp4v44wcViQK
3naY4odPSYSx1FdQmULX6hjeX/UduTqLc6Z1D/E8WNiuovDO1IBaGoqEm+S7kiz5Ea+nkMEjeqWF
pkcsFYxHX4miByrGSw/IvNRg+uZ/jJcVh5hD81Q46ju3YaZD9IAaFBwhPj2LZUf+4IBKx8K7w32H
3LHv4nCMkxsbbJ6skR8DKuletpAdUrJLRFoD45PkZux5kpBpwZKcgaq72ia/YU0gMTqbC/UdKhcq
amG8dcl1MMgwdB1XnvojK6L7c26g6PkTbSP2t/b4YidFXOvyoe5lHLWJmg/bSwx1G7gP7G0TZKMX
Za7tJkoJkPrrrlipoFLoVwaCZLclZ6R6tqVs+D6Jgv0TKijPhjgywwk/Y2vzvVmXqpGlHEXLceWa
Y6NiF9dCnFzD3HK6NXpe11If9ieA8v1RJT6dtiZwzF071CYVl6O+kCEziuWOT4hD4rCVyU8B6fHr
PjOT2tAI98nbkPri4bWAJuitEXu73BpEMK3+4iX/jmfwt1hWFqKUwDNsmYYoubxa9hg99R/6Dk3Q
y4bmcuN763gwGVNQ7nBM8/eUHGpKirB5ITmKWEUzwUv5uujEq2FKsJ8tP2NF2oQzXObRwzT0ZNjy
x/kecaNkR+t02qq7Z2s6dZW+CiTIXgI+Hw5BwpmywVpGlXS3gth6vX6hi+ifvb3mzFYZKxC3Uh7X
L5kCV9HodLxg416GobKJWRK9nwY6f1aQ879ne+5q3x9oj7KwV9aaEHY3anYZCZqfBPCw7/JhFMSU
aonYKTZsztHwKYmwdlB8maAaLFFYExROudfkWTIdoWxjHC02UvokJWYiHMeUldDNApqUVie71JY7
l7PSO44Xtp7Ye22nXGAw1EIkBH10IQIi4FFgxipq1WqdlN8aJu0jGqv7ztte1YH/BAgOFW4VxruV
LNS05hFWYZ4hQJyi4GnCLM2q+h4/D8MUSfUstqbdpcr98JeUyNsqnjNLdgLORZNH3pLoxvWHQQ0I
2vnvTufVMVsM+OjAKDyiFX14hYmiE3xxgYfa9FlCxAqa1C29C2H+Fl+ABdXWmkshABDgVFKptJAt
So3szkvEFhUd3TDzB1e4siQlrwgy4TPhm55cQgu+s7LYLwW0yf9npMNia81Gil1Qg55hZf/foP1K
PWbRnEb5+vwY21QDlS+QAoDh8KM5DyYw6vKCrthu8rMb3gBOU/ixl2cbmz78RFtje9Pmg+zgoAuL
azGslSpPMkG0EpTzJpelfMVN6cU/E5PVVp60U5Dkek6Gyprq+MmDdsQ3uAMnz0+5is2WZ1LOa/o5
pIYHzQaxeNxXtm3lwR+lfMOvlNKzPYA/1qQwtzTk3EWy6/tYuIDUuF05I5R/MjtrXmoPyun+xuBN
F1AGxdQkBVIdOUdkMYUk9E3ijy6vFIO1jfwPqxrDbpSL1THZ4fzrIgzaMdcG6pk8NIiynv4GCDL7
2prGwmV8LAwiVLi2cpFQcXqTgLQZ4kXj55gytIe9oX/rb/g7lQY2eCRRLms9JJg4nIwPNahODdNO
h4pmYbvl3LJ1g6sc+fuWCQdRF8R0HUbHU+FqDF3mCqZUJr8tJSCROl1Qdd5uw+mo0IP2Qggs7PVp
xaoFTcNvfp23qBURg9ixy4loqaECyscsJ3LWttvdGoMPXI5D0LMMe2XibgT3099cydvCcDWN+ZaP
rpoomMlGYHmLtznsPXqBPSFtqg2oD3AOTPYJ2vB1/cU519DvS+Y8c3WAX3kNIwRg5B4IZOo+rslb
mmWti1Lw7gaKEUsZyZi/Mf5JnBE09FqDUOqeljI324o5xv0NJAFMuQoEVVlkuijJHYMYMatwV/cu
WzcsuXP9WG9GKPNbCq3lZTc9VeWSDWb2zMJ0Ety0IMUMAQt+I6ns+VGSzJQUTY+u3XoVCnr285/4
Rvh7Q+vzd6fJlXAaDEDsCRvMyxX377WiMumfJHMFCnEOB7DQTa95LMd4vuN0tcntuWwox4l3yaCC
CcuKm8nXx0/WrvM7/pFlN+fkXT+sz9w82CmAZTm81PXKltSBbjmMacII0EzEOu+Ji4xrmB3yefXO
lhBY1NjZEkRhw4Ud/Bb1UjCUh1fS9PmBaCz02VT376u9JcCJgtZbWwY/K9K2q+vAuHceLPk9UdxN
znfis2O8nPweXNZY3Aeys4p8b5hIsC29OUSGQ558JOzTmQUYftZWy7bdEB/8KelSutu37Wjq5bB9
/rWCFT3mOBxEB3ekXh565bTM2lp1DBZ2AoYmRRSa6uw3Wd6G99LMrAC76NcYL9QzE0UsJUhma3Vj
15tp15zcT3PlBqqXKYEilpAJ8nO06YcLhLYHU15vZAx/yxouNJWWDd770A/J6U1i27FfvlZclmtg
BBx8if/1yhfCRjloBSUYv8No75xXdJTQunsyifGSpjmt9qw55YAM+dcidQ1anrRDm4PNSBIvfb5u
MVdirOwAAvTFjYm4w5rCitidsB37yCT356obKkz7PTtsrKjHaA==
`pragma protect end_protected

// 
