`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23024)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0INbis6m4LNo5fuoc/7VtaFb6U
0+5fXdMnwe75smPOBFJPEC7G1jJjzTejAYkTl7IUTkgZKL+qPo9QsJV8bWnGHQsxi3gvlQOIaFQc
GeHAIu5kCH4qdG/Rd7Opht+51SV6MCUG+Jzw6T7NCWSvcK1kUSxl+7AIlS+WIYISlJ+EKHtGVS9i
EwJnDml+BfWpTB9xPafHkbwEu3i47lW0rm65e8CJMpk2rTZCK9mOmdVwMqdaefo3r/+hw7Ca5b4h
GO7RZdxDr7GP2Z+EcrUoas/wlmYFktCwFO6F5IYzIeSTLltbWIALvXpEcIpEK2pndXosoqvAB265
qH/Lv8GiMDPvfw3MoWLM2bgMXMKaMevblL3WuepLSSIaWF1lnvE4I4vL6+dUS7tTpfWZmJQEwbOS
KpWHTCa3waxRAAe0EidZoUrUguhSsqaMz4NkJNlTKjH3pJAhZ/g4+a689dz85+TcC32F09L3opM9
Wy9zjTTAzqCcFhOOGIh4juGycMtvW0MSTWyRRzuzDW7buKVBJJpDr7qfH12Rv/lEsLY7D5lG8jlK
MExKGTSTmasBz00cAI0tEQTMlLLnm//PkraCwUb/mK12wy9omkU06oNqMcm/tAcVAjRj5jjFasjV
/Orj4QXqIMdDosmAGpTn2jgEJqZtqZ8EZy9QEsuHCpuH1VPp8GXrX1MfzzlF0BsHaS7SFVC6qAhh
tJoli0AhDAXHyyFPLFmJKHZvFVR1TqYpppzhalJhlih8I4AxX4uz2ycgjcmAhaxrojlRnMpDQh62
XWzLrwga20FS1q5vnPVSPKMKm7uwfGpj4rDQAiV6jp2daVYm1TIJyPdvtUVHrCgzkccxz0V+Aq4Q
EUPL0TKWj0OY8kmViD7VKTEamTTYjq9LQ6dnPE7Bzhq8+jR4rbOLxz9g5sIJdbTehWuE6Y9LXCoY
U27VdK0VhGASnA31U8ssS+bCni+mYFs8nc8VEIMdJS+Si8iMEKtrt4bF7SjaKHuVdYbQuZS1EXZJ
07YuWymWoaRfJocIz/AzJx1oc7D7kvBWDCw8xL3gE4j8QIimhurIMRFQWzSe2vmXknLQ/jzSBG6F
8/1z1y1hMekVC33vEZ9zBFAakZFDx+Vjo6TUn0x/5MxJcIiX/nIh9Ch1wsrtyUtEYZ+tfGGYmr4c
M2yuCMlGuP2/alLR71qLrSlCVHWs7J5TUQTJPxGxm0FnytF/tRQ4WfSqtMOxkf/rOOuYeXbLOF0N
2INRd+a575x3DS+FuTl99leiICuvn0pkx/S3/eWskHGK47fBkxSLYo+y2IKOyVxnlblthJ7eFdNV
+atUradytMnSBTLXIL0ZLh+DSqWAL+A6lPg/0f1TzR72O9mBEY3yjXZvMkQWzGJ8V0clfxslG36/
oCglvOQ5oYClgsoTFaAkAEEEJzchyHcPEYMJAiZZ7d27e91gXa5OxDmKll+4dIWDT26TLvAVAeuS
nOp+Y5LIa/Bl9eOTSH6GWk2qhTpcRlTh1/uOsjws4W2sn+eYQ3e/49k6U8dWxCSGRFYnkmvWm8DA
3sSOIs18/b9zUFMjkJj9wNF9Z1YFh2qXK8lsVZFjAxUsWLFcf0ohXEU+8YVkNNbXulnXrZK0AJ6d
vaHQKUYBw9gdqrpPm+2EIFEbAj9qa1UyvLGUHbIzfexk+mWrcsASp7p7x0AZM8ZQXPWGAuvZB0Tg
RcRgHXc6VnsXTxx5cFfQ3wWndozHuGoOFCkbWKHiPgv9rQsCE66y6fikfjLJKBmVrVvTfwwew/IL
3hF71CfDxdZn3RjwwdeSj19wPd/R6rvoojAi3zdDgilAD8jWn75cm+ywHxFpeu7FTkB4o8GMgMlu
phw/l/iNN2vap/s1EdyT2d/ZAtiShow7oilY1nuKmVHzstj9Lg4sckSIN+b6b7QSpNrLsDgFYumX
STI8B0I3qsnFcYVFRreuTUDSqVTfz9uMah6PLt+RTJiYx10NRGsnwf+5JPeN3gFz6OPpSvLRlWzN
d7RQriPkuSejzhJoHHN3YFcWd6DyxenlJnuW/PLbY/uXuHViCUl6yremdzkGj+ld1UaqlcorqVoL
0sakOhz7wdarcd5RIExslCgYfomN20SIr+exJWlsQvBTa8NBWzAZuCWdHJyK6BbzyRpm5GSx8xBZ
Ao7VjKzEqigtpBrk+BZi/L4kZx6yRPW8mNx9/YNKB4FDUqgbsVaTlcpKhTO0LEDorN/hSWnfed4a
5VVv07JJpXJm3Ysk0bsjpZbYg9u46V5He6j1Zr7+h7mtgavS2Fae82K30FcYnS8mt31yMOUYau+x
i1e9khKSvmprI3yFdnkOQJiER6zYUlkAn/E7uyz3LjWzU51Bbdk4tPt53Kmj2hT1RmZpyi43Pxfu
uprk83ywG/jX22+ep2TctAozN15oqsg1oTR5BsE+EMD6HPQeqGSL2YWCvQd30DChpgaTOwUMcNhe
jIfMgkQ5pBmFz+pJmnXGAh9F78PpEHO20eriNVUxJUErOel7c2eSCC3nqndu9ejjho9XEWutY/aJ
2SBHpFRQVl97WtUUBAHEUWaI+COpBomOMl8Yph6nOJAT/cRqnb35Gko0ff15Y+nS8uUdhqSbQmcy
LACz9FDUBxVw0uvTnJXYetxTT/j23CgK+7W6T2o7gfwBpouuitb1SxZs7K0ItsVFOEp1h9zIZswF
sOTalP5ZmNrUFEbXSYInCrgcJEyEdfWL8DP5SX/1ExlFjFXz0BrciY7fj/mC4lY3hwkDXUqBuDEK
P1m7QzasZWeXbmcZt2RhSuF3TUTb+75FZ7KD1Z0LOpnMJfx2wKwcJEX5Dv4fTkkHbx+HbvKqXEJz
nRZUsgRl8PQZ4rl1ZKQgAS0XXx7fmvTKQ4uggWLkiomFHXL6N5IRUstgx4KBlJXrnTUMrHozLXrY
meUve1qdCb1DGUx+UvgEAOSmiInf6ZhA+WVm9uuX3Bkt3p3X6+mx6bEFavWGQHkqONFbrM+Vgfuv
vewOOmA8AYC6ArcQmC+JqggWp1keyxWlP/zYHQPXvGzWzr4JiEhWc1mMc8HIhKYeIKLuGUMbKuHY
nJVlMKDfzFqaPNrr2nDQDBoqBvcQxcW8pbluCDtmVT/3UrvUDheDAK49Gt5FKcJeXPH8qbWYyRlq
56tjRT2o9BUJfAuyPc6mn5TgMM/BeXYZ3mY0TyjuPxdqNXZjnTcSSITXCuZFT5PGyozvwUFFx1H3
TbKt/xKIJrcubvtHi7Od8s2M5XgKQP/76KbJbqIEOzv0bqI+SNh5gD9RYTk9kT/dqvoQQv9dWb90
VqhsVJn28H+fsQLvSL9aH4yGkOCBcaZ2W3WenBTFlZfTHv6FWYbVOSFwvfdGk7TsdwqzIEzdHzOn
1ngRsASpDn4weRUg7/NDW9AT9tMRkt83CZOD3g5bj8Z577DeVLy37B9bf8wOuzXZznqMeB0ydZKH
RBrBg6iFgC5sdxjt/vmajqZ5SyW6BO9TKJthJRdqBpxI74lIO3LJwM/ZzhuHnBMAebfSkzm1i6Hw
qkvOasPSIef9m5uZh4TaBNJ6w/xuZrgbj2DnVM2+UHNVXyguHKxPQXElqfBRIj/Ei8a3kNz0PIXV
XruNkqECntFLQ9VfiYfwAF4NL7R00tru+YDKthz+nzG45sdJrXWhph132JRirX7t8mrGzRqfJv9M
W7MqvtXs3MpBTfoZxi8Sewcj1KuTQrQp4c/WrVFMZ7Z5MotlVxH0S1DIC7e5QstENH947w8FJgaw
iYLgrYUan65PjaslTip6uCWSxKJxH8XGnwqlFeGMrhlqzy7wEBoP8HaF0lKfps/5Pv8nyXy4Ohtw
XndWZcN+50XKH9VwVBzwPj1GcdMlfM0Em+CxOfkQiLTbcmx+yQaBrjCYjad4T7QKTJFppnZlhsO6
+eT3na7E7ri0U8kmXisHnbLXPzpST8pqzHZkn0+graIMHXdKOVDRRSTGSziM9RVDltWQmkmwI1oM
jdBHNvDRSTIGp7itxbB9VLJsPNieFQ4PhMRtW6zJZmmMNKpYI1PlnQzQQoLR+vTSv0pNEy5v+CZp
ZAGjKVQ6yntuxwm9ZdrJUe6pAewExVYyUsSS1fV5d2LZQY+f45mx4fjU4MFJmrQAbvDFQzeQCVCx
eBxGVYX7grRqenY3pl0YPhXw4V+SWiuSii09ZuOlIGvfoqbMD33VIfG6jELWhHkQhPC3WNopr/VE
aRpdNiTi5JGTROdya0UDxMwZHwK12kFQKOdVl83cc2S62K2IXoXucI4LOk8I/D+grR6F7tvD6eO/
OpWFZ4rD4GQ8Qn57VMZHE6eFgxGooENW60OkoL0KZvl0q1oqe+COqSqeIxueE8we3xsYyQNyI6CK
XRo6XErgF9YCscdb0kqc73dmlgfxXa5OuvIuygx/48VKVczfuytn9+eHJkqRr2pXnS3ZMZ5pdQW6
B/XE1ShVfGLFCCbeGAsr9qqp/nPpmanHiRSnbIRR0PynaSPs+2wb8Y1pFlXgk3piZ5Xc4GnAvCgt
wKQo57TU1laR+2hpKfeoWI/bGdrtQTI9J7U8sHxpxh3BiP678pUTiLBGFSPnEJIyPsOnJ/KmZNXo
KCnjOb+qvbBJLjx5wuOf4UDqIp42ypIOqxvfomO9DlTuZlwGfFhf3A64ko1kbn1YG6/JsVwS0okf
PqOQaThUHLrenDzZr5Utsaj/rbG+tPJUclTkNxTJl1inVvSKZGnCHHcMeS3vhstOwudP+DEyHkan
HZjhEHE6jN0zx3LtJIR21FaIhF2kCDEoYurz+Xunq6tUoXHC0wG1e1tRow5eLzeKu6UE0HW09e0X
IMdVdqyFBFDWUoc7igHX/321rlPsErlkhL/EI8bDqHdjIsfzRLa2bcPi+ZkB+mrwVrku0SH7nNfz
zkZGrrdCzVI3/3a9kf4aiOSoiR5wW288bd9jDQFgO8Sl0JpKOaPff2tPwr3yWwAFZlG+UNUI0R5h
Ca1MwTxyxfkp7HNQgcV83w+BNgJmrGc/LcG1VQIzd5PkPyQyzdQxyDh7CtzB+kYmH8P7VF5wXel8
hh/VjbKBREzCoEBdVuiW5cMeBjDoiuEU0sB4CDE3bKfX4GfukfAFxZkzZPiGs7ZPq620UQd906S6
XBYE3/bZXa7uYUqN1kg10Y7ijTeECZ928r9nwJbMApsUQ+PaWExnEDDH2IWn+dK+VjLN3VIbzFlm
I/txEdS+PIi9NMJyh7Ux6gjvR40vHsIOhgg69E4ARFJ+zoiFLroLHtGZSRKc7FF2RGv06IhulQPT
TV+05nr99w6N5WvaqGsfLpLUJD093Eah86o+AgUwWe4/8RvJmuiRRMEFVrHfAzLt4kvVKPRPYRWm
YGQR97LCIXCVGgUTErV813VYh7/zVRhyoOlr5qxgWmwYV5RKSh2BqGZOVui1prYQVcz3YRhN/myI
c7OojEgV6pE5KUH4uYuQx0EwKtE18oDqUlcB0prMCFFjjraaGfTlGYVnXR/CjHL+ccht9wRzw/kj
SC3QEyQuKnsvj69+Jz86YMxwugNhdSear9AGuss3+FQ1tQ33U7cpll//7Jf7blN9rAZfwlAvu1CT
H5dMMn9RIRUnA0bjT4yQzRdOM1LGcFsYgpGVQi/I6sa/Hg2nKIghJlCB10O2UFUnZQCBqViHfX4m
emiXvM6Ra4Vpe0jJDaKJSMih5mDGQGQwTLW/Cp1R5uvphZlkDwcsj2v4LEdlFqwSWpv0TzfJ56xU
NqWpX9ombRkDnVhZQ4DZ5uGPXOicCG1y33aR1URHel0CSxMl6lwFzcK/3Y9uOVXZ92CQy8kTy5NH
2wH9J+Gj6MEUwmSZ4kfDpXKbwGQHXvPlbwqvPnOhJTOmu4nRVSiebrmBJ9CCMsUIRWlIQ5RUbU0v
sGR+WY8ylihSibn6vQJV5zmQw3eE7R91JfU6xk/2zMyDOvqGc14pYd3hmM5VV4y9pLtQocmmeTHZ
QSTEGpNL75AF87zrb4faAVkJcUHil3v85aeswWo+ldWG7Zozo3K9HsNJ7UGb7jsHxSJQSgtc7M2Q
aIM03bPm83si9T5e8t7JG9wdU7ofdVrhQ5kIeHOGNWXzGIwls4nspmh9wvRnwPQNvgbxBBI7hFfU
a1Gk74r+TahMiejSY0NB5HGJQV0DBLpj0Czk/JEoQonthNGpL2yuWNBqbu3dTeATh7AHZ5YBlbRT
evK4ZryCX2EmuwKE534i2cPoo+UkhzoC2DcG89LmoquXznEcuDm1zmAuHjilLikZQI6sh6fBJjq3
I4E/ki8oTqc7dstOlvtQecah9flY5EiohHjaB3vftlyx4atp1Pqjw0EfrPUhvM3DyysD+0Q4TUvx
GAvYGQfLxs1Paxqh8g/DqQo0hezcyOFIL6l/TkpAbnXb1S2jFGAT+knJVslPoACmr41mG917y4J3
Xtv8d6FqX/ybjOOLf4lKdvgZvP5xlotQrCn5Jy/d6cUKCSg6a7+LkQsew5n+Fwn3foA3W4D1PUpW
f6EW2nkg6/XCmMO1IOksk4tPzvb/AmMLOLJ87LV15hVJ1HFv1ByX9Nyuubljy6mw4rqKw6M1GfDG
WVmGT7jfr8Wb7cBPg4nXDTibas82RQ0Ugc2vhxC6+8PV9zsqbu+q96hsRYbmEJHHJWLoZJZ+76Kj
7b+4TgdFpZu7x8L0NQ64n6LHOHCXnCqdqHRblAFmWAdzd65wvGKA2R2un/spgDWOOnX26lyw6Wu6
SsLLQ6E3XEyEmpmKGkRcrozFp7XjskYXee0q75r+nyWYAyZqsgiLQa22QCGcEJJ0Ezfb8IueqKNd
8rklCkvjkCbOlCmJGiiGsQxtbf4uw6Umyi8s5uWHivWgUVaS3B3jKRVUW53Vrqnj15elCkUDLRkN
4lFXHGSFMroHIFhPpxGcIbTgh0IvkiYhLGjlOMvqBWH7tjcKZf9JJKVwSilUUzoJyKh8Dzo+yQBF
n6xi+XxWSzIWRwK+o3cYoQzi8tTggRYcJ4mYyXpE8wBOJj2Akm0K1K2wQ92cWqokDci7UF9QBjgq
82M1xk9VQhzKahR0EvrluElWu7oRsuZr9i+F9g78YUSTtOGY9t0NLGj9kUxkXoCSyfMlsaw468G/
b01oQ9Tn3lItf/e1KJLdkE/uEr2WFVlAjcUTDMBp86dusRYzJVLlzFbGw/i1cNf7wzLN68WRZde4
SOgMBjiChuYqN963h1YWwnNV8VRAGT7iVnEC7M1+VrMWf3H70pUBRadtRxf9gtGN6j6U8afL/phn
IRhRpRTcGG9oy5I+nLjRClIJ6+WTBimNj2u3elAVujUque0C3/swdejhpgsil5uo0QNWOTRpSPse
cYl5KzqMQKGooF6ZcuXKUfAgFUoWybX7YUYyiZS7vvxdUHmPmBEtUp5OmjuSkM0Wu+wvDzjnBPtx
wGSLB17+HFmlupxZeAKEZ2QDts88dYJqSu+mDTDToKUAQM8Zf7vdNsisDuhlijiQHlaaQ/x8IiJO
WLHaprLLoKoMt6fADgXdjKbpNzJwCk3zKJOx4UuFvd2DFrERT7wmiIL44umPAz4reeyF8IIuad7x
dkXzStnX7wjAKPLnNITebwMkl6fYo256ZYnm7Ioi/s5M/G8oQMYRAi7qfN6ezkEci5dnKBvQy69o
SNo54q668MK8yhcNf6o+yWf2WzOvjHprUO1wyF3hHYO+pE0M1tS7nes0wI3BiaYUFjE1Y0RnL0Gi
pphAtTU+3BUViGTVuGJPVLTSWt7UmNqimiAYN4/iXCKqxHUYlBucgkxkTu+fU2luEvouDBBJO58w
xAIPDIeuEMkTRhzxsGRT8DM71ejd0MIVXOLy0V9o5m/aaP5+ek8qc5aTaW7k8xbOEmKjN4TpkFw+
e9lLZtJGG5Uuigxzd6BgD/Df5CzPNLuMXHntePdWZEhIuoFsgC9JdcMXBuRrqUmZ8zhti10EFLtA
0r8zBFVgUPrOgICgQuYcTjvs9on0JRuGJ1UHoy/2A8aBj2T+/Xd5YbvfJuUmL4rlytSck2G6epe1
LfhjVf6r2/5cro+dnEQe5ukw5HkRWy3pUQrtB9LBd1XamDP7caoJvSM13A4nayOyvq7TcnCrZ16H
Tf8bFEp9oreYSE/fCWmGVLe1KZ1rU+pSPDhj3pZ7ai5wptMtDqG+TJ+J+6qlyilJBiPcZayXctE5
XOsq8V6SlK8BqsFoHV68/mIHTXVKl9mzIOyIYrphJf/JAgQIfEKJGv3F7O/ix/ZJzlyUUHfnZ6PK
8smPHvw0Z5bjlDf6Me/orCMsRgzfKC8c9N19y87oGennj/mpdDiv86uCQhszJqELYaBFHlV4VrY2
ACox9QOjh9Zj63bxvNKEeEvql46JmddhxHC41W8+SiDzoqzZ6qWneEu6C3O+fZYMXVuSEmNMTDFF
DkpKif7VPUM6cCR5veE/krrJm72njQd7lEnEZRWzFuim8SDfj9fu7xqqxgeHoxYmWpch5EzgufGb
+6rrfS2aB61NDl2zcIiRfaIBE13MKrs5qzHJRNcGzQOLn/+fC3GXNsDSH735wPIjcB+oBhheSkjF
k9FOaKxy69tg2E5ZjB7CUOAezSewk6CJ9HXmCNjDDYOwRPjRbIP5UkWUAqpPtHmfG/LmOIVPyOkj
1lVahkkph3a6DhcHdRWk3cU3xlHexvIIQaxdVL8vIaLt17+2zDRS2rxmx384CqCb+cosb/dWzFL8
EIMwLIK7G1+MybT56ZnM9Fqpoz0ELnpwxfE5WlHIN1eNtFOlAk9vjcK8D8lkl5cYIq2HxGVAhpUK
Ik/F2cqEVFKtztYJC83eoVaYDPNECPhbAjBpsWUDKAsIURp6yE+MH3QOR8Cnm2PmEadst002W3Zj
KVPhHF7qyXnUEbj2dEbF5C/BqKre7UR/+qmEIDMyBV8wogfV+Sijj5skI7dYm7rDy3HL2OzQioX2
p3xSvBgYtau7u8FnCnzYu1QDoPa/vZV0hzCQ3bx/EwPLICPweiFROJCKH4OpeHRZWj4yX8vzyKpo
Q5jX956SdNs438nMVp7tDcrncL3SybbHpDTRi4IzQlftWcXfjQ/1lGGnqlPbsi/NhgGYEEP96daq
KGmbgQ3CAaXmOcMjp85s5xtMzb1rZ3P1tJgLnDdxctB2NqKX4qh38N3jXgXSvbFNhxkocp+a0d3r
1Q6IcDaUsuUROmVIw6If9E1I1i+SV0flXPLsDEa5pMVnVmeCs3bCPdVSVOLQTPQtxPA5MALZd7p3
n3sqN5XGU4nqVHOzDJ0gMFTaCiJTYkbEo5F/EzTew3mCrSqCsNAv1XINtWRkfhSWgAe1QzhN92TO
XHG3te3GQL7MdsGGAmsCOvBImwLgvRE7+qPu+3sNNLVOdqMfVhhKtL7goiyKpI9os+BqYFUvLfgx
+XK16sSx48k98XEGrFcRI+LsKcT3MEmEHPH3w9EeXImZqltmFqIxNQhkB4puVknU33HRoCrTaYRO
BhbttCx56Tt6cuxOjgy2eSXh/MU9R/QIkJrTqya6pbx0rZPZFQVt4PvQfUrAIm3nKGM8+iAFJVcq
M9NJR685vwz+zEFC8zACeRQ40DaozvxEIqm0tYv8KvnmIsSYQAN05QlWtTSh1E7eWpr5N2YXdnck
ku4vnehRet6S9TEhpIKQr+Ri8ZN0RUeZQTKA+yVIUljwp/8esznN7otS9XdekMFcUooDdJiFbgZC
MvvtjSptkP+rwTRJaZaM0+gDYGNYGrPQifAZEYk2g1TwxxFy9Fj3yWUhntNQReFZeEZPFC3FKc8q
pxezrAz1NbPM0o3e864ySD/z0iU9jchNIdzjbiD+gvF3gLjGZVHX/Hx2/6GGD6/bEUaS1uiLD86b
cKnckNPYrduGTtTVrkWe10MQWeEN3OU+phcIVjr3T6ACb65cNFh/f1GKvjHVdXtSme+LDPmABysz
zh+8TlV3NsozvjDUaGrKqprD7zebUljwsq6TBjRRISYgvZzi4PDy/zegJv1hLwqniike9xmJWQNU
8zMP88Bz3PdQsczYo04qmXvQMYVeDXMQdfoXZxRPEq4s1pnXQJnGG0hD8FDhL3z32ONalG5uc72t
o2L57l6MQbu+QjrTYgfthBv2f27chB6/SYjXulmpWCPkEyFJkxtQ5XuoWCzFKcqzEH3APsR/lMnI
jkAviRH2dqo8U37bl6M7biXbWlZDOT1jlNZGGj9/rssbuvRx8UhFNMq7BtYPe4Ai19sSzsQTekbz
/PDE/a2+UsDh0BpnyoWpSnFF/u+TTKTV8fZrxlBl5YTf+DIf0AtALnQ+dGcRgQrK4PmztTLoDWRy
heDMeG/iBmD4V+l5RZZcIFWaRcYukLcCm0AwwaiQ1q/t6bqTluI15mTA4GElL+VvFXjiQ1V/Dtho
ndtLzrtBc6vtiRX6gfFzmJBarsY1Fke2mmr2PXb8kuSucUk1BybE5nASw1OQCxkPCbbD73TW4/pH
zjl5KnKBzV6bFIkZITAm6jJBmrSKrkn/5sU18tqIL2F5aiWZixSTYmCbySwPp2nj+9O/3FA5xPnP
atFQcLdZYa/YZfHPfAfJ7zh9KQp5+NPqiz4RvIypPWOlH0vR4iY/d3a21gHcO5Hi3bCkNsA416d/
dbk4FCivkWSs6iQqYvSqGkFkVQN1zQuTaAQq23e2u9gYctHmPv2kNF1cKNBRHxR93zGwV9tV0FSu
QP3Zt8ymyso6no9fF1jVoe5Dm2OOzGPUxT0ajKDHkWNVRzEDu5waZ6mmdfUQOCahi3PRDM88gEoR
L6Tb+y4nw65XancJcdCRaO4uG7svZKE/83ASla8lRFOxjSkdqFxmpvcR47ZT6RyqUVlR2LNLrYTd
wdLW6BLKbVK1ifkrPfhJtNznX+E7Ze2TxvUST+W/N4edlRwKi5vgaxzBpJGx7u58Rm6YLCd0W5Ul
fvactRO5pLzhyP0Yp6UM7gX477nxG7IXHNjFRMyKWPve5npOiofBIuag7229QXNvxkAfSnq3HhiO
n1+5Yzp49x0eQqNp8w0bGawxgpuUjD5XyNKh5/tJ3/EWFq32XITGo85Wsp+WihwaFyI8oq4PDr96
DOx0czbMtyMMggeqAtVXj5b4wNYz6q/48zyYtZALq30Tw3AmNIUsyDYCKaAzr4aiwbwvRFnF+2Rh
6yjPQ33fiz0/nELhM9SMoKDv24f8DIH0211exYyM2ZPOs0SgBcNofD1K87Z5hacYcem2Lr6dyHq3
OVdkvqhSIVPS1EMiXEYi8++dA5vW0qpZ0ZQIIups2uZXEaq08Y1SCBLJcKNZBunlL49XOh4/4ip2
uSpQRX+lCYIJgSmEsgM2goLyt9vjrNVLSh2x6kabE/Fnbj2ja8AXih4fVdDfsZP2HULYMjNbMD1L
kU2dgwBD9/w9buTeAr/NnKVWiWLxA+uOs+4sltFdQMwCupPgZhoH4EZLFhXgHk0X3TOdHraGcLWu
CBotAh4TfFKoiYXABKColMXKWg2l4ZlyIWt/R6h+lLWUpwD7mL1eSzqnepiJEX5yu8geAAt/B8Qr
SNAsi8sCt5Fg6xU+IN0ob/dkjtV9BdxKeoTOAag4RLUXVoCh+fMBlhOSWcwUAWrUnG4y8kcXxPEs
rMKQA3Yu4xY1Tr9xzPLHVUVZ79sxWqkCxvMbfs1YotNxNpj9MJm520WjrNqCLjwLT8n87GTRAd6O
QKXQisX7DQ4x5w/hp1/eTi9d9XbJVE/eQV/mrJ071uaVmDMKQPzYQFWsNSRP82soZFlIdVLfZfHM
r2s6odE0zZ89cvexm/OgPceq3CTfDDTc37Irrm94f/WwwbeYsLZX9ocJs+Iw/gC/vlc64i4fR7fF
XM5ZsG0rHH8P6OxGE/aNH+bYAdEolkF2uTsCm6EVNhl8mXCG5ir/GcllHqWgT6qijSflYEZVeslQ
YRDEIDqvEfGSjUh09mBcTohG/XzMkG6bfmq3irmcXBYaX96GtmUXkI5T33W8vebTDdwDuX7geAAt
ADF3d3SDNcevv3CkiUAnQLo4yf2IbEd8jsBqcuVtxUt76yKisZXnjqcF6sf0/STU3hbOjWK2PuGz
aMwtHBJqVvvdzApKv6q8ZGravM2ujU3jHJum7nc7Fi6xx4PWzxWVpY6lvlZdrMTk4jDMWC0rLoHm
WnnXT1LYbnX4ZxQTfKjHXS52B18ms2aY2opwCniEwvI/HpWql9Oe7D1FKh8Kkc9ff0JyutQfjL0e
r23nTVp9pTvGkBtMaJKmw8iBs6loWmGOGsrcG5UI8nIekUGnSm4q2SSxcNDRXtyzrKX0WJCKT8H0
b94gTPg3MeRxzoffKGTHkIZReIM94/g64xZEosn1kxvcwFzrWFRDbbqesqjpRKEputxIa5DCMBTn
+/vPwnfV4ifY9FJ+Jl31QHVvUltch3OtV8/h3KdZt779e275Zuy9yr0PQuXxpqOS+mtstdTmuwXa
eI6qnX9o4QWENdqAY2qQ18tg/U5jmgoOHEFf0jzcpUQO0ihazCG30OmAp+JsAfBN2BuqsR0w1Hl1
JahZVK6t2G9HqNp30XATgZy7+H+8Cl5Hzjs93n1tXkqlWYcfFYHXmmq0WTr4qXVCMfdCx8z2af7e
360fRzUJDtrrwbkpOXFUhrB9tyCpXJXdjI+IbAu00vW75C12kiy1RI5r2HJ8X8EWoB53GU4SaHb3
4KpN+HjW64nvpNRbIXiOaHUCMWjTAT8V+epJTDg6u7uj6blangXlFxK9if77oFEColjAEj5DmQha
TBnklfPlb0RNyn+ARYxZRDM/lJkntTF6BG10De+v0tbHDGTzZkdQfBtWMt2P74XC9hdrykqYxKd2
ZYeRWad18Wnzu+K+otCQxmxgBPYgEp36dx+W5p8B6Ix4fIMFg4mi3jFbf+wCMexSkiy+LT5SeJ8X
HpSoVAZOa0ejvWRQfPAr9lguoVAqr2N911lYa9Pc6yFamdQXhPBrcyjAfuz/hqsZocYwMNBgbYWH
mLxByu+UeYrs1CXvWuLrKekFF0lap/dPLek1d7V/6BUZeSjQWfJFbwvWk+FWhzMs7Vf4pg5+1G5C
NF034+7P1QYOiiVud0kmxo+m7KyGkawmQs/GpvKclvrM62dNy8qemDIcG0aSiBTqPk0cO0RJE4DN
zMuGEda9tCMgir/HVi7Bvxzw7RzVcOVcitUG5EfvKKYcN2rJqc6+pGO7PSo/qeGnEbIdDWjSBQap
W+o5UzWOgFSfeXP+tQSiV0VVExwrB6cm5GSmpXpkgY+4Oqyreo3Jem96OB6/Q9KvSW/eE3hPgL8N
ZUEJIb8/Ls64AmLMW30O6lLoYzKfEXFDd+ag/4Cwb1Wwu9qYdSdLhefg2wk2zWVCenXHancckIga
WUJKcUaxqWrhX+iNGd09zRoY9CJuIOE1csn/Tne0HSBmoi/CR+u7GQ9UuiULAQzERbcSVISgKg64
Wfh9OqkHRFebl48WKmYlelJyy+kM3tynBLcqwRHdumJvBdiHG6ccwUjnvvCSotc6EPJEpPUJ29in
QujXb2ZPJPaBdt4+FWat0fcLavidjEk5jDm0s6qc9j2BbqyrOWdVxGI59312TlEscCqPYxtKKYtg
q1HZlzI8mXkV8mhDTK9eQbLFsIyaMnHAg+MiYkbW/LXj1BXaRUeEWJTaWDNehhM680Miil8BkYvz
8Ljxjf+7i0ThjOcNpH+olAuPFsfDQu5CsihL0GSteMiF1dY14UvcovKoziGGt93nRmZfHrduvoIT
T6oMx+nc/YSawtIrBIZmBLcAKqYB91UXQlACN7ph0I+LA61yG2ed5eLAa4hXlL5pgKw4XjPaRhxb
Mk6jq2yQXxbqLS3TsCgLXZRpoJy4eNcY0SYJAIYpHwlTq96Fovcog9fP1kOAEl4Kovkk/+OZaUnj
AV29pBXdbCLCGJdqrhuEWDQEcFdeWj+WOVa/EutEpDhVXrQh0giNogJbaY5faWpMTmxC8Xix/mBz
XZ7WF3a3quEfCO1iUGpw1TFX2iDUWwzAUm1d6mdpPhkULYyJ+vPE2rb4Pz1+h4hHG4tfunDtjeHg
wg6YzQFFBIbUZqN4saByFdnexi0xk7ui3PqdrLsRZ7HFXHW7ZZUml9Nghl6CU/M0Jt0of7EYCxVD
oj8YCdTfUFHU0yrNN47cYY4Bd5ZxpuiBR/Op21f/FK0xs0+qWr9u5V55QaSiDrDUC/77gTDKGCGR
frlMdoZM/CuL+vmAIP61+CHSmkbUykY9ZkVoiPf8KrFHXi6N5UxMV4xfvkfSPVvQSlecU3sYa/4F
pX+KOYTxYQ5lBDG8REhkTYTfSh2RLPI1OIfoQ4uInDfXgz4cEfXdRd8kY6BSewd9KFMNgUWleAbB
H+x5q5FVUjBwrV919h3KVitO+lLmMFuaggvc3+TxMw6nOdzmsPdQZzs3c29Z8YCFwe2khnCLdX0z
jh2YpGQauzCCwqxghI9xqNyv+3CNwfiS42oU4L8BZ+ELUizqmHr1oQb3CdLWOYPggqXT2YyYeV4x
hjcsdRSHaiB4EgXNEdhbeE+gy5jFmNa6+8H5t609NI38iS+17mvoG1OWE06lYGhROOSyOW8KfxOg
nEJFWUnnHnna74eXymmsHxAsebU/+yFo/hn20gTJFL+AIK8s/PxkP0oTthtrEJEXdCdnF60UyJ1l
+2IpOTLMGDSCswxRihtw8H9nSk9dIiJacwDoCxK/HTr2nSfdll/24iJ0UO9lQfS1c+hCE2C1zq9B
ob/K9n5tNDgS3Jz4IxOPvPm4xunq/W545NaBTak2Nh1CfM4CRqmGxyU7VGyWrlWw/YABBkiQBZ+F
VQDMDBfUE2z5HTm0JAHEwk24yxOw7JlYKAM3vQXM9NH6IjrWI+++Kf+yYgjZlu96LznI2NtKZIYZ
obXWseK30BWG1Is7FtuWuSSIp2KbgZmaShbdtw69rtgb7aZkD8pOetA5Kg0oRdEkZJIBD4IZv6bM
yn7cXPciv767DdsEywDZTzjLdhL7zyAGPoxWU6v1V9ZwHwv9CG4Y0uI98/n76kPZT7K3/ZA5Stsq
aJjyQd4sWb7O6FehLgwRSfGe3yX7NOrvhhDm28ifKe34yz+7w+b4HSw1cnY7Y6X0wGT02+3EJArQ
1hGwg6mfpQBGrMy93VwSa0LBpoENHqpBpyYNDoBN5IKptFzUHvK5D9qc+zh4CHzMXw4Foe6KPqdR
GjXC16En0zFuoObclt0htExHPAAgi3fy4eCM8grofhLnDorwGqw2mVasN4lxe9xaAKxxuEfey9Pd
OhtCsewpN3mTf4QXWFM/H3sn2ZWbCzeM3phHXmioHdb141EhyMHdcjtzIG1fulEp/3Wx2CS9Z+/3
AAt30gpN6LLQu9/jrPDZ8kiGqAmUN0qyK78Yv6vbK0fRCLQrQIiFn+UJW8KcsRH9EUwbXd4UgIGr
G048NAn+Qkqo3jG+7hQEK5CU4jpv9/D/hpTuymnO80P9aSVK9QnSgzoVTSRReZwFQP0Frx+weT+9
XTlVtooWkb3v8zAAOM2h3ERo7YmgedFUE6RYpiF3BwqpuYKOO/Wr0vc17pbrUP7sJvylgB2MG8Bi
in0npFoZzb3Y3srzJdk/+XIP/E3e9fiZ7ry5UCNrjKRoGLhAQBpTpw/8bVld0Q1LlEgruwAbqpD7
0M66pPYiswUXbnB1/qNLOUz6JsMH+NL48eChbOROKRw2Wtnk7XpkANN4bD9bpv826LHajtJ//BHI
+MBpFFOk9n1HB/a5ihU0lRxujIT7tybmEV7YgsWYJBjaKHS1+2k8ZaVZId93GKESJqHFS9Q0sCnM
bn8+BNhzqiaX54oVn3AyjXyLnMF70bNBmjWvIp/fHY6ZK3DojjYTHz5iAkBCcjlMYKHtfNuwHg/v
VGh9YatXIi/dH48HVkpGCE1mZ/AhI0AfxLli8XhTZCgLh4dWgDQihnTD9kfe4iAvdJOcX+BWn8oT
2g3rPOsXYWe4XwCw4IjmIvw+CLwtrjWbx0d6kPUll/GzmDSYwO3kDq3iwJrQhSf2cH8Z2mepklAt
1kG7ncp66m3bH9rfPrBhLNLzZKeSqLxg02iUZ/jFTzJeJ8YsEvgR6wV4LOR8kX59FlUACdV4gMRy
4BEEwk/7HgrNzNnIVFND5kcdU9BujXd2lISz4sAIYiOnvqUFYF2pCFaIjuSUC8/34Vu+bFsZ662G
EcNPvAUmAowDgJGYDdvVF3Kv3AmMuu1exe2tFsGxazj+5KPVrNRACk2uot0eQ1ViUZYOwZfEyCqB
iYvYL7e3aZgYivQI+1KpiWLYCU/IDtjL+KLhWXtbc+y3J1GxuZQyNAtkv6UX3FR2edXLVitdIZlJ
+yDKyqfWIORWJbkCTlRVDof3Bz7RPhB5uDhTzF36GphWIMPj/v+SjPwQGO5gqg33nUo074puxDZl
3BqxXrLV53gwToXkp5w8pt7/xIe2bkxMbQF4cgb8Xcc8frKvZxaEvwz01RxNe3o2iNtAZdueZw5v
IBPS9pMvk5tfm0c4ybuHEEaatDkUM19LPI6pP5eFZ8vezzAgSEwYEbmH1BFjx0LLYqfsHAhqnA7a
JFI2XEUC03MXG1MWY2Gvb/j+ouPkWR2vQcU0kk2GTPkJ8NTALPBQWr5yJQ2Foa+VchQR7ngo06eI
ml5zdB6KD5NtsG3DWkG7QwwDT2mICAU3ttHw4ZJHWwI37I0PG8i/9q4lJebLkTCzmjp2xzru3CCG
NuQDCJk/3TXgimX005JUi1t6i8+5xESTZxRDu7x9x+Oq+tyv461PdPCNQgs3uWnMosyFGCfTJtd/
Fir4L7kWj6UD3qaVeR4d5nRqk172W8U7e8SGZcqKj6eeclxBm2YAkPv7YfibGWuNO6kbfzr6DCA5
/xL2yS3TX5lY0ryQMSGH9e5EncR9NHHVBGdG8ZjcH5t++hRGqu2DxPdY2vmGyRU4AkOEEwQhbB2L
cA2jExhgkegHcGn7YUlVzHNG1Xgx3FvYCZtUVO/CUMlnb/gHdQ9AhxrnYs4Nxb7Pf8LPTU+ZS/02
kLyHkDUw/jOS7WC9xOcd7F3Gyrj4Yzf+SBZ2+tnL+0RH10tczOw3zhAlqDyOGiWwlPewTOaXiQEV
gOCTmcpT6jgxzAiMpUNWQ3htIM7fLGSqaxWBBk5LePXMZ4o1wruFE7x0/acE1ZM4K4CTx/CBmvnh
5PMMxtbVDPSd5xMkVjRmvPlQ0HFl4AoTVWkN01UQFXB1+A1SC5AjtS5hw4atl8EyVxsnTY6k+aFO
rjFA3J2ibJVSP8jI9/7G2T/xn3aUFHOnBEa5BR6WxDw3Ai1ZspzrNDojRP8fWdhl59KFxThXH27b
f2HeCYpfIO5A8XoaGkl25YdnUGtJRnmFU7Ml6uFH6IlEVBZ6+eIz5HPADu0P3oLvR2aQLRCFf1FJ
/NFyzib0X3lT3nS+RBt9MRjFoonb5l/tWefzbLEZLWCW6byTmUZpjQQXgeWCCdUsEPGTW0L33uRf
/zE4qY1Ut9yy0MMFnZwKnahXxF4EFY5C5vQZVjy+M9EP0MzbKov7HsLyYzHAkScndovU6L2k2HVO
c0W930t3yJlTRemhmi/TuPsdxXv0YihKoTI4/eyNAUHE/oCiRxAzOy5vURvcobSHJQuUFKuljtZh
m8OoVIwGy27Mx4d4nT8Asjc205nWghgtxC1vioN/U/WwY3HXaBCVNuD1frsfypqvnjk/ezVWuIHL
p1cL2KEah8f+FzHdR+eqfuipqD7RMHFnwVSNtjSURmmjEk3g2FYg+M9mGPtBxw7MjSEap6oDsGMk
zBBEBcGgz3D9edD5iOrOuXaBSL/4RSYvuEBecO2jeeYvsstP/MnscxXz6QUToEhQpoR+R8TD5iPz
T8q23aPGpvtcOwWQqKkr35zzoCIOh+subQpp4nDXqK6spARsjQwwJJiDNcqNua49XEBYEg9mqJS/
n/K0NJZApXk05WyTUKJXpAomCFPPXX5vDsHnGKuYwmL/EfmaS+6aUsl/ql6/5HEDo7S4ljFvunIG
110pBL2seGrtVwbBAKUjQGqi351gGU1yoExR59vX4qolR+ckeaQFNC+5g6aJHo9bmt0qJ8F6WtvU
KP/tj4w+uox80FqPNHBMuvMf+X58Sbe255ehGPESIEhOaC2eoyskJhC/gLZDNHgECn0jxwTuQ8HH
JvRIINgk/9L5T6Q66hvqO64oTZ2UJFNb8T5f6udXZlCJCanXDu01Icdg4bEjKVI0AXcoAXgf5T4t
ASxzsKDCOuiHWiHiNyus7QS53RjX5MiEMTXcpJGqWZn2eqkWQetr1it9RXZ26APu/eyfPOVdPzJ1
GO/jg3pce2zc2Rjw2NwnikntZMggM0YKYkdP+QFB0dsk76QvpUeQdFoUbNCw97fyvCEDS8XUn5XD
ObfDRkQHKJ5/xTcFPkoH/7VKFMzLA6urGw8pP7mEVsA3F4l48x/eaSA41UFhOrcMz5xxpKKym+vf
ARv5wgi7TYDypvchndBp7bpBg8itQGiJvEUhGI7FMwztgUTvC6P2T/mAdanw4zp2VWssPvA0ym7b
bybgS4urDVuCnjYLkse3yv7BNolB+Tagm4SIrhKR8mhflG34cuRi8aNaaulXEBSI/uA8nwy3/Pmi
P6XAR1QH3NouAOyOhaJRwKi/bFGkgTyihQwep7liQ69yAIFkFqw5i6Wjl6qRWGTMyzgV24EvHhrw
YlILfJxFChnrpVG7zHCWtAvuOSy8ayriHr/CaKl57xkM7a62RmVOa/UBCzpzlhiHMNyQpRLSnihA
0IhaQy/MJ5R0o7dWygZGM7gviqABO68sc0kaXr9OwWQjbtPVXwVN60QaI/rUfMrGyLcHyvSzbLx5
qRvABrdoJU8ywqE+oV6WSKU9OkK6zV7SzLrbgKhRSVXfKHEGtXN5nZVgxmR548y6jyAKlzzSJ4Tb
O5R5Ud89vZzkoHUxPYIDmfHPg2NP31SBs2m72uLFhG3PGnSoOuBCFRidigsF1Myoh5bhpuNucKZS
tK++ssc/Uoz5ZabB7peEA9LkPZgtOhQ1xIVspQyhAhl/Safxnjd38kXDqF3Gm4BN4etyVlJUJnGi
0GM3U2D5xg/2LdOaqSmnCg8bmn74Ws476QpiUhDhFZ3+Tum8AMuuN/TFRQqGevL0akAHz7Bdv2cx
TeZDZhcM6IvN4b98vDh6cTypuJpFvqTZycHk66Fs3GCXrCgq/MooratFYdFY3GnMCInzwZturxxM
af9WWiguhBNHo4K5CM/JL6dB19KGh+THvvcUurfGhgvkMYBAB2GGibJUuaa2L98QKcGatvPV5UXo
g3q6IhHX8+K/OXiq/5eG3FAg6eM5ujy2YVpG9/5Dvwk77P8oKmQKs/41djsYbRXYTqV8aYP4RtE3
Ilf6lPXfK0mS0L5fmnUN/m0okNhCQk2cMPH4s3ik6cefhpgdPkuVtncs0RKveIzXtL+JuzNstc+S
SKZ+gtyi11S6nYezTheZ0CYDePILMaruLLNjMIUmOs6txUehTEYy0OtX33EyYw1SAc2xsBMtmpFP
MRVfwVOWU3/SvIE0ncSYokc6vJNMq3Git9P2k963v+XQHHDvqhYpCvo5WCNsjgdDA7eK5in/wPd9
CMmDCkbz/EGupIYt0tCJcpN4K9wr9QZOsPLKHftomCW/zLj1Rk2crB2T+goE7IRH1cpHtf9IbyM7
ixyZ2u1F/ZMsl1ha68iSTJaZIBjWop+oGJUS3NL0rmJr5pWrYwdjJI0fzYocQuS16seh62p/wlLt
dvrcznxqwaGgKa+wsXR88gRbTtrv4Tiw8pshwuhtWia4sBUNcNfVzlwALlJX87BI91DnCzyri22/
8l7bxUH7yRH6Tnb+y8mcI3KTUTNVly4FWyHFdCG7mOCZcLNvHWyag/8lF2Y+/H7rye4lyxvQHviR
zgrlKSOEuZW9myycfovgzQKD+an2kjklwxnY3/F7oDqG44yZAPMX1TauywIx+rKrJmCTcNoD9PtT
Arqbgo8lAh+z7msSFnqXGCmd77RWbze2OGBeQjKPfpHYmq9YvFRUnScyFdEK3z3O/nAlnGnFKChu
htqHxEZcAI49+FDGHB4A0b3Ko7VHsR/VR+Rp6uteEA77MFYdHktDcYIqJbcY3K6v4JC2iyCsq7pu
nUfZYYc44kCcgVwnXLhK0duT4oPitP+n1aZaspF4YU6gBXAhTkB3NKBx1K0CyypcWO8EG6OymR8l
Z/dNXJv7UKNHlkHDr8BEmk2sbfL0piEi26cS/jYIgV2YApCgtVjJp/Eo8s7OFer63qerPA1xGjCZ
rA839jAaUvopXswNEusCKNARYmNNlV+EMKsnN4Ci7c/ZcQJ+zIzOV0eEY9vUbsQikr5WnbrmbtGl
65XprU897/Aw+htrE/IlJAtKVvCA372DJ5vg5XeGCEBJFZiHYIesP4OnVbdsdxa1V5FOSmVz7vgy
903ku4ek+HCyNPPTNj2wlAepjbNsuE1u8gbtPlzV4PcSOyc1tN8e4SO0AcK/jPa0DjMPW9UsMFnU
Q0l2czuywS9DvVz3z/g0Wg3m9ltuZ1ivNb8OfM3URVxZYIj8RNQSZFEKoEved5VPnLayoVAo6Wwm
xMlC/Vw1lmwc98UMCqg0vXamVWih3Kl23lLtoJKCZ6e2JABSX90OQRBXL2REO+Vx7bKRx5w291AS
sQf/eROyzaOELLtnAmhM0+BX69Lt45U6XVxrDRNLcaWZYliBoBk1kn3INYeQBR1deaogtyvYpoQi
60sg9kxXCst9LX554gaZ1YzgHmyvl7WMpZykDea1KolM3mTJucy065vrsn2i4OOoisYKQOVAoCI2
tdZwGaEpmYMTiXA2HFD47x833VEGR7XLZ0KilMjNKMey/cRA2yBpHTUHkxfuKnMJkiIJcBsCo2V0
BPVAKOtQoIW22O2C+t2VYDmSydVUZlUkfACzRj7nQ49yGaln6FC1JA+e5410Pq2w1bNgkqgizWxT
hSAQvh46f1LGk1Qxwn2tY9QqxLHlw5NWnLV3FTYbBWyqSdMPN/UinUPuzAl30rGH2c9FAygOPEV/
vOiSJn3UpkV4l9RdXJMD89Dg4ZEYNwFsA+Rkm3RJbiypVaiGq9XxgcVOqbIgWtPWXK3fb6JY8fsv
aEF/SPDuGxiVmkcGbOjxqfEQEs96tbuVGSnzIPoU8uqNUZGg91PtUYdRLffxzekjnDJU+jpaCYhT
q1DhT//1lHVthIHgpsVgl+v1wnOqTjTGNorvJsd8YOBlAy5gs3jdgO2K53Q+yvTdq71Kg7NYFntj
/hq5QHabPKUqg0KpDnBfLnO8warNF7PRUb+Z0Aailm2VFaTDWKNK5Jr4v0lJqF5BoElNZWR+BL0p
ewZ/dKTnwIbJUKaIdbjjw3ZkS0BxPopQ3ijWd1Hpk8eR4u4hI34pHtCIcNSbD/+QP6DG3Npe7dnv
K43ccv+zLMlj+ygJyoYDNlFBNb1htw8bPqIWp1o419FWLdkINNNKpfaJFc4Bl4PfJkWJrRecVcrk
K9En5FNz8esxuXlW+UrywyK3e13NcxXYz0yPcK6uSmy4ZdlSsWatAcLM4ojWS3PWRmzZyJn2QcKn
Fja9yP7o/cBCuVa+FXdRQl+3Wd4adp7pPGnlbxwejrHxyQJw7aJBwHPVDR9/+o7dHRJHPhtyIFLA
XF8hW7k8SbUHKhA6SrUT3+513yoJjzNs7SG7t3ydb7H/Hsb60NZAFeIlQEtTLibqHKZHGm1fKPJR
C1uE8tx7CJSEW3p5rrBjAxWHKAWmA+1LpjdAubebztL1FqPI08ntUCrD+EUiYnO6avjJ8KuoPHEC
HPgpw65xTGwOXi9gER1I0A2tF7rnhK1ijyynznckIOHTTmtn6+mX5B6J04H1inIYzQPguxZQKt5e
KDPaN7QdjZ/O3UIxB16ha//pkka+GXegdR9mJblcA2+LShErs+aVi+oJcrIsSZoi3pJRBW+rY10r
ZkZ4VvaXMpLCktLRHwUxx2YvPaKyjmZ73scmys2ycIZruhSXGiYhae0PiwYJAG5eerP4SbnvSjxm
kOqbFRNBwaUB8vz7N/4Y5EZsd0Lw61oq7ggTd+m+f8zFuZJBIxs3x6vDTEarP2YN1VGZaiVNbYEg
UqgWC/0q80gaVtMJeB1Qdgy0Qmb6f/vbxvGq90XMs/y0qArQ9tWiPJ2f6eWiNnUft1Ko3dDuhFqL
WXHLKdn+hfLNIgX2mVOuYuuUUXeG4pZIZBXDTybaDI6F9dTTZzO6IrLIM+f9gVleR0OX3dcoorGd
Reyri70mUWQ/t6MQI//0m6LNpulTd4JP2m7NctWdAtkWPuJR/MSLye4Rm/8BzS0Kgn4PJ90P+ZTG
3e1QZUTIhI1+TwRxXYTD+/G2ugii/ZanXBp4Un9Dn1VtsH/heCeRKp0ruHbLRkof+5tsnMXHSG17
QD9AWRsDSIMjbbQWB5j0trPUPr/8AINHgJVAE2PqdspastsNVkFPIsFViCBv1VRBMcuIXAcxZh1P
PoTgJjNAZLwl1B9GiTHv1OtNVID383/bOXuyOpKo3AHYGnmHq2xiA6r3Cw2ppS8lZOwr7yWKMesn
h0bbgrY/oegbZIqUgZjONxCG4+7q/RHYOD8Obwm2I3MyK/XQVQp2w0BTu4fhOqqo8mpuSjhk8efY
zlzXQAaYlPlLPTbrC3cEiyVdiEETnk5liRlvFCGP3pJadMsi8UwQcLHdbgyMTC+VfyfTn824R7cn
9EPOKeK4a+/WUWDAjufKcavqt4EQ16sfk2QH/1uoG0W09Vegpe5WdnFtjQaXM4vicuw9g7Pzuoe9
i0+ZsTsDJDr+Q4MwB75FHhlUFlsvoUi/SiH6IeEg3pbqXj4fZhxeFve8FQntveN0TJhkJLoEhF+2
CREEwZxw72GYV3TWiXwsljQW9lsZe03wg/vZLdcdiId7L7J8N9h06aAbXi0lFEHa3kwezCbtrU3b
dcVZqMw8GxazohpU9ru3++lkf5qCmryzPNfBfnsBIbSiNcXCY1PT9eAXWXZf7EKsIQoc2iMmFaQI
CyT/Ae4rYVL1A7TEX43KIqE4aWy4IoslBWzXlTlgeXH8e9zZEZitpjLyXeWry0Vu27q+AypENs4t
2C2rEV8J8gsUSmSbNmNO2kz1MAVVu+bi6Kq7f/jnegHq2yNUxSFRxVcn9uFBZS+izeLPF3/A7r/a
KFTk8KnKFz1NCQ4cD7PAnS8nXTgBBbf1YZEAFMv0upRp0vcEXvHnR8FqogI6fL5/lpKLfwk8AFgD
SuWGdsspKr5iG8uL8RrQ+Jm924otLzVVdoSWNqj1KGq5qOv3dFHp3xIZSLANexNfEbcTK1oNdm8p
4ulKzQTfa9vJjqbquDthb0wBAMvrI8Ah4bFfKgnLaNCQe/Bo2gfCKU4smxugqKszzvkENhvaWju2
aLXcrH0RBrxOafYFqKda9QShXLjbu0c5xyOimgX+JSfcknxcLvkv0ibxltpo5njja2ZBjw59uZ7l
UTG5Qgy3jmKmP9msTRrP1hkKVax4J4unYYTk2+nrmd0ZNUgonvI8HVRnxZaTPswZ16zDIdz6nwA3
E77XkJfAtPCDfYOaJgFV1MsH4JnN/tugq/kgkObuFU1+73QoziU8UI0DMdrZpmUpRvurk3fnmcCf
sCydf+i/BRFY4/VltT+/2J0xvJ30ta5eY/57UBuGvo2pLCDpiLB6/Dthbgge7qv7Wmv3RMSL+Hxi
Km/oZDEV08ks25DdWMaQ/hpDSLPVid4p0nejVuWgBWsYCpNrkBGnrjmLhGo5emOonuCy27d9XBwH
ycm6XYpBB16rrySU6jhKexop8ccge+06T42jmQblzD+MBe1xq8NeMP5GbzsvYN+OUGUOhrfdR30q
4sXc7lmHGwLz50J9zYymbagunJbegi0450sXPPdlIIBo7ujmv/7RykQAwrP3ppXDI87aCVpwy/nV
/0+JpNqt7w3Ee5G9HOER0ynQ4w0K7pAVaPKfsEayMKmLvZUKllSV2xymRM+JhxSXit2AIk6jktou
FHTWmvbYUZTkwYOGZkKILpDC9Jvg8nfdbPBL2wtIie6mQpIebZH7BR2cx1foT4r0F5htE3U+n1i6
80muh3HCu2RoGZ4KuuUL416zvzJIaVFVPvqCOeYKgQcTkA/Xzem2r95djCuWd0SNw5MPrjkC0+hY
V6uFOnjPFKpmjHUJOHv/sLjDrhLO6Xyt9Jz2AMrr1SOu30S/FcNhfx5eERZxCjzqGcLFJ91wr40k
wVDysIlSh94phCGx4hncul6J6OYeqluaUVavndmY8BF5CZH82rdkQxnp4FmhPoDvpDTsw1Nahrow
bkTbMICGo+8LNAoeuCvRAU3KFs/g7Yccckz1BEjJWkVcmvb+YFsMVg+AeoPBWpZyhW25tWBOUACw
9r3CbYgxJJVXZetRIozJHIjmf+qJ2p9S3/TiapRCsVlw57h3blzhJ/hul2zV8gMyfMQamAav3c9Y
aqNVj9VrmUefpHLrcjcZ9Wowq+YPodjNXcazz2AZ7Oo3FBr108pCiha2Mahi/T1xYSSOP/o46rzS
TQ1OBMr0Z2BMlw5IfE5uxOvo6xyFXX+fpEhjcERzVwStkhH8afGFpGoxrvCWyPLY/RzTZjEqR4Xn
Xb3lJd6UtRxNJIObyBtOBvJ1vKwlq/LyOYjVqLkU8wD9Xjg0mipZ4427t7w1Qg58PBkamCGVowFb
CsAcCWL+TpHEFz5s5uP5WODO63z0zBZE+9cyJ1aXagxqjH4jZj5GajeCS8NQgHolAxpkcflIFWP7
xQh35BA56cWch7hxe6Uy25clAW2izDjNk9zX+84gl3aGXgTBuJlbob8POggP2dzo7SrQ6cYBMuGx
voDTzsVyPoQvwfoN9XMUPCKsr3DEc7R3C6KPDtpItSlgD+nOkqxG0AiMpm3UNzYx56xOscVDY3jv
cMG0PuRcVghDR6SOhVmwkD3GBtvLpWrRmSaZq3IVhMge2y5A2ma12S/CIiTD6cPslf86x6A8xIwr
JEn0I2qA34ZZBqzkjhUEot+FHU5Wo1Vm82JTotEIlHqhEeEFbVwrZqV0X9rOcn+DFhM3VGA35P0y
uHssAl8XYIHb2DsOADI48ciIqcy9Q1OBuLYohpywaPyyIoaVAvZtnSabZdr8GRv187HM4y9eovqu
NlDAD/GuMNJmTXmm6QPmMNJVRpj0yJANMFmbQiW+J9ZNQteCfzzTK+pVbzjtU6SGe9aqQvmhXpME
UngHLtXzLQmEhN16MMLPAKMEMSxCGuGYQlEHaCVz5bcJBQvKvZDVBwTJ6etWlPFA8JIcFt1UP9H8
d+q45sNIGTPrHR4psN4xRNBVK3vNr/ctuEzmxFlS9Ouwv5ZYPOdp2v3UFD6eZLkLfMEPfCBLOwNO
siW6k2E1KBCMUKqEvoaRmdkmdHhilO1V27Dvs0T2LojSEugqdFjou3wt9fTyXYNpPcz7Ct3nviY8
bWjuJ67wyQHypZY7P+XwVYUDqCXVZQadiJCZH77xQrmht3f1o7uhWWo4F7XwTxKZNCa2ugBa9pLw
7haPC8OvKKTHDN9MkzYoVIAS7wtuJFrVfNBjYhG88Ri6PfA9BhOCje0fBWQs763jE0bend4vhSud
nNMqZN1Q4AYPeA9lY8kQe0GHbI03p/3czTA3PKYrPromtRX702P8KRlJgvVndWPgUqSWZ4lf7ewx
EEStz0MHhzIsUpuvjIcEyFxQnIxqVkeh1ZlZEtFz3m29d6T0lcRI+zAJoFe3FuFEzpcywnO+O7rF
BR2jBGFnPSH1eUVkxZGUB8rnh3dFPa6gW/vB91WsR/ROrWcfNh9hqFl/5g4dSOQ0MERwZS+JPcys
ieGUoHOVnE8BiaSLBr5qQ2WQsbCIMliB8kBYX31ORxWlSAW2xvy9ckN31mxX37SJpffxAjhJz6h2
6UNFNtCDcQRiv9f84Gw/4X71QQNllsb6+18LYXVSpqJ5DfkVRcie5nI8pfhzq2NlkIFii/e/Mkv7
7I+RZoqIB8+L71IggGGzT1SSU6Ai88fSUfRt2MJSInguWnGK6ZsejCAUViaCxB9yjbOEqz/+8Ogu
9G5dNMbigIxhGv5qYkHAafqlYp0FDMzM0SpNS6AiEsxYDQWeFuBrANgOR+XBY6OrN0joBDRC9rx4
nwWLRjoJVVabK0S8shUp1HidqVXFH39YLqHCWl3YCCj6LrJCFngEQ5icbpJFFiktj9Oxlb4cUWxz
EKQ9fbObwNYajOEJIYwqbBN4d07XFkoBfUskkZvavHx0Iyv/QxAQqqLuvdX3/he91ei+quQx82Zg
YV0JtoMxIlItCbkxESCpIPtO9GuPTRSKmGzd94zPMUwc+rzWEH/9PnM2RBCooYApy+wipAtHPJoX
9n3czZIlYN09EOOBu33xbzWvq2HwQ36qBkGWtHEVRNoXVdWnGJm5Il0ttd/S5iDEy7kni5432SJm
WvzC0iL1kfcyy3XmGhCE/Bdn6u4f/bwIetOgbCwOetaXU1NBih98f2dhr75HWnIVostXsl0IWVJt
TF9q8uLCcr+YEed/724VKSTaP+dCFtnQq49lxcNLzm1y02Yuyg/T0CKQ2Xkxx7qvg/gTL3fhHR6r
3Ry8Ccjbv1M/3xoRRoHOIHxHm9iaDMyernvbGmTyyEEPQRLPRzHKzRIrEg3hoTiACeuDVq+iZV64
Vjg7L7S6KLIyYNwXBP/29UVx15j02c+ltZ+Ga6fcN0ks4mkwKD4gloSlmTucfjSLdYqPCiMQXlaD
vjm5VTi93QdbveZsJ1b7yYv/y6wkEv3WG/Sp/bw8ZQ+dNzEgUt8g/pYhwoVoq+RnOy5dCqkvD9bU
9uZ8WlDlP4Z4VTRfxPvNSS2gfOkyLd9ZHv2Ta3awrqBF1IEPO5nf79JF+D7wG3Bl+Fgd9RYQy2wA
XfmoJRfIB477yadOIfZngRiVD0pmFuTLTTWG7/XWmlBRmM43nEiBKuryUi8v6NiYaRZYU14vWFaI
8/GUdEWXurOteuCiOa4SHhqK3YxbH1m0f+yN5YYPRbNzIa9I+ZCAiMLfn2ty+6PV0yVia+eUiQvP
8eBZFAbwxQW3tXo0MUWqAQ/yRTlQZ50aA0YeCkByH1wHrdlVl4ghJ0oXhuypsMJpe1+LkUYkTEua
hGj2WO1q13lqqFui4G6nSxqMXRC1+YWq3PMs1mKme/RzhwmZkU1bxsQop/CXsOUzSA3ONtIdNZ/c
A5COTO8YB1O3IAvaYAzmvHJjitSjQreVu0RNAScsvd4YxAGiRbQDGKNXL4zrGNRX9oPLAbAoXOtP
6VzwgXW+fUxTGZnN4msIuF4LoxXTflHreLFxvST/AC9sFzh88VWT7odnSkd79hll/Fkasg1fXFpu
bpFJLN8pYhW9H2O6srftraE2es1ucrSsy7gFWJoi9C/gAVNTZISvZJG+rjb+YbnkdpXYbaUb0QHM
oX8uduoMI4Nz0JYl/x3x/Izfm2/8+L+Hk5bXBpUBoFzZ5bt5G1/bmkbluQUBPQEdyMn1LUwOSBDL
vDcOgV8VaXqFmot15/LHA7cTT1X5AMNLGcJC1sTMMl2oZtscKIoJP6PZ+oY++KV8hQewZxdUgQVf
kAfoFEgVk1BogfFifBNla16SnrOC/yXgNIIgOKFG29RpSOfaeKqz2T1J8Er4LtMlbXWPzQeAo8yR
zPxIqteggWCYDUeuNbFo2fo0MS2LKxpbQadT1FUZ6PuNZido3PxA5JNq/oSd2DWBS11g3q96d7mv
4B3Ea+O17+9Sh4YOHiLcP9p95hvh2PQp1v+oo/NsX+zzTbJw0mQsxLSNtqmvZ/qnIpHnarGl5zaw
KZVY1hPb6/49X8n7uOoAmpEgMOq3aZcMl8LM/D9kNkVC4hrHvuTTSqk6C3sThXvEylYWuoVQ6WOd
cKvGUSUpBagik9iSdyBqYJ7BijceceswWMxJMyqKn1m5F4ser7IMOL7TZabVTzKehf4CgNB92ASe
HomIap4//gAmazECciEKZazT39U2j+Z5zj9bbWjhNll7VmoSdYUH0M1mfI8glxKomWV8m3Sq03lk
SC82IUR1+RbVpGca58vWAtS2exnBMHpWRaOrjCCn2OEQFXxsjq6li2ozdHw64BXTPYOQiqO1chYY
tGUHCskxkVyYq+1cHr7l49OeThDPkvggqJGduLPB2+aotTUdpCutWl0evMa0CG47bEHx+J3zBzc/
/N2WoKZ1fSBq1idS8kJYorj4mc0qQmfODAlEjWBpGF3PigShiNkt28lVgIpuxk/UE18BHd8JRLEv
xwUsacA/yoKCE7Z5gi/qLh2iXELs1yICfjxDO8tIrx0aQZ96vA3uaM0eKlGZUhFRgtitx2wGHNgZ
4MFiFSdIen8IqPrUARaIx6r3bV8BulJg2VxDG5XWkHRN3i7N8pyhPUCuqIucOkHjdd2fJczl1D8b
YnzABqCNe8iHiMLGKBgBFlwlCHUhRd00cqP1VufxeuGDE2W7az5m09tScxr5XpDAGchMjOyg/Nvt
jUniq7zpgxF955sFTikVvN4puLXS4k6O3rETAj/DDfzJmCE8FUnQq9f9LnR9+HbXuBGt8nubS0u4
EPblYd8RESPECeNpc5mhkA4eeST5NtXxCr7Ih8S+tlJMFdYoIUHxMfVFWZYY3VyBxnlrisI2Ei4k
d5jiijoocToVguo4YH1ozOcpCvBYxeKAQNKPYB+q4rq727WzEKJFkVEAhj8UGPmdIhILycDdFpmp
v4mtUzrsvwdHEwr1zJSObx4R551u99mSWaXdTIgXyZJ4A1KrUS1XQj/or4Orkb51X21dBGU+AbfY
gyQ7WT//8m7bwWuO4j2lDfJa/wDvyWMfnf0gSe9C444IJ76LSmYwnVm+mc9V3dEYJIwaA44vU76N
TepI2cg9CrhJMFynmAHcHB7IXeP7mZyHlY0alYKf5QdQfn2md62H5ZL5aJ8fTGFlSxVcLJcHozHC
FGRF6ZvRq8jnwKNvx1MXot+55lEkSvv+6+eYSIh/OEcfcGTJMHfsdT9ahI1D/EWToT/eLi17wpQ+
kU+iMGxBe2MCEMOqeujLqo85mqLQYW8nj0UZ9dqNx+Tl69HYxyZIG1C8Khr+WgcATtNLXiL4/TF7
AkyxJIkwr2K6NrTJO1tMnei/QZam7aqO9kgCU6JJB4KeT4jKXf+9f1lPdjrgOu+99+bKLg4d2sQD
ibFWOY8EqEiebwK+TfJGgSK+8LJRjjUtifX7HdUCMkK50vKNe2xieri5pOFVOqQFVGT5OxYi38N3
+1PE7VgZr3DhMTZKxx8axQM8b4PgYrjW9m1avluq6pnYpjVGBDmCkCwozORJ4ywwtAd3Q4iyaH8f
2sVMXnL3sKpWniSX0H/rswVd4jSb9oLFfdjFksclbQFAhS/gcn9yOFgdUP0BZVVm+kgAKO47nfKj
RgOYa21QTswst8HKsHYMvJK6ZRd/GJj62z43Uqqa4Rj5xowt7bNOuoZMXVW6mXPZvHnLnsv3mL+h
e6pk+6I61JihO5tMafFxH8THObgAPrWDjEeNpHnDfaqEWboiIUXuf8UzaqLgrlpXg+bd4aLOWDew
x2yUUCVwookANJsRHMaw8Hw1cbob+0YuVsp9DTdRZzcgA8EqGLZi8jL3qaQQ3Jfze8VjROrytk/P
GztZWnAnbiZSZk0ATAM5HgWSXabGMoUY5rqI0hzR72Yo48A2k6ZCOFw1Dx/geG1hwf2j2HUVf5p2
laWz73AwSHpOw7v9QYUvJkvQ/mHG0190t4aDwl8GK25hyQHJmJ9gztriiyqukpffeVRzO3ERpczi
jZG2ic3gq+/DF0qJJRQcV83uaIWeEZgDUMz+D9ur+Fr/ekATQq7EqWaK4g7VMF/dOMIjFvCronrB
WS//irB+9ctA/b8KyFYms7PJJOCFFa3kJcCwMCZMel9secqEVdounH6SnP+VZkOzhDXh3hs=
`pragma protect end_protected
