`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16032)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrM41f83zxdpq7B9Bxc+63s/ThO5
lR4ebiIUudrMSnsXzTRn4negwrrB4VipTwcqyfoZbX2gIf3gPwkP3q41DFrLyf9opSDFSsyylvuq
0tfuxhMWxI0KvORiuv+DLG15sEi9Zilc4jLqmJBgxaj93813ixDm3VBlIU1BQYAYzQ6XobruGhlp
W7l+H9tAQt0BvNuSDNd6KHRHtkpbBcXPwpTyA+6hMW6u6Ccsl4qsUag/gM7FTpREXGWubujKpgQY
rp/IZCyMTpGc3aB3VGl9Su3mHPexcA8bFwc/WtJprApfvCcjuNPHSMoRig/QdwYvW7r63jNqA6ay
eE6LoC8jRjjzApFYT2QXhy0an6uJ4lRzdqq8okg33mKXD8LTtEuwkjvIrFP4TMRdogyRsLRwnCUF
Vl6pZC2ALOMmYC0mBxKTLXa4+hwCpkU8IqkUAtiuTwJ9avrQGEZvAwTtBEL8erp4/uPcQqDLPoG3
Q3biWWvhp0EbP/AMJfIV2DlNac7A50H7VDpnyP2BhrrcMebZHnkmzQYYbOFZDJNtP3kSzrjDT7zx
iFGBakrxdAqZ5B2WBiiYrR+dPLTApaH8rg4anz9+Op7d+eMVztBC3MlETutkH1nw2AGq4M15fTv2
Eu8yvgvC4JsUeXzbFpniZggYNol1TVPyk102TDzuin8rngqIxjmZPirVztCcIKaWCYVbFngY3KPf
opYRI4SrhxBUjIXREEgRH+RhJbvCBypaGwYkUgTLu9BbqMiVvnYw98BaO8Yg7z7xUDqZ4e3Y9M3S
v7mOTAHAVRZeGlPpcu7suuP7TrmGlRObj1chzuhe9e3ngdM/GDhia8R+7rjBqDPcCPM2sZ4JIQ3z
x3optJmp83akfu0Z49pdR28gm7nyloSovbp9EbCQcMPXLJyyjzg4498Kj0iAajaBUMoUwXaRM8pa
6zgkmSUg0VxfYGn8K9lyd14UmGpODVPaPawxDoZqR8a12OalVWdOvGZecZ/rU7BqQvLhTNoLZ/7I
cuzugJ2urUWXgVqgdYg23l4kXV4MM4YzcrOW/0lRqYUtCHUGkjWojt9K2qI0QR6b2abi3k6jsQgF
2YYYmexD+Q1I9SEZdCbj5oHbnQf5uc+FMdd6KLaKI7IBI7miYHdoHcz34gJ7XSLYOaV4qL6GGQ2u
8l1mN8is6WtGT3qBODeuNCDkA1Ptr4P6Y4SQInDZ1ijzfeYkCFuhdtiZkBv5zBZFbEafy0FZItZA
MCr6AS/QduJdbZfrUGlvRKlh8ZF9SrVgppGJfPv9+H0WWWGyy5t8nbFpZdNRS79kNPr6dxDC0XLY
S8o5VApfemIkxli+KSjYhYq1JPBHbQkMvEq1rCFl+SBRpiKltpFByzp9Ywc5I+fnQvuJfYkhwr0x
el6+rTCh1nmOP6rJd+j8rFfCSdN38BggNbxG9FhKXosupkiAgM2/rw0akssKpYuqtRMwCA9dTMt4
vZWM1LL2fIO27ftFyHVN+gTmbvXYOQ0VWMsFeIgbLM6+OMLE5dfSUZvxe4tyMjWfua/37b8d5Rfo
croUPELNS5jKcezFYsojiq9w2ADEyNZeUwIeFNSpafrB327/n7JNTDKzQa83DOT+R29Ek9Te7k/t
B/z6owO/olZAIEhYEySBNAl4pKRN8vMEuGu9E42EJX+aESbpS7vh8iJtCsLUko1cAp/c8w+V5Uh2
rqyY/CTZbAj6QWpVwInmhaWa/f4iIriecx+2BRrMjFgf+hlpRe6Mt3CLUXn5r8sqkuL8ddOnO2IK
xtmyiFYUZ0vpL2l6iwmd4BZszQoxPiY9BpJ17rOKxLRbHZdbJFhFFIcX6oi9aCpatIg+Q1YuHZRq
M+g73J/Xi6Oyeo2/CiZXrysjyl6FK6YEyl5LVejZk+PJVFi67vkSjWrfxZC13skr7DDNtLfq4jXI
c/7RUoFQg8I/mbIQngtgqK5taDA/RkjXSkxg5xioH4JwCqAnciLXy0OxEHtwXnsWLLKdf2bizksK
omzCnIJE9ALQtAD6vGJZ/+0tgHWxLgE6DoZQW0YfzO44xZWB2EFW1vlNHwSenZLrUMD9J0ENQQYw
MIrEOHmZBUTGuu5wurQlkIb1iJgRNsuHDQE0GAQI6Fli4pyCk5ZJk/ndr9+hSqhfLw+Nm6G74O33
65gBy+nr15GulPz1cr3RO5WV5bDd9QGlsW9wIfinl5EYFXrqBXa8JqyoIUbTYeBpKca/Pe3dHMW6
d8iNmWxSA4HT5OZ8AndxrbYXU+k5GT6mh/ANlRe35sZ+LItGwgOV5wKJqfvXvjCxZti0FzpcsruO
BnB/3VQhbt4wjvqugqu2L0QdTlyZUxjCT6ppJG5m+EwW6bOcoQOaW4O8WdiPPrNnmlm/09xddt55
fBYczGrTAwf2Q43YzgKdDwkPEIzucj3yIQiGbp9xgrvikspexLGGLLG7RyYm+QnLiraXv5aMOhr8
9D2Ygt1erNlLHcwSxZV6N5P89W7B+HRAhia2XFPDIwwyOdMZqJkWE0qsm9xX7QyorHZNjilyI8CF
vzLgAE1TNokSMruhhLS7wRPjk4YeSTj8QILlf83AwzozE97mWQrsNFt1FbuB2n8CabOTKG6NQ36X
CWlvedzyAIDCPGgPoPvcd1j60mo20p6Yn/NLI84wPg1ZgAyEYXWfex1eT5Rn5o+VDajWAvTWRjvx
0IlmsfdL3yzK7sw/GGFaLzl+e0eCzZ5x2gGJyDtoYGzibMJAbax0wk2s65Wa8zOfzkMqA26LOfLq
6LHZwIfS/hHCOkS2ntb51UJGU9qRp1WYjMMSQOMPr1tZavU7mGwhgFGkFtptVGs/ws8NKe5e4NfT
zBcZr6/a+RSCvl4mCQdpM87kCKaYCHfSMEJmbzQBZWGotHNo31HDPmUwxfoweoTXnyEuyyhR/r+d
lqhTyHCysFkS2yzjpNZWA+PD09C5pZBkLRiGlPkbCdUfTZbw/PoXKpOlPVry4kKBpzciBoEoJx4D
/+3IIF3jTNpDWZpQVNuP494uA0EzbsRfXcsWQK+z0vABPmxRPh5IuLSlwu8Fv67u7cMY/J6l6eL8
ngnBljTtbVy81JEF0LrjJxYs+v3kK5Qnc96oNiCuJY7BiyOFp5fL6GrnVecRFf+AAlDg8oEWHooo
ik126NSU2ZmOyv/BxDgBog/7LkNdm4vexdS2Z04onUJ0LtZi4BRiPQt4abAvGQbTmLpCzbKKxMnf
3ZjewI1+e/wZDAtmTURS4RhPuutslTO34sxjNcWLVzEmrm9mvQqB1Xup/dHW2eSf8IQtoAh3TloJ
xHpH2qpTj1j7RlFe4F1dwjJEdzyzGEs5g/YijS/ZlYIPseMmpytZgQhiVyxUVjaMv5cd87T6+cuc
emlWmSiGwfWvlkSKGm+TsB83WiGEIRyIai63fxCqePYfXOcvt79G2Lt8OfwL4CL8AyRXsG/VZ0Rz
YD8kGFZFJqoOJDd2BePSxDhTq4eEsZSQQhpdl1ion9X2UepBdMokJAEwJRoR21+PmcRNkH788nGu
LT96un1pTI4w/53PZWxfhD8ESBb4rEKKz4ZsDDGhKky2bP2xZY6CmsdLV5/XT3xX+iWh0ZBmutvr
7r9WFpAwEIBXlMjGXBeO4GCPZF50WXqaSm26yn18k5knW1rFwJiDLGQH9fwslSo/wYVmq3IS8Hrp
Bew+Ap9fbKAc3HiJzVDC3A4c31oLlJwHfvhHRCjVJqqj7ahn4KNP4a2KFB/RT9AVmTbsvVfGqVcV
1hExOyqXUOwv2OopbucCaIw8pp0szawFPJz0LPjlfCnuMKn1w+YTbOIFEziaB72BzKlSC31GlIwq
2w2MhXiy0R1B6DaMPgrJjOGbKNxu5h0XcBwWWb9xAJieFe1DfKssQ+ZGkxRWhWYUQSiUvRmeuu10
KirRbTQML5JTyTXxsbzowqfKij7k9x7oDCNHB/u9mEJRk2ydxL+PWKHiudwHRz6uqEE100wi4H4l
Ez4XgK2LBJZDomalyyLQ0+Oa7NyqT0AvK8+asuhWZaxzdaMbQNvPBXwhQ7KroqbSu8vt4i5Jv5H0
N/0bSh6ghsC6rLId6GdosUMFjpjFqVxmDzuDaR+rhGvHku8xIvZfKT/Foo5jKPMFwnUWGbwjmeNW
rQbzJI3t33ZH0CShklQCMsF8Kd3Nj329lWAtS0WB++cy+Zg7C+T73BXQ8WLu9BjgwseZNybEDYrT
pVajZgwVHn9v1HYamJKHVBMsamUycrfmj1vA4aKEwFuSszItFaFV0w+IH+2q22ppXFMJx3d6IG39
7+LayV3zXag5gELBRBjAJBIL5aSF9xIHutxnWCHkEAXN9mFfYJaUVKs48vYMTKEQJgCderhiK4L2
ChksLasNGYnTTvRgEJSsBVDMltEJinSV0pAvVPv7rPruvj/UyIQRzNHArBjwaqMV3YjsiDUX+vLG
XAGlZGtjYqTnevc4tWYTRH7TmGpfO+8+sfYjPaQAs2dg0eEZ1mKYyA0zewyYQw1N6rfHPxJf/iEq
+WRxfSHdjqkDWRlL9jQxYO+EE6zKzeFx3Lkm1FIv9oj/Ap1M1DKtTmd7BbSHny0n3Bn4X9WGcaSp
VttVKnFGi9PYptdymj201sYy6bMp1HKeJGwArqjVJDVmQo8h5U6OA3hQQeWZIgg/6zAWIiTu94h3
qRCPYRtRHQMY1HZwZCgC1i1vlzDUQbIxC4ytRmsq74gfHIS8eFs7yZBTarAOqVWeA4hqg6dc6SRK
PQlM/jHYgyD94msi87y802vtCdcfVGI+Pmgx2nfwzxj2jCL+Tu39nQKUDAIHhRzkVQv7W7ZzQYEz
NZf36sMu3mwFPVXesQwM5GYHg/bd5JZoJM5SUoL9MWp5Op6wPmG7uaiy7H0N6AhBEsLOh1f+Itv6
Tijr8nk63Sfvv3EPZxkkwAsq73w09vDlKzNq8VYakU7N8rTtsvIc6fIaJE3dqDkhjP4bMLZao7KB
Vsy/53ermZgvyx+IXiqpiFYlQxfSYufGQb3gOTCCGLLSsxTrvOVuaj92ZN0Nru2sGSouVOWICMSB
8MeUdc0HLiu54E5OslvjmPUcxbIAGFiMb79j4o2Nd2jXQSUQFivZDzlnc23jYX7s9HygPYhxzxH4
8z24hFFMMOZ+hDmRns2RnkMHfEdH5Ahm78VEWsdg2hgUq/9a+oj5R1c9Jz1Qy5fxtlWTRy4V0Qq0
MvfdLLZc2E9uZFrUaBZR6u/xw5l4cptZB26TdQ46VV18g70niGgnq4EuSn50Utapz0dSkez7MNpj
AJS0ZerJHAG4RV9gq9RjvfI+lKpLTCss2nJ/9X7sIHMDNYZDRONtKS6N17kEUbdtPcLOm4sklfDH
7db2922kqw7x270oLFOlCEZNanmeG+E8qteDQBRmSe/K07YmN4i04b9fUPkfF/3thn0eC8Af4JNl
zfWlkojzJVuxlc1vh/s38nz9yLigI105FmZNAd/FfTtWSfJaUzAR6feQ7KgyXaMwauCBp927GtsU
20cY+sMygYk6nBMYIicFmwDyfIjRVPtLzDLSgXt+8sx6lq9ozjpc8qgYYT+gKH+gKn2cpLWXf/eo
dP0rSRRlrCUg7z7o+cmQILhyPRDEv3aZX0eAZsJT/xscsRyJuYTR74dhfWApw8nX749CeHkHYBXE
S4lThtLzdEI+BvodI0vZWtKvwOTRzUQ+YWpDnfGF9nSRRObviAJREzlmzUnGvj39+oiJRGz3gbJq
VHcZNBDefvw/HEibHEfl59PymVUvxSnYoVIvS5qON70XCJb5D3pUj9A+AwL3Y7efzzPabMffQelp
2g9S4gzqY2iZ6Z1O+peQo1zYl602lHWJCW4l+ujD8TnsuSe07Ug9q8KXBq0Kph30Bx2Bhj9PVqcv
+LtlCzYU4idTBS+MYgSc3+c7LENbs21d9nzBL6kVPR8ixeD9sKzeuSMr1eARJ3xK9c3TOxj6ZGMA
x+/9h5Gje3VGL8XX53qZAdsMLoUPmw6wDljVFbD6PcV3kKS4GxTnlL6iDU5nMu9Sl0T5X1B4LzZw
ynD+thHvMrdDJhfSHNxT7rsShiy2W5t9Pgbe5PU3w2mNleUDB8Bs1O6B69KjgRW924kMLl3aF9EV
DVeJeqCLIrwHK3KdJcs/dmgq/8o2qz9cERo1lu+TbQn3yiN0Dxjfxej7hsBLlIChVL+C4Lojd8dj
O6euO/1kBMbe+qtDlSVkj2OmorpUL1NpJpAYSXWxH7F9u06i8ZVRb/tMhbsluinxciPOqdhGWxxX
vStlr2MXm26rDKwI+ey2X+ht27cfTFSE99hJfFghUsSxYibe/SEXHm8nGqX6hsCoQpcM9EG+Ogk9
HJEPdp482R9q03xZrElthg4R7O4E7Wj+m0ZrasKahlq+syL+zE5RwC+4ZNaBLeOa/m4x42nDUCHk
AH+sRBFJMP7kLt3OyoTIPELKokWrPo+kLo/+6UdtMPRW3/jUm4WSSee4yY8zNvAh6B5/26GW1bG2
ixJX4koGy83bHzVfaJyKf5nZwKpYDHxuYe9T+Lz00Q5bk1qmEccpJwaTjobJZ31LA8eFE+QXaTBd
F1eQ58AZJCrt0Zk/7EDdz3cbx8dTD8w0ZSzigQk3reBw3rbyiTrnppNYupt9SUGXcuCvyxBxpY3D
Rn+4KjXL7jroxI4wrJh1ZHBugmnungph0WsVFtudx1ZIJqMxTtaBdNM/F4ttqxGh2OyR5lkU7vlU
qR+kUXZHf6ENBFOern/qZOZqkWUsTuM/R3Q1snGG2XEHJtNFrCZFpIMWQ8bgf2ygoVnbzWB6cw1G
OsKhbdrVFkp72UgwhRv9kAi8rLI7GVSzjaxgFzyp15rwS6fe6d91f8mod8k+AoCwjJ/epakNzNY2
Iz4HtdvEn0AOKpiKS3tISfJox63TGIZA6oGG2QnRukZD7yPu0Kklbwb3y/9Voi3lkaLJlu2jMr9J
SZEAyH2yMZgFQMqDcAnkBmivExwVLeuXr9DMgkvfQnP4oXdSM8gu/rMXeVqTAGi33ft88A5yAzU5
ECgw8+Z0ABUL0XnkVtvwaktnGA6xZnVAQfeTojReAu1P/4epbFu5OC6JogASLCNHAFW3nnGQv3SY
572sJc4qZNcpbr5nFJxwrtdFTrvYlZ8PXcKXk9ug/QxMjtZw+tFVYLsxSBtZIYuoUVLdioz14FS3
UAvSpIinTasS1JOmCSyUt0Gn+oD5ikNrWVKopkSLWSei9esnWF+czlgxQz2i2/zFnFMcql70aIPy
g9icuSnd5civhvIeFggeRs4UHDxSzac0/YyeVewBr3cm7BU0FHzyjno3IR6hjhJQPHwyIMnHKdQ8
Kua5tBz+hI4h+QyZ1+/Ix/RtbjG6H9UEdbSjJs+gueCrnAtFLcc5bc6h2lfzh8Gj6xZa8qMjmpNM
o9GUAsSMiX305PDSGSlRgXz7f2NcWL2cKUZk8OhYSmRvqGzWsZxUhJT4KaCJIcZ+PW601++2NOEa
n9oxYpHTxc3FmAxEaIhPgsHwatE0PNFUkxhwuvYQACLvs4ujaMa2mVpMlyRztqVrEOQZQ5zAsnGl
DR1aa1cdjQ9kLU+bWgNYdlSFF5VoxJmKowH2f77wpX6tIYsUSde9OzMyMil83D0nTXPOZZp9/QoN
/pRFLJes8nzJIoXNhcczV7vxFSgT5ioQN0e4rjIe6FfaGKkL+vPQ/Bmi+VfLkqUzGmYlZ9j4gtHN
s9Q7fNgXo5kPKogRSvzks0/V8UsydkDWxEMUlOfPoqJCgf3R13KvHX/U7uNyqLu8F6GJZZurHpJf
CKVwmt28F2XvNP+hgtTf9HWE+0JIKvW5CcYRSjKYkZ4dTYVey/g0CejYsJUMn9bzyCkhOMcRyVFQ
7Z4qUuxNVT1Ossl4BOWXqSPT2g4emW2kUBWAhfocQhFi21Q3cHzwATB4o+znsKDPLPOS2dzNN9CB
xZBg8g+NT9rHKHaFHOOSIfge2bfhueCXyUqnlDB89O8Q2EEGnREl7LXvJR1UkHjQ5QMEodrzUovW
+LCHZrSkMDmcvd51U2ZyWsSaqOB+Ez7zwV19JIyxcvZlhREV0CpRzqHfI9dFhS8SRgyVpdMUIpRB
kj7DuuTsR5NP3f1zDnLX656ZDT3EwB/QQKRpPcxfw7Q1K0QY4g5sKswvWQ3NqmGv9pKrWToELoBw
+puPMtcBlTL5YecDEVWQlI7gJGVfUrHdyPTq49Ic+HYkiBfM5BjEP/zYeTewtdfxZW0G1nF3q5sH
kaEPlfLYt3AiRk4RIeD6A7UbVhNbtP5I1Kro46VCUWmUIT1dpYbQMYthEDI74LUpo4rUfhIjE54p
jc25nO0oeKvr0/5pr5D+dzoKsCMuhZMql3WjihsLu23ihFwDHpoxuAbDQ23rZ9JQoERQFmh+2/QV
n4BsJ4S9AP6v5o/i7JcvbkM5IHWHO3/cHVRz+gz7LS0ALoiFO5ftdsvs5M2mQzlwp53mXT377tMa
9vtHq6LXytxVN0uLgx5F/1i2g80G7W+ahhsI2Si6kBhZ66uNNawy20p4tAoDYupGxt4P2+EthUNE
FiXzfNZW9ROSvUG/U+n0GcrKdDavxevrQDwMjnxjGCYkImoTTVjtU8+SzIHgz92YyIMN0/CIHZwB
cFBy8G5Z0nFO9BSUIGj2DMzogeOikk9/SgjDtLYdaoonhVzESNQSZMFHkGl5r/nL6zVO0IXwuD2a
xeiE3vEAXcQE3ruHniiyFO5mah74vcnU/6TPeNFKiIEn17FKNgFsgoPAtY+5LW6aZfcONOZY69pt
njqQNbRsiT5W8J8jY+ohCWZPOngTA2PgwNABlFE99lUECeHAP5L2DRoGPmQBy7FMZptrCj/vCwKY
KJ4Ch2dXvPf8wFnWUCpTagNbmcHGjD1XBK7Hro2CW0p4ASKbZVbvLbeR6wDnTNSCR7CPpntrASZs
PnmxkbNSOZo/rHR07nqiPqnPDZ9qqyuFqV8Mwacb0eiFd+1xXhundZuBc5oqJ8rkcI/8erwn/jYo
ZO6SYXmVWMrwtiYRy7CC38FAaf2uxlQOfKiEVwCLoLA+Ufifb4WNRo7i8nZePwOsdcuwHtUXwETo
dBJLpfKkaVLDuo4kKSkOedeP9jtNZrcwKTxBshOQV7VBxrTSTUjRU5muL0W6vX0bl5yE4k05lGpa
BNoOTNwBnvhmBaKiPaBeMsIHj9v/i8ujSpLfUdtKd2KBn5Q61wnyvKW4hjeMnnUCXGJYWnsdPva0
jpYWokC3ugGkhYN0Jx9aNkVoaCQjrVpV0pHazl9CR1CNJiqQxhf4MsIfcJdkmn2GXzNoQKeLRN5K
JHXOmN4E2vvdSkod7ClrGmDQzuB+YHQ9PgQycAhYcgO2UZxMoOHSCqCV69UBpZhfF5v2wezChG9/
vn5S3psjT8RM+wA+yB/tkiMvqx7JWdAHb9TFcE4/lTMBVW6k6nhMdm95PDcWSg7Kbxm3SfeF4UUA
XvdlwgjZn/e6pw8CQdNbV8UmHt7zbbNiz8UjHZfbh3oejnSmBLb3KRMhpkQYGApVGWq5MasJvxFw
Kz2qehwKzr4DCEdENaufCmqIL9ypK8pu3/VQkFMa5ZKHpV2uCrDfnj+tucqUS8Dnp7R+JW/J7e/i
WdYpUSdrykrB9xEoKAnS7XL7Kxja+hhJGqr3YKNUhEq4ieLZ92YCERndHV0jr440X3gDcDNgzvxt
hAC897zPVNFdkcBpi9ZdiNaJ45cHZqpllwEuiJFh2wui/YqKoQ1NGBJG5cd/jspaDM7JqDO4VsFN
u4NDpV9IXvUZ3Ly/FZpsPs32rwRbFRAatGa44pHTmVy1jJrmDMj/GF90S5bc5DinWRvAcH4IaDzV
ySUi/jMBKGkqkS/6f3A7FOuLQcsx5JauIL+FhEcWNUhiX3D/bAiNu3x+G4SCkgf+r7ZFyRKMSYkb
XIHKc0UyyiEyA9oClIsTk+5b+GAaiS1llMHQ/MeKiURYb5TDSvIgNDTMSBw5cWzpJ9xRtqmUpVSx
KYMZPl+gYxlRC9gUqVmg1uOPBWHGLq6alyu0WTlLJF8vAxCGzTUK79T8oWeWqdAhrmPfxcddLxTF
lfyDW/S6QfIg6eTQ/TP9mFA+E2giJ4/1KkJpyDWgIKotyIHKRTV167xCU1a2gfQ+vKZXXgMFeKeA
5I62LnO9zV9N1inlnQn8eID3c9LfRvQZX4WlXWvCSKNKPnwxID5Z97FTP/4OCghvjjHe+yeIbzDq
kWEeNisoQ3bxsBcAmnyrsbJnwd6NoF+g1duvlFv6X2R7vnxsr7kf0hNJ2d0Sp5Q3wXp3EzWPS3rs
+x492o7uyn6Ygk0j1QEWFu6yvppux6huDPmregirwmBtlcGZvot0sB9kjZ656c/aD9EHFGR5PEpL
6RRuvZwNKuE4gs88IoaoJQWcnyNC/XXBmHBea14Hk4nxB1MRLBurUjMbdOuPqUYj9+kdJ4r34rx7
K2+tcXoBtGSzEPqHqCSlYMclDKraoOnfnmqR8i272r4Ozm+v6nZXqFzI1zHPtgXmy4UNuLLCWQZ1
bSk+toPehHBjee6Yp9zU8OdCFBTyd2ZkURwgN5WaPAxB29sCYJ7W3Xu2smvJH6jDmxmK8nNCkOGK
eiwEfTuFTBXZ2UXG5G1PuOx5N7fgPpEhZ/bwLshau0RAKqFN375NtSW1MugUDdXKo/YZVVIve9dm
TzNKHOTpx9cWJrmDscqAX/PYAP76OqvbL+g0xiMdske3us4bZxpom/5rXFZmjYpeTT10RuBJV1vV
MnNw7jGuKwKOoTV8DO8vF6qBoRm/88l3AvVLruzp93wKEbxS5KGwwgJRJrgKA46+IEVi6Zzj82bv
I4UWe6/XM7AlpRWfW9PhLT55hMPqmE8dT5tKAAs9FBfK0vWJG8eGxqMBoVpyVjXUHSAoClc12Qj3
w4MbhymvliEpy2UUyWlj5dbp3CCJi56zURZV1g56nvmb4IbfxCfnIRmIwa8wxHmrwSYMwpSEhG5m
8s8234J8RFc7SuzW3DkMQp41fOI1MzKkmSJNjOiGcHgUC30hJdOfp0nBylr0HcHDO0vOeAQeD5Sg
SSVyczYXm6l68JEX4vwb5o3TaFUalWyYXlyh0Ap7mUme8hH3asMl23+s6+I+3G3WuzZZpqErkJG8
GK0WS+fFcG3IAM2BIbMQHTIixhG0joY4h9ILt+I6nKoT7ltAn/Ai0I1pADt2KobzWFWSuvF4OzZt
7VikRRO/OftM6JchC67uGR/Kc59UGiYKoFFl8Eve1oVfD5Zksys4OU58AylqCZL59z5nyCECDpAW
j+9ZXSBWt5rp3RI40u3ghrFpEOBFlzugw7hyqjnGIjgw7pUbXmXQbY3D+3f2BHj8PqXi6DDedVxN
Lam6uDiu7BQ3pLvqdwGxegAyKckjriqBswMpHuDeZyFZy6LRE2YjeJQK9l3X7NPH90tnW5wT+wkT
B66CVywnNxwreL9S+Euxa1MhDf88YoAEOx1nAVWKv+OAr1mnrXY04FaTN8rfPOB6oUBjqFb8secI
+D33A/TS9Yh9HxpGg7IFWL7Kj/TISssW2FIV6Z6sVoJMmtgRoZwveLFN5T9fNMziW6TlqNrSKQYQ
qfjvURJassVMVZ4dxgeqXo2E8lE4Dpb88ma/Whc4J5+qMjzbDEKSp2lF9AYU99aM9TQrdufFF1lZ
/Dj0yRSo10Y3wbtEaL3D82X8F11SPj9wX38/bpyhFf9JCXEguDElIwJdPchSN5PocXsJk7Wq2nlu
kDj76kyAJ4SCN6ZP1SGQC4Cvok/Rf83gCwfAro8RAcO93JgqERINYs9z6+BzEl3W04Hi1DksQfHx
EweuR6Is1aP/irYwq+3eTRbLKR/36cEBtKsRDc10CODQ+ycwZZCodnR72rv68Thh9c5xm1j2o+U3
idqaOpASKhCPXUp7Gy5mWxW/uuORvNu1MDcSEOaIY4b92kA4awdQKxMpawK1S5pjkr3linmWlkNP
zsUEvu3ACa0TWzFVszKcrEarg7/XizJLRNrnyitmToAl/2xHKilCpXTVrney2FTlb1xYvW2Qgnoq
WbtK8z03Iq6Q5o5A9d7yl2cHmw1VxfQb4OhmdnirbWnN3BcLVZWkBhtJ//0SNBrbwsIKSAivI+Nl
9U1XTQcLAIPghyImK04ED7eOGz0aUA2Ib+szMLR+/uANa31A6RJcCSY8AG9STvGsSeiUZtNpEEP1
MFP1AuhieSsBdRk3fokpsm0mxA/JPo8AjZAIqwjU7NO9nDKZ0b89B46Zgi7dkIvIdyJvUe0SYmfA
e2hLBS9uq1gFIL5zHmRuceL+BIFFE9ZXUV/XhySwNBCyDJ1MEh5b8juteqtG8MC9/tEPy46TTGNB
eKMkbkA3GJDZ5VBMW4X/xC1f50EFAjMaLirYvh4RSAMIVfyzfJuLpS4f6+SRq84z4hIAj3eu4Ewd
X7mmusNUMAYwFN9o4vCUYKiYrnF4s+AZlITUX5uwnJLQXgmbZuhBjPi8LwPNGmdOpEHTZGkvo6Q5
8RO64y4bvJDQbmtORd5Jlg07zPU7yiJPXk4xqQpJKcWM0Ej1UINKIxZSzsqID8RfckFUpWR0l+pz
u3ihBBcWlP+IvH+8OS+hKkZ4tQvgNMcBkYjPaH03tBomAQHcg7LpLQZqTih4doPvXJVWuD6w0Yc6
DPX2PBxbc+szGkiFXqX+JD/yYHa6YABt+suDQwBjKDRBe0XnpbEIn0tihxqNc4O7jdDMseb7SAnB
alm6AwnwDAm7kndd8HgsP3CbmG468vsPGVbW9fHdz+mQtz2LYB8rSN6BlZSe4r8E7m0a+eyKDDAF
EeuOq1Z7ncSyuGGhBvjGKRK01i1ueF22/ITmItm5iawQSMCLpjrjvfOYttFwbKldfwyxOgrlIGwX
mEjg5N+tA2z3F4udN0Oiex/s2IM84IYbwz6//bd8u2VNS0QZ/ys4DpLWUWeOTPbhNCWiWQsCvSIk
LcMxLU/UBKqDF/ROJRuYNRsQ8+hIMhgh199zKgBv7FypyECaeVBcC52y3vmFXdBTr7nGdXkdyNNe
k5aYoo5jlDkvimjADuMQvABmcNqfCIyIUa1cGfsiO2/XizfbsSMdFeRcBTtGzE8K1LuMjaHVkAFQ
3Dic+hG5YmqCuv3F5y5o6dKKYpNwLf1VJf5ONGky19nG5FjmCOcEcUji3GT3KBRTwktpTA2ELyjB
JLIyfAjTmIW7ykO6RsAVSVSrbwuXQvzhW9ol47Wp9X6S4WQ3Z+evvtAe/jSdPVgM9T5I3T2ZcDmg
eWTh4h59KBJqx4KcK/Dmn9xDpqNjQYkT4b7hjQQ2jg00l3FT5VjiTvXJEsU3CQq1GHEi+FGLZKky
zzTXiGQd/3ueGA7Nz4uAqWFh5cg7IMEExvqTC4zyNMGOqa4PtQF4Iux0UT/BUSapJu6EGFzk2P+T
VtVyqph1m7vSuQA1TRSBCWAhdUw96I7qSpoFIG5fiNi1kJtiUmxlH+wWKwvBLgRv9kT2PRmxrMv3
DheSmk7EEiyW/kkjG3YU2OGygRvziFqe9drYrzF9oI8JCP2jMAaqRtnng6Dl4u77qBJLHr3rShxC
03BkO+09m7J9SXlRNEWEtc0If7nsU5xqewGFxlCd+u6jh1ddERYa/CCmAGEmbOmufsXn5qKZaICU
QY8o2h4ES5M38+F4aG+NvoaBYMEQYBl9T8XUqM3TG9a1dzPkdXbPQAQi2AjtcjfTeX3hK1C7NDPS
BhUXReLUp/SCBdee2cyQWv5wpLvzm0fAeHpozy1Z026jfXXVYaUsw+g5/nQG2XHCaToGey8+OdcS
NB214tX+iJ74dZZezEQ9zzYyluVyENHy4yN8qHwWNipsEO/Z5Giq6cZWHlGwPFTdLsiL+X3PniRv
LVjwl42AWRuOsV2GapUtEz6jmUdkgL3Wzl6LngPzyUs9y78N7uJKysIsmZHYjZnqNToH0tDQIy1c
wx40Fm/U8/kzjTbUMqNPdhEXmMhAZbS7uD+LSXT/sbJTFQyrxGCXYNwTMGXrOSLdmlPo5rF0BZU2
nce00zf832Z++tIMuNUO73Jp/VG/gZxufAtXoyyHsoNL2AkCSo61/50nEtD2M4UTuSogO0Y8rCv3
dl971o7Sf01OL6iaIE4wmbggm+ob0rX/7ERSQgdIKcw4BmcPfyMS2FEz7KWNAk7GRaM+pgzYflva
L0szOGGFhBhs4q6pWj35juF6VMeDLU+VYyUQbSnQHIA3ik7o/znf120Nxi0Jc/kiDcsWpOKh6uqy
BiRcI05Vs3XKER6oZ5UqvoxPZd0ngJsrOD85uAsGSSqcpOwQVf8OkaCXbD1+bbzF8uDph2mWQxwr
qk8gnBpvlII8cyZVm95sbsf3OiKhwtIJTu01r11dR+T80c/gPKjyFGd5ewcbWtwD03oFM1wQwSWl
0qZicoZQ7Vq8Dh/kgEzbyTwtf3x2oZVNIUVrIBRh6DPCqvl6Kt2TTeH9pD5RxANbQ/aYXBnSPeFb
9X5Q5J1nYz7Fk8mK3m3VaWDBRjmoUrGwfR2UBnZahq3NElqA7yeC19NjsU50ewOhzO5XVFV0dQEZ
cqNKk09JozpFcUbyuLZ3zXJ6cGtLemmbU7wCCfohYxO8YNfqQgxdENy7SKXxo3AN8WBcv7DnW8ph
VWhB6TOlXJY9LX+TM+8gsMWaY0kWJWnVIX7DVW+Dfxw9CCjkejpaVGCIb8Ffoq94o8UrHANVY8F+
GXVLmIYmew2q/EXlwWqkhJ1I8doiZZkd1x/oN2INxG8Hx3Mj5MTxbbhxpyT61a6fxlo6aOOq7DyQ
ESiRsv4Ad5YxWuDUve/KFFi7CWPQP0zy0LeM3U+jQbmVXy0jEGd/IDqbG0LUzSE+ZNI6UcEpmGdY
wkrru8tQYanxcwRXuicbCxgqofbA+1d2JSlApYpowYZZzEvgTQii2NqZY+r92IiqM1Fob1Y4grwi
qgHNTU3kUIPbOXJ6+14UvRVtEgxLw0iKMBpj8TQwdAmAiaP8xDrGmxsQkLGu6mYWWJ0EnpHV29ve
rR524m/VQKLHm8mhJHQGXtq0vPL1X+h1Wibk9cxw5Wl0M0YJO9Fl2MJZ7u3foHSY0uuKMo2m6QI1
XwUaP7hBNHzeqcSlLaHjtoZRUfzxwT38F7jTC8rutxrB9rsEspcISLyNgJcpVm5dlFholMOP/Ewc
y5akt1NmEGuX7lbfjsATgy6ZJIAEyFym7JgV1WVSxKHBUtAgvw63eHQLuRXDIYuphePg4seT9FSP
e+IdyO6sujeEimuLQCss6eJIiqAyoS5Kp4CgksPjEhLoqhjC5Rte9bbhEQlzWQVUnHrxOCzTgsLv
DaTqbEsTQNqvv5IZsTY0zcGXRKBTT4u0jC05Gqh9mTlqC7VV0BtKZnpwprjlIIYkfs3jw4fhuCrp
06c2/fNS/VDLdYrN87x53+A/Ew2OKl4bhgvpga2mrRUO8it48o14SoVKw0klhYJq4nGEZUVQRR4A
jWcvYkj/MiE5SCSW90yqQ/ZD3fbKaSo72xHz8ofukp6URw0K0N+ui8svazn++CYRJExpJ6//XmVu
mM1szJP5tAmmdLiaF+4B5y4tCGvDmzDtpUoV+vZdvx/zLg0xgcmQZu03ajsAQgEZjykbljQ7NOoo
rDxydpxO4DpgL4P0/DqfvKc0SbXA4kROJAuWTP3ekyUkEy2JKSJiTd9c8wvH+Ka/hk366rNT2hKp
e6l9ivPcXYFdX+JkArur0c2eLv309ka69ScTAiKN5SVw91S326x3tts1FWyTzxyHbMYGu8bFLy07
udrTnCG80MUEH0i4EF8Iemsf/HSwbLYFG4CUDwm5taIx3H3R5fwIHg5ENvF17t3lQipJwWfCeYf2
E0wqBxsTlbWQ5ATgkiiI5lAkq0Dbz0V1NtFT0S1Oo4KzuYU9Mniad4v0WyqYb6QbWIPJ4Q926vHp
24Y5BU2n6ykb5kicccPos0J6OkCkM2EQqQl68sDBPbbKiDYhcgWIFmPSm3gYWQzvsid1T+6l6wiE
v3win5OR/PDJpba/arD/PQNH8rdIDFiAMAKt6fnlaRT5O5HDEeVMLwS1WdDngRu3K88WVw3lml4Z
XAfuWYrDoi6bfLgk6YpVuCLHMZqtM6C9sqwQdWIoSBnS5udYSubO2kzNcL0P2/dpEi+hD4FnVgF6
BvUykaSyhxGv1kZJTXNZtAnaFQF60AgUv0OQBSAGaL/GV5kW6V/XuyVl23+eTmII2ejbwuanrSxc
kciosziNBrDtUgxm3CFyd6W95GIAflxD8UDMsnlazqfB9Hvjak4JQUibeQgSBfNmMOi0wJ2JKwTo
THtGAAr7msCRCzBEjfAmgIQnZ4v9LRt4aJHL/otmFR2KOa+6V0Ppa39Y6Vng4tufRKlj+uwkZ5gG
jKGGmy5oDyHWfRHVGVWOTTdgn/YlZb9Wb1enrrvjp5e/E+JFVbnYZ9861xNyBBYMtnrMIte+Mxgn
Cn00gPR7lz6VHE+vdo7h/sR2F5eH64MWZA2Vu/8eKqaqP0nGZ1cLwzxTV9I1oJ2fa4HG1VSaQfue
oVEc0+fo1s+ZdP4Xd/3XfMuxswqsc2e10Yt2LMXHuTI1QvIRpKtSAKv3gww9z4XIH6JU76LYDxZa
vU4S2J8S0Dgw/yN/m754w/ZMOJ2jMeVGEkat+7hpkvnbNnPRRxsCYDfy6U1sM66iIF/P1KPWkLRS
Vq2KFpcTaPRHOT6/cS6SXlHWONTZgRTpbR/qWx51kx5FP9iqZBVBLaYR6bHTPq/6YTJ8EcE2kNL1
xKf1gXJXc1gUxrwl+CLC/EnZmtmHqk5hAudoUAgiEVuqCelLbyn77GiSRRbJ4aSIIhidbqIkC8il
7F/T2ltcGB8890vMhkd3rky35vtlr9uGz4gWnr3h41H/4Iv+LbCZcXpx+VOaloN6QrTL4pjZFCMz
7FcKdb0y+iz9+MCEgvPM1exw//jT3eWBxk6i6keB9yq2eF5MCc9BZ4BK8HrHE6nECll/zGeEcB7B
tenYElAGDrXxdMDLTGXLWACKJviPP6Hy28Bl6craHFVdJ7DsDEd8kDLrss6SVaGsDyCYkeqV2iW3
1fyDvADFJQP60idELTS5EmZ3HTSLjsFx5igpCOpl9WloNP68efGM/OszqDOW2eRS9WnmAh+OhMFK
h2G4BZVZOcXsXQFJu8LVKID/voo6XZnpld+6eHdt6pssVevGpQ6ElmjetnMWLBy06ZcH8/KHLyUF
BLJ1BaBVhnUUgfJBeLT4LYrEYnAvvlnq6YJXBHGAhxzpPVbKhGhxiQg6PN899EhH3oXD+XiSrY8A
GWlKFd2zAwsHcQ7LC0xYEIImydXj73rnQKe1DnoR5Ir8kwOVrEN/RHSZ0P7INLuKASQSI2xa596U
O8KT8CoO95BWE539gIXF6mU3AYazfCOu5GPyoBeHXwFPSW1CqMo+oW+CcQ5JJzmQA/Md5+VLSBoa
32NKyuYhqx22lMAPgtiJhjUW2morkE7/LhrPKBjvaWIm9t7l0lQ4ZXGwrdZGkGY0EX4HTaMgTdgG
6jPpHJCXU4yIWcaMeXp/a2Gu5D/xj3h2IxOPjpSUKxzSdVN1epG6e9yR/2pTgqKG8R+uO4thS4nY
wTkQMHXQGj4XhGY3H8dVgxYWqCTkU0paCw+sYD44hgGEF1zOS2bICozQP6W0CE4uVkdzrGgxvMxq
Otc66ziyAAJAm457UHz90o6QBpt4acqumqOEBe06iFWAOL2MW03YVbux4a5iGTQ+1hPffqyzFXL+
C3iGw1gxk3vs9jvTyQd3EePcvbJGNFlLdAqfzIUAtEnhwJavWr8jxmnlQhI92eo34bgcTd12irDl
tHXtJO4ERYGQ9ETMJ6+NyqXvyqTFs5rXTBffjLPy97KOgiCh7nyWw/9qOqPalNzDZpVbHIuN3Agy
Rbumi7NxX86SEeNqH9MMCVKU4SuHuujiyl9ubRPXGwoKHv9JEdErulzaRGhWWzfAyCoUxmpHGq6c
LsZ+eSfgOAy/eFnhExXxWuGOZdbjyW1k3jaCaCHm62dHLNi1C5eOxYTMoXLhO76uH35I1psvozLs
J2E7pBoTa5uPm8TR8EVUx7tqWgJk7iCYIjB/2QMuaki3R0hpuKOWfAASJxvNN2FlLNFna7s0b1aU
LJXXGUUdVP698EARAIBLH/pLBTsdo0fEJPanV/nl5w2zfMjccvMUCvJKPMqo+nge7kpxsXHjh3zs
oy89IDHe7+72yaHfRVQ3W9lciq3BB/faBq5B65ep0Pl7OZSjrJxFoDxdAdtYu56ZKpHRYjP6CkJc
JQHHZaBN0Lm/Al6a1O5PQg0aemyCgm/Voso7+eZbLdfq5rbSVWKH0IbvilOzvhNwA53Xnm9D9Ul7
T9+D9HqpfpJroc7hTmi30Lcax0en2u6K/YalyW92MTVt6f/V/4mnAsaA3igQzEsjKJ6aNC5Gx5ys
IwDcIEqGArZdMMhpkGDFKTG4ND4OPz3G5JijNVD7fGichLnTRTfTvVuHqmY0hX6CNw9LxTXXkNQ2
wj2idJBPsFYvMus7ok2ARBTsUNGvyeNF8rO7G3ChD4YNh6TvVdEDeNvBeKptF3KuRW+4A5w896Hj
uzpVM37b9+CwB2DTcsuMeVdHLEcpOLmzVIkcs20dC/ydX8IpLgBbO5t5jfuEv2l2aTViECHjBPBX
gvBu8P5xQev5XA2IT56qYyRAtC9xubf9d5uWZSyTbpfkbnOMyK15PlAsqdgw6eUlykUG5NBsxanl
7uVkeqqMIgcTqm+0/HkMUNg/b7+z6hXCa6nixGtIMwOaZnycypEk37DD5UvL0pVo2tTFUnmgmN+f
AqUiSTbHh9NJULlNQTX5S8spCaoEaCptgFpLgHdIXizfJA7I4FUUElswMeceALWOggABAnB5dpwv
dAgOJcQwoXaokhZ3Bl68UAVls+a6Zrd+/MxSH6Cws1K3/ySaxbgoFoZ6+DNYXii9Aqpqwhn1u4vR
dWkmznA2n+fGpwlpQOR1+19XUTK6VyqbGA98pmlYO8Bq/2sl5kzlmlDu+gDxZVyzXatNTmtQoX1q
iFn7LGoq2fjFycM24Aegb25Ulaa3tmFBNxITbhQL4lCRLnmEwdtFmNh3Rgy4qehsZH+urVQWb+5T
5d5UArL/A4fNo+mRPw7jJjuX0+dJsGu54Ot1kglLQQsysrdtlNf8Ro5KTBlu/HhtZ746OZmcQgyF
9ZA+Xm0oNn2oJwyKbTLnyXkcMm+UdPq6ImP39Z32tzJuszdfPxQGonx5IS6SGz+zOkXcp8o3pBOP
CafH+3V1jZZ58a0g/6fn9SXgMQV2XkHxyFVlvWIf4Pu1lvNgUtkByFu93j2XvElQpY2YGqupvRJN
+PsMlvS81vX1UdkkXER111K3CcPKhmZdFmGZ8hLrPEOgyub3BQfHT2txzjol6pTOYTuxDpwAzxxy
OXp0IwZEdHsCEYa/QnsUnwj3wUBuwv/Ucu4jtTmWzS+CXTuGthI0m7v/owgNO/xRifRa7tt1b6ri
wruRJOUttrVHz60AvIF+rISu7Cn+GG2otX9UZIhEOz0I23uzpZjTPlhF++yx5p461nW5okUebE7M
pymv/ssAvJmkgA0IOp1f3cGKQmGkWkuEROg7o1C+J0/NPd5aMKqaDUok0yZN4J9fm1CBn9y8j10u
FUGllO6cljJnTqEyQ7LBuTJ2+qZGFxY8D3vbt/1ZeLq6CAPOpF3ACpFRmORVIo0oJKJ2jQUIgN4S
pgR8oYU4+Lm2oJASUsEE1FplzKevVWBs/tcHwcKOiafM1Ca5RrL4aujhNRbpagOjLIM37UtOlL5e
M6oTD1eqypiejv22/b5sz9ua5y0pmSFjDqAA3ERd5zRqFT4T8sUCFfMCjmnR79RLaHxTE2GEavD/
ny2njgd7zYS8BQlpDCDrqDG96MWj+oHiKULx4xX+aCgba9fdj5NA3k3IYTrUlmz4k+allcI20x57
spk2tG5JcdwXuDZxz2iTwSsZwXU2oGGUyHicRKegokUNHy0ySELJEB0z1lyZeSd6Hpyk0EwBSMX9
ftlHGiVaC1AAAY+kKeiYbOHrHxTn//14DPC7LOr3nNv3jpgeaPttEhAYrb506sMpWX8MY7XSs063
Jvh0exw83T6EiCSoeRRlWABB0MLGe1pkeboZ9vNUGIOn/k2P6uykdE2JWp8aSKinkipBTqcL0NK1
83y/Gh4K+yW92DF2TJiJ34VfFFwYCIHCoXkGLsGevTDUC3isiUuD8Mx4sC9dW8izAQ9AUG3AUtHA
36hTiYyjQiFww4fS4XuyUVtQMUwlA25UjI456iVqJM/WqC5K07AQz7te84/YxoGWBohrVJAwadu9
pANY7ga9J+vi3Z6xn/VuHRBlJuMzvMnp4P7z/vBTAVDYg2l0k92vGBP+leMliKRg+acZKz3RHPEs
SNTQuSngNFQYSMzDcue0DrD1CXvoPMCFHKFEwL5s5HMT/F11bC6YiGMNMoa1PvJDI7AaDv4pikmR
ZAWvogZl9P73Yra97N/T8aIFs9Hlyj7w8Jw61XNkB9WeYlbc6N3o8O4mMYnp4BwFUt/Lk4WJ2h1D
EvO684506Z9OExtiZLzr
`pragma protect end_protected
