`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5648)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPalcIedAIZ6PpMM3qHb6Agetv8CuZwnskICkRFDQV+HXyVeNKALxYzPmu
b3s2TDnXo7GhgYkPcgzva+tV+oaLfDARS2ASfW6GVVger7l0N3nM3xW1j3GZyZP4st7cvPKm65hj
xaiy9Xi57xLEfC1KamWI3ftPZX1GNzfxwAt0kbYNnl2xb8Pm/Rbw1ZnUlJMu7Hf7J+ek6OmOtl8m
J12kpkxa+viNkU7tMrFM8zkOS0ix/MuzFI4hPbZS+BcrPncGHgRCF0qPvWdYKE4ESezezSffVnNQ
lH/OHay7UKqj26zK+SjpkX4wPMhe+SK2YFDefxkToXPvFMi5GV+G/TPFqMpyrrzZRgHJL/nGHVpL
YUYhUpDUl6zuBKlZWKduqz11Vxl4cn3S/tdEI6KdA3umwBKK8fDMqbQAccl+N5PCoINTWPHiDGF0
SqTXsSiOA4AS9vb3fvIxioeFuNWge0oyOXp0xm/nbQblRTV6sSf7V94Yy0LkW+ydIY6vHxjk/Krn
yZTgDSRvAml60Eg2pg2Ww3zbXXDbmlyX2pz2EhW0yyl/ALJWynSqN/6z41D7J8PCMAvZM+kruZCu
AWn9zTlwEuWqvgfwyZNeN//uPGDUjuZAmQcoV8TtNnffK6xNXTWzgr7lPkA2t3w0TFHHciFdCYHg
E5SqoEeENTrLuvYsdEX9uWYNZfbmry6+uvfzOnSiger+e9f8rpkE6HUA4vgcbP2PZuDuVGiIYyEK
K16q0jPxQQ2lXPtASOZtB4VfMWckuchZnoquZSpBjVz3IbWWRg4lONBAQl7olnXGJ8kaIE9Z7D9g
z0vHXaZ6HiDptcekwRGWINlrtpFTr2bujXxOwCg52iH1Mr17hfVok/l/Blj2nDSYYt0bYXLUbmgK
QNptnfZg7C9hJ5eNI9Ws27d0m/qhd40mf+OyYAwS8N/b32XBddclGbbI54TTjl2NkCBmPcJYeU5+
kKq/wqa692PsM9aYYqfBhIODUSC/T9uBie5Oxm7zdPKjHOKw4mI9i91x9l6jhpYUJW1fYeBAmycR
ooR3FClt03JFSjTNhxwD8nt72kCh17hYfVF1abB/JBO/T/My+JpKBZ11S8KYnDw0Mux78KRAP9th
+s54iRfM/rrXJRPdC1xrF+m8FkOQqjR3zvSyb+o3rSWWMJZ4o8CYwMdIVyrfozag+87rIN5ty7X4
Eza2RVNM0+rL9EOn4mRsIHVmOVBhGEBExRabt6rHqmC/QQNQV7v0c9Oq7ZQRxg3rZtygv+3GX++X
f3T5w8ikqRynUrE7ko0LqB7QOFDYjPWyO74GTQ4g0F3jbDAvkStMs+c5bKahGzc2swaQXywuGugI
mgfLQFoV6tkLl4I4FHCnKHPl43kwF2DHP33xY9pxs/ouIuhOrScTogS24N1hkNO3Ni1dzspvzpqH
l6kvDXAUHu4n0Z4NOGRggMVV3rLmGSpc//vCQrmJmBKM6fKsP2/vkPkq5PSeQTuOxIL+TR6UgQwO
41TfpokmAdFlAEPzLI1oHACymz9WobWX17TEA+bvi1gp3sLU/no7cU4xNoGzjzGvSHJ9QmwFwhwg
ARlmZZDSCfQ9dYOSgWBLbj86IfFdgUwwRh8IHya4/vsYiM4zCXE5oUp+LxUEZZhueMH/lPD5bWoC
UyiqO4UjiOGTzioRdqOk8fKHMDO9oDVWNW5GocL39hXJc2v0C/mL/cOIYohrO8aWR3+tkEg70XI0
EgDLBxIdRfNhXxuRvDY7O5X1UdLsdGREFd6Yno4Et0S4wFhrcHD6dUDCxIRi2VasiY8JfCX56QY5
xAh0VcK+8xYfYzKIC6UEWXVUzEagHC9+eAHXAZPJVJFHzUlJ7JB9nHzyEkqstOrQ8eTO+vXSnWmT
sPLV+SLywUpbuwbHXBT5bByNDv8zFT2hopMxntsFCuOw07JpvYf3J+IVx/qng1uJglg5i0AcbVMy
tq+C1+DHQhqEpD9hol4zvPSEG8N+pWEPe/SeFHGLYbROTAJIVphCXGeWIILpr3XHKuvfQXU87ykU
3//PN7qCUYEqiJiAX+rIla6VoualvMInxkoKWKJ3MLlKSveoETBQkllArdrWFgcYKCzQRBDkWgNh
e0U6Q7eg+dFHi9wndJkhjqienES8w6Hk02Re+uqUopEOW1G84/iofgXSG6uV5C4+XZFwF0I0zkwz
5rrSmAdaLD0pe/JMQErndChBA5zK/TQt6/aqxZ48D08mGLiGAkwQL37JcklCJUxvpcll/PPK72Xv
qJDk3HLatrwuHlsdHQzufhQddbZaLMo2p7uy4nZ1t+NOWyaKy/0c9kbLN9rlfcH7Tre1NxIgQQ6x
ZUnbjMyEew9qx4SPEm44h8Yk4QZOQX1HJioNfrj18BUHVGBEDPQ4KpCqVHuOGnnNHadgjDouA2aF
agnC/kA29EgT3elFgBV9tB2bf9gLL4R5lB/c0HIuVEIJp5HnnUEasjbBkiuq/34YQfgeH3rG4xfw
ntLLfHV1r1aPEsigiUPGaqgL2UDZfl06vsmFU3FxrPuaTh74GTSeNRO32kyPpjA6vhKJg0CJi2Ob
ZQ9QfI1zEAnkp+SvYEHhISEY21Ofez5pU5Jmlwgjigo2ghe6G2E8awiqTa1uVrBcIFfpjRlVGUii
SVAkX+YWCP/ujWGk07A0McIdgeaZacPRxDBy/S1bhTmzWehJHlRPuiDO3IU+nJ5zvcH77+QvJcjD
PtalJyFYOZNzFvIXkcbCTSFwcEgs2J5DCH3iXT0S9+7pcUGTUvpToJqDlthhXTLmPsK2uJqZVyXC
tj1niq070lcV4dqR0S3M1ivne9gzXEdd/1M7BSDodnM/GCAWUrhh8IjpbfyEKb3XJ8EnjoszYTDs
Z9245GC+e868xJXel5vAYhlKzVPLIET7cdbmcxZdANNYh5xs6G/CzkFfXR1WfoatTPGMEg/ewmL4
vHWNJVzG6lPFe17XwMdaBMoqaKtZHRyyctbf3JWsc7zsVGbl0Wwx29q8fzBSngiRj9+ZeQqn/z+b
zgF6FzPeWZCtQ6IOdcYEy1ikgFJCZ+ikncNA8FzbZqrA4vH7D3JVCuuppVjnu18Nr2KWr9DkSHoe
RvQLwVPvzrlXJPu+a/OmWSQ08yPZGvTI23xjnn+rIT+19iv5p0v59xW3ChVjVHV/m0wSrYRptROT
QYmLlaqT8xz2bSvFzMluuDhlczbhNDD5u9yCMDHZ9OM36hpDd7bUEaaPls01esr9KsNSx8RGViqE
TlAc+1vUL0ybTALdM4f0fd8xlBj42x309yiah2yQVHCMCDGRyzD/owfoiwo1sPnQyy/ki8V34EML
KqLqKf2VWVlxZ4CMad2WaFb+xYmqwPFHKkwhcAGzLJRioIhBFORdY1zuzFeb8lH3vyMH58tHn/Q8
UHfAFOUynDo4hO0SgQ3zyMINQ4ENLgu2cn96nUDigSs26nPsftd16KgUs091zDrIoV9gH6CjuwSk
0vccDTIc56nxMYEypFbMz4sfmBJ9fTQ5JDOTQdVhoS2znnvMaXBcYPe/057c8LhdfPGC6VgG7Eex
/CSQmlOtMn9B5/z5kDjgVjy6a0B03ZamZaKFt26GJAdSJtF/AoojbWDXWl/6TARxSI20sVOIBfIQ
4L6UgsAlmyr5c7owIP9V9rSZP2+12EXvUqxsOlAWybTEyQhq/+Y/xQ9ggcAa5sxLY+ySnhsTW+rA
O6g2+un7tOBmNK8EyOwCYWHaStO3EGBYfc8yRqfa7MsiSt6wXhoJJbhLF+nlV+Vftwi2Z5ALF+sR
CJPM6qvh3dmyQCD2EapTl0ib6Q0Hq6UBHeN/hQCkCyAWX7PJxoWc69bXUxQxLnJ8TRlznoBNoQcP
JHw1TT/eVrcjkd2sg0dRNS5Fldg9G9I78D5lQDm3vvnmMHQlfy8F+Ja4d/E3uyMn9Nxaoa8+nN9h
D8tVoI9PYRM1y2cdgOdjCb10Pr6s/IPS+ZaoWaE+3oc9DXlUBCvKZFbWDzt7V1vHO4Bd1SmxatU9
BQTer6eALCR5zDLHYXu0sR8pQ83e8lFUBPdihzekPkNjh24PBxkOTJSxWxJsRl9lsWfINUAsMXSW
AbON7tdLv2HKXTmjX5kGYC1v7Ce62eFWop83g+NYqzgwD147FboZQf3HMLMiJcrcgAhoyMEDaxAU
l63E9B2HHQvBDGrkL5jiVHc1Jud60T5eLfZAQwR8AxNgFJhha4LGV+uj59R6NBLzJsqOON4tpQKv
FhQ7nJY6VOVuvNxll+7edCRCJTLHQh7ThxpRet4Z7vgzy+fqbVQ2SiGCi8MfRHwPquME9zmH784k
szr4PBigM0tiyI8TS0EZIDJZxPGIPaKfI1Y9DGiqY6BRKTY06vBdW7od7YwI7R/MKtOmFz8XRvtR
n/pPd7WxX2Ixqa9TCMwFZHFEqS7nRa1oTwpek+FV6YkM+oBubSKqPpg9pBSCVo8EDSt5S4+SeKy7
/VsBvJZqONKHh1FZvHVQvoldfia+7MEQ4YWN5jJnFLRi1XBB7jwelCo20AiHjVtWbnUEaJ2frWr/
ByuFSwxGuufOExQI1nZpE+D+wxmgrWDtzWRW+wb19axOOdNUIt58m6LxGxNW7F5B17CtEkz6Ovxz
vAlIEgIHflep3w5Arv8OPycjeY9+EpNKhKFXm9uqwr7WX0jYo++fXsA8iGYbmC3s7D0lKx65+0Rk
QI1VOjnbBhwnBFohtQ44vlAWQyAJq2uVXFZFpNFWvk42UJR0imH6pcf0q3dTwBKGenCXUUUkTYmS
sPwZBM7P06CygjBpzb40QDqimYu6yF/EOzdU/Vutf5xpMKMXcfIJ96x1NJZ5p+Q0vsNxe7R80Xib
Eb90WusUOU2CwYUrRXd7vBtCulxmO/0qa11qt4MMnKEqCnnN9og/WpkJ6sTS/JGN4Z72zpF44cZt
DR0GVazr+nkKRKCJl45/EF+EjMjiA0R2Ox/S5AK6b3AEJSiPKNeT0b9mnYHktlTuM9l3BP9zKfhp
CQ04Ubkw38BOB81BwdXpTUR2h0VpRPYnF5Qud4prEUei1rG9dy38he80c6cy2t57Pqf3NQ3ZDyL1
2J2dbnSOzH1aYr7XRaqtMsGjReSn8nQEU6IknFWCTxOXURD93Sn3bv9aU/RnLxrdnSdN2NqX9iGF
am9FkCNV8SPxdDpnDQld9tUwRbyNbTEkHoz0PhxQ2TOmSR5K38U7V3b9kJgXgcZpWbYSXweQhzLZ
vKT1q7GBOHsKmhJNAvS6Uc2gkUNrsErmGxR/kdTrjbFH14TAvWDUvufq0vMhUwkZzLG47iXiqmx2
oySKgPLkoQ2JBrHQ2hTH072FmKnaZFw2ByAsOUQqjlZYpIxgzJRheKMmoFK2fyvQUwWyitTRvZDJ
y8su0q5WUBo/uJeTRwMqfu/1uhwKf+nTZVdtgfk3wo6N6Wn5fAVyqb44s4cXirGOxAh/aBsq1Vlz
N0La6dRX1zNJhJU32oVucDEL3bERXG4oCEEfgyMCgVcDwztpTisfqfkCuFF/RF8ymD4Dm9rQQCOl
+dzCKJ7+dUzQ9welpwo+9C3Qil2GPGbeqKsEfaUMn8+mbV00x9cvVHGVXsoheluCK1WOqGxy5ZK8
hoFTsxaSDRl8HWkM2LRDxMMo5dSoaoakIElE1kh7++czfEGeDttAOr3qKXTu2Ucatd6yIb101lWl
brdYJ9XBUFnyAQD6sbcAI7F9+5B9KJ2zW8jEDV37XGjJZkHnNH61BsPQaSjiMC3otHIn+6/Db0oL
TJwTzkAV3sxCLWEpGF3zBT67nvi/q43wJWAixKTxMxCUwVEAgLa54HYIkumBiLNO1C7ZWJucI8G3
6aOUDitPYFhJTLmwfPFH7KDgCTrMX2q67/3O4FbcrsyP8bpq2GBZJtNuh47HkkdpPKOLXHRyR0N/
mteNP/F8ls9hdKmfmsOUvKrUAGdkMR2vcTzt5TlGeFi8o2vYIxxZ05HVFaJ6NwJ+FT5N8AJBk3qv
npQJ+z4crlv6D9pm8DxU8jrj3t2LCVoR8ebnz1ncPtyXgYqliE2B7Ib15jdHf2briMZJ8GoqSQsn
DePRuAZLZe7z/fFnaBcymuJOysIBDhqVga6/aNpE/v1qTrFhfwY1qAx2e54dexJQBRrOMt2vkZx4
qE2I45EoKZxv6JX/JpWnc+2S94cTlGT+0d9bzpS93Rmbf1LgjMr0UNjxjnQw4s3F03vT/2xerCc/
qk+CosmLSs+0wEEA86JmKBdgRH3Q5tWpESxvGYRdXLxD2Le/1NPBLvm+ZbGWQG+jSQiwrOwtWFig
KJAhmF4zZua3zZReeJT5c5CrAGL6lb8bPVyiYSLeh5AcoitOhX9FhKaFcbU3+ysIoJuuaoESXUD1
PvNRMpC7ZC8Wiw3SCgUj0GAcvWZNBUd9IumiBIMad7gOsLH/OvrL0vOafOgecF4LL3Tiu5K9L/ba
cEq8d2UVy10SqAd7iqwcxjuvlFdkKwrSiXa2YQgSVMFQfR//vgegzVebmFCbLL0PvivWwe2omYNj
SU26kyWmYe8sD7J1XITzcc7SwTWCUKKlquSBDFdQPpvWeTxUW9iWuSQHqzaeKD4uWk7xQHg3cr0S
Vtox7vN2NmIsn7ziG3EGccqhBfuZlL1BUoQqHHA/810uShGU2Ntnk949oYQ6wjSw5vP3giYXg3oW
+3NPWeKX9+omRw+Ry1wdWqFggefnIVeP6nxyZkolE2zlQTnb3ugjo9ldSZ3oWTnUo94tE8l1iU4f
oMUCTEFmTpFU0oYBJif7MerLMYwY694ed3e+6yweIeRpkd6wRx9QoT/gi8OgBsqGNVcikbtbxPVi
oi6GBV0uBqZGLaWaCLGQJ9+pmcSYi/M8la0Ogx2KAg2A5cht9MFgQnRhsTiPN28u+oH7A8Piah2m
5mWjgyhvni9RqcibZLVB8CbvxeRakGKFjrssElfmLl5m2WcTy5yjIP8v7KGcXFo4vThCWFI5hZBX
Fyobqz4D092ZRXbZ/mUClWlmp7mYhmfCFYQZERalUXzszx+7e4zvp8WwvTIN/6Q31cgew6Bq5C3F
EA2ofHKI/OLQhzOup4Fk/DWlzvNrohcnMcTocvZzQ69oVuzLOMd0amQW3HiV/e45zofj85LzBOnr
Icfd/HbfTax5GDUniyvxKJNxGKOo+SGZ0bNUuA3JdxrEq7m1GIRWTWH/hnlLb0qlsuBNpaNljvfZ
Xuxsp2BUEnmbvZAaGCZqsrnmHBdcfWFR22Pbtnc3yQbBZgUkTou8x44iaRx3S4BWGMEd+DW7DH3b
2x8MXaY8lS8eW4sfwGBb6D8J2yo5j3cPFJD2wzAofMu+Hql7sLRoQiuDK2yI8PcEB6/f9/yBc5Ao
HkB8vSUMfofASl9g4p77+x6Pebyy8d/DIdw/jRs/3MKJgYoCGTYZ5l3epAtTp/xhExLFku39QMkw
fIH1gGzTi9C48azjcZnoejC3BdWoBmvWsbllUp8mpa3JI81utxGmolhoFn7TMGgjufydwVhhpw3R
QGztlws=
`pragma protect end_protected
