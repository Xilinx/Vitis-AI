`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
AQ6j7dsgmtiWPp5nzvx+howzaeOChx4BUYKmrupV/fxIRihKV7lhSsxzgfpa5Zme5MJAuPg5du+Z
YzQ7mxX/DcQMuCqu1emgXe5dyEPyZOKcTJditVkqzJ618iFlwuYo7dx3XTnYS3KWa26xP+ccwZQO
S0e55T1IMLlBSEhphrFKTpdQiheViyxH/Zpj+jNWhtxIPt9A/A/+TP4qE3UxPqHNdDjQ5tXLGrU/
HUKk56M6ozfVuuTN80XejcM02DZNlvQcyjYSBBMA5tC54O2G+ji+fbMgkXERUz/JbMVZl1kX/if3
pEPzo6JEJ3ncZWuiRi7O0SeIg4rC6y0uydj4Eg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="w21JS8XT8ZZQagEjgWtJBmHo8J1Nqb0FXAC2WNLNFR0="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
ubHda8TJ0plrSaVcJbVhfhWAx5tOj00BjHFdRVcNQl9NH0RfdshdMJUpZ6dIFbWOKBbOb2GGxppu
cjtwe02MsXc2wPF6ex2W5pcB67U2TsWNyBpct4VqKM2AZDRQK4KunRW9eRaCFjV6EG1KVek2xS0c
hxyRgls2V7I2R5kqF6L0ulcUr9vn28Es5FY4Wn+wH06vljHIFV9HgJTxJCmGu3YuScAVuHzfysGv
odxUrQWOrgjIdexTmurqx95KgWPVwboo9xWDlnviSmXyX1YI2UHQyV9RsW3W8CA/DD52neiQHAav
vyLabFATLPHlHqXRotEjIDtjttpLeMUisN2eergjfNXxpNXZokMNHSPzjzGpaV546PkO57MG3yY9
SHub5cfwbaqK0IZiqCKtRhR4vkR7S1OpxiMHJdI6/L2rVUj1GxGg9TrBDPDQ7iv/eUwFWfXdS5pV
PeK6O79NXV9IR9dqkKXDJYjnd1ztiah2iU7nF3v795EBgLEIyA5OEYFy1lRH9QMemab0yIgkk3RU
+Z5ovHADZNbCGXYLx0QY6FYpA63X2XGdH8rAOEcAc2QJ/Ey08+pWeC9EMGHZYGqRPAvQHL5Dxqy0
9KpDGpLon9dFI8pHllC31H1Js5gWAyzf7KK83fiPFUfikLoeTxV+HRfUT0EGFpNf8FqAwWhX7ljU
PNX1pDrxf+DJK5NvCzHzxM5d0pB/xF5sfBZIyWERmrKkGLoR/UHUe/tpfNqHJqckAsvD5sH8D7F0
wv4FQHSRTAKMveYIaqc1xd/FeGkUuXDjxjNVCh5NjHoK+G1fAL0lrmxsPK3vvoivrgBAeRqOx6Bd
02c6YQYiCKD8JE7vrYE24yGKX7BvLuWnZwspi7G1ZBlYDX0qE3wcncirxs9LkOM94rgYNY/6Vd3M
zIoem3ST3H+ybFI0GnLbVIp4DI3xR9UBDT1835YnvI/P6la7mmkKrNdMWulAS7aVRENzzHCIZXTd
kM1qPDnm3eryNoOAmsd5jnC1ZPIZao18YBcwkT2qXoiisc4SdNZ2VCeSjV5/skjr8Nx0I17qU9QY
2C2zMW/KrHEKecX5AD+PhZzPvOE76SuhDkseifowsgNa4v8UcllcPTA4C9m07ekIH9j2RAC8ifGD
YKbjm5ZqSW2vI1sBWD4L3qxgPaLgI324zycRv6Uj9DYCdg93jIuLY3amaNFyfromXvsfDopSYy+Q
ybnkfHrIp2IEOXLwide7GT2ERUJ0B/fY23rd7jfSsTHhIiZ8XxfnDmoZsXAePa3rGvJbMg6Snkm7
bOxvXj+Jyi2iqLAnrDmTpUG6w9QlPw5RomoeA9MrFOZnFVkngMDSg/25qRFHmOlztiybEdvzq2B+
ProeNLOdzhPzeKCNAVSsIAPDsrLdV5U4ZYTxXkcZxBHcK+dXA9JiY1z/1RMrcRRiPqTyxZ+8Rdpn
GhpkvNOsXVkZa97vUJ98EbrH6gJ4ASS2wK6FEemNz03cCa1R1A6ioUIos44zaii3xzsSsf1NglFd
8tPOAumKUYh7ylqMdlccANYKoYZMM/iAYwOo9LJApRHmnsluscF/ZFIa5pXrsMnw9GnTAudyKTED
IZOZLj+iAYAlqBSZncgDM+imtpQgr2ccj2kzZ6TGHIrJ5WboIIGQ3SgmFY7FsDTQoLG2nBbhuh54
UhF4jTkg9qNAoVurxP6eQVZjaWtjUocW9K8tAXCBMgY8i+l7PKBpaGkUANB/drigYd2QOVA1Mc08
jjg8iDyKLGJo9VXmB2fYmOD22ivk47B1eBeUIPALpSgw7COrZdR5eKhAMZJiNX2AWzUh4JlzbrbQ
zAI2gMNof1225zKVmpJzBjgUYw2RVmPSb6mJbTn6pexkAer23O8J3hGpoVBQpf3PF58Nkh0lsayT
3AOeNv22jeRqbipBZ/SnaEaAqrLM87z057bluHVhYS6ljVoBZQ4fKJ2y/FdwqOOADDOBt9Mda58/
KrQCVxlwEZz9d/pwN3cXKmnK4L2L0zDLTx0k8oMncLpa4Rx0YLODmLYb9nGsMqXfGkdFzT+S2yzN
VP1lY/zMl8kJ5qImAPT8R0HjHEzXSf7dgs9CWlfQO4Yf/DhRKu5Wco6wmSoTy8vYuo6s3tMBpIQr
B1596//KOemcwVdM8NRNymsd655x9C0iYQaCFIu5eQpb6aoEBW1Th2GWKvEUgH/l0HA0aZsjT31V
d0BnRq97OJLYh+M5nLeimlSEp9rv3d/Eeiv+k+V/5MCX1WRj02P9GIBTPLkvD+RJzKUWYeApxG3Y
M/9XsNquI5oLzrcRQsml5AothtC+UjealH21dMS1zql0IV7m6CFXcrZC8YkgV14iA3ZbzPcll0X3
vYiRKCu5zb8CkNIboytGNkmaocP0QtHagUR2rQxMtuomEvWI8iYn7WComIyL0CBmDVfxuo7H/w6g
zdPjkJnSa1arcpXGuoNn2GQwyhb9tX+b/dMpxiQcfUOOyihvsg2tr51m1+iDgDPCyaO41svRBsTA
H5tOkapIHjfOr7xlhQTy0xnR9kzyi2HZwDKRm/c2oUKoNXn96w1ZxCmkozDi+qodxVLQ0yUGe4OC
cZDcLtLgKeEV5fwxj3KIHMWS1LfmMYEJHcR2B/8hnQCqUhUyxaI6gSRAXmByMWznNOr83B9tPmYs
GjieoyyZmSozOic3cy8xweQg2gDeiLiAlEE/j/rMoq2V2bRUx18WCnPFGPdoWsEt7bPWHnDrawYd
3XYgjNKQwC7UXD3yUbzEhwzX3Lm8/eGgDZb27uho1hz4Dw5YzTohu6v1VGNDctT9BYra/jeFp4A5
XouvJ0Bhg1Xh3PN8glFMfmv1OSl7SPfkT1Vt9Jch6wHhUfVdLLRVmzmQ4fIjIr3Ns1ezvA19QrDY
bTntZEdKbbAUz4Kcz1yl1ueawEh+yTt4IlNf6G0iiu9oCN+l529S7wBaE65VHddGf/jQpyTtM1qC
2GxY+PJptpuyg6EtNZhtS899rBuvq13ZRNHRz4uykdavVEVx9CuRjoUjuLoFNGHHH4ktJVUviyVI
cda43pvgZ3YcTgWhzyZreFZ+Dx8K8rT+p8mVP6sg0rQftvnj+Tvu7waWJW5ekXZbasvGcF7V1LNs
zO1Q6Z6J+W28kCLHbk+5OFb6rBOvDSVi4YHbdf3Rz3hlBJqpiWXvdY0CL5gJdwcaE8theZywiDiu
sFSwRTdQEqAe3Q07z4Wk2+oiRzVgjzQl3guwsFMka0BF+kFjBIOkpGlV46LCCdZs3ykFNT7X+X16
FprqtB+/2ym86rjTgJgVCCkQ7CjyvaHxL3pQ9gUIQKjWYIXxx2VjsshzeE9DB3KhAUW4rnSVw+F3
kU7zXOOFwjn6dwAjFWEdOXNpUFuWeG+A8nV0NtiBF7qOdrBxvVuvlfIUYL23fSKZSKPNXMRW2fdX
iMTuUUYVkF6HjdgzHn67hchPaSMcYESYnn/4OCalCVI8h/1ZuiXZiS8Kff5PONTJjxjzw9V5Z1RP
hsi2srdUJZz/Ywer8EY32+DFoUb/ElRLjO5PWKL9z+k7Fyg8G452BqFbZqByOQg6WqYw5jdw6VuP
bzDhsUry1hDtZARIsOdEF+T0vn1x2BpcYwLSpXfVkExT41J3X48xs31wJOP3qz6Ey4VoS9NUBS2X
aAAgbSje/PrJD0xVBdET5Yvhk1uiepkXbKQ+gmL4pA926KedXmui7MaukTUUDzrNfDMUB5tSHWhL
L9JeEfPn1J9uas+nH6H65Isj2VBqvAv1j9FDICM0/O/KYRU8HeCpEFbnHVkQebfp+XuZ9iIE9Atg
UYG3pWxbXx0z5GESDhJazoJO2D8pqgNpbScUuK8UqMH0qec3m9HEl6ZrPvA7FgKfFa5x8z+Jf0m6
POmGL+ACnR8TpThDEW/H8BqfpVBuUyC6wWGCmWDrBnpHAdjL23mty3zfPAJKmgFBXG7dZH2AGF1g
lUS+caSUNlwytutU2JXRjigBkd8+0gZOE29Yz59/X4zGpvcQvGviy+MhMhskBFQyhayH3I+Oq5q4
6j0pOIj00ey99GJRK7DMQLLSGYRNqrL/ckCfhlF0PzYESQkh0rmlauJS0DmmtPkpSlZ9ryaEIELU
FOfD7oyW6+zs671d9dVwPfG4fUiyQsCFTe2Eu1AgmSpaw4QKBA3EVOW3HMXWTWKFC9SEObVfbXoK
rRrWVKMTuQNKGz/KpGmKDhGzieoboTQyuL/1iU8MgtpCp7fMJjkbsqO1WCiQTurGOVmrtdrk/vq7
6Mn8xvI7jaNWouBAkIkBmqzko9x7PE+reeqq2Ly17wuANJEJgCVQmMvLpb0JPV9Q50No182KCruR
ETYbHW2Id9NCNniSns8YWZVhW7PB4iM+H7vsAweRPbwwLirph93pS/F6FUtnGdqu7z43ONLqJ0cg
MTBw6T9UyKXxZjP+tJwF2sM71kGB1XNMpX2TPAENpA7K9T/BwDqcZd/dyY4cHTOYV4YopdXE3+2Z
iq0L8eG1vBcydbG2qQGyAR0/Bg7Vhf6NsHNucOBXkZABC/o7Aw5n0uV+d9p2SXO5SczzuXLADkGr
EqCA9X+8Xj/XaOHyRXfrEb2Auay/qxhPpaOvTENzKXNrWrnJVCzXISGO/H3BTWoYC/NQDvOmbx5N
+fROUgpfaitBMPvCL8ALeepPnA/NhInzk1xhObWtxXwShRapgjGk7KBz8SIEUiFl1EM3IBg7Gboz
61qgY0IQvSnN2Xapu5DUwN6+NYgFl1kfWqUY4enJun6KVyD2OU96raryFNTvRJt4j99NLPZA4q9a
7u99Qdlk6000sO7ON4NLT0YEzn0ejKqJHkNiRsvlskqUNwlI7JtpJJQo/Bfii6gWrDnCxsnGbKVl
Vj/OXkTQ/6PhNG0qMQqGmau4xiW1jGjxDoyUMue4i+WurZCWIrVFj+DfcImu/l4m5u+EtxxXz8Bw
GsNqCzBneFkocziMFaehttolmkj1V2+xRz8xpeFEd3lI8pirmELJUlSPpg/hN4Zvq9iMlrCaVJMO
O3Gsj/E8wH/pIeMq1yNUREHiMpnwb15Ml/kvoyTYUz6eWnrkptV90EXgY3fFHD4OvxzICt8Dd7Xv
+cb9l2ePo8MLQwvLmalRXVSydYBCtBpucTqttSYztMFGonR5w+8SY0hvkarkqTHHo5dFIUhBAOMw
C6kS4wRlVtf7T1M92dlZbpZJULzaNo3reXy4CPoCh8X++HxGSwDC3YIqfgvcYOUgnQaKjdLUBya7
QNnG4BEtdvgMj9a8gcciN+oVUUCZ0YGS8Bf+8S0NNC3O7ly+UFUt0xehDxiQwL8WxZE/0czHqtir
onGlMc+TIx/FmLkewYKmpvjjEvc7In7bWo5PAm24fcjheXmGrC9CKfFcABinJyLTiu2NFKyXfK6m
6CxiURmQEbAx6/qyVUX5gd6tlSvI0YghuGo6GLYg048OIwJdA1Eezo91YO8wcHkIH8EDkeV0Z0II
rXPBJn8ShWR+RLg9qs8V1UU4gRX471pD2GP6FNKUD52sFr52taadbqiWYFs6vYR7i4ZBsweV31IL
pPWUENDCJhsepW1UtCj8cN4jVvZxU6wBlwCJ/HZskkRDauXqEeUhlNoDTOX2cuVfnwKS3rHA0s4j
iunq76XeVo5LRdT+3XFhXQTCPKM5wRM6Vuu/41nE5DF54IETw6VPqMSEkr9ziiggXQV2f97ePlOe
M5WrVG+WaDi98pvLq5qgda/UyBTY5xhtYsgzaPIoij4VGk+YTlhwx8rKZpoxTe7aQyrm+0BEkZBW
URiGDpNTLmolimgPv7mzjPKD6N8K6rq4IpTIHL0tM7k09mSvf5MEhLfg+Z1UVFuVIJJBq0Gwn+Dp
p+4dV7JqobmVUZfPxYlqwI7jrQfonUF2POF50joJAlumsE+YD/Qv+6aQX5JsetmOmrByQgwzQqF1
zDPezzZbYjuJMmAL3AIHNqjSVwa/dy7Itv/qqTr+E+W7pE3TwiKY16IufCe4oOiCkDut7iP0W4jC
tc4zGf98GRQZhLyxQV/pkVvQJzaEw+c0o1z1l4PeFffNDrXCnLFRHySUidjo/4ZXgchJi2asLuXl
lx3FOMGcXF7S/D9h7i5KX2w+MJHE78SviNtEqLKy7Pf2qOzcm2bMWEAxcJ9k468uJJGLtuzLL1E6
bqVnOk3Bxppm/FBT5dH/fG6QXniz3e7eJfoUX8LecvVXLMjdwq/pDP110LmvYM1DccV6hNrMrJrr
mG5C6KCGjYLyqFVu/hbGzR0UbbGlVgcnkJFuCcvQp2qWJFSgcNpN6wYYpf8GlBSBY0NO/2HbGCY6
aTjDUjQFBIUuZH0eUUuA/28OqNz4A9OeLilFXAiryAPal0iu6BuwmOAyGaHSW374Hctd2Fgj65HP
lyBAVB3cp2Gjc/2mCtmMafAWMLBkzXq/GofxaRFjmFBv4KwTauTo2wiTgTh7J2HKawZBtEG3YAkm
UdjuWTV5jlVaZtBqDP87RMdtT8Zvp7DHRj9Gm1z4gaKkpJ4nOF1n3mqTW072PBifCcpBcmMfNo/8
dpZ3Y1/+8mbPTVoSd5vQ9YuosOSoqO7blmrcfrdof8CU30dqcqpMVpq2mj3W99hLY3/sLKorfsmP
j2dxNrJGdO+Z9e1pjbd9b3DF0D+iLBI+bYgN7rDsKKNeXKU9tdLp2T76dGBTPwO7TonKkQGh5kLF
Xvjsg1xiqnnQcDK9m2Tfu4YeIs8FRzjtWCWbgapGdrGCAm05OWHZkqMq0YpabU8V/COGXuENYwwK
9TQb7Qd9YYlcN/eXurYVBJNMexcO1kKylgy/I3jsl9C0ei/darIyy+osDTD2kqGMaOrckSk4f+uE
hv3q6i4dSX1uXW7KkgvwJCOHxZWooYsUIOz3Om0cfRRjyOhHoch8n8O9KLyFwNdfRTm/IDmRZjPn
QWJAWcTPRfSqFTPc8rgFAzLmG/9l/xgELdXYbk7e/gqrY0UKae8whELh3UqvGFuQTgeqFEByZQyS
wQ7lqAnYwKTglYorOHaWTBUZfIP+HEVSGbRBWtYjzc19O7brV2vz79qBrIphAiJKFGGwxl/eEn0m
u6FzaMzA1Kf5+uJXrLcHrfjJAHRAS149hRs/fgNqeoGjwPG25+Ik3kC6TKzGx/lWypZMH3J9y2Pk
deChQs27HAqUe2UbmLHpdPEPUUEpQ1QH8sPMKYgAi+SsFposPKyMTbngpaM3z01wOnZAoKtMp1Wg
FnyvtGCbz/9GPYzQGXIYJnHHrzsEF+j1ietB7v/87+O+/wcE0GPNifQ7AxKPBraH6jgFdfcjCiAN
M+ScwZSCGedOuGZVLq0wvfJvrOWnSL78T/T9u6ZecJ1UW8MqZwMtc+5f/axsnTWXffimtmxeFNs1
cEwNFCSJ08Gnszg96YC79daoprFAy9jkOFVvZy01p3Cwt9UoVr9uz+dzQG0C8eBX7qFVtpjdPQm6
BkXKX8KRIRvjoF7c+Tm17cGdPMx5GLFY4v7/TzLVPRMyeMDFSVzkmcTmi+nOcg5FZnf3RcnTZLWb
GiJQnS2mmLOAnmqmAaPblLTh708rg52VEz32olzT1FTes84J1BtEdSwBu8/FFZDJ+q3QisH+u6/O
iuirp8IuCUchcluFG1a9f7Q7zHhbq/mn938r+qdhbai+DGeGd+R7dOG2KfVYmLq8rUaI8GKQp5Tc
qtKFmk1ZXXaKZgxCG6kMn2MwsFujzqEdMSZp/sC9xjaRZw6cJ3aYcjhPG4pMq9hozch1aFqZf/mv
YmicqSop1IvkhOoxChpk7T8C8nM77TUrsjsi9hb1Lt+HWpbhCyFT9F++XWMFTGQCDJEROfPmKzMd
xygFflzJdoRlFMnbnG2kjUa9aWgDAqDlGON3ZceG+B8OZA8onb7VW1LKKIsTgFIwq+deviPUNhs6
oybJSfH9MKDNbAiQVl07OiEk/2OyeK/gKcvUFaT+qqYs5gxBCH0klqK8VrYJFpUkuIxnPA8cT59g
CDGhNmDqFNqwa66aKPSJ8btsY2K9nITzeqeVNfGjH44iBNfKsnIoc/ptOwOWDS3EteuqpKCs1UV+
QL+QmbtaCBkUIeM/sJ5Q3Gg0QkM7g41vpZDG4glWUzgVPvjGBkYnQZuAY+7PWUrCC4/TawHBGwQS
GvTZXUjF376XQ9COOCYicNbRgat03FMU2jEFxPG+wcUrDecZXJ9W0p6MP19rpWARjFee02kgYw+w
6UdPIbobWNbAuP3lEJKTpdUuQbqcoUanrG2JOyxx6VWHh7mJ1gMzUBelPTVlVRb4uWkdW6/Be52j
caGbiQq1TMmwF2e0D7II/OecV/fgWYHWAv1L2ZBfPxp4f2wOya0LxRykCX1wrAwddcc5gILi51tO
3syIgZSaTiFTq49ZQEVlXC1ISyYMhYsWcJtrSmon6FAgm81tpn73dHb8nOsvNwxh6Beu25BqJHs3
KA2w9wzMbS22XjpwO8WL8/zmoyKagbwKqUOxb7VvLZ6qtyPMhO19SSugPCjCeT4kRvw0+Ggl9J84
HUwiU3cIgdvwolaoeIVdQGVyeClL3MX+7ten3qk60X8575zGVT/30DtFedaXp9GOi2i+M+RAIjQM
GN3KD56qfoyd9TiePxFra2QWfM0mWTvuhA3rOwkQfzE7V4l4rIIStPCyZF9+r/7pal60HPjcKEqF
ruI/aYB+OhhknxOtaoWEu2hpopcoSNCG6PBNvkhPmD3ldI6dqCfSUug/yG5dtjpVuUdTTYIHilZb
ECsOEr1JT0nzydaDi8ivVrm/MKsJQzU5/Op6WpRKlO1WroSwiSjKL2Q9cdVzadn4kguvYCI0k2CN
BSsheDYytztGcoSVH3n1m/N0+UuU8VtY/XRtcAdA1RF0fa+JeqTAY9803+jOXs5GaEer1GpiMg5d
JULLbndWv1gJJc8kzSOHtZ/jw59axBZBVWxQI8bJhac0bawlgjjzh82wCzQLmvaF3FoN//xeWw+h
nLYabGMQY/z4yNqn48dqmS3gp0d/x9IeLF0JpF/eEgTU/4jpDv9we3urcAgrXOnPvdOiMzFdZq4B
iXrp5yxtlOKMvdouxH0R5cv3Xk1MnairhJnHYLibc5ZMXfm7rkwg2FgyakLXG4GlRkjSsnSuz6Dr
81m51tpLuC0ducHY8OMwt4oELITxyLDsz7rbzEKNsvht2nV7JuPUQqH47r3HJ+LKheKmpYLAq39U
eljJCUTCiEq/M4K83YDV9UIKoUIkHC0bVYnH9dmlTqAqbK/foXk4CLT/77o4EdpHsd9uTSOh3BDF
BJIIp94xw+YvmZLNn+e+iXMvGGKwgarYbTyPriig5zZd3iRNKNimWaFuoCDltq2QIT5mJTldcn8T
zQkSZhC2edTNrHolGWTkXVGS8j7IOWYTjNOC0wxTtM3bUC2GPAK4LOOLgt4dx9JGWdFsROqiqgbu
4fuVLYafjRFkL3JvBzaebR6cHGDcfHrYRx87EAU+bn1OTs+zPLOTWDh+KwyCSrarx6E8q4zPV55R
+p5rWvgx1tIHNxccbjOFzwL+npndHtZY9ugiBkRCQsSkedhw3Ngd06nWxIf7A8Jsn5FxTIJikzdc
bzE82PECGiM8dXZDUp/Dl/H3X6f967jB72vZZmBP+jLexcUz/UKz1A+07eq71/m633SHlT+V/eCA
2KJO2lpnmG5FjcT7mHUv2HaEDXyHGy3f0AnXYNDyyXsEiVYLVcR3ABq8KG3rgxjC80sES6nI/gxG
pKuyPMw7NC9OuhIonE70d5XAR6/LyXxaM1/AO1ELVkJT8TOCI7IQKMVuM296oYC/OZevQpab8xkH
UHr/foXkvPb52uucL5vP6/QyNNn1HsZer0Um+2dAjX2p+Fml3e143umZrPMw+xDHgQKX0QMeg4wU
VHVbCllqsZ2vQmGp852qkSYkONK3eBu77nDKuzxt52oeF944TsidhxvNe+0r7hfCTpylPapmAE3s
zaEX8jNhUlxLr67f8HSkNGJFzAZs+mWpgHEIkzQisQBBoCWCTLndpeaFGd7EDkG7cmIudSzm/AAU
SVJUATW1MEOaMKxUZBLXHkduiRXJbSXE3YGT2bL0ZYKZB4ChtZoWvjvm1+rE16TqYKpZZrtLbxZk
M+MiuLc0fZdVxGabN6es4LG9ONQyI4vGccxP34/0xAmlGNfYycNL6E5lRJrq5NLRYXsb22FIfWHe
KtgpAFXm3DMlk7aVO77sYn8Ctg95g1rFYKry1/k+tYvyrx/ch23TSgJ32bwFeFJx3PczxGVAn9Sz
es7EZUFBgNMooqJdocOuzYSw/O5TXFUZDnamxz+1VmXJndUKQ4li667PdA4wD/nEAowq4D5E/sp2
wK+dx84KzkYJ+u2DF2Oe816JXnjmcyEanNF7u6Hmxc+w7pVgdkUEK62bUhkOVMugpvsAxzxPLcR3
hg9jZ7fEpmv5LnShsK4XXmT6xrTaCYvIrLzhBWotPhVNjhzBenw1k9rbVFzhKPhFBRNCkiZqnEh7
F4aYq70+5cnkJwIiZXMW8UUJxFIMfl+DvB4wFgxqWSHfAdLBh5uORung81e+Fu8T9Qf4yPOXYXfh
1inbhDMawxrcSp26y5+LzW5zGdKu20KJZ7FE2m5de9G38ry/JYiGK6EeWbQyFYaCwKT2Ha+6Qqgs
RdSERrcQHE1RqeZMuVApUnoik2bkKpKxV6pV0FuEjUtDKFUHcDsgC95s0fsg1i4uFHwvETvef29Y
Ul0vgKr+mAcMPnhDrx4wvUj0D6I0LXxz4UgEX4kNfpbsBEtkt/AdLLJlP93mp2HiwETYN/Sh2kuJ
w0ZfxlUzWiMHmM/v7V4UStj8KC9v8z8ni8pd1IY6KUSflzzSzrR+Fg0WGFUgq+dPWQjXiGbnbFkL
lRelGXFrfBRJzd56vuFz6DDa1Gu8PwaDGClrNwzmzfRy7ohgjXJy1PQIs3zMaLYdMVZTuplu0ch1
/6uoTBGLXF5UbLDno3ft3wMQP38BzJRXeUxog6a0dtqRf4rCxGCBUb0Pkpa9dmpkDI53TebhDgDQ
ZiICdIBUp32Qht9DvDyTqooEHlImHqyrHJPbO2cbuW6A6oB4q20gWe52bTfKd1d6lWkz+8tBGp+J
GHDQ2QISUNkkZeDCMkyBwv1otik73GC/NRPA8poo74Hx/xjLWwGPnjhtDzC4wPoqiK0vvkYcSzBM
4IIZxk6VD+tBB1+f+Oq8W7qKtOililGs/WHNEKShiyUxE6VB2HG8ZZ2ZJGa7sM34GASkbfTOh1zX
R/DqpjOGzTsd1/Q00UBXYDWQwtRpibQRMzniSAYwsrqeV3ja3sdjGdXyykxsI7t6eA3cZiJLkGTc
ruM+ft+kI7pHlFLeD3jYnvxTYPc/7WrMZbuN40A2r9XFwz51IhMV2zTqVwsjb2MmsFd5JIlxaE2q
GVXID5vR8NIFvgkWH/Lq8z1lsdy1wpTV0HhpGn5u0FUTK2tpLCFi8sDPGP/fvaJejwXfZZJThNsS
oYKV1+qyohtLypPOR5HA5H8vFv16RuWm/ZVjpSpNm7ze88Ha616xiWOKp5Cz11qD9CHhAvSifkJJ
enSsWDkY7avLx+uNieS5pHfy6bb+tyjaHASP8fSGhq8KbAdGCgNnfQiJvLup1q1kQ3FImkQfBzKw
Op2+Trsil4uqeIvAdWb7Q+SLBRmig+8JK0zk6i5eaMExvv6mv6RFfw/68/0uosBbUyLHTDgKuBfD
0BFsDg42rnhswz854uTUC61WkwuE2MoJKDUhoMk4zk6aprw0yNtQh7VALpnTD/GDx5cX/JCUqjNO
TqXGyDQ4BYhVhoeAZbdvbvW2yC5gTGOOjHpBAqqer7mCXGGFsfD3PHwvMfBHg+C49kH8X4vpUqJH
SWleUo5VNUnVCPQaoy/RX+G+B97634ZCBohUw18F/tpbA6lj8/pDg3b5n7TjGydq0t60YHNZSm+J
rKflcS6XlVRqjg9dUagKWfLPbpawPgqSllsJNVRA3A2lTQZwfz289lnq9RfpuCAc1Zi4i5GPmvpR
2Kf26TBcq3FYykqvVDzQfvpxiBx/QmSw7BgJR1BjZBYH1suQpx5rep8Zsz1tCLOl+Toh5lz5vpfr
jjmuX4I3wcZLGiRApz2cPgSjEJ/i9NcxJFjgcCjnTwWJB4stabPgeXdtLaI9RIFUoODFiug53KHo
VhKPn1NUcKGK74MteG8tinENMmTU08D7/7PHWS9B+JFKLpbXUdvvWQ240S1Xx/muKK6las3jfCvA
5fGdfkHreI6Au9xh1y1/Vekda1znd5tOTS+ZUold2MGNSMHSBXMgFU+08NRO6/Bp2aLyN6CMdPr5
uXcuaK5aAs3N/Yr7fwkWw1fBiWHgU9vphKsHJd2XmXe2cmsvO5BpCiJomBm8YFsNXkPY7yugJahK
RLwES82V8PuFUFb8N/nKBXkTtaE2OOVfYlQ6qG5ARkoln7V3+4ESUo0dPc73jcJt9WyTBE1Zh7u8
epcHxEAT6X0q0aBSCForPdlX8c/a5p01p2MIcOkYnlXYb4k5kikK9WlIDp6SobRJexWFFFdGxiY3
kS6VAq4WakjFXFGCtOE0ARCeOfJzoyeyOu438gogZ+O34KWCuwzk1eGAbdLjHrg5y1iMmex5hLbU
hf/KEk+qZtz54W+UIoUVyN3qV21TPWtCIiqn8bETPkms2362L1Gl0UbjF4fjho3DGjRUzYGv7f7X
DrCIkB5oTXvBQ0wxqYKplVkZr8b7l1NLsNvQg6lSEE6Gs/C3vSUx2l2PgcZWco1kA/HFhRmWfC7/
RoOE4WoX/hF11s+loJ1YBxQS7h4/+0BYhfRDBOfrqtX0vp+DdqbUMSzorB5/9k2wIr1Una1J7WSU
7el79X82Lfjcpz6jk1dUtxkG3QGj26r85CnC7shCtwo9DVqn2f6oDFajwX/ehxUAkpnYnW+qVkvr
LgW9yMXH2shQ4X7Qhb0N9i0EaOLj+vx6mgoVqg61187KMzBYtszDLaYB3aQivknqWTe//vfmmHdH
KShVzOxAyZflzAg5a1LdoxMQ4K+ieK0ti6mV8id2q5MxQ01Gmf9ZH6BCvYB1y8UTldLChsBp0gjg
iUnzYtgSAc0CHVKgu3xQy/8t/N93RLIcNJ09HD5mxv4QnirqzZ3IT3+C3GtdovDLveNfjcLbjwvf
C2YJrXIEvnG/Sp8rrcqxmIsaCB8FlQAOFp+vX+/RIR603zrwvruGJBp6GKzFRlX5TSukacHGRTgR
98M/HY/CF82ucJouErbeU7b/8/F3z+LKnORFFGDSjn3bB8Ytlyo6nsnv9qKFFygtTOGBa/PkX2sZ
mfgAQQZie6z6/qtY04S1P+VyHO/vyFR3qe3Ut88wJe2/MhCPvGDTahTdXcXh/7UxJLvItRFQmdBG
jDRlrrXxXaBI6OyBAwAKi3LwtYKGJU2bXHCOC5zFHjcSOxEQPoVWYjXGKc2kXh72rbZa4aZrQxma
fPQ/fcu/GSUSjbzLo7uGPcfH9vbQ2Rla0Z0MwUAExExGYPliWHX108W3Wm3K6bZQX6865g5aJCTo
0u8kXmUPQk1BZJOSymWYfsDaf8PzkBoQjSOWmvlGk6Wzc4czt0tPYpIHb8K2qIPzOlzgyv8aw6tU
BDvY4ly4cX/dIN3O4ae8Jx94TeUlN9iSlPjUFWeb+ws+/CWHxAR5Jpf/8bRa1boexWPuey/tOOHC
zwhLeoSviz5QcnMqmlzgL/5WqCTBvshagwKk+dkCVMYQRrBPZ7UM4yX3jTPy7+Ugj6yyQukjQrtj
MTFTEJdHkomGUX5Xz3byVMHWLKxnMfuDy6Vipocuh0Kkgk3DdnBSL9U5JrYBdAa3w8BLvrm36+xl
kbMd1IVjabwxITIWu+UJjzkDBpsmTZyX4qSX4Nm1g1nt6tBtbS/ul8AkmGy/wXDhLCZ+kaStlko+
0tBDDjXeH8PQEnUFqa9eOAG53NST8XyX3jqjQRd/4zbvW6RQX+dvrezQW6NeVynJdoPEiSf6DG3Z
pXtnGh0BmGwTj0OyR/nTeeGWNi/cM3Y90ojs1EqXQH2RFQzzfknCG9feDaryCPS7u7gMVUnwAD98
HqfLb5ArNwluXPX783R/3TpKMGKSzoh5tPD7GQ3vN0znlnx3S0JPeSC+e4PoXemQeBByOT5Y5u+e
0rc83zo3a6R8IP+Ut/l9kPtxhLIFddAQEza78q3AkMJn/DbSB0toe0AGWyi+TU+DA6PiGfmWAZk/
ajcrXqH9Tulr0UtzqpamngzLJZFiroM7uijZnVBWQ8JJ3iKkM1ayBe8GvPAxxfWrCLQX46ByxBN8
YPlTSaa327MB7EAuM4tZnzD7Jt4YITN/6IG+xqGDkdfTJh7DPfHrR13aJtpVRi9WZ3XRBzBpIQxk
wVIhb4t1Uaw8zZXyFqCjYPKgVMIfmImTGu/mW78JrJcT/DCnrtXDDkuAY5vtAMW20dM++KP5GWCT
H99C5ZW5qug32uVNcycW6X86EkbCvUcTjVsgo7raU65H+2RKZUFiK/1GSPWRfMz9ckLPYoBtMqTo
Qk3S12jftnWrt/8hAU1zl4LxN2ac3hy7jorBu1Iw614FCxNWjoQz4zk4ZGMG1zUqUpW1AepAzqUe
Z4QuxaZCvSFE4HXaSLhShY0Txai+d5VmqQyEHSfStmU3YyJ8M68k/FikQ9mygzfC9TEDvsybaJGC
5cpyZSixTbfxKmqNkGuVhsGuunE+LsY79iIBwwObyaWm4Id3LqgjQS6PnhEk04EEvLIclh7p0sXm
MHUtqyD73anMJPN5Jrnk1lcVUUL/hPzd+yyuQ72ISnoJ4OCd0xhruVsckPoiyUg37eGLooOHZ1t2
BbtjDultD7r+x3daygHrgzpE+yEe1QiH7iYw3hce79G5NWUWj6T/cdG6vapPL+D8XzERsgz4hHnI
dNbl6FEkHWnDB0cWPyaLrKaTVpqeYU6ys72DTiFw+U7P0yEmLiKDBtkd3dXixFB0cFv04ecMJKXU
b9/yvAUSr/stJVTp8PqlgOmxTplew1ld5FkjddLoyHSzXsGhi7m73QrEgxx1Vj/u5WQJsTTM2aGa
qrTAP4DbA2bZPXDQWNTmqRTfy4dO2rWWCgZ83j+FvBUG/PGCNrVMd2Rf+XKnHVNjcB2AG+n+rrNJ
4bcNj9j5K0NX2lrAwqq9j4vQfMlVdiyV4wR1sgX/7pd+Zj0S/VrSHo0GrWQNPyLOM6qSdUvT8Jpm
ig+YchLb7OGmD3DwDpPtkbVhMwr1Y+T4qA7bowvU6bQ8eX3S3ddRLTzVdHCxkxxzxZEO26Xp+I1S
fOpbSRpr0t62qSSOCvKiTHFEmHwZmRB4xmz3MpPCZ8XsoySyI7AUAdyoEceAzOYRb5w5z2hN2INi
YkjOFTHOKwV0wQWxoNw15M5f4SAvbxJH079Alr3TSReYnYKbfm0EL/WVzD8y77D4iEkaBtvW9Apj
gHVKZw/RebxcenU8BkxO4Xs9DbopJezZ6E7VNnnBoNcMiLqQs1QSCUFWU3udYC9hQkrmb4SFcjHc
rN3s0ZVRSfxZSTn/87S956CgTHmzoRTsGjuTUu6NFrK5h/fldIq1XLhmeLiZF2J+wXaehc3uwaYd
32EMUh9LQmAWoJkFyGjQxZnX+rRJyKMCAQUCJGtxZ0xqk91omhri3m4/rBf4SF25mXDcEz3aPTvE
tMDmjhFFFTmpb70tj5HJ6iWDM4/O+PVjx0zSI+ujR1TcAoaPUKjH4PXVfbyqq+eAnoB36KTfVkqg
YEvXGm87uiaaeK+gK3forxeAlLVU743Tu3pDSWuR9DnHCdXnjCXPbLxQAxnzbzo8SvtlZApLNDJq
UMm8g3XUsvCl53rOfR0x7dIxnd+JFC5WwxDED+Dg0fHJD/1Sz2FHz7YyYLfH6gswvcQfj2sLLqXW
nDg51LHqepInDZ33+ylBKdMU3w6Xv2L+//ACkJJBs3EdIaNfONCX+bjeY2s2IRoJD8KQWQaOjDGr
GLJizqtOPJL2lF4f9t59cofD5TDAo10RzE53nKm1ulevvxoEDde2MGX5sL08uNbMMvAzNmFyJRT2
RLhp5+38OnbCF66KZ38MExrj2LSvu0cQTkNVMAn9geekwlUoF5Z1ho3MAiuyl9yViad7d24Q8Jvq
Pve0Ne1+r45aFrJfOdIMcEN7iZS0ZCKqw2Hi/vp6s8Yf9m19lnYiWqgyBBLaeKS9iGDrZO/uiUmf
XXOMyqO+jL59CXUFiPsFVCNFv1aV3ZFXHJ0dXDpqMmX6hJrgfbS/s6YvcQhDvv4Le/tjT5cJJLgG
3JxL2IgC1swdQCda+2xkDWX/pqy6qdBBVOWzRdTprELV+ZlXKxAX+fuBT9xFiXtFhqjEzNtGa+xo
raSh83+RmeIe/6jR9s0Pu2Jjpe+5upfT2o5MWx7TqGvRtS394I9JJlX10EqbE6kZKr+bKyc+QTXi
ruTyVUMU0P4fvBp2plFNC/JOvZdSirKpo9JZMDRHwlhCf8nLBFZXygWQStdamhxw8HNPS30g/Obj
ZpSjJPbzbB0K29Euq24TCGweTr+eIKE1f8LWC6Vm6Fr2il5pL/erwJwTJWjRLkjY0Y4N35D6DJ55
segnF+Q6Na5IcIF+FOsqIpRfu8r8YhH3QsRh+irmCh8rwzznk7Rv5lWqfn8FYNRBZ338tvrgCc+2
h3bmqydpDMPiXPSnPkoZEg/9Upb2MKn4J2MGQwJNXhFbga8oraIWswT8n4zQsIqxo84tBK/Y7tqn
WX3n/OvejqeY2+FUifg6MyanKlrObV907I0+5qf6WS44hmiun5Q5deBljO3THZjKA/mNNvcm/Cuw
3AMsa48D0MCrgfAZOf8uocqUxbD4UweDjIm75IJqjc9PRJ4U+clVMy6rGH6dgoxNa9VyB9hfaq8k
seRX/wuJ4S9irtApbU6bAvIm50EuMnFtpSmwwd+kDnpJzk1V6Zn7hrxng3y3H6KocgKvW+ZuOwcD
e/fdOkNRblJyxbKNaLjmLfOQWl4XkG3/KbKwO6VpWmdiLUfc6a6ztHx5PoIscDPQykMMu+Qw96c+
lfutxSQD/NHDkkgDuPOhEPS3g9un9nvmEwhm4tq3B7+XP19UB1/RMnWjdXkX4vWaSSnQUxnd/t4v
bjWcbxIG3gPsOykkTFMYIuqRuLNpKGU9t71Dk30BPifyhb+2s+vlQ0GWkDOF95aZQWY8l3sVpqrk
huaAVnwGj3TUUo3ViKbFhLRwTJdoUH3TTHZ8u7YShVLcNokhN2Sz13miysBs/cp/esLBKvRV2Um+
x/qphU57YJHoW1luwWIPZv9OIDf26dl91EUn2rbPqUbXpXIHf+TNcxfDf0ytd2WZt+6L6vkg8lR8
2bvsqwhuUVOnVBrqGZox4/UsaQhD0Txft4y/C5KLbPom7VVPlAluXphQm0P39MaBaL0co6Eebi1t
Ly16j9zZqblYOJcTCUYwvepG3/8xA5VcMPYa6YihYKoVrA0CxD+EbNIhXI9GDCftogafmlodnoPQ
skWGXv1pRar+FCaNyYxoX3BGigJejgpiF2FAXxD6yL1FsiW1zC3YGGcSAnWL775/QVbQLPPv/xRy
/cMzV1wonclRaBYd92LX0S05bV/5W//mi8uvsh3r0ywWpDPwbRtu/1etb1HMGA7965rxYbPSOUfS
G5mX42vgvuzjlst2J1YxUf+w780GFA5IoN8jhIWb51Dt/mdG3Xm9L922wJzY4B8x7401o41dFjUv
qMoIlB2qPRYO/+PIiEVvQUa6tJy6wU0WNQPlPWK2blmCdmMQ6NTl5h/n/CJGIH8SZtFR2bDHxZhf
YRCuS5OIuTM5sxenyBa1b/kwE6oIGjFsp8hqT5iby/heSFGyoI6xUUQtI6B3+dwOWiY21imrmHfU
vLpdkaRmbI+TGBaAh84KrochI04O/qM/+QLyqe7HxUIpDEGSJ7F+Wby5Nj8BrII/mOyGmhwR8sP/
cPILUN2hMyuoTQ80D2W19fWuoWY1RxYhapwZy5mhO4k8R/PMGke86FUXjvLfIQanHZik2Y1wWtFs
aQMfmGT6FSrfRqnWFAVxC2AD5eL/X5IoMB9KE5LGgvZ3IClWqtEJHte+i4w6npwwNJ6aAHNXNnJ2
pJVKImgeYLyN6osgrMXyZLriXXWFbYZTIWBOvJaChRwLa1kbFlXaxiOmS4Vclj5XfLKZjSRu58xZ
E37ItHOKc3MsKlfIVz8AKykkf87T7JvoPtv6lor0FcwGhOq/ukEzvJQlPJDk/E8QOlPiTvvtWwDT
WrwnV4SqpzrFZxidI2UwInJfcvVVUCK8bUAIQ1zsbJOSoyYChwz6u8bJFB3wB33JmiYKCNdw26pF
a3UyWCR0Ot/E0tWEDDX9iOd9XPVRaKfYIj2YNBfOFVysg6YgWcKVJFXKrDHokC2PUT+PFvh4Jp7K
My06QVVr2T0jX2lnElBrcWaQv4fseZxmYAy7dIQuQ/K5/8FPXZD8h2By/TkEv7goklvA7tplrqUH
DO1k9wdvnc127JphOcRjElSomVd24otg4e6P/gmk2bvhwXh1aki7pd7qY9otFiU8IOFw56cG9J/9
PMj73WEB+BG3/x1pmg4176666YKjeOwPoB16coMg49YrGEz4etTY5lYdkrZuwPxIjryiehynsTk7
16Q6yJGDU6BebYmVBE7opyeJX27zorRLvBJ6XGVtl4fetLB+xdy7f9xuomaJEKplQufzLhdz8l4+
qEbhMcsd+AkEEOlV0hP+iswOqGuP2zpfiBrXIXwvu8iIlCfB4x55Xg/7JYiFBeT6RyquBlrFFSIu
ORE5IeoFVtfzHjZGMA6pLXid8pT/nhiBBB18p0pwx+VLJOKFX2Sssi+2GXcSZ7mwH6sf+pmd5XET
cR+muQCMHIAo8TmSYm0CRrp7IEcSBMJj9CUv5uqYSrcxESAgthBJmscAuOpMCoHh5sssFYhvfA4m
6n+TLjJyxIeqMaZQ0otWDfAjwD0gUY5J9taJvGpj8yaiq4+Mi8V57XZbYli+mvXTwM6/NT4KnznS
2rUgXk1Sajt2syJ6Tf9fAbVvNc91UMpWA8Aa1+DvP+KV52BOwn2cCFVjMiGurYVmmssDjCLuvNM+
K2T0od5LQs45UmvDDRHlms3XTthLFr9Hh0NFQVzfK9bBYfbyypqCb4ImzFfD37fjC+wSl50nPtRs
NozQD7GovxFfaJ5JOEbr2yOaAderI1LFYT3v4d7+a34UpywejhWxTAuRCjO+Odh203Z5+xcs7vce
VqJOvE8j9Vo4xyfxpslpODbvtOWIbsRguRGHSctbr7eRo/4LisZJpeR8P0TkRJWuq3qH0axlKS2E
coelBG3adkJIdO7aiJWCCKE57hT1ZKT9+yAaFr3HIazngbgq+zHo/GZmsZuef69D6Hq84PHrNM2m
KaoaFAE/J4CsrsZRMruwcv7U2AmvZdNKDlNsbHGIvbWCkS5HX4gKOjBym0KkFHDbGsNrRtwqXp+v
SfmLGK7LOW4nLQcUgTnRHSQBN7HxJwv9C4WbdQOFyAiVrDJbKLOPWhx0Vu2d/t04461XrLCptdKv
19Ne8QpCWGg8W4SSV4MH8H+rDf8QY1CoE73WpFxBCUF2oynZ4At2z0e4lxGf4RRAqeeb94MKO56X
JmT5YaIYbLpHZaZqV/pOZpfeZNMDjGNxzvOEgQN5E997WyVquyrPUajk+//zD3Othn/ZAuFLcEG4
NQIv6de4xRYliPhNkq7r89Y18bm191SezwEkb9hgKRGTu9h7Q+DrMj+KhHGe2lnkJJbf0Ae+4RL0
OQz1pBkClDG8cUuUDETMA1By+QxJJuvk1NbswUf/rAUuYrk1WNI59u8AgvbPXJwmwjnZYTkKIsuy
tXmjCRtpzhwqnto3bHm4nLHR4Ovy1cWOlgyLOG9c6sEVc1oBVv1KR1hlkMDxbxItuEVKF7WvKtGV
mHWYSdvs0uT6si6JwfIMRJcP0ioQxZoFZjyAcSgvlW1MeF4uWnmgG1kEMmmj/BTJ1EfS2MEmtrsV
2vIwD3aBXRI9Br2gbnAoPpZqLHsVi/bKtXE3TzBo8072XJLHIhIbyOMybaGU+DjGiqtbdsDq3/LH
pPWhySR26RXump5VMs5VPXTlMH7SNKsIp6uhadEooWb4EhmSIhGKxqOTffMWwVK7XLr3OlPluw14
oYdSHRlK5gkvhlGrvpedQ+Ct4uJe2ro0J5ZZ22Slo3KBiRDdF0D3eViG7AdHVUzkVcldrEVfkLRC
VF5E0VqOnaBj8Vf7Vk+666Myjpsjf0EKeJGIFxdkJ60BEOyqjSATKUBY6hpqhbZOv4A8UqaCDVd1
+7rUI6j7aBzoR6hH/5GkxHkRHlhp90TQYgOC9nFpmDNSsY4KNJPgIYqMvreSp+n5vtKENNQ8OcNp
9yiimVP0Fh33t/9TOhbwqRi9cr+xOeg4Ku7hnSdG4NDIs3LJfd4/dQ+82mB/ExC7jMy7RhBezgjN
J8PP+TC6XtT8f24F09NoJn23bUumuiTDOfk1ZTnZKbIyWQFJQkp1io5jQ5B4iUQS0JxuLKugQowG
gu/u9HrgdpiD3Qc21qk59zclSl//yT95QhGfXqs3SYbLCX2Pv85CoAceN7Vx0hLRYof+RYc20Sl4
X5fP3DsaEJQTbdRxLQjpWyw8JUtO3KT6geTM9sTCKeDOV07sIRqdWiZeGm5XhNrLaLyVVrDP3Ej1
9nNw/HV9vwWReCx81lzJPLi+xpXMUSaTL0dgHW1yaYgGu1t70XVm1bF+PBF3UTBfEU4kIKxlTUhv
RpHHClP1RathT/C1ysUQh8KDw7nZXQNQlZWnya/63urT5eG9bWrlxoqC9FCanb5FEZZNvDO4QrWJ
x90wzg8gFCj3rMYUEhYlhlNYL6eTSeyCqTYKYirrH/URyS4THp3/TGrlZ15v2BWGbP8vCB3qwTPW
b+PIehchPWFbFPqmb36tHtleUCJGQyaSFe6UwGFFReVIvxwyMqhyj5TYFDAQ9SOlFZ/yA+fduX6L
90hZFzroRCopbdhf6b+n5/IAcMhM+S6cmvdtDi3EB9zxe8qKeDHBS5laVLCsIVCJOKMH6w/TKU8y
4G8G5+/6cUKKKCYBS+tO9RE9fwsyZVzg1SxacZypSPOfXHC2aIPwmK0+d/5ZHKx2WsdNyuByvmdV
FpTlu8lY4G16BT69GxQAcjK6VYmz4VjDrVVuzYpLhJdZr59CSPWwP8/M7GKPFXjlaL86+ViW1sIP
HcSFJHqqJ19cFMMowx3noczj3ciysei8d/E4t0/Sxh2EDfyy3YRg2I2JFHmvymFKpFuLFD98RfVn
aIC2ai4jvDyd7G3gTVthwh9T6wirT2xiV+aen1vKQVdGwpj4zGS2p4lvPKmVcrfJMYALzbPzf4OS
eO0KhDkxr6E61db9dhz1aZzO4eCfY1pjoIEX2r1w5FxEAemEJH+8sseE7GHuO+KYr9T5KdUwqduC
peFLoniPtQrlmGyPuc4LzTOW8la4Du8s6TsxHFxyiks7PmTEdhdPHzOqbUu9DosdJSE5UkSPU7W4
8iMiIyAZa+oaoEF2mNckesO/F2kS6UVyYmrKexiUzm5+Sl+O7REuLDcOsQKhnIsaX59KGuQp8TYS
jeoo+0mvmO0U/qTD48fa4ipZaqE8c2kIqKd5YjzTZh5tG41ap6z4w05MQa8Nit3/lw5KkfDB+FLF
bYlb3tBmMYnwFS6tARkeInMxhcHAkkENgQzhBzCrTmMwp4q9q0+fOg6Fh5kVfwZPSCuo/kUTPyqV
4G51JOXsub8uTPcvZMshC547Dne7Ehnxy/9TrbKEM5tzF9CWDmyedisxu9dYprlmRCpfuxHFQdpJ
Qt0OfH58SHvsrm1YvS4WEn43CvHgnmP7bhhwGOg8p2s4gupkJzlhbFE7oN+MHMvpEbkXVNuB+RY6
ZuEXCUsoBCMDhC3ojyKCFVfG15Thb8EHVdcVai37WXiEsrtNSLXly5xOD3sC0Ub4V4PMxK7iAEbi
uxTgJrfnHwxuW7WqEZFQI8wGiXl2y2pgrUksdek1btJLnPHtMtcFOaUAi/i2MvdwOXVG4BOJGAst
PIIXT9bg9iET1A4Xvo26tLoZdo6cYqS9zOfzi/dcOEoNaxt+c9PphZYpZCx9i33NWusokVF8OOBg
RXHMtO7KtfFelgUH2addhjPLP9vCv4Qlc6P/K+HlSFxK8j5kCs75nAR17XT6TcUjoKIXy39bHpoX
nGAHzXpuiTi9PorSigjgE+MTPlNHI2CMAOEw0LF2odI4EmtWwaqzbO5vdpBWy4EV0IOp5qwJodlS
WLAAZIjdysbSCDm8VXAqtQXVLK0ZBXn6NTAi9ITu5PZtFWg2wdJ+YNDn3mj8CQxrN4i0OveZFaul
NH6yToMELXl0dIbzKWmCxFjH6zCw32jAJaQ6+71X8dNn+2HAl9Lb3m549iKPaDlsVqXOnyBpvtmM
TrdM+Lu8r53ubGW0n9sVKcSid5V+LRRVxsZLeDD6KbNr39IXJA5DbdFPGSBjeGxKbP2PSOrw7WaV
Ip0rIlAsrm0mHBQajzXzwBebjTrjNzF2HEIqJepaNLdqpEp44YN9Lq496CeHQD7psl+7Yk82f+Xk
ASYtFQdpQRgRaNqln4MxgHKplAtdmHv2wNu0VRJA4nRmh/hhh8C3gwYdzCgatdwtANkpx5eULkig
55KUCyxefVh55rZ/HNH8sKlDAMshPee8GeT32ycAM44PQjNYD/Rt24NQGKbGoBdhzNs3siZXdUnY
xqF3eQ5J2JgZgG81mm6M3s4t0cOtwqngDvfEZxQRUDfD5yCFoRiAQZboXUN/TrmSMY1X3+ZJp/Fn
CQOcj0ImfqsbrM1KAt78+0w9OIuv9QVgSWGCuS4AZm6z+kMAuu9yz+Ily0wnVmOq7JSMmWvgqoC6
vAfgnIM0HnI4bkh92Ed7kzJI4CuQHOKKFa4c2G3OD5rPn/HDmIYplmtkX+pPs8fuvhsqLbCbwioj
KbKJHTrgHEKwJM4oT5tDelTOPwW5FaiQCZh703Hh6rSuAWp/M97U1LLNp63U5VvRKVO1QtuWA5Fr
Z5qSwy8xAVu5Pd7IJdgGObuQE8/ZcNFCnePeTF2YADcvibUf+c5B3WGNMWhE+lXPkvqZaXGwdn+m
7HMqgDJV+ZBQuE9uYEX0TBtzq5pxwbhurYybtOScI1VOCI4pwVb3L+Ugq1lPRTeZaHdbU5Du7enb
D/Z4qTcbq4apuZVN5IMp1u3lXp2xAX+U5XOqxe37XRLclU+RGyRuyEOjpWPOFWuWx2SFyyWmV3kJ
jvlv2yzsVFYRrWCF/ZecTOg3ud4D0HMvW7kIvrqp1QEHC4zmSpuMIVNawWoqTaMCs5JdjKTu6M0k
hhoxjftJJ9lU6EHuGbHLkqYbZtxnNYrzof0vRlQWKzmJ+KFeNO3x/7ENwmbkmW/TPXxcsHD+PWBv
S5Rjjv9GJEIcI/mUuQTnsPIVZoEh+oOCk/LjcWsl1ZiOIxO/P+j5h9pQdvwl+wH3hgeqfBennb3q
7ec+LbOd5Gd6Jf1q841iybOJZIbiVH0nZncnU26jB46TvmKkfzYO3Q0+li1g21c6J9Gbiz8d2kSM
tYwEH0EXAcjJjzai59EW4TFPIGtGzJcvhCt39cNptKkDmHn0j69gcAqyLQkEKnRpRNx6atWL/drt
qEwxlschbq/og2jr/XwwX8qY2Vi8x/PEnlp7c6BpvkRBlWKHK/nDH+L4ZAZpDXBY2xin4nyqxl2W
WULvwWz3LOPnkNJbgPTYrD3HEVI7dSQfg+aUDOKxL1el5lLn5WB/TWLgWEQ7y6e5z/Ya21qHpfNY
aFiimNTGAYxOkLwxcc08AuROA2XB/+yNaEHJn4Xh++fQ6vbD9JP4SWqMKERNwNzCcaBuhYrjHuAX
7kKb5ZiMe4VKdXV+Nqa/qnD5ajsFPL5hyjBvguZo0NKlyegwEqgJp5blFUpwkH11AyPfzcwIMc4r
3zLwLw3NpMy7pnijBJW2mgTA/ZR2J4g/hOH4HhcDEIkM2Ommcy2k5shswd73QpzVNuRQIHSBblLa
978zPKi+XakD5wniMOl3ubPwa7PMc31DhLKroFGvLie0/Q3nM/Tzy28AfuJ4pducQgoEb9tyRmYB
LcUO9r4YnZU46DNGHI8NABSYWhXYSS2B/y5w2HVWLaWwono+sVoEfa0uk7c6/FYunC49ctI3kHfe
JnutKDoLDiAksg/6VArpiUHOhdF8BOXiuO6Z6PneTuOFILRfMdKZaDa4UqdmBsxtPpW3S7II0ZiT
le1YROWLwuMSICVPX064ZtA5+QQxaV8tP3PBAUbRlQqgVnC9VyvU7p1WPtuzhhz8e4JvLlJ/wNvU
qrs+x8Ek+kUs83MbWLRDHiDjBWUqg0PTnHo3TU86ziWnAdlA0XqzPJ4jVK4Jwrbnvf4W2dLmRIVO
jp070WMt8qxLmJIrg8YmlUpjLLteArEkebO8sxhjoeaVsAlQn/ftUUqGMWiM1aEPHuih864OMcXr
5vzhGqfsRh7wJjfdI32YXMpcdAyc1IhNychLmU2Zi5bQh9xZtbY4aKWsJhw0pq7rpz1xCRjCd0rl
kl0jF2Zp7F+HF8gAGLXotR4Zbp/y64QOWd8gaZ7xnIofwHADfevNjPy9vx/9OKXboJfMJDT3V89x
dE445eoJI/yoLNY4SJNxWHB6jslJT8C4eU+q7s46jsh2Yf1bFVPWJU0kh16v9U70/4ovCfwzzwUi
qiP3U15/zKXsEHK3LgBkloXqK1ILBb9smt4+L0K4lFFhUWhWUFez1pVM7uef3AH5vXX5BoAbrDL/
iL/VEh0/U5PYupBi5WU5T0PyUywjnut/t4gYiwmnxsF7+AEFjLp6ra3q09cGHYrKCZKOPLVjssI6
e8h5eM4PNv+pgxYGMIg/jcDKve9/ZxeErjmymksWW6iFXk2Z60nRkp2/SGwEaRRTDHr4AIvHWmZx
dqkF/P1f+mSDyWFMjjgq9VcjRXG6/8L0UtcCRdGiiH2w+9u06qRGrNOzhzZkoIQVcAXIqu5a8Vmp
lchTsJ3lfmwnGcaN2NKc4vYql2tZWGwktAaSNU/o047lS28D2a99wa3By8HLNGJLiw9Jc3Xo6lsC
1/wbUfWrxApyNa5NYkVGkbp0bcTgqMIT91ZTU30mlf9qubCZ+bb0kNtcqzYzJ6qPj0j5w5P0iHuf
ARmlqSJ/f7Y7yqrOYLEV22+PDuaSqXmalW8MtJtLWNCJHIpuqor+1H8VJ1FL+A8GVPYADE4pXJun
KKtGPezaeeogo21NMqn8EZOJSWyy4UQu2w/O8qlv2geL+qlwr7GSCJY8oT4EFBOv4fbgd4uuTwG4
Ino5rAYOVqeOc6h/HyxQoWl4ig5GCuOU+i6QvutJXiLCfvdva1607u/khLrYOxmrVxIppH1DXp1c
ZhkHR+ki8Udi4hWBkkIbqQbjL1dapFG3ouK18Tnmr5OJDZ3iiwnPLxKys8+EvXF/KeTyABwZot9M
Sy+ZKNNldXRYkWcDNGrG2LorAz6Tgo48Ifx+ruIcPo8FZ3Ql4HR8yluTAXQV625WH23qtRpTRajX
7XFqiT7ZQ/Ar0U+eOwaeqwIdv0vE4ANP4obYRQ6z0q7icxqE6rgYe/fjDUQ0Ki7DRE9yHeKLJGD1
yvK6xmfqVXzQ2zdktrLKN1biy8xFG52cXMsapilA1ELFdpq21xZeXjNOocu8aTao1HddX/dfXxc7
GmRCXXYUxkWCDYVVimGNibNpxPlXs7Y8HvzbL28xImI22ekauB0tZp/jW+4sbG6nlAX72Jh5E9JG
JU5kkD8mY1hbtQlrjyNpAbYYhqwnKY+WcGjw+/LGodQCSRK2/eUKUVshYvJhfeJaj6pB/xoNX0q8
+e0L8x7Adk5Tf7esE0tq5rMZPtV/Ermh27QiZQaA5UuoIafdMd3hSECQd+PU0eZPihMDqblcNzmJ
kYxwZGQtM9K6RiD9X2YF0nGPR1Eg+LYCP1vxhKxSWbcuiNkQtkOPN/RjPW9PHbijiRofb7Qk0YV9
zHG47/kjoU619ECgozoXFk3TnSElMXln9FKrvdCk/Ku/lRu1vwhBaUxQvNrO9TtS8O+r13cwv3KY
JiBpsMv3Svf8eeK9BMpGddXDjrWxAspamKbI+PSxHzuYptypip2eUMi6AEkXhzqGpvNSPTaA3MZ2
y5w4ENVYVYV8ZhUCfPAUqfkXsdytlO10aWNUodk8vemUXOvfiUBIQ1xw+8cdYZ2iiGzd9fGwAovO
YSN5LXkyDkDD5of/WlTV7z2k0zbRXUtpq7R0y132Aq23040lIAHX7IY4n1I3pSZdMLAtHJ9q7WUW
v480MFAO39TgUYzsdjCMXD5XkqXMRVKaAxmBeARz/QpJ+OsjjT3Ml4zxhX+CAnixdtPDSgdjMKeg
wUISETfFppMcQ3UZoXxlo17tmXgMnzNGw5djuYcfdIfNHHkMhahPKt00uqB3Szg5g0FRvIQRmPVC
lHwpI30icBRef1FR6mES8nRrpgTNiGF7OXBf5Rp5KgmwiPadUSln6jwKENl5FvK+SaPlNRl/JtZj
KhEMWJAQCoOQrObV1TTDPWs4D+gsOjLSMKnFqduZSHjtunJopoLg7p0ms8kZhemq58bd3EIIEmKT
TR/rFyEvSWxQdnQeDJukVkBfWiqx41Iucsi34JzS5/F48DRxuZTxGL42dqeTYgnz/HBek1P4lX8t
MMexhGrDIb+HBL5ONRntlkNPH2ROs+hRd1o0w7iFKN2H/dZJEBFqVJ4rYls/6TrK+30KtlQfTcN3
ocvISeF/TTYkeegoxuEHptPYsDwCgFY514Kl4BybTl1H1IKQuDU4slkilT6f1joZCaqowqvcuICp
y+0+7YHnPTzpwEbWVL2xk2wz8ZXV1oGai6jHP1R03ee+iHQ7yYaTBQvJKMX3rn6C51dlrupeU5GG
R//L81kzfrsC2GOXy0eO6wUXAMWcfM8iae094vGIpM9+mk2Gm5nppcleP4WG4sWBEFSpRCRsQQyV
ZHIx8dY3v5DShuhtvD/9VcITyyQZvoV40yXGCEEH0bFlB95Abw8cIJRHkAjzkpl9IilPmhz061GG
TNhTWBsXsnXSdNY94ZJB2B/lKZdc8QeiZFrTKnx9Y+I8USIR9+lH+c/+AOV89EIu6Wt6D2HUsQrP
PROGhYbr3rPm+9FLbVO+4G+98bnTOYcTgRKUyscy0tnhyNn82Pt1bvmijJZ2k+iKEGwoxrS9qaZp
S7fjo5jN60qFAlR6wWIdgykStBhBXt1xFtHbMbAIHdw/eFY0kVBV3isRhNFJgba3Gwrp1qrUFiVD
dPF2ibDVWPS3w0ZsPO0APmGIFcECRRKGFTp5JDirIEeoE1xvO28WGwrBYtB7lRkpi6JWYERiPMyK
Cm1sA8R5fGUAvj/h/1B/n7PsxBGMy6WYNPAkvNLoclEgPG1GBo9WLq3ToR+DjSDvBJ+QveJAgfNy
5SisL885WC9jC+x4tlioWhrhIwKdiDMBMXoWu0xgPRNbOYS6H1KCU93AcEOHJWpy37DSx1eppxrl
Ub13sBj8aqGgH7q/wXYEeNbhGHa/VXw/KpZFLMxJsXC70uNdsBr10Ff5lhr37o28Z/qyxm70Skdh
7esaaeLW8lRsZ0a1NB9NpGmu2+nKqE3i1wu75JIULmeywi0bISYt79LfInl1n0hRUahwP+llHzFA
GlyqVu02I+rClAHnhh4pvNf6rh44jEQvqPbYINyYMrr5byGjQhwoyLuRDZpna4Ar6GDe7U49vT6t
3CWkCONEgsA17ToIfFqiSYbDeQ47WHW/SQH/NX9s1Qtu95b6dLIXIm8snIkUgYAGmOccLh1Ou50m
g5SIybdyYig35Gfe+ngcn+raQBsqCLsZi6tW+1hN/JQPmk/oyvfBG7hTr5X6BkxJWLOHTtwf9v84
rMsM9nrAAxj31LevDm7GTsk/3KmqD3dUBIWq5si096E5WR/MIIYpPbXvyv35MWOPqPnNAWx5+G0H
eJnf3II7y+Mm6lpmikhf3GMFkuyrBjkNDYX3zL9Eyc29BSHZjzAFu1NmPvArkbftWrzaql+T6BCn
y224mh1Z6WDfrMydWY9LCZ6PY/rTDKQY1s0djICITOg3wnQUNqhAuIJxuVSyiE1pustVMlg3WLZm
53GLEcE7/ULcbJXp+0/sZ89j+RIYARt11Z3tdj51YVGea43LOvkln1Av3buHsP+mz7uS4wF9bk2g
qzTGIc7bhSgkLKWRddjcIgUVN2B6K1fYxsIKMatw3r1Fnq+X1QeQxHhe+rEhn5NGL+uWmoWtSYSs
HVMVWwxozW92Sgpr/PjU6EsOGAU1IZKJtpr4N1SqbIesPDFrr4qXuMpJj61mMVdyjeigy1kNE9xw
5MNMin18xS8ZGQHXH3pYBIfG45UQcIk5mOdzCosF3jj0Y7yNBrieVIDw5UUYHH43FtZ+HyNtPhYR
LQZ0uKlLSa4f71aYfgEgw5wqVs4OsyYZvSj3cd9MZLwLtTccYj1ulZeNLntGyRbIjHgRMdecFPg7
Vv6Ybf64E6AXUf9m+G9qY/CY5oE7EY2S5U4ryasTl2onMdOX4ykB9QWSIrqX0m2ROd+Rg1rIcYmS
h4LQpIzMdZna4MolLDHwzVhrzbkb3zHGVXMgNiagesSok2fOERNnBMLM0HAKuzh/M61U/Ma6U1Ln
P7U9tSWdP1h+1vKXmwyA/G6zuxvs74qs7+FRBj0LjrW+DGaQwRiFY36x/I6pgtAa8t8FY7QRzl9L
gbSGwpaAZ0IpiGL2dsRhxF1JttQEDUQZrEIXB4z807Yjneab4L/XNbPnKpM75PnTa4F6lvSC3jZ4
oqOIQQ1M+9v2q7h6uYCEK+eqfefySkMlOjkV1WWV1zuVyx6peA6WWX7KNGRhi46LIyMSp8xUxZgm
A2w8+tZUe9owqsOJNIB7tPJ3TYdIho/tgXKQ6uso1o3S1oEjdqYYDIxEQiEBMHJrGxdUyJ/D0lKP
PS3O7K5owKG1e4uOENt7JZpnlPV3gDjDE0tKVj3CTsp8Y0+5STbs8I2nKLTBH7/BaOesmtTKGtge
wdhO7m207l9v39pfRMJ9dylBTrmCWP4FfQA1LJlftPVG2O3/0j648VX2si0J+RAL0KdS+Z/DWkfk
j6f8jUOVc/1nEnN7fkLf+GR9UQkaDmeWZ6O87h1ZSahbEM3xAnnKvctcsUvauKQkedebeHEB/CLa
yP01AZOpZ3LV0v0xZTc8HbFVImeFhVUOZmkY4RE8vNVbKt61pjp5xjIYVIBfderPgMEUyF379wh4
6kiG4nFo5/dQy4Ix+pq42RvZjYVP0ryamWeSU/omWbvKHSlxS13DSBUXXDC/HZspSPwqaksBnzlb
PpDYwz0JtVFu/rYfEB/6PBc1lGwDqkkZEv5FDR/Co93INim5KNLhnjY07UlkZoEbUKxSBz2Z6uQZ
A8XljbuQOwZoqqd8cdO3uIlYnQFnNEOTvQWmlvp7yPICTuRxIepmhLzPLPhlYwMRCh9lxtN5TLJ0
f173mOU1u63+o/lqmLsNncaEdrcIzlicZay7hZywI9HIXr+y+VzNQG6KZoO74iGJeUjCu/q4gFIx
V3X10+CDTuU24PZa7Dqn+3RwHUJ54cAQFmk+hvGPA9PxJIqwQURlY5jP5afX0xklKe5Q+i4uRhHX
z9ScsDJ/Ty6ew9CgikytkOURhSvDFDS58ASafqeXrPClFEt5fkVTsnSmZngpZblOxbudxMv6pLKl
DbTr1C9XSNxYVGeW0PlQ2IMZ8PhDk+IrYw/6Wv8yQ6J1Zs1yh1A7/2TnqD6yzmAv/nK8jpW1pi2R
qSclkSCDsz2WJc8Aam76X+zWGdXqHd6ezi9G03IjYWzi9NJH7R7DoRokktHJh8p+W5z3GvsTZCET
BhtiZLtsMavS2YDIerSCUf5sw3Hzq4/gaCkzuQmx7G5+O3dzt3sBg6JQW02/cvme+AcDMIV92SUt
Mm6jGXzbkM+NjUDDbB5mWdn8zUU4byEPz0KBNlLUk8CJAtEiX03LQl4EiifOK0ToeGpH0Rhm93OI
o5jWJF2yxPfRaeJ61M4Y7E3jYs10kUXa3FBK2yJ6YIhiC7cxGglSdzmsuX+7CxRNo6Dm7QWob8Ox
vqwrgFGDiHVVtQgPyjezmtbjS5yzi4nmHW58Rn2LbiA9F5T1aWbWNpl3sDgdxj71HRMCj5EcdNB1
IplUse9aAkZa1+/3qoFZz/gPoHsjz3GACKY5XxkKE4rYqOd9Q5N5rzocaxxdsWUti4BjQi8z1Brr
jZEdEmmpza4ypkGOH5g5xrXQETDs+RgWS295oaljL14UArEKFV/tCdZqHGkXHf6DdsJBXA93kjfu
2oqfJ1KLVntzYsiQ1Qi1kTe3cyMqmDMETHQUO9gbqNN4BGCaNxymCoJF7wFzbofkcvegUT9iP6qG
QjSfA1Kzkhyky50ysQpmeCDKGMcmCcguJjFxF3qWLvQZTbwsYmiR9G3GgnyXYsXt/WNyI6Rp8FBR
XXjXMQa0Bx3zowPcalwiadASc6cbcSrBmQwKUYnc7Sdojl/AkdR7+9sFjVu5Ns/1z9RyaXhTHkxj
FouUWpvhpRYkSTZ+zbZySKms2mlK7VuFqdX5L9vjBY/eYeCKjqXUOePUQnnduptIhTrA9GhL46kc
t3SE3Kug3L3AW5wyrgwgsY60vKlIc2H6XiBL0QNQ/YcoPBR6M/3R5j8Qj5x3EWQU+A8UxgyFZrWs
iYh/WYZBCqMfwlsU53wTpT2fL/YuoLh8tvz8hV7PFFg8v3zlO5gXYz1oeSLUt1IUjoRqncgXORs3
u8cyt6MDwaNBXxWbGvm+17/H2JT9ysl+vSgR2fuLadOkmOlnR+PesZiuoViWjuGVywyR5OoGdRnV
AO0Nd8nbwrVo3dvsiBYdRVmvRTOfQkUS+ZhjgNn8Ln6RlRVKJqaMRQ9Nec/XCX8hoihk1k3X5XL/
oG0sKfTox7qnbAEE2tsYXE5UPs3FwmM3i7IChwmYX4if+EYiunl2LcNbouk/Vr/2D1F36F0mO7cR
jNAB7wQrvLnlGFvfQXtdQuXbTAheoPq3+keItWG5HVn4+Bl7LO7CUWTsGuVrk6ErGW4HMVJOm5Vt
Iu9WeCk0XOe5KYRaYI/WwICbIXRsnOYHt9wwiXpFQb56oWrxeTa7lYY18R/uKZc/ICjTi8PQPMdq
EzI/voNaennUOz9Jlx1NYDR23z2feF3hy4pkdjr5cgwOUQXjJuJIkD0UwnLUjpmajs7PEzud8rw2
AtlYMZKHHKPsTKwoLXjwH43hIm/A5aSjR0FYPyuOY7OeiMEFx4KLalnJig32PQEPzLugc8NWvZkb
O1JUYfqPAklqoQ+6UrZa6zlHLjIXI50Blnt/YBRjvzKjZzYGkgSfiTfNH/Q07Sss/q/QLmqKIOny
3eF71XujxfWcDPZL68HsnB5LsdVB2FRUHLKIFwi7NQmq1gEGZFvzex9VBwNFNapItuucOajmFyJu
GEObSOnuz6vadQi4ZqyYpQUXovX5QlI91iT+Dp4bJD0Q4LgZ76WZ7YnNWA8aJcKA4bXfASRWQkxQ
MniodumY1vAFdy+9CI0LbLrL212AJxD1tTkF8KZ+fIRC7+B//zR7xuRerrAM5tlgN5SrhRUGPEK1
GNSLC2cTSNr2PFhUsBB535m3uBPexs8NLh7cmsuq/DkcLwPAWmMwOeGTT82Gj+k7bzFx3O0gbtDo
OJ2WudnFzHGBvTWLoLDHBP75dNgcNiY+MCZeOfRSnGbNUzY4eHEql38QCaCBPwXLNEBMqBVTIlef
W/GYGHzMHRR74niTAjo9QW3xXBB8Fo4+co3MX1YHRl8X0UoEV1/uUccCew2eOU8rW9Ijwt4NVlWr
Lxck2gVGF+v0QCinBawxl9xY0oAdV59Ih0jC/SO9w2xY/T+BlJWMfBDSsdS5gONENisFTXB71erh
3W3TAMn1aPkoYdRno7swTywsbWMxxRDkU4IY+CbKwKaAIkjHtUsBsv3hzJr05gXdMQOkQfUo3r6O
d3TxCjGjxVM5UjRtR/9rqs0tFk3pKV4La2hZoNBNDt0P3N4X95Oeev0wxq3pneQdjNv4k0of+hgN
6mHpxQp+xoLKsi/Px9bFixra/V6Ec6N6LcEvgCnai0FMFm3PGjZh/SmJ61ACbR/US/jsNihQ6udV
PyYWNw20AefWr2K5YwFTGckS0F2n4FzRy07T8aiOxedWdEsBcMnw6LLU7DDaH6l2vfJzK+0/cVeq
K9h32ZgONsPIigpkYnBrUsHtyVtYdjns/fnc+WWvLlmehkdYBvSzEEEP4AOmAygtklMXQdf9DzgB
kDbZvVJH843XnNG715HcC0CGWg85Ts5Qp2i8Tvf/HvWLjZkZGfNZPMAe9lppb9V6GfkaIqf2DUTb
BkYd13ECGeXeTNyvk+88id5caMYRl4cZ3CYcnpoNnV1/K2Kv3feH1vTrua5A//am/YxFmj73rRa5
YrnegCrhaDx6PQ3yGPCvzlDxZY/qmInx3hLdSkuA5dO2IP1LQwRHPQ2lH9Pyt1rOOwpATmvQYG7v
HYhSYwOb7DwK8uDB7yLcfl6F6iZwdSD9LObfFwe/b0I5e4DvQ4S0MPpchViV+tyZS/GygSEuYr8d
iGqAAH8d7ZU9XO9z9x9wN7GDpnZyi7TuDAqQtxuY6x5kPp4oAgg4KYMbmUeh4FOMa1AyL/9LSQxE
ExPGMWnZg808LGlXCgRBMPuR8b4jmWj0AyaDJhPTOySK4KvSmjh2JZC7Mjlenke9Dn/lOa30jfHm
yj2DvG6D5aNLdw6TLOhso6s1Chmq2NYNAgewM/cBkh4mShEDszdFJo91+x2tS2BiM0hCTfCoUjaD
h7sS6Evziwr9xqz43+AnIGLRXgdmBIeMXPsBhyf8g7MKl36U/PDF7lPZtjYsivUpnIpQlNMu1E87
PJdx7D5/WQ==
`pragma protect end_protected
