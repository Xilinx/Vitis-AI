`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4368)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeybh9y6pNmr/yLVxw7bC9T29argAiBsrLigeOX0pfrhT5qyqh7rTUPW8zZ
jae2ubgHq4DuHjhAjg0aorlD7NHIFHeonxWrZpEQPqnHnklJQ4aZk6nZMfuYaV7i/Rdua8DXx27K
bWrkVMex7x9K4i3KL/dIsWNfrACYY8+GpZ6llYSmffaP6tTBaHRaMGw4jh1cjRsRPdGHxdeGesdn
LyzFrR3vv2VIf3z99S9xvyrQ7IggiTL89JCNL0p16Om1mWEqn1D41RWIAe/axZnQm/cYaiv5DzFU
xSVTPhkDRZixYr5x8GbLwCH+YRDRGPYTwC2NBEb+efVKTKBybTNY7cgK8EkQe0Ae4MWOtPAP9Z2R
O/a4UtvxV//9LVrV1c2nINCZSyjxPtGtpjtwiTE4jA+vBStPmoVkbUs/XGkakwx9F4S8HzT9Hucc
5/VkV4VKqBw3pdFVVYJ38z936ScC+yw5EVQMSCLe3/Vh4HEcIbnRH8b2xfQ1H9hsM0StyCU4VqZj
/T5A6enr3qekR+jE3Jb4HYaj+2JFBi9a5kbuFJRf+0H71t6PgWF5Q5q2wbE0fQBgX3TQQGjkkLVZ
9fAD7avuZzx62dcAnmdlWwZtIVHSx4nJ9iDrtehJleM7q6Kbt8ZZxACY5ZXSpXnBDTjZ7FdCYN7I
fDfsIWV6hLAylOClwXK1ys0+/dLdFvNn3VlebfgQGgl9LnjSfZQrLHXYPXqMLJgxJN/s3twufg0x
eXm9WL4hKOFkX/doCL3leyQ5gzSZOfX/E7DRjpxIAPhXhmTteudIXTKuZf8fCK7SVZ0FoudOQkSu
2+AjgeE8vd6pa2YkgVAhhmj86724N1cVdtpxcUXuqKf7YSyYW/c5R4FpvCukqx9tO0CQAlWB87He
afuQ7pNJue7pwssaUxAaVU2weAvL5bwccoNt+MtmypHdkgUP2PZzJassXrZuUHCpzrQrGirmPqhi
C+WoOGcvFxC8cNf/bkfaFDpGzvscgzuHmycGArwLbJAriRV0d18kTLEV4JAhN09RgBwnmvkusVua
4YHnR3i/AYDSReIu9Qkt7+hu88EA4BS0W3usWW+LbOYd5pOKgRbM9GlvfXxVtdlB+gvqqWmpvvos
dEgKzYwHHOIuJdLzl+Y4Vfig9yV6wZkr8xV5milQLmd38Mb87FED+ePLZbDWEgZ9p262ucm2dFzz
/ihin5FrnYTf6Z+hbieb9aGQFJDd8iZ3RC5pkiIJWb4kP2kWNI/LEc0MzGeXIF0jZYJjTcqFwK3g
t59FqI9hBkK/PnUZ4+Q36QGzVPSsVmi2LpE/G1b0VH52kX8BjCcaQnnCTKSIS9uLALHUeUDb4Ckz
njEyfxOocNR585L4LowILbjjLkCe8Z24kYzg5GMp8wql4Rz59q6KK/PyGyMhJVKJu3PL3itKgQVW
N4p5VJwBNIafOMtx3teQqFRNmbGfvMoHMsm0HWk1rE47IDWhfFvDLiYu94SUGLUYl3epTECHlMs6
YJJ25C2PPHsRT+fcrBmLDd50yi3KfUG4CHNSp1B4XuhiXK67/3tAVAPPi1iWkzXLNhNaoBI6imzc
pUvQM3B+/LTsVYbjkMpXM6A/NfmXD7NgDLLznlZtdzVyDkIJqLJ7fu4MBZixZFTji7TdQtU8M/9T
N5WMm9PAfdhFmw/Uk3rUfuC65c70UXNUHf0mqjM7SLqoyzaXwPmW/3rgBURPiLGHB6vZ9vxDfAkJ
m2zXHd16rin0I01aZ3ip/79qRsLYPDh8COuw5LnPRiqVrSXz0EFyzUbeQhddVHhkOGnedz+ZcpLl
J5inBwgj2tzNDyS9mthmOfDpx6A2G7RwWSmfkWufip0os6SDgQCsnWUEnEukHb8UStrXhbzvQ6Lh
Wa7mdJq+7VqE0uSCxMZkdZJNdnqdjJi7oybLMz8/QKZH6dXTjaUzBeTzLIpQKUO50b7+EEKEkMHn
BIei4JAC/pBpLGcF52M2IiXjzzOYctvQnRu3pDOG3fArGNjYi32KgdH8cxbb7wnXaQHT5T311ap0
c2VRNgUh2AZcNg0i90XLFSo6NHSosJjgpdPe0hZTkn8iwPTA3Z5fWFTBcUjdEp7BYN04Ed6k/Py5
fvbvfjKgqvvNLMDcLPTUohc1M8mwiGHvlZl5QM1xw+jWOQeiwNen7+guuMSkNK7/B+IRD9tgvu3g
v5pRd3mE47DyFcE/tzmvlYV97hECKNoH+sjyWcpDhl3BZ+vc7K6SQe4Pp6NnLZC7JVcKHCZB2H7G
37iO/pzBWw40NNkZN8l8EtARVM4ndFrf8LP6/huYCykbU4pTSkJ6TkzRH4rkyTe5w75H2loO/hvy
NyWDvLDEw+8jLJ8E5hsPwUd5SNr9IS+M/ly/03CWkGNL4LY91m6rRRZs8qNYQQ9+nDK/1zpgrJmB
7Q9/MlY96dWgeCwxkBgssHeMWP4CzxVqkuS2hYUjbP65qf+vnRxIL84z/+YH+ySIuTjOKn5yfpZj
S4CmNbflcDkroPu+3yoRbfz/Z+59mMDvDTVouq/A2zCYPjPjfc2wHjdxvR7SBSlLyFWCRZZslglY
s0lcebr6BBp3hdlXPnrypcE/XzUFJaX7okLdwPmLS+pXwch3VFk0RJx7yOMFbRoYOkqBmoMSCmnB
V4Jpy6ue3gajwRpoUXmCPGmkVbEAgWL1Bda+QPBDqexe0+oOr6jWjGVn7qtnvoai8OAiT6fP1y+H
2rVd31ivPq+IQA1MyiMy4iF6nZUz77XiOVzJQnUDKsGpY45JxOP6ZdmwW5Se26zwC44iHJUU3/0L
KqdaGdWIvdCmJJf5//lg5UYyMAY4e81D5OlrBNXwXPAg9YU5hbzSxGoYIpVZrlUyDPpiFWr5Ze4W
JxK50LYyFbD5G3+qJnwRpy6yAao8941qOa4r5l1s17Ozxd9e/WxIRSMgFyPUckp736Xz0EBkHjFL
S7Im4Mp5EbJofdYbdIKR3eOspUHzZ6et+ckfzj4iHoDDeNSX6eisVbr6onp0PK0s/GysmFc2F6A6
Q66CT3EPoUZq1HAdVKicOSG12Cj9c1YjgQBEkGxRWyI3wIcW51/J9qiUJE40HqAsSfqJz/X/yM2m
80C63B4cT+JR8w1qXQCJ5tNKB5nld2ReFrA/1bxitWjLbl/7SnNEOYPeP3pMWeAAfHay/wCR9ctH
/Qw5txF/IFoppE5FUCwEJpAln+mKxRuTpJNhKb8jGk2rTM21YKhsfGC7UGs105RtaW3FNT5cY5wL
VCJBDVY239MEAktd+CJi4X07HAE1IqeeomAVw79SzUf2LqKp3vkv2ZWwB/kdOHeUbpiBi+28ZEbi
7GtSfZSLuNkKgrUIHpQfzV94e70Ez+2+jPGOi5WaUJJ9tK5fFWphI/JhN6rFM3xM4lvEVHyWFvaU
nsPtnV87QhTch1+4rEEunasHt/WninrLvb76DklUE3iEP/tXcnetUPYtYS1Zru8A9AdrSM3xAcHZ
Qrn7JlBWJ+fm6ZUaoiYLQtoTAI5s0ANboobkEpYybAWXwBWHi9vFegu7VNKHf6xD/atC5Nr8KCNG
gkcZdw8usC+nXegFE2xvFKlTvpCEIK7VZBoxSOj2Ddx65GJxUUYChFqq04yoJVYTC6x7CDawvDRj
K8rSLDGy2blBczgHP5V5DkGih4I6fIKnVlSUvMOWsPr3P9bBDIqrnPnP4EqOkV469GWI1xl/JKHU
Frd0rzrJBp8Kr4vIR6gc8+OH2fQ0fcD8lAPTLo2ptXelSckLnSxfw2IjOhmXZD2gGmQX0osL3rKp
ghLp+KRXBsFSZkqbCouIDkpZ4DN2vABaShj8EtXzSC7Y+0GurVDwi/UYqCHtYZ/FmmRC7XkxvzEO
bnbNhx6m/5eNgQ56CvFabDd0oor7sVJijTEPLFR8jFjj9HpSLD3ZFz66bZLIaH+8i1xSm1mUMifd
vg1aF6gj92cJ8XevDQHkn/tD4nqlkzOvtXkgpY3Evc6kjL41BKvhiDOz9zhRGmC4I6bXo9YTtQx0
NfF0YuAwsD4qeI3QHT7UZr57HzUkTp3hhBQH5J7QjL3MymX3dYb8cQk0DaMEe3PWpr2hTjsMUZij
MEn+ggxQx9hkKjVF+IR2kWxefqe322srzoqSE4O87m6vBuC7wq8qs6B5zBoP5o3V62+2jIWgl9dj
m3kTGhT9Pbc8cPBdoklkC1BMSaTS1CI0QzOBJX3xA3ITt9/+iJ8pLPbVGW5Fsq9v+ey4Z8NlO0km
9DWQ12UVLtg6U9vKb4kLOc/HreYexz6A+dDb5pGeFyh6dIKZQrQ161I7jRem6egbpx1A4wtSKRIX
ZyjoAPSWu3h3ebZnaZbN3TdDRpIAuUmVYxTgevQjx8p3IYv33AWj7tP2bX/cHZJadN8ec7/6lita
EWl7J/h7aaEoB9DwBJGp1U+sL4mo4vPYb1xOfcXwRpQDRE6pjVuJYRcpxqPzBbMq0s6RasuZoJAX
+yBtTQ8k4lXmx/+YV9lh8z1v9fM9WmUyzCTHHPJjwR1t/helST11kiSM6rm1ZQdjHE4A5zA6u7YV
Z1LCrLhAR5Am2gBsxp0J2UHZK7ObK8d5OxCzLSeoqI856GijznvXM4Br4QfFrjC15TOeEHpL64PY
LhsYHHoxAEDQoED1JRuhDUIGkNzl6CVuG2KPkcA393oGnL0StQhX/sECuZw+/v+DDctLtGzUU8Dl
DFuOl9nMvYeqn9ZRdhokswbePHLW7JebHdj0FXtiCQq35zW6MgYGrRkx8lWHd6eH7gERJnKS97ri
iIQR2gipsF1AoOmsail42pBnxngZLYNqPflwGPayth74tn0Tp5GF/T0758gshTRxdSkmgjUDjEUg
rXQj2O4aF5zwmPJPFVEZJpkQcVDNndT3SRH+eRQEGE2LSjadMXbeSpLjWWGwz5DryDsZnoBNfXWw
+LG1eJ2OsV5GbTHC9h1SNrVPS7yvaDO8z3TtvnhvDfqwAOzvk8ga+k1loEOWP0byBrLOLOrVTNC6
0yHmD8/t+HejwMj7Ulh06tSDUzmz0xYvus1eiPsctiIqwldIOsSrdenr8e/fRUFKa/iS6aqaMd65
mlLWV7nsyOYGw7+1lR5WzTgQ1Yu4Rvg5eok+Ff9w2NYN94FcmTm1KYY4np4u6SZd4Xrs35K81wuu
yqadNDSQ8riMbkCB66CYId9D3hlrVAYQHfxsEQdNk6WA5jJ7iN8WU9XKgLlWKzlY4v+6LAnR/oaZ
Yqr+sFFAFAJ0hDztS7naDzfW9SToRFci84hq/LZQYAzAW/tM6ykMAUCWjlbWYPoxq9lh/spUWzn9
7jTiAcH7O2Re1187362jmP4uOmcCbULHf9gmYb7s8JDwD3yizJV72THf+XEQ8a7ULkdvggVgl5sw
Cq44dAKbc8Nrj+fBRkAtwRwBKAyAh8Bg/ZNSEOtLfxGAh+IZnxS8FQGb43/EnroQVbnJPY2uaBcw
PxpBIxhHytNUdEsYoBktMgPKxXFG4ohMAVrN6b5WAEJc/9X1V3VKwKY8SuHtv+DhWT9r97EKJEzr
dXoqC5/UAkrRoI84nu4DfMMImpQm0QyHnTudLC63YqKbjEIYtVIIBGbPlc5PUbD7CPKEm0QLLLCG
ty1VyQu5Y8DLkUV8L/DBqR0/HoC4aEVNljjOpz2HFTjXocD8hllcZIf2BUj4SJEjL/mo02fdCO7Y
M7iHbzKkfPtVo6jd7ZKuGqpiDJe69ObOuv9IwgzHyL2wXMYH0Hpb+XhU/yfL7GpxNblzaSSYj2C1
/ikPXh8aN+FVG1uNMSVTbvBgg/30Ap4LRvJUsRUkrFOP4SXC
`pragma protect end_protected
