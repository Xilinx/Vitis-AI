//Setting the arch of DPUCVD, For more details, Please read the PG


`define wrp_CPB_N               32
`define wrp_BATCH_N             3
`define wrp_BATCH_SHRWGT_N      4
`define wrp_ALU_MODE            2
`define wrp_UBANK_IMG_N         16
`define wrp_UBANK_WGT_N         17
`define wrp_UBANK_BIAS          1
`define wrp_LOAD_PARALLEL_IMG   4
`define wrp_SAVE_PARALLEL_IMG   4
`define wrp_LOAD_PARALLEL_WGT   4
`define wrp_UBANK_IMG_MRS       1
`define wrp_UBANK_WGT_MRS       1
`define wrp_RAM_IMG_ADDR_BW     14
`define wrp_RAM_WGT_ADDR_BW     13
