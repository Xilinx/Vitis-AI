`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
EAL1KS/Vw38wD3JWW/68sgiHXQP5qqpYKAWo6DWGm0jqTLeZBNdTfjK6OxBXBXlszX78G3hUm/g3
2Kju/T4DpBP/au7EVujl9Qy+F3OR5J3nSHK0BgiTefxBc2X+dl+/W8mMSpDPmxH6MQ2VyLYaxeUE
GF1L9JgVmy1RZ2MNEfL9mK4papGN6GpHTSomOFs/5h6S8MW1J7rINqozOPR/S7tJmLSmlNC/2gWK
BfaqY4BDn8YoJR0JRdE9Rt32WImbPSj4OjmikH16/9dcO4cTKe47ANPocwxsn+KUNL4aNzDVJKBb
HC9oiN3QMxFeBa6WMegNBMbnULA8bkld4IvGcw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="MgJGPigo8pxsrJH149hqMe+FRRdi3MlBKLz11rq+4oM="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
Hl1gS2Szh3WmL3gBASBPam+r0bfONaOhbtqrynQ0MeCzW5UKIPLz8e4LfEAdjNslUAGpvunhR7e9
1Hfep61o8JM/UPqGOw6m/2KFzqofoQoF7mmhJP+eBKYHiaNM6S+t29BAe0qqTrRNxDI/8obTsmhO
C1tO1k51esI8hInNV/LEqAaD8gmG/JhqR1lFhq7zbgHJ9zcY9L1bn+0xezZVFalbmIv0E8ExKBH9
lat5wwF7d4/vF4mmxAlYwbAxLQpvEsKrvWbjhOLBJD191sE+poliqxtjyz8RvRhNYbPWBOxMzYlh
l7EUrfQspcepEJfT7Wy8O3CVnRN4ezaftQvxkdrMPuUTEqc/ng9SOfNNaPwjrHjc/MOkRTY45Ed6
RAzRyD4Tdx8ZQY2TurGnPJGaGOwTTFpkOJ37Z4/QdW1kRFB5lfzNVbpt23OCr0hnVkvbUEosiWW8
1i1C1H66QXGCuAmM+b17L576Ay4neR5w1W7X0fH6GAL+4oZ3jeTwwU5+j8Xeiv4pK83sMQ1Gn/Fr
PwDwGF9fdILQW0J13GQ3TiE5RpfRMsiM/IifFt0lOnJ5a/U68IVemDhVtw/PNENjvJr9WfTRGkGQ
M+4PwgZd+Vx5J9EVR8vdFbaN1ckoDxM0m0YUEe1zZVXWxJHlq5Wt7DWrwwklpTflRVEFt+Y9FD1w
CBk6QyeekcUjRD9C+8OmH+HmIdA/BF/JOuWLT0knl/f8MLn0oV5DKUPQJW34R+p9N8MhaG/+6E03
vdml9YyBtXNWcebH+QPMcSVqf020U61T/CClMnYvON1W2nVPFrN1yBbYpqk8Z+ZmCgy83OeYGwji
4s1ZY6tAo6oJkA0CcjzS5be91EcIjt1USnGvJFD7MOQWHDImOAPYsPyZngNZFlFNcJEuH2kiFJBT
9e0+AwbZVCFRpnu5CFfh5BCv21X4jWQWbSwwn0g3Yan0tfSta9pJgNmZi0Qoq4kyLNcJP/GxgiBv
2ntaqT1PlrLO8GRIxDSWpAyr68dYCgMR1XA+7yII1LTHluwY/JtCgQzVjenq9hIcgJDIP/FP1xZ1
N163e0Jc0iW5PSuHrnegxxVxc7W2cUk1j3gjpmkDGZEk9lnUu7NnNYeWATrrNLNYPHjBBn9WIWsl
u4JnKF/EK3fbo2DXddIhGan43jj6zoA0nx+UywQICIHJPAEuARUO7Wn0s0s3UO6QLst+dAhCyDx9
rScmTb716VgERuBRY5F+7wIKLCU6WACHE24l0mJ/GJJtyUHHjdUcB5kEJoHzkE8ig+3HnVfevgHZ
6caWthdjOB6J0ecTzxa5WKb54ThGiNaE0bulcOsiI1K7/I0z3NsWA/vXIr0ppy5LYcxAWzXlUQH7
zmtUC52CVUdP2ZAogBbpcl/xNuSAWuwvRchxjgsHQ0XfPl1NZFGj9LLNfPiT1HKEissREqZDBfTR
oqDpd2weLDkeYRw4BjuvXw4sCrAxDlr9Vb/NamgESL7NyIGzyT2jpx/YisPRMJopD4Qt3B/B8MY8
4s6riNyhrTpqt7Y5XPhRSfjy7wdXEsC+jJMreADnAAAqq9VyF4riqT9gNlqZxuBcmFpEWXvk0ztl
98m8W/5uiLWuIFY0PRVIZ55z5OlIQXslN2eSzeL8d7u+X100t+dSMcoF5Gvm7YC9JTsKPDxOgN1+
H+ZlSIADTGaaPtoe8CXaAM+KMEruY3DWMXwCYTvPSiAxJRBevVSoeFkOI4f87WB6BipDMoU+l64V
qovBSNkkkc1ZO6tmzJ0H2RS7Ks/M5nZyHK6AYJQDuitJ6RdBkUmy9zacEauEQP4IbbxP5etnr7/L
fbrTMjOYtYtwXlA+7iV3chCYYeUpCd56v6GdvH8Co7/SDGXNw2hzwiL5lu99WqZp34b2qdiEQpV9
DBELUlh2xvvTYl+1P9ap7fzTnemWicKF4DVIVc2W4D9N6nUTi5SZPMPI2hEMr/svfZyXVWspKVxM
vZq1JqwKmO2Rv7VoCIaB61PLbCDX1hSxVXQU+fHoLcyn0USFvREi2PPbTCneGauIRqH0sDPeKdSq
pBAbBVy4Pm9OSipza3vOTrU4lySSfBZqEipoUcpvhWY8+HmIZCxWyXqoGwnEmsKHci07xE9uFzNo
P6cO1NN9Exp5rmmzVUq1I/YdNudCVFLWC9nYWrw6QJBs4gnekbOZGuhMxJwJ/NsQGUlHZYvMx4HS
dIgiIrW8BGizSkDMAkkpo1kQyfB08IaSJYtQPNRm8dV7JNbvN5TEWJFeIUgrvkFLM/RNEpNnPT6M
2tfSaKkT0EVM7dLkR6QxO7Y7bIo5B0PW2MQWXSZi5g4+ctvONYbkH4yxqK0UBADYjNc5opdcNzlX
jbMeJre/8p/foTpGUC3mpwGDLo8VqKe3Mj2FPDe5LgqzNh2GBqFPQ27y0pEzEjCsENWzKLmbqsdb
kdpl7ldQTFoJAGf72bRD2cMjHS+CWu8xSoLQ567AJYB2cbot0ir1zJTtIdXqFvxt4z07TFtqyfTD
pNdaol2nRseGXHg6BvaMlsxjcE61NtkEjPke56C4VTcfaR8Q5YdI0UecsxWYc7ETRZUEYoxDZP9l
mXLES60pBff48WCNaAsFbsCgDphJtbXyZHfDoXXDj7nDxeMebwAT7RtgcfC5CDZnEezfJM6uodzK
abXq7yr/pxa3RxhG9J8vAjob5R5vO7p9GfEr/C0Lv/dCpKNBWn5i4xuScZ/rp3pTwcLm1CNysgrp
A+4DL+Np84E1CaaP/EgukBCPYxzGgxsjYJMicuOt/x9s2nZ7BvVs9rQeay5+VjotH4mEL/6ocCPE
MBxYi0xVJgViyV4FJSrDzca33wX2TTfCx4OrhVFHKIEsh1BFtDUCCIkm/Ux0fyYuE5oryR3O17Wt
3cPmi1r3Cutz8aqKahXe9L9UdcrThONrC/Pu9ViZamxiOdvMptk7Yjr2hE99zy5SlM8p6uu0nbc9
u693ytxyGKI/tWiTjwyz4vh/DGlVjFmcblNxjQ6purNwyG4GdnuovXEh/HuH/YNCOUw3inNAjh/G
Tz01ysrM5/PkvrMEpVQL6qLfx/FHf/Tw1WnXAFwE/TXn5nd2bryZx3AL2cKgOWFkJB4IOmbDiNHE
Ah8RjEqoRu+/caZj/UPmukJ5cJgqKxkktY33X+TrASRFl7NV40k2BQmVIxlNect6EwnO8fmbNqnV
mSxaBPlYUKKN6qLmNcK2N5i9PYTdtDu0Wr0F1yH75Rw9F07X9haNJR60U9llfBd2iJ5/xMKw9tD8
rvEvJHV3Zp54vdegZDt8O/9hBozJJ3MawOXplnrA8MkCBnyKKgRe5ZCjYkjYsn6QWAa/NTycr5ka
M2TQzDODm17wcI3fteNEqs+2u5+XnmRpKykCjF+1kW0szs5IQfU96LDhgyaVGASF+V2Kwh/T0pTi
9QDbVPXtjREqvp/bmY2MdW2ytnoB91KlNA4CT2kkD1uiONfzbRJVaXUHeiY7Y4spC1o+0tQWZoJH
jrY32fIwhKTqthLH3UUWAtP1r30yK0YDmPNKSQrpxQ9ixVUT34+jBhLU+50PuzCWzsY65DVxOYn8
Qc239P+D2M1fW7MFI7THdTAzMtTTIoseEIWsAG4tM77oMfkSLYpfaPB4zyPpbrWwV+TjqXqHSUX4
lvM9axNQ27d8Qd35OfLGUq7ufqqpHcdk5JKPXLD95RiKbhI+L56/OKhmS6XuV8HUyB4tHNc6tvNc
wYlo5eA+6YoSdBlt/OVx0cqIapU3hyT/tGyxiU5Py0U5C3vJrHM8YiNmgkRcWQwdELuzR2ztM6CA
s0ajyro41Cx6NmE41DmtJX7W9EC2LPpC1G25UnoEJj+oat2PFlRnz8x5KkUKei6ZQCKdPGCGD/4c
TGG+iIe3Lele2AK8IuQSFg07xYcZaax5c2dni1lDkFde5vPIdxE/0ilkhGWF6HAOPumJAByNaWJ/
IF1FX+eL1sftwQQ4vZcSbee7x4a1yHh4U8zrqclH5J+oBKscR8XjbQVWGntMDjECFRsObxhr1+RP
l83w7Iw1VrnBqzS3ERvfNTwmsFp6PS96uGzj5Ay2cgAhIkqotYPn0wlO3bmnVM6+Av5GujlGpQyR
1J6h2LlkI087gBuJdTrpgJSIQvse9YdkFg0tKVJumo8KbikAD3HNd5segA+9Fah0uqB2znk+i4Us
RQchCanouSx+tgzEoZm5w0YBE/ODsWaAfwwIwWfEsxxMj7oNMACozDioJUO8/RJeyAI5TfJS+wZy
YhtwOpJIks3rcHVGYO+mATcYdQG6L9HOXOZdnIGM08Rvy9f4HJTCQJTuCw52VV/m+QhWdpOra11w
1TMycnfC7oq+f2lh4vGqwuWAtvsXN7P7GLUqc4eXvM3bYllkr+4Axnwc4YyivB1bDmgJbaFKmdSm
nk6I/wHvyVWwmmMlMndMS1g1MRz7aV2YaYzvplU56640tGYxGvG8I0baEnOfYpvOWebC8db+MiNs
MARHAb6B2N8rsIYkg/F+JBw6CQVHIKwx7DmJ9YbvRgrtUUHpOI0mPkaJQpbvglqM6lHyfnV2TVpJ
1S4/zU9LA13Sa3fX/l/aQjZ1P0AEqI/pITvHxSr/mLUsbqX4lcXj0BSbPv/+XixQJpuQMjjt6ROu
QyFoK2RBHIsSPTgBzylSYXHgQJkZADXtibv+WH7DtqLytyF2kOSMhLSWrPzPpymNat2HsviFpWZk
r8juspdykFR5CjMH3Y+rnCNaO2FJ8lWWCvjV0KOB9y8UMgQ5s/MXWpsD2Ne31KV0go6RNMp42l2l
AgniiYlaXnh/uNkiGfgcIJOyDoHqAIQ0FKLvFSA52jnwZdA/udefIKttj8z6ajYCs66QEMD+ImtL
Atf/GQL67uCSnQxUvpO/BaBQui0Oy0/tVxK/NynKYexMGruvZy6J1QE2JiGKiMCDTwP5cE/IxYil
+BqNP5Dv0uVSumMVXPwsbQEHS5dQrIAkZUFAyrOB29pNRrxu+slaJ/YaVpdZ54LubMp0+EMtctrs
xWzF9JVhbePLKxjgkLiwaFfcNvROcKB6sgQtwyNBDr4RgZnJisQR1P/5jdtMtlFniQaBqOzB7+K5
3Sk6vZkHJ9UII7RQPYVV4vFUSXmNZez0baDldiN32y1Z79edcmjRYLNfAWgyLFKVFIdkz8q8YCOB
J1bDG4Orv60RwRqCwkr0K/CCuHwZT69Z3fNiUqv1Ej8LAxuECJptK+OpFRLq2ayqtDpWF5+kkDJY
bAK4XG91qepGAI4NiFMitFEu1lkG9JLE722N0QlzBzsG+MgoBqAUk/abbUC5iWiRIc0aeceZxw0T
8CJEqfNaCd8+emLhRMvQllWw/1l0RKLILuoOzP27Efj4MnHbvkz368y7HX+JbDoV0sbcFMpZTNYd
iu5/28KTwHWg8dN1FLYaRUCOlq5CnUD0fTYjnk+bcwtF/2iOza8omtF2XW0WDy9awXhTE21C1tGv
BsI1l6ERLK5cz3nd/Q8XldOb4zzUXvt+Hl6BeVwX+wxN6xko1C9ze6b4YsA0KXhdh+bdxW5ALgbO
/eMuFy1POCxn8E/LDa8/6n2/6rz/1PLTyPgThuBCxMqulXmDbgA3c0NkzTVu20K/5Y8QtM6U4Cvz
AjpL2SEknzO0mCoMuxYglPCRcmO+hbRGAy1xJ4YMitr8vlcpqN+P4knjpI2ABWSMUivdx0m4t7Mf
HaMlQMPYR7lSSm1C/q3GB2efvPzXRP2CwV+sXMCAh33B9w6AuOxptLzpCPkRmb7JdFo20jzNaTwQ
3b3WNFjWyc9xE/N22AQ3bkoFHBo3RQSdpjC9j0EJdzKS5lpQP1DI188PH1uhmUMJCUDsOeoIo2CF
timklRY+rIpRjetRg4s78W0iWacoMwCv3abkdlqtBA33f70mO2w/UnHNK4UJkVTmPpLuf/Vuk/wE
VxJlgRLdd4ZbArLt6WVtpYycvLUAXNqoFaGpo02baXs02+uxaMR1Hj7bIFU91/f5RmTrMVC2BErm
uYRMFl6p9XnBdvu3Z/8T5g2Ijeu+Z7uuEIeOAkn6yF/RzktXmOKd9CzU0cPG9x+k/fZzMX7ez6OE
oiJOyi6aDesc0rJWAYGPiwAiUQwu1jDdAbvqNTuui8VaiI13pEfbK8mhFNbIOuldA8zI5hxy4b/u
qedZYy9+FF876lfy08G8CTjO9Sp+mzsCzWLcuLqu1Bk8XbXaSGRIqSabA32UT3qV2j5hTwoiBm7C
hjzBSEaCpid7QUvnIxnG27m0UBjEASMW+oLtyCt63TRJrzRR706GO+DTyxyuAS0IlglGcm77MSAA
7BSto7SGNDzMuFHCYU4ApQiLfUsPPgtdLLqcE0oApCcJYsMEW1AzjJm0jlrJyyVzbj9RbCnAM/fZ
o/2in4YMK9GezrfkRP+3A4y1tdOZnDWyHqcSSHjQQSmbVzBOt7AcFiFHxKQK9TIicXHP/xUp8Osu
v9Hb+TnLHmYLcDj4kphuusaD7/rIOYTNHevFo54uPZ+lSB8NyLlz8YtMUaFJMiFu9Twv/yX+WxXi
bWRpyL69RrwFfzZ+wyegxnRX3qcCuYSCWEp4oMKHjSMRy5syzzlwy5kkWDTMteIP80huh5zyBI/r
8YXzd6E8rvDVVx9yMxk7udYWhFuAGbcY3yX6KHOd9/jeQya+c25gBEcEehk9iA3Is+gsmSpLc8Fg
6RL57vA/aiA0O8XJSyX0uhCXMjgb3d0sYdVFustereMJrG5YZDPbPNTo1kAURNR1+E5xqyMBxHJI
Jl+4wGITRf20rk8TX5Y/fiost3+E7PZRbEN0gjXT530qujaCB9xz9xneFayLo8bFqqyGoUY3RTBV
ctn3wSVhrKBtEti/5LICzGqAMF719eppx5PXIpB7C4ypl7ADiVQDNKxjBzunmbzbSMhpEorHLXJp
EeSD78GRcwvnnyek74bqdDHZpn48eLNHOssjV7YatyT/y62dKLOqAnZbsbHs0vwcoWpsGGO6WGTE
E9r7Mubw1FOyUJdey4aLpoJUr3yRwr2nL8pkZ/wSViuHJ/QZ3XT315PsMFRl0OgGAE/cIOeTijJM
qi3E4cSv+wRcSBI3rCRWIS+/j4uzyqJ4tF3UIpPHxcYpC7oZWOhLqNFedXv/Ty3lNcic/Xtfl4j1
d7CQApk60TOA9fVm3ZrQKqn2ZyhZaDxSVlz1cB4Cnm+juNSXgVePTQ+bC50FnZjDL1qKtRfH9hSy
49LKEdDlwwVMVsPlh+cN822GdSp6qZNz6oTobiGG1nK1l/LzBz6jGkCVWIwrm+0rH7g+DQSDQolD
rU1CtlgI1Mnnp++TIJP7XkMNisynb5g9XJwxuYdbjY7giBzoaseMuKUuiHp30h5f6vzrywEWnqMR
k+2TpyUH7NfToxLy1caczemCemTe/oFQtj1Qm+qmTvTj7zRKRFPLkZjmriY+P/D6Ymw8M6JK1WpC
64qmYgfR7/ac/uPTAqQsF5Yj8IH/arpCVq2jcK1H4cvLvlaFv04h2ux4rALa3syPXhix84PSN88/
CvjY4qT3a0IoR8A5alW6RduWpIz2NJv4DKirdfApRnqmfZ69PgCF/9scCLyzKLzODpelTfnmk1+s
CZGEkPfJcU1dExi5EeGz+V8IhSTGcL2t3oP6nSDVGdDC9uo1eNRzDptjLP1Z5tKoRQCkMIlVhDNi
ZZjmomvsWx7FKsSjPgC4dd8eqIA6GM63L5joJ4L264jbM5LKJD038Qjk+81vQsXur1CezefSYUnf
pu5aF3kpXEzwxxXOIVOVvd7Q3prBlwkUYhGNJeq4UqzlJnZOyjMiqUOKKESIYSTbVSadzP107rz9
EPZ+Ndie9HxA4lfiy3a73XHUH09yyNdNYLETS+GcvibuB379XGGC6K0OJIH2ueTHgEhUaspIGxlV
2S5s2I7oBYrP1HAgqWHgGxdS+ZllD1amP/mb8ci8e/gZSTsKaqsR3e3hnUdIBvAk2yAVNTTCep0F
8bl0QyKD/zyudf/Jx4rLkndzs6S+oHF4JNGxCu9/BJgJT9fTTI1jpLqCKoKZfCuCnfhkz9c5e3CJ
JtirTzobmoFdrylOZHPUW0dodFeGtNRxFb7pbQXwJUyqLndjpaSYqtF9/3ahu//7A5YmxGa4c+qe
9qOlW3icTTZ2V2ornaxXeQEY5Y8GIFvEe1oT1dUFiyQYOLq7zoMGiul3WqZtszyuMGabBNBLX+EU
g3ov0Detj6HdeHaENG9Dkc+HMChlkypSHT9s9B+iaesOuaURH8Q32A9QjJUxi6hNW2U2IPYlnuGc
TulQL4SSnGoveos0lJ0alObuQkIJm1LQf202e/RMPMmdaY35y+5906RI0D3rHh3W1mor8k7MWwEc
DK4uKYzIcNF0I7N1kTk5UT0MmNRDLOhKtFQXelE3f6edAodQHhvuantt/sNnHgZYcKSgD5HGjk0q
Ap7b8LzaNetP4R6ft+UjFOOOQM/Ms5DFLWxebUdhZqjPus2CN22JB3jPv7m4b2X901kLFlPDAPin
0cUUPtcjKmCRtVxfchlMkQ5vjPCCfrQrs3hxE7ht0MKM/sOvM+UCkLd6nOfsaE+N8aO4Z95S6BFY
RaQMHp7MWo+lOMu39sPMArJAzcUYeame4wJxa45VtPrwxD6w3vsyv9z4vtSiM6ZQS2S/ih5naDnm
wXPZ2l99SLcYSO0kV7Rmt8aE6GEl15qSbhFPk5oKPL5jhFzOdGGhm/3026eJZjeZM7BbOvyKhm95
Ko9mXeTd5XPmLQt0k9SkPXgMDzg/Lzdi8YCu9kdF9nslAUxU/P2Qm5nLsxkHiParO8XUNNUPUm0G
Cq/36wI5FSg2mraQR5ZTORpoI4UiNNf2Ih3igVNHh63hFmssA33xtMiZAZnJxHBzxgnuMpMg2m/s
BAVkbK7WkcdITbs4c3zsMvdsUBHCIhxsn6kz1IPL/63F6ayZpA/LkKCe9IJUXQ73mDg2ejngEoc3
BitWPQMnhzmIFYCXR6eb3gPs/IjEBPAwyCsbJTa+VRer/8/xETRXc7oP7gbVPcyoTQUx91sUSAqH
E0ZOjAorsFdnpZ2/iPqOuOsfG2G0ymMNgi3RoJv1wCh0e9WiDP30fMzI9v8NH2UA/TwwBJdl/uaq
w/beJjx0HG/IGehpqe7WFVb7qqigSbvjGqlRjoN4uZPxUm1g1kBnQpbcWrNDK18FkcU/Jtil0ga9
Q6BcyhZk+8EjAQRmVvPNqFEqlt4VuJUDrkWtPhaB62bpbzJVVPfmOCoHM9d5rmfJccoER1wllXyU
6JIC5ysgYlu5wv71atR0zLJd+Ag1SpEscvCM2yKs24ygttKJzTNrUu5WX5geLRynUr4G3DOSl1MZ
3s3x2bWZFTQMQAnQWOrxrdeEr51PJ2eADs0OmRhxS5ckM5BkbaBgQMBqL3t94c7Bh3pAhbxrMTsk
yKVKpF9PhpPNsunUaZ/DLJ/XmmYi9PrjRDz9SGUM7czGshZhXb4WQzgGXle1b3XT3T5o7FYZi4GX
7T/DebxEEpYqr+CCnPa/tCl9F2oc3CqiDZ7A6/GT7A7rGKaRvvmiM1y3QTIIYjqnG6GDU0hbNUdM
D5cmWWvVJC+m0XdyHcv/pF/8sNCkN/6k1fUAbutttnTIKP8L/poCn+9kP8V0Zu18eK7GOFTadnzO
oKD93W4a5u2JBgygJqHD6yfvjWM4L00L9gbhD09B2LQwzgLHdl9H/3aNlLiWfXerYEaAbPN97cpb
oEwmoXIfczNXJVnQ2oHFnkgaPS3eBpxf/nuPMO8GxmpAdS5JpuXNOrL0lr9HA0//fP4sG2WullLp
zqKNf+LO2b9Z4RiB+p/+oRt5Z0sRHbyvTiCJXoG0s8ZX6ihdyf0Ey8X0gRO26ErL5twwpIgbV4Gz
8Jn+Moeb0Asvrxgjsw7nE0BEj8jX+n86CXVwVMl91KrLaLhKsBEOexjyeormSIZUaoKkmzsGOczT
ZSfEOuQjdx4GjyWHhwQUXChgXjblRKJgTXy9FUBEgJPeCoYKWVFXRaeY24ua2QvDO5yrPNYl2l3C
26KuKB/k8tDOmjKK0iyT9rh3CwW5707G0qXz8tFfYEbtgqMkiAc8/yOsl4fciATsEDDySkCmn2Bt
60+bBWnATOLHlh3dJC/vzqs8NnWeAL6+briEQCspK4LNHhF4kC99aO7Mcn4G9mWdM8WLj8T++kFI
0OvnmJ7QT8Q7Z9YNBgYgAb6NRn+WUgZVTXgEmZFV3DYat01eLj5zNiGJWJsVIP2IZS+nFIAdAbYQ
YuChJfoeGyu0jM+YEt9JFiTwWXOngcwbLH1wqBKkAf1Jr1ytmCk49moqdMWi7jZ44XYGbg1sbhqF
d5Bbfs+oNPbVJ1Lyq84tAD2HalTFT2nB29bjhmYVOFj+uwWBv176Fehb8YrmlWHahJ4gT4bTyGOj
iz7hU7H6HXtHmNTUdH078z+cruOU2j+lZjEBKjMNC6Y1vdpgSs0t7U95Bach9gAoh793cuy1NKIs
z6CHuUuEGPxTFBvPMi+Rg+h6o59XwgBEZdA5QCUy04mzvUoREcCVQIPDKUQD/rlsBcNlV9Yaukqw
LdSJfSa4sgwLX8BF+OpquVtIR5hlm1V4zk0ejkaNk2HBe9092h81uj8tKBOuLCzB6z01IJDBCSH7
S0fbLnLuinEWXE5xbShCvi2bUtw0oCxtEXxzfWQAQNeHrwV+9WcZ/3T1i2r9WUVgA+kVgmUsA5pr
RDRJAGkIL04QRyzu03JRNsDEkwM/UKCiZqBgUfUG1eKKbCGMRLq48cddB+YCQ22Ex+WBaB8g3ABl
TNtyY32RSo8ihiBDMKgPxSWZN0U/FJI4LQxIS0xol99SYXk04ZCERWWNN8UcdDXpA3kpFdDCcwVh
ZRlEm4LGnqiz+eQgsOjVuzkbdRyp2FTpbtMQyiMwk1QjzgrsWuaDhe+dspb9XoSa5oIlvkNnww0y
Dl+1wcqzLOhr7Bvga+4nGkldGBtKKZf8SIKEqqLu/0UsWPefJhuL+KN51yI3Ng9HpfBkrZvGAOd/
DlIR2gdLzivMBpkWLzW7kYBxazPsBxYzkNmODNQqzTXFkgplNYH/gXXHMp5trjMFugFos4rm2NWd
Weytuu2F3zE98GqW/qM8FqgjYRLxg9dHaxfv7thRtQ60by9O6rMfKMDivHQBhjJzNT+TPwaouxsI
AMpNkwaGFlkHElC5hFdWoDV6wd6L+2R+leqWxtSywd4fiYH/HVAmsr52Oe540qF8s7VTF0SQWGbz
ZBwz+52x9hiTTBRCdlaXA39uDLBYnD7h0yNLSB7dX/lGczr4HGkEQs0j8+Jto1Lq6YHqEYntJgp3
V5XrGXSezLLRbIh9JHiOouN3or3vIc0h27ybpzowE+wx31cHvaE6rENsYVMtPcAoRGVWFSkT7fE4
lcSVFJY+hafpiniW2JB19WDEScXG9VTuAhnfupHOPHKWYXBfSwxC6Hq4ZTScK9K6faa3tfhrTx6C
DJXqASKjf7pwfXUujGpalXaI9dUwP+L/NGRfhk9T1ZCnMZE3WJD3LF3wdnb28tvzdVE3L5AQZsKv
m2GWFNqTxCMktMQPa16vzNrvuzw+cYIjmC7IcM1N5cjJ/Fs+W8XiQ7uZagbM0gO3INgYMhxX5qT4
wzWwY35tPD0PjfHLgjcMy4EnM01UfTkGqbjRjOs+lIzt101KnSmWNVKzMvkzwQubGgI9HUd9yNAt
hvlwAlCS4e8fuu+Xt5YgX1hPIty5NeNJUZd69E0S/exzL3IvvRxhIUoNzrVfIm3eB3yuGl7KtDVm
PjxlCe5uzEvHdQPek133DSFBZgH4nia6wCMBqc3oGDZv19FN8zWAqOSlGdoQh5tWlkoJvWQ9dEfA
WxvmomtkNiiPLhK7zK7JnD2XAH7TgybzAkhInIsGzGNH5yfhsEuYH84zNXnQKnHGg2feGId1AM1K
pJiNlGaJ3DYE29cGDGnGz+crluwINSZ7Agb0u0OcrnDF2qwF6372zF9/Dtrj171+X+jPpH0p6ZvB
TScckoMvOtHqHN9Rsg37PEp75JYQuBMrbOImo8QNqax0e3gSaUymZSgqkd7t/X3M/wryd4jYcp1G
oVa94Pr8T9nP7IX27KJ3Dp7GogicdKu2OXECc/T81E4DqWCB7gbFSkIT3LeX5B/uKfmq/pdrGZk7
Gv4l3qjVoW64+zuLxN8LD2Y37SDeNimGFJyT8yac3aGPrE3vS5MzHpFG8uoDECaGlvVUBBfNO/om
9tQ4PapogJaD/LLVOdd+S7B+Zn4+gTc/orxGKVTUEEasWa+E3atvWZgLZHHDn/6fCHXlwxMB8WMI
SjRJcuSIj6ET8iCb3+ariMt+oSqGWAxzEZq/KfbAofeTUqWeMolJLe90tSGVGceUBfNkPMFz49Xg
9KqVOwkFC/E/HVbQ0jPnVp8VE5lBLUl2Ecamk3kMZCz2aUl7kfRH+ebpBqQ0oAZ+JS5v4seHM3cG
ULhcoHcGQ0PGDO7s+3TaGTRS32kjrboDxdW+a+3I8HtVkjZqBl+sog+r6WY7RyPc0O2Hdv/k3/gF
vFArRB4DK7Q43ebvoENVfl39ATQFXbd5pcpVwnqqphaCq2jpldTmnTsUiNfxekM/Xe+zRVHu89cJ
bZykrJ5MslzycMbAqlvjps2fZtPwWntil3YfmB18kzk73ynESYlYi/utKI6GUUqqSmpRdgvZMLup
Pg84o5RtS9KCm9Ba80d5yFUcD1Bvi/2WnBPKI6wwZMXanxVjWTDXPxXcjRUbUaZfjzNs3xHla2PD
Q2xC5rtZk1jJHDUCQQzBeJeE9F6azlEcfO+pdxR9p080uz3J+lcOQZPniOXZ4FUdeu35zAJ/EH6O
aiMNnxpN163jJgBcbCcVnZZI5dn/BioRk2DuSDjbV5Rs5tBl0lpYhzopx+TTikdA3I9by6Vlmj2v
N5P2okrSqdat57G7+UkfmSGpRsbDSSupwcg8yE4twEJBePYZ27wmUBbGM9fcQBJN39lqtk2Mxu3w
DrfQxwmXrvqaKBly0JaPILFHsKq5IO8rbtgtfvU7vv/ENbehmc6nTXJNbKrhgPrbrFyNLStvVT2/
SAcgupOewXxtytm2ez1Ybvs860+zN62rTxXLY7yB8MObNJUDtbk7862xsBnkqcGq40C3M/v+a9b0
l23tBi0h+rT53euhCXqRZ3O4DPCc7HlGGrV0+vJ5HPOn00qXQUer1790IqoCsNxq2AbCHQqkzuNU
H3i3wcfm77MBCRG4e8rgWWc+HjXss29PKig8jLmxjFS/28Lra9V3VA3WsREzzn7EZDzaxh4fcPA1
nYBPSxROn50/kC0sSNKYxgm7LLA2PeCFAv3r7Au0lVZz3XW0zuhNfosgFf6+xd0EvS5jYuny9fNQ
VXNntkCN9ZcEFC752Pw5FAFNIoX8XVR/7gqKRvSwo6f7THdv6VQMRrvP/c1ifCN9WvMkNPGOnWuC
bqwKuKHiDK5mRFFhRk5IxvzaXh5+jnSBeoM2Kyt4jnG0YPy3j46ucVo3sZrQlGvIRT4WxjzdfOMp
lNPiEvHOp7knsMsUvXrsRRRzw33QM5WoGW/bMl/+a5SLduYaRinSMHo3S4meSTXRz9+kBZ9olUOI
mHVGmx4CJQbP6lhQIP2BwKCnVj4Ii+F3ei008PFWys/rewnMlEAM+yummnrTcTW4QZgpCNu78PKu
dqFCq6/ownrmiWr7LxJCfWZWvyPjbHHmsBMi8HsPWLUDTkNFm/OHpmmHgl926Nk5c6CW2lqj7cfM
1nmwQx7+xwxemCWkvxa9IkyAZtwh1dD9BJ46wlFJMMglDAnXRY5ERgexz06LuybIPS1rKJQRATQy
k0ZPUrnRNHuDDgMJszPJB3PXB4DYZMCXZib/RK2pOjVE7LPk8344UAOAziW2UsSGCbfc2Dr1IZ6J
/m5OAmcryxNqlxFG1cbfTYeOUsXGoqw2Dfm/1wosM5tUpGZK794dIvKG1Ek4IMBQ0YNc+n5fNQlZ
56TPAg2zHhLk1J0bzxth/YqXT0vSjm5g/dp4ge+qJomPzCE+oxGKNYVm15+d46C1XkQqeYax+KL0
VkwJvo30nPIlSpIdjiOBv/iO2btrUX41fxHtdu14SF2nXfgHR6aNeLtj/V/v1Ju/ln14mhLxIliz
v8KcLmYNmkuub3nSiXDMan227mWhUgGQo89Et4RQxt6niMsTAGlxK5cg29k0IOurPw2aml+7VltA
zICTcypbl9oRO2WTSTgjj+7YRm/j+nb0lTXwkpGJ/mq0dqYt51ImNWLrVHhEWkhoyGWN0o55AzTM
tlD8QVa7RF9VfB1f3g/rzrPSOJKpvib0x+IXXtWLdY/krLG8idhxfjK7rQuGwWL/8DiF7lDFKT9Y
5iXooyluA72CyT3Qtgrl4OZT8uhFpLhycob9NdbPUu6v94DMInw/G8GyBiDDxgq3WdxldBmRsXo7
4wR12oO2BL41dUmX6ag8+pecyjIHWTB6URZDDnrnv1mTe3vlp6ZUu5c8nCE0bl12WbLpqg3eJQ3s
CYIF45KpbNNRiPfFL2wPJvA07DfOxFgK/pRlQOKzoKqFbrX8ElGSmURDn/A7QPg0r56AEOw58egN
xBHm7LG51Pyxip0bJAxn4ML5iqXD8oAxmYEvmobdVhdn3TMwZRdq6Bd1EsKJAL/YMTmJom4NQ4Sh
qgT8Wp5aNyFvtteVHHX3+VK4rurgzf6ok3v1rJva/2LDW1MPQzWpPLC0fFB8b1Ht2s1Vi99Vpx78
AMZnZ/89Rw1JwOuW6mgNOZLKTvQrbx7a9ZQRX11zYwFoX7Gy0Yh3jckxI3CKDWp8TiYVuaXzfMjK
nWW5FTfJBjWiHSh5bhqQKBs860wBeG84dugFqHmvsfcxcjloAmvK5Y43F6ULkdLsHXfkcOnSp8aG
163L89ow/5zm103Omi0R6hthH1Xbax+n7sIHRM03Y31C3sk5WUoS/Ovf7Ana4fVc62pmTACRup0m
QPPR8fGn1SpTXI7H+oqYcO8+QbDuNfOIsmkLpMEo5SH3Cbto3hG/UFFmo5Pg6fAkQYjBg0u6DPBy
Q5TedzRIZk8MbBbck3KZGqG07RrqSQopU61hI9nXSQixj/BpeNOAOLVyCE4nfkjLv4PShdokPDEC
0JAg4Ihh2fHMvXyMYXOELsQU8umDAn7P64ADYACGIVKtsfBzaJZ3SykplXPZ4+I8PPdH1z1kdfmJ
hOUDbmQ0y9Fdc3gOrTS8L9UMBSxcJR7xZQT0hFgqM9XRcIw4wu+xwN73kvA314+w4HV6RqimoDGM
tT2Hdkcy924Ktbq1LejSEdyf6mYT9AQ7opi7EIMxdZN64OocqPgOIaAjdg+fZdwUl+9aF32PXeFD
UrqQpNq7eDnOcCoK46sfrU2Vn95tRYfZiKSXcWlFI1zc3rDaUaBgit4Zhb/nQzHNztaPwnl5vHPY
Qps0h03Lea0AmxnBSffiKXdtgBEmFdLT2ayWpXjtX+JtA5DvWqgK4+K8wJFtrwrWCGsJXh6sMcMy
Nlu39Elke3SI4z/L3GlTGdI3Etbh8Ieh4qRqDYdPotbUj2OystU8Z33Z1N9sTihyJ4q9swsUxmjs
8Dwa31GvRsaBMxGzPJvdPn4vxf3yONnKL5XYF1sMN2ny4HZvXrERqUYQfW2wwz/+2cNQBYMMe5C/
eBw358Sxxr5RFG1A2jWQ1v6Vd98Wmd+D12ccT50iG2YuDxwP4hxLAB8sKQWzwFBQcRJQEgYNYQsT
A3BNV1Jfywaw5oDr107qlWS6/3XfHWAPDqqrL1CUOaMDY4Fb+QqN0NVhF3sp3Qw3EKKEk3q2RbB2
1Tz4AnXUJ+xEmHigLfOo9Bm0LdOTPLL/2Giz3S6yiL1USE+xrgeeYwC8EZ9EsUKq+e0bwnAiRra+
vK5G+9XilQCjvH12AwXto69xcd4YiVEZkawsad4A+gXMEvJPN6MWeZsRlUwROT+K/04jzNEnkcGd
eV04EZ2d1SCheaPRoPsgad4vVytQAnpUUtMpV/7rcQ2oAGneQWxTfDRCZd/WtfCbk3QDnnWun4ln
0x2QKEvQJMjjsmZQw2H80HiMiAy/cMZS6tMd9NrWmB6yHTXXHhhNxJ9nzqgmPrBMzhf40xZa4ScW
Qg7/u13pOSB1+iDNvmVLaWt9FQ19wk/lTXqyTG7VHR6gKlsdkuyW1p1DknNOwCsgVKMvPXeGcD4f
TOq+VyR/2hR0RzdIX4QLGNWe90zXHh01E/qbEtbQzUW83v7DETBF013bszs2DVF4aWUFozCQyPhG
zHFYX4OyZhKaS1pkn+iXRvy3MO6PmcD4N9cczwp3BBO8Gw+gdK2IZGDCl4Gk43136lxnPugRnZRH
2sIfUVNT2IfyJJymlNE3nwSt31F1XyDh06rmDg5m98BTsvi8ClKdUudzXTBdsqgXK97i5VdLCNAO
DNg0WkFamPot16MVviUCAvvq+1lXWJb2kTQvUX+m70jUxT38B3SdNQ/LdcEouhCj7WRfYNj81P5X
3MVNJbxIeWMKoG2pZCgJpgGcxU707ZKECvbYco6Al6NZapm+7YUF1CHmnEBN6pvCOxfgNO3XH8ZP
6ehEUN9adfbTfiRLl7J6Xxz8j/2paCXPEEUiCLAWvJ5bdjYebj5anrX0IySB4huWnVVmSn63T6oz
EIeimcYZO/7Iwp+r5j14Xk16ohUyMxeRUk/2NnJHaccLXYBngaEJFQ+dDlLjXqrGfsCT5Yj/TZvV
2F+Di7rQRz9fTRWuVP8DO2N9o2xo+jZuBz+3LhF4SPcZVDF8krT7iV+xNhf9ZYI5W59kCUZfCVPf
kf/rVNYe9EaTD1U5eDKhfRAq6/JwMHQV80QqG7d7q3Gwb6MGvR9i3UQnl4VScG9vZJu710FncUz3
D3Wl9U7zhA+OtninP9+l9kqBa6kY6UpQRX68WRS9KnmnKA/EvdPAMUslIt4eO+C9qrgig5MWJIOs
5BN00liKiTOqFeH/iiNlR657rOXuqDz2MkTNNkiRcrbzbHn8rTPss60fizT2vHbViCUWe32OacZp
GddNo6Q2/tW5vpkApwuYFnhEJZo1MGDCDkFpRRmp+yVV0WFEkbO5n6YmqEaJLTytC2fv0E5+KxJl
8qrKgz48+VBuBfG1kJlMGta0cGKefTOk0SnHpxz2XD1jB+9XFdV5hQHAKw0tUSsCEIAs9o0DYo5R
V7X82vULplwrRnhbqwFRycI13XGgoX9banNUwVRyhp9Lu3mLk59y+8MVIt6CX7StE1c9GWwTDOO4
y+5ZaqvPOYX8HVGUgAfnTYYYoyOfCzou9RlXIuItpXvNo/4G6LGdI7sxoDzkSuxrBeQNI+k4pR7x
KIS9Bl9ENEaPc4Xmb5S4KQ2YY+srxGntDZlSpuJ+FVbcfAhv+jldK5MhjcCD/bFeSIw9s+r34iTl
9vpZd1WIULGY5RnP/k8ayZp40Wzi+AkTb+vECRKOw4ZK+Edv/dKTnGMschgbVz0QfWalbrAZe+1o
tUNxWhCjz1DviKC+9htssMT2WJ1UZN4PVumRqEjXSlR16MmtJuBn5xh+fQ1i+/7JFmLVrO/olXYE
gZpQlE0ZqLPzsKiRHsRd7Q2UYPbcbxEFuC3MltQs3sdGEVReXN+G4lttMXVeap0TEcVDkRbrCNn0
1iIiM6Wb2QpRx+ItC4NqAb5RhZKUJD6sWqzH7KOBaFfP9eftNg9jGAWV+Ba6HvPL4rFq732Rh2T7
j+NjHmkONUq5H/iAXbCfbpQx75ylQlO8NS0LxZT0NSAMTQqVxJY1N1fxjARZelULOpNZCWSE6b2D
y6dbjnsbXj53SOjVi+R2bcoztuGTp/rkAB+Im7Vj5zU7NCJbwiEGPn1l44zNH0JEnj3ubu0DmtMA
7w11yQzqi3yW+Fa1Oi1LYorj4VGjJCdSgYA/CtPAg8h/vpbMcPpgYwKBPhfBK4kpq9X/QwFSq+NK
VRoH+RfdMbIfBY+EPhZqLcXyWKV+8E5xrvemZYqcc8Q2YfAbrlR3p/YWB306A1A7yypeqpXy2zse
F7NZNv90ItvqwCyHV9tzJdXANesR0pjIt5y8tR9jzSz19qQ/xsNTcaJgs25DCmzuVWaPGZF6lPl3
RuDEZjwkqbrHskEnxOYhb6wTNW9OsQrP3nCYTd5CoTpE6CybPou1wqPwcei6Qr637VqgEPnnxAR9
pCGozjqyPrG+Z3X9VqTqnMExwdzPr4OboE/HegUBEafxPSG8m8kF+VsrBJMRCwiOcg+cOVyAbd5p
PfyvZWDowUrIiXWESPhHo0jGK3CjnqDYA9zSb0NoOxld/Lk7iz1SlYc1zcnMYhPMTvzonKKjsL4/
NERat0V4jGjOKxH1sBrJWZ4siP/6DikUP1atKM3tcJCfXALuyhJOwJuowt569r3Vj3B87+gQzAmx
wBBuVxImmHpCMR0tZCLx7kvVKIPcNjPM9EW6rbo3pMft7xJo1FIW/+mCKPuPCgLS+r/O7At/mGd3
VglRzJlyy2vWsbsWwMD3DUXt8rTGm8+vejLx+nC/FbMn++Bj2rGT5vGrY+sdBJ99atUaq1asKXOz
k2GXAmKHvhJ4AjqQSu+iw+oOwAgIlUx5+4b6VAM2OY0RA5aXERlQltELXJuhIkx3LGXHs3HVfxFF
vd99QfIZdAsHKhatvXn/B4AlaUBYx1lE2p3Zb6BKd8hE0ZKPPdN3f93yFsYteVFRKICtdcSCPff8
xmd6MyOchiK+v5PvsODBGptpTa//CKvXR0Luv8t0RBTyLWvlpuBlp6RwySX2AAjj8iqtoQLhzUT0
hWE4AWll+XcQ6BU1YhhlcE2POvOhouUDDvq57VyeL1Iq3saOsABZpk68hIVBMrraunm9UcbvlX26
SrzHcENm2g8ArQ/2SzJNCX9rYDMgQmfBPg2q09bjxLLgsiy7dKVrexeGzB3JiuBfkwHvfm5qo1Dj
zkwcQ4UurlESzajFF+miWPw0KZHQYj4Ou+Pl4jVi3pkbgr+LyMqhacaVvjASZ59YWP/F2mPki1kq
IgZT0xryRYSL6y/cESQ6gxCtI6PJGMAjGILKfUKP075Iyi6xuoNDW8BQDslRR4FG2yIFEklpUx92
Nj3QQ4r/AUiq34VW366e9/BaUwxzwWr1RUT+1clOps7684AQBjCIlz7uObWOH9B5isVfoLjaODFO
Hj4mvRb0jrECOf7X8UOS0d74XHStUUWJ4eD4BHe3cnNTwNqrK4+N0tgyJSqz9he8z4E2prQO2696
KfUohUA2HZZJ84vbMmKFw1+aN5lWXNICPaWiX6MwVfna1Q/0EMKETp0EVUJsBMTLDmH15jbjZdcX
Cq+G4oIJdgDGzCVE3w6/MCPDUVkaZLd2b2XEdZrZP1J4g+b/7nek6/78NR4Z+L/7Hkj2EUbN/jsb
9nA48F3y/yLHgBrUROVXNV8JIdT3KjiRTk2CJH2OuMpQIXgj7JNQp5WlO32Xp5zVDl76skIFyKec
KOHgsdrX3I/FpjV+S3LM6S6uOZiyS5y8vOFz4TnZLk9OYnQhPvd7ugxBVpo/lz3WzyI8VxD0Ipxg
CBb/9Z1WO3zgmw68pAFc86rqLHDtJseJR4NoNt2vb78whHhqdESjlma7+63pKnefSR7RdqMpbzIg
wydm2y5Yud+yWa3lazUml3gtis7WfEhoffwCZ/Jir164hTnD8E7GGJMv03uPX+ro8NbfjDoYOnNE
OhhXsJp7/qIcpZRSfEz7kFhfDG5oabAbZZmaEtYzW7q9xUL1x3dhsB62ouOGt7rqBqeB15oQsrkv
U/otD0nCSIkfYzqZF4aZvjxEmAeovzeDuqNxbMkJpb2rOLTJBstR9ipFJrAqICgIGJFh2b7h2T6J
HRz1yA7j+UMjFQi2X4gKb4smW+Cou9Jdj7ku7wNNfasfrnm+16D+2NW0r6tnMP0qjzEFCbsaNHE5
Aby243DOXU/VlSZXfmjCTksFDa5mVuFWRQM9mFsHQ3rWdRWKjoMfZy89ACOmB+98UE2/+hdgdNii
P6RPvDkyHm/3f7FFDBmOvmsJ5R/fBlnZ5Zh4ofIJMP5kuEPM+q8QQpqVf9rSr248RC1VjLiFWgfN
zm+cXVLa6r2pOSWaJ9cvZSVwR7G/1rhi7zjLIgmTq/uHNGOAJM+BucD8CccdzrFRJUzcmAGuqCGZ
MQMCNc6Zxkzay8OSHrFAoUBe+aRotGuiPsFr1QaYslvTRT/2htkaZCj79p72gQwlOVll1ap97AOo
AS8A6X+VgxbtcA7N68fsz2nZoMguww66K8s3qftk+fxmqf5HfateTOdw3qtGcJQh3Q3gFxx4iUvS
l1vKLHfxmRo1DIYFSUS7e5fcv3G6/UuETJjPAowcdMGJ7wPDqacqU5kmBdvZ47P0rp+Z4JMAsed1
1Y8iRm3+ARtn7Hl9jljAGVh5GlxyeG1VoV5HioRKStNKzFBFbOeWSULPnOmOPdrBUMOSPD/O072F
gxHTDXo8m+9lNa84wc5qh+rCenKCh+m05YIMqbevDXS6lpcAYWQXHaid4GiMgEP0A6WuE0nA1Fpr
u8Ac4jdImUCUBkdT5FW5rgxGux/rkvWvNcNse3uBrL8+I2rtC+KGuli3gjNIksczrhf4Srha2Sy4
70gqsGLmvqpIpA/NZdw79oy62X6Hu19xpH8l/Xl0io1lu+T/DGW6dXcnBiUY3MNdd9B7tvXwplS8
dPsvIabg0VazFByoJqcNLU0c1uEPOQ81P92RXsJ2uwSZxfkN1dKTil0SMZGA1nTHua+NEGYUjRiL
jvrnfDtRZMn4fPV6AUxXSDMN7P/0G0gJo5BKHk0rENkcbL+hljs5eCS3+v/Kbf9hS6kh5wl0w6sf
I/AWpwlDq/7Gba4NmhWRbb3WdDdBmNu3i4YqohwO9hmnX2tDdC5GP+Ios2Ypk7KXC6iDTCF3fXYG
Sz0x+X7eap4iyWpYk8dyEGWuPDVk+dsbsCErsFgZ4U071CbAYY+YFRI5WgvgBzBZzCJYWC96ydIj
Wjk6twSf8+ZlDVJGZ/cEX+fKrcguiVdXWm6pRGS/4I06GE8kCLAVVb4KCk4jffH2BblJEWnH5Oc7
HJvzIE+6g9fJyhJZCNAdkb4xi24jmTtpovxBiGOvvNznwNvuIVDY2NbWQE9lhs1jCy5ABGUppfHL
I6TsKG8AUkMBHPDLzuvrjCkW6IkMv7L/t+jyGE8inZdEVz6XrrRlZXhSExmnv+ZX6CGwvnYX3JSN
0Bun2Aal4jMkS1P4NrMO8+YABn4yYWbjBsqCsKzNS3zq2fivjDOV8WjIOq9xofg9ktP7wbLGs/bH
Dzj4USEHeT8NXmMw0LN89+E/BvNiBZOu4Y+GuLJL0n9Ws6jej250u73/DigdA7LgcAmu50rvdo0h
i2w3t3YlkzDfaH8pVCUkxxjWW0yWvLCw0EzP7Yk1kSnRIS40ZLTAZfwyJ0CWGn/gT8AKYs4Rjl3q
WqXyCeXS+kywSbcDKHjDGqZfVnX3Q4mSIoMp6S+YnbFH6x4SZGc24iHp8TkOuzuNY9MY1rBf0fr6
QYg9iWrOvK4sXWXZPDdISad4WUxYL1Ef1tZpEvVM02+l0Eq5MMA+xOZih6hVeDBYiy5M4p3MkyW0
BBkelJv7xndtSMsNtDy08fM1xDAx7OQqZ0fMbu65h5ZJWMSEYbxDvLumWkaKLCW9JZZpPF2QG3vD
K+LyaB1xcFyqI2IUvmdIUJsd5E1pnONzHgeXGxWuAF2XJr2qrffvUjt7PN94kX0dnvbrXBhDptW9
wWvHKdpLmGpBTwzVRDQWDbAIYgrwewQamXFtQh0aVk34FM596A1lsh+7adAexyppGo/yypCD61TO
AkejTNBtfMb/wIceZwj2u3naRhZjxSFvpzMM7Z0MHP2C5rt7vrz7Qbm+4esXWnsqHoDiopMLCBJq
W3yYSuQ8T1RaL1WynVWUe2vfGn9kkopLszA2h0giGz9CiKdN0NdeV8zetFagijHjnZB/w9bfYZm5
zrEXGZXu0C6Cp9IfG3/0/+YGZpZY7EwYal+/mmof38ZfS4JnMnLy0Gem15H1udhU0AUhL/LB5gOB
tn5hbGnkr6tGqmIPvqkIVsbzhx7qeFAM429HmBr1ll9DOMiAN+/wZgZPVQEshtbB+20Yfjtxo3Xl
Hyac9QhzvShhADOphE9m7OJxYd4Eyyq+48i2ipd9j3ZNYX6MCijRfTKr2Y1NW0wsOwX4efUYkwij
6S9BVK6Rgqz0pneAmsFbY337UR9r+w9hdr6wLoemW9o7kqtLePbg7ybO4dzXEMUaVucXmwPuuUVQ
dxMT+GZoeSVkYx3Htm8JxV9KaeARtdES/ulopjAl5c81S8sa4cbm1Bpuroxzv1uQanbWo74QXu3R
+BC9wE/gidEzIS9NN+qz3TRZY4WiEm2amFr2Sgrk4Prtcxhy4rDYmfFptcj9iyRxjcv/t/Fw/0eX
k4pTKLxslmrqHACR0GsmG65to9Umb0UN68lFEnWv8iD8CXB1FOS7BUWkOIYx4bRUk/3oXnqL5Vym
rOUUeowfMw5BqIDasT2kTYlIbmWM66iFnrECKNerd0X9lDnr5HrkaPRjSVsaskB+TNbAgOu4Ckb0
ZnowF2Ly8DqpdHBFjx6UPNnZNxmPoq9KBw4URKRjHVzqJ3SwxNSx2zl9RuX33vv16JBPiOfEm+vx
tNXjiFp5w1aJcTlXxUvblJznOm8+741BmoVBdfhkFYRFjBXZFQJ2SxSFa2iJ/HN8Z0J49SBzxfGG
U5XrYynTbredVlIwUUaVXjM3AQyQxn69+YjRhbjeFGmjYJwwGBOVqKRptyWsEI3hN7tdT8oe0jSV
/wC4uN2h6zeMTb9UpG4ND0QEjl7Fou4h40IOJ0r7LX4MwSkm+1y6/JH5RBoYN9eij38E2U5FmxEV
qQSkdnNoyvEfHXAPUHfN3Fbuv+vwf67jJcxdIjh7GPVydpyiyLh8snbcwnH4xReEDf2FJimvHWaJ
CvXDNVJrIKj+6/NyrInQPefrkq1Yeov9vBpTvYIf74c5PCU4p2ydR1N2p9wrrrkcq0vGn+mXsi//
3zsrHV4ncoPIRd/NvRKZFjwGOxjSWLAeix+j1e7OAbBkSF4X49xQRQHcbzA6m/A/jz4IpPsFlRFs
sfEegfpde034MI9uVwudkBIM/pzkt97Uf/wcVAVQzouHwVZwgHMyfBPjThmdTXzUmtM5EdujXwL2
JAbIV5qN6IyYhgxqXSiEMuLqQa5X78ozKnxYttqi5SpGK4NnOIFZAKh4IT9U8hXkeID8NgRKuua9
qT9900S04H5AFdnNncCBuc6urgSUnQ8h/fLJusToiNBINfQHjgRDRipvOqG8HuI+/YUGTAM8mMHO
vwgGQuGn8jewl2xilmA07qBQaq4YM+nYtS9tzzJ4JXGz9gdOp7dr3PJJWRmf42CEzeyUnWwwKeoC
oM4bM7OOVvNlOa+v7n3LJwc9MRHNEAVCxV21tXUIK0YBptExETz+4+8QVqkcaHYfdhQTiW8O7vKN
PYIn9k7qtSMCbbQ+ER5PnwfF69BWLG24kXe1OqU+5W1LrgkQyuQ35WKTnwPmJsSirzt0PrYeQk63
UfhxPvuPDHurZ469UCCF/+Ev2LFYpc0vw6m5o3iQLxcKzx1u0SMfzyCvBy7LHyB0wfwQC08jT2cS
3co4bFXBg7LtgLUvefCx1oaUkFUVt1Ic5HCL19VLjuc0KJt4O+qmeRurnrJUfeFobNolNALM15ri
d0SSKDUutqsRF3IB6E+i3tRLQgcDNX1r1WwhXrsgjCmxcdnbRCVTRZZPdwiYHwyKs3NwURkSwU3K
7NPBgISiieA5p/vEA0nSIgtTMqVIL/uShgDxpsCHk9i4nnrGKYa9LcPrGg4+vsM2/Fy8KmeNKJGa
HBU+kBWVK68N5bI6C6NeHGJ3j8W1J2Pn2LBSTfCJWR0IJm4J8dkH/Ig6FzoFVQ4zEUOHT/9zavHG
uAs8/KYztQxFEdvRIfrFe1DmlBrOL79WS1p+s+20rjkba2UM95dTq0flp/74alyUx50Zh9cdMcaW
OZYC7KURf8rRvk6GFYodUSllK25IS0gB4R4aG9+pR4n2UWjj+779PzKjcyNFiJBnfHkiKS6syZJY
Mx6/5DK5FLmjcwYTqH6hqje0plWQCEIE/H0hu/7bvQ70pZ3w9RhrJPLwDX989t+Ze8EkOOgeNJkr
JmJqaPVi3mHnxfl5WmcJvCzD3RQ+gFwhWQH++yU9Wh6ci/Zfy3jzeMHG5p0YbeHj1ZsyAMdKhLD5
nR3t1Kj5t2iVOqCpigr0UUjV98ceOoJk8HAtg6r3UPyXRtVPSD7X4Dh7s2k0eN84Tgwrmrvl0TMM
I8M/Kpe61XqKiyQxfNCJkQc3gFvgXsPMbRlWe4P9KPenHLFMYyKNCAsJ/PSYfXUqcd0zTQBZb3Mo
La1r51c6VXNPAvN9Z3t5+R2JDlnEMwxCIMZGFOZRv3DCL9tAVbu9P9dZkLYVV6ufo8rhhchcsF40
YxqBhs5R3NsDXYyWwquKHpPIYBkL7y1EXqpPgMOKTIrIGmL0FH8kJWi0cK4W5HZ5ey17MObFDoLb
PtkZnirk3ZdbEbMlp0s0+7Jyn6R6AOcK6wXkZBJEUwEvbSyQowC1f5pA/tDwv86FISFJcW0kDUDd
6y8hUKqpxvH/SjznWTrh+wYIg+4HE2iig2xL1c2udjS/SDkSEgDsnijxEMZ/1tg42tzADqSkIVDt
fVAfma3O9pKeyYCszvjx7Qw4VVG4Vkzg9diP/wdr7CNEAMbewiD2OpqST5U2BQqCHb4F/OtR47q/
zDYb89BoRoNr8p74zgv23I4wZJgnmJJO8w0Msg4xxPrN2bBGHjlpgUtMyW46oQ8g91xpgPvtqY8w
i4hv7zZcIInQKdsK025X8SslSrsOQ983AZbwPYd+FkDDeRXdsWz/jcSjxpGx8mZmygWXL33VbnVu
xvV8UcoGw7X+A7HWT1WU3XzcrkA2NUTCfdV8fyzfJuSLfCmFk00ZkSNB1FEOIMYyJZ9sgtw5jZlV
SfTMyQSzf7hoRDvEaLS6pP7cWJeDlJQjBin8eC4nz9rbPamHDVzMyhaUOAv1yinmWCGKoM+Y1Nv+
K2SQc/pWrRTrAdAuk6+vxpT7bwLQ4EDfY5ydwgIeDryh9WEDVM/YOjEVdMinUAKNrr8IIr/fTUAp
CDwnNgZAI6YxVCHQV5cYXDNeIgH7KJLu0ozOujsF5QFmW2lJOc22PGCaIml2xs9nsoRJ4aayXUw6
wB5qTl0rsYHsGnCnw6ZS3dxSVjUrGUrRiptJE/G0t4l1yigXxuTTYXERUSs7WTa1GvNBl6cfRgJR
slvJx4RXjbTR/zDqBXGtqv5HX6eh2oc/K2EP8TlvYsgzfUDl31tpHXkQSpuLGFi1VhwlAAK/mqWF
pax5boiVcoKD4v7WCSbuPXWFckTYvrptrPixlZEBWykLN8twOOjllap5lGRJANhfMsKDsIMdwqxo
JEomeJm4Lfa91A6fe5taMZpgEFIV/eV6rdVj9fR9yrh73qR3809uyhcCx90jELMj8ph0snFK74+8
mXdMY/y7TAqZkDiT+c1k/JhsvlphyRjjeh4FOxc3QcZ4ARB9fuGj3eJTF7xHristCg8eRXJZFguL
tHrR3AK5Do6gL3hCvG2sL4TfNuyOxrWVAylFjcf1y7fTze0vdAnaAjWOA26RPHm6wXS3W5pfh+52
damv9jvTTE0011Xvf5hOjTc7BOCXVEw0AYPTLftuh4IzdzVfo1KRdT16mj5Rrxp/e8JOpjpbJnkm
nEXhaA8OKoXvt+KGapfVouLu3gyw0XRhYSgQ+wZuVvawUp85oYUjBDKmnHqDb6FyzP/IWoYK5nDT
DzzQ67HYyDmFvkCmBHgjzo6et+wdTrXsDkMbiTp0iPkQQlFECHJ7ygZFI164XurjrBrFCTq362I2
EqxrU51hcqFwcoWixh+WT0Ui6f2YhJQTylSDU1o5GSfIShQQqnvA8VYJ9uLY/8XfZP9zVj/hv0fA
uqcMge7xUCXpIjwz2uSWKf7knqNuawDPvR7j+9fDdREBhkgKEDVwg4M0fFAN47Z4pheKhieQ80hh
LJskaPcy8X4Aj9QobjTWa8mg/gCtP3BTWtM6gCruLQUMJxa4Cz3sH+dBftXjv2iOdGBQcX6Zy+Vy
dTQPMseWtwzkFvRtpprYJflt4dbODa7DhAL8t8CvKG6cOcpILKYV3/8KwQ/GRkIIXVdaZVgArs2i
PPxbquX+jxsWgn7YTBbt5kAcVm/y/oJ7NslaUaWantYWNmDr4dtKWhN9/+JZ9axp3lqVE0ueqX57
wDHpNNUY9neArbyG6UkhYqWQ78QIlrYT+8reSGI+vr0PJgulWpNBJg+sgM3lRud4ZiXDQVbDAlec
KC+X7QqIY4DXNocbJV+97RybhOiWY3JS8PNztuw2rPePOQSso9vSTuX5OYd7S7yZzX6vU9UNvA1N
yKSXtnksIE9BmxYPRJqOcqXy6n7nQKcFvrZv+Zdv72FokIOq9FwIXnPkduwayaptvNlnvIIsM9EZ
oGbxq+ksPrHLzf0DXThkVv6sQ42EnLPQcemvJGatBlH7CTZYG1PyvlTxZ0NfhbBA2kXFtD9C1BrY
WxaR4kFt7IlW4FIt4JjhhTV+JhHgW4PrI7RmBybZrgFsFw8ZpJC7KptlONS5pOVt3mITqooDmwsi
+9DFnuzar52v0pE1twGSmnHjLo8hgQlPH1r0dgfzmUglMTm4H6zoIPnkG6eqs+3rbksNVYG4q8Ws
+uOZXvOiXJmcXXX9on6qnn7ytHe9whaqETus0tmqLzvW44W4ydPt2cZDAm4tPbbJ7z/gcJEkFdp6
C2ZlVHqpdlKE0aZNz+AFOvS/T6rHkAsCn8PS/9vkPxgtp/mA+ZPbwsYwG3nwMoztzItMZRGLXOfA
fKmt7pheh2V0JAcMvcqKNHty6PpnUeczZu/sUTSDksOkhh76SDrNOGJAfmXrXFfStCEUSORLPPWL
+1BbxDYs4HaVA6D+daGjJcVnYKgcWfqxrb80LAAUZ10R94zRzVX6CN+KNpAefU/CXodmwbVYjHpW
NL1jlAeA9UPTpP7eC8BkWsZiummewd60B+hd3u1bPlbYNxJbXHmXnZoZLf8aIjnU2Yuq7/sH0OEO
qhx01ZrDvPgXOPdt/OrD2mpIGgchvej2tDQ0wIGM2P22639ESDeuJKKKLN5KOa6HSa5hsvNW7xFT
IOAB23/AfZopuDk0yRsQ/Zq/FoMbSKwYD1b0uFvy9pTQ5B4n/j4VCTO+AQCtSjqjPZtlOPFaciUp
hA0+ecDz2r0Ed8p+l9ZcmzabVbcMRJb29CTjY0B7yYYkip9ratslIqPQ70WKI6ZDMWUSZqzGI/i6
x/edlA/wyg2D6IcG0MfmmI61SjEpf/qLBrOjBrg6E/qccGNf94AbyvbTYBjtufcjkzTFpQYhc1bZ
J2AEk9a7kCLOQhQGO8SoIg8Gx0KH3VWGshouSTSukX9oBVJmABFm3TT1fN6Wt5Xbpf0EU7xuVW0o
NctJG/5k40TFoSFUMZsDdbQdV586CApp/+/hMUny7VlSg8ubpp49RY0x4aGO/DhiY6hLNoFsdaKL
yXl/LnHwUgx2YgE9Bo/QcfAUEhhgqFiWKrialYSM4XzeneJ8Cx9WG4d8W6DxJoLQRYKse6NO3F8q
E/pJ1+9Gs98wt3LuCc7isXfwuIy6SHnaoFNtufDYUKTRHvgUFkqQcYIejOW4tMw5CnSX2yyQzlOW
l+HOwsSFoChTNf6opa64P76zs9xZVHSh/X6i9jPtxjKf4DiZFM0aXptoNv1XZBjF96wJV1b2cioM
+gxK8ecKWBx8Vp5TT+7HmZGjYp+ns4UwJ44/Uw8mbnuGJRb6cbB0EXTBILdAPnEDnkpJojd3jK98
l/dR3PXPAcyf6dJD2hibgNGNDEDMXNbHDr6MgVr6NP7Lk9MFkSW4Ov5Kre5oE56MxlJ1wQ8zU+OW
XaoxNyoFiVuHLR93myMDTiK7I6d/D2MYtrfdG/c6SfZH/mRz+11AqXzQ4GCAFW29i/OE68qffCOF
lcaEqdMtp/O9pz/bj4Lzhqdc4m0hI7ZaqrHaP/wq2/ow86dmtFnvF0meKLwYPaZ78aMZX0A1P81K
9ziNsM4+HUqIZqU5P7pOH38GPOuFDaLQZIuxEGq6zYnaDEBS587JmkfEqK7FBjt7Ny0iOpTNUdcm
8iBGtBr7Vho0XTTn1toK5L15WgW/JxJby1eFgo5P9H61/xI/5oMOI3jeuivEoaFwkPUtJ6JvQ1VF
lr6fkVH4li5jvRHm2n8dgX+mR3iehSWSZp3utPRAkWg4fkFNMHKIpZr/bvMHygsyLYqRvLbRJ248
HxLi7OpaFRZGSVz8iZtoY80JiDk8AAA5g706JvvhRCARrl26lEJgaa7Q6HliyL+2OiipXRnPcG5m
HJBKoxW134cl4BGJ9U0fsDg9wq6x5ArjGO6YLqSRu86xesScBdUMqJc6Bjs0pVt7tDRYqpEEjJ8n
nm7gjrWpE0mav/ejv40dMg9mbE9NwOvJyyzkgQ/Pqles6O8XIQKBY9ew6H15JBnDaVyG57Kj0UGq
Xk7BMSNtD+Fw1PSu9xYfnNR5VLTaXVDaxj8eA+kTJ/xc5P+bs/rfRoHo57Bj60cCaTzRDejO1pM+
/HSwbwN9GHJPGB3FqJxCUqfofkTZ09sIbdl3EntiK01Bz4/wl0NBNaPGGgENu+DgYvAhh2nHFNgp
GcyRbfZBI0cf4Y5KDkHdlVFJVbsyFTJwVjcmQg8NIqLxwSBlXN5aZzaS23wnTnUWVoKNGRNR8JRU
G1tKpZBKL8R6GImnrdplYOtoW1+HojjWLvxmXZ5ycdd9mRPBJ8UmjobC34uPPSRDgpW7+m8wlIvR
PCjHeDpud4kbpNBYQvTXZwv/V/sdBNm++cmDMXhjPtt72wvBFimuRn0GtbXINFVQ4EVryBgqZTO+
LauUESgshSeYYAMA09Mbwz1oTsKFzIYNQhFbciCUUHb+qNOHQinhpF8qNsM6emQW7rIASO9Pa5ER
JvDIcfETDHoy0pENsOPqDauPSkIO9IQ6Gs6+kDYSiprf/TNfQGM3otBrqyeDYGvclvrdkoN+ZO6K
R5yj94Yf44CznkO9edIpFu4nFevBIsgGjeLE1H6WNde/y46wo8MscysxarTia8ZW7N/0BhBDSb78
hLR26eQ6L23LXeGT7Bi66wwHSB7HA5d4dWrfQEGKVp1XIvumYseosPbm26/vIToxo3eo2kU2DI+n
6NY1Mxw9aOhuBTx2NsZxw0dnh/MVP1BAA1MWGz1mO5uv1fnCM+4I9yVJABuuBgKAmLo8ZzJOnciw
IgDczQiV6KF21hUmNASkGIcEtm88zbedBL5b+D5A3DqVK6XsgIVdNuDaES49LosM+epT01qMQ/uH
k9cZQWtrZkyMIwgxeDpuw986zexQvuFTL40k/P67frB25UzSmuqAvQXx7dxOCDKIL0g2R/CfH82k
AkmxU8tY1rwDWc71VuneDVr5Gaz7yCp6TKMHPQVVBet4qsVJfN9frW2yMEhzGs75wIQ4HEizwuxj
B2KLB7Xl6gd6vKg/+5THG2Czma8AcQP9GD4wcooibAfhQgQsRGti52B81o3bhKvnDjWzqB/+c8fk
ShMQKxn/OG5cQ62VPA9OlQUE9hbLCureV+RKsbG0iph22vZeN/spa9dTczWVUk1M+B8h+uSMpgZv
n2YcIKjHGTnVoqQqZToyoyWhUhhBDwXmbS/cb3ccik3edWGMXfzjkh3QW/EDnXngUI2tETaM1eu+
8pn0FABPeSogtdUdR2ttHsdUAkT0T+fAxRu7PhieUOHDChNz9LpltoIT7B1AHzdneyFmI1QJMRrQ
5PRcKbCvYn7Qkj2HPUwOdxZjjSD6eaQsGRUytMJJ8y0xCF6Uf/wNTYInzUJkAfuJWLlDIPsFr3Nt
1scYCxzZ0yMMh2cY3R8jsbDCBi46misbMUfHICoeu3Q4XFSu59TzpLuhWRVJ9pPCWbNWrEGPlm8v
LcHOpx40ozGxYzO5giX06e+mMTexo/fqh6lyCmoiunaj0RbADobn1jCqSZdwmRS/FNbCI6l7PFMK
iFRzqCONq4T1EW2ZdwC5hywB7jgCAJeNwTcNnBm1yaj5MyoadAsXlRIJDYTYO8fFXmtVAExoWszG
a8N5EY2+jSTyyeQMTqfZFokCG+PKvOyrKo26JUR9/Zpg/sM6Dbwgv4s1SOjZGY0LvB7eAPQuGUK5
y0PadQ0dIy7otZsZkhSDrl9HSX7FwTUH0MhxBSNuoM4d8fo7ymE/5V+doNL0t7VmRLwJ6vvvTO1W
7LTiXMhRvdGAVBIloA453z7MR/vY2poSdcCPBPE0+26KN/qzoy7z8FVkdofKDrvR4e53VDEhvbxq
CpGKskk1gcWHgDmJPqg3kEX+jqZ475J8fGT43PKxj+gg30B/aBAGFUB8hFzuVRIV2II48lWr3Pg2
W49nEp1Eg7FgBdf9QJSihNWelGdr8gp2IMaDr2TbrExwvifdCpX3lR7TrPsrVmRWLmnIK+D3WbSt
G3onnEsDB3EI72HLnEQkM9xEZmfv9vVg3nOCoqu3CYpu+YY1pK5lI/wJioZpxIZWAXwmDcF/s4te
hy/vzUTdJQTIJHrGL9iZIhdIXUdz3Bnbf5sj+lKnND7UUP+nwchkHjD74NCTYylztp0JYW5b5PiI
efM63wyKpo4ryRf5+Z5/OBkygwI5AGuyzyRu34DgJQO7VKOXdKSc0MRgJppcHAlpljzOrJGKNDdc
aGmmeYw+YPtR72CvpgIZdhscEhNCqE62VX6pbeZ3p9Rqg9KIXFODuM1e+XSPH4gBHD4TQqwocygA
sTPgvd823QsWaz/FIk7xMlCzH28F+gx3QzTNlz7R9m7NWTEt9NlXwnJQ7/WCrB/4qpJGTLsvXkXn
T9e+qv05vIP7LCWdAsaESUTiqdWtGvkuK335TV8hHWsqzeVjBwEguOUMnDbNb5xOuRh0mem/nOXS
EzybOMaaMTLX6qbxFynm8AUoy581UKSdYNuh+3fhI7xFx6WP/+cm3BaKA6m7+cHlzbN6FJMuocdi
WTtOFAfWOI0EcHDpWur7ljsU9h9pa7fnAT9zpD/LFCI2Zl80PbfBkJ2IOAl5KvbCnChl7lMZC8OY
Pi5m4+90qrh9hhjiH47I1AHoWBI3RVgsl4Pqh71ltjlc+qaKjVx0UbCFOuAM4eFlH1207JohVypM
y3R05xVJvZQdIHz4wvgKP4LBnOWglIhUYNobk/Mnj86QTCqZXUEqN1SqmSdCqiSwdRwbFzw6XYWe
Jc5CBFEkRoebitV7lswNQ1/MrS+t80EH38QzkYmqXdirlUB8mwRC5dmKSem2z57bLImn5D+1IfG5
QZvrv9rGxekzzox+ntLn/NKrKhNYMmxLrKLjzb1fqj+WoLs9iX/c1fBkFWVtz0m4LArhlvOcSIAB
9vBXazYQ2dWRE0b055yY26G2zgOW4qU26H7YPZMmjSoliC9Gj3K2peKfGlu0d4C8tDKuWXw+hbMd
FqTBFO1vf3HU3xMv0rukxvZuEPG/G/nae64dRMAPuW3eRsgqsdKjtTZUVtxgzCcphz1MmD7WcV2o
u/9pJUNg6HNo2qYRZ3v8yyqOHXctEBf/6FZcQQFDCWD6JplFXFAzYeJNeG7HOmllcHkAW8NpA02+
hfB+3VDFLXgrl4rR0wVUWWkkj1ln+xDRa8eOoH9FYO3puMoHuK4s1OiKiOtyI6WzsulvmqUOwH7R
Fm0xrvNXxDiI7SEQmjJLljFe+ubw043WiofKoaTG6cwGuGPrG3ylT7O+650ndEGp25KlKeWs3YA5
J5ETxCE7NifVS46xonch30P/AIqo/D/g7zXa/kCgwH0GCw+ZlFVvKXb1SGwxh89zKuPs5PcukQzP
vZZ44y7gSmghvl8n08PhUKnRdZXfZC2J9Gx4yJNS7nVKzOiTg32KnnE9Vunocj2cOVhI2i+R/nQh
KicUmRrQdqf74YTDEggv3GLeNP22zOsfdCqoLsJtf341iFscs4emfVyHDmbQUEA0rN3+H8g2n9VH
h2QC3tIZ2YIP3LfFBm0rQESqnqnA5Y97Mk5/ZypdU9/KbjLsxZGZLSiKOCBMirWNbbSEwveobFa5
Ldaonv8eSIoWJ0yIRdZfLoTw3GnAGweNbL8oj55IEW9fx1WEsDweLRgOhGuhIPxuGzUbsHSo0DJc
qqu9BQpMoNdaw93AdzRDYhfeSjSwUc45Hi+IoP6KdRtEnSZylp6RI4XXkLn4DaOvjkfjq0BjEKRI
/AkSM10yQLGXG7h4qvQMS/ya1amFbkjoRr3qJWhvbxhtzYRHscXhtM95mql0X5bb/G5U+Lvu8Wrf
YkgQt943Kkd1cuEFF77Kc8vcTONOy0Fa3jlg1tedQQnLCoMWcFLs9HHKc+820FSpehrnBK/ek47R
O8V5feZs+DwXu8TYpXul5Sd4WLbxiW98c3exnEDwd1eyBwW52+fTYjzEDc5U1erH398lnPcNnNIf
57pWwaf5T8y8t3kCKpzuZc9I2I+ffd414MNejWKSgpspKmBjPODvLxWQaW61CEb+gbwhrSDu3ry/
T1VlGLd7gfNgzF6pnBf+hyHLaumV9b9xoLXh0NqWeUNCqsFZToiRWYO1dQWmYrhZNu3k+Y1NuVHh
0IpNMM7n7UuijleEya63ingdXh5xKKLaVisNmxGIBHI/F54gr0IRlPyn+gssnQfnrmRciSN6C6Za
QySSH4mujoaIS+lkzqOV1NNqPVY9sJ8SpI+OQhy94P6Oy0vu7uZLR5AuT6KRHxxKhDh19BnZtnBs
jApRC8SMirW6M/+20ZodyvSajM0wi+S8P+gyXyeQJqKNRN2GrKVNXNLOSuVJ38nVPMR8GoW7oDVa
JBBjYL6g8w==
`pragma protect end_protected
