`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24096)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0ihyhG+RjxpRi2+lE6Hwejnk6V1emSVM1XMc0wHM24nNFo4vzdO0B6vu
/7Bz/j2QfPta0fxXtKofEqFMJOVGBPh0dxSVeXxt16eHsmNt45lM4Ph/acDRMOcMDVvQUo/55il8
fuakEr2oi1dbz137NkmxmCUS36XydQ+Zbrihxya/PRAk4X1Qi8iGzJEgHXVasfwZHjYHSbmnx+bz
kYxHKFc5RIsKgQz6M/Hy5T60kfdorP/dex2CZd4en93qPx1OpQ6MhHa+FU2AoWbEPJhWVBfsxMl+
oUr2vYRJVznDiYGv1b/pfiG10wYrK9KKoqoAK9Fmmb6aa3YHiBLvZF0bymlhshLVdQn9JvHBhebu
fkBzuOuxm2kg/6EaR6XVcbsNmwWOq47VC6b2mOh6yiQ/qry6isGLF0MdaRMgdNILzVNwOdhN/lFl
4sWx5gxF0IuvTg4s4m01zQbpq/z95pLOes0i6snoMdaXT4u/ld79o1GnhFS5hlslep+v49I3EU4x
zOwmaJyq374vObltO6d605qNMKQkOujwXqo4IesGxmKFH6m00FHCQtrdjY4pf8Lgrrp5q4YhMk1l
BYwQOd+KfKXgcvcc5BRRPrzjbm4OJz72rtGrC0/kBSjSzdj4pgnviqsfOSldTtbtnQmj4HcTRRbm
E5DRVhQMuIPxjBu5jWm0tGr5KrwGIsZCjFy2zAwPY3TtS37enRyocFZJ4azZM42Y49/SPGW1/W/5
iBd7495hp7FZWwmiOm6U4+FxXVaERXQ1f+eBNDQ5SRSG6h3cHANrZoOkEDUj5diohgJMTGIXLYAH
r4c67K7BaS/79zf+sJHU6YR2M+Tqhu0VaD3+smfVPTmYAiYFZGljAWJLLwM6yV9RKOe8NOP1tuMU
m/PuJpXhHIEh0X24K3d6kXM/5CQmK7R4rRGTiPWGtbabsZifoLBGQwYk8IQSKkYC3s+vsoKkbUZX
gfqwhhwskrOEJ1Nq3ELYWAP2fulPYUKQf3N39mFeD6L0NRCxJS7g8DvEnmY7mnkRgkbLQ7WQ1gyB
TKv/fVIb9jtfJ5Go9Q2YZpOala05+l6ADoUMMxkvzWPHcDsAVBiV1JC0q0VUCGmXjZGHQUHEaRQz
4IrgwHOBFz+caWtAxQMdgxwGbckSnMaiZmNC/7rPGxYeW9Wo3D3PtXfIcy44cTYJ2LpSd6z0t9cO
7Sa7NfQfJ26w4ZbcNYQ9EB8kroMqIcqS3xMJlvHYSFw4gTObXmS1BKyzfYi21kONVqS4ir2pCKCN
P9eZhCeUlZmeP+MDepZU+6KcTnDyYLQA4jW4e7rmrMz1bXVyPyMdf08M905g21FcR26L7Em4GFxh
gGI1HXayWs0wWzEyJ++mA6Bsf3ALZie9aX7AHUx3y85Y1LvbZfrIhl6JZ5A/Yfckywyyx24nRwAQ
5b/yArvLA6HYXgF/sDTp36FuZy83skp9+69TYJHf+HgbI+yhX8gGGqg/YF7bYDkz0pshXIFRCCU7
z9ihY1g66rQK0r836hM3ShJK+kFXIf+7A89QsdY48OsMl6aJp2RGfAJ1jbf7Rlgb4aCwf+a38EUH
lvzMFNcCU77sQVxBE0YWbXBGKRidNBo0gkO8enuko/JIN0MdrLkIOUo4AlHeUcg1LE/jfveCGRCH
hKmcXQVxCcAfcCpugjtj5tFNAV/jGnlQ2YttKlt53LQU166qi/ek870bphu4bcbdbWTMPs737ZuU
8wyzDRKhP2Pu+7cVfxr4ss9tn275M30TzqCck8k92jrRn+dFLTevmX6Kb7pu/5IWfpVNRQiVi4oi
MqFREONkzCPdDGIFlo5MEA0ObF/uWOK0nqUWzYlDz+Xv1tpnbsJciwIZTRvhyz+CGa5h/LvW+28N
RUayKcVifY6sbVzJPussFuZxPHtPNWZKgcOHeLi0tKgwQXgx0+qN6EuLB0Xb9UABbwBmFKiCaAtA
uy0fghdxbPp404oSbsyiq3KRf+lprWI5Oq6W11RlusHRPoF7AJdJQZOPyq+yoiQF55xW/hFjtUq6
WJUAbOkJljXxa/MMVlxr869HrcCcdJf7eOwRX+QOg1M98Fn3dn6y8Kse4xAngsIcaPTMgFbSaLfy
JNwVimDI/E6CXhsl74w5kewhPTUWhfNh2tOYLHxmGfxGUPNjpwIarxyUHqy/Ia+RVTN9BRBU0C1T
aJ3T10VtJpVN1GkP2HCsemLSJxaAU0aRPz8NoAhu0TXpmsGCriYdh47gaCZzI5uO0PzvfK8eoB3/
sLs4z1yeuXEH78Vmxoiz/YH/wG+QC7Ty5dXvAp5PAe/4oEOupe1lmIc88+VSWp4+VGs5GUmqH3ju
uM/pih01ZMGj+kJMbWw9ckNitapWqGdfzFt7bUvuTAngWwfg+4MvphpwXou4zlecLuO3oPHCAvkE
/dtEJIirFaitQX32H3PYUjot4NOTPy6rWjUip7fw2GeRWKyoXlY6YXDUnCxextQS0S1F19WY7S5L
asO2rbpW/OMQGyqIVysh3TMVfNSXb063wXzRe47dXzQ7iARaZ/Hc9R1yWj029SsOkbVA/r5cA5Lh
3o9VOcwPVwpzpVcVmrYMxuBeCeDe2A/msSaJClkcvnuKFxSgSrW76ULW8PrXX8qrG4kUQvaRVRFH
BNq3U63OZ+XnVr8J8M5WHVdQGd8i6lk1nZGGwrMXAsJssp3Dbk1DvVpsXBgagLuKE3enzEnMHIDt
cKSk0YUUNjB9icjjv9ABPX372slCrBkuzHaakZJT3l8sHWNJpSvIG3kqkY0Mnl2u+/yVNpzoJwdZ
JGbx/q0q/C+AGFjCWLfCpZuIdOUEIeD9DdnGMVL7G+P8lAjSWBSYArBsx5Ndn0jRcpVrEliIxdt6
YSx3y88/Z6+YIRqWyCUSXrA+HzWNHpztWuqTGN6gjT5tl6dTTp6lamQfN6/5W4amwlDynj2mxdip
EdmV8Jv5Ts2YpfswTGC2oqallqbCwVj0RQvPPJdbUslGKl+OJcwi74Q4lF338EsgiXZR8G9K+bCa
w/izYDoNJA7yHehT7GmgmMbugG7RWBbAE3OAX3cOUv4U9tHF0k64juroMIIGwGNEOzCo69tsbcxM
tyx56Nh80GTs1oLRwsi5F/GLvfXf6QzD9P3oKkLtg4Xr3KRFhKOt4N2gf6GT9HLv2e/6oQxCgShe
EH0oNT2IMGuBEktI6Zj/4vKH7Z6IPWMf/ud/8cmqNV+4MzFNefURq7AjJV4ldZgXm0KS8p8UIeHK
hMyFI8KmPGZ/1E7+vo7m9iChPIT0BV/u6R/L7DOQlApQve52vO1YjdtRO6xLi5IAAjuVEJdB49oo
1NXnPFgT4yXP91WioVo+5zQJUgawOrOuVloU9nZZajHaHXc+Byc9t5iNPbKcbH+vkps7kkHw/SfY
6UUxRD8oTbS2jEZ3HhlEZF0m0j0MYQ3pWIR5O7Zf0opMtFZ7rOLOj89BI3mj39EV7kWni6MCO+SL
ioCoaCNEndfZCQ5RX6DenRXMEemqQAziylYwBOsEDphM+zrndYvck9G0ulhC3alvnNrY2XXk543n
7GknZMLCBDArLtalLxMnpXPDM789bls6yPDnUTFGjobxdX1YofdCDKKM00aPkOYGnlypZCuK7KJp
ui25bcw2NxORokFg/k72KwgnrEy+C1TkfCpHateUPlJeLZZJI3QR/T7IHgn6j0/gtSTIeMKSAwUi
RqiuUgaT3ZAsjfyG+MxD521BsIUcftCYfs/AAqFLeTlL2xSaDO6nsH+4YDrGed5m6AQtGGpdMyj9
POB+EwRU9tEYB6HgMmnbOfognKGMDN1d2mQ93lfcZKFtnJhpdLdNil3GrbwB1I1twSJ2fOfvmFS9
eo0v2G9gQK0fdJNJpDxyGES080PdjYnEzkmxqwpJfWoa9YjurqTr0Yf1qBw4LCENSIXylfzRe7mQ
t0PfOO3WhadD8+UtpMR1Au8x5o2lCbtVTtN2/lCLF1VU2lFQaKUZf0GSosJdpQrCDwPs4anVF6I3
vrHusHMMZ2EDQ723gqVDe8ORKEFAe9+31FpTZRykKz8MpC3sqCSp4F+iWUoAGhcmtV+hoeXXoUDQ
5Wlt+dXdyOBUScJmxI6qcIqYYAlGJmq2E0KY3s9Ock9/kBtmwoqzdPDjmJ3xgBfuKVDhrwBODs2l
rKVd+PJXP5JguODLyO7akfxfFhJ3bl//L4UMPGyY0+xLO5jEgwXoUx7Kb9d8m5HLGUWoyF2I9cfP
33slW7HVl1k1kL2c0WwagDP3bpK1ja1noP5pObCYQUuK/wJickQljL/+m0GdPAJdRXkg0fAd/t4y
reaedKX0379zXCHJYvy2PKpVv6g9HkDLfOxWViBjNCkcWArLGLYx7h4KOacxV4AOdiQu1qbMRYMz
liE62vHkWiyioKnEP9kYxTHt1jiMSHNUaCUU87zq8IWmJHyZT61LEg0gVOYioNYLclh+RibQrOff
SA7GTC4PeKeO5w1Xbzbyyv93dhtifKDszNA9GMiANRLvGmB5swrjcJZWdJ9esbF8nZEmYOnDMy/R
hvxE2e74hnKdv8azqAFjHkUa9URlEhFxUpcw4xFfJDDpsLXea+xHF5djJD6BzJXhJaJCQkc1jSP5
zBDDNgIzBO3+reCDv8YQguHMbTUhOLE4+zEtgBWDJfiT+zptoSpFkOZCgKo+5qpDj48pX8aIhdGV
hzVq7f/lEf/lCZAFwLNEwH0CuqhL00m9UcPsdh2Xg2RBPEwCPNivENVy3McToicn6wdLlzIps7M3
hi1epk0z5xDP+7owASv0Phy8xNB5IiSDbhE0a2MUPTDEd6Kv0I4g25PFXmXqMfh9/Bl+YFkVRFhr
a+rcCRPyrBDGFRBRiKUQfrNv+xL84HaMUgj58TnUbU7pU8gsrxCD3vPjH7j1DHIzPJX4O8ZYiy6s
DxdK0AWgHQaWaweMSWhGY8bgsWGhwsoDUd7jqOz8Df+Zz+JLHrWTf1/XxT5TQud5lezwJAOS0/4f
kVjNMWDu+ygCKGH2tbMB1oRcCqb3XxzFMPOU8rChT7oIwSgN/rrlu7hTCQ2/9iqlqPPaOVXILj/Z
17FwdvlZaJpcG5oQPppIUMChafxltx57f/O7XJXdKW4ITdbQwLlF/c+MT4vVZUcg8H8Dz3Wgu9WW
qJqazDXsdtNiGZTE9NdQe1fb6eJDJsUesfzfIhY7PBHoUfUTkSuqM2tSatAms4aXoLhjCYnWj4SM
N7dVcfx8Kta2M34opCFWYO42g5QYDYTfNoFgif27rJi1VOcf1leIbGcNEePxie5CZNDueZA/ouo/
kh9LcKXvx2qgtwTrCuNqEoyEbFQsJBnOO5oa0FwIhD9alyUh03UyqoK5matf1Ys9adWJwsfLyPvA
5dE79l2E8LOG/2IdEIH+aZpVd1nYoaheDlmJxqgRj+BPxoafeuqjJRo7Itn8twm3LEUBok7KbVaX
O51b2qPvEvEd2voFMub7Vb6wZX/mM4huScBvVFk/4vBau+d+UwO1EbnHW6R3yh8p6CoYPsKcT27k
hFpve94pcQfEW+CgguEMVvftBRR0C8vzcOCN0kbhjgopk+VhOwGS65WPGJE1wEHCdalCf4hfU6bX
IluzRuZfLAN5yjpgd2h95iM0IkXo59Pnv+HFqIQGaHg8tMxoi1miTl+9foeyD3mDqN7wNQfZMS5C
d5DZWoIF/4gLi/GPkzTps7H6cCckRrcKfnV0AR0QLkghsIlHQePsMeZrxHoy/HEpna/M7Fabb/T8
3AlxN8rzKR052OWK8Th4B35QWRR7SKVaDsJANR08pRqX0gMn2R6gZiR8JYhBYvon3kq0WnBc2Bx0
zeO26wYaGOECEU2WWx+Trz2zj5zz2G8ESupJqlczLoWyWw73ah6XxfkktGyRF8XCLQPxAjEzTeja
7NB9jzF2O9cXtmLfOVAnTolris82x9NDcDtegoA/ZlXcFFISb5amp3uk8cMkgwY/EwXy0DK6lGbK
28EeNRRybVw8+fij7ax6ohJUqFFJILyz0wd8Aykd/SzfZGFOre8ijEh3b/B2OHC53x/wNlDwMeXl
MKfuvxNtkNrR56bSiWC5pFOOtPo6FLWRzLYTrnTKGOuRGQYNFP1Oy2uHoXK1pW6VQ36uhEiglZ+4
7Hj/dHLUR2w0jDhFXZ9UO149C8mah/nb3sqwez34mWUwyp/XQls/CQgqLBj5R82afR1xT594FbNf
ykZ1dmMNfUx6OF1cbu0pn/kZGTrF/hqpx8a411UwTiC0J+iqsK7QAvV/6fZgmkK7/X0eVatTrRxQ
E2y3DLclMBKRwqPPWc2sNsVyfJ+f4UhPr7drVYadYrgSKmmtEhEv3MxLltHVgAsu7e4f+o0HaEVj
oCf7YlIxnmsZicg92G9kqiB6j5mTJu5LFXBLbXJ6HRfwirf7X9vBgNV0a+jRN6t63Lc3c2uOUvZK
K2045AdeHq8HPBpxQ8TZI2R8ppdJAUbtlslknWae9W7njEwfGvTR1kzra1RsfxMWoD71C0L2QGYV
OL8nIE1sGldLwh6Il8PSL7bzUoZlpf/iwwQB7bjU94v0//PvoPMUcpq5IafY89aQ9SkY9ErctNiA
ioLAVlwqKqVuJbyJUdkzLL/Y6vzMZll2SbZiWEZP+JD0PV0wqMLn/Z3ZSgrP5H2qxDHkR0Ls6suQ
iqAzomktzpwxpAqL5ltq6W+uHJQrzKXME4WPgrowEjHXxqV967Bl3O2oleM6X2ZPjdATdc405N+u
o4eMED+8aQi9tonK+NZfuja+UrhntxaE+T7CXkwAKZ4ct1v/D4FZXg5jebiffJ9knZKgFlOfPbO/
H1nHRJLiXXJwqKg7Lrq6qRmmiT3i14kN/5OVHikvdgp+rPLu87R2ZK2eCSKZsVG/QiJr0n+DccWX
AZswMn1fQBxzB86vD8hc11kAX3MbbenuM2G4YYtEe9rWLSTVqQhBnBU7vTKz/PcZXvBNVub5ZXiw
nYFtAOfEaqkPqQiLw+iyUGC+DcFLAxy7ApSxSNc7uVG/U+oNrhMVPMQFUgplUmMoVzC+5JA91DAO
OnVxdRwE/oIsgwjlbmdCnAVycDjZ+qf6YjTbSSD0c1ioOh/FDGVQA7p5AnkFG4XROwv3OvQC+YL+
+CYSLLvBbJaPcY8Yh0yPiEvvbLKJXK5Adm0voMOfsPXS9vdhRDW4nUn5NFKUv4FDOrEJDngthGOY
Q8FBaNTg6nGyqgNkQJM7g1jnuQR2KdWrLU1t7OOI/PXJjugIpWuP1dftXanEGdPq15EdfPB98ZBL
mSUfAevhsMsXnMqvm+yueQvHkXQ7xPFH1TSVMjSVzAQ4BP4L+YGD4UQVzY+maMqXX4mcoDUrjdWp
6sMB2ItDE8oeeVUZjW7KF5HLsYQdJtOlwRuZ4gIOlZ7mRjTRpWE7T5jRtkbF0X/V9EXMDSojVXwd
Rkum7trII/HxlG4Z5AZje34CWNuC7Rk6/4z1HWvf0aYPH8X3st9o9jMVBn8Ns8oMBnajiryXe2Rv
pT6lH0iKN5p3Hh2MEF7ftIjew4qzUv4RTkdBsdJVkFk3xcfQFvmZWbY+vu8iSck50POqnTBYx9WD
OzD12jCIvM2ehkun9aVHA3Vx/ua0BmpA6ahTXOR5m7rg6vipWtnXOyih5u78BD+H91XFjJOFMzBx
Y4rmbaaBLTB/VNpjncfr5OsriUrmNmTPFwCypgesjwh1H46qtcDap39cHgE/Q1pE7JAMwSfXQ7ta
3K+VX6eWhZVjON2/OflcpXcp7UfOySwJ6cD6C5tzgJWHcZxuZYuPuHgNCScsvZDpa3TZhNe9wlAC
OStINrb6D+rlmOn+a4Ct8Syu2y3Uqmm+PfHkisbTbfcjGf7zpOj4ppjHsN8lD0I4rq4ZkdydZFEt
uR0mGt0uHdP4CwoNKKvgPxxiM3EP4D0a+mxNVv0IPuAD/K7KLMIW5P126qEWkP5A9NO+6+TxOz3G
TZGLFb8rdNoVQGyV1/eIvDGI16qvCr8v/tAQf/xSAVy9WgZthNBWDVJQcpiwEXkipm06N6Aw/N7D
Z/Naulcd4JiFX3Cw8dp+WK3qN0naYQFyAvAJrmAmhxXWTznwayIIpCPAGjvjhpqHWOlqA9XXAyvt
hCC9/2cRibcOXz6LCqt34SeWMzWW277MZs+Sgqx7p7MKwMi2xy5FdxbuhhWM2VUyibrkskV+1ZEB
0ypTvO3gLGny0gfPqlnPgnMh2BCy7BsrC9kXoHOhZpWW0mwjzyh9rmxE24NhlVzMFP7/GqreQVx7
nLaVBLLjzFBE0ldTBZ37mE6uHu7cXZ1x2jiPkfNemt7Qd3pjk4qUZo8ORsZeewP6yPbMDs6z5gl/
A1KWkCx/sZ4K2xhTs1KbJvE6xETnoes4inmcaglo7kTMKRWuVgTdJOZH/BIvffyNVppvPjISRiay
iNSS6PuFGSaOu+GePy18byulpDx0Emwczt0l6vxYlwEby2QcBUuS3kcO4pPBeXjBFl9FLj+8nSsn
qq5ITaXIlm0yvy6QpvuuVjZYmOBUYw4naKRhygGqKJibSfoeOTobweVnAJkxmdk3WTIjtZ4aq+nh
4ccaJCUjOdKtyci8wbxLVA7C3fnpbQ8jg4rQQ3t1/CP+s/GiODv4Rn5sgQreE6j3grj1YcW9d5TJ
7SZhuEMXJnN8oKAWMn+I+V/UKrWF44qcSXBhf9daQQyrQBG2h2lIhgqChpNjrw7KrPVDU8HtPrt7
IXu9MFuRh9DyGnpJQEwKwV9JvUbmrnPM9Ucgz6lmGgZaKJMjK5yi5K5qI3fzYUMmWeOSSyKsj9w9
4MgEYJjah1PtvRSG4pvot9QnXh6j5LoQRFgnSbsq+I+UfdkhrRsdBY6oR2WadItXv1x4/tNYnm2h
TEFqbhOcOUWeihYMtkl2BNpiU4rLCJUtpk1htpzP5my2ritegxHZlVHt/hnemedaDzuL7We30woa
x3LBWu924rcDv6KOdUzZibdMWLpKVLl/BNmXjEjqiT5j9WeqsVwuZZzjD6PJ4keiKn8yTCU14r6B
19Wo2xs6H/1pL8sC9LoljT361XaFjcTLMJUQ1aKPAooKkb2x1XIpmDPZPExzSAUgDM/679YOFim4
4YrMwnqYfdgHl1zDxZZSJBASn6+5+GwSLKaFsHjehpgCs2Ax7zwJVrbeZk4r+5ZX1g6LFMKPdED7
UiXE2Dwy0Chn9nwBprW3OdbOIPhqZ5ahRvgw1vssA2s69h0eKYta7SSY7dslujqv+bAuEK3uQreM
ZzrL/Fxd32jzffZOuKxlbgQC7Izs4uLP1Et9hWYXf8HNGxUWFgH5Ivg3TxxzttSVW5f5q6xWHAjB
FqYOoinl8q4A/vWuhJXkU8LD5wH46VJU4ZDH7kqp0FE5fMec5X7/E2EwXTgA7/qKZlwW9qoe4YxO
390lecyG7p8IYLRoFjT2WXKZMuVMFDfxkknsW1EM81xWP4aQhlaeXhcxp4DWZ9dR/57ZPkMqtPZm
whF1YR8YMargKEAw2DBTzcmLKDlbAgnS0M/0yJFrX/GfWz1X/k+FZGHGrXmN45lL17Q9gLYO1zho
PLGRtZbHpnE6aZXG/eKe+TklOgO8M77BlcGh/EGWAD9plQ4shfW5gj3cQB5RwIKUIJIH7xvrfBal
dAjrIjy+2XI5JuYkEgJ2wOfBpl/ys3Zac/8gLpT0t1KPiEeefpcSY9B4h0cUc3Cm8995S1wIoxub
/ysCIDDO5YUdCgq8I8LLB23caeKVN9C+OmHzqcylvnV5wlvd8Jh9bUYLKXuYfJFLwNtDtEgsllZg
R/VhvoS7B11+iaZM7awk6/XfV6D7IX/HrZqQSW2xvguQm+Yn5DjRC258mX3YZV4/R9H6RHLV6AGW
B4EYaKJ48AvkHwWSNWbTEVqdTRMvXOuK3d1rKEwqrppcN7C83WBgZ8x3jQuIVZ+cQ5Py/2RkElh8
2dTCOTJYKSSiyKU5WMATTu8GwfNMP6BMhYAwPOZgOpPiSeYCKo61He8zqGkCkE/wNSAgwNSKSRWC
/ZcaUcUsIydyQnaj75/wAiLt+PWoUQARSypjfa05O8uaHW0Ko+33FFYIgAQmXFohiv17l42S+Q39
JRd9V0CMP2em0xlZgGPcwOptypOyBb+A/0Iijkp5GmE6JCQDv1ariyN4ejOcFJtZaapOxYwuhpYy
Lb5QFw3FkGPJOYZugflIQt/gnELJlJcUdzMaOW4efJZ5lc0g8dOUbbMesxyk9T3HnCUuuY7FsK3t
Z4pttYCf7chnVBphKi1un6cJ35YeAudDVxB1EKbUOuFHS/jrS/6y4pxPVRA64GbaG73wT3GJv7TW
6lCrzqQhoF41u9a3VUutvJiE3WyOjxsOnjJ2MTIrIJve0JYPO1slQKpt4HXgNih3sZct9QSjhSV3
x8xlvgk3mQECGTLIzC8XOZMCS+WrS6/YS9DbzXxmLL7FOdG0mG/6plIPW1NFzuYaL3VT8gC/wdek
kCihvnxXQPnz4I2JcT7lXJGRenUBZn9+kk5ZsOqI+iEG2+CQImmKfZY68GNyVLyS8HIdVfdU6liX
x4r0LJN5dTkqGh/ipzhOig6VAD6l1VZjg+lhm1zU0wvbuHwRK1PJaMiqAlcJ+DaE1JtZaf7TYIIc
PaMszn9BXMBgW0FghsP3hoDf7CVGmOmaBuxVxv+qXdJR8EcFm1w7zcmdrk9oOKZVaQDMJemJvuKn
7rQslvwhukMr426sO5GzoJA3Js7dBHlk7zuHVFzkf4eagfQSgU+UohYGw5MFQmqXhmrDKlT6HnMQ
7910VWBeUymIn4kbW7YuYKOF1Up2N5/NAFLHyWme2r4o7kuPGzbvK4qBhvX1XNNTaFCGQD8J07ZG
tjbzPcBS8dRwMTq0t+dcczaKBtfabg+VpEecYD/lbubVcYtu3H3oCRuL5lR0f3o3FWMcot9YXhFB
cplEhj6+m+AbWxH/+9yl7mqmvMj2yfGH0Wo12wW8ws4R6UZwjQrLwvlaYaJy6DYkM2mIZ7n5K0mG
EuOm9jisFX0TVGDWKS4Wo5zE+H5L5PxvxxvjXlznr+MFC2gqjrtBxYe+2TmLX8heBYPPgm46Gcni
QFoZf6UtgYv9yDi+Zl48Gx9JgKyhvoyPIHwpxwMA7j5St0crAYIyZT/dFRuTRe3YOEM6X/rADoww
d9ugTiedonkO5k7xCoLADPFNlqdff55Wr42WN+V1+PDkhWGCz/j5DK1NEKoFuFvplMjSpDCrQD0o
ZHde+QjZ7cx4gzFcfIJjac7U099rEj8E5SfKXRLQDs6Hc+IPwR1pzavTYc5EgridwMOkTpcd0OWh
YrapjIl0uJ2IoV82rBxVw8D09QYGh7sPqhdtoNDQVgMrgIbuOKB+/rBSMhfh8j6e2Zt+KRpeWzz2
K4SiwsTaeGynzyR9yDAwkxNj7UU4Bey2fDLEeOt6OqunbCM0F4g9wUjA/89SWELbUyJyTiVP1sCQ
hBnkkS7oGPB54x3RFeT9AljOJ48dUg+YXQILYtdtGwk8pkZ2TCoYLozoTEJjDHaOQ+zKzV989LuS
b+FLS90Ra8kFBKFqrYOBncU9+bVCL8923GtzbohGK7di2OBNiqQ3CYq+p84wVUnNotywFMY1y7as
rXiyJks3T41CnrB+VE3aLhVG+AVJr4Qpqxc4//WSN/Swvl1GHuHqj99ELSzuEh8+m54qie1BIG/Z
6cAGyfTs7CSuCz/18Yn0rKHH7zizJRz0G9pCjhqa0jZ8daqbt+yU2z5t0w8yFS9SwE6aCQNfNh2/
mH/UkpKjVUpG9SbFHXMB5sUZNkguO/lLl1biSA85ayNH2Uz6nXWzAXf/9galsj0NokeMxdDjByV5
MVfyghUUZbUxIRTAzBEZIdB1zE8LJHheSsbhyX1zMvYDjmss2j5KSevkBfd3ke+BatHkhig0wYSe
pOrpUZAcQFQcAZRpW+YdetR/TmTdGKkBTGRwIIH0t73/1GT4YEEXZe1Yid2fon+/qc7BX8cVK/7f
MLfprp4p1InHwMkVnZJQG4bI0ovIESTNQ4rzaoL9cSFH+eS4mQm0C+Ewt0KdYExZXY3/NQT9CIpy
C+OY5/ynN1ddAI3kcxeU3k0+kPU/zFKI4qm4PlBaadqXv0AqG5CFfx3RxuIeNzNAr61FaaU/jzMx
SS/yLzznoULZ4qDBsaD0gEP1yD9qHK77qcowfEHLOD+VhbdT4rjIQTq6r1ck/YrQUnCpe5698ruy
2TzCcKmb1qmQl91VbfGKJ0XqdWbtoQcIXt4+ty8OE7NWHv9wrJc9Mmpd0RKIYsKnWHXag5HToJ4Q
XbSBUzdNlNgcmwDMv6eENLr1Lur7rT7GEHE2UINgJiRUoTSUnyMSn+wxNpYthFKbEf8wzSevXEsd
/1oOaBw1DZqyVRK5AXOUUIz00pBhbTDqvGCTGmcMZ9ZhdqtFNsuxeXZ76r6tyzRLikAperaVTZcu
lIvn4Pzkye09muabIiM0GTwUrFUFARAFWpVc611lsxZTaYVsQ/kdPyGL3kjYpDaqWU4caw3o+d6K
zsdhjVKg0fDV0fgFs3xZ3nb1/4TSLYOTGySvR0DUZmjxstZ2XtD3S5jPStAAHGPSJPUr31qQ0Bua
F9Nrbh/jPJ+S+qG0/jnUDtADaroK0gWtbedPauZSF7VjD2IsVbqB8LwSKxEuQGVjEZNWwB2PZJxY
jbK/fQaXbp1x4l/kl9J7QPAIO0KiO+eFn02f2kaE23NKLorlW1EOyK6xtp9UpOtBBck2P82jZUyi
UeYRPkEb9J5BL7PjFwpnC6x86e4DDp9qx1FIRVmmGYMzXFu0q1RGg9B6cz6ZI5e1CuatkvxtIs3l
+iMTSDXqzc3yV7CPilUCz9gXRoP3PH4nzIl/+rtIWk+LEjPHTlby2JgjkvhIkcuaiXKEXvkOdPrX
WgKcbAw5w0/URCi86f+k+oECoWFVu0oHnn4NaO6WSSJL5Ij3Hwh/tU/7C912RD4T0Ez1KxHg1paO
J/SInn8qmGVZ/LGO69EwEa0ZsYMEzO8NfKb5vL6hEbMwmqy/0ddyDoYzr9F5NV4gwlMOIjPVMjiI
uAvlc072kFKH4p24dD625yf/wbJgfH4EqeNQ76R3J+A9MBdZYOQWwjIZ4koMK8gA3osqeQysr3nY
R3YVKTmEkSaJ9IuCUKtlmCgSOHgyybLfrkEZbSdvttKYQ3YPWgorauS+vWs4U3MGUQ4wL4z5K9hd
4062gp4AYTjuy8Iamhz67KarJMC5ROhP4ViZGBDx24ivbCIoibpDzNufMBt/7dqfq9E7WyLns02U
ds0fwf2HRkaBRyla9q3TrGPhaiYp9yFy8jhN2pLmcE0xuZpgZIQajLx+qzPO1at9l8uC5LEj/qSB
67Nkxk1n+6UdtMoF/cbMJU/LKY556pEJYS/BHUwlU7XAp6rnUEHzLPbhRJ8FAhY9gjQWRTIu1equ
5uM6ILkP6lPvTtrX8YG7Uxacdf5EFmYs7fEntiVyR35X0OY7zTpwH7jgZjz82gtq0tLlN5lacmUp
C28jyjZPyj0IEPeVmLdyzn+dIr3Gjs+IR9tbr4fZwnHoFG0I2yAD2p4YAuAp2E2E/2jvLCC6UAUP
y1zdiu3Flv3M3r1N9mwEObogzCBsb8QSA/GMSCPEO087PlpI6xlvPOlxw5muGLxq7GhA24h3VW3d
XaWIXrs57boui57kLEt/vORGGvfdiXNk1olhP8ygauYJtsRyOP6uXFhaPsteCH1Jbc7Pfs5WfWAz
SAWI9zrDKW+9ftdk3whqOgA7K37dPodLWFU9ph97u4xm9dRVsY+c9ZHPRqcVvdEfwrP+Y4hbdAB8
dyiYju2BmzDNx6T9zukWqU9sr7SyI479UCOO5bc52IMu3/tcRPcd0tRYZDNOeMTnR5sl/9d6lSlL
8p2dnPRXHHLd8GcSwyT0JPrm9yk9zC9r7RtSMj/Amve0p9RrD0L5L6LD6CXMowpq8ikeMoy2uINf
6gxQi3Tb9TTmxFHMQsGwWs8bCFU754338Sy3AxjGbCAG4QqH3P3W6T73KzYjiuBnLajSNwllN94K
0tN4Z3NO0ok1pkoSQ0Grup6nPJ1PlqhC1y/fWuvxX9eQvj28jylZKLs7rhsOuSpp3E4R9tSzW/l7
cEBsXxhXsq8V7P1fgEIPS5VZHzvk3WbLKYw8Sr9FrX1Uv+Q/AqleStneQAfgEbmwlV5hFOh1H35x
/cC1H0iWZwSE2C2JyTVM/CKbqh3oLYd//dox3jDTleglt5PSGIL9cHkgbD0HCOx20xMO1AgUptXQ
GniG+IZa+/CBHiSYedA15IV84w/RYiCltlkcWGTEcxiyreW6oOQtmBIaTTPYuA8uzMg62F2IsNnd
MQq6Wqw3UABgfJD/XGBSZq28B2wjxNK5ewgFMKLYdkFK5pCod5EjZZBifgG4og6V6yc0QICLyI2S
mLBLBMyx1eg2jOxZVG5TBXXNdOMxSZiPLQumGyCvggQneOvepbcHA4ZE2r4qX4vlvgDBZBfjWCWc
1lNqFzMLO3N/79YRxgGOiVyS0rFOJlLsMxs6FcPB8T9GgN7Ho2IXEwL3JkpD91yKzJ8JfRnWpbYj
rwcQcBW6Ca5liHZWoD74sgScGboQYCATVbbZgPK5swPVI+H+3zc9r0yHLGaFoZCoLaMPJSdp5SxV
KoyusMuU+00Qv/4pK56CIG4WfiTsZqNTF3zKilARHAS7xiVlz/42iivt4RwoRtv2tNJeeNtkYRlz
Pv+xxUHb+OhvhxZggl7N/3P3INPRrppYDjKzKdJ9Ld1P2gYbyFKEV9XaWQ6gCwshKRBL6fIztCnB
vpllIy3cz9F7a+PZJZtoXni5cw9Zf7vN56nJPfxHHj4BH9b5em49D/TVU82vvgDIOMWogLwxb2FJ
YSxDjO46k/Z3Z8N580eciX4eybNBuJwP5orLzUu/dFvnZ9neAPLv3CMFBAbsUtc2sja6FqGmLMtX
TXWx6S+jbrAwhxXQpsRTeyE8kHHoF/O2yDEthXDcD5dBPTDj7BcGtmMAEDwt2d3uSVMqg+IQoZ30
AtuffER9HJL01bbsLKAGTrEms5QTfaUTnAt5ttKaMRx6h93y+iKDdEtBpVWDoeWESOOouy03kogH
Pmg/olntXYkSoALoxu4V4lEAz1+5QpIGzgo3sDu0JF1GFf5JOVlaXD05r5pixsHh7cZGPA+tPtar
OV5Hwxngndo1yzSTJ9JKXpsJLfsUcyNGi4w4GiG2AlWZ4mAEo6FGI8vS29oZWaV0s9FS6bYLTD4O
jUcl0F/Z28O78uPHtWSmPR1e53Q53NhFKq1S1zdEpdJzCi4Ffj98j4zjGd++Vc54Pqry89DxQlkS
T+ETYSCYnsrdkpdSwvqqoR1OBEZ/Ca+KEUac6TXUmkgeIhSgId2afkQeIMVJWKgFeaaNgnzUrtL1
Q2ps8GfqopZjVGfeK0HdM8r4GAVSPdb//8SY/lMThwc5CmB/ox5s96RSOo3fnIxQetdRhzkrAxVb
Fp9ZYp5rfvtQMBHmmBQo0lQ8WAYIN2pesUbfLF9ywI4wDgWflPlm2KeovPkqXEWSlVJhSEl0ry5X
YzJS4CjEnCLLyJ7ArZE2KmHB6CXlTutJuj7TK6K8h408baYaIugyOWkID6+kNyszeS3hHkl9g2HZ
ekxQrm6J7WPUQzXcrMm9R+ymX/oyHIZZtpPYv95SLbzZkf2U+P3jZ5Tivkh6+XaUvkK6PXA9SMqy
eGBJI0dUgc1j0eZKb5mXwt2zNuCcu9VVMgnqlcgdxx8oP69I8HqSZQA9yaakZ5X+Jheaj8UpZOjV
gQMeHpqURHZ4vP+BWQhq0E6DqRJycghNpNVe6FI/5YmQd8/9G2mos+Mlyd68HCNbW0MJRL0yyd85
MKYYZjgLCe8iFHMIUYiNUq5tMY4EjjAoJm81rOR61sbW+NQhcrrBWSyAoHiC2bHo4MET6LsnnkdK
S7mWKhXwTWqIWG8WjOBK1Fv5jGo2zZEHSOz7M7TaFuKLEoPfOmh8oLCIN/yaGAU/+ypagF2bWIQH
ccEjTlOpYtrxPamL9FXr2YIeuapbnLDX7aTNHiueKqsb/Df7dOmuOs3DJyDEO4F0t9crOwhmSmB6
YyHONSGFy+fRRVHF/5GddJvhnJu+M35YI1RbS1I9IdTYuRVQzutwOL6TxbH9qfnGUcO7vLo2CMVp
MM1s/5mSFFmBLT7/9oqIsycUcXG7MmUBeN2omh6pQ+eObi1eh3R3/G+5M/m+fBdT6ZuuadW2LZcR
Fiab9Kz8h3JA/U+7LNP7IXmD4AXcbAhIYL3gZ6+O4TWjiJt/opvElHf7+5oHR+M34CcchGqPtlOv
BNQcVt4Z2sE+L03PRKeeoFAx1n5+7um4s7/415ZsbsW0Gnlipmcoh1LPChu7IHuQ5qUspBU+uL9e
rMlvZdiDiCNNT0p7wPibyPGzup09+RVLuP8ZChE6eVIGId31ZrF3V/3pSuw71OFPeNibkP/BWwkO
eO1Lyx5NML7nmrm8YzhFRTkD1S1Xv9tjQ6lwxmxpczRmxg+DJDX+lbmarvb0zqE4iuz2ZHTyBDYY
FBUjJkR1mFhTJIK3/6oF5xmQomokr8IblNw+B/XIRiLabEKB9g3vRMnokdRfx43KQcypmDWb+AnD
+V+lOHmplVBgm8JCUbm155F+mtYVg56Fp8PbMvILD370N6NMw0RxNcWXMfDy8j1TYhQQ3Bc5GkVV
nkMQJefK1io79L+1klBIPs5754t+A94XnmCW5HCuv5Ojhs+tIvv6Bw0JyVYz7EDQHM34KS8Y0buZ
G0brLsTaeQnLKsMwQEUUTue1QuoZzPgxh0ECPBT23VOFd0VF2U3rsqEW2XBmhJHrRiXN354foumc
UV8bYyxnooCdmOKoFX4O9+Z8NLBAIAdQ9djLufgQ5tZG2Y7NUGx/oYYbeOq7PGjH828ibH57LR9b
QrRRkcy4iqrRBU2gLNrorzN9ppbQoHJIK/D+UyYOZSkDMTBnI6GkT5uDATPKY3VRFvKS/k0e3ewt
BnFwdsH6/o4kvA44+xsqu/b1QPRCC/EeepWc/cMo5vPrZ3qtZiZFW50lNJQm/lAgaUw+g0pnrDLM
2x3ww1qHwLf4djHS55YK9o3mUeBZWlEgR54jK6jok0OQOf5oXfMBaHZMoqD1+PJrPr2ds2o5BkQo
pX5a0lB1dKS6tgJny46eXMx5vrcnjXzQMOkBtQ/8df1GQIixPdGTfrZAn92TwoInZ3c2o9soe5fz
cCczWyLakTQJCWaREz3cjeMiuF+SkCHhFXF/pk6xkKlWI4NrXqS48nZTbCa5NYZbkfdvs2ORSUok
72Vfy8ppHwS4Aex8y8aupUaLC23jhakOZW9zQGHlDVsr6ImiDyB6Z2+RxN9gZAK3FfCSdFmGFwrw
4bopog2VTXU55z5LLFPnKx7HD+b3rrNxqbe+ZqwQ0mAJf52UpU6ZImDo9Sb6kMKUvmxxXpUYJlcE
cyfvKjS6Z4fG3KGSIUePIeycCrLXngAc8ZIK6MkEh5nEzm3m609og1/8A/Uhr0Muihma5DraFLPj
QW92g93YNmG3SoufC55jRorWFIk4+MqkKgLLSAJ93bmOIzWSeVEoCSfILMnm4Sth9TKR7xEzkjrH
0+FyEwLECMlyAGnNtDvpkElfqtOooUL4KNFtB2rtfSEQctu7qHjkz6DYwaQksqi3y/Bc23yWTsGL
Pxnidu7wuuhaZ6twsYXM2qFsy8hK3txIbT595hMHvrxTAWRIweh/0WOGJhI3MUWInVOgxG1zdoes
moZhsq75LLuk9oGAoQgJyKJBZxsPtn6YoFUKlU558X7y1ReJvgcXoMF9+AHjFxzAUkGNNaEc0Ml0
i4AWJrRWRWrWX8f3XlScgT1gBjY2iezI7n2hD0YNQ0zU8XOVR0ZhGf05gk76EBIfT/BCYurQ/BDb
SHWPUaYyTxnT2Ti+7J9jHm9OKilfzMyutkwaX5vJYCGCwAh/AF4VDSK+NbakBvopYvilSmLTrLYN
Q2Pslyyn2I1ZVBDdZerM87JVjLb02OXSVKTH/FQXrCXfKYOoXR6TYoQ/ZCAsmeVxCLpOQIcAdNm4
Oo3dIGpr7hFwyF/IN+cIsAMf9kZDwWOLKH9O+wLU0kYmVYP0LHztiupo/LumDEngKTgc6di3w7+G
l1/h/skMih/k3xtax49WtKNy/02rhbjVuVY0FPmNIgqlRRvqzVMMignJvdUswkLsfLGyi7eYvTF7
Fx36gfbo9JO7Y9QewQi6ZBaK8e72w0VPUM3R/sGzw7tkK7bCS1sb01uz+Rmx8AI8Kg2s3jwpObCe
Paq16tFgzuw/rmjEDv0URlVwjuIXmmg+EFPWQUXF2CZn5wUKw2JkIgn2ggDZabIXFcJ9XOeQkvI7
IUVeZ3Jnj2cae/MRYja437mEW12Ea44i4aKoRNyTXvNNmgDK7oOx7SNECl0ujLgqrMZnh516omA3
NJHksS5t212ay5MCzcjElL9buJ1zuyqbkQghsuVpeGmfdJmPgLhoEJhP4/Oyivn6fCZUCFnF0wgm
uho2UeupMPVzPf2d9tycxu7MeQCNoCV2ICrOuAzg9sNMKWAGpMdQnjITDOqo6ElM8FUGV2Z0tsRk
QSYT8Iuw/vO5oMKMm0Pwg/W2gZ6kWt8jw0d++MsCLfOuFFQtfx65cWlSj7kaxnzkYktTS1Oi1QVy
pPsavHznFcyr1V22ULfqe0PUXPTm/8+kCAhP/XewFzjr4D0teW46KnOEbsXZ6O4SwPmMUcomuEtP
ShMkSmPmDUBGBRRlZm0Fo/CUie5PAN6kkQNaViLlcuav2xXQ3VeIKmNSwYoxZ2U9165IdnbkeS3Z
Tz41wz61S0Vq3sSpjNpI7+0Gzp7BrAQEThHecg9ES6jlAImjf+XUwbjk6DnoMscU3BlifWUYtNSB
ACfp23y/aya+/ZJe8sH4J2fR+wNrgvHkcIKYax5ire8AcMfiBuhNLmtxJ13SzctCT6WO/oSslLva
8OLtBSXo9aO39IP5LMZF5QtV5bDjVmgnLxmcf3EOMFWN+2ikLsdjwCoQ+im96XT/yIP/SH919o0T
+bsAk9VCc0qHWNemffeQEnT6ToKFZv8pRshhSz81BBLB+ek1mKbzzOCqbtqveNc28YRdFSTeyG1y
we7aGEPP/26XSAcvtfLxnsqtodW4NIOGq/STg7dT1iLUqdwPbqsPSfXVIhiNSnphb5pK+MvUxQ3H
8a1yC4Rqa/p2sTHw1hMG1MoBRvibq+wr7SiRW44JyEnac32QkYdLbmmE+dCaV8u17UmwSoGpO8Jb
seSUW3Kk1REjkGjTjhOgt4Wotm/AZiICYxwZTOZAhW5zM8P0fEZ4LRktjXx6OqE5cqXTlIdQPWip
A/opN1MbUeQ3jSY+rQBb+FgsXOHhKndk7ZikvpDXQ9kgcUfgI1FfZVaxuKClDmnvWAccBU9/m+Ir
KtJz3cAXa0UtosnlbYITN0uvsbVWqsFbM0/6r6yJTN4HwWkPkGNJhA8Saam491/P6HRjMqttMfm0
KCo1NhroU7fwsuS/jqYTMI0fwvzcNBOUovOl5RFPAvatX3A1ebypoF+ZaJQKWkBIYuEEbMARrpsY
+OgbkfDRRFUW72aU3EpFluF2feK0sZrdfS7Jr0oti9dv4rYVycXZYW5LJhh23ludkQLmjlwZEBSv
tD115ONUnhcMIKtezHArN8rPaSW0SnpLJ7PQozaPS7yUsuMIuUJN2J73Fuy46ahqocp8m05NnEyc
hvWA/exxPCZunkXO05ohN5+kw8S20G3R0kfMMtpjnUFwOi8WYzJIsUjMg/GkLmfO88zbO5A3+UYM
/SxA1WBRuAJyPmYyz3qXnMJSevA+D9JMnmpQ+WXIVwLcGGs+JrxYO57qbPG9CwXgJV2xr6bPLMgu
pcsWs0TnfBgDe7RZMjiiiRuwlIhdbVrgU2RaISLGiiINzuFV6NvPFzwOzt+tR5A450FkgWCSGy7K
c7cgB1v1Q1fdV41jtpo1UziW7TV73c/ZZCTrh/rSYjczVqqy5QGnqnBB8Ib8yqgiA/w6nAImasM7
TT5HmnY4XjUgq6ddiGukoWe33HWI4H28XjHL5qWVTr4T3SJnim6GSsNYJCsBADhGjatxzzIVY1Q8
TcW1/pAtuvlnxpLVwModLKQs8Bm9oOUtLuFo8BDUmEwDpLpGoKC4U+N5y97W1fqyETiZS4sjCkIv
3F/zhiT3dPrHkUL39bugQhZcbBZOEtheAgQ5IcSV1ycTYVBNXagRSevmf5EUV/hShrVTd5EIJj1G
ASj5waVeO8pJr/zO1vUbI4w47RYPr4Y49EEcpA6yX73yvv4gmWbBsaNCAMXu7AiSGyPApCbfpUfb
8JifueE5TGdaesJo/UBXO95x5Cnu2Aw6d701ic0Jcqym4IEb+s6xXMcW/we539MoqvnyXHWNFBCJ
IVbd7ZxB9cud4voHaawnDOSKkpuxnaI3h4fI1JfxlL6Wuk/xJn5zXmn/OC+3ToW5tk3rvuajIRok
ZjIBHkrStmGNWK87DqC1aL2lE/8JDj4oM/gpv2/UI9qzX6YCQueFuYJP2WK3GE/vJxMG9QYJ5hGt
YdRrhjGNoK7MizvBCPVmpZG97358BN/Lo6O5wMeClQo7mRNpQyvocF1qVCal4uaH4ny8ZOLvNw6X
8PRDIo87YpbCQ1VRo9JMXsIpvNj2s5R6FLFWs0UMyiMOOCabMrDLIcK4l4z/oftz98RBsuD/XnzO
FETmFdxKkVy9uGvtXFMZT4TH8/Wf9+bK5nVVU70SnmiPpHaMko45lwpjiswXM0GZo9FP7o+izeN4
9ebDhPzwaSEzmdXmwVq3qmCdZBqcYinHRZo6bsX0S42oPaWHDuFVHkTvurAwKpQCsfg7NhWYzmgY
PFwPKlxoN4rdoHV100sBACuUVWwBdPfIgfKJilp057IB4hZy0BhkbshBYz+hvZqCISh8fBWRJlwc
QJYpZowoyDOSeHsv7m7J0Tf3BTJPFqi5edAlYAQSL9xYrI0wSdYE4e8jEn/wlWqvzGzjkW05lEZu
ynvZ615r+bTaGspEnh2q8H75AC2BZ+2LN2/rMGZxqKL9m3EruC4TZIfP34HjkqteuoFBotoXbRnj
G8vfxMwBWG6GYdk99KioNwyroZ3K7Ju1EPB1QNPx7JqFaCrUYCYB2ny1ovQmKKBxtjDde1oXP1UI
M+EOoKSUyK75PDU1nWK/94NKPIlRgxfFTYg4yIcHe3KR21xoFp3CAR6OrAgVAOEIBAS+kA7pIPhy
B2LjVUW+VPL/Tx5CJkBZ1kj8k4noTSkT8fu6PEWvZnskI/VrpE2sxWF8dQPcJxz1A3xDgIfdS6eF
H4HECqVaz+hCd7ZJSiKT9TkfaEqEGbKKZibGsLwRrT9kRgwPB7q+rGkXOyNRhqQc6RY0iW1sbocX
CXTMUY4A6p5SeHVHWTDyN1EZPsZrOpKtbAXgqJeoDt0ij2drWVluvh5khKy8AU0Ck1NRA+RxC/sO
HJl66rYdDU+b1ukYNUdV0Q34GOk7v49wNF5qqWqvgcCR7w5EUK3jKYpXQY3OIt1DXNUrdazc6eqY
MewTW8Ccpgq1VEwN8sYZe9rs4Vg/uqRdFCVmYzaMLMGq24RTDLcpVe/PtHOGpZJJxabyOpRc12Yq
s2EK9eJ5lt1+NTqd1xuOGPGXYksseFZ93N1eUrIEsLy2yWBk+yKjm951MteGBeIL68wrBcNLjdqt
K4z29buHTmYv8efXYIhL72eRKs2tKCpQIl9jA5YsVvuMCwz1h8vybo0a9qB0Wrk7Rx2UA/Pdg+KY
+w6QhDUWyK95Cz8HqGHXfDsvfQUdkfI2le1hei8FWQYsgU1/nFt+LBOCX9Q8MNnp8O4573hqp9r5
M8adMx2qpV0MLX+12pA8PDrK++w9rWdWr+26ATMCaBaS6MU/cwSKSzLOccFRKlQoHZzkRB7A6Bq3
/PKbGWMR/ITfZJEIcv1Szb1hNdyktnMZVkE1Ldtdcd+gcf8YDtan5DKH4jZii1Mx2lDx54Q/fd0P
gMQ7yik4jzslnZZdo4+GWfWJY5KkuYYZBqHnhMnD+FdtQo3eNDUFz/JMMH4+GgGCbntE4HoeipCp
iSC+3h2bdB7UVKn1z7IXVCiPW3PgSqG6PeEcYf3PyRpKsljGDvRx7w5wF4jP9psJKS+KW+uMoD3P
MGU+zBl6rae1zJRSRdhjGw+E4KS79Gzd5g2fMN7icH057duSa3qZCBamjF1PD/hWYlC9bme6nPnd
MccXXItQejWcdrl5j9xGEP7sLJ9tYUBlbjVYzmYv9t9Wz6JQRmVl/d42jEyfGVrCmWH0PygwOJfn
EpspZt0WY6a/E0TY116qKwqwKjpuRJAygm5hj8phvdH46o+inFH+9y6URWmqMFpHLG5PpSn4yAaW
MEDJhWAth9pRwN+9dgiJtg2/rdqnuJ9Pz8+57vs8C0Ls9q0SeTadDlJqfTDsQTjxVaRacyLfnssC
dxGK4Um4PoaSGyLd2fRtULVU6oMd5EsmZbR4L9v0uuK3bwYh5sm50dbODcIWN4ZZx95xCfW8GrFC
P1/u+d0YtjRcKf0Vm1iSfHDOJ2Ft/ejFR9xST+M165xW99PAq+/QL2RnOjCr/4m/Pjf9lIZPR0Jd
G27kuHzPjdV/fj8dW5NIL0D7Ax/HKKt5WmuicVC+6J1uGpz141E1RnWfxsj2eNcW9J+cHs+BddH7
zSaQkGO1EXIH2lTgY+LXsEOa7G0DyuaXSD75PA4zlEtr2I2agb4BpQhR/hVIJ8XkIUOBM9K/gLIL
yRp3HcHPRu5ltjfQEZvZ3xkKV7VXIZ4k3j4XqrRXD9zmUWJeh6VyhV0DUwxjYDtlxnxAxtsPgsyo
sPTBxOz77Mt5t+tXwRlD0iTnqZD91gWRmXfz//SsdB5IZqE87X1RXp9p/3fvl+ArHzihJzb8f+vl
XXNWJiiRob6gzaFQlbCLUdp+gFk1OVJ9oUx0pix1HFiiYv+oMd1aNcPMTcBIx1otkSC6XqEZurij
Kr73eO/U+HgPVWSPd7gZNfdnRMCDVJWC0DiBDdPXjyMZ8gItXx99s8qZakrPn+NKSu7huB9dgZmE
Cay33aRadp0B8yuRdCU7pV9T7TpwnU+bKRp1AiwdKApVpeqgADnYxQy2Oo7czb6pOs796dtefJD6
6Ir6ztX2SbFpaafuwavon6ZKmTP74NApjpLE0fmSdTZYI8bQctQt4b5u/b+OKMLXsOhtu/6MEjXv
1ZPmQ/lz3mRsadwiNcuS1f2OxIx/J+Ziv0uTsftg3dbftk6Mz/wA5/iUqEqYjNOS2BaxVwsA4IqJ
eCNo8MlL0UnYoEJz16DzVtmTjeEifZppBbhPmCtSC3b2HX7R4elm/5hNZSgPQui2c7lVOD0OfRyt
09t/nXRpy3Q6gx2okjffBTfbfEsotk4sgPTrYLdUhE3ScL36XLIvFXAZz78lO+ThzkHC0uKfWexO
B6h9X8zRGT8MW7cOc8Me4rSbqBoR2gHIWIkNMO79oytJroRv4duNhh++OmaR71MjyHeGpL/OpCOQ
HNYmQF52YEsLJH97ypxNDBTUextvpgrzwblFjXGuZx+dGgaZioj2r3XvmBCQJ2j3ErhKY2e+mGO6
ZQtOJxxRvzR5DNpxSFXxVYhRhsq+Z6i7b66jXiXK4URv8KbpmMSOt1/0qOFj3C+XjbyO+/hEmLjC
uGi31TbzyscDA9vuUXf4G284GZXSQj8NJXbMoM42m91Ut/x98R8ojoRt+TcF1YwNwblMKLzrJLhv
z2ggqgyXu0S6gy7iyaAEf9tmtAN5TKedXxxVByPXZ8xY+eiCSZOgUMs2pCtwL4NysllnxAFkEYZO
V+L/sehFvFdO5PW+gjsFjWj+C1hf/KL0zLPwYdT9vAEPrezxMWtgvYrVhRiuWF40LdoxqYiQd2EK
vignaS/5gD36sRwph1SUaUrMXMj+4nsLRFYRKSoZV0Xf7awHcBaU6Xy5qbrUjVglkMp4pOH5jdGs
eRMj9ZssyZvXkDDZvAt9U+MuxtCBJensSsjg8g6z42o5DQKJi2QU4vyjR0CY+IOiOTLSmRGgxxqP
2DC+IcVREMhlVfH2nVZ0CYxN1UaUmsv5+uPbTfJorkhiHuK5vamYXusQd6/QLmSvdd5SzE7oxm4u
eM/5UtR/JA8+giYzyeb4rCYy5gQi0oEDGq9M0gKYJzFJYwKElDz9tD2ya5NIyQ2e8XLsJqQXuc6D
KQogS5WzVr+YlrKuSj5JuopiSgA/lDhZ+3/PE/I3BfR1SUDpeY3Ng2uZJgF/pfdZdlljNpmpmblK
lZpcF13HPC85tQb4FEKG/g/JRd7iVKAxrgB+rwSbnmiK/v5WWbNFpJl7mXn30oiTAKE871dEWMtj
Ue3A2HZRjfC7E8mva2QiquC3/+hfV/NJDts0QTkEhd+0aXiQlwTjyRM4fuzVsnUeBs8aZr0ajbI9
LoIeUOZUgb/1RUxmxyIwKPb/AdYwonyGL+KKn49/yf3ZMrXRFIJbjzh4WM5VadbR14x8TE+9T1cX
RGk2HxvBbmYwYTMwXOKnYx4ATVAgZGa7qNxEa0e+VEazApNTlwsf/94s/sQ4Eedp7t3X0cHS6VoV
1HevB5rF8E1QgY3x1AcTZfFjwW+35EBfyGwzqAVd3UR5oZOVIAS6iJT5JICm9Ffjw7s2SYnQPTXG
1XAnRvlAf45mxHuRzaPkEHt+FvFmoSmlPcI9r0q2sgne50aHYZrk3Zwi4aZefmDUCVw7Mf0p0dAL
qSf70SOsDlaLfptORZv8gq4vwYqOG8CILL9SBTx+bpYnWVd2DLeoElYXTNGj3hJ2EIpa9MSGawOZ
rGlnVR5ZTsTOZIvUFj0veOmCs1rb1ZOR1ybmTJRsONJ01bbaXpUOqiTa8cTUW2oA+m1WVzYsiTwg
w3eJ9B0CjddU2fnQEmZ+3A65CmR+3hHYRV6QMxN5aAhjfZzsrNgkAPc1Bnh7u3jbJrpQ0QzMQyW+
ggHSTJtMTHNKQuyhhSkd1l9lLwtQAXIJKh1hdza+NOBsSPftiRQlcksqPDJFnSuLk+hrTxZ4X576
lsUjrZ9GcEuExNuhrxVcbNdwWQbMHkLztAYD5yvASCRwID1puq2fWiCFy2bbbaCZ7cr0GOcjVuHI
vEZ7Fs/0SAXDRwvI1wTuGm//jG5REL5l4d+HKJxwbg7ph6QniL9NTSS2Zbz2ADhRLu1Dq7cBy9w6
ec6h47kZjUyjApqU9yFO3Q25YhMzFrjJq6KNiVjI147haZ41GigYhRxeMXbizndvr7unLnWmWwst
CcCjBlyXYmkVZk434sHdFEe6noR8jC5+Bg44I+UibVX6nJpgkBXXPgeQQWoVyREcTpm2asvaTBGA
BKrtTu5bWkBrfQcc5IXotSShEJS7fEL7Unhh0UI389WmzFQO5c++jGddlD2d5X7eNr1FGVvzIXU8
8owO3Kh3wkZoXhbjUMwTpghnVOorthSsbK9WIII4HKz47CeTOaqhJqZvqlkUt9qoGQKMTdis5khS
SLCMhjz8UGBUNmQZkCX0WfeLdkVXMhc7nwaXrtcPeO0eDCTySxBINJ28cq7+dQDJpjU6PHWM4NbW
yA+99v7lHAHvx8y0kso6NLg7OlWcAOADjOwlXHfp8WeEkQvvvA7ZPz7vFlWpyEIAk/hGtlJwQ+0w
9D7uJglWLWGU+dM0mNGHhAEgwCzFHCjU6vSY+aKbkusipvmxE2oHUKe1kB0AThPQnjYP+oz7fjJY
0owJnGVGg4MYZXcgCBTOT5huCgsCP3yU7KilZmPVabU6p4K+9Z2JDqwuW13Y8ygYC9nWrBd8OqWI
e7a/1bLw7yVzssEUavPwNg5a9i3zB/wbgVhgv0050Zmqqs+I3f1RI0SmYzRPO+Us/DrzQ6Rz3NbF
e6MvcWWD/4Z7JElkq4a1if/2NwE1vOKkDvInVpm1M2QuatVLnKMgInT0rR9wh/arxcMe4mmMm49Z
MjFK03tLtH/LTGrYKGFvqTlEMopQyGSyC4y7PrPTACosVLCvVII7a4MEhF6E+und/u5yAsyoyN7u
c1k6fXmcHp6RP6P0m2Zjhtq8ERf2NhB44UboH5PZCXBBphhj5JJbUBX2bKjFDUWNgdLtrjIpKbOo
iNVLkm92fuj0VOCJAbPe2UziSK+7XGEN5XAHT0Ynn0h5UsF8Z0KQJzLi1SNYwqm9sDZFLG1EcPzG
ad4unyQa7uiqzo+MDZEGKTXHEkBoWVuzYMkTUtmsL34KMdQ9HiYbuyKHujJEBzaOGEIQ3wNSYzu9
AQZf04K9zU17zWI5tbMDlgdQaS+gZfp1wlsyucVH18qQZIRSr2LRjAtsDdPQoz7kU8PJa3oDD4Bl
Fcw9f0xKwSzoIej3DlKjIPSKonUhSlYGsb392aHst2A/CZ285rsXwrBUFTryEd+kdMWKoPSKfLOF
x6AXVKv0vpri58pKWncL6b2qRcv3gL0nkX6b+hVUC3O2luechXac5N0ruGob8HPbVqUc9BYDHsV5
5PigsynQ5hmjbd5SW2TY7SIW2PQR+aTe7cj2P9NrQsT3wzlb8mbIWyB0h+dkuhKd79A5R0ETqUHA
/uEq0tQ0FfSpnYcCaaSBDp28X3c0rcq/jKeygKsbXZR7kUcEdpqfMjeV83+mWGmiBhSogIz296Kh
H4qGuXjb8nmFrsc3LeZieW3xj/oozcAQ9+Iq6u+Iah/S8avPo8ty7kb5xgHpwADk0xa7yjynv2JH
lAgJHFc7kfB4JjabiRZck73enltHS6EFBkQuvJ3wY/8Jq7zkP6ojz86RH/rxblJNLrJmq5LOrJ8h
0WfDCM5lyhU7GSyc/lYxLy7n0VS4WM8xNXaE8mvaZNqxkCi7REFS7WV9jaUSFVlnTVaZ4J/LCDAS
XC6ZH27LDpyVXFC8IWsKRMetGlairXSTv6r5eYFYHsUDUqvvfc4IVkVlhOjobnIhnrVOdir//4se
hbJiGDgq/ns4uhFFs4hqiCrEFqGxjALmtGD5TJMqd8QuEIFJTKnikgIyzjXOjnDjRWworqTh6VNo
J4BR6tar1VbQ0weftOY/v4FF+KtGuL1Z3d2XteWOPj5htwMf63mrubjiBiKKBaZF2Uu69TtfU83d
CdTARu0z8T8kWJj9Qi2ZJtEJ6RgYtvGtge/BrxvuaJHh4sZKi+gp2MrOm5VLAeyGtPD6c5WfHGY7
u3Xdk5eZUpZZQ1FS9QErl6w3BKFv1xl/pUW5BqARqje5S3y6j+t9wx66KlZFb3xq7FLHMNjye2zW
ZYQhY4t0dHnptRcLy5sBpOQ5ZzkzbtTBbmHec6qKaE12zDhj242ZRDNDdXlXyRZb+239TRAKc3hF
CE8Z2IBE2wYhyEUCJdck4SCzqBe8HefEwQRRIJJRFBm1qIEgXLs0q16MIU8wa2eo6GnUuHlrLytb
N2bzFfzKlH9D4HiLnx34kx/gnt/Ki30vqdH2blt3CLddyVKWjaaD1iha85FAl6dfsb1rRCP8Zz/R
dyhJqYfMtgkdlMSaikFqA+wzEveLtYMDupdgWPbTGEsHdHmn8Zsvs3lsKlCZqYM/6QNWn8DSrz1A
0kn+rTAQ+RflxazQt9WXlGWJzUzMw20BIjKwR5eFr/fhcSmmjVgGXglD9PfA1gmbAzs/IUUQSLmR
Yb+fehoZzFUl0lT2CmomSK3hYdLOYPqyjVa1zUYRET8MnxzIRmc1JVEo9QmOVew6AwVM517RCeU3
UtiOtUXF5PWT9fJEcQF1jPUMl81tLC8Kpf9ASwp/B3Yi7D7jTSC2X2MOfsiVtCN2KZ2J4Kvwc0FQ
xhnSpbLfF/+0cptoP6r5ZtJD8xNnhT0NGhQnSrDzpSR7mX8rw7P4/gx+R3RvcMgN8nqmlvylq2NE
EkUxOUUt/aUWle0k/prt3o7Zbu5ndUguV42WtrixXezCfoZNWRpWqluCg7hBTFDGnScPMa7f5Aq6
5ur3fTgLUvC2Xo/lPK/VhStId0zECUltp0bfdLDNnCzNwsCBsPsQA79nzHTZ5ioF8IbLMVlichE0
eSO6m0y+3RpwpTKny4rtE7uC9DDMdMQ19lURJtczJVnhDZcSbDWBfn4xOaImKm4yS1Fo6PehvS+S
7+RZJ6zZPa6/yd9fZRpO2f8XDnyINLQPVzwpikjsiOZoKG/B4iqTBICz+g4LsrddAr/++FJK4GN+
Phv4FfWSJVSKp3N9Q4tqmNVqGVJgCjfzCJsgOA/WvscGcC6v4Oz+NuhELbxG10AmLlNQbzAVE597
kciaHrt2cLUg7ixZmydF1s5ELsWnqILWHhPvBYlGOQRoGqL1jSuKeyQQSf10hJz9+BZ58HXuv2pe
/MXBtgk+EjzV0k8slxSygRtmx6VYvmXiiIrqRY1km2pVJu7dH69WSk/czyZvXg6LAgp/P50VWpPq
au4HYzu9kDibhM1UQZa9VKQe30ORgq1Xbn3tAMz5V+/xlMfrWLV/x0kf8dgt0VH8M704FcAR+xCV
t8MSEY+f8GkDkbGs/Tog6uh/mdxou6G/WaU2kEfPiZnZo+FY+Qkt6dftn5BRc4Ftyl0K8juKg7OS
MRqsDfEtRXasXM1rufIHTVM1B2F/cdc1m2dbKQbOE3aCFrTU97FJ0dOajltqsgm7KoXR/3q+1zNV
JvTy/hcn3gEeYAeSVGaeHno+dHv54qmJ+Wdvkxs4rDDgKNAKTzXjpVBe3an+kb0i9V4323qAzapH
FTA2u7pjkK7dXUZYOJqcqep4Z2tKcPaFzejMVp/kJPmTrBj3rJuZfYndoPaxrh4oJiNC1LxXR4J1
62GS2h1lPc9UuMYvw3KrmvlicRFtISTaplPpWVhuIYmbWAsgsctEijPT6Q4XpaUPrjxgE9qWUJkl
CZjL/Ymm9UlBEL5oFyv0OM5q62/hQ7wli/gQ/iRj+16xm+Vv0pq02I5lY50MxDoawxquNuvt2lum
h/qxNvKlK1kK/V/LvExVq8yphYmaDAs2ertJQCsO3ezusvQN74HYPMiEQJVAzb41NwsFGylh0ti9
jbFU1uMLFAjZfZju/viCqgIHVUQLaiN9p8Be2DATAtmPykO8NGiako5d5Xv1L38UlhldvQoo31r4
R2O71WNMgjpnolW/pI2oY4My8+N2/Bb1M136Ljvo2+tJxF0OQ4LIAhgQd/gVvlJRifq3QJpSU/N9
QxAKmVRvQutJQY97wxX6w/HvdnrfLYH9mT8RO/1CYCdym7NMyr/Y7MTRPX+3zBgHciFqjOQflB16
FlcsLps4+RlRldFO97enh4oNEAQdVII72ZOl1wRlXlgLtq9a+EJqbV5RCjC+zmJBKStN+hmQ9uaT
T2Jp5bivgF3757PmXWuNz7KVaznsxwiNqAZeb/bL0l68/7NjV040GbzagnyRvAmIs6N1kEYVLCun
Rri9nNKS6djkajC2rrzVAKD0e60O7VUKlfrMTKGZs7akY5cI90PBhuisrquKrfg8TLVsvm9S5MZK
3DWhFx2tHuDe3oeSTbDTYJVsiLBSwSUAH36vJULRbSZgUumY2hHiyG5/X/7fOFKYbLOtex0cX5aP
1KyyNEFxvMQV46iAONnLztXSGNWRGqfRElsn4Nl8WC+M/qgqcwanHY7RB0UWOLsClHdD7ganFFTR
z3Vm1OE4HdDo+qYKC5rrcz8AXecL609oK1BvM4Jp1TxaGVtBT4seeNMbzNurnj+w8hNnbqcYidVe
IWc4msZiij+4oeloyecDu164extz5/+P7HLvrhwt4vp9A8egt+KJgx/bdYzHWVhF0f3qotZXuHYW
lehKT++eTn0YZlQIaE1MNgPkit8hiX3eDjAlgZ0x0ZBb0F+veSJFKlrMry7xBKvTId7bpFSiqLiJ
/P+YxBpESYs/D6SHeDzOeaO/R+tXUm2BAwYr9wEzuJz1w39KG2tcB48qjpk2r70z0cgSwLykihXb
pQProvpD13WNT6WeKZwOZ3DVWppCMRiOYtCH9hPz0npMAQWniIfF314c+JTgz/YzCk5z37/MRM5I
kD3wZCc+OPoR4AAAtzMZd4KRUfoGcaSCcFnWtD4Suofm+VvXEd3+CqGA7c8cOwVua0JG/1sAP/Ql
VPo8pKdVnzdypn9UWjdZ70J4ePB1CuPLhW8cSUgmN6bxls3hqBXbu5UrDyDmGL5n650VuQzWlyVf
EA/3jdjAMx3EzMJzt+TSS2LriKNhG9uxRxOfqu2FU43AEWFyXUwGmNJgmEgicN76sm9/9LeQWMoz
N9zUsj2G/9yNwE7W9BwmJRp2QppeuGanVNIvulG1yknMvfsUmLmCMBMd394fqXBOFXNjOnkAxton
cQemt0wQLfDm/za9ucaDj4w2Pb5B5IUdWYR4Zai+jCBHsQi+xqumTpJpMJ2SMiC5wLrRzG+pzLXI
JB/18WrurA2fCeTleLxFmdoh7djHAfnTsYSlkly9osO0XW6CBm7qwjFlAfduOD3HEZyZ6HzqOjFO
xuqc0PuSfbB2K7BUHw7beDGxFLNz/kSS2eHCcf+XTOxHFx1rBu+vqQ80t1xs4HqNTqtYjGKWRd+I
C+/mkrSBEzjqf5Z17OqubjNiAtxHmO0x/mh5fk6zVzkKxRGCeiHikusCq8JAmX2sPtICGNpTYcO9
wjcuiF5h0t8Be4fGK3nA8b2r/Dz4e18AWCM4RTYUd2qPnP6JGF9ShN65tivkdlmzRpbQZurmRa9p
zBmCOXkw7XaUUybjZzK4ICb0w2IWB7m4JyBUuXzOlQRTYHV0ubVC4Jy6ehT3yKdTFYbk+SHQT3UE
SVj4eAvDx/hjCfjzXph6GSrOqzEWgLHwcvhEWTurzdLqntD3KVAqATGqEZKOKvZxaUvPVkno+UuY
McR3T9jBEuKQCvfk6pqwfEWniIDhhLcknGCfTcuEuNe+AjdUI7p3C3EVjmT76Z4FnIjsLCWlF7/c
leBnCucK9WuoG+bXbVj1G1TUZcP5fH9cok06svKkACL+vwK04jluNs5Gbu1syFR2w1TY1j/316sS
sbs5R2d9nsMcV+IUf+zIbpzK8ANuABYkOFSxX4EAw6zUMEWGcuJ3rX6UDsuYL92lCVrppQ9x3ous
KaJ/cbB2tGedDPoPzallh5O+nST1n/m+5aBAZYk93EUfbBdrtzT8Kb6kecFldwOJQlmkVKtjsR1+
LAiNYHoKuB8rG0+dTrwa7ylhQLIRSfhCAw6ISr0LUlpIKhoTUMetbPHWGjZ35RyXLxP+ODfpIb8p
GwZtDYaNuX74xoQ3/PNVxZcC0DIVBOSCXVKQ+1jamLAY5FxTZ7hAEFAN1LTZvam9nULH2LopaRVZ
ves0hSzcaZCV6Yb/ufUg9iywUBCqQ3fpagW6FseVQRlpt8aIejR6+mczo40bZLQG4gDlOoz4labW
NX+Udp9hnO7sKN/IytC0SsejmGNQPph4vzocFkUV74UB1jeTEp88ypRaXwkt8IhrE1U5AOzjMYRW
mjB5auQ5HfibImlAgddzs5XkTibzWsH23HwfJVjfNy4Us2R7Id+nAtTXGWT36F9rh2hsKkYYjiJK
L0FDQVu6+arxufDYsKQrzUevWUABMWneTcy8cssURQvVB3M4S7jhH8O5uoJDQ/e9nAj+W/WrCw8f
mzFbez9ofJMs7m4L0fcjqixhERt1PihwLMGfGEep9lIxEH5e8vSNzZwEVVkZ35aR/dA/JZ7lKQK9
7hMFXR5HyB/mrgVg8YhI3iFvKCjmHwK7XrL59yjqcM6ehJhQeTpnALOneltEqHGDecsu2YuwGXVY
UtzDzExBJOacifsi5bFdC2YnXwJwYLYiWbTZYljkD+NMHvwtblz8gfyJ7Pyahp69K+wIH67JKoe4
gyoa9dR00kzizWsZ6IQH/lyftlpIFxKRD3YMPYyzKbQOTRNfX+OxW2l2Wxm7i0DuuXoJOX6yMXBR
Y9jnlK96Rlzbjt27/9U7hFx5/grnlcg1+hloX8CGPLtefQamkxsqqk40HSDr1TuIDCCDmNrnD8KK
8qbgxQvDLEA/aIx4RC6cwa5GV+P+QzVIwgSqH3vFEU+yV5jXNI2tNN5Rh7AGkB2+8zx1xqZhXfdT
juHruiE10W0hfHhRg6djc9L7XG4rekp01Unhcp3+2P/mohS5+IYx0KNO
`pragma protect end_protected
