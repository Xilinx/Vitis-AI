`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRkcajQVnMQxKjPBaLZIaR7/J7zs
kEF1+54ixDuIyNX+QBxUIanAUk7iqIQDed2hUG0kfoXoL3vuow/GsZ8M3G4iHfWrH7YjpZpxAU7u
+39ASljNjmhxyj7sp43zFjND7KB7yDk1EnS5RQNQKgSwY3fvRC0feceeFHyy9eiKM0+E3KW82xi5
RDh2XoenLekPW3PgKxqpPoG+gCC21CBlAB1jv2k6OVsb0sJjvmBbm0nN4wPphhhkwJPqYyPtdgZc
CE4/fZZVZGZnsaxeuw2e5BkftS+Jcyvy7TwH2EXFCj3+LCZDd+5i/jZOKxpmhardcB6GTekMdZ7i
B7ESXKl5yXBMEiUrw1/krFisIqqoQwQyWbQHyK4mQW+7c1kKlPjP3I5seY1cqMXtBkD6oIJ1Hswg
yyonui4UkCxSK12sWrTP2NH44jyydQ9BDklzMNU7M3uy1MSVAE1jBy7+bYrAJhktusP0i5yY/xyj
h225O145vWQz5iZNA9o7doPEv42QqTbZIQg5E0vIgakhEOLS4+esQ63qi0aqS897Z+JuyezIdGoJ
vmGHW5eB/qoHd+TdqwJQVzHrl0F/d8mlhGER0yxHsTpMAJ9yZHq7jiVa6v5zOGVlxMjwU7tYC3Tu
IgPHJy/NgCnIbOpCGr3zFWFMJwOkOyHX69A6NtABkQirG+klHGVAP04TJE5Rdm221B3823+w4si0
B5A6n/sik+O9xHTxrd2okFGXvTSCqpazfGGI2PyfjCLhJ4vKrG3wZwhhC5x5rYHPR2dCeE7yDHYP
RhOAc4Kamnvay46GdxxsIVD2aO8yszJwTg+OmsZFKBm6z/N994XoXqMOFTu+cYLc9vo0Lw8NkT03
PRZiIQ0/DP5Gih5nQ7RrbKGGE4vvN88lWGkma7MD7U3r6lGvD4CuYeCQ/rXTL6REzCEl8CgxsCms
NPqrkZjwPGvcBDjFz+0hH2qQqQv6mMBkpyz7nFccKAoQ0AqGo84EiteI7RPQwhMTFAW/+6PqpaPW
ZBiH9xYzOjvpZj2jwpJz4RhAmd8rCdzdMd0b2nhMhT+G7imvBOi0/sFLmufBxPP/Wt3E7yJnUwOO
doNv5/cfgRzg6jlgBIyhFAJqFiZ54ASJRYKcqPQeLn4WP9sLP/rSRtYT704KYV5EfEpEwstd2OLO
Qs+hOZe5tRBgSgE7LtWLCmBXftNF2Obvad3NUOXHXQGUDKZzXFmrNonuJB5Ynezb59FEvcztmBgh
M0v6cpeqa9oZtaqpZgXz7ULNMG0QS79zgTN68DKQICjvBEJamb7iabtnJycl9Ef/ZTksqvO7LMV1
SAlp36pmFep0Jq0gOrxgw4Bul/VtAda0fTeWgyWVwUWrzbqBJsLTEkA0fUqA4V/Sd28/8kOh7bYe
AQgIpvdVHv/T+6NgTbc6hNN4cIx+H6mMWcDPS3/Ur3P44Nnl4Sx4EVKmfzwtu5QqAgv7yW3X4e2P
+qgXrQWrtcn6pr+h9DIOR3ZyQVYfe4NtgiSLQgghCjP0z4T7lCLGEbWwJ08Pod7PKYgsvIeU2Lbc
6wXkuQErViSuLyff7+7PuQxi9wXA5WV4FpjtZqbgDfiXwPaf4BS9XmmCcIrUjRF2ylxtSOLibMsi
jZDmngNCGn5/RMgbKZEWmjdLvDd9V/PTjbwsV6RbfsmTWF8Wt/0PkJ2t9BuDjuatcvDsCjmitJm9
n3m5o78YiIPDAMzqjA5dRkgS56dJRVEtKJWmoOlhHlFMRZm5MRuae4txkCBdlILCd3ckGRuBRgo9
V0hq0kIlrxxLseT3W40MsRW7SA3LGcW9TWTNhNnr0AGQxwAyGrjQYyYcOQPIrz5zP6XKudaCq+hv
wLAfUEyUfDDbFiFumYr9NLnP98Qsy1TBfSpOBxeXanurfp3/WXGyb21faTyl7lZnsfyTfGKYamg5
Yfnl9ipB6i4NB3RSqMxwr4W55GuSVWba/3DUtwdiRt+UB9Nwr7I+YIc3cZUyr6CDq515Op4pHGI1
vtwU1Ks62+NZ6jfmuIVZc5ZzWoCpY9bE4N+Dr9uHVvloGezZpwXRc2YGwOON+KSS4/Z/CqFRTxZ0
SQYI6Cmg5B5A84RwNkUC2ll6KmztJOUsxyf1V+lS2J7ilPz2m7F8qU8/HkPOJd8vAZTRSkgIXybh
TG3DUP2p6Rn3HQdW3rOdWCGmhKYUUHAGquwbNmawXdOTS076pvGKp4EJki2wjwZhiTb+LUMrxbFJ
Nt3S8RMCGuFlo3sUz/rSwNZROG9popw8fzFKmem7XCe3j16beLiIVE5AsDCXZDXgGRg+G85YIKyu
xqIqIslXvfACIbiVTiQsMhMlEOuIjRbnYuiKXd1tXtVhApbKBbSdkYCcrjbls7BG5gLDrKLtiKa1
XKJ8rsIyieWaArUPGR6JebiOa3WGNPH6rpMEiku+6923zBS2fDCi2xWETO6Lc74GmeVFMYpzj9BR
YquaVIOlkhKPVjjZzrXT0W7yJTj4BBqdc4UkxcF20S0f3IjPDcRHxCFiot2+9tIR1GCAtTPQaK0y
hRhLirWz3eADEvtU7vqwXxAlZGzjshRjRtgJjIh34xLUvHUL3Z/YKWFnLMt0aCmhXaiouylut/oF
PyKKdE2YNIOI8ZQXvuQckB4f2swUV6KTg0MAyX94MpEd8lh7wa8JKkDmNWeJYnTaxS3tRyDM1vbY
tlT5kLoOUtsaNomzxJmfTQsOZKpgYXU0ymGFpVKcTE2ent3rc+Ig4bOw1/u6CiegyxBJI8WQTkqd
RljWQgARZ0bnidpSMBIV7LQhRx7AOWuJbpoMX+uieFfMyHCk2xT+S7S/Mmp1znyMhm9borYlkb33
fKrfSkSup6FrGfUBlLta9zkzJbBiFquhyZNghB6z2mVSFwTWewVRM13+mv7c4Aocho2gvg9knpHG
EQxGnHOZZyzbGtOGsB1y21VARzXK55w1gZkPU5m68dOOzAFxgcth8H+8EzVhluL8hdb/1+KUnm8u
4aT5Oe934DFFynazfTTlrppXHlmhQZhK9H3CVBwwCviTAYvB8c/l102gdSBkoqo5tin8fyjq19MJ
Bzi3Xh1rHUbCTS4zX4xDsfmqczWZ9MygQA8YqXsEWfA8JJ7P6gDx6/n7k4xPd8khJxbN8dJ22Ot1
YdxuzCl3wMqMlW0OeDa6dhCMF+dtX8RYbE5z+8ON0A/Mmf4fzIpY4yKZTXt4ViYvzO1HGmbuHw1q
PqyXLIc3k85YhV0vQoM818jgWnrWWLSpN/bwmoNLQsOVNqI6O2/SmzOCuuCZhVfj5eSBKC9h8ZW8
BMvcTpiitEtPlJpH3zsopk6B7uZhIsIT09gSXAbx1PsT28MEDKwiRFGqd324gf+mvIuOLjxa+puc
RNzNXI6FjI2zS+La2oQufsJ1gUyIc92VUxljF7+WIce47TQbgv4Mzu9g6Q2XCJe4T89Tx4cKwlaG
jzGNdl+3NfGk9yrNRyBJbPVfNSBeW5It+8kmMx9Xdq1bbq1q8KuqeAvZTJ+MlXH0sUmRoOLLUl+6
Pajvk08a8b7IUuIj7avxYwzKSMvhb8T+6eP69CUjcUURVtQwcH05hfCvVAFh4RGTpofqyXDbFyOg
eqlnLWmfgfQriKsuuU/RNn6nDTvcR106EFYvuR0ImiaJGAcT/OezzQ/+B/+jxfW5iE0lD0jOyYd0
02TVMdUHL6bqQ9VJmxvPROt3SBZPZyYI6ARAbITaQ3Hd9Lp8Grd5SbZddxL0OVPNsbbgUhwf3Ng1
fMQOElqvykH1GXTTARUKqxy9RnFtuUkH9iWsawyuZkgJ7uspRQhobSG2G9Rm6Y99rkZaN3gKHQKl
SRIiYkVpx1i35+jBImFmz74g+wXe5XnKx2/4UFqBe06yqCxFgPJdeKyKPUIyS9DsPFQmBBJZz7k3
9gjYFSCTND8LJA8PwS29eckX+gDm3T/dCnx0yQC92JeskOKirES8ohnvXXC9AOmNUMMUqRjsq2rP
1AqrBcqT8Gk3V0sZnX+cyoiGENo5pa6j3sMSXOOrhzj/D4lRmLTr4ntc/z0BRJwXloMNKmV57dkJ
ZjaVdw6WI9X9YfX6jbuKA6CGYQwcKvmrV+/QNotdp9WQLomaST7Gune3/9FWyl8YiQmkZgADO76c
vfxO2V5zi9LfWcZSFsd1ZXVitWluTrszFaalWXYgX3gHcYwz5b2V4SsOZAWkfRbhrkqeGmLwH3lj
5QJLaT5RanyGeK5EFh85a790PcC54n3V1GI30jfAj1Nq0CXFNMdvyvAn3XyRD9DjgukDEXVwDC7b
X0Mn3TE252zBTTL2taTJ05Shy3V/6L4+IoxMsLFKS+Zzj+FMnDpwMQgLjk/qtLg/Tecxqk5wGSna
JtwkeJNLGxRDMC9h7po44S2hfPIAPSh+PQmkgHYDAVDGsjjJkFAsFrqdR1PCC3ALlChViYLg3vIB
myow3VTqKZr2kivmwJkC5yJTOuQiOqDaovvhwMhMAgNkKwXi9jlo6ljNe5h29nNhBTdPWYE4gEif
HtbFap2cv+I1XGGf6YhojjATdLa7ypYpsOiKLA3M5POQZTeB0X9fL4dmZvdJeAszm8qaihiDCWB4
cXTg9DvD1tkgoVPadzj64CrO/Ad7rA4TNMUcSuthJ1KybmbeUihBnI2BZjT9coPmO2FqweAwUALR
9py5D1lCaRoG1Y9tZL7WRPVur9CS/gI9n03OK2desIiTtQM/99tCdMSVIY6rcpHpxcJxucLrAAa7
/H4VgYVM6JudwNQwZobWla6haLz5PHdjokJ5LoaRddOYZKovKz6TqjCdgbxSY5Vg9fijQqW9eneH
GIT5k9EeDWliz5NxpIHy8fa/nb5LUqHKbvrtEle9Q2OKGuaXnzUgWoRssqrVoppXXaZAWk7WTjgn
BHbVh5yvBEvEqVOqm0ZAfW9rOuNnDR2WtQQuT0UkVj065oAy4/1LHNXLKNL+gvzQPBVM+3w1COOb
pDCdXlZ3fy/kL7MjDlQpsHtF1uIRH/P8tfoD8LGgwjmgOjreR9bq6Jgrnk4Zt9Ta82YyujAS5buE
Y/qIFbukdGoisst6Qq6cJVEoVsFKMTQGVWhwtPN9vOHnhsYPycaXZjWEPAmAtNTSPa5wDKzBQP85
aHR4dFcfRIUIUY6mNA/4j2e9gAlJI5Bv2ovb3pg9uRvVibOFFLPUc5rTYSKGhTSOUMggbtXtOsxR
K7m+RJ6Ov4BmmnsZqCAywsDR2WvK+XUJ4a3VftXJu6VxkW+rigtwRA2VDkqDnUqxTTNJEuj++oZn
s9pFNDC8erarGSJKOw9juvU7AiZuFnfqrmmDJ6DHUHPI3+WaKkeU0x+X9NtqueddfSQFsQzxz1jO
80l1/H45gIKbsJAJyS0mj1sBjdI0lSf6XAkmXRqNolkFOf/AJceoHdhh5uzlP11vb63Ty8zUMBUX
X+aSQgkLfeBjR43SQ6DONEUV4s2dQ8HjBqW0hdy2gz5qZBIcu0zz3kMtdQmBN/WIqX8+8no6MG+P
XOLNVfdfM7VQvwr8YUB8ou9tui/njBFHr6KKgLkPbz0XDWK01YI2uvaCKC0VEzAegY8qFQZztKzg
QRtMOqDtqV41BvNW4hhLj0yU4rOpBEH/l8eiFhx6l6zCazUT8UqREvXDOOg7lz1HM9MVNsFT4P92
Wl+LNLjr0eNBU5wLuJ+Q1p7YWqeECeqtwHeU2zjKWaVfE3ZmHlZVnU7bZylLx2Ymi8+DoLUIqOpF
EzZOtcGzJeQGSsoocblAPNF7E0MsheWdD0RvWEkH+r5lXP0TI4BSnOliAdDhSMjdI/FWKNFDc4qk
McC6EHmTTfYnxJV/9ho9rYMtIVU1bZY4DmW/vgmR97NlWYNcWUm8D5e/1OU0IzIwfgfAURwG9R6J
9HKhIVJ7ci9OgsOUqEEZB3kxRbytyX9sR9/GS1dwcHK7QzHRl7fdRphz+q84yRA3bClShogH1yxi
xjAlmL/Y9yhg0MScLa+GkMr1iXVOdKrMDUS7U+p4egwtOHBxbcXragc3tgD7RWhZNTxkSfEp2rPS
i8iawGv1eABs7fIBUYqqihJ0UUrt8+Lmv1v7JC7o00a5qKISOp5EvGw8D95e0aM0J6lSiCeHgnip
CODKUaR/OnPYxljJXmyObhz8hBlbDbIIR3DhUqVME+UmhcCbDKIP9bg/Vy3beir8Mh5EUXhTTwCs
JyovC2k+zNUYkN+cjPLIkDhQ9WglrSGW13rhTYIhN0c0tmK/qGW4FFL6xCSUyY45k4hCf5ubuHn+
oJVKoemLg3rYARugchcA6yrwN2yYI0EsbBO1SQuUZTyvaC8WzMU64KQ7q2+29rqTKkL8/9V2z5xE
j4rxq9r457fmDNyJs0tSgnI5Q4KRdCWZvr0xh8ulx98twhGiCSiQ6+ZvA5SLnRsxudlEZDxBcuYL
bEAZJRVaWca5BMUJV6uCDKC+13YT2i+6YR24JydmccWYJtebn4fGxdKX2RkV4gGikzXlI4MN70UQ
EGTOF2uyr9r4HUH/7k+hnTOsledWCpi3LTIeOTbsxbyD9KXJDvYWlEb7uf3S6HjcBTSf3xEWjcTW
7DZnFzhLbo5G+OsasqJjuLQpkJiTvTh2sLgnUkdepnViMNiLaWsrfDbLeTBYNysDQRhwPylXn3mQ
DlSHIgpZHOw8PljACGrrETvLlwk/81VoG+KO/k2NMNWJ7/b8DnM6jHZOzpE9TqBRC5BA+Sgg05yH
t6fGgU7gFRt/T5o4OmRoSojoekLYVpv/ADy/H/cYMDnaSPKrNIm2naKTrA71VQHyiTPsJl5S1vb7
On712APTsBm3EneZhz62XoF7Vf4DuCGPEOp4WOISJFQkwpW0Od7n4Q6d9ommM7M/4uUfWvcyM1UQ
DvxHc/VC5mWEM48VDN/DE8w+J39BNQZnQmszfIAX9tlRVPV0XeInmoBpk6mOGQFU1mZnxUbsCWu+
rqDfxQNRyOepXbHpMpPqk67SjwvrQG1mZwNERXLb5gY9v/ULe6tRLDlMUExutCkE6XHKnnsze+e6
zfkHPatYIRy3QAK3BaRp+JIatQdt06R4gA/dTZh/KE7Gt8eeFwMFFZ1XQ3I2mpwennh4GSKvgu/F
wEt+girDL9VwY+ZgCLtVMt+HBP9cMGm6zoGdUZ+ZdK5XfWZlK/zwX+neuIVgUtp2IWFxi885MH4C
lb47O4ikjO21QdOadgXfuVH2fhVWnRCjoy0flwuAH+JnQvAUlndhbxcOAa0cCHcZTyDrMEswKUWA
Mo6FxILkHLYDcdSdUd8p+pfzT9jiMkpqV0URf7/rbGSOCcoVnk3CxMMSRzChqeiZr+a0YOdh2gKC
hwmd40oVCARaBsg4bmRcsGRgSzXZveZH4Gh3dMMMIzBaPsGqfcYpRq/28okoeqPxj8GQmVBXct/D
ydntytv7vZi/A7fTah9Ckpvvt8b/hYdpAEcA74x5zXVKyjxkrx/luuvhdb6Z2WrDCmPZWPZkQLca
MNoWzGoUnI/qhwx8U9gZbvaaCDSvDXndRjXPu5hVy0kPfWVhcn5qL/QxOBQlZyBQa3cW/WUfDMeZ
Q/0h7e1TK+4DIUnE27q1+KEFLTEaBdpL+8JNxAFuYJe9EjxNw9DeAC15AhTg75TsEt0Fsthp1yXH
GmzRamecCYTVoVJo982s6ZZZWWgL86GLVq0B5n2rFxF1o02wGAFfmciWP3w95Q5hQAY9FFw0d1yY
GotivbYYcHkSsnQBkLbHHyaywdY2ZrvVEaz8pqTEgbUP58tXO6Qa8RZMkHHhpVFdHGzw/CaNJeOt
dNpXPwhngEoiwva1kLdnFkyw/NqSGV3Tzt1VPuLmGhP/I5dkSL4is/ndFNP3B35Po0ZG8/lKaCd9
QaqlyfqNEppwWBwoQjSS5d0hAu09VpE2BtsCVZGW9/2S+Ex24GpLZKSgaV/om5IbGxvTduMzOPRS
LrabQDpxqZ5X+VCbs0aa6RM30zmoA3FKS9BMlWlyuw+NENwdedLL4i+kg0S74eu8VnH9S4rMEKwg
x8ibmLBXAcfK0oe4UlVeiIbNhMy2XCztY9tzu/+IqzTosaVv1S0svd+e9g2XJZFNbOD5bs4j6Iiu
Vixz9sp1Z1GUAVrOp2ikzmWSV/mTHDgUt3hPQ1kqQzoNqhBSkMHUXp+yKeM+u5pumHx2PBCxG72Q
AyUTV7/erP8YZM8rbgLbk7F07crNxgFWlvKhKz9ANcVxmD7IDfrqmEklhqIripCIk/ZLZe4w3rVI
1JIuvEtVWCJwJB70K8hA5x0Z5WOL/12prtsuGsHCjARHHFfLv1nh+GVY/SHPsMwIYMGgF/G+87sB
o1p10C3CfHgDUKDOSLd1jxhfsAwNzhzINhop24OVPHYlugxHXSCtYG1iyTogUKW9zAf2j+O70mt/
qC4y+umoRNB/GoDHO1JQkCm9ncVvTPFiXSha+1s7nvGQNEhUTsdp+Ln50Ww5DPZLjN9qVrxNmcsE
fC9iGB27+PF4E/pcjL/XDmLIk57pdIels9KcXhvFOlVO7VDgeB6jWdNsXAHhwxL0qJtzEDpbqKxf
BIaSxoCz3X9WKJ472vStVdW3xMus6sNjtpqZq7Fj9keLN3SklDSFAsqTsbdpxnGnnXXdrbajfbd3
cz12B7Raka2aIXLN5TkfpBtqLVyj6f1TmZdcIvrHYVZQcpEhEIMH1lNbrwjvxJm0ZAWgDAxvaS85
Yib/N7iBEOhfysnVxDNgcfpXkvVA97ZVvj4wKSmPtROHuMlukuMBQTD01wsyOpb2SeMUHoCZXHBv
D31nuQn1Csy5b4cgWBBiPnwLFN/eDENRCdzU/iSPgnNGI+QqT8V+EuEvJUaMaXqtR+H7ddd8iwr6
Hixc83KYLmeimZANZoymecLxx464TPHVrHbJ3eS+qkeEoyFd2/1Pb2TrJAHlgkSErCezK/jFYUKB
RN2LaRJRiu0vJy0iTCTU4hjGGX4MTc8+uDuvm7flt1Xu18yX/lp17M7tnoeAR5rWpH8ID3ifOIVi
32qQkev+C1Y9v8iOVgpXFaPMyBTyhcVAd1w/ei/dxZ8jRVO1UdmeAvVb9i4khTWEtQLhRCGEPPVE
noxq88ygJ2xf/zFMEDgW7oEEFkm3L/pwlVg+/EvtwJTk0Obt3+DFvcsLDkPYGZVgdPexMgNFICAH
Djt93sfP0dD/X9mCclLqG1tSbJULSyGBZxDG6uTD3XZuldBkGV1jiwmHnmpVCOOtyv52NysNvQwA
wMnG15EVeuIbbZzb9h/fBus3kmnDOkbd9SvAnZQRGSRfN71/jPSa9SBOoZVhxMBub7e7B2o/7cuQ
wapOh44KrTRcmB8mklt1f5zzUulKDexfjy5uCE6zUIJVI2gKDLGHQOwWPP2CK3GAGDrRdFUDe5GT
eD2jTZrzFKUa8mkFULbO4Eg/8kxn1ouMdCNs6HmMXnO9lq0oUsBmUPWKNWfhLrqBR25sXehB7oQB
JdxVYqFlxcElz/xB4gay8GQOkMimuQnRKb8GO+aHsoodUSNJp05f/v+HaIgFhhCvaM3gdylXEwFf
x5HltTR31TLihariSJ3N1wYxNxO7Pm+SQRjf+pU6KUBVdMruD+qxP4RGUGR/wktNSL3SEwXOen1B
20+y2R2zj7kFgK9cniKyiIdreCvlmrgq9mJRXrdk/kch4rMpK+egi8nK3c+ME2bAuT+8ufF9F/MI
z0D7yWm9eDS/5tYjEGpQ8DAlkqQbT0tJ3htKv2BT0CjYRlkLDU11ErYlP8cSaCBak5NKkvJHP+Mq
tWZE24cWVDhWir9wuifGQCjftvezn+T5c8V6AORrSLlITO79ovcmdwdgMIxtAlOpKFGnjfd+/BM0
KEQLMsLbsXWy5RGhom91DDtLR0kUWG8QJq8KN+5EYgHOAD6QL98Y/42DrtwIc3EYZKfuZp+eSpU1
RWEhYXTT7xkMBf8CHSM2/tvAyrEVQ4SrcuIQjIP+uBvRzovg/VFklaNGsBnWKk1bpBIWfn28O4Vw
jVZyExEQ+8QquPGYRy48YmMW2++naL+0yjZ/yz+UJB/zBhgJO2uVy3sXpeyXq48yxPkKsgy/zlDJ
PTWeBxpQRmG+OyalSbJyjLWiY90NgEMHo3SHuOOywXi3vay5plm1tOe2E8VVl3METMKJwiz4jwN6
nyEATsx7CNa5pSkPUx/2lOQ4PX0EeH+yK8NrLXQlHhyiJ9pgPtOcBV8ig8FAdhSyBwcaTP3A8POh
8MC9htlGYnHmmdlxHDl0u5USk/D5MtzB3NsPZE8IYuhdwS38a0aKdeFrWW8wvhiLK43kHRp+VSN7
YPmIdsjcdeAPqobzJrVorojyzR6HPDeOtMPretSA/6ykrLt0MuDX4zxPZjeMjfUAwnqpbDtM8urz
8Ns0OdqXY+5pMIjD6vDlKWrSkqtqSXyQmvSfQuvAJSoFpYRcPapYfdusx+xKN+7k6MK9MePDl24n
YxbhUBwkmA5Wo9WGh1cWEJDZrarCMW0egFgUOATrrJljyG/V7ddYPpHDEr2KfQScyrfPc/JuRMNX
iHhcv6cXRrbB58Nsr/93HLi1fQCPpVB85xz8zjbMlavppEGbxrx5aae7QEFlJ1/F8/6a6WdNoOtx
Y+zOLTVbK6OuUlug1lAsrx09nEagJu9SjcEurnXXPLg1cHXVAtDLZQXEM832h1OtuM4lVS4XsOM/
d7XM8V14NsaE6TtXdC5v5Wjdr3B08bsZa9ZzMba771GB65/1NyaCkJWAd8yzcyBDWUo0eIN0839l
F4dq0eAX+TMPvzh4yn+ycYrdd3o3gO0pSpDQkwgKVD6MePCYSaQpArE78mrCcbJLa0Swj3GvVQR/
LUYOQwD5Idnqgjzz37rkbS5M+BHpWT5m6+ngTehuG02zNFZuhwLGOvejjHUISkw5X649gt4tXcuI
TlP0A7gRHuLKhEkyszsNfybjpy4yb0UIX2eCpG0i4zVM9qMSyL6nurqslsD0Ls9gSXeXJRAr5exI
TWsJ0h1MZ1yoEkJW3rZRL57E87KJB9ctVLDbt6tcbLyq79Vi7Rm38rMnei86PkHb2rorS+3ZpcaV
BNVq0pHaVGvv9pv/xeKgTwIx322kTvG81lfzQIvg6QPdi6ETZN5crj8mxaq3J8NCw/UXZFXoSWtA
0sIB9DlywaYJbjSYshqrk06wc9U9v+3Kh/1DRdEvegJrdor+UO/p+yyl4OM1+1Y521n8oVz363oc
KbIZzY95i5AWKhVlN9RzlSaaXK5LT/sK/SG8Bves0PrR2BcHPAyZwou46pTEV/V+BlfX/GGqdwuM
TXp0D8HfADUbP9oVrjpI+rfkgmOqNq9T57aBqbU1PCTqTaRUCsuzXeQRSgbcK0Lgj2Wqbs6SvPrO
DxxGCFPg+JXRnj9N4pcKgRMNXwOZ9gBI55kO4e9hI4QDX+mtbAkfLtXLE/p1blLoiiwRwvU4j0sG
hQrhZ58kGHWaRYWZGNRTXH6Y8mtTVxy1SmwywDtV8S8E5wp2UeaXdkLkBH6MP5DGZIs5WP5SUt+3
b7y5tPjFacvcp+6zHMYzjkip7qxquQG7kBOzeORfsIvSO5aAmvcoJstwoe7vuaaE5FL9dN0mHXml
gZIgHGiRR791YmC6/ipEMmHQxDnpg3eo3aSJVkV3fBsARe9VoPTXecmNHryjsnXidzqEIa0+9sTx
2ySt7qckbD504n3mxAD7FYitbmogFDxuTcmglIdQBPi2uMSRCXj7571PUPgRupCI/KTrJsF2k5Pu
sPeUDys4uuZkVPLiNTPKkH3Wr6/SqQDNEfY2pu6eLMXS0MDjRKQPtD54+TOxASwwWV/yWiHv+nJN
qsVM4sNFbyXatP6soi3Qpe8OZY23MHupbZwRYt2Hfctlq2F/kyymuoBkTvD/HSVrtYKPABZi9lO0
1zSxCGEPE6AjOlbBhb9ejIMF2kntmT5pWFfDy/yD1wreRIilKRfMS3fvkmir1uvAOw122vORiH46
OjwaxZXvqjgzv7TJuB+1YL0D/t3QcR7DOG4NEklPV/L2HO42iSMLV3N1J5OwvOi+KvVl6ehPAd3Z
7lr4sDemGfwEJm1cgH0hozbMWJoBjmYeZQ0M+4t/XBVfru03/5pXDlqYPafhjp/tOdflzpe8Wgac
FcFrLgd5bBSCEOx4k/dkptNlXRFBLZqusBO/MXMmQcg8a8o+qTraGeGp85JgM9APBp2YMHBTMDuR
jXDeENDuRGgZ1lK6JFwFR20E/Ia/jVwyIVw5ydi9Nbd6zqWS103DEZyeA1PW0J1yZJOV4JS0v52f
UUxPcqnvihxNIuMpzgT+hhIKAUVGXASkBa+c8wPq7ePncj90PZx/WPuQVkN44/djBcvLKU1Od0Xt
KplaSqf24qPAlgf0iCMEyDPYe23Rj/voowRRSkpEZ9niL3jbiPrWEoIlYcNo/ypCgETZ4ctMoABT
U/rXVjB/5A8gbrlmQZVuHHAXzJEUwNELaRT9cvjjnjkYKNjePueYqkyqZAGa9FOo4i6yV/h8lZaE
AGqADKacd9Lh+Wt5UQAfCE9RW2ttetYxsdPlWi1K7wbWhCeWovYhg+dU9PhI6vzYlk94+/BLe3zU
Hsb9Fn4Gvj7AyTt693p3FHBY08Afwi92UPssQXIdMMojCVo4/1B1rCeavsnst4RksJVBvHd7Y8/Q
yZp2p4sdozAgFfuOUWxgFLzoc/VJelvx+lkILN3N+hU7vQTXDrVlexGw+zmTLUwSDM1RQ4b1PewQ
Xk7DenDEzDxj/9uKjanC1BOMs/BPQohSjB0rjl3PA4c0xOglGEQWMZElo8muEg9XDLs+iYXWKlBA
S5U2xW6u/8rmkCr3PdEAe6sOf0AldKPaxzKzef8tUtgTh8BgIc4Nk7rHKHMEf7MqNtgaZOmh8Tiy
UiMWNGkJofGa7LebyWgcg1KMfO+oaU85jMad092C+Ho0wnEqW1vHSEgTlFHA/mgvDnF3B0dDgt4z
OJfWMwoDifhQ5fm4crDEw45Uu/jpUULQLIodP3SCz5b2XINrJRVpIIS01EC/aMdFnK6MLyhONxui
cnNBmtZ9uvp1EJesi++OSEvXHE9WWZxYDUiYpSDU2ghHyxMq5rNfg2OXOJ/v1SKwY8sO0hi5Lp5J
oK+5S0uVTcQ14MEu/60yhaYuBKWIHElHqpq6UdXI9Ytd4+dTWKkAqm0luGVXRBJt135Ns2rsuIJt
8RgWN5RSIvK20nYQW2FDuR1QIKkbF9VtHuI/BmaiFrA89DxFkpoVQmOe1H9qUoFhQSVsgwyhA/AE
bGcuAAzpY6QOS/T/BY3jBWvL1yZdr+KE7nbFY2xVSdG2S0bK5FVf/IMAdDllFN5LqgvZPT9MphxM
XI5Me1uucTqgKjSAh+OsOyl6LcBRa8IRcL5vXxGnHkYcoqhFk2ZdFYZ8CBh22rND5JOKHxKjo6ZW
mv0KeGgVem4/CB8CvA++FpUVYkVlNR20f9M5kZAZKMxfuyCMmz3l3NiHGPn2xK4ek/rH5bOJGtHY
YSuRz85mwFvGbBLOXfpMG4CfjuD0FcE10hptyjdnNOpvku3E5gN7TFkLadwn1GgVp9bjTJ3IA7FL
9cxJCvbmGWwDL7kuvkQdWA//Sjq6VCfhxuS2xata4jbtYohUs5C9/PdpzbjTr1/dOrNu6uLiSgNe
ohqY4jB6+J367FgsoflfpphzsmrsBSH+n6O3eAqz3nXEuha6/KhsIO04SaRFdUHAZwpzcMRhWbMq
1F7q5fGZ+s8BdkaQP1Qb6yefhYA4O2YbZC6G52eXQij58XiWXy0Mnwcfkrdb0YEZjz1Dj8CJbYkS
clOKkxvubaoncw9kQGEilrU3xEGRpLXZY+K6qC92F+pRAWTwgSUsepOcHY+A4sItvxnccqp+9a9O
pxV8o98oJK2/2H4RfKMdmPc6Vp5r25NA0wBr9ovFB2iyIR2j5fIf8+ve7dxiZWjwbSwVtb1e3xut
AgRBKb9/ZOjTFAvpxLMJykTBv9tJteUtsX6MeSqmjpXt0GajT2+XjG1ZYePDs9tpr4OjO7mCu4Ez
W4LdvGTl+hdELII6cmPrAbSIHf/Xqk2Jle9iwQ38JnBWbGq3JFA3QDW5dNc/2EAQRhiTRyN0bNXH
8HoOJxCL+Y1XC883Ao/JKmNcUQDQXKYHB8o4dsL/BXkBrasbjGqr36XvaKCjxQJqOsiofb41+83n
aq1EwMfj+4LSU5Vz1pdO33R+hF5w3xgL0O9VCu0GiK5DNhgo3G9WbAmYtn1cCEUQ1J8CgGjk1xKX
ynjPgRNsVe95S4lyT4R214acwCRhq30BNQxyskKFCv5Eux9/EMf5wYQmRowPz0Hbal7jL9MLMIkC
Fe9jqw/hTTaHbLnsZ02bNE8+n0sEnjGyLsJnQ5JXVGAwSP7Qw1efliE/z2XPax6YpSIuLfBBLOVF
5ZOL429TenP07XcnMAYbw2BTcNkY1ueqzaA8rT9d/Pw8dkLPkfJv/HCy9UCIY2UkxxzXdMWKbmKD
LdlSEkAfd8dl+KBv05EUIYUCrgMvT1k0LAkxWO4QOw5MUaKdPHpxJRdmQAZ4rop9ZnxT4fOHGA5C
IY50QD0ToDfOosiCyADRxGU4b10T4fNg9bjk3a6wk+gqFgoimY6YVYoowuIwa52Y9dU61VN025rO
Nz817HCVacpTbxOI0qEx4C8SWZY7NEhCHjhTTmcAqlwMfw8TuC6DzWqXXAbUSbi3KXekfOHUsLGt
YWSZkg+yHjL6qMIqLLtZtlaMc8s8HnULHyn2b5lZGeij2dMzshmmjqRfavufbpCH9nPR7ra/yfYg
7+2RSMSFZaGWRqD6AJT8t964kj+jFi4+DbFwgsgFseevrvtCv4VZBHZl8S3p/bcJN01hvxYyO1Oy
ozEQ/Y/+QjanS3znDdLCSe/woMgIobU4sRRzZOWV7nsNMuxQRxvQJJGNyiEwUBQarAo1NG9Ytwaz
5YK0QKStEg2lBKQwE2VzdCeIN8PBrCkVgm209p76KL2a+fiA2EQXgUVoEfROqYnrRzZT9pijUjJS
sMMw+xp/L9D1RfYHy3pEaHX098dftFBq+dALVngP3nVP4EUnyzRnbd+zxuRjp4CCYcyWMbf39sIs
PPaoH+q2S72nkCSLo2xFIyleYCsCGXau18WqCW2H4nFPprCRj8vFzpbO46aIm6jAn6BXgremcS/8
ihw5zfiJ8m7TNz1lFksDt23gaC24X3ee0IniyVlOTcSnI9t0qEqrt6qhJa3PVIiCqgFTg2BvCK1l
rVmOeJRbi8cd2LYWovATv8rOfBJ5K5df3Bth/q7tqeAh9kGO0kbTX5WQbsN54fjedM90J0auENge
MvPO/bXAp0jv6BTSy0T/vO2vJ7Pq+0bjLMWyfyEDl9iVSEhul1ulJWFn7hUMvCQgewsL2t0UGh4m
Yh0ELmHIbjzZExN0ngLCh1Eed1ohKapFEuIe2vV77gG741kQ2mJZAg4fSMsHgb8XL7Eyh05o6DXY
pzPmoDnZJ3/SdtuRO/7X/7Vqs2MjcEdIZCLL99kqi7HXn9mw7nCaQTWQfuH8SykxmCRsYlca9mts
89PAcPoeUKBVZndm0o8OBeXBYKTAm16DV/MBJJDAaVTB5yNd/aEXL4dvKaA8WtUG1zaygBFoFTnW
ngLrRs4sFMWi2TtvOouGycDhN3BKsvaVEfBp3GM8xSQPAP0MBnIPs+RtOraZVgZqGO7Gcsv/TdA+
aMqcYVchvtJs+JYn9/pyVnKvTB6v4/JfgzBMrQoOo95oEPB5IDeM2a4fGN5vC7ua93v2wv8uicY0
IOPg7F3DQYsNEbziy3zBmNoCX7CJT8MNTp/saMtHyS0U82F2LaX2UaHHnoanVZaHPZJBIqVhYrBe
Se8peWN9+b+bqdzzpIkCjnIB6i7/iYnBRydvlfSroP5Tfj2E97gsnvVOj9Ivz7jo7XmlLBzUhwEB
9r3eQ7looJeY6OrLZA5o5OQZKUIN5kutYmjEh5DBCHpvmjckRqZanBH9UeqB2e1p5L2+DYt34Wfz
Ciqwzarr5DMGNrE/VR+9QZb1FcYI3cFshj7bLEIy3OxabE6b8/r9n8xaSOGkzR1Nj+WLahIcxcLB
zDahBmRSbBXFO1BoskucfBy4TxDuRty+uieQWkcdueWNZxzwkvxP7pZQxYbma+PINeKsTYUg+r3m
Y2NSJuGzx+slIcwJWSuEcD8QQGIhVCYHiovt08kNJdPOwRbJujfoTlazJ3w0sXk25uxt6lXhp8AA
B6BMYb5+a3MrN8s4J5Nme9h/tE31SBqX0p7RyD060GKN83k8X8qWECtgeMsmgOGMiz6Hjswr0mkN
V4EopdEAUo/drPLGHoLI9yhNfbeVifUbbI3SQd0Dd8dCZu3ZnLHo2RhfyD+bv+sPctxO/RZlGjjG
KBBaRg8gevOFCD+2tJMtpdpQCcBA3cMZSKzhEAWa6NN2lDVfmXDFTvNemLJsUvJxUMZFr6EXN055
cfXiGbnV+0iqN9v12ROTQW+ZEgvljBKCHN6iaof+67yCevuUXiQtWt5LjDK+kj+7zzX+AHfswLS+
36gVH+kPrwBTGKV88qIhJsNZ2DPZPPBtuLIFwYq3eE7aB2W/794GmB5vEpYWYJpyQF9tUK7WiJbC
04hx+kEHCw7B0mlgHW7Ks0SEwDwQBD5W1+uvFgt3P6GqMOUL+jpuZ47HjdZhwumX07nm0Llh4wJp
NF32KUkjUbr2wVFO96Il/paFpIYHtgczpVOQ+3uoBTjsJp4XNt6R5mtecoTSYlztBRi9H3BHfocn
YJfyFrst1W5zfKgCViFMaABcOKjAaDGXKOo+o16RjJ1McbUTCAAdlrxqcVYKGuFhVODucCXi6cdO
bj6KLdKnjDUQbUy7iorg5oT9hdeo5Hs9RtwGWAB1yiYjiS+ZyDxbl1XHu+g4mpROKJkz7EHgplVV
cawERUS1pBMkUVbuT0C0cjyLI3LvqKwuK3z1McdtChoFqYErX1s/h/UEcW8+fMmhVOXv+Z71Mib2
Ix2TiAG4IRe+RS5H08XVRlxW/gpZZz9u9/ekK8FeUh7HJ/YR4h8CzzXLfond3aggBjc0Vh/7riC2
jQE7rn0tZlMNsistJhmV33BoCpsSPKeHSAoM0TrrBr6eFFKlaZwEDMrHt3/dHCkVvK+eSo29IUCR
yn8gvdjXp02Ml6BCnacnIWY9+JJVLfqZdyvdhEgMJ6OrEWQRJZdpaDOeCvf8/fR9Cmd9o7N2tRXl
i+oCU+ILb9uv99OiKaIqUvLs7OqaNJs051sMvWWVteSbTwQ2C9iKMHmHxY/8MlsKLqpWV2GbYSB+
l5GjLAoBYrL9rbomiU/+kjbE/CTW+hVIivN0g1SIzj0Dk68CS37NZnx1ahDQLqYBTlK/BV4bqXfC
tw4mIPcwQvR6Qarz18Up1+DXt3sKOqMfG7NbeS2ydXv/t/kyhNO4cPTs6zC2CfRTA80w6UH8oPI5
UKC0LDoSZsCka+rqjmDCW5IPJB/HP0n/MCAZg/vCX8Xlr3V9keu1iVmCSFxWz1P/4mjVkKZg5PiR
gYJFhojM5pM8ZBgboTMhpRYdZ7L31YWekwSPhXStRjuB6p+GK7NdF5IzqPPQ3mAtuNSj67FEfsVl
3EGG8T3Qyg9iLA7lt1l2buImknXxntp4UbnRzdsQMN+YMTKTpycVobLt+cY+oxUJ9GIe2Rf/Tx4A
mZzdqffETZGYZ2gUk6mzRfr3uwBivn4kqtcgNt5th7ssVJwSq9RU4GHr43pMYqY6/mC5/bZq01tH
IaTXaE61dMI/CM/D0/tdht9mFfYCLLgJbHQlGGM/iHhxTiCODj/QbnZr+FB9KLYrqf98gli/Dwzo
zliFL3ksHUyUe5NpBnNXnq0YBnbSqibGjOc/WsDB9aiyXeIv28uePx64qM1XDjpwGvCfpdTnMsi2
zZNvNlCXmEPzHRlPHwUshZvD06t7bxoWrXIm2Bai7iZSXzmXqXNZdMbYOpRUQKsCQjlOG9BuW0F+
lsnRbNcDnE2V+XNso52avHzSj2YuakFUYwtXQTC8BpHmrrmU3pfPgAB76iWYCoYnkQ0Aqs6VgZSh
zdEwRVBCY6ys9tIVEeDD6xxWsJHCgMWT89A6z3zbcJ3T7c25EihiTZMgJbgChurpqVeSsFJCOAla
CfMP66z/S25/tfkabvj4gUhzvha0jV/lLVXKykhh0ax7/c5zwzecGqeKnb0ey6GbrHR38jOa2o+l
UVFuW1A1XndpEOU69RO4GzNv5PVNVWUIS7L4sVOlk6k2DbU2CE3tdWepCMcgHhkFdQh1JtU1nSZz
4F5m3bFqMdgoXpeTAInBpWOPOIGQCuDCQ0Ru0ySfMjK9CKGUdwdk1RtG0ZHafPqgZzcmFlHpzRtK
RqEkCps5SMdSSiJCEIudBjPyUKhIKPC9flNPePnGLXR9HmWeaxhWuly7UzUb+obyFoqp7ORss4yg
fgjLCAVbaDhxA0mpt5ivyrzUeMstc78tGaUCM3gqmbE80ih90HNu55RsOGJRasFDcp5e4qWMXsS5
P+sHNWcwSeDCpEP7IKXIvw+CAW/uB9azc2z25kw80lGwGbq8aU2p33jSOxfsw35BbyDYq0Xn94Jg
weQSpxePxpnUkIYo6R0ffJrZgixKN8hrMP7R7L4SRSZVsNHGU7MySRwZbBeBTjKDLcABOltcPKyb
CcllFF9HIb3aUbfRZmRP+Xhs+oRpHMtFE0H27nVKnMgzuj1/sALUpFgs3l+IMmhtVRdDeDoBvOlx
vCwzMsHaAvGNu3u8GXYBScwLe2jpw1tRbt3eWZF5P26Palg0H9XSlM7AksLaM0q7h3Kpy+gcmb8o
oquiFMm3LdI+kqPPKV0DfIK5KXYXEcTSXhFeJSQaRMaEGe019m/EuJGZIr828njVVARltnXlkkab
J62SG6eQZ6G6iY5fK98TrunC4ynfYy276OCnE6vvlqQ0+guWjdNA5l17PpS70aczg7QrEvo7U5aP
oUoqaipVtj+WRbAqxZSzyMb5h8N5hGpRqTDKnX6nLTrsGtZWrvacV0LdYev2S5bMkED8wOumAtML
jC7BbZo0OezcUXHujDBm6YLi61tvX6w8i1+PXP87f0Q7F+ugj+kfVH4+9z4bHXhvRi0hy/orscw6
rgc29cAkJfNGEMz2mw1Onb9xT3Ejw5zNM0I5Skp4MhwV525ku4r/Uz0YPjxmALX6lhTA7Y4eyMQ+
A18Yx57L1PkEvLBpNp69ZyqVNsLB+EXsOuJY6fF2O/zxSVJeRxcMhfBfZJebd/CCjvrtvvR8dgiQ
kncLFsEjJWbWD1NKu8e9gjW5ce9FPn6EUUfRLf3uQqM64msEOTZbMbZcXPKWBLtim+Qk1uycfgJ4
U2AWK5WkxRH9KBCszKubc5ZdIMmD4WhsK8QH1kynAKU9F2anI6ftuigz4yBFNAKlxUbqWZXAlGVs
RXp/6jzeaJtrh17/oFn2gxtOqQ0+zvNtP8gEvrZF8xi3Kcu1rsiAf+zVt5xyEk3lku4X0j/hhJ2m
5CzYkIiBPDKAsVJpQLIaVafPLDPmUv8WMTXeAzdMIIVJDOWdEMi8nusWGTgekYcSjqJwJSfiuL3R
fLe05jZreRQ9fQERcDUZc6VXRr+P37Fws6TR15HuXMj5TntwoPKj6BiNXliDaBJpi71JiJVOiW4F
d7q/N0nDF/JGng5WUg7jmAFvK7MGiVblZaiLTpMR4pPSSqBg9xBYRElUMqu08isNB+d4qhGGJYtH
CGob52MScBpIj7A2BqFt9Gj2/slCmRglUoZHIuiIEKEbSjDAfdDiBrfrssuaXXwdIMsRWLxflDhQ
+Lqn71WnvlqfGPimcarpZT+c5flvGhGwgm8JHOVT7UwpiQf/B+BIreo49l87ROD+GuzhEM8f3/zT
3pEz43VZnqJUC9nFjKRk+fWxeVh4iXLAh+TKw9xzVjvH5cRIBixr9ok3fHGaDiWkeCvVHa4MFCB+
V2K1YuDv95AMAPBEguNWof2wJPAZP1Xf7tc8SOGdBz5j9T8/pngit32S/OnjR9Ox1sOLlemDET+S
a55FEFQ0EJbDuHcvmUjVVf9K0dT81+ahqOJLwhKBnlzmx7YyZSk2HNR7xBBKWQnG9VbOhnH3v6av
6HxtyyYBqB6zYyyICf4W6eClmpzIMeasnjR3Kg1HiZJdxx8CT2svrt5FsC+WMJRTd87T7LQ+RFqu
bo9Lx67WHaNLA2eWx1AHvujedtGqdyhZVqBs1f4qy2OI9DlHcix/Y+kdyjhIzWlr8ztQ8IReLjdO
7s17AJxRDIBI+CUfyb8DmbgZBDmkp7C6e7JlzSPljBpygQgk5fXeicHdmzuBJt8vo4u49DT/yRPM
QfenNw6wBEW27lu+VQXutxsngwFzYekEEK2TDFCKi5fNkMh7F/50rMJIKmpMlLnv/wHPQMyvZSIu
Q5cOFDVbkWUvsAEUVG4PIeHJmXUwh6+QPeuZdf7H+fZJR6CATQixUYhFLYS5XOnQRDE4GXSBa48I
yCMex++JYpaw1/9FMQ93kVnrnh37YaFb8VKQvda3bGR9tOi6Hob/xjf2afau/SnLu4T0zkapwJSe
j8PU62HJp6xX12+oiV8jEy+A0g24zmFMbo4nPIaCFDKrQGX1LYw8lyGPJqyM/oWSE4W8ddBsfitM
0p4usTh8rMVK/C2Df/pB53QblTUpAK3IXkeVfX4p8B/3DClk8HwKKH7dgn5oqiYDUZoK7w22hZ7u
kQwKenkn/F1yEsrNpjKHBbgH8oTOC4/+HWvKzTSv0cgQvmMzCHHrdUFhM5EGug+o739i46Z707Y9
t/WEGdp0YUFS1nNKqqRrr+nqTCt11gWwQkiFP3aH2SZ1124faBemPylaV+I0cucHXkXlfCu/9LF1
Vb2DuU5tziaq16RoyFIcgM3vag0B+YwSw+FbkRowgVDynHwsMGVKzO0qCSDYRbiUbdHTNtk2klZB
Ti4C2/RkztcFtoUYeG4mHt9aS7JN0WuIdBFncga9DqTV3UyfQbzbw/LsI9+Vc1S62xVbqcre7KFl
JKT+Ryx6nIVc8agYlMqhWh8JVGiXRCM1bKMEguFQGK0PUdv1aWne0LgaYoGkCH+Bf2C9HbNKXpAC
yPVDUgb+7Yu1boeAXyVwg2wMslXlDNcm4Cqtp4FyTAVRzw/em9VqKvj/O76qXDmc4hP2+Xes0cOK
yU0G40x6K73ml/KJcThC0BtLv9UhZUuIvJoNOPXbvPERV/DCRBUmkEuUlRI7aYG5TgSnkAapBE1a
SVS7SU7wPZBQlDObtEd6exGQwfWCjnGWyJBSjVadS8A+c3xBsJlnccmxW3ZgPZTmcsZmDHThDHnF
n/4Z8j6CBNUSVM0VPamjYMvCjy3Mr2z90ieRW9HlBiF/BZGUKq/SqHYIcBYn/37pqV7HOTDTLWKJ
pzJu5KJCELlURPvcLUb4Z8QHAtQm/CveXKXuhFKCDrR3JFVQ0aHVltSDFVZs6gUaMtiXmW8K1v8f
VNpy9t4ndCtSExjEIYsyDlsxxzaBEos/BeQMHCG/uvXnTjYvvm4iTciGM2Fr4oUsS43XTivhjreU
3tAeOpZdmHdzvXyqn7GKTPu0VDuqY0KAiDAca9IG6vMKY6u8b9AV5HSS7jVMAX/da++El6DDvU8p
y94zeERoNpznk2uWoUZa6D86Y3Zhwj43ImrCKr6SrR5c4kMUcQYvzs/rBbFp8Ex/PZRH0AHr1jL+
KYnOaWGrG6ckRpt+9rGU4rAcq+ozUQHniXJ3iTVefmP1S3jaKl4vHVN7dCL+Z/6ZAB13h7Ws1I8k
+o7M+4SgkYYWqXQ6Sd5KGlMZjEckh4V25AjGubtf4BLmwF6n/sYffZijsTW4AeZ0tRAB6uacFfNE
ZyZHTcHuTWDhd+c/+WROIL+wNU71gTig+eEXLXIZEls1HBBMyEHyJAkDYFgA+G3K9UN7bnB/fFDq
+8YivFJst3pTmYgVk/57my7BPnZvQbiThSreJZuaP+bQI3Ri1ONE4+thVwwRP1Wkw/2vDs9V9XEw
d2Rxl++Doo+J5gYS7cG1DXHjrEszOiVODvZI65GLPZYQPz/eaH2RXSqrduaMJozQRz0bGu3YOFbe
Y5UUyjTnH715VpXomp+TunEpv+SgI3ioc4TQ62utCJSSrSvtiQ606mihGq9qso4J0xQW8LouWIwZ
yD3NbGQohj7BBnUJDKARkXChKEK2SglAjwzwINnHy4zG3kBauBV2JcX/KSCtZn+ZqSZ44ajkGbH9
OPjSjUjiszAz/KSLguA1VFPYSTLm4T1mwvjBb7Y7N7ceJbCk+JtG6TTQurVX4kuN7Jc5lArPRd5R
svtvWRKEH5wCmj6aOovh/Gs61/r8bGKyaT3b9i7yS1GJr+M4Hjzn6XNubpKQ0iH3V8cgrUCZcSiC
igZd6Mbus+9dJ2NJrnLegZ8o+5Rypda4xt1mSehPrxSJilOC31RPO+SQLDBqSOOYm5Xqq+M/uVV0
o5lDR3uriovsHh9IxwphhIxpHd1nywtHzcAx/oQwlpibIf+h4oWgG0Yw44nyuoEL5EPW4Zhz2unu
jVMhujm1wlTozP2Jxg+IynkoQT2nwVBoQNGaELWORhm7xK+N1ie6Y0WWm0TPn2FaesxlMBO/Pmn6
/68b2re1mO25dLZpuJ1osCNB7HiZSmUVyXcE0oPeX24CqjD5QUhdqqLbWAKx+oCljSOucT/ycPYM
ifVqlANqXFbinl3ivJPurUcCz2wkM6+nzokhPUp7lU7x8TcUR6nrpMcdnIcEbT5HfvLl0FsjYyp+
Ywjqvv1sAGxguALtx95XUUCyVqMn5WKy64jIhO0uOsl+vwDJPU4iCPa58uVTevhDNSQqGnRx8xse
pvIahIgDftgOKnIj65lgR9ISj65wI76MbTvwXJ5oy2s6+92oVoQGMp5yJvrdFKf2MOolNzv5OhD5
IfzNvmSUuqEE0jmu0U49QxfXNBJoe8AFFKsHcx6R9peOaVFv9kLn8Dx3r1kQEXxvnZhQr8jzLk+J
evt06eeVQcapufVV9oe6DA36JGz1W59SpZR6PwqW0FPmCPli+FBIfvvDZQLgcrT8xG0FvagaG/hy
oL0exZWchLx/toCW6iGAjypvIMPexz0V03D9E36SPdN65p1YE1zGqkaP9riXpfwPC0UY9JZFDbo1
f5S4rgocmSS4UZ3bXySvn/u/d4CC0yPIHyHLL/VckBfBhmrQBIDH5LWQRuVFvIYlrBJSumbY71Ir
XU3gN9Yh0dUVidpn/Ga4QFpvgB5Tv6EQgEnMOem2Tz4h3G7WkyeklRTH+mj1qjxC7Rkc4E9TV5E8
F8j2cPZqYBkrV1YLWltJO63a9lCnJmTccLDWtVRvnK2vY0qnUDSEVkdWGmiYhHAQ00S1cPIXcHGZ
rITCztZ1c08bkicoK11L8DDq4CwhO/PxDsaEGTEWRYBRfIVhwyL7u4BuVVNwJ7x09yextz++MT1Y
+6b7Flff27wOloreFYLOirT6hKnnFj3L2YQZVN//86jquYprEzrH4GaUy/fn6D+dDg0GDFVV8+c/
fTpIw+Wzpi6/9KuarEcvTFrsoIeZ4Qo02VfY4GAEzLbFh+IR5gC5VAh6vue0sJPbZrg1Lu8JTqM0
C0zNaDKRpn8gK/KwMi+XMBd0EfLaLBIWI9aTDNpL0KU3wsgFrY0ZIbE5oBF0SCvj+FcGnxQJ34tk
f05bMApUjTRV57eFOItpOr2Jhj4FOY9kh8XqLcQ3XjniD83PjkkYMeAlRpmPykpdiACUfAFVhKzc
naz5b2RgFKaaNdWBt/1IKFM7sKzRbuplhxETD00Y2te/K1frqJBnUIaQ9CRZk7vf2t/eXfIPNll+
HRiG54qPH9xxp1F+oaZGq3j+ZusNvmV4KufA+vP7SC3INiUgTeaAyvHydlSkO192Qd0uycT9PvGI
2NKmXh82FXEy9/WpA8d3gJEfO1eX/YR3V7C/0vuBvmZ3Og4vC20XEe9ywOkLFEa6HiaeTTyauQyu
VnBvPSKX1TDqp9hNbfQT/f2u3+YQ5z7LiUZCH6i0YB2DT93LpFW2Wlnyvy/gndp1ZgRqg3u2qZMX
5VyPW+BITpzTR971sXhgLd8IkQxiGdeevDIjkc9Oz313nKCanjniqm7q+EjmRpSfj2Rh8ex83wz+
A2qlGplCjbMQFLyiEJ6+vmhmPJRnaiOA9a2vqeyVWmslwxhUmdaoPDTa1qWSE3nNiWNAuhiHR95e
uM8sJGR3Ddvyc0CcHz+07r6Znz/jl+PD3IQuhDq9Rq4YJYukTzHCvXqXuWUyUs+S4F+Ns4KbPnK5
2TuhrGLBG9BLV7JTyeS0RrNnSfwybyTCOTs3K6wnzxXHQHp5m6bFzGHoshizzPAkaQz1Trxf5q7n
nkyLHzRKxxOEGEgJnsSz1JXWdZByuU9X9n6M7aV1S1xuvlwKl7U2lAJzzpBR1BG8lJm/mkdGcpbo
r8cnHIeWfMwcXgHvZUcVD0BI6jYJezNiWlFMUw8EzYcGiAFSwhp6g03U3e4E6abfu6TqnofuRo9d
vOjiBHcMZhKSGwmisePXXsKFQjjTktQUk45EV3MzC2bFgPsvQH97aeZPYgwyrgC0HQQOmBk/4jJ5
hp9kjEDjO5Zyt6l9SDMZz1j5pBMa3DT4T2vg38Q0AJwLqqCNlWKX6Mfu24dm5SSoVLjAIcf0OIF0
5hM/29OS5CcXua9OeBwRCxypBC8sLzTiYnXpj0urcmLzbOvnZ1VQ8Y4gFAqzPQKcRzZT/e8/3Fti
ZS4aXZdTEnwADvglXqg96Ibz8wEtYr2fRgglgQuyXWG64hCkj/WvdemH0Y+rkRr9PRfvqeQ1PDJ1
uzEV2gTLESGCtk+31i8TMvNUDSlvZ04L4Ay8RCOzqqsqkwGausaCtGIsGXotaFduEbsLcy46LT8D
PGML/CQXbEpDc7eg/ACkPOSqoagWAPYOzZuMDGhaOX62fmzZNTJeFC4CU3VTiSmVhXm1sC6rVPWf
kFPzmwjf+aoR4pKf4K2CNaVy5fBYoKDhx915hzGXjN9aUzFkIDalIy2nVrEnIwDjRz5HYUJwkvl4
7iERv/dJqbHqUQV4k02Dy9+uhtKsNRDrYIjcqd9UcpX2peimux4Sr2YE8l9PZoBi3PKAFsNerEoM
Dn0nrjeWosetA/ECJ8aAPY1v4gaWWbBUjTwHjpQP/kA55ns4pGVzy/CAWL/YrFKj+u4UHtPsq5ZJ
6ZMao9t1xAlIYuPp4uiVfExtE3w0xrSaXA5WN6MO8f2mcn79U/g87dVABsBrF5G26G6CXS3FljS7
8bdT0IJdOhiZjAKIq7BRryl5lbvPDmVh88y2mbOHDjw/ePgQ0s7eL3JyYacwFycOpIPkLpSrfLnc
YbFNdspXFstrUtxwUnpgw1zhdtuo1NR6CvlhWRoXUy8tgSPKJdMckCtm7PHRRSXJh0+MuNdiLrOH
189d+YRUFIvbu7sd19af6RTP5ojf+liMrvpejK9aR7FnVyhXbkSrTDrH7NsQVTSxjc7n0DmE/4ah
b25Yf+cYjtpxfddooK1/GEvTDxlnnxamQiZdE5fR8xOzMEc9tD/7itbzs+pKWDTdRc/PXk5uhZkP
K34jgAxXL1/pXyRl3o4i2OKNZw3d2YeQY5Ml0um0+aS1As5RKif7PfxZUajY4/nVnzcFOWq+b5VM
9ZcEp9wmTEltsYy4WisKlGeMCEeJYlPG7PRC9WCtkxd2Tda9GjOo3wIt/I60ayRYEyTlA2+FQb4a
gpkTS4TDfBG4trez0x1KvHNnx63tMeMXvJ9aALvD97KRd8SGJHhebuw2FLgwYLxD06SL5nwtVbN7
HRMtnlqctxGOFjVhrtCnkP3ESIra75arhg6cAzRHZnnRXcSDapDC77boNXpbK4jscKfgIMX1WoHh
f6OAQLtnbyg4c+yBWb3PxvXpfPA/VUtJ8M99aMTkUtfpizMpkzVrKE84pAEdjlj6FeBy5LYVYgXZ
l7awGvaS9GjdNnA/scz5vhHLVEk9rXu5GsvOp95W/M7zVjFvSD8DRVu3sDIYluHXICo+iQPene/o
oM21s90zagkXnRfMb+k4FBVoEkYqEV2nxOrgcIuQQcy3PVbPo6+XDi8TXNfR4D/Zp2jhdf9d0JsG
HfI9lQwthstAYBh1NDJWqjGnRTfWgt8UroMG8JYqYJpABj5fmRY3cq2/7S3lnDwE6Nztgw6a2F54
Xutx1tRB/QCj306i5N+kSu0xJgqvbYcbFiqw9mgRNic24lB7YtKgZBHLBnFD6WC3pONJAwYmggWi
aKtkUhG33uHv3Wbzjy1FlbhvSHS53XGtLUCDMUapkjqW2HhCmCerNg3HofKLSQfdwAMZVDZm6Ehl
QpiNnPZml8GzTQ218K/E5BTzmXb2/ulEtW5bpyFXwsnwC8kANlXeai5FTLwRHoIqSFjdGcaVU0VU
a/d4LGPpg+my6xSX1oPdbPcxwOZLmCiYr2NFsY1vi6AX9A1989wOj4PqmbKLDkkCzrNu9LXhFkKK
H8f7p+8YbchkYj8jQlDWTgDZXu9h2tT1cMT1XW9vpCeBfrOktXzJ+ILJCfdzPptx++NkgQaHOQ2k
kN5IQdbFl9vMsO96mzBKfuC+sHGVEORfWziiG/Y4bWrTbGWUKe0rvG0Sgfch3WWQY8mIWV9A44Xz
FumSARjJ02e9Xx0DP+Sqq2WKr4mbEvSiMUbyH+cnp8T81Lex/+o5q73vEY2Gv4c+o/7FOEn3etC9
TB7os9xsmfXw/DBYQmRV5Nz4DgRyLkV0MSC3OSYqnCkB8XZMR6YjTgdiRzGBZCilYRbfDPZBkJYI
h2N2Wdkeu+bFG4P6otpkm4afRt6sRrujt+S/W7PJNWFIfuZuqmVnM/6hZwZ7HnpclmPdo2VLt8qc
C67MLNS1oeR7ActNwh/zV1tnNeNvw5Rjc6h2p7KgDMYKpafLmrzM+I986MsqOH0tjZNpWIZtGQWv
StRxde1OB9R1uM7B3Q3IzcgSd5wfpMKB6o0ksXj9yBcJGbw95x/7aK5DazmE0TrUtref376ofrzK
qyESTFXgc9oxQ9fpSoXL0TSDN6v0Ky4qVT3YvFwiNfDIKpucrjTJncgwlb3ZFyNqZiM0gEuEBpxt
s3sW85ui+szd+TI3B68zSjShOk4QKiej9PdAssBqGC2B+IiMoIg5oNCvC0svuFnhAu+DZYKqck7S
V0T1lQRAxgCDkhqoE2ODqGyBsb29GxlIGMr3lzgnXNC7ngWgIOb9QNSNAHQoDzU2z0e4gRaNBRd7
bDvTLYBIfpfzrMt7564qPRoPmBsQmJ/tAwO3aDyf+HYK47sGoNcfm/tTrQWypCjdev8W7MeqcJO3
A5uOGy7sFwL3FDTeZrRJus98x8nOxdLxGFap07gCQ5QJiUFMhEjLaP8zhV9/84CzD6FMOS4HCAYV
+13G4xvhbCdkVtVdhPpwu+INwLWJP6YeOC34jV/DBkY45FthIb8dIKwzpKkWh0Jk2ddilJzOBj+J
21zAEzbwkbqc+VCXQhNhFM/rAq7fDAcv3WNAEiMrSROujxpe3RSCqHe+HSlKXc69E32lP/vT/OdQ
KPgMInqqthOo++G8zXagXXRQaqpRDXTzrxiWvG3chVuBr/YRARMqljh0eUKuFY2WV+CVyFm3wOie
HEbSmJ8pepfeHfQ2XrHDnWNo0NORPPtyg7TNjIFE2DCVeeP6/GORQjKi2pLPakQcMqLD/3Dc33mB
SdgLF0ca5crX0wawXR+zxt7mP9iQnh88EDIHsdwJIrXErpG7QLS44tJ9GE8TFbpMjz7ES5Ph42wg
D1phlrChKTA9cepyJ9oaKYFqto1lVDVXkv7IW9oMw3x313OD0Lm3oLDt7QXPbXzKh5IZjfGns9+g
5zFcigmly2+ryDnntBKrJBYH3J2O1efvZ+XxW44+stZpvZ20rLeBOh9bykRbKNxsBHoj1YCMRqd4
DFA5BdThKPVDHcgFgUB8QObfP5d2XrkL+I4toLjXAkqpbKsapiB//kCTDzKm8lrRu7rFQJ6pOOjk
Nmk21eHhL261an04+oaPAtkkMI0txn8K+5TqpzXsiJ1LJ/uTSZSOZ02wNcCvpm08xV1sGAhK7E6M
F157uOq+c7DvxyjeSG083X6IFF291bB1r3p/49sd7q5q09KISVo+DIgstMpVBdhGd7AsUVZqFg1Q
ZpUIo04Ql0BAV7z0xYKOIR40PfiWiTfHVZ1gd/b64S6xpahMPeANJi1DMHLXbETUXLUhUA6l4nY1
Xd0eJle+Qrx2DP9HUVTm5S0jA6TIG330Hq828mmi51jy4G9zeQevNvwkJuact+WTXyXuG1cgrk7h
Z+EZT4zUe+EAJVvzL1FEkvT8wCeoVDEpL1WppipibqbYNEs024B25EOd30rYqYp46TJ/t3LvTv0S
2bkbMIF/xFbBOSGGJwDoKcLhfdI88Gm+4Mx3HzCN6rhpqZKIvqmbQ0q4c2NT4dtQxIKBvawtwliA
TdSqCQdLnyfzedRV66x2gLWVgsUJMfh6q2vJ98YheRrEarcuixAZolbY3QDMIgbWZ6gOQTTUUJvU
hc2xzgA5mbi26wcYwn/8vkmU+2L7jqfdemBnmUHs8ibl3o5V259tuSPrna+kS0VrCnSeuOCO8jvJ
ep5f6bPWGRrJ1fptfEXrdzR1tXSoqzaIbwUJ5P3lgfRUbZyFaVZfGgUa5VepvQ0K5Cw73fQkxWfz
gdPlYYRXAS0TKu6S5u4YqykRA4OxcsfmdVTUDipYLcMh5/qPpen3ZZ+73FYQyXhzR4uKCztt8s7c
0ZMWAtZYXhUAez1WM6YzIpqkLUOnlzTzkLhSv+1HOM1MGnbrNkrIpYYoCTHOuByFb1YYAZ/+mwqS
apTExw2m5UpWONlXZYgKpbL9S9x8JzAEz3w6u1qROCrbMsvHSrZkgiOW4J8396mmNYueWXs7yFhs
K6asoiVJpFRXYtJ/JGiEBIhxyzKQnBq2KgYjftnQlBDpcjBJCM5QQb6eQiOVPW0Vn8cpXsCXZacB
curdcQuBAdF0a+wJFJW3FTGrZDzg1KAVNkM/Lu+40iEaBK86tyhXY3yiIqJM/oDDJ7IR4wJrFwoG
ljRVOd6sBCxBrwUMa+FxSwjUYpdPPccHfkBFZ3+oUlYTChAsWidcpp0Zxx2E/CaziAdu4MT6PraE
iNJ509RxQpQVcENI1OrJk+J1bjSO8wpH+u49oTwyZwGngod7hQdJHcP0qAk4S5YXJIMBKdtLa9+/
x2/HDRHaQStemSo1WRCk9wLPY1QSvEB2UTR9YVkoCv+uXw1L0JDtBUh/PmpUxfKqzUoF/yi3dF1i
Rja6MJp4iHm2PI4QEXJmjzENfG14AN0caI/Whcw++hV3FO4ZtBwSQCa30z8Ce4b6eh5uutLoZ68I
dRlP2bMODfyEJdPIdLbvMdmPX0uWXUvKNM8VrxsUldq9SmPsmRlhpxJzF8BiMPKENQmpHSjcUTgv
a96+FHRi7f9YFQgrPuHJMhZgAOUAdbvRiTpFsJqq3R1vpd/2AkKQgWTPaTr96Eh81xNZQK9RglMm
TpzM296GO/0wVl5RWSPLVzaoPHWcKYgzbLjsbODf1qrcYY/CZlFUchBonxj4hvMeWaVyJOptYlaX
KIgDcmulLa5u/iIMvCSL1HxEo1zZ0E8JLiv/cfNT/fchr7U0W1fDK8qo38q4J/GKctwe+XSiw1kz
by7bmb4ImFECvbD7GXvMkO7nLsFQHOZjDrG1NPee6v9Li/wfI3Y480NGqa9yL3ePmXh1m4GZ6e3B
ehL9Ye/chtAFDkRkl8ztJ4I+3kUFQ7BGo9+Eavw3su1X891WPQDsVCEm0UU3BgGRDXIA5XC/WQ0A
SlsX+o5yh3DIc9va0UEMo/noOT/itWP765VLgX9NeYNsCHQBq1FHs6heeRoz3GMB3aq9KHL4eiO8
LtqTyDwSeaRyEuwBw3SH6nRgIqUWLAk8QZEreLG8ynvM5Qi4F1sq5O65ItNaBd/QQliHQWDg7aOs
8HrYfWJUgZ8Le/7YR7L2zwUn6gjk/9vCzGCIJFDyC1Ci3KveddrDtHTlemCm3r0O+YAcXgIHzUMG
2I3V20ddWVGbGx4HosxMXunJcKhr8mb8ESftMV9hJOQ530JVBiZgr//axP5OnHBmw2zPqEbPqkaC
ayKKF2t/sB32lJWXQ9N7LNKsUQKOHoAqMfdElNbt4ZCJ1EvP1QSmw1k2Nkb7K3+YBrcGbIcDqfNV
xXC5a24gWU/Epv9/8LD1/Egjdtn1JCTLJBZbqjGT9cwdW6r2B23Udr3BQYejPvZ7CDuqEuRCRwkj
ggIRNCyI9naOXqCeYaGM/Awlsci8ybHxLt1vTtiGR3Z1MMxUxDaDarDubaVPIwbL1UqqNFu4do+U
NjXQQuPU5Z8LT82ByYEyN+nh7Q69GjI4ar3otsR7M/O0D2o1W9b8Zk7Fiv99fZMBcXArEBjMBli6
b/9gAvLGjXmlt1sbavMxWv6pTskEzNh7E6xvqNw1KC2B8moL2nY+3bCdDvpm1tyMLyslwU74Q1Kj
yzte6J11SZIrxfwfm0aX9j9UptpTDXq1qbHW5aUUXqTHy6pdzczciKWmjQuRMgfNq23T3sUeaZlJ
140w8RF1sRUbP1MzR5b+ODYXgln9VFyLOVkokAbojsGqjpHcFgdk7NLOOp35/AlD7SDf+erZ6kNl
5FcDEhnr4iptPNPMGWxOntYjjOH82AfbokLCrIwMtVNCRlvgo69+A6gzoWhsknJxgIEwqMKCxGob
kAn+Nzgq5J6lS1UcROEx7+ge+b8wsy1jWOL2BtKsG+mSNG/x1608wWsQhZvaMUlQKD7nrX3AU5FD
mgJJ3le32uvf79raPoiW/G6pQepZQbVu/dj4qFuYBFm62AyQlvsLPjVex+bRirR2j4fQd0iLBICW
4AWQa7enTyyNF9GtaYgvjMRvwdD+s0b51rfvqi+EJR5SzrWW16EUcMu6HPCjBfs+AtcqjB1Rgun/
A6kxEHbg/morcfbCgppwk3K0j7huMvJlcgvSPPIKL2e7WhboAjqrhZbJ0RQ4iNfFCWbcjRGYheGy
T1VIAhcGvz9+KQXuvr2h0TR/0EPA14QvKDs2f09oQ9ek5Om0W1S0VgqqgUbGF8boDWM7uhPQilCc
jqBVpON06bQ85Kg1gjowruFzpOvMazYvi5sLHmn2aQ+5r8PHQLwopEsBqhIDoUt7LErWR8a70Uq8
qh4tLwHLqKXSIc+3/tI5AMJFJkisXtahU7LB6z7kcPD7lMQ+ysVYkZMaRV4pu7s74IzvreYBjhIs
0y2qbUgGz7Hlj0kXZEYAodiu8Y9uwrKSqejGVoNjSQfBBcZrtotRkMTjJQF+mnTBd9X99+zdmjSP
kKgjTJ3fUrQ/56kwlKNpel4PdnDz0L7GJA5EXguQCNX79MR01zfni/DPplTsd5K4zWHq1OwbgKpP
1h4kffD/Fyc/t+P2bt+weLl3NxMrXwswM/A48AmBwLRJNJHxqdUpFiGI3zZJIqJZ89ueVLTiSK1G
xEgKldqv9J8dSCBrtxsvinc+l7ITSrLz6bPFJ+F9ynVv9Ir+Ld3AIulXVtl/3d54zsO53bbS4S91
aGsWGLGpdRd6JHA4NjPDPM8s9Ewa7SrvRrB2zH1vuscswu38gzNCmEzUaTaEgwCJ9f9MGsYKrvU7
PmCMXgy8mTpbUX3KG7nnfGU5b2zSKkIDxbJ4vuJRx33P71nTxaT8E4dsYlTx4ro96cuzAZpkHpsj
Aa8AFHGUndUo2SuQG/8Vk/ja7TYLRR/XHwiFY5x1JmcVPSm3hYdTCO9kMc5jZDcEKxOHcOlUMmht
qkRN/v/b69jyQNBetNdo6+Erdy0MPglg6aCF/wHSgo6xxzrbklDRgKFAy5KSFxKXaorR6oloN5fx
4Xnj4an7xDhP9rq+ZPLWaX9sUO3QgCCuGLnU0RMMBbXnsxLEvie+97idzyObwaIaeLtDJzXH8Kyb
xU856CxZFFmWe/CKAp3m6TNNwPuFJXLvqS2KOmb3ZR8XpFvuwlkT6JSmhrh6o1FnvK8jzKmFkCy9
C1HwDO2vnaqV6KtHE7GtXOGdbz4R04Ie7LtBxfE5AQynukbQhS0lClU2Mzh7J70uOlrNSXfV5ibe
UlwqihnQ/6mEu44XGHGtneWo2Plrcgv0a52SDisobowTpxRSrAvneF7BPyph8cHw4+2FnGDw00LS
CnMUtmLriwqn74IAvoUd0WxpS9uWhzkQlsx6ds5WUCAhn0Nvhd7mxDUcpcOa5Whm3U8x1YNuf9IM
T9Gm9qyUAH5GhQN4YlZl0T7OY9E8NHxXj6epVCcq6q5FFJl24vbBNlfCPrdyTq/2rOl9qFcOm+PQ
UQi1W1zv73IH83W7oPKTLcPhCwRUOMZxfrGMM0xwSLpW7gP0nxj2PL7/lQe6aGjH3xdHkAbmzwlh
GNb6s/PukcDmP3fenWdDr+/BblArHX3zhx/iKSR5UVbUO1Nt2ve6VSoSzshOsMUW3iImAdZ2XsN8
Nx5EUjRfPubV2PLhBhV7Re74Oqf0Toz3AzgqiB8JEBb7uMM2yZxfaSSMafTfFJIaKpq2c8e1t591
rBikXjGQ2rDj/l+1FHF4s7xVBh7vzz4eoU7jADCLvj9dU598Pg7aukb5rUsSf+K2D+UFjF7BRMnV
QPxQ9M9qiyk+CqEqFNebjOmBmB+DpLLmmW1KdmMuMp4g2RN91QFyfyvW4AgsYR8zPCsYI4B3SH1u
9gjQnS/HO5LbdW7ib6vHgJVIg3+Jv3DU8sCRmNPIEMI2yB5DYCt+2bhSMwx18aluv+NufZwfNECB
mAJ1ijJl8TKvBXp8F0E0xV/morVMlVI5UKWRtjXoL/8WeFUAurlb9N/un4EsioiboGTdvMWuaTrw
DQjyeHNlq9rlQtmMT8xuLr5kjlvVjlDQZBKsU3+8T7zQlWg0K1AsIDUq1PcYVLgl2fzCk3DOsdOM
W2GmIHdt0usIBeH+9du9r7/tKNJQ/udIJ1HGoAPP9S2L4od6snfQjEfuP/rPVN8wlEOzxP/YgG8C
NAzcOlDmmsDPt5pQaKQonBmuPkt6fLZAoBXzsfR3VN2KikHJv+kBdNuTso9Y0Eb++Ni5f+RbgWRP
KYQ+OgKmIuFUldvLfjrcYicAv23p4aalIbuPsnla5wIAH8sazSHQihRsEDCn73SsNN7uAzkDw0IY
dLpkB8hCQ9+/chTakVVsQ+fc7qi+XHL738W9piLMLRZKJhmCGPkzdlb6isTY+XoG8RVcmyyf0g2l
gI47ONXrvxyuyzurwdYkZOrDcNy/cBZHp47/6/5OqXdoAhDKy4oKbOA21VCgSjqh67rdIfYa80gd
fIwSb//JYNFlVhGLdrKs8RclDqakAuhBBFFgSvKwX20/bfv4txQ3h/7Tzuip6yUorYmfrdwhqLHw
46z5IjPsbOHb8zsMIa6j4YwmHcJ6i2IYNKD2TOmCuyLUbb60X60zCApVGnIxdUQOuZDw8O0VpmZN
umxHc5ms4b5/u+dvfkOlBhPHlc8F7rOwXGW2qTam42TBODYgYSqB6MxRh9MXeFKlDY/pCQJmyUv1
+RbYuT9n1OeaREMWWCojEx+iFuivkAjhp1oqRVmgzfhMVUMkdiEIIjq8lEYVQMPOwlQKXu4DSnVw
RO419gE2WJLnhQcb9/dY+1aQcoMqFQR7/hDpboj/chymNarkB8Cynbs4MJN68OT4E+R+K6ipCW0i
TpGCCiV1m9rdNBGJ1iM1gQ/YjxiWKMdfPzzQTrIpdynJfQ5pGcwZlH5Cjg4ydmDUZg50EBwhDUN7
1X21XZx9Xw5qu63wk/5ErLYWkRKb9pYlag/4Y3RNHUIiRxPf2ShWCMJimpaWxcIK+URFNacxFmxt
75j39bNffdxQSiOuN0B+rJwy/KJbzqO7PPBAGNZ++dwwv+4zXxeHqKWqQ+PE24hAzU+mERd5OHXD
GaJy9I/x405owNs5Zgdn5cSBm46GFanVsuv96slbNnL5369/hE+EDV+jDsvGlsExhiUD6dRwXjCl
xif1MIdi/rmE6835hzq9gpIsvVLxqRJvyeuC9WEw2OhCuRQQuj/SF7F6oEYt9cDsLqvosiZwE7qe
YHYRv+XII6HC/Js5lYPBtQ4XyLYCYRybetOzw4VebBoyZewaW2icaErGsIfMmbe4aM5svdUupci9
SakvEFgnP1Y7P5+lgrasdjMtvH7LhMjuDumNEAHaz9EpKsQI61arI+SqTEs6q0EgUzkWeXW1RkAr
Hsi2suAMC5Tw23qwQ6M8pD8t2jEDtMbNlQzbwqGDDK9OVzQyWneVkGlUomVTbqvVQ+7cjiMdozD2
IpbGWB5NqOjQ7r5KC/RR+GwEnxTlb3QLJ6SAb4q6BEdTSner8fBB7zvSkH1kef/wpRKc/SOcBPCV
ywr2JIZyrdXNcDCb4z6ygn+cNjJpaq5T7vClLtK6HE79V9t/u3wwKTPt8en8QMKe69b3v3rpCYxo
ALaqsQl1jpgInTMNfD5VVmeG/bYv3Y79Hqj64s+7OnfJSm0X7eGUlgxbhy9jykxBga8CEhVLh+TN
grn5FoxMcrU0uu0CH7FTbjB8mSEx4fD+9SgTEPR9ZGXPjF6zUUXXif3jA3rtCwhyZ5xldvC9mZo5
z5J+B0+/NgloWUA2fTjp83t7Ff9Yr7AQzkwFzoL2fwzzKBu6ERjFVjaMdJ7xBkNcf9Vhb2ic0vH1
mJHSdZeq9OrVI3Qaq+wsD+qWOswHiQuMHwJ8Es4iiLt5CL7elGdMQOElv2hyOiQQaLrXZrTStyda
rcxleZOIB16aM5GNUZOfnTZVxjfx0U2Le1eLVdDvhKj0xxYRLvI5QqsiSZBKJPRDoxbTEaGbCWQK
2eZFEXY8chZ7V7rAz9gLqthAcxibmJmsMDFwBVUWbWoSmVy+rACqMdPuzWZckksH92lJaPyr43dn
3elez6NDIqGnrW5mFDJpSUKyBFhx1DJsdLgLwEwRFDNpUNYFjtg7cQAGQB+UQYE3a5pPM/8ubWmF
MD7tmYp7uf+N6gfTvw2+sTpdUruX338DaoJ0uOpDDE4zhM6FPnx7TogacdlaQehO9SSLOypGAfoq
1NiZ700Jc0t+OIyPE8l51pEQkxiKy7PnUdj5mmWZKXF7mc4rr7T2ZIYrDPnkI5Ms73YPbd87TAg3
tKS0Xs878J5Da5uDv5I/qk60Qo6NF7XRpAuyaSGLqQNtjMpCVbWm4KAi85fqLWapPSZnBhN3cbXz
R1mVmbTz+PUTNUfy+ln51Z727VCPmFI8cGVFX/me56qvrVk1GENfbqjdA7csUr1jyaBLkpqH79de
mJz7SaFDmtlmJJsLLAYYxQgrMBykkad/KLAPQovFUIJpqWLKcpVP4YhCZyescwM7mO/p/pe4xVJZ
UAqq1RyZIcV2oMWgEecvMw7NPj7/Qqm9U88YNb/J9i6WF9nbolmvPUUvAZVKVmJc/xlO2bjzrY/u
vKD/hxyvlr3X9e2eeEeNR/scQwnmuRWS0DbNUSPGHyqmPKwopAzOThq143hUAU1r0HYjkE6wHHrz
i9rENLR0fyraWr0GAMmWNhLKxE+rdR6e8bpn26ePBdMR5gkMvuhyX2FP494pkdvu+cV27J2S3c8j
z/GuxMTD+WIvexuLPAX/hLWrua1xlswhA0RvzPuh4/FbV9UTdkOjRR4eXUZRBZpG7prP859qqGq3
62jzSWGpXleBcFrZDUiODu/gbk9P9+mQcWyO20Exa1iwlZJYGbaEuX7BAJmv0L61UPKkdgyv0ZRR
5HN7va4+LpsAN6eTJ4RMeoiWm5+koEsK8MRbh8SE8/W2+yklOpEWAcWm85dHdGfVeHHF/X3ito59
uNNgir+U5CNaAio6B1dohQjKSzsgojs+rzzWfr4c3XoeDKDkCfzUIQjCI9GC8R+B4Vdr1OJ0fS77
XdD88BjADwkqUEwtYBT0e1nqc7MDzluttAK8SwxRU95lnSRfaKfTW469XQM1SsX4zWpoIcpJVys5
2A3KwyXEtS5LSR3Q+TixoTp5Rymp9R598+UaKuisdyeSpgRtpqGH+SGt/k3BfsK4ZTsn8+CIzYOZ
er2NFOxK75vRmxnFhK36HE0pbd6BRw0NqVA9wgp/Y51wzygQkNBIpvCc9Z0/IT8Mj0OO8lUWbBVP
VvcarGgT1aIn2JYTUUrvAH/Ela1jxRMxLPyu1y2KI8pvcCbuBH1uTAuKQ/wBARdaN8sNs+XFGEYM
T9JtMEVcGlSbOiTRsW38lGTijPNPIVD2Mgk90D2B/qqEVeikTKc3icBnmbNRNVPBDT21KTcQ8gbt
13B7SlPoIdAeN/cPm42QlQZmwjkIRdBB/An/7D8Cq7mAs5ZmP6urtE2+oqUbXkmsNi8w0NIuHhaP
F9ldT9DaoAczxehsGmVJBVCtCWGAsVDBPPO1Glt5p5Omq7LUVzeC7AXnPujgxbePmX8DnPpStJcA
S5UN5xO3+LgAbRtUbvvFJLwbUzClPaeAoZrk0SAXxUWEpR6eEmXyVvcG4+4OajxPtXMcAnQhvatS
+Eu5EPmTEXlJ6+jfYuaRC/4XNk0C3Gw6gJDlBKU+8fJGg/ege2Qos3FudzEWUGrbJzF19FjR4hRg
5sLj/pGxOvZwh3L1ENhy1w0hRVvdFGxdeaL7+cM0niRhi5V0SEwhV1HC5Lw2WMtitd5ZJFC3lP6c
mi8vl+d1iFGMwzTFQaPTKTsx5PtFXu0019rFbjjfuv4XzBZSjw/WQU54ZZGKLn+qolmo4BnH+jQI
j6zgUCmIdjI4lBrua1Th7mTH+L2jx8xVrmachqpLbWc3zhXUO1ffv97ufyJhicRo5OwpwUcUGHeX
uJMhiqtjVeLgcp+HfrG9dMM9EzquNgxk6LPLrWfc7uvolkazag9fVi9Pslxr4yftCYz/hzV2uVfx
UuYH5vbOP45IYztonUhI0KXy5C/ie/t7c75g9FsGbKtO3JfXxuElB8Pbi143xUd4R98gXYYQPIGr
w3KGVBOF1LxyhXaYk+dFf1EOf0LIUGajK+ihy4U214qMAOUT/V4s2nOL/4n6dipv1cmEMZEIwtvr
/Ka3+aWvPiqJmp8jNfKtgnFbbyhZuH/ydR4H7Xbl6l8+nEv/dd+mTZJQBXkCzEM1p1kbYcvB2rSQ
38hpgkl6kDVrM1IYeb+8uOrnzmpIFFc+LKFW0AmtCnUM/SMYPTL7SbDxZwPJiPDKf3QAPgTwVCqm
otFv+RdW33MgnQEDt9aXGk2vHDOp6/EMhsnklciHwL8c/1QmzwTwgcMSYSyVOu5qF9vTeHXgwoMF
S8blrZQTD9gmmMRWOmYNzwyYz2dfD5kDvAVq2TVIgm3ys8N5YVT+yKCWQRqCkEJFMa2eb8CHszlF
qqv2dkk/qD/IkqjmQgYl5Q4kN6ONVTJpC7WlY6hGuYz2C0E7s3XwwbJLAUr2W91w3x5xqHHJfFsh
nvIFjcmYBSjmrChtYxnyKyDQ35A6rMziOIf+z0zSUJxAiOFJWbR6O4h8TpJTpVJbNueOJUrmaMxE
f3ypUYdK99J79r2KrDkX53ZdJJ84+z/m6XlPzNPNPnmQr3EJ3LF0ZctexjAUt1C+cXSn7oiz0aST
wYS6+pjuQJdSwbyhyvRbaFjviRRpkNYDCDhyMYw7/ugxa0Yvi/zk21GDZS2sbQKP7X0rIcjsQzzK
KS1L2CyJcgQFA3+LbRlBiYRMb49DvOxgQtFTKa9ob+T/VlyB/lsxLHjeaMEG388GYZnI/QrA6W62
UDObRWTFTZnnnczsQfxda7iMcWQMuV5Xls2RbmS0Prnih+n8dMjlAeTrsn2W3EyencD/nFKKuMZP
lcp7+U7MC8nekOKag4jGPddpZk1438ajDTL2c4GETKHAnXeyKHpWG9p3Og+hb+ZnL1ChqlnzyVtd
WWzzUaDh7x123OohHJWGCU9xYzlrvr2z0kRdZ2fY0gOIckyODvfv1mvoCoMe/5AfzSxiJdr7Ygxw
gYOswUpVDtp3JtQ5dg3orwLl3GRJE5i/wdSHfB5MQYz0FD6sJD6M/TwAjKqa8O0zl8G1SpLbm1aM
FcJ80MMkrR2XjiBcyKvijoFcAiLw6h+9ChBQaThLcM9RpYF6p454a9Ze4K7HJviJ1YorMkJ+YIpt
yc6+9Y/dIbK7gAS0Z11wL6A3i+JoXQvqEaWdpq3rDiG74PkfKNMW6jseBrW09YYGJi4bmsE3vpOh
IHZkVZn2QNZZ5lDG4uvFxIoBauJJkyat/pYxzXZCZcgNdQFDDQny2qA8BYfXjUM68r31B1EmZgSC
9sZT94HavI/j+3fqT1EQNI7ABXAhezZmc+fcUz9r0JKi/YyIHtNiLx/Na6cvb1gOvMU5lSUYZuR0
Y5u281sx1vHXWJBY1c0hxjTgHDJSspscfDFgOTdbXDKZtk0zn5p/bqbbE+LZWHTde+y3in7kiuKF
g8fnh1t5xUohH9lOnM7eIZ8Af9GfZUEEuGu6fDkX3Mar5YG2dfSVXzB4IuXGADO/uwaLwuF5u0Ab
IA+IMHyxt9U9Ype7tLrDrHtTsqwYkjtQxMMCRJzzvXB2aqLJlT4Bs98UYJDWa5CQ+px3myVlBuGE
htkRJO1v+mEXr7ipZTD7c1ymSfNaKFEsfRsO39y1fGHNBweilzpua8re6m5OLnvOjQvdYZJNNIi5
HuldcKWWog7ZcTC381u8GVa/uGj4dxoqnwjLzdWfufCJXSwVTcWL024PWUdRaTkt9ZtoT73DZFlm
WRWd1wLQHp/t+Q/+zgc0Z0kqgxald/8FFb8arXXP4WXP8gY1fE4ZtlRi7QHWoSYFuoawJ7Z2TWfY
TcwLOcnQP0ACFSNusizG3xoLPotf9LFCxDlNJmBQnf27FZpiIs3vsuCR0PjW8vdpyKp/G/OQB499
AfmoKMCm7hZPLpJbk6Si9jz3zsQYntrJyQA97z9SvzNhbdhGYtx28bNRUg4SjzqfMLgrBt4O9xLD
po6y4zODrATbukzfOTD3rtxpuQ7VRvO1W7jqAriqUATQ5itP6XNZlO2oMiTivXBVzsHoZ596U/CG
UmVLXTFKtfIQKl7uOoSyjwU0rnGhYM0h0WZ2cb7czLWtym0+MJF+kVRChy+WjgOflZ/PlN+S4djC
1lwL/UzOV4nhHhXkB5qo1wbetIdFlXgd2+ruV6YvYypkF0g9SeM6lD3XfbNyu0npvS0m8ZWmhSQI
UU/s3zuytk/GkCxWnM2hIrY+yXNN284iPG4/2mCLCN9fpH7nAc/RMHzoYa2BDfhhcNNN+s3QZxBK
ePi2xr0KIJyYDSTFnOJDZVDqGxPbjC7lKQH/yY9bC9eOLXIrVyrEyxEYbyLUVavAIKCLkivpJQPk
KhWKVuoAld+RFtwF53pYhtfi6o0EiZqSorJ4qpK7cPlzrMJKP+b9ZYEWrAzpguCsupd+v52ZDhem
sLQWNmv+FPzVQcSMxF0AJb75n2s22d74xbE34M8wR3nVd+VehS4KcB4zWW8rGG1AmfdrrzKCEPOw
nCPlhs2VZhn4mZakBApLvDC0gMEHhAskKwqciAdpXwFC/A5h3F6W3mdVR1sxhPDXAWKxdWNVGBeS
lgoSv0Iqs80x/9wE4EW3Js3Oy1fYdQtH500KGlCdwTiJIuuppg60DM6dzxQ3nqiVByum87s5id8j
utsjREy+JsmeeGT/kDW5AlSO7oUqL20irFb3VHWVl7qQdW++wL7G0rlbSy9/EWO1td6pF0T1z/rV
lc/Lc1eAVZJpQo7oASqYpN1UjQ6yH5mV80bNdW+8OvUrrj8cDx2HA4P6SWLEY2VmBhpeBV+QyurB
/jniafVBPimhg9kCRpC4nNZOvDoxB1fNOM12JLaW0+mybzkSoIMbbu36Rj7Q0y8io5/pNHWM3EeL
UyJ6iF86hUzh3/FCOvU1dmUQTly/fVAJhysAG/w7V54qIsvxGBex+73ub3QI3sfAu9ptAgmh314O
O/eYLYoNyxYbOZM/NKrSDw9DXzTNqpKAn7jsRHqMD1NLz9jAekvH6zAhtfo9+9cDixlSNdDMT6Cy
HfJB59cOwjRCVJEfbSbqcVnBR+UauwnL5pgb7eqH2eQa7Yt9CLrIuHXuh1udP6YZ2ySFZ1o8Y9y9
grmxbHFFgzBkWEXwUqJ5GGncmK1af4tMfoAscSoXfnLiRaYzbjAjUcbBXqbLcl7KrlJuHmRg1Jbe
KreoroCxfjyPmmqaMwFJYuj+WMyHygi/734fYjIKdnG1UCenax0PlvSFjR2eRdrsIyTXkRpznkJK
hnf7F2JhtTHwrNnE2kywbKRuBnH2YV1LJLmOn0mJx2AJBUEuQwM3PjoX8ZhysogvKofIdsansH1B
GfZUfo8zyyEO5CWxbQSXWGWxhm4fKXIF70wuZdeCwMTgWhb5lbOmQtDH7jP7RTH+lunG2zri2JhM
XtQ7NBIzH5nQn4vlL0xq5pgPJrH/7bnlFaAHZmUTBKGSL81qbW4neMppRWtnvjfeIP0CWXaAMKrL
p7GlxpA7CAR8Moa48FGvUMHJg+4ZqqTHcbV0hpHhVaKFRW8s1f8A8BEm1X9COzNkJ5fdmS1BtwVG
j2ZeT6H7gncwwtIOUwyFZ/7PA+xqQjTiD7vlE618EQITbZPop0O6baJEVtmwj/4FfKLZjFYJK4W3
RdjSfDDytPUQDJmkT4tiXBqNfO4fGBfGiMNLSxOIySczEA4AZPFROiatan86nF67aP3R+bSwJEdy
xEhdb92CnE2Gt2uLSYBPE6+3GuSR3f1iDvQ9hULNObet1D/Yv9RuIbvcZOFfpOYxhdK6CMVz8lSe
3gh9UlHozh08Ux2azPbsjHkOzL4jsqNmGFm44eZ1PQ0HRKHsuGqKbdYRlUfOkp8vsprJdcl6lJaf
ighxWDJZO1n7ZdiONsreb163ltuVnBRty7nlGyzHzQbpSWA8Ep4TFHgbrmktPh1gHyIMyMA8KDR3
JXXhew/CFv/n3+Z4nnA+gJLh0/fb5AGNpDtR6vxkR1aw3wqSeOGoZOWNq9Uk2/f/Qvf0C/ushX1b
tj5JEvez82rUjQxcWXDyjq/NWybiBZ2INLqdDcBiO85UQHCyk3bSzhOHtHR+jqePhPlLI/8cVT93
Kh+AMFj+iK+M8Wgf1giS6UN2if8NPK5L56aMPXe7ctikxKBY9hAqe4DaFYabb589oMBlV5xy9Y1d
FxCIIqSYbEtw7ZUAr8+y63UTFogNP2EnVwgVH6m6iy9m3aOgAusEt0T+SrV6+Wm+NF1VPibp88hs
XfjJO+HwBkIdMNIwR48IF7Q3n+Ey71J3g+8wV5kU9zd286iUApdQQE93sA79ll28O6BEit3/FPTu
U7xZMlOV6g3tj7/rCroiP7HBcffg8uW9du96nO0nAzS1q2QYm/+uMibsmW2dx788Q/THACGfof7o
P4fo60r87T0sdhmkB/WOBhsjHoDgcPEJ87HO5ZPTcbRzwLYqvkrEwVBG7dgIIZa26tHlgtlrkNRO
CaVuCP2J0v/xbUV/+nyHwXDcKStwHJ+kuK4vsYtukhTidSt4MCGAbN2jo0/WXM44kig+ZqbhB8f3
5vfTNwqS7fsWJXpvE6PDRO0pfY/4IW95r6VRL+giT1tZ987be+wg9WCV+zGhmFtfkwbF6hequ5le
JT+2qSNTK1TrcPnYOZr3FzO40r7/hsVzamAYyIf8H+4ORG9L5ghn5IR+hRZn/thFMeHoqXEvxWde
aXbuIyZkTG7XgFpvFCJ82DywYm8Y0K5pjjlPxHffKN1Drftfm+wSYx7Nc50B5AoGNhmeOnbJg13Z
wLeTR89bsJE47KXlvLtWW+U3R0BhWn0XBnp6qgmBRNo3rBIjHwqm9Jvl2wlYvaaR+PtRzBMnVBGq
/I0+5dMCqruAZyMu46MNOjsW6KcpCVrsBaqHMbpXS0UQXzDZXF9yeOTQ82wim/6VO3FTDmCa6V2e
hJrjMUQy0pHKxXg39DEGUlm94IISy90MHdkR8T8Vd1uuGFaGSY3+cv4p5YrAYNO1v+ZhKxzn6jHu
8oHF9zDGmOoivRDasY+W/eIRmDUhyfuMh8g0eUmSOREXyOERclzCR4ENqxD1I9YbGcovkkAPqVpf
uRtLvpoS51U9CSIhkLg9uX99xy8RjArrUdOaNsgiUHKAQQFhWB8UFPVEidncEPQs88KbOMQB4+76
nhxFfZyTlKoyRYuZBfi1mUgCyQ032VQf6mzginhzdceYP1cucv98SC9dUDaQEiY8QCEIp4HikucE
u55AObjlO/LUEdmJKZCYlLCx0gZh36zEsU6yoMR3MwKWV8wS1Xx9TLw4KhWj0p5NNM69whHtTLUu
jL04RtJwscMTeJjgwWqAPKdWr+io65wzeJb6DwHxZKBXZaD+GU27gZc6b/HHXWJ70L9iHmanhQ8+
iPCkWkpBM6J50qE3erVLfJsbQFScDrht88y4BKgTAatG8wpHgsZGNBmhL0EAGATg7eJX5TOdOMeX
n2BouQJemY6exIq/P1TAavO4WjJvL8nKzS+jXgnEcs0Yg28QKXlDYz28DTFsWGiSyDTqtaR6rFVo
PFNZXgVAzOa8ZpzDnieKGjQqoB0roZAf4Yp5+HxwmT9kFKdpxADpRhrj3j0rHtmUKXPkpx+7a25w
66TZp/jrWSRoZTiiZzVgJG6uXjcinXKnB51CskbHGnP3a1qcVcmjZ2Rsn8OJKKnHWIPGEMccc7v/
QWr/q5wfq7sFWA58BY5XTcLEJZA9KaTamtdT3tsOHNDhmgxxpAYzm64SdRjF33CVtMb0wnCKUt5E
9ThR7OT2QBHm+lnV2e4Ucgcq9ja2FpUmHm19LuwyIHKkd4G6UkP4BlCdVVL9rrcQ62YyQBph5CF6
VHKNL34urK0ZCoWXIy684Cd3n6vOil5/57HqfE3TlN5DC8QSI9m80jZ2NEixhMtvG1Ga/XfpJ4rq
y4TnyychtaJAdo49dgplut9wMOVsJ0Xnn86r72N79rt6/0d2OyJ34Ne7xgqwSOfbd8sxwuS83PnL
whP3KV2lsjOGI4fXDu15bOlu0YztfSzAYaSyQajZOuDnoNYAL5hcpbbWLmY38Cy2QAuI2gKZHhpC
m/tVEi9K8mE/TEzBdTiJ6rHCJK6SNHzS07ORe/netW3j78IaxLmzIL+SPPm/lJxcJZ1OKdOz62wO
dScbbsn/luCih1xbUL0IFy+AgLw4qAn1WxL9ZLzMHEpi7EA6jEs3628Z7wV5cpL/rM4mA8FQyAX7
u1vWvKfd/WjrBp4A0jZePS5pTKG3nYqgmZbnLP9UkpvIQZFjhnUsRgWbeV/CzHpAmer/jes81YWt
DLTXpFe0VYAqeOdus16slrUAKgHFz2SdpxzVuwcnV0Ee3Jra8SdYZhcXIfDGn9HjKZHfkv6sKBbh
VjaRLjtWOOnWF55+DH4TqVqp9NcXtEKM+QhdZ42qLZ9Ya9sqVxW15nnrixGqGep7C7UnAXC7W3GP
1gzqio3GPbmj6hfuJMTiAl9f+zZ8n75ejHG/0cfqM+skpOLQvAgs9OCV07yI09xI1ZcDAf+4OKyB
FNTQEe+I8n/Mu2EC6Kzun8c+AzEspKHbB3B+Pm+HCN3p1XXACdJ0RyLGLkoOT6qRkJ8akN5wIIhA
r+J0uOQir5KscaFapIyL4QrsO3KygAmflm3mIfm9LbzCxItlGzs9ImFi9KlIhJmgmv8+CSrDhOL7
HnLemRIPZCI2bJh/xwsC7L/d8NOw51rTqP/oMozvWaoc/0kAaWmDYGtUy1fmVUETJdme6VA8H/No
04r7eD5GObofaxOIs9rpUhE4omg7NUe412S7jmDG1zpTaONVCE7hT3gUdMJ055qBm0pBFd1m2Csf
GJMcDBRAS5YQOCuanZKfJadriR3LHkyLkDVaVlOoWSzyOfc8zDj6qASAsi8p3RqcrcnAFB4E3FZn
odAy41gX0Cm6b9C81pHsrZcrG/4Bfnwqm5ofMPk4ujZf4xw4mV2dVGTlMYasDfI8G+lLt7IlXcc4
a5cqxRH4idLKXDNp7qXowIhz5lNUYZGV+nIKiFyV9+B5dx6kSRpHLGp6do9CA2RMeLceCrXi//yB
BGxFzc+xdQrBHeRZD9UAjininIuZ9MQqn5qYqdugt/yiQX50wuJ5HolqyMNsA5djrwfUYtQ86HQv
s3iArtTZQBcDevDGObk4zsJIfJUaVFvLXztCKCx9zTUR/HEWvwh3ykRQwzZItFHTxPoUucvb+OzZ
udoxNBsVL3LylRnLX0gBi63wE4H9Esh/MIw6Xn3ClGgQZ97Kyw32Sc87eIN1WHaFbcKNJB4PHFFJ
FHh6SahM/S+rBNE0U0lYRCkbJJkUKftUcYStTPss4RhyWLyWj6r6QB6vIRr+BqfwBCkljswIpcVl
dWAsX6591Emq812sP4eaM4B57koU6lS0EEWTJ1R6hJ839s7MLhwtp9ZaEa+OysbL5XR4RpK9AVWI
OP75RY4waxN0q1BDM+r/vsoMFQDxJQSZfyw4m1oTtY8+1Crl+cXa5o1jIdhQF94nxuyw+QEQXo8I
gbls3K1vFKmgNt7iYcA2Z+vw8s9LUioTII88FJ1Bt2PxaFOAKZrNlbzp69YnsoKVrszip/fOHOoC
7oBim7bvxDh+OpAA7FUoGEjs+dzw98SQ7/IuLXzM+2XIpQ6kvSE0dqwZ0FBZe4GgFMt+1Q/rYuUZ
1FnCzhuNwvPaK0CqcEhm4CVdumpoQ5Yykk3PoKPpo9bmmY7sQv1GMAxLdUHQ+ALF0rsePTdHju5K
uVxDX9NHSnc2gUmxIii6falWuTR9zy4Qkq+vpsc28+ZbwzdIoRRktCEt4aJmVzKrZTcpYxJWwZd2
lKiiRNbx5v2625lFt4bf64p+MxQN+C9L8AXOQ1lIlqrNggfjWNkqnpxepLS9aSsL44qLSN1dEor+
k0nRr0nQrSJnuQ9a9plg/SbnF+oRedDA5j4XPqBxlfl76czAAaOA2az04MlTxCFZyg3AzzA8C1xU
ZZzFJa1PlfUB7zIjz+rcS6CGM/FCi0wI15A/MtbIxzGChf9bKQjVgjFbhjFz7BKgIXGk3SbMijqf
j6un79p3w45LWjKVbTDNHWPoZLuooWJcBS382GvI2yvWhtLWxtxlKsTFlNMQ0Tzse8RPtSwAS8HI
tDPw4yXEGpDYhKu/kaP4qGw4jYBMeQcwjlREcRwVD5kFzSfhEGAHzIvLyyilL593Dikk/eoqlEC3
JISXB185mkfpqK5UJXPM2t+u05KSdYZt4s7rn2MhWy7BABSDbhAvvnZASCMbB090DP1kLglFIhlY
4LsoC7Y64xrDI3/hnu7yQvIH9QNRXQf6lb4MiNwxglQkM+FvtAjAiXmHaCfWz9MKJwv8eUm5EVwm
3WVM3ONH/ssl4lw0diRz+vOF6hRpT6A1I+xxssiaFhgoiggOuDg96NDWxR+DXcC9eUatC9GepYmp
1LQX+vJecy09W8s3ly9VIrZ1An8DG8upVRGUnQGMx957DM1x1c1gfS46Ajx+FOBgHWu5gpBcBXs6
mvP2xMdElMJQXOj1KSW/DdHgpN1g21xo+2suOOP6MhjXD63L3NGotg4Ev3fA45UdUay4RQmg3ctm
2e7C6O2iozkoRNjyrsDQnudnRTgx+qJoG59T8fi3ZschSnt40ftSxrJC1V0IpXH2jkIXo0r0WVaa
7BtvMAPMWywA6qZygWBGI7hWXNxXq49jyUWWcxn5UXl5iCxEM70JBT4p9eDxuU8YW0PWVfz9VbRU
fb2UhJEXOl7TadMCS1/sxkC1j9t/2PnM6F0hXOUdZFweYkmWBnpmvWvaoU9FGPUTcBAlOpJyrfgP
nyWdS/Sr6cSupm87F3A+EFe5axTgOl9+i0heCn6y+pE1sUqvhOEFTdf+Ep4MQdUuJNi+A+fvREon
uWrPDnpWd2nnFqPOu+sFlYeMCG7RI8CSA30oupMwfpWJ/VC+dtyzyKfSIx9hO5S8O5geIypYWHxY
zMjXnSoo2iihlB+kEVZsmFHz30+xkSpoVqScu+dypzRLksD+cy0DCHvqTFDTGjb/AiAODLxKPgr/
bnxuVSsdMbcAyx2CcVfLp6MQHwdlJJVL0szEoC66QejtuEM8PXXPIjZex1aEDiNlGsahXPeSzCva
wQj393o87VGOb1nsE/rX8BJ543rqoXOBLDxr7HPbtRQZm1HqFXoIZDm+vtutgIqZG7rPOVpS42w2
+eO0m64bCfT3sGFu9kkw2vm9bC3/NylGnKPQBra5gjxsbwTQ7zt8sHzHEJBA8wRuAJaxL45U2BHm
MfhiWoT8ME7+1w3dnHsy8MVnESsdpRmbQsDOGUyhu0rORxRPk2kHrdyeXXDJcWhi7av/ODVTXLRu
K8AjZPHDlyBMDBYnHgiFqtnTrME82o1aAqSJFo7fKHABDh7sspagyzuXPMKaGo8SdgI2u6QSY9PR
z/Y/UKJqo6SLHG4N/CIQ42NbliuZzsU29c8cWYMBwlN70mUbJNn8MapH6i4TGN+G/VjEgWL2wqzR
Cqz9xu/zfxy0OHbWwvQKwZbOaisVq/hhMFkeYb7jCVYVKVb36N2FzuzHm0A5Akl0OnmJ9XENxGVB
TuRV06HO+54XpbC68eh7PPh8W4rK6ijx9xwW5/9/kaYfb0z7syWF8cWyIlvYXCLqLbbqdY3cwnye
G7+7ZmZ2DTW0KvClZC2lV+/5QPttjjHeK6JKb6sfil46S7Q8ISlEJzhr59dER0ug+q7dMREnc8t6
A3bkkRAIH6EDs1VArk8709L0FZm3M4t6UA21joacC7SPE3Ss7vMd7Yb5EZlgJb05KurVK5tWz67G
269mkmmIQ+tgtK4TulLNWF2ONK15HwkGa3DnrvnPFgN1ykvnQl1cBf/xWjpIMmLOsmLsRmtSmAwg
/XKovUgUqTdeyWY4ASPmjKwAoSFSBbFJP9WE9PtK4HlwCaGsN2XNG0eIbX5a8buT1FPjp3l5AR0J
HXyH03oaTcz1Bd9b2Jjku+Lm3H6Mv594pta61aCLio2CkZO/brd1Z8Y0SkyrximIioadYQaqjdZh
jCfAOUQAfKW3CZSSWu67/Hi3p3B0ovEKVx+49y0RK6JE2cXpp8DVLS/PfG27PYmlCG7cAxRsJr9v
Z4teUfgV7BK5zpqSy3kCjrT0ye6N+7e8mELeuNkmCk1YvZzW7f77I1/mUeGJ23097BldBUt9Kevg
t7c/a7H8OqguEHEFoB4z+XqkrPMUCmF/C22nAHYzRqf1iRFImQgZJGjgPKsynbMdHm8C2gmKqJQP
bIBZjWwF7ctkR1iiNk57/NQ6BIPC3ydRuJk/vNx0OeeVjnrH/LxCcT0x9PD8iU1fc0kmQSSF/P9g
CVstYyqTb+K10LAlGWUzK4OM7wNulKmyuU2x66G70yRqSV0lzJVrjqnWo7Wd5q103xCcA1t6Tb9w
zmYvXsFmoD4ldHYUQvTfig3WDgz4OQ7zXArBop2aFkFGKPmPk/IQRsiKf3OFDZ2t5giOOJyQijua
P8u7kK86IH5CKtcEZl8pUw60azy3M0HxAPh02PO+Qq5ipE5M1z5V922s9aBUoMiI2THVyJdjmGFG
wLgrTh12PisT/m0IPpAoKin6Lb46+LLec0tnWBgbbOMJTjnWGjrvX9fxw4lCF1y2IGCfzovD5o8k
RNz3BlLSb9sy9kr7VqEd24etF8t+z/tv1Gs7LxFxkrCkQp5g/BlArGnG+fWVHr49oemGs9dr43mq
3eHwpAEhRY42zpuW1NlEdP9NQDfHtSYcLit5WaJWdE7TBwwX5M7ErP9g2keTauI+7DZ0FhWFJ2fo
Qvv6igp5YjKbHeXhmeMBjYOcjBqtRZn+MUW/eQ71U1YXptBJDeTVeMrLWhdnfdtG6xDhKdXH4mS3
E6eWdHf4nFatjzA34xZKBhTNf+cT3Xaj4Vlv3RkyrAS+omrPcJWhxSrL56s7V2IKmgA8DavhXTbm
Jx6EgUoSKoRjP87hIZY4vlGasgkKo3lKUElyxF6KRZ0XG8T+H5sRVwmiMZBUKtGlalvDiH9kccXg
FnRXmtjMfGixjnLRH5KZeqnuvYX3zaIA+OiWnp10h4ayOdxs2Oa0sfeOJd/HAmherzAhm4RMzaim
bTUxXsVJ/SS/Z/XNmluFyUEgw8+SKhF4ZGwwGirGDxeT+9EABkLQ+QFvgMR6B8u2y/sYdLJrJwdn
yYZo6kr49OeNr+pHKsH1hsJUjQxVb1i4Bk3FJ/B0nJoyWI8BpXCue9ZK957J7ZYv1rr+55Hymu/G
W8/7AbWWMPUQUMq0c6y034NTKCelkWPS8FpuwBBiQtxS+5LYY/kT8SHw2RANQ22J4LQqCpOkZSyZ
Xuahknj2E6DDF79hdLY5WEUZDCCngZFyv8l39j2TxNVJpRsyWL1NG/jlDQ56ofVGf+tud7sgRLhA
i2HfZMLd2FrZ0jk2LCotN8YLlTpGwR1wns0knhgJj3+qwlGNiyeIakdp/xpdtTFepJ50mAkEncOV
o8qJfgD2BNbqCylLiJzsYLUXo5fRYAXvABvhUnhbzqvCtzHOmtW7L46TbMccTG8rzP+GndnA0/7g
R5IjZKElwCYvw0X3m3jwZCFI0Ehbcgpy2jhE+A2Q44Fzoehmzj224OYZROo4sojLeNBM6cMrwNOH
N1KAvut1piJho33Pil0jhThSAhFCOcLE6QwbJZnSLiCymkyPFxxjNGMaZL3kMLF1ygT46zVz3oXQ
7XHo2qemrKUyopDSUfo5UNpqiovxKTc5hC9mPZTq3YQTgnppGyE48XFHTvaD2jt2Bb1jA0PiGort
MlUCiH2ozPs0pcaD3CX/jLiH14E3xIt1KADFQIoPEtzjoKl8T3x5loEt6EBhjTUo27/R5gqCTjhW
s3y6yPx5a12IKT9rONS/Dxl5NPdDAsAoYhvD3FBiX1Epw+zCXgLnBs/UMaY4f43QlxWwVsZlA3jI
JnzTTHAmDSulukCrWkTqspPAFR7/0RifCJxZ8HmwLDoTmxqsM3wUXBDE465je5LmdjbcIgzA5Jmi
du8lYKh04jNyIv1Afz5LzysBa2q++6cpLW0ck+XauBa+M9L3JYSCZCSUzXWJ9YuCsXTkqZRLog4l
G/j4b9e6E9ujdI3Ei8vqAcozZXushhc7f1Gxg5Fr28CXjDbmte3gn06XQJMpAjovGYlUz1ulavon
pFjd/0S0RkSACZvWpszEOhVq0Bayijnjgf/Drp4+om6zML894CTmSTs/4psBqve9oAYldUXDLrzv
IWIXL5WHI9PV3pMFCbx9wLU/3vcHZVeuaFLYFxMdtzibrlWOlvmFJnkObTjRqd7ngqaB34mPk9Rh
13wZB1bxr7RZ6K3bwb8mjMyYHCUpNIBoKOaNha7eljFTsKENgFBruf+dY3plpKXAoOHOjEdfbX0b
AxueK43ir3cKICKX/sxiVLMIzZF03vTzrnrYu0g60CT7Rw5YmXQSpAereyUFpaUDb/+TXxzyYxo/
d/xpDQ3/r9pQXqG9SDZ7zJJne7On4HHCwh79UYdYs4Ufk6FBzZ2ee1vR8e5To8y4Rm6gytR9wAxb
nCAqIOG+juBAmv9zgH2CRQtW+2DZlolUsdu97qh6liev+4g384qWZqwAvxOnpOYJz/pgpGUtyb1G
ZrNUU9X4crYYf7GwDZ3ke3qeeIW+pfMuDg8NUozEz/UxCy4JO4ahL780xnRRP1f4/VeLeeS294pi
wkxnl31zfvEWbaw4S/CFJ6YQUZ4QpPdHrTn8uHqMPDt9pILGFByKCYhIGqGBve4uT1N2gcDZ3Lxa
Sw4UoWREPWAliqo5UqKQrKrjcgxDtidlFh1f8Gh4ONIEjP5v1O/UVA5aKUkXBYHKi2WRzva60zLD
sFTxMEuHnBjlvhhpVCNqgIm8ZUW054rHD1Qx5vdRpkMQIR5eDvUCfyHxqYNxmA7rRcuV+rs/ltcP
WZr57aBWs5PvzvbjIbTkV6nb3CS1WLU/MnTTs1UiBLSOWEF71Eeh8s7oLFPbIB0VAFRWtPkvHMq6
8J4awe0vva0EAZRdlv/sM+G8JMDtK65O/zPO7EHXT69AFBWeVzGqtAF81P2UtcJh/l9GSaXUiivl
4XnCO7SC6eY+6jfpJiRnJAP77oopREX0Oya5YX9IBwci3Cp9fZh2fMjQTRvYb4BsR4bstNi4304l
1NMOu6uZ89Ri80sKIb7xgmltAK4ZuoG7XfDp5OhOOfs6UNMfzonwpcbKz4UlDSAIZtXJVMS5OafE
HzATAfnS9pOOquFZgMACHIRwMeTrGeabll7bdhksbkop/Xv86iU5xvuQt6ykvLwETDo4E0BF1XI0
h0GshNYbaWhNQDKPeXMBh49VJgRQfQVRzRIUY2zt2wkiI8X0hhS5YJ46r7bdzF2LJv38FJnEtY2+
A//hnncOZh7CT+JnzR+aLWjjBTa85ZJqSbKEfBMDNhCdX0866d/aUc8GoSxyrhoTYMXpOXpuzOWi
78qrA0a2tLBQF4ByqNqvWhfG2ODj8cldMp3y8bfVmK1QsgOuPC+R2kS/l4XdjAEtrWxUEp0ieU4u
zzh2POTI0Jn1oQwGOL7bllMcvxMisqC6Wq6JZcCpbEk0D2MW92VCOEfgYeGNHCYyXFPkOdzNQpud
yTHHWvPvPEpMlHgv3+R6joaUXUbEBVHg2Xd5+RNOka9yLcQzR/+i5nFNGOpOiO3Uu6TQBBvNNyid
gX0k47b7lq3tcjvGRcYuEuDe7jv6vAjBZF3TdX1U2VjvjvjkwuyQqfwGCKVaI2kqqYs7xo9+P5GP
9vTuk+4p4yLRqEZU2oBkcM6cSEt233cPTliw6CEw6oYaAdjIhwzjKOlZiEHjaV8GgYLmd5KSpKm8
4dsotyX4+JqM+Mb0HcTF1niD1pIDu/NOl1QNjmqOI5AsbIxxhoe2IkCpZVDl5nuMLfjZhW9YfTwh
Eb0aDTwtcea2FFrZgZSTU8BwZhyFZPGyKaGRhQ4tJFUjDBTgt5Ps4iQEpsXpqcS45qwxWSzi9aW1
/B+7ajjfbEKqX1oFyvDl746qehHQIWHurkcwZVYHCZb5GbADkCN+Yl+2bmmDfZhh5QbhyG5wcJaz
L8A0i2qyrnlSuD9PFvdedsfbxq3UhrqAY8NcqzJoFZHNimZXR3QA/LnM2JnnshBNaou26jNMhYHY
+1kSWSR8d42nUj664b042PqIibWLZAKJVSeikXrKWY5a1ORNkS+ep/HJQ/R0v7d0fpCcgUv3FclF
qsqzJT5YxTPCBz//vK94brjO8lE92LA+g54cnLeJklSIDJndpNq8cfr6ZF50e0SYrUAGA4RlUZMS
SAO72cjjt8MI/XXmPguLxilmClUKiMlDx2GmQg9vNISor/VAQEPCCinshpBHn1TlknIkTAnRD6Rl
6B3inVWJ24d8PWoWMMrD+fbWQFHo5QKo13z5kyC26HxDvJApmC0Opav8J8+HpU3bMsnZh6+ZvXWv
XdGAkUsMiDJNvcXRsnGB1ydfzME/lzYHtX7VTSYGOFZbvXa2OFFLqdGyNNzr/Ap1Avae84ODe8qi
i6bL2sxw1DoYYAJ6BlQb1oa9cK2rIapJeppQ/iHUpZK5i+SYuBqCOJGY7LqPAkcuwDzsISO+GyfE
58240U0RgctH99OhJOo6qSLLQVKWF2l/2aRvx65iR6ngPeWb1Hn3J075Nq1pOISfeFBglh4X6suQ
exImDuIcSyOLVk/mVd6gtMuym86qpqKQApgdxLc3ZGZmSJOhKMA4f4cG5RlDITk8PaIPlzgmTVpf
yxSxxo4N9K2UMEJ6+4qOOodHnEPqPkBXTBlUXgg74mSmF43UEd+0E0h8nuWOb72e6bX/II4SbXRw
an54aePx988Ue6dZcDgA3Yh4vn2uUeRVYwzutxzF/oqv5Zf3FXQ7N8uwrNpCZ8Y+7QwfXKJ9v9i0
KcQ2GhTfWud3XdGamCkP0V15I191nZmCV6JG5wHHS3H0TPCllk6A4nmxERCMe8NoenimrzSUj9+Z
Uf1sqz2++04Q/QYFhp55CLnNcmiLceQ48i8SGm4COqJuVYjD1Bd1J9LSNZ+2y/iIMUQeSE7ZDIkY
P9UFSvaqzLqkBsHHgt5FWlLRc3dEYg0938Vhuo0YetYnTR62owTaBL1kzJF81ShPOUK1f5uMoFAo
JaIaYAPtwxJTE6MxfwlVMKUh4bmPZJbDbWCoySvThvklKj0tID7wv2XHLxX6cGo2iDHK7BSIq5hm
/atW3tsNu+ZOrno6iyaT6h+PqhSy/VGEzY5MIzqXT6ysRlQv44GUtCU1mkEtqHFiImZndlDqM7ih
bFot0xNCFcq5Cvgo9v3rYuyzwK4UzJebuNfDgnW66uJHdq4Z4OUc0YyxmHaiwRQADAsLBqhRMuZ3
z5kTOtfMkVggP1RU7bZhWhqYnrK24flTxj0tJClLdPdRRUuyBIKVwGcu3FXwakVnLEMvdGjolPnJ
ovB2F6M0EBljN/gk/wAS2fdVsPI0iaDf3Kn4RA9osIQQDmg+SzLvwBYFX8f2KH8ywsDKOBSbm7Xg
I0b2Yz8KmuSqMiTQDPqnn1nkx2PmjoGRHYyAAH10knZmYxC07BeEha4DMDUxkl5uxJ+xVOQYLCk6
qz50XvxB1T+bokiI3itU9Wqif3iHwDsruwAsqFtiGJdm0uQE578q3rokbubgZTvgTkGviqLQqeEg
zcpkfSvBFR+rPqChhCcYPLr8JJ4yNf/jY8hbj+uZBA6VNyez8E1np8380tCKLBqTcuO6SmwKMWvu
2qQSOt6I9gcXWADwTpQRvM/uwdz9lMzABqQNwTC2SqS/3NzpR8/ww8rJsZF45RGVWT+nhn5HZJqO
OiSsa4jAiMX6dfYVTXFFhSzQnZwxNNTA3ShI2FwVSN4YauZ5l/vZhm5RD7JsT9/CtoMC8wIYBP46
KmrgVHfVATxE96HP6v5uUbgifhBxzH3dYgOqiFoajcYhLe1b0z7bRisBtDgTJE4+zGWhcxcphFh1
Fg+RqZjaTqj5iGR3qtGskH6l+Rc3kOGlhybW5a2szK9gR/jfPD31+paxEXZM5VM6s0GtrKL/O+W1
mwzUBt+pmeP9xgf7JqEuKnNojVFrUr5vJoYqiRc/voUGaJPeyjbZNvRi1tkMuIobdQ1ZVhAVxoqS
roftTxM1QCFAkinscetl+Mqew3AQr8Q5GhGDYfRmpbUdQHJqX6X0doDn5/U5T6UimfVo4m2XMc4K
OBdes32DD0MU1TgVvZnSBe29/32IzqV0dxWVOdQZR/AkTAJqLcb8xzBB5zl2p61wps8ky1pmJZ9G
tmJRUj8MUKkqFmAmdx2LKqRsNC0PilWOhCjgFoiTF79SS4Hw4OOxYhUCeADXYn1HFNTPGpqZg2iY
yLq6nELFkVN+immdPoqCaiWhzu5FIMcPc1YD8QZivmmzjfI0n79HFiF4VImBoOBOguOQ3yl6xSxc
xBCoB5zXxgXZRJFUp1ZY
`pragma protect end_protected
