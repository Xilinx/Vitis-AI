/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
c/7RnxbTBLBfmxPe17mJcVsuTfXstL6JYod6sXIR2GqRyG6acW67xZZBckjxeey2BwNcWEiyzUF7
2TlI9yqQIRtqyfZ28RnxBd11ryhK/mG8Jeivm/7pPk7oGHPzc5WNx9o0y3yxvZKYVUr53xW+Dmvz
WjAjJUuRM92oq6yBbwP6I8ojKVXwi3dk8CT1hKgJp9geR1noWwq9ydjsiN0RLWcsMMPz72r9cfAn
rHgCu1YUqR557bMUVWznOKitvJ1nQQneO6xKtvyQIKQuFKw2xgc1yzyPgFEI1G+XimRHlit+g6Jh
a65KSkf6+Z2BE1Hh2wgwj07T83agUkMET4LpuA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="h3z2bGIO4pbhp+QeehJ+b/kFgDlGqJFZ+wkTvaQEnxs="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
IlbOgh+gaY74LJQCY5qLAPUMPKfX48feJPSDOmPsY5XlGb+Sbf/WmuCndbtT50RcIqIr7oWR4j6N
EhYR3aurfpVzllcJWoVfD7POl/uwgdn46Ea5d/1c/0PQV4KXyROMTreDogixYs/qn5EttY6CAx60
1/AVI1DbD09OdH3EaydPDG5pFRZ+pchzuwbsrIyng+1uwjxXxmvo2fKm+GQgdhwqAg9lasyztHVa
5w7X/QmX30etIi7beFDMO+KObIPDTTLi5TlcOAT5uyPr3yi73wfC27lIjtOnnRT6XiLnTEL/oj9z
JAsaJiKxCBssB1O5alwGtMRaOYTAkbku0478zXY+n2a4Pkod9lHQhOB3F4xwUEXyOUFQHRyh8PzU
PvBrfX9S1J/lMdQdnqApZLuo9QgyU/9dSNu2sYGQPwooHd6arqbDiW9HjzCG9fO++Fm9JVaSRYzu
CXk4f/1VsvahrcK0e+MqCRKeEw+wYTgCo+nOREoh5sUm1YX5HyVSMbwSeU65nqma5GWe4MB7pPiO
5FLIwI0ZKc1jibVcm60s7Oh9daDmO+vaGstfNdnQ4/p1Rdjz1IiZoXMsTPSQjA6tagst4gU2++UT
jMdcJy6cPqgXAMN7JETjG/6UJQkMot6yf775KcrpyM72n82LNbcrzy7u1697rpKFLH4kxr3H4rff
GkgWZEiaeddLpKI+UPMEe6bYPweR3rSKaFFC8j39otmhXJi709Pu3oyg7+FvyL1pTZKDn8K/VU5u
3AbR609y4yXs5bRRCqyT56mmM1xFa7k39Ln7eYy/Pz616kF9pNdtNU4zuO5QIhR8whtBDy644pyc
GRmUM26HjL0xlGI5MvihfMnR7skSZDFuHtqu0D7UsMK1KTPFBWwiNnOBIYQAZQ6Qp0n/gHctoT/A
nCHYV7NsngFBi5gfPpY2lgSkDU7gexFxGVmfOBP+RbuILJQ4FGKFcSCQ4wEW2hwiCyqsxASrPKPc
WawidVtK665tv8yt7coFkSgZoHL4e6Kc7cmIL0YNWv+H387L3oXKjLlTWbcii5hxmi7ka+IlEsiE
OaZi0WJOVHT/x/z8cmAvK7o0SVdT5TYre4CriyAFoXUzGs068wJfkx8W6UsCuzUuk8jDeYvDHTET
n9QiiEzmdKD6p9gS56ZZHqWT88XCsiXkwOsuUDjFxPX8StZan6k+mB0TIEpu05bfmGzQ00Dh/RAb
DGyblYTdnZu+qtryzFogbkcXx55jIlrjcA1xOFaSMpfLxY6T3W1qQKsJ1ZGMbHbh1j1nUJFPfJ92
VbTRrOrvlms52VEyECJSgPG7qR1AlYwMItaBGQshKz2T6E3yqAzXoCAnqnkWxxwZ+Ag0fH3JIpy+
sM8cYHNB/rABOVB/iEoxdTLfCWsc08K54Fbz6pKEYixYBvMa/FOZAt3R1+llB0GFmSeGt5fR0FGM
O6iX1GZxnD/P+Dyp0ofMF9duVgjiN+iYr20fidBiZs33OW9ypUkx4EcDSIsy1MZ8cBLn5LQKmctw
ky4dJlDFh365qlh0J9AwRxtiqt48jzb3/wF/tUbo1msfAzmKi81ZLowoz2Yi5uRWiajBRv3mfRSY
5j/wZrEHdpHTrewIkO0pGtjS3lwe1qxk9zjHbB5+359JnsPVb7PLMFjkNW/3wqWKWaYkgXJCoA0D
mDuFx5F3IX7JxhjnT5KKfhD3oMGB1sV8JSA3tuaZmbQ85GjIs3hpZT9cMuyE5dhnZppZVfNikjRz
xvvcuLOylpuTZx6lUjLR2TzreEwAre0GDicJkbKsQI8d/qRcgodX41EvUikah2TO59EQoMs2qltt
IfNNoKVQZi8B1PTDW/9XMqqKnBTHgVCFncrxl15K/MorgOJoaWMN336+adKCMz4cWCzPIUHJblTP
Vq8DtRZSBOAht3ikL/Wf3jri5718hb3b/li4Y65zQL2hC0SP14FOVRrLlOaRiFeIsN2RGlOH/2+s
6P1fqc+6BZQf0eVAPYtcj8pXaTeSM9Vu4srRC1pmMMJ/l3fJe37VO86hwINSemHEz+BHvICbxy8u
B/TaLg+Wy3JKybx9gdVJvqI6CeHHe4URmAghWq+IFIfRjlDc1j4pRfBQPb3YdlEZnzA6crEVjh4d
Yrjldj2y3UviAAsQcDy/p6zkTHNvHQNKoF6lWcZFIumuc9A63tlSUf8SXTzhZhxO19rzPDL0dNKU
LrYpKIzCrimmxJEreE9kSnW0IE6cFlKAqU7Oz3HK5BxKIZ/Q27QWLFsR2RzgQu8mpsxEIH8ptfM6
+RM++o0g7fX4J0+g7OGW4vky4+cbwJpil9Imx6hGqRFiP/D5FqAqTtKFuDWsI5NtSipTtPv2lJB4
luMKftCcohH2w584NTPgA41ejN6IL1NO9VVYgr+HTrk3i2Er3h4kWflNusuoV8zlmhTKMG1LyRP9
0+sn6ETzhwu0oa+k2Mq+w2aSR34sCOxM5kxMNlQUcstxclQackhiIY67nEm7OBxgSJAWhgDeuX1e
tXsJEDLf5/dasOCmLwNkOydSyh+xQVWimwKDuu0fycRwghUJCEkU6wq5Fx7zHAGfXOo+UDXS+FAh
XIlXM+mSqXjQF7awdyWKnuNkqprqQyX3EkWLtfY7dghv2FZY2dKkqo9fV9J380/i2klIDt2Wp899
a736+wg8xGeAskMLAVR4oHLKCcz8H+XU+ekNFgbYmkYK093wmVs7DRweNpm+vhFAquOHpQMC7cFa
uIIsJ7Fu+7R9vTuctRwIl4LVodqCzfWx602UrEMJnoVMI2uDALqulE+pfJE6wwe9amWsChU7y3w1
zN5JYBgZW9E8VsCjeJAbgDgYKIUmtxmFZteePIF83Xn7nV7kCd7BZey0o4VeGScS39ma7vLIERtY
J85K1weI+tRVvf/yAxMXAJOZ1Uof9nesC3rEdp9PhKPztKF8X7GZU5dqxCbx6/dlGcf0YTveMOkb
RV9y1n2pBQpC3FaFmM1yzalqi1S50U42aoiw0JNSwRCUin2Wg22UFJDeH4tEAMtJgUJ9UN5fJrjs
7LPPA7lKp/zoYHjRdcIXmaelaS544zo+qz+iR+9XhMH6nv6JsFYgLHO/Dh1pRekDZD37QL9FfqN9
n5RKiVAOC9o48m5W9CkuVs687R+GpW7IoWanhGqz0Bq4jwXdAMQ+2E+u78XBRnhCMOnqPXpFWhjn
C/w5PtlqZtrVdNx44d18CEeqg5wxmLIerTBTLQBs72jwsmfxqxmHnjiccf447NJxFgDUSKCQiX4G
HfaLy5u4/6+HjO8sojb3nzlA2L7RTrananoYhBedVTHbbuOBe3jGCw5JkTqHOnWx7Hd9JxWEySFl
q839ly/6X2X7IPbrl22uKR/DesRnGueTLE1LHcO/Q00gmWL0SE1LZ+er48pf/AHrTLFBOw+8vc/l
zva8eDmuJpvVZ9IfraENEWVl1DDT64WkFOnfgtOldJzsopLA1NnS7VV22SHH8DfhZst6qgLXcM3z
4W3IkVWYITxwKbD7H+sY+/xHAfeluCF87HzW+Pz0BvTiZ4ZSNfX5+hqUgVLBwqtDE85EzdI9U4+a
TgafVRHuyVZxjhpzQ7X4yh7ntiTqhjUjLygshI0SSqDiqKxBpdJ26iESgYp11ZshifeRZKtsDM2s
fR4jvWkQ/LUpDrNleCjUEdlYl6rcpDhW0Tkhdg4297ydKqtqok+x9xQWHpgyTKVzxDTZZysmfs3R
9LDKrapP8l9/9lxbYOqz7Cks/Z4dnNGmi8vhWruet2FgQebODU87YVx2a4Oae+La/lu4XFBQtepk
gLa+GHCNA3c4YTsbmvJw1it2WKkwoDW/FeZLxB/FLL5gF0UlMWGV9eT2aDUJ2ypije7XFxfty3ai
V0I4pPOqZdjwbEkkq/qVZiXylHmEuhgLQ3leKIXRgK95fS8UlDPcHpSCwldJNcCM8rmXbvn97YZt
uw6faE6I0gQ6ZEwaWjuqZi7AcnIy5Z2T74MLWtKgrlt2yQzgXS9hLFBtb9vAicykHrGqKMyP5gQY
fKIIsE21Q45R3ksWuA7UfdmdSDRvRCZR9cN0ye0s7QFfp/dj+20UxKyua16cTqrDtqHCmPAPa/dr
dZftVgNMmLVIctLNyEDDxPcjcTt5djkH35Qgdh+qbCEJakgxTCIstoNC2wsL0Rr9DsIUUGwoP/q7
aZjcl/3YSfYLB6EdmVcQ9G2+Snl1sYlVR3zkEnEZYdpaYlueCi02HxSIva8AbtzIT0e0PEx71VTV
BFcufNPYhmcCc4ex9UTnpllz7Q+rlVQk4zHML/P3oc6V8qIHFsxK7FhGU/xLFYDTpTA0eU8vLmwN
TaGMPQrNXkic/ltletSf8LzrtQxtyw0y0ibEiZaAUvUJtM2QOMt8EXNJ5g0ArkRiuYGtQHTG0NC4
V1RH5zyTN9Aabzn7rn7hQfwakwykFc72nF98jXfFZ9tbZtdfBtamKzLs4j1m5ibw6Bhpm4JXIv9+
ZntEeTCm8G+p5GZrPhLMObHLUF6Epiwv9Os/E5tTNnMNOBnrFyhQYYIkRJGP3UNwqMDMOXi2obZL
zQGAv1E2j228yLp3lIjSuH2BH1bnazQXtzk1xWdGBWOtUQRjySJtPcjvGJeMj6EZ/PmQQwcjCBad
s2yecwFkNh3fDAnNool9mhV9KLZo87W/TWAKqmwH40nJNNN5Hv5j2ViLpcMhEjgnHHAEg5YBuFnG
byUyVEW3YYvF7hrgiVeyZGbrCHmzZQ238J66MMhAFgTPdGUXx/CxX/jkrUnKthr2+t29sxvLORwZ
JJ8YaPzOq9rH90EX5kS/6DR/ps2HbYwKl+W+zUoZBm0TePYJLqfcFGRfBkWM3gkt3f6lzG2R672v
9gtROFPzx3cC0+4WcGjKfKbh82uWnYs265JHp+KNitNrCoZMvfazgW2wcCeZhSnWObqGZOc29hEI
glOfo5BSKANXSX9X754Pzskrw8mNiP1UTdIF8IHKkXg5WDuYau1tG2uL27LYDIuKiYlqcyugaULR
I0wzZrYde7u7cbZaoYOvWYuBZDZVnK7xOFZ5XQ3dWSCmNIgCc+zmRmJfRkd3RM6AyiwONcOj3pDZ
3tpR8w89/Yi2VAxuyOewIl8WQ6zOyzmpTTJayR4NjjKnj9xE3QzjtCU5KIOiba95AvWf4Lwji0Rz
GDLu1qevXkgBD7HSttHVxSZJPa3hi8DG6PQRYRvql3gh2OBe2DJTghmFfvVbUX1rhWs2kiBMtiDT
Rsbj9eOZEwBkrBWpS3jUklDwgh3VZs77/WuoOtiHn1POr+T3vCI6b3s0f4jx1jFl4Bw5BX9+RlvH
Eld3YO9ADb34o9ywvIE+/TLVaImLnpBlMMKtcNl2GPt9dwxL56RzZXA6PNet9rOQNSoObqtaGYSJ
S1IjFCAbfHU7EbP48EhMBcQS/Md1YMhnFuMZ2FmLFT7SBtwyt4/Lu2i8JXcPSUDXAx8m7obNL9b4
0/A7iA0GAXkWwC00122iYcAmrB8XN01KjpkdQY2SidRzZgMvf7lsG7173htkPz8zqPdG66I7L8bA
MQPsXiVZVMEafvEqEZxDh3XGKAYdAPnZl0cq0sSgNkBOsgwcZDpkAiD4iPPpAsi0iE3+gBAkcIm6
L6xAhw7D5eAqJS7F4x4ubTOOX7fqEt/4M25JdsLZ2gD/t/rEYvI0YHHmOeh4DaWbpv9hr+pa12UL
QJc2hJ8WmjTteXWF3RAjUQfKSV94IxisJR1fQvqjdGUqtUkys/+x9SrgOaCi3EJCtr4wWlSQAiCI
nzTzEK14Bc8AMTbTU2C92iJ0jOl/7y/+2mOP6gVsaCgeU8wMv6DChVbda4rVAn2LdpWUEG06b5FI
dWXOCXl1FKqKivfByLu+MkKUPcmAzSK1eHngQIMqiYFn6RHk598p2lgsdzOgoPItQr8qhMiVsFXt
mYTi6hStu8bsKh4vnxVNege9GBdF3JWZk+8/Ht3y9JElRQw1888fI5z/iTHp/xY78nJ/k6mDNMi2
UqidwH1wqp0tmUzoOcVDcVFGtgC1YM2tF5QqCjebqSpyFz9VIzwOJgnqIA10eLYCzF1wczTZyJ2p
XzmqORRT44iX8GIXJPPxvrMzVYEfTKVo069KNMUIdVZIjtJ8SIddRfHOAVCe43pdaZVb+JRI9T2O
5UfStNJMlpYCsLwhNgX8/jAqMyLF43SzPxQuy1pTGXIoFeYlfi7Zvrq2Wl+UC7Y4/8ClpnBB0xAS
UWZiUiJZ56mBGotw2/OeB2LiG6Ki8MGjMIQCGq4/rNP8zCJeUkJ8D7oAvnOUtdsw4hl30wIPdGmu
vSM1mLHWCqSn2aUSUYraWLLxYX/mBBVrg1xq1qJGzBwZkOXWfPpDsTMV/WWXx6RUe4wHZ1vcvGJs
39tQ6Nhxk9DUB/sG9X/opcv0JvLhTo4d7JpHN0zp2AnCq3ibzudcliAiq++FR68Ibpt44PcfSB1F
1rfdRkqdR/BD7AdxXJSaD6eDI7aWoC5mM62xTCWSTISSxnrEDL35QFob5aB39k1Q7Nebb9blLc+6
m/EI5/5I5mgWaDDdZryp6c8l0klcGIYKBcb0U34MghVFNjkiS8YsdK3ElkWDq15siMIEY5GSoWVg
d1/Gh9HUdU7/yKIP1MUpbpoxT9q8azCEKF3Vt8yZqw/hpS/ycSQQTKchwlq92wcufhIPRJlJUmx/
Zr4xxX9g9R9uj0WUODzU8T3xh59rOAfMm+ffwU77lYU56Yle3EeIw2Cx/Bd+IhNNL+x5eU7Ylxdh
8e6cPAYAjc15c9oQIjBNen+o7yn8MPbIzAk8J3WQMyzx7QieoSkFBBjreJ64aySwz0MlMBDS71r0
DkH8S2jKkrg1hccJm25+jl7Tuc20GJnsk+/GimLTfQ6HfFGbmwA/3slPmNGGcGjjKrQQLBbv9YGh
ednbWtgf3kGZXVw1U6pDEIBpztZU5uuV7M7Iws0Sw5ZagMk+pfAW/BVqzSZvGJGunAK4dtEJeKGG
RCrUFJ4ZsZnhDVzgIE1XaDV3SVkvuHIVaQvFG9u/q9fXkaUXhMhG5DfxPvbaiiDB45bzOuiTtdIV
6iQwdY72eS4ceBWbd8Jzdd9wz1oNXc9q3XxrOzKuU+DeGjusRygy3EMbpQ4ErD1Oy3V1vVhlnIxG
iq+Azp+hTrJFedOgK85VZIkgvtulgtzWoZMaKTXuanWgAX04r3/qwHBCQus43WnSSIMmzqfRBb3O
r97UtzXVX+sHyfEajkgtqKDzD1x8bgApZRmH90e2KbHDSHhTWjlYR84yxw/hKvyJ6oGdEi/4Vmuh
ai4r4tDG+ahy8KLsBiUy1XTczR6e3iZRQHPUFRrp38BabF61dxk84y1CreJoColjSEQp2QQFMKHp
2GfkIv+DW+B2D0o/oTtUk7Bwaf+EpBmQ2GP7GpXxNTeyh8wHbfAB6mdglxwrTMAbrUEF1GudTUwM
Ueh56aUovz+fhO1r8k+aK7V6CiM9IOqqV9Edh+BwemD3ywQyhdUK8NMAyzNEE3nQb4lhkNTRItqR
W2ir7UZnE86ck0chnpyMyJHjsssH2G+CO3H53LTh6mJISRnfO0xVIgUUf6YBFg2edk/RA58GSKVL
EB6UbjEkWI3zCyrMA7W/IOLtINXbJe4b8oSOurJiIk2s6F4YkrE7PPD/FdBPBpoa+uZY/0cbc54w
bo6njkjxpo3EWGOq4XQQT1qwCAE4Ec18en0q0e1E8TSgJ/Kw7XFdPJbOxLdLyrQa4Y4KFS/KGLd2
qlT7TUQCkq+5kBpb9NZoBTv9K6xGfXGynRgq4VE+rCbwyT2u0SA452emfrIL/FHthaIvyMk4/4gg
5XE8G9M09PRxwMENlansh8V1iSotaBmTWny4bCeJlphf3WLxk9T20B3hpnjlURuZyU6RSzP/uIzD
eE2m6/pAwxKl5o8uJpRuxZi8o9JDFCPYXwhTJiT4DlSFea0SggApQtACYIx/xNbI0omREoj+lGi3
X13y7SCcvfY/W53Gs+3lYJ+kRH4C/wSm6tZE/9xni0rYGkhlqDthLPDIypbseByTMzIn/9RoSilI
xiquTFWl2vUvtfft4SOZNGgV4U4taczvB0HaA8kXyeKXhT8IJRf6OOZUOqllVeD14jbHPEBLewsQ
ej4s9BYlk90wgHPcc2iIHk+pJa3iG5sf2OHAtNKMD7gM3/EsMLNcaB9fGFPHYxmEIHPJNMSyZVQx
es7yY0jncJdoOOwOwAZnpmD1GeUAmrPWwlYldIOZ1HOevBEhV9fe9SlXO4mbT2ywksTZ+TPGCilc
0t7R8UI5lalPXBIXv8L8mBD4rsNiPzeDvBAJb8WcJkrtv78aaJ6k7ZQMopjWDa6g/Cx5a+IpqKgd
OMVEAVTqHTeGENSxE3crya/bBqWeIn3Ntev7C0Oy5calGRdlX52GK5ifk6xIbUdyJzfwbfJiI3Er
AfAA16N/pajNUWWkuZ7Qx9t80iyOBIHE+kamfzNI8lf3zdU3K7nL7dyy0AFSN9mH2WGX3t5U8yUf
vOaN1m8/JE74m62FyXM/ATqdCtBUVlBfkm6Jqx9ni4ClaRQPe/UhbVbEivd1qaAXEtmAIHkyvdpM
JG8zHmEUSLF2lqBzmSYNTfG9MBD17NCzC5CwG/+c/isqc5Ri6GsdQ/KC5W55eNGQ2jv+JHgWeVpd
d0KEnEu3TE7wGkkR+yzKx5XUdGrBnmkar7RCC/sjy2s8GZSUFVQuDlSd2T+nAabTkh18sS+EzspU
sTQJ2tCkyVVW+33Km7Us4dVs+8iOux29T/qa3ELqgLOdCagyXB6nv0oIJ1N1dJsA3QqB0LZBbOKA
g3Rak98L+bn63rs2pmeZUV7oqsNhUA2te33uEE0ft0WIG4xtsnADpRy0zpAiubIbZ/+hs6NtMYth
KgyPiakcDlj9fyYf93JRHTPlRNB0fj2EimPevRYkCqM4HPNKMNrCrvKV+gHGJRuf3zuTTs33a4lN
Tb/BB/V/05Py+jSflN0Lfn/lXXl8ISwEGFmmNTxhxt14N846pkppsiw3fTaAD1FbfJdfOXe35iMk
HXpsJiafQKYb37hNcVF2AGy3fA5hOhxPfteH34Xv6oW6L2r+a3gAiQ1kxJhUWIEu18n9odZWrAmf
VUnGDFxWAEicpNAE8t7HIBjm/uJ9eV6V9TtuZHsNbmWqHcETBZwERSaQ31yLCQ2kpG7lGFE9umH0
zMLAke2JVqq4iMLDD3B0oGKXS/rqQaCMGkVAYpSA3X1xtwxfjALalYCoo1J1hnyUeblffTk3boeW
FAClYQkwDbCy/xPFYqOUi9Fp2rBNiyJo4FCOo6lISBkuRfhVN0owSop2WgimuUTv9K9KxojfHc/v
U0F5nkL9LXRT/rRvu1UOhZhP2fowWpCbl1pnIODMYfjFcuWAqDnwnBHbH06Lqgz4tsD0MZcgDOp6
0uhYXU8djXFFO5RPc9seRED8JtdtbEPE8P8x+K+B9UA/rLuf3zUaQCo08TWfEhxDCwZxzEpFgdcO
fdUJwy7dAQhph5WpvCwDCOKS4/eMSsz7tu3BYxER48G0XvA7FS+lOlCbFxWU0okcH97cYRoUG7Jf
rvU9W8B48aWbdGjmOsM6cjG9XHQ2S0vHpYDa2lyFcpNUdQf9tvrMdt1h+pNLy6IWd1jS2UBSgxZZ
a4FPipLowJMyudB5YzYJ7uMFa5yL2n6f6wr+bcLCjufSyMEINY1nvWNMslPx/U8KXWT/0XO6M9qo
PVL2DdiVDgeZnQB4Ezg+yenofkRMQW3OZH/e0FFyRcpzK+9Sksnxmmt8qG34BxCijxBa/eYC9uld
GQ5ItdeSSRT7A5NIS4PA12dO0eVnAzP4/EBc1/4Z/1K2BsEEaIJtuVYK5//Y+9POLiKZiXuPevk5
C2Oxj+4SYCocnZ+1WhiS7ZobPbsnkjGV1A35cQWgToKhXSDYFXFNCuwjVUrTntzTy34WFBOWQvI4
Ko/YtPZyj2U/sBFbJ0ObWdDG0N6BDPghuDrmJpbN0KMi3K5KI7tjCfGa+i9HL+3/6s8r0jTdEYhG
rtuq/dxwC1TwO5TCdebUsw9if3W846kejDZ5VzrI33m9gwXRmc19AWMrm0VRfcNdDFul9GYmhRcj
AXy92Rd3IafEko9RiStVYbpwgGCRlDC2wqa1hb/44YBbW7teNt0M1Ob/dObF+dH+WukyFRlmE4vy
GophXbfCsZERlSpzCKq7JeAEtlX6bNbi+/6N9JrWFbjuhyOqYELYtLgJoizGQamocKo4K0BIkNLX
uXKVfJOBNaE+EPbLZy/Ro3PKeqEnRDoEjjdiMaIDy52Ldhz5vjAn6nzT+g8BmgUyGxlWNp1tDaH5
ynedJSx/7eSAjMG84fU2GbVspoAw6B2LuuMwJFU1YSnFAxYe5oqNTalZRlQPKGnFkppw1AbqigFF
Ag1EMt3XXhaIke5tIaC0W+nFEB8KwYeJPWydtA3O+Q/vQN6kWl92S5mqHlFYMAQBORUWkOZ44+Y3
Y4CSK3/VoaK7GcGNvqDglhP5KKWGtHPl0UJ5Q3EyjSqngnITJ5Ct0bpCczLNhLpFyvGnGMQvBh2y
4H+OlI3x95H3L84DUPHhyX23RDw1CFUZkNYwr5vhELFX/zHxDflJ9gWucihLCXdpCSnVxE8VR2Hg
pTdAupbmXVijpGvYtNQbu3qxiNrOZ61RGycTfHVrOOSB+zRl25IMnMPrN1I8la7wSHNS9UEyFC9h
LTC2alGB88A2EoVCG3VuNoosv2nXeeUAHS5EDZ5098v7B2nP2AVbSnFi357sOSDewJIH07G+2Bip
1X6PkxmMLCHVpvEvbZKolpytDvRpC2zmOEZuAiYcHNxH0pXdgkmVdPM7Jaen8pSCGypl/Uvc+jh1
QElOk0Ur8GiR0RzbSPDKSF3lwCAjRjW1irigrglWcxlkrVNnhf4zPOxx7CrNPfqGlIaCuWX/DDUk
D1Aqb3qIXOylEnCAKo2tUWiHMFx91RO4Ro7VYCI+njLldS66TgzbdGryMcAt61trPoR5xMzFPxYl
QqpIpXw7+vnIPOhYUBTfdWUg9By2bjwn75bbc8Z7004yGdxEq9LLM8SWvt5ikdBcXxDsmG/Pys2b
cz34X4ZWaoDLI/a6Ja9iKU+8mouq5iK3HKgFqkLLUfR/V1ALdO8PrXNNv5WjGe0vUQZhOYLGf9m9
BvFhciIPxfIGpeQ9BjbnizEQTeA1vNqCMCrclO2wUn95RXSBbTqx7kyKn9t6OiJ8RM447fmW+IHR
TGaIwSj0jo9J8XI+o1q5UXizG4jtRH/LYL+AxpP27GrjSjNnt/uFfDmkdF1qqH8qe9e6nTE7YBgH
rrKE36MVzFRhcquf5X8CaymZVmhjx7zDSTcMssrKANLb9o33NUbKpGTAdWCtDGXgFN99wfHri5AY
h8SwChlVx1g4Lf23OycrJWi9BIdScn07eH87T5DRgFJ/mIXFqCdtH3swG8rbn6EY5joWhT6iLDSJ
0QmB8dYcbQaNJm6Q0i8W9J0rKRLTfLQlIthT1R6ShqwPBEUw4rLAZK3kvta7FrHbL7OvhSmM2eQ2
B2wV9hUJlxpDYek3f4K7CFcjlZ14wNHhjFgFnHBVd4jXBoM/pDh1afDeIDAlmnWmAZ3OyKtxX8GG
mEtRJr2oDBq0akt2h73Oqc+wGBszk5nr/NmVcm1pypf013Jnz+o7R/GQuBbPtGyNPjzzCzH4O3Xb
B7rWXnXuVL0dN+u4++ccdS/qyipj4L6/yyiQfBemkMLflA95Zo62C4biCA0F3UvdqVJXZzCnBUb5
ah1OiztVciP9wfxyr+Ui11nk+NPiH8R3wtsiCDKug9duXsBjpqCQQrXig2L/CshkTUfLhTTZjMcM
1pk4wtuDN7ph1ZfWHBw0pvUKhrjCEPDk86S3hkU6qaIlmdvKsaXLb9588kKKJ+UcYYQ9Qc0X6/va
Hi3e+ts3vNruRGSsnbs7gh2XYqcQoeroH5Qy0/sxoVl4PG2KOj1463zDO7JVc8rCLE6y8m6t3sfL
6kM5ycMQ761K0JWYjpUPKwuJ8P+wGlRG/CUfb7//bfwbZyuuFAYsDDUGfwlrCCTIik/Z+5i3CoGS
56DChrffMMqkFxht+WGmOt//rbENwTxnLXT5kEjk/bfhxDiFL5CupjJC8leWUfO5vjq3Z0qi8ffk
nEPeKBuUPOpb+pxjG9sOzoyDLNJu1nspchD4q5fz7CsDyndGak3GkgQm5pUzmJz86PIOvtWIK+1L
TAzGrTaq0Rpok3gpPdxN+5Z3+pRluTgKeP7rmRf6b7eYEIt47LnHDhhG+nqYPfg9d1TJfANubLcV
sN8BTGZaTQrriKow1APzHY/U9xNDHbxn9LQdW/H2qFAMkfMDBSfvr6e3f7N6HUSuZHMqF8Q5z9K6
zcCE7h3H1AjAgCgyPV3NUYKhFiDGLFsQf/Syw8hu9LW7nRp+AWK3+n7do3Q6kMrtJQeWUqPPAj6K
25MsAL/po7GSTQXK6VWb58/RNqb9wWMREvBkPuo4ydqFYAipZAtu0m9+0XabRn7howAf9l0D23Zc
r3P15+UGhjNU5ZYM1r8+R6AZNH3KgXvQtVudPhvsnbmPY0JL/Yd8tKSnAksWw4cCiaR8MXz/jVeW
aSp2EctkkiqkZpO1ZTkez92nVdTPYv76sapQwxjHeuNvR1Wn9eXzBKOa+SHyNB5e6R4O7mHuWcVS
CibxP4ToiyJUuEwokT47GRNwuwPWpDUQAN4aGOF54jlD+FIiXrOP2tE6O93+3VP65m4lQwdm1wnM
VQudibXiwGJcokn4/wyrcwPqUqm6u/EtQ8vQX51eq5BcO2TEo4ODEgbyKCNFAtCdM4blZPWbTcIF
V5V9WLn/LuQ14A6imRckKpL9Na1QNuOZBBs5fD3ZZZKKryeQtejUBQRO56H5knpYVqglYiD0vGcK
2wv5JsvB4r7ClZOywDWJJWXpMBkXzlPBjGRuN6Yt1+kX/yTapdj9l+G+8zIIzoK9WPhZwBH865qj
Cj+XCdguCqNhM7IbociEJxrmCT6vnhGs/Vc6FkpoIKSBz6T0efgzskHZ3ncPnfk7o3GDOooyG9QW
cs13ctwL9KKQ5mCgt9b2naQpmrXlV7XVZpolC57G/ATbuuv8VAejumbFkLQWB3fdwswFrp2ymjeq
lTS98QnX2Q0lmGSgk6osTDrGu0mByuStye0CRAqBPYLtd7onDdsHb95190/cSRzax7uc7BgFbgrd
P47RzreXC26zOIu/idsbeAv0m3WEICV+286k7zSQ2vEML1n/6+9LZFoN/OKcoF79X4Lm+JzZ/hqw
8M3L+kEvaXV5vm0VqKXC+gtePaMSCc6uKkU1OimUYz+peQngeTZuiMYd2C90yuS7CmcCl/6l+2qC
5jx3woQv69MH8tZ9j/t+9S+sdh6QO5CZG0IpvCB/dweRCsDc8z5Klh2J0QdGRPg8cfp1fpV1WKFc
WQ03lTLla6Jry3VnabsyhnS4MCtu2ozPHCi0VMQAOEQM9ozO6zE3lapho79rJALxTAPFWIHowvYu
HufbKNeXzbyM8mmPuctrLICxq0dNhLXmcAkZ8WgZ4k1s5FDIL44WUgZVc6IcHTVOmgvwA3ghGcIX
Rxl99bQ0LOtNqEaWCgIhC5WxoQ/F60F14pnbjuKZFJ4Tsel9I5Yxo4eO60LH3dN8EbyiwDa3E1La
2yXiH5+bKpFgqrO88r7FkVeqRRGIZEumVEmbmMxvxrjVcTajLUPM5YTWUOCkQlU9Iu4AekuPdTVP
k0U/1aodC+/6goAczMu5LxkMfxIcoEb1uxryZDBFS32Bj3/lynYtroiDN3WTHOnkIlJVVDnLLdyv
1WwVNiThf4objG+0tEeHQx6G3AslZ5ihiAQD53itu5CPPjFwy4Ge8yJASe7DW3izIwy8KAK4jo1X
+3FOUfnLMGJbP1OKt1PFqA4nTS4+fHtLDjBaTn9Oe8kAtSe7EIY+V6oasderzbryuIX7MO3JIlUZ
Xf9jmqEN86pyd8eSU+UWqHiY4LKIGbx+UBB/M9007zB2Elpob4uytu26NuIFoR/N8Z6cINkorU3Z
jz6x80PcV6gMgjvXnsZx9yVsjcCbGq5nYMQi9XmuvUoJDXXVb1zxuJ7RmDDEmc+uXNjOrVyfdHXj
ATFaUWM+NOYlvidEphoO50dOWWHpDygONWQGouxsiBBTJGX6zI0Je6TrfREDHc1NGjwPNX5C7spi
OxP1MdXZmkn3fAS4AyLg4BQ46ss14gOoLOukIZ39ENzS9Vm0esOPMNDDzfPegfl8s4RbfwEwrWEO
8RNF+pouilcOIqx3asSKGUNEeeJJKN6AflrnITCiqCIru6jveW+1keRZcoOp+/pQfgO3VBjpjLIX
Q5LMB15pmiwT3qVQOVfxvekhoSeZY8cNW2fP1teqOt9lhJfsFK2PA69lt9fyJrPirI8aiKSkEX7j
S/xxuJ/o8kAtmBjhWutbFq0gk+weEXyAbfEVAjClsSszKVvqledUY5FPXnqDBurbgjqOjAopHbvH
HjKHe/oGqBNLDVmO2uKoM1lgoCHtD6LsrECrt2Nanqua1z6Ky7kir+EzUDj615TAnPRTCk8I+9c+
hxuwQbv8PAshbxSOXmN+l2mDO5KfoUqfmwAr3LkOZIqXuuuJEXUhYo0K/yqgOvNyxCdCWFOUpVST
L9/N48LwYo3mgf3vDUt1Nt7iJNTMT+ep9r5vagmDtTvtab7tTqSaV3barVeS46fLC0ogzZl8dm5c
BBOivYuRx3Zve8+Pei5DBA8DDIInn8UKx0wHGLjVCgli9b6O/o7+PWY9pMYvzRNHkO3ue4ysbiu1
SijVjtW2A5O7yExNaRFj3Q6ckU9VmAgMPfOtwRlDtIwbr8VqJZVAcovD4/H4zE6PMFRDhfayZX41
GMswyjCPrEbp99Czf/BGBzthYYxvLmhnMx7DRDgk8L6MkBJNXvYg1rPvw1bOaCBCSiLuV9luH+iV
xC5ou0//dF9uYcdKARcKblPoR+mqplx/WbfctmCziwsZnTOJtIjsX0fyhYoX3tY9XqtzMIagQ5J7
bF8IhbPkPwEkH4Z3ETO6fySxRmsGNAfyHpl1exUflZaSUMijd+63y7IxW0MJoT4nsYZhCgBbohMJ
b+NJZ97CIUOoW9g9vWUO9GOJOADMLWRyLNpIcX7xiVUIjD38U11nDXSGYRVroNgeR4nu30WMfNuS
avmeUcY/fgU1rT/weWbKw3tbemAkWhD9ZQkFIVpOMfXqjl8cRNoivEC3jK/UINwCNG3YiV6y/r3a
9HJ+3M9d5NCbCaydk7psdGRWz+cldFQa8DODBA419Gn+iprE4t5/T/5bhJlQso+ImzAMD8ifyYJ6
VYZYdZ7UhG4CbguOi6zAu0emmQ+/mUci3dz8g2DJpsmSX4ts7tqH3bDjhZt81JeHyeCMYRBPGl4v
IQ3WlVYceDyCfNCgnJA75/FFnJEnAxgZBdKVWA4REE1Ztz8/GOOSUsIIZxjD9fRdPFmq/4MxHNow
B0/kVRIDrGuPo3sbpYia+2qcHD9qTfOIENpaU/SW7MNk5Bu8aqeuvXWZAz1PBMwTKWDwBVqtKBb9
BZbDOGC4VqNV4agiRMrdxi5S/mapqq9zroRDtfurn8+ksX0+vtzGmS1l8Dnyno9v+Gtr74Ps+H/L
UzWEeGEhDzGPUIUaqUF2FpskZMAJLSdgRztuMsOzm8PzOTnKr9lNLXYHxoItQkKxWfJ3x/SPBn52
RjHOh9xgaFHUdYUQ6fI7mn/GlmcFCtILNpvCLR+yuwy/QyRgfGRY8rOv+oRrqwyIr0wc3tiTz0yb
NhsFP+WDZBw2eTMu54Dt+atenwy6j1l7Bv1niWts4pkS1+HNojWSSvfcGaUasBvZQ4l4v/fdof0y
8y6Bx+qulV659VfA46MZfwC/YyNQB88l4IUPomAdfORnJbB+9LBDtMlHvuaaSeCzU5wiEnmEjd8E
OO1Db57m67pmAwmspXMGx9UxLJXhvSyrhkM93S3rJZvtyKOuG0dZLpb37XMoPSj7ts84S+eFXv3g
bO9YEyw405vmXenCG1bfA/pqHzG+yezV8gAFrEHhEuKh5W1+lq8MsLqpntDQWdqpwMWiWwIDyuER
Mk1SZLki3jPHxmlgJt1Zqv9kU3kDi7uTF3EtUP2IzKu9WBzcV8i/jzGrjSDMYgqOmgOT1YiHhA1u
0cpFLG+AyawKcnSec+7HoXmcdiFVie3R4IfPh9AEIRtHaYP9tzY5bE/7pvGKEhEGKrBQ5aajMCgV
wjYsEl7yGA3ssXBpwV2+xLQdzJ8DrWMG1+Vj8WiB81/2SGzQoDUZSr8//Y2m54c6S57ufT33IJyv
oAs3ysrVzygQDI5EZ3n+7B3RrRhr6ipkRKm5cn/OopOhYi7raUjrlk7AtsZLgeKHbTZc2o+CeQGT
EGAEnPTemCJasmXeuaJeAw7+iM/zBJ50Yhrs0LUdY9ybxFpmCJGX1rfi8Y9rgEO1prb9RRgOWH8i
LxFDxUqOSB4i5Dd9f2HHfkMfwDc2as4aP41lMj3uURNJnq6Z3ALIWLAcYhYwXWysRzohfS2W9Eci
Va8DQVuNJJQO3Igh7PPGoyWxI/iZsxIiwD9kcEtl9Sr/TULBJFO3ahDLFvPIKjgakG+2JhU/Mah7
7OdM6bImIy3RbBmJCUkBZn+Axb7wxYxyl864WHMv2cP/IvwJerBZnse+SWLgI97eW49THR22sYRs
9wfPgVHwM85R/lO9rXeuf5TDRiLupUz9r6j1QkjGTDozMeeOI4Er2z6FH3t/fvSREJ8+4leui/Vu
XM3sr5GM/OGI2824tCVNlynRRdfab4SLHIxQgcE8A2wCIssYNeoxzntN8rJ8erW5sx+tE2gnh3dl
dqCVArOGH+63zfq3YrHpJrtSH9gFpeewrl3mis51mYG3xXOkNcUAiDd4JLATVA77hXWhWhKHPu2k
fiMsf4IN7JPM+mS8KfDa/RIkRGINFw4Hm8+25LpXJFgNWgVYPXAhAJwwAGvRVqZ4nqoGGMXOOFdQ
ZRs6ip8lTqkWK4u/Tqw/TOBQMfafGrxqJA96x9qneeyniKX2cNBoeJQUrHedCghroFFdItVPxC9c
KE8gUI9WnUZMs6Ise5EsMc226/j8GurjrqBfmR0fUV0j+/VxBYpzqzRgF2C6fJIMTsO7PK9PgJ5U
/J7gCkOOROZ638T+G9ar8Om9CaTYUB2jLVD7nN4/3NUzk5xeOIbNdcW7gl7oO17jA/q6thsug195
BO2QA8MWwDY1nDRQIUHKsPuf98KncQv/vF/tmYwVMbBT9ASpspbjXz3X6oz9YUBi7n2ErwAeyRiD
Ni+JBOZ8cfQcJWgbId2HQfOMRh8sxpZMBz+lMX0YrNSlFv5j0/bXq0fAu0tN+BjR7pvn0VRx+Oqo
gUegvHxtnlUwAFsi4eItVmXpJ09kHr1bbk9/WogWlzYiJotj7pmm9vCpnKpQuqAGgxKgT81nJaj7
s0P5opks8O7Ku+RmMO8+fHBTfVVVVYsTrNJesg62X53dR+igZWhyPa3qBm5jOY833GUetINllv3l
axVfTeTblEos3d9qKV4QZ0KSPcL4f/Ubf1WW6eNMDAbTE8rhUSlTj/bHPy6evnMQ72bBi1Uwpv3G
oG5FRinHE9siy9mKAA+cCDoUn2swvVXEuYIuCo0MYhQ7f1TDRCnKSsC0yyFHAEQeGwvBbQ9xFKlx
tLT/DyNOcT2hcMP9IOC48JJmsbQ9grNNsPP5ewtsKRwKsYkUx6gRmGYJ24AjOy6ndMYP/0wQWvxP
7W9WJDBcnK7+n2XMaTaqh+ublL4OUrJVxR16Mmh4ZwLJij1Za7XMNDbmtvPvZEnfS1lNkogV16eM
m5/r3LGIt6UV5EYQStaCMP9nMkfQmcZ+0B2LuCVQia2U4SHePuUbKGpG3mzKLlYoRUZiPaCdVH0v
/VyAiA/BytXziTUTuwkvvvyvcBwJ8T9oXtnM6A9BJrVJ65ivpodnEb5TvzxPggWg4KIcdOlWupl3
x7SJrBTW5tjyX08wz0ippnkoPRP2U3aesz/HInXx6TXNAEDVFlhU/IR4/qmHRq0H/CS0TXoaPQeM
6rVeWqHjCjKEzfCX8C2sFXP7ID0VXg+GUldfo4+HY26DYxXE6voKCvN7mTLj+uMsx2/+tWELeVqd
pvat113PKQKvb3Zzi6Dbi5+hk9dNGhLXTI64qW0NGMl6KQ72X/8UjKhmQeOqinOVh+3ZBa8/iscv
Hjf3OmaSo+YIqicbQivIdVRRZNWme64hKDf9at6MKrLq8qMpdW3U0Etzc5DOkOOW2d/WGsJtP9RI
EhdaugtQKdvFNUTcqwaScojtkQwxDicrmReU4NFaiimXfsQcX2mmkAJ7Xt4HuhWJQ1QRmnJfN7mN
gk1nxi3BeV5YMKDI1Q1aKWhMoP0LLqxRR7AwGhGdqBk/Xa5sZO3cyrUC5P4Hac9CZYv3gN15j5yB
x+KM+3v/9wRNDqufrrfTx3mcLQ0dd48vQNjPrJkXBsdRgVzIKNvQQLuAx+gUnKAR9RPIhtNH5VOi
Ukz3Q3pGLY8JkAxMdX5GfJ5sk2RysQPtLxcZ586HJcaimFBPyo9vxnhzSDp4k0wZgJBcMaPch2fy
29laJZqnzm8fUKdE2TVquUeGakeyCzXDMG6+dEitusUz8L7I7uFdG6g3d/6PdBpSRy06pc+7HYa3
IASmgHOz8BZuY7I02ARSeJzid4gB6JJLSCbuxIhqBLb9UqrtAFkJJcPeAvQET0kUz16/IHq0HXSS
9k0vgDmnSXqqZmAR2OjXHiHMVPPf7nITOFZffTadW7Ro7vszNHdHbEFVflKVpOi7XSzhnKPRlnHI
4y9NTlx1edk3vIadMMRzA91Z2m16LR2RosW457wXZz/jKv2YBGVxbyClHfVy8fnCClfKFdaAgUkX
PUOloPY6UEFxEueiiStFQ+e83/2QrINDbp1XG4KmjvmISmYMYVDIqoundD75jhhjNoXUQjGMaT4k
1kG2QwkFkrBr3NDmvtmG0Wf/HyAtC6rXleC39dCV8Qy5gaq+s3qqUawSTbmVMnHJ0ayqVFBIE+YY
R38j1sqpy8dDAKlsE/boEga+Oa7IhaZt1c4h1BcSTSXsda5L3hlciL0x3cV4SRbx50srezXahU7z
t9zeFrlY2IbxB2ZOYq/jhnlx9zVLPsLfTeX6t+33cKaKV/JmN6a3IskzPY9yTH6bIDp6jXrkiyd5
NEzwVcuhESal1Q56LmuxOUvTgaJJedzuyhvuOSlZdt0jzCLYjtq6LHd5Oi8tJjnfSLodVVjovApg
MaXj6qs2peo9Dxj5mDXvXVLqgU6xCKls0/Def86a57oB5yeqZJh/Pw9P/fJWvUgr0t5JJSzKKGCN
OBBNbRd0UbDzQ2SEvn6ItA2ukG0sRT3sKQx74cJkXhzdT+nLw240/ovIEmXyk8LY9IFNeG94xrK6
9x8uh6CvKfjfITEerNNk3IR9cXK4P4w9XFDdmGJMIzwxCn/FJ0dGtq0rDvWtAdZFiJLqcFXLePRp
Di37YA1QIjRH3zhxgsV4bfPW0kA3LvbxfFFAW6l9K0u8irxaq1ofIhVJgJnlgFUnrMfo5ho0yOp4
/UcKgZbQ3oABCF5MvyDZAyvoWdUDXtPIysJW/ZIdtqsovXy6+SK9NZA1rMatloPc0A+AMgFKGx6C
YLQ0MNyRqtJtX8rJbeoUXnnxredm/9hmWULfbm2uNXFK5EXqM5aSXCURnCf/qhhKnzhlGomcAlLx
rXPHPi0ZLyxpxbCfypwbMb/FGqh2wcMtKfI9vdviZRUpJbTtXfarUgAn7ZnpbVslABadJPSvlmPW
BZZXknCS//hVy6dAuPfnCZUaFRULArcyoNNPd0tsipBPsiiQTRrOf3SluNamZG1Xs9X7z8fkbnM3
qqg49YHOUzNFXF8z/+QmVYamTdb3wbHJaiIqetM68nEmceYc9Cg7Eb/zZ7iUblqqKrCaoyWBxJH4
j2wxGN5Wjyvz/jpunn2YD9kbrji/Z0zOau7G64nlTh/KTwmQDWXRSKkih9KHFYg0NSsLpNwf5ZTh
tW87lKoy/K5Teyx6BeuLoV6Qc5+/U/M0JoyC4898GNLbr0kN7v+o6UdogpyGLfhcpt0048LXVDPv
s+A34tkdQEeVDSFGsxiIp9YMyzeHKmR3sznLpdIx74h6BEq02pyaSD3ku7N6/Trb3HFePyAneAzL
OUvt4T3MHmoLsnDvb/9x0UwgQfZS4pQr5K/ea5R0iA7EN/NmLWXODoDogxE+WCiYkwZqZS+QzI4/
UrtUBJQEOlhLQ0QuzBWZIsGSic/jkZvLh4cH2WRkKYdjNACgkYO8Di3xk42wHv/zcdRDb6B7eA0q
3gXtaZiTMtjtfSU91avvWNe78MnROUs2yqxlewtbUVuwFwyUwbW/Vb7FPqtzELjPTVK31chIl7TB
uY34ye4TFEK8aeNtokIMgHKFp0k1ZbTcdSkaOqX9JO6sNpos8mr8+yMVk6djspnqbijDBFAeJwge
51B+TtC6o7DUtY/KE++BKraFGIX/fveZ5TSL4DEnVN8ZcS90TFLlJ1xAQTRZtvif1Bc6sT3qIWtH
N348B1c3xQJswRttyWwLwuZwiHs2zZSR6/OTSNk5TXtOLeTvppDIpnxBoRscDtVx2fwRBCHZmw8w
t5dTWP9VrT+TnNhszD1CAxiB0LgrAbHwMXwuWoGsiF2OGZzLGx9m5eZswu9/Ro1gVqaeXh6TQ6VE
5j/tNxpvxwnrhO58nBB5QIkKcPpH05UVvR1CQcU3IEDUEBTsO33NthOsK0sTRBjsJml0ft1DLgDE
1sXoR/QjMO8JSCHz6sffcx6bJkwO9ocWwFNpaAwR5nb85Y80uAvsEQDirLiFvm0odrCnhn0tZBer
amTEuXR5eEJOiTBLNY8UzWsUt188Z5Pi4QUADcc8pOcxn88hLyPAnndWaF5upzw95TZyB1sfoO9h
f+uq9UsVUcpjvMui9jbeiqP5jqSTEeqnNZ7BzaN1ZevogL9s3pU52XYcXJBRq0/YD++Hy5/Cae1r
mBZFqu0LOxcQj7nP9ItEIGWZ109otsE0dnlnqZqNLuyArcobA3f3n4O4LaXrtx2NuILZxKPqC6bM
AE7/LUQTSTYIgCtrpU+qiNh4yuQB64+3ldLXwOahX1fVfs8y4eabT9MELAwX7NzUyoMGalDltKOI
GSj+hzQVxswwvPMCJ154OZJviBXSv1IbcQ0ISycc5EEax3VN5+ELxFRLH8aGZAO1dFX5LFSfTTjc
mGmhlnKzNV9nz0pqQ0wCrY38jLmvlgpb3+cqllvPdi4l0H5SgUjrPZyHXUBS7RivPlCpYEbbWr03
5+7wYDyyWe1jKeqb24pEP9GkV+4tH+a6TJbcQGRmTH9P/wzbrEWhw1sYNhUP04m+KoMjWHEwttEg
avWdjeq6Jzuc8u4dY7t4Yl4yaq/OLx3j6R5xGH0TUsnant69BpxCrPDk193CbTxSgft3ui6emBxt
aaxRm1gRO+C3V2ET46N6+q8etH6wUKkPZtIxRyFL0ntJKFGdfZhnr8cvpOVeggnGuOM2y7grnD0Y
HzVeqS+nnueFjSDjdZEjcVMFni+gPM6eEQ03xzAO84YdstEQMGMCSUgC5DmgsoLPE5eawo+YQrWg
Gs6y55KVc0olS+po2H78zJ+pXEdCPb+ZhFJOzuT4ZYvk+YXnVXaYLPnNRIez55jK8uOSJRQ1EbtJ
Sg8bHS+RdYp2PRambB9f0N5Xr8LZUkUTs1SUgS9SLRMh8YCaqhMDibVU9jsHf4hPj1K7H2DUiAoW
JyNMxTDMR51OaTutrKVGU33byDjjATn72PGMdZkI3oHdE5xcSS/zftieoHlpT2+E3GX4rU/cnxtq
2noRCxJigrsiXacC5QDqzt0mmX4vBYHUmoYLi5Gcp2Jmnbq3o2tXKJfWfqACZUAnH24e45VN2RUU
SaqYyC1v/y9nuV1RTDEZyGkoy4BMops51P/RY9v0YhgrQxi49DBgUkmsCgCiWK+qTYVWcPCsb6wD
x1gjmf3A1ie/4TPRcY5+HZEWEuL3JXAi2sm3bEUZ0BFvQslV/dm2JmjYvhY1vWAMZLllS6xGtwct
4SExDv5LDF3wKwzySIrR8tszp+t484THa3KSONrKHiKDvmLg8PQHcuLCSS1avjqbbvSSh3HWc2xA
vr4WsJ1p9QC22hN8Je8XMnYLZiYLYdfrECF6dkhus4vm7SNl4sAynpEbn+X3Mn+nfrOvCowULYWU
Q6b7NU5Pz0sTPAjUqudu8ng7BJNZ54SDCWbtrd9iEpcb+6HkplGKOcrJVCIcQ3cYVYGSG17+HV43
yI18ioQnT2T9AwcyRv3vA/xa46swwcGjFocU+8vW7u/yPFfZr/PUl9HZCZ4xlln3rxGsKSWZbpfP
WnEgalNeojeXfPyDWufKI5u9XZp8Q4UiUa5OX6KGseNEim0RBZNOCgpj7rkI0EqcRlhf/WTaaSoX
zWHfp31VYIBAQJrR7hVYvXz+atHG5CP0LHX+3E6BJkGpIKAPiyUx05pc2v9WEJ5re7IXDoydjRhb
cvQ/gUhD7Tl/sHJLwnkL29Fk2Y8E6jA0GGuqPX9wUcsSlfhOaUEzq0lu6dLk4aVG02T592rAVs+P
obLYkCRoQ3kmY5d33r6rZcG/RVYxyddfVj1A/bafuYm7rxAR9hX/da6rjQolnLJciFpVrPU5BHu3
6lJCPogZs5hZ76rmNI+HLRX0qS9+oGwW3Xy92utifp9fm3Lewz5kdl0GXbPS2G11RJFb7KUZs9QH
oS7d8Z9FRTTKv8dhqZ68yqltfyZoxf/g73ynzYPQS2wRmEnSsY1cSHYL8gK9KQB5BrRHKeK+LAB5
vS+zBipm3NsiuKStD/WkE02QwzveOy2Yk/AI5Olf1OMo1+k2tKdq1JNSUURtdze804ZZvkretum5
3sODOjBfkOduapiwU4gsfS/cGXXfLBgQbcHbqJEDI3Wj5txguWK3WE2J9sESsObM08F8VKGt7691
4bN8S8gXVhhbUnGfV6LhICawVJKk6QutTI7baFxSBc445xhweLsJ4hUvUtehmeG/9ZAyE7W+7tqs
NyCVibj1dpYeZf7o7YIVPvBG6VRGbR8isKbS1DOkn+AuLfskxu5u3AOF2g69hcKIEBnlkkNPZpUB
drCwYvxDe+J+iqwQs1BQYktrQNNiamOdgyoOpkMmugTIugCNcpXswv28GpYHAgqalGP+Qat+08px
fV0dO3AF0lci6urDTOWE/5zIhTuyeuWLOSmmE7SRytOntK6RDfdycKMle8d2A5UEX7MWTlRhS+uR
4nTOeg9acbho09y3kEfxaSBC8LXQ16abNR3uLTuODOSo8DVV8mkuwGiuvea6MIYL0IV4oh+DxCo6
OpnCRxu79mATE/yRdqdmNg1srVMcDuQ1o15IaYOvNWdss/r88KIusTLGnDjE8C1hEd6IpfTo+pv6
UpqjjJ7ufHixBN6WKNKe2eXgmrhnRYc0JoVtHfEPDnmrnn6s0dkyW0Vy3vP37bi1SdXkdGCr90LL
WSoRoZmbln2SaBcjHvcel8PwVXTepBkaX5VrMBO9vDwiNamlz8kRHz7lvc/fGGAIFW3geOc+kAUo
aA3tcMYsbh8FzrhCY1OASlqSCDvsYLvTG7/olUFcFLpA5KlX8dSyWfJFrxGKd3rR7Ls0LfJyhQua
TFCDZP1WFsXLP6w2dkNgVpD/nGO8Oo/BYChFm6PBQ3kiHdi87yncaixJpdGKqEHN6LBnzQWw05/R
Zgc8wkCPTWjo7f76fD1m4dXchp++W7DWFGcOsTen/GXlYwcc/HVIjn7iHCCZgX4kJKOLs924tIKC
o/+qtpHD06jti22zxC25e8R7NU6iS1jzBHOHIcyAgiNDrQu/nlw4CKtLW1/+kzGQLmjEJ9L0MhgL
y0wZZ5/gzZs9hNXO6s8rmgMP8tEpkkGuXb55NFUEnZzdl4YlIy+yDfwlvrZdhCHFuSIHk67VvjFg
WPKn9EPSfNYq0QgPAV/A0abaqPQCDn6T/NcXojG3fyzyHbdQlWhDJ9V7qlYpURvkl9rSgGm40DY0
YbuHVzbJ87z4D6fdBpu9aaq2TAzAIo3W9uhRmNUf/+TytXjq9jy0E6Y2PHUboCJlou+vtrjrYhTn
gxcm9/QuWi9gGFZZ53H1Zo3QW8u+vrXHtmbf7FEhny7j4/Rl4KegqAa0JkVY59m4a/5giSgaI05x
LGHrkKNiEoSh1C5krwm/qnrDJpHcwcws6oPGbemttl1RJ1Wx75VYSYnTLl3hwLZnIfqpkEWmdZ7t
wYnG7BZZ+wPdtKu7RtcygRDA8IA2FMW8MT90H2yLRsUat54inBA1NYeVW8/q3KoCrZ4dMTAvHQMX
fCRG403cUfjAjPqma4HKSJHQqeYl8ZHXnKoRN7aa+5lo8vK70lVQE+iqsNZXfDFaQNyk40MyJVwI
VO7T7TukuFT47fW1PbvsVXif/Lnu5y6GZHV9sY9YdoEJrDj2yBrz2dYa5TKRAEVDdVVI4/moDQhZ
Slt0iD9skrseT3/WbqQgn99njwJTLdavw1s0ky718GOrl5JSXGpWn899EMYrod4HIAyiVxa0N4YZ
mR5hmESKANaWzI/RX8lJq4atBuqvVZigHk1CPM5vXHU4yvRvhm67zFaAqKXorsU33dRBiemyDpfH
gLW3T2ke1/Tq0Va4f073GoxDIwtxw7QIXbWvaYmsiAI38/st3ymlvbMQCspX9/Brdq4DwWKuNJ9R
PQQZBYHmmwph7XE09wiQVMivOOTdkTWLkd+6tNpc/Xv6mQB3HwESi2UiJbLuFnytn9PRJJgshxYD
c2uRjpkpCvZ+QVVxBakrB1TQro000dgOTXkSPPzxsln8HrquP7GZeuyDbiRZdrYpSFfmxON+UxdU
VNCXHOegSnSdkBTiBEJVB3sn2QjcQXyfKWMsw0A6mr00sWsyhXhUKAAKKx2Veg9OEsZ0Zwmf2tHG
/G8nsdt3thi5aUlQnZAcA3sPsE3Ez/ceS1duiZYflELOdm/RsulphKw/cdmko58nVGqs1jwVgVve
MiJKZVQvFQ4SEoepFc3rZ/fVRHpeLixa/TZ7kWdkc+kibUNPIimeXoMhjvrxaFszb/kyLr2GKNXa
pqmANjwRTb+jNogg0P2GulC2d46aC2+kP9AQXGdM/owFyEWfy2+8c12Ixr7Hn6I6bR4eaSwxLp7a
v/93RBZT3p5bfSnqxF6T/4swv13bM/YlNspfQN1d9uDaS6Puoeiu7c7YrGJtVMh+XUsH1ywLMt37
hc9WxDtydV0HAPpD9lTwVAWKL6UfVA3FKYrprhvd5xTIdOoE8PnNG21k7FlEE6vy3UGguxLZVCiB
BDyiVN4VRzx6UHwBnKBya0kfWuZyQwrzXPa8a29I5kIp3npE98CZOANpXTZ4WoOuVOz7/J/w9IBn
OF5bFCehD/pqA8f2K/Wr5mXxjXGg54q909heH07V4CVYXYDBFw4krQYhP3/eumbpNWvst9n1quN1
Ag1eAsHqGSuSGl/GSdfyXrqdVgoVzQBmirv+3C01AOQ5Ph48p8m33NAM1uowpJwsEA7o58mXnAzD
od+krpeG4ojepH/y5eNpnz7Hhtf90UaT+4MDW5kE3BwbfdZP+ZiWgP7Jgl2HLY9jy7bErKXH4IHE
58dQc9i66bbdXxHAvxJ+7Fpf6V6BXRG9AEMSdxBVK8WwL4YoXxnzYmTPxxyy+9Bgu82kRgWDprlR
WTi3zG59ei3wjbGWR5eow370mFqvde5mFEyYoLXHeGqevJCM2RYIOtsY2M7oueJQEkFhODGN/Bq0
QtfQg84RqVkHJHiIl9MOUWkwZi/QjqG13D6/79nKhU4t/j8iVDvJZlo8iSu04jtpwNYG49vC8jJo
uOSBx+4ihLc6i3/8Q18ZN1Em9iMq4wnNSs+UbEERXtrRBQkcJgWhRJMpKr5pP4u8nItK9rYf8aLr
oZllG5rQMoY9tCip0K3AL62Z8QpNR+mwShY/3FeV7TiPR+WXKDIAMCQv0+tl2WeAji38qy/aow7P
zidxvnnkquO+IKYxjahEpikuvy6M6Nwf53upkDaB4Ec8I5R28o5LfDHu6ZDutgbyJRDHBmzLN6Og
Ntr2m/5oDSGySz6t6qw1qRXwKOTH0l3wYW1lAotdg/7iFklqRAjW+pTuh85QNxttLq82qqMyk9E8
fHZMsoSlR9hghkaQNyOjW2Rds2xREVUHwloU8n0Jqn2bV43Xl2HLcnm6ZyTVomzru1+gg1FO/Iof
ECTUrfrWZlvgPO3qbKT4hODMIDZWpIenaSZAG4Da5476fgfyG9sVPqOqaEzGJtOv3mEyXhocw0hw
EKRHSdc/RQZBCxG+BmR2kBYHnY1BpI/JRAdzjTatJwFELJS8deuvgxG+l49LLqFtDLAHGGY/b/aQ
0xGYw3FzymO+E4bUjTuhH9vIZeH0GBrunpHmmGRtHXdGpROYHgCV41G6Hja3SRgHtzOFFgNJ5a49
SIMiDiVGGfi+Ff3LFr0FF/Atcoff2vChF/u1L84iPDmwH68ubPY9U+N1BUIFqzV+EGkGcKuLsBHC
E/GJJJb77Ob4MfTCnlH3SnBmXQYlk3MiQRb5Udhf+rx6PlISeaSEpk44aI34OLaqKKR0vM0G4dtE
Sctgij8vArfQodI2Nl/Ar3l+kCZtaAPtj+3R45ZMFup+9AkR6bSd/gzRoFXV3fxM+lOj44vkHYnU
rf4LJq+FV7r0/zZfRd/0W4dd3pnt24invxPBdQHY/atVGiPGpZnGX/HrqkvWO9usv4rAI/O0hciv
WMg1KVKUjsxLKS5JlKK0IHDYjZ3CzHBsGPbFkStHjuK8V32Ux5r+T6D13POGQIkr4tEk6gMzAacH
oYX+8tmq329lW47WKXgUNb8aX1PZKhseimzkxa9n1u6i80DIJr1pY6tvHDGRvxu7j6RQulhqHthU
ONduzIDZ1fHYNNwBGiH3WsqeHkCzlH5lr4HE/QpbpkTWUCGxY7aqREscX7JniA/MP/3Y1mxA4dZk
PUJAYzGDmfft7WJiWuBX0vv/ylcndFAw8DDPLIB9XDCrhVA8oUhfQmEFdAHjsQtgn/A/lHcUogRc
VYyLbAN8KyWW3vaKhnF4zzuCUedkWqDLzH9XdadQbYuphriTe7pCL5QPf+nuD/TmMwOlLElXkbyc
5Ye2TcIFpcJSGKkNI//ksbvb4NFbBP9dy3DcuVOc0cm4zoDH3POAaZutZQvkMraYiwLgrLv57c7T
ETZ07pn5ruEMVHnoVV0LAYFZmHCeXIo5M4gCqBOFxJ3sdmzsAlUXoG+i9kbNZzHRfkXorx6BpKHF
XTQYHGXrDOs1v9BGjPykhYqHNOhVbeT0uUN5r6Uh8fEY5+25JSMZ1x3fNJxg6ADx33F0yNZ3N3/R
F9WHYuKv/Ddtkr3x3IdLJdYDMmOKB9xA39wNH70nU0Aq/nyb4o5cwbpo4t2MyASQod9ZRPhdR2aG
bMzwCXJOR03xWqYfWhdd/jJ9JYbB09tP+vcjBOOoxEIwvNG89F7mtmt3bDIC8VKgsmukwvfmfwZh
qlkMnQFBFzkOd3YrVxAsSQODCwYIjTx5RYcsFZ8/GdTJBvvy+1gsR429TVwUsl5EnQhicJC8l8ic
1M7uN0BEIzSAab15poLrW3hktHGjYw79O6V4vIY7S5xA2hJjr2TN+OJQilnbJhLPfklY6yyNBNZY
cEd+PFkDfH3YOmHIBBdI4MyHvtCFGQrCHmAjof7MuGNDqVwbfvK7njySgtiMr2Cnl5DTVJ0bsiF2
q+RYtdJsXTmJKWmvkwpsahFUTNGDKBFeNZC/vum5p3gXynEzEyAc60+Kbkw/4e9Dsm0H5xwkVZIl
14jXpqFvy83mXYvE983MHhRBYoQUUV08u8NMbaKtii3SA6Aotrb2QLWMs92PMMzHrIUjlwWONVuG
yh14hoeHXRHScut7HEfeJ3C0bL1wErEsdm/ZbHQLKF+9yv31usJDGniBssKr/IaLJae4EutlhKXI
AYpQ4h/5xsYyw/Yf36SKQHzcPOaJk3lPDPHppGvlj/f37e3ttpDQYvV76wtllB2CA7RRX7Xjsr16
nM5PgXxxJLJjC+2dJZYS6jP86lImUzB/DvXy9/tniGb20FtjQKtyXh9I8ZH3Mfhpr7dnJzz/Mneq
4fOjAryPf03YoEjY6lk2clJuUKSMZKhPFVEUElmpI/gXY4exZtzL/gdx/kObwx91/NDhc7DZ7TXY
9JxgCCeUeOQlIemHUBYhsLTEVvJeGfkh2vYc3zN+96uuYRPOqBujDxS+HjZ6NYEd+4yOHGRZwb3H
aVPyou2QTzasnH1+p2GTArVb4xQfiYhy7Da65eBXbnGMEO0FWkHC/jhyEmG57cUTR3FvZUx1Dijr
t88ClJO1dLJAiGlgeqk3kKDruW624bqW7y4Xd+64zvwymPm4d0DiEjUFo0DYlncEuOEXehvzO0lp
sE7ljiUgkD9vFBdoXsMkIiWW7hLBhfR74JVOTmRmHllTpGejrlEYM5THrt2qIZBTvg8UWQz8LK8C
bJVoel45Pe2Ya3T2nFgVv+PLKj4Mzk+rVpol6BzmelpiVZT+gdf2iORHGLp4I/dQgfhsCSTgTe9p
zBO4nV+DwC2mOR8vxgLt4s2MY5Oi4AULKwt3QuTjCuWmwTKugWjqIag1/fUs93ledi3BghffH6LZ
u5zSB9d5ivTmsW42qW2Le3XseryCgtYhDvAcztj3j4IR6O5emaCO0PW1vlxG9WILENmB8z3TI/EB
Wnpp5UiDjtgtgPqgnioyn3CU+nIoJ1Ifl5ga0sxu8ahE935cDeKOEZeefLMARVYJSx7atjV+/DKo
wfsyz9SNvEMXoEhMHl1JA3lL/RAzK9b6D53kJyA7ZTgs0Nu1VLt43dSw095tbw4OxN3nwm+6fy4G
RqyfZR/1R46/rpDEa5mL4GiOBQKR52Sm4ZsjnG/eDE8wFjpwoHP2YppwJ3Dtp7i2oBwoS0RwLXMP
YE5IOpgymh8x/CQDpis+p6XnAlR2EaVmnV6/BG1MmI2trefk0TpS0TCXmzls8jvLmWBLDLXO9771
4PLhcOrYFSM7MVGmLqyF2tYkYUYK3QIHPzk4D9iWwB6Aq1CRiRHJAo9AkbeMoHbCUw5X+j1Bqvtm
Th8L+FfK5c0TtoNSSVcENV6L0/UxlfqVYmhqCYuBH//9ytvW/2SK9wefvu4f5J6zdjITmGQtAJDS
6C1ZwkOFw9Fq1rwCbNd78Z1CvDcTKdfailWWu7CUlOYvHsOt2Wh73p0ydz7ALIyf6PfhlJYRoL43
Mb53zxTi6aMSMwnK3B1emOSehFUqEqjxOf6PX85D+IBxbTzZRSJ+K0BnUoEuigOkGvsgKZAgIieK
kSUl0EpcvA090kLdj6toXkXxS48uXca2jwh3S46VMwpvhmokcQyH1+ReIWopMDYVqyRiVSUJ//h9
yJv12jBWzfHHgpnDyDEQeL/2CT7CcQslSZ20JgmuiZKbv8MN6ZP6PLGczTygABtltNtkWkzHH90W
tC4H2KcQhH66xgSkqaoopCTALGfzLJa+NF85BwSrA+Ww5ppzeWbgOjh0E0sehOCO1d5EHrK34sYV
FVBhcweAS4KyQfNpvHjYk+dGRvce2DhbTJmQOPCJh+7QxBRYvVJGBgF3jElQtJbb2HZ+H7a/RFcs
BNvZnBLW1pPfz5sy+CBplgA4PcYS/u377rlkbp71t0LmcJNUkeQctJEeE9mqjMYZsykj3g1w3qUY
rQ/m+AlpqBRZNltiMh0gnG5ADsUpm3nQWe8/QLp0FmrMGlb2a+hZMDKbwzqpJLHHJEQ8shDjaTY7
amf0cTIChDdpTY9pEhBNYsb89Dr4loxjOrpXFRjI/0BNmqeJWaaTMl9m240PNG7fDGlSFhTFuwqG
KwMYevk3vezBqTDX0xpNtIrqLeiWoy0Bd66TH/VTI53xPsMIBsYJKmgqn1jppZHS98yaP4qxkEG5
ISIwbIU7jd9dK2eZI04Cuhbqh6HT+o+hSr10JBLgi5UjGVvPCPy42smp9vU36YZm/az50Xwi9R6w
pBG31sQ4eCRCEtgKeU/QQ0CLyAPwLnW0xmWv3fZsYsH0MonxL6go/HE3Uxm4IMv2xbvX9g6svwFV
0ltRs/QuIwsEdft5L2r9ZdwHwxywrIg9SQ3bbyDx6aQCAAlhgXz/HZ8DyRykBd+NkAuZTm/5EmRV
ocxrOqCqXIzxfJ6rTRlAgWe0aUL+GdLdo/S+XHbr7Ktec3bWG8e0FYX5yeCAGOrLzkjM5P9jvOqo
ofZ0l8qQ+T7XclnVWTEqF0Uq99Q+YxnX9jHRk4ZbsVZsYXzgz4+6kMdAs5cgQDVEhe+p8f1Rwu6a
drTi7ItRI2npPCrLvcfZCvondAkw3ZDVuX6uGTp0ql+G4tD1oY5ODvXYG3V+uukBqtt19u5iu+Cv
idFAfmqEfEcde1Yy+1kjLe0VrBm6Wq6oqxNJFs4AZG+CtcxLwMQi5mOaojQxm3S9sZ04nV9N/fhs
jydu0zDdV56JELMJkNQuYCd6DfiljfxZVubcmmV+eUphupk7WnEo8ZyetT1F/VML7i9GhgODivo5
3iCmywtkMT4A0BHlJjdhJsESQ7fF6kcNXHfIeffaxXt4axdb3xjRzcwyyMObdKhpvF0mSl4f7t/a
y7bHC+wcz+ide82qb3CNL9s6XkaG/LD7okQdaMWQHTnfkA9NksR+jLWXBNQScGni90TEOsVXJ1Yn
K+8mnVUT3R+9YZz613rjFL6Fq0vgNfnt9XzaRdA9Mi4ukZuc1IcsfyRfAhnbADaAyW8e7Yn2NnF4
2HpyULGiO5cSljM+w84SCjAWV6bT4R9s8bI65l79ZO0bRKKN4y4Po+6Omd2IksaCw24Cg1Jgln95
Yc5lhnbnmwztKtAmMKUWa9xrYfy1X8MyJQg5pQaEZWzlPPYWdAzUvwVooFHVTvwrFE0Z8GsnaB4z
KHr4AmH1u8pICXNCDuNOt6YYJFf3G0HaXsvvyOXybOo0pXXnf43H/w9peEPWUes5xDC8U4z5Kxj6
+lJSNE8SnSemI6DvOiaHS/QV3rBIrSJWZ+ydcfovrYi3zuL7y31a8oePKd2DS7E2rnt3ivtl8e09
a7asu0wE8EcBPN27Vzr1OipaQiPZsWI2iNUiedCgtlUTPDYTLy+b+IPSK92XCbqFXQ3NSloPCbXt
nH5vZ7qoB5+jrE7gLgExvZAIx52nZRuQ2XaGz+KBOK7qWnliPaZ+f1HRSqufQzZQS+yAX4pNDfMD
ltbWGCNdzoRUrJeUWLgwga6puWL3EJNIP7vKpdko49grPLLBg9cJY847bjtJWB/MErVCov5DGa/M
H91JXoV1nXYgAW6Z9kf+YKFgSx1e27heCauDRicurzSIcgonlNisedM/iyVh32CWeEzy5M6oDslQ
sTdMvAjdHh+li8H7tQ4bp99aNWW+zcsJAx+UYbWGqpWQUdG4IgRWYToXsvjU+dmKEOYpKKYLLW49
oDHnT7HUBbYr0UAOeHSDbtevyzsoH6Pe4mX0AW7z4a94k8PIXTXLRVU2+SWf0KcHATG772Ah2TTg
Jqagpn+kACFYvvpUTNOyBX6Rh8fztkYKvRA90Dy5SMfsC7Ny9Z1x0xgGmp2KQJFDXoGk39vnmJiL
HQQIhSR/DJNTRVe7ap+9zSf0nJca9kj2bUd2aupngHrGvwpEIEoKL1kxaHDknwasTBRUdGs+Zvev
K58GCfOB7tovrEos2dh++XRx/hXHFRRaa8NbSgwEHuj0bpq4hlkYInhXHHoFtxvXC/3cKhA3TVEa
J+0ftDJ4bV/izwKtZGlu8LyEvGw5Q7XxGJ0dROYhm1eVwb5sMK0r9iMW/zDNKWt7MFy6kFoaYKTK
gaZ65mLb9FuiBlIL1vv4UVYZAMoTH5d80C51C+4RNBj1cdQT6UCUOtfOg1/+LXs6+uP4Cc+Q1Pp7
IUBQpLvuUZh3LRnuTnhPhvSqy1Z/lJPWx4IE584uXmap9iCFROl6e4ZFH5fBWdEUVXsRaUwDV03c
jYBsnpw/b+lFU5dwccjnqUgVDcVkKMn//6Y32dqTbWNXNBJSqcMSh+V+KM0gA6hCPLAtVgYPX8gC
I76AeG0tqE/IFRRTRIwBobKfL89S9Scfn8RYn9+QgPgD6vYqQfDFiKeTXUxvuGFOCmoZ0U0pIqrk
sG+SpAooXxBHKGjlJnZc5TUtXowZnmYZw6jfeOOTufzVPAmJrEjG6ahknRVgxzHF2FQeEgOOr6+v
rsmOGmiil1Re+4nYgiRZ1EMiOBV8J79yaZoFlBjMMOqjNZ5cRJkLU/4IHtqpUXml82pGrbnVSLxZ
S0QZy5tee9nYt+dHP65Ggyzbww2fBdsIMIoFaOouIaoDC+XJOLT81hjmzpVw8UW7p8VCbP/yXfXk
GE41WZ7vIRVBAq6lduf0JknOIMkZoFitnNNq7zKTe4H68qe0oVHwTLzpjlVgkee3c6fVRsTVYNzk
1o1/bf6e4aBY00B2QUw8SVUDzv/JAXK+Pvlez50rGlnWiY9WNwbR+Yd/NiF4ThA9YyMlbksjsfVV
sDEU58CKutcYfYfBexUywQvwwgg4YfTyxdreU/yFtYAtZFZl3M4mtBXj869Z7/lyotzZP3TMH2vv
3TvifQZ5QhYtqcz9EMJ3V3YA4kqU48tLVbJIVUxNXkqML8jlH/PpyxxrIEM1Ndtyrp/BGTwJvCt8
earvDbHGWW6lcs4sNpNdJinPAUpaCGh0ML80ZCd6bJ6IOidwnMD32YC7vz0pZGsaNjlj6Ou8mUcJ
BJ+CYdpAceCCN4TJE/XhatpxLgp+uqsc9l2cJ1PtfkrDY8dq9gAeiap7mhbfRHITgv5MKIebCc+T
qR1TCKjXlQ9XYp3eERcUdOUDWXq00P6tvLOMxearOfUEQZbrhb5VZF/wCt7h0cexBQTAJMpvDiI4
RR/oKyoZ09YxmlBs2mqZnOdZD59yKbl4vVdmqCVVtYIZ+8WwNHOBJJp0rCARXMrlD/KrXpkfhihd
jEMloOcuJ788Nk0VL3yuzYmNet8uxkaCuv4nqak4cz+6XVn2lHj5GFzUbleaniaDEAoACl9LqNet
bRB6JWGdoL8CAR801gM5iHwfz4VN6lKLxTPTBw90XjStg46LBJtVJahoHTv0MaUVS6K3YsYOgYfj
i3/rgvWM+6cwkTlFZp1pvA2mvrIxg8eNekJMrAfjg8ewu2BR5iusJLGPqWmIVcg/VRu5/z53oaQA
ehLP8cbqqwhfLkObNNyqWXSK7kEM8kmuo2/vIq56ftWjGZ2bxpLfLnrTG72Beyrw+Fn1m6TNiJgr
rhr8fXB+n1bEAP4WTDdgeBKNJqWkfvfXCkQaSocn28JeN7r7+Edp1XxCeo97gfdNkvUDor6ClQQI
rezunkzX0vOucs1a1R2zvlaV4mxwxF8NxptQxWQ6kCHgD59SwDOvRkX4DYoj1UVOYPNq0Em09Gq+
84FbN/2mG3ZBuQOp0XBoVIUmZbapqCYtpNFnvljK+sEwVgceawHBZb+4XLhDOi9SNdLhGhaVzi1H
tLK0uhnp0wuMcpP9aAm78oJl7WTtnhtYOZpPOq6Ozq/qveP5rl3T5ZGrOc+Bfo68e3d25nMBMqwr
JJ6a3Y3dWGe4iGSzxbUw9JE/O8nsr4Z+PyBx+0mJLu5j+bIYwjZ5kdysJC6DMtzuQcM6wOvmphRn
kAQdQmTMVIDyeTByOK4mXFmVDIrvSx1A29YSCoJm4eIWk0dCHQE+iS8ZuKNGFa4qsBdAko3NvIP5
FG8PnPGEa9bfcgxHXMTQbKxuXj2fIiT4knfMCor/IJuh9GKzmfwBEilEDx+Qi8RdjkeswRBo/WJg
5A4XVhiH7EqWQVlkam45ptW1ojNlmRscumuU5bKaWb44OM9DPhsoMD8Yl3zTboU4Jmmggp2UqGs4
y8lvOtiNt5Z7AIz8+cJ36vnjO40Ac+8+u2cdgRjbzCNIubTF59tmE3eK3lGEnmtyFDy7cIDfm8P+
SWJAj60GRq4XdSF5WCicH/fypw0DwOZHgRwIdnc2f2KoR1jYjzKfaAxynq1ICGnsyOHrb/EBZtDU
/Rah1T4bLeT/PypLsvRHw8jaHVvbTXtsJtIIcOMtnoq89ikB6JsngWGUPaeDIfEGB1lKmVb0GGbn
ZezjBj2nZ1Kk3vzVRH9gvOzseIXq5y4cnbRPGGuOjRKD+7uu0l53T95SJHt/b68yQ/itLswA3nEi
JWDwZiH2Lo4vhEwncHFglvmKu59N3uC9wpFTmLsK/u8ltCIcJ34xoVAPQ6rVaDOvTomTOi2L/YDZ
9q1p/ZAe+Tlmbx5TQmDwNwx3YIFJOq50pR98e9cMNvuNJobdvlHa8zr7nO1oFZhFJRK6ZEcRpN3n
kagjVFiptbTiATsjsur9VFmVh1N2x2AOjf0TVE0lgMI02lTVBwoNc/d7EIqT/edl9g4W0wghQlUI
2jLk7aDVG4rYVHmIkEUYCUVdo99tszGiZ0L4dt0Nh2cdVSnwoxJzJxP9ETGZmlYSjCXKd29idEAT
+jXEbJ3VTFVZsPyHSeR/HcI3rvtcNBj0mjdHblQvoE/bohLQ/A3aDXTsEj+f/cB353dR6629sARk
xw2YA3iGAqtlJl0VO23pzuBz8rnwi4+4sqd9P2iiJ3pBRHq5Vjwa7nqGWu8v/TQ6h0+VL0ZUi2bB
AbC8AjRMkifzA00DllTRCntAMCCXc76KDQgdspGLvrtUNdd0mxBrLH8WXUIqDEKj75IWlRCgWJNH
UZBer+wEpiOL0sFoMMRdkj2+QOtWUnZJI1x1ZBKv3HKY8fOG+8B2oU+rMp/wKMTtZ2YG4r8asJuQ
CfIWXi4YRfrIrfESIG1/+QMJ0djTJhyPAAJN8K/ejbdK2+Oe7okx8zC0o1DUJ7xzMk6F5EKlP4B7
jfZCdEOBuYeBqk+y5qyE+txVcy6F+CPSUkcHnXP7RyMEsCSSMpS+N0Y9xL7Maod9sHAUbT15Ukg+
ua/fF9qWUEbuTF1SleEoFg1XPhTcTb8/siSRG7K1lhR72GH595Tw311j/ypONIgttFBjEXVTfksr
ftkMu0TxCgvVDboUCxy31ToTCHbc3CmNFdmZ6UIFKJKRg9OWqa80kgbLKxPzQdSL3qM75374LtZU
lhieoKoEin+b+J175LjDOVqTUk1OpXahUXb9KwXjN9V/e6cBUty3KfJ6MUXcaT3uigeFxJd6oCFE
rF6GBhV/IBFENHblc4/0qZpdnB/Yl9t0b3GppOalcfj9GiVdrXNQBBszU3RP2h6pxs3iG3IUKykP
4JgoPEeDQhSRkGwpg2yfL/xmSM4EC/ztxBQqt1GJzZsvfDtGpqY7fQboQRkZSwR1TgKSnz+J0Lqg
SmwVdQOLJ3sIgaW/KfEmZwBSf/Vo7sUjldlaTzavBlSPHjyyRcDG6Q/Q2h8i52S/skJ9Fv1eCGT7
uCOwR3VfMSXlq2z9KuiQthk45YgY6LnNKZ5iTSh1BOcvYOOulfq/ujqhYTUbfDpMVcSfq4awNy/R
Zly6tb7a2QIsNaBFWGypMV2NKZJzUkD4GGQz2IqrONUQBAoUBh8XFsxA/KfMZn/eMgWgYGy1/QWm
Ig9A64m+Q+F36BD1A7fKDTlEgl+DMHVD0KL3DYdbIPwdOqR/ODwN0mqqRKTrC1rTPP20SCKf7gGT
5FobfMswTGaRI3y1XBQzUssver5u+CpoSU7CUJvfS/z15I4+C8l5UUS+1cB3NMJo88XBUEySW0qh
V+fVOoEaqoLILMO4BD9iBLSoF5VL324BK+5x8eUoIKMn1ngzABCGI4nkZU/Tchb1ABvEyueSGv+t
uCvT8TH/b5zbBFRsyV3d/pkg2QG0hjCKR4XRgAyOYsk/Ku387q3B4181QJa5prMvdWtHrCXRgjU8
nyCNgoDt2MLUE/i9UnjXhLCEfSQ+BZ0p0TvkXI3q4gToYEXbP/haL3XhrxunKLG8or3hmjCIo6we
spf3zdh67dUCcI5SHIYiNcBrTvQc5VneSkUt1xFs/4TC0oQAkxNqt8RQ3U08S+p+uP8cnVdNKpDo
AGKQ8FrU8jdxAfDzd2WPiGtyB+FzD+ReeFCkhcVsmQmqweLO437BBc0h4r3UZpWFIYYJhpVAjnO9
1UZ8WTBghnmWnrY5LRG8r38dkFJKdN0vSooPqjZnhccAC16zde2Nc2vNx+Vn80h3BvKANp3dUpTQ
iFMbxSKWNtCmOMTa2cGxOuGAQaemvaAbuuA+wTzB8VBCdeotbGSF/clwSmQR9Isu+IxzDtvTzraV
DzsyTvcW6JONcin/BHcdagrC+zezJR+UNTaeTkrP3MyOuJ2cDOcvMu5nCiMY7hPPHyNV8kGX24js
ULEdAUXT42FFstRudlK6f1WyyRyZZ89zwS1JuRBv9AoMGvH7aBtabQrEi8txKubp2Wmdus57xrkp
UaZQrScEJsDffvQZOWZ6CqzY29e881L/H8KHFNwwhwxcWtuan+Mgo25vi2U/LLDy4zSDxlwq32no
AQUShMU5lZ9+PM/MlVXs2BhCZDIiWzz4yPQoWF43WWuRFMWLc/tpeUZWNceWM075I0vXIQayqMAW
JTN82c21LzLmH401jo8+eoO4u6MM2WrUNnVCMjx6LSfWZyZ/Rc3Dr5T+8FIx8fmQsjFGj1RZW5NX
WYlrmf8/5EtH+rnSoL3LYAsheWnJr03N0sBks54ITxErsOK1rmaoX296xoUd1amDEzkto25/NO+v
iNesds4phCvjdGEwUDqiujCvQ3h1kUJ07mUSeCOlVRKueggy8Jttrw7fKuwQ/9ajgJOkCj4r1HLN
joeG7nBgxEngl3V4aGx4zg65QKwkv0umhf5XcbzXPiX/jjn1ftOomTe3CKg6rdTUBOSApcGm9joQ
/XLXse7zaNHK4pLppvWeVAuobfc8doUpChpKKjn6mJUpbip8HmnQVgo1CxGlBxbJ/vBbAkIOqC90
btFzQpxcK5efwF4S/3FyYB8KjklFfpSSV6sRwskSVd84kkm99sSO8y3M733H63904mE0J7jJ8Jhi
dqAZG1pkXmbqI6ENKtJPXHrTp80MzbDDUcYqCOD6p8RoeBv1dHy5WdUoHWFfw7WJjHHKU01chEzh
4f6sJRECWGqU/kcRPGwI5rVt2qaPvEWosVksfYwhyBTgabByUSmviADux4F7Aev+iwMaYxkb86ZA
rqmWIPqSZ8gaSAIS663ijpIKDRJzkuLI3wAeVKm6VHYL75C3iei84FcwvCmkn4zLQ0E3H9143ULZ
zjJUd7mAuEPvKj5OtR1n+w1+UNgJfZ50aLqJoVSu0b0ASSOa6xSvMqYTS6xNlM/pOLSg0PUidi34
KWww09VcfKpSlsgrs11xJO/d0RttdAPd2yPkM1vtVj2kdUaQzS4dLeHcgENOhbfEvo2tyMxiAbZz
A2kdTShZilJBq5XSn8MYDhdUHn/TE3x11JFBxa17zBrZgU4yvyweoTMsO+RZo9eS/wa+T46f85AW
3kPBoT5GkTnwozQ4J6f0zQyaeae0KP66ynZLxGHCBMmB0SdaVjdloZ2EDW3N8c+xf16qOZ7ZsWWs
BOKsGgUY7bNNkfKcWtu+TfUzCZ8QI8dG7Uz2OEoDRF4SYzrxJbaKHSQWAEg5igeDpr7/T849n10J
iQFgeCIHcJEW/aQghvlcPpveUFgNjoVJjDGQmEsEKvRbOVb3tW//jcq/DM6HKFACwKLNJjxz8brq
OgVsOxiKOHU/jKcDjiZuRRYh5AKsf/MDWzdqVpTDXnBfU1uyflVu+rXTWICnumiV22HfK+DTSztp
gAW1BzK2TsS3tYC6Jnq59FcPsb8+V6UMS6Ec9qtr76tWb2PugqBPOynlmU42fD7vP9XS6CHWvDZh
18c4U8CKjC/7EtZrbADW/1zwyxe/dvR56vsfGC2IG2Yllqa+ebkl00r/LfRs7mzrbmwzx00lO0mm
O0PqrJqnIqEqZ4ChMafqn/rTbcQyBdIhqhiu4tOhsnZ8oo5MdTKn0m7zjpoJn4tXWBqlYa+32RxH
QUGfVwpU/l0Or5d1IAUMWqDjGCVfYtBqmxiEwgYPl2gtqrd2YcvlS+7/3PyoD2W9ZRx96prHAV+6
1fcZZSwgp8A6TSctwo3O6QNP20NdJl42djBei7PDfK13qMlhbaI/QVDEeY4Lsu/HxaJHJOgo2D40
DuXj4QBmiTKcJeYhC8vBoV43NcxU7PsZ0yt0WU8c6W9KmMYKoiC+W4UlkEZziQ/oF6v+5XxyUgkf
4VG16yLFK7/otIsS+t8dEVntmpWzj/ZThL8DQRmO5NiZ4lIbxWmLXGqaT+MANeHffyEYYXXBTAuf
GnGn2CJIwLErnd0A4eJ11grijzEPSN0H8mALq7OgAjHXyXQC/vZleImBZ3TR0r7v2RgDu7l3f49R
RmccedIMS9sjS0AIxzuSqg1G6RsB9xl7YUsyZmXUeZIMWagsZxx8TYFJdmgFgQq95kGD0orFQNX8
c17K43mnbWeb9xVUQtC2viZ68yFsGHSNI+3MrlIq1V8t47HHYgJIxrFlLFR8qraqBWJCpH5smxVG
09EsSvMcNFwOCeZR97wdWnbEcaiPB3kqFL2fiIDY/y+R9adyB93hQwoRaCx4GR/DK2Q9KKJC+Cus
Chi9ohaudyP8tt0TSOcrS0IrZpzEfVWTrUVuTYMIbTRr9pyeeR7T0btEKgkvxzlVzly1hWinAuFU
kaumJi0EaI86Oc1tD2Mtns94c5E3xSDcaZPy+jBYreJgrRFLO4tWnnYFhZ4V2PVn0LL5ckUzdPHI
2Nm2KA4wfiIuF/twLGdjhio9U3qX3HThgUSLLvRRBQDkp4OdLaXQIlMErMXpQ6iur6P8EiDv65sn
rMtVh7p4FWFkoCn3dZxvppidCGORp9U58OhTj2blj/xf+A2Z3Yzj6M8ybzza3/9Za9PvsF5kwEDF
UayteEyWH7EmYmDrJgfqP0/oCMk/ghY9sUCXQp0wSEb66iqynEzNOhlDbHOjKbs7R9KmUcJmTSyy
cxpFsaMXpB6WUdfrd29tTZTYC9YE8vLanoHROg9yN349iAxrVucAhxQ+c2I9JEMhDZvC7mTLwAw+
sYefs9yTB0KC7BaoaWXxchy0bj93NvXPtT65mPQJOGjXITGMGMHKRFBbh7gwXBgV3r0jFKD2ASn/
pg05g/exq9YvQLMoCKE7qkIvm2RonKyioVX5Uh/a8N1fMt6pT+2kHArGkzZuZY9P0ZMcwd+Qt3LY
QreqqkYrJpXvpcMRSUcKiuoXorG3unyVxMRC+iCxT6hEj7Ui+cWgJYYDN2OYRC5NGDpipFjv6vuq
nftiLzptcbHl2Q0UzCqhQ18mDQCcjX4xf//jj/q+5wHHWwdrRUm7nKBtsyPgh8YWsK6p1R8oIEUe
P2DcxHIgh8gbcw91ME4C1ypscHIr4aLmc0M7fqf5Mu5ZX96H4Cq9XYVLKQQ3W48CSEbjX4V99G+Q
AhiamAgWYfzvqgwFI1b9x3rRgGn5/5dKZu1Bv7EtLsQC3PhN2YL53AtWlq14/Yn0j8qEHkgwXBMz
HXNU/KdeF4T43qIWoskgOM9WjSDePxbMw9obsSSRVeVaiitgmiRYjoi5+ZviT6tT+l2Edb/4heQ9
xoAZ6MV3bolU+i2eMp8nTJfmjclu1Xs08t8xD9g/1phFhcOfJ0zgkyC9ZfezxBB71cjFwyq3kxlp
uOEQWZCTQnqFdS8Ufti1KfWnULWJB/u+W5QaDhBCm5I08xFSrM+mJK5D4++xW3CZ5ICOkiOMtRfj
YLgj+9zNmoq6ap4HZSeFFVhp6Uu5HY9BXC8ahxiEiqSU5cMwhC0/FSlfKs5aID07ImHEMElXl+Pp
KrcVtRTur2LCeNy4SEHV4Ab/PC7Vos8R7z0vDiC0CnGXzyxv8Y525V40U7wGx9qZRujz7FDirsO6
VD+7htxQlxiWLJ6ZGaZOEAA7K2OLSKeQKY8RHG1po3EdDWsR6wqmsWS33Uo+OYuxDt5UBy8HHlJv
hIv99kE+Wp0c31XL6LLHYHgTFToLVft7VLKV+4y8rRTbpQRvL36/eOEbsohCFSAhatknwwFJM8d1
xZRx+Cbb5MdMFtzWWe8McLS0s2sMlTrvoHejepTIFQYx2gxPwmnDl2X0EcTja/wkN2V6ydGXW7ih
wcLbRDIQIGdAjbjAWlRxAK1yB+Tq4cdon5df7JSUpj3sYZuBywggzd9vA43ANJfyPdBEJcq4IBwk
078zXGK1+uExdjI1Eqp9zW/frhUdlkUSgkfCAMwTW40F55vDnyXa+MbTdnt2epEQym4FPVnQCNAK
O+VYz+C2b5GkZsPnVHhP5lpGoB3tpC87PY6NwFkPnPFby4b08M9LhdRyw6rvIbCb5PrZafROempb
fI9TEloBEND4K8cqjXiJLqo8QUrkMjFs/Jc4fd9nmfDk1+0+4MQZ9UsGks+WUPz1FcHQp15uIGmU
ig0W806Ww6L+7f41z9UY16HvPeePtceneXYAmuHQfjVho4YSq5BjRkJ4m5Fm17AUzWJgaYdZT7tQ
Xs50QUo7HNS+9NOCtz+NSvL6SKH+INEy6EY1kJXwyZYoBykcOpmylc0SQWw+KSnEjJa6hYXIMHjY
e9BaqgcrOosAn67hCIQKe178JbFIeKzdz8FsvR7W++fOBzRpdb+GaE93ZUfMaiMkMyZen5eyxjoE
uTCKzWojMKlsgOQNTXaaAFuhLgPIK1sdqv7ufHir2tT0c8BE1QZAoi8gNY1CLgcJUjVHU2hbdSS7
z2XJcZcXU5ZJhtBcELgW/G0LydlrygCNVCaMoiFq31nqY06DqKzR6txihk5A1Qqo67vjBcf2e0L5
1fNh1EzYyc+jh7fzyble60YBa6y+zGAE95vP7YCxvYPTyPSvS5ekvtZ2E/HyKdf0Fj931Bp/TOSt
QLMloFSqSG5P1DRygz9G3vTYJ4cGEJzfhu+8UJMUlCsd1kFntt48olkQxeXylSUucE7uOhSAjFH2
tmchtHvFQhrJTKYxUwfvsJ2Tf2ro799Yylaoi518G30ggXQoasJdAKvDu9w0ERwYElr/ck0zJt18
hA2TvY5/6sDbO6wpUijn6tXgasMXqPQixgwP6CpmXox5lSaQ7c1vJFuSNoO3UFCUh3QHq5gs6A5Q
pplEkSTL9zcyi0rI9u8pxaRQFuSG84FLXyDaC7MTfn3IK6Fg0I9tbwxBoHZ/xJbosGTXMoSqfUIi
WX/+I6zaihkXBpmvB2XHgbXcBMziRRn0ByDFW+kgkHu65KYX/Q6C4Lm5EJ/GHYx1PBp0N113ZSIX
He0acUTltt66p16d39dNGZdnnUeuh45fhO69ukIMx1d9mfqlMa4nWP7kL4PmE5/Gpnnhn9oh1fJd
s/CF3P6+gjvg/bKMjUtWFAeT4mHNofs6zdAcO/fhNS3JKJ5XsgnZRifqWydL8N6ESqEcMN3pfIxu
jIJcL/LBd/J0yJ1QBJifNr/pGuJbNbjQA1jpX3cl5RaU8dgtrf7D7tws2eQSa0RCUKy87FTqLNda
6Vi2M59AveM9y64X+/T5OpJLwrLtgnVwUWDTmhwSW7RTqf8RMAje4yB/olfeC/YHEdFA334+HJKT
+c8jc7PGHWLC2Nuuu/lrcfTLsh8U83aCrj6Ii1u8dFxH+Brx+Mq630sqGEqVqlBBboOB1G4lTJ70
kCtuhEGoM9V/wWGuNbP6zWj2fnKeT7jLDUG6NGMKkyfODx8h20iUwKPtft3C9J3vS0PJfe/9e3nv
XiSTT/4zpVO4ryCahaRvkFh2vc7YWH9Uau3Dy1Et03MAf06YnmaRVw79PIIRnBxxkX8mjLr3Jeyx
PuH17TUQlMtOj3VCNTXQswbKkqoL9VFo4KkfCPLSOqQ10ACCal/ZGtdc/kVQOm6hsf3+hGWwj4ea
eRMAuXk0bwSamuBHVKM8YxwDrT1x/a1Ssr90CE1eWJZAyxlsTPbg1+rwPpWq7KvAiGqYGXkDSVF4
eAzZxc0Ev5I07Jg9p+gY3iUqZgIuBM2/UtR7zkBDUt60pSZ5Efg9pGq242ackUuhouTftyFU3ySS
VFwGqACd26iX+HZrbUksTl25y8DyFxu5AzTMtkFhOSSTPZAfY+fgD6lVE9eqqjJKFmBSe69UxAO2
lXA4SJJan+qlLkjZR+K0w01F3pVfhTAQ6HiuJiP+LrUGb26bcJf7Ns5EwiTFeu5tj3mh6OzFYI9F
3Pnc+LB+uUFaeRy5Wj+KN1+2lLhHJHY1fkcq2mAVxiipV76NmqYxYngiE0DgEbX5BtxdDCnUZbnp
uOguRz5rafjMwtneCoM6IfD4lUChoX2NuvdPtDuDuPJCsPecL4plD8uWvmpA4azO02GKP4M4cqHq
MtKtZiLlgk/7/f7xP/hqsnCjrW9schcGyvvVJ9njhNYbSdB74To/XWxJoQGZNM5+rBeHNYfqUN/c
KJFQI5BDA7IimkTRprG7yhGdwso2R1obUTe4PfnnqD3FKw2ZD4w/fa7LMV4WHKmLp0NLCj7voNJm
FRogSwQjMAG69gCkHGfq2w5gXMcqVgwfnIGs8ogcC6jjaai04/RtE3dLQ3fZg1zzhnwcEI1LfVmM
uNO6YaqB9IoyqVzhWVXamxzagggxT4YsJ1+IOlLHyqqoBj29uUEyKx1xFo/LDGHMXIakndDHwQYx
TZfBFx7ouQUjYaF+3bqMMzCNYmfKyTDlnHJ7U+MNa5NuvRCgTnZLt+nhtAdLINyrMLDsnc+plSu1
XghvScVu+ozPYpw8Db+9c9AFOombGyderlMIwQ9FnMKjxGdfgUDJh+l2o3rSDUlAE7iMX8xrm5rB
bHWBHvm1Ptb+ch16cwxGTCSKCpitHizROOmNr42uRcZiQVXxctbT+E/vvIO/IeCqs5Lqz2QkbrTu
r2PJqIFKWl8w9jrouaPi3mNHTZSIf2PuMernThSK72GjNjFsdadTfLnR8u+dcnuuhXyGzKO0/8MQ
yHRoiMIhAoEuoOFO0aTP3Ne6L0K+N6d4GZtiStQv6svDwCLfPkacaPZlI9gtrAs1/rYW5ou2Iswj
UFbXWR3phzUcad5NVbqU5DMzFCGoau0yABPjwfWWRmRzJppigYRcaSAbtjxLCuQShqVF1aM81uOT
dYGdcUrEXwYspENs6Aw/S28ii0rpPv1F1cW3sUN1J5luzi0ZWw3Hqs7zm32xwL5wRhTSZyD56W+a
YBgXf0EsMfBGKEhsHZSumZ+IeO4BuarhrlQt2H6YeyytiLFneDDG1RGL2+zp1pAATZXgRyqYAoje
hOhxZrPgh2OkIQwMHcpc9iekuRYfElgcD19diYV9701LgMIceC+Z/t+rsOkkzRWua2WmBgDTopUv
vPlVpcK7PaE0RclBEKUmVUsz0Wsee4MmNro+CMgKJUnlCCgAvVsz0rcwfG/wsDZN9ts1XeFCPfRs
HZ8r8YewhZiX++o/OKylYfN4Ii5kHgRVMqdw6oOCu6z5Evi1Wk9ppv1v1VjEvvAhLVJKk9GO4yuK
vM9Fx7myo44CgLi6IAoQdj+5LS5Rn5i1LGeTXisHYJ0zcgowVWGhDx01FmhwHc37rHhhB1EH72m8
8qsQ2e/hdRQyBwxdAaDpQjuWBsg15TutIOqnZGjv60oW+Ve+EOFG8//+AA02CzbBKlqn9t5XGpH0
jiLbper0uUn8DzDAfM7g+soxLjJDf0ZAdHD4+yk9wwLtf5MJmY7kAcOWAVQ/G+2kQNT4ihqZc0Ft
ceHs4aExmhXK23Fr/CqCOT07Hl+q3ywCkaEsDX/VLMlsmX4lJfo/Ufek7Eiib2F8qp+dLNnAf+FD
fDpKLQO1FN3HeVYThRnVGY7Vh9SyfvhLVH1d7G1REEUK89U+UHEmlKN3zQfDKHSSLqM0apOONkaw
lJTOrx2zgFJaFnufYgmTSqzEj5QRmyNimgyPPB4N8ET4MtR22HxBzHo44STE2wf/uRFerl/QW/o/
+kTPpzeKCr+19z1DX1rpfls1gmzLeuqyjDmwJxBwrVxoO52Ss0R2d+K2hIMpBQ5w+7sfmmtcXxuU
IjyIGgxNvitADJy7338snGn0OFbOzUVPsc6wGG2c1psZs+NWckmEjHKIPQHZZOZpFR9oF1qkQsSu
eYdhzpxtvQAm2ur8kxWV36rS5IGDGTEYDYMZI4J1jXLgtEK3v2a8Adt4ioijQoCRjR5j+loCTfbm
13KlqMNsQUICEl3kMQK+bHtzzwFmFoVKmI1RcD2V9hZkHB83o53WMywfpm0UsPrkUCoABD94RbQf
JiKbhpBgENe4r0lP1g6y28EQ6Pzg0UCkTRUliFIu/hNxCX+rOy7/qc3G6/R+T1kZJZDjS3D/Gj2d
crYt5m7kLymn06/ZmXeVqHIbELTB6qjXUAfmwOE8RnuwSdkwViQEnjRrCeEGS+eP+xh7mideWZay
4f1Ve1qVxJEK3WKS9heVIetiq/jGf6ogUIW/BsrrBAXXDtAwlXNxmtygR0LTDsTk9Y5+gHPLh/TY
idj9mVtFJ4PGOU0ALwpXmJ/43wspwt1LHAfIhf3glSxNONGPOaIVdrMR0L5iaOl0/tGT5rEmG7Gi
KUgZkBb+K80CKRiP2R6+KjADkDDia/3tQOP5bnFByNll2AuD0jYat+dYd2LAzPbLpZEwq1BOvYQO
wiVA1MnvIcG3M6+7JtxPEj3im0tZghyt7OZsFqT8Nj0l0LSmpSyQBcJLZnX9Ta/9a+muGfBkKsoR
nzfvp2XuAtdHX6UabF2m5uYM45iVPk7Lf/YNJdwO5zB8tTxCOiM/Kdj++DtvM4OaC1FJBcmo1wP8
o5H4GMUBRRATu4THEkiFRIhLG54PB/ajBIen+8btZTH+h/rnJI3mKG2sIhY9UpDMzgqCdElDxmvH
EBjVLbsrJfLwsqjbJrvVeO37lBhgDBsT8aFeTMlFmJJ1D9vlRBKHVgIKaZoQmFTGZ+FEhVGGOJrL
rSZ+GwHyokJqBlvC1WU0IUiOES3tw/n4PzwrIVGHdv65P2vElJUN/0dRYRPGemmVHlq6SRdcYXkx
eYJ3gvs/j6jldwA8/2WVoxTUneveyjYpW78Q2JCX01UWywkw/D7Pal4c+G/OeCIGDSu0nQuEs+hO
rNvBOCrBEtCSDygl2S1ynT55hLpTB+GXjwwsyaP41SyQrWrwu1sreQVYM7tb6ADfAObjqu45zQC+
wEAcHSBXoTogM2NzNY4YGT1/AqeERYpgVTtPiA8fHKNd8XC+IAdkUQJBM0FRMcCRfkG/N4L2oKP4
POKYAGw8sDgbVSstWvfci81INwlVUImtG8XXS+zNCbWdSeAufckSvKyruzNv3RrV5MOJXJfZldem
R/uQxlP/RnnDFnY+dXE5OCZUDGvur0vYBXtVXl3o/1YrcoVpspoeAyMdMe8BjTdub+g9aMrVvOQ/
fWNFAOyUbWUXOIPkxikaeNGs+J8KPP1swzlS25x07xWVYW1hSSx8O4Gry4I4+mpyJV2jIX4BY6SY
tYeFcZ8sLN60oUMC0fnHBzPmOkRHQMbiROqUQBaT7ui4m2gRm3EAxEEZGqSkLYenSJkae+CnQ1/N
JV+RJ4SX48VndFLFBRjTOo75GgeYlQPC/Sxo7pObn1GIEzVfxtOnW0/s0Brir9RJSvrHenMLy1ap
owqJqLox+6D65SxIGGRt9H4YxKwuBjcWLtDd8gNyy6W7z6V7HKNXVrT7xYze722vc5v2225xpKeU
uqkHL1MENJysYx/TMlgexMrHUYqsnhk98Xvm3OFPGJEwkdiN3eWSZ+3tZMPEdHCBT7chxZSr76U8
/o6H34hf0KLCgRZN7bJt8B/tVeHbeR8/4hn6eSmRW5lAuSMkw1SbJUcKnK8kBy4dkHdX1Ojek8Ku
Y8f5iPTIpyzaCq8nZNB4FLgo2gqR5EXFCNmNHzQt3OGlt/8+Zd4pdZqjKk47XWGhgnN+e1h+GTcE
xngC2HTsPC2Wt3GM5R6hjokgpeMZAEdE8yGkCyj0KkNDiym2qYEspbdFCvzIt0Atz2OSyrrIu41Z
rFMibK5xwAONfstH+WNszOgCXWA6YNWOkHw71tM3fkXYyhEKkduEY07JL7e+Ul1UTUjclgOZFPav
gVFp6AKXAbgVjAT8gWAQE19ecgREfabsdu67QZ7KQieONw52yoA68C/dCwen9Fh4pNUfNKEoQv/+
pzmVNdiAjtZHyqVMdcdYcr279YnZ3SR3AGv0OX75bsqM0Cumr4jvKoaXFjbpSd0lVKsKQ5l55s7j
Dxf8T+LXtIUJhMyCeVGgIf0LzrGp9GzzGmhF1FxVjt2qypDtNabkTnl+5fXUlC/Pm9panmgfqz21
i2mgAasa7lmcSI1LBLyZjsullS4XvNSqG+oqHizs3NTr8wCJR/t1+2thhwml21XHqymkhmLUfnmU
9DjUNNsRYZ1JhGOt/UIksrgn4IVFimvu5cS7sCU4srIyoVPvdKYTsqk/ig7wE+QS+yMXRj2tRhCg
cSg993Gv0rrIKYl7NzuNgQ2rWY8yCHXZiq9Dr4LClMxVLVcGBxlOhs3H7u5W9edRJPu6PKOfCJkd
e5qJOZO+9dthOP0W9XNg3pFkFbmwvv67FgdXDN23bOaDPJnknO+EABJInn9onoef7amtz+aZtvPj
bxjBNu5m2eDNroWxet2fkjX2aC28iDTGUG1GxliSQCmV0YGKpSsUIU26PpuahopXWjyYY8stk95M
pP88Z4nAWRa/UB+t3DxNqX670n9Uf2Oy13shbauOD3baUingj6h+KJQSmjGqxTk+944h54AEa2Ia
bf1J5Qlaa2xk0nRxGcaJ/YhShzjQd6RG2RoRqYzSYunEmuakbsISwWZdUTOIIPoe1cqR/n0pjPJm
vexyjGwQ/Nb7EIvbO6jl9lyTk2c9/0onS634+o56Pz0JTkQ6M25pXjUwKyTQyt3tbO0TRVjtTU3H
gAcBOWLu4+AtSufd1ZM4XG6Xw/PYPtQfQrKs08NJWaNlHpWEO2//nmzZaEVrwjoZMPhZCC+n0AEf
oKPJKv1vJJNU1kfDDVWjUyO7tmmTM/AFCA8hDefuIeV6gmN0R3Ptf9T9saGIXD7oDv+IwrVrq4qO
U1Tg7x3RkkJp2bhD2dS7owfWoHewJKszOOgLX/kfvpmR68aetLYGQmf+OH38irk08S3voep0Njya
EENTEgGlkPcJriT6tSaxPB0kRMZMEmX/ruetsRSR6DluYnAOqvNOUZ5J1RGMdNzSQuhONSZf9C0g
mXJ5beqAKJsFqdBcDRgLyePHKOesMTJsanY8mTN1ywppqtNCB9+OnB3tUlcmvueEiZcuuOEMSbCM
hVGIdAkkDW2AYZZnhH0U1MbuWnZCUZNvT3b+22HvRv9liftfBjX03JK73Pgl1LufXY9ZmzqXp+3A
IfFYj41EOy13lAfGWLjcokowocX44FCRQ1dgM9IaIcwEWn4Cw3Pv/+H1NfuNQoY0DyBAzE3TSjqU
Jri39oAx2pjTajpqjBDDLLn9alLTL7cVsYxZRU2gSA42UOmYMZek7K7bVmxDZTDDP5D8oWKAA3zh
15s1ghlVawfGazA6yPy+i47Jub1wCW+bvnCYmWzSObCNXKtTAnFYeVc1vhmK5EFOrX/xLt//t3uj
POaX3BnKp5P8dBPtxaH/T+KluHTuCbQVVvyXLu925Oqr953gj9faW1RkrE8c/8CLlj6Fgck/2xa+
vv9THU6LK1/Wj7l7BhQ1Pdg6aQw6rqWOwnfnnT7cqfPQUDm/MmjoLVzIkNRjNChnbvMVGIn8BTQF
in9YEgnZdwc11SabbMns9gt77ZvZt+EC3Npb+Gy3sm10GpBRjHDTHpDJcnBJlmTWVROp49OSDyQN
fFbvblAzGssyjqklU5mm9xje7L4ZGpn6hSruEwm9ZFtP4qQY1vU6CQk6xNsk5+EY6tAOSeRglxrq
zJvM+LmgDSpOoulf0DcU3cao44+QnLS/kX6LyMwR8q76AS+dTAEAakDwPgHDvBSNNi5xfYZOvPjt
lPZN9RjT3oLoLwD50ae2Y0sxEXyUO/LISl1T8s0ENsEpJNK7Tut7PGu7AaQ9lPpy97AVFMgj/Dsg
H54scGY+C8LA5wr0SIVfe0ErJN3pygZCJjoWNHdlrWnoxHJ2vO3ejKx/XY7SSIatqxVLJns2ZKM+
iB/oHhY1SWjuZMYSTKixCp349CXYw2UMrrNTAEunjZH/1e8XmGk7itmZ9y/yNpzaNM5W59TvzJEb
qQn0GeWO4xbZYUJcwxzhBRaFIB8y814UftRAeSm4RG+fGtn1WTXtKW6zUvJCjMiROksF1Os0ZOUJ
BaxsMDsJygoN69HTk9JJxur400RGQtrfUbmdQl7N203RsD2cT6z9rRYZzIUwhDWOO0YvRtHmd1+K
AQSssUvRbW9uCf/ezvX5Q1JrmnBs/VSWi3Uioof/NRQGm8CWSB4FuE/schOKOeN3jdomin31Ddv+
oQq3gCBfl0JHuISYnycyKkyAmH+C5cjoy8Vq8WgB85WdoSZjDO+7MsK75meyYkfXXCgYJTqh+x9d
86aClHrOL3bCac//wy1KbOt6/mEWM4BPZ6c8QrZFbydPLJ18NPF3WplkvOV3oYP36HlMZkRIb2C6
tOdW7GMUQ/iUrY0R1kfOJUv0/90UqA8/LQYWWfaeLXFTJA64YpZA8iUKMI1Kx9FMyThqWuZ7kK4H
pFUQPWGTTSZm2IfzTuH+ABGGZnPPtZ9yWNPnCEeF07dwTSu9+1aCvN7unCcDfFGUUAG+KOhWRoR/
WUfhp0iFh2l0JezQCmb5u4bsnBJd5a2cY2XNiD8tMZTuzvYFNIwG60AioFGrs9N1vsuPR0GpoEy8
57kTXO+s0jxczf3x6NVnqXSECyGNITkVIj3sKjt08AVIb59t74NyQJ9AMUqKw5DnkOU0kxQMZ05+
US27oV4FI7Xd0EyDKNrq7cXPv9UDAmFy6qZUCRMvYGI0b8DzU1NNYn0G7/A6plVFwoNp1pbQjlMW
1TOaLD94Ik+j8/N6ZAxpQzhWanMfWkKOWgWW4TjPsGznxHdtsHp1NGOcyog43DZNG/rWZCMv4prd
Gp+mxGt8sAeNP6IDzkqIjedgqLvkOp99AFqly7se74Qe/dZs4fi/ICnaYKu7kje6V2ZNEnozWCzr
6rwDvRQ9VdqUqIbEylADqQyuy087JGMzcYfVTkpJRYW5hcOV+I3xvV/KQcKPOOwJltfLNnrIMyg2
5VB3g7ElQywkN5FKzDp780YS4naLV7BRGcR3CN1fr/lbOlxWPFhM3hlV0HDDQYnmsUUFbg69EKl3
AZ+Zn8iLwX/V9m5kB6qOK240QD8d6C3JLMq0BFVNildLKqcEs0lx9VJP457ot2hfBH/wkP9z3hTk
Qh8FxFkKPg/LTFPJOSxZeSOMA1VxnpmAnKrlKH3DxOvGSQG1jalCGI8W0XVvn1tRP4dg+eULE2Db
T70jPgrouLpQ9IxBacNJRjt2qTyjoALb8Hi59UqaRK9pDk7S6SGkLKgWPWhFzscnvkKPNmQRxZ7c
5NxiVpeU3Uy9sYElNeHEp7UWbR6k1KsUwM1Cn6PClywcKer0tZHhOoKhU2XT+EBZPXtzQxk26qTD
Rd22fuz1LhlOktunskvUSs+uyMuaREYtplUWz2rcjINNY1Oks2dWcHzMl5jXFdqCJRnw9EmjtYKL
gNcWUfDYOIafErwaBcyfH2x24ca/9wV7vTS9eGuMaQ6ONgZ1qaa2iOi/F9MUoAAaLu4d6uckoWLx
sPQPR6zOKCkyc5KD/JYmOM93n+AEy+/coyj4wYrd2s5IV+WgxaSOFKOwrKGNE8VPomH/OXpw7eJF
SefJZMCyfSXs+t0r9QaDbXEbpnieEU4W+uZRqdAoPSSW8KYI6OH3/J14NJ38cnTRFo3UklZXykj9
eJsmhD+IxxGJACvGumHhuWcK1k2/MmuYcK7j+YaBs7G2vIc5WePeeXAThJUNMz+BNzFR1mkAhMtO
LijJUSXQQnSqqNlMy1jTq3DmgNRC6swQTOoa3ZqqGtSyEqDfMKU5l1sor13o35itqzpQSlle8sK1
BCjMaPq7/SHr0fbDy1lqIm86I71wp5ZSqnb9dFxuQ2BXPVidJkAoR7PNdfCnu0AhE8eoB9vTGzTO
GzV0oe+WZDt5LOx+rVSfLIYJ0ofAkQ95q0gBh0OcA6U5UqAcqqFawk/4nOtwlDkNnCkkD/Z7isgj
WYhLgiuGcGrRoTRKFUmhxrSPD/M1mJi5Knur+kDx9YCsSoPNPWJfNOeDwplTB8GCAj04xukvyKJ+
+t+Yt1422ZBmPwznmmVuU4enYfzDVovRPStAuBRpk/waWy2nir4W8CBJZVqCaoQUycH1xGr1NE0X
BtqxafDgS0/89m/hTx/rFpgCyQ121cgH8MHDgp6ReCDezTzgMOVaGexQ1yAmBDmRmkJFpDGyzVn2
yUhhDi5fcn2CsGjEMIPA9XUHr+J98v9LHNeKmlfRyQlPOEhBRLYjFqMf3h7q13AXHuHFjhEu+zg8
CmWOD2/PMQy7NTEdfQXv1Qlo50wXGMPA52Z0wSpT9ctjMK1LiMSF4mb2QCG+mNFgqjsA7laZgnSO
KC46xUsYiv7/jnqrB7STc0So1bgqujKdoQrPRSTC0KWpV9yF9qxnU1zmBRfG5Bq9RDMxjUCUMOuI
tT6KS18D5N5IMjh3KWZmtJVRa7mpHnZEJXXKxUQpLe4elo0ldgXoJ8zHpB/2MDTqWNqdWuIYNrWM
0HFZmrTSYfq3d7wvoaBPqfG19RXK95tIWBjuPlphd0lXol3/SoVlScA8Ud5Nh3iDrWHMsekRsWkh
jxnEE+W3INp4th6uXOvOEJUFpumuz+VoiunQ80+XRVrJ9d1/fg9o7eQj/rR4cVHErk2FygxKu5kO
wmW9DGVGRvHWWD00luDnKX4oL8lYvsgSjboSsbG0gqivje8c+T16DsZcy882xj1m9rFBS/XBA0o9
2EgXbHvRibZ8CiqgiWquBYa4aON5qRPohyGp3LISQnnQOPK/nM8A2iGKoOuV52RRLa3ymrVZvK69
Ue29mx1BOPVNF6rhfGXw5eOR2n2b4owf+zh4VirTlk4S9G+q6DYWz0nq0ezA8C6xf/QjA8b4FPgz
Adw0GaZ2owjUoIvCHh12Mcw94oqVoNZNfFgKAvIXgedWCndH8qWYjqjn6D3qfHWEYlTPIDfeV9Dd
OQp0nF5lEX+4RMNjUaAeKZCrQxh2K2LhZSRAwUF/NFoGkcLnWlJFpzQliEPhoFgDksWeck3CE+0c
Z/vVZzk101j3j0rp8/9tSr+2rKxX69iqLT6pXhzmfIHv1ER5lX/RviWzWCvE6X0p2qu5QFYOet84
31nmBJCljWeI8cq7GKcAYTsbKpZR+WasIodJNJk5IMlAWvEsDj0DuoGF3LqeK96HOpXEH8bjrzxz
DmcZH7TWNvMo3nD1OjHO36CdoWjuKX2G3jIX+LOgE2hYDn7/dselAPlDBAzE015srtdPsx4M9ACI
5/HLPztDbQmccbRQ3771hfxxVqjdtOaiQRXlCxXG1KTjJ2Q/6TK00npmRVFM7TYl9RbgwNCQhw+f
eNGRmpRrkAfcFVAgU8SlHKNfCbjMRWZqYHbePeimhqPKvuYaogbj72Ty8UeSRBI0Y9NO+6Q3Cz/b
ltQfNeWWNYqH//5IsQ1jSWc12cdlkK7SocXsRjuETomyE9Oc3Y78dzLfShR2KHz8WPO9m6roVcBJ
mjFx+Hvva082t4LwNZstlEjmbR28yOREd7vM9+X35keqbNs5aYKKgHLJYPDnKftIi0OvBQ7/4hds
nkyJdTWmiNbEnpKRV8soc0gAt7Uyz4Do4qn7Ln6eEJ5XfnanAY18ku6b3iOUQzsp9oC2+lfxd1lE
YXPhZRMGMtgHYb6HKBuyrUFr83jTyWLeansm4kmr6o36BEwCIdXcTvveKCM+BAlO/DdywdNmo4y8
rGYA/jDeavYvbDIXpENlAcejj8pua6D4w8oaXDqvDNJzfUVZi61wPKEksnrcMq0FSS9pf5y0naeE
hJ20yBqtSDhNfF9WwVXO0Q85pFBkHbHBffgMY8BZodpU5quS+/uyY5E8j3RRTIqZtgeRJ2B6TtoZ
HUKycyuM3uuCfg5hAwdHkfW0YYJ68tQIvu7iQzm7k8gAPPQ41MQC7scxfOsW2S9c8ATFLs5nswpz
X7994yjubplzQynBE0wj9+qDLCnCbPPK5vW27aIC+YyEIoc0EMe0ZR2xnRDWNAdRTbZhzube1oAD
Pa4M5UtDwXCkK4qz9LwM1k43v5NJROdn10o3OzPdW8n9VgIimxzEK/7wDTFuJ3onDD/6R7PaaI8f
kS5BQSje1QsAk1gpe11qBbOuw3FcUn7FbgbttAcYyPzmaVTNXs/KeANvy9owqGmCgjvT6K1gTBtu
giAOnVYrEbi2LMlavtOE3uE2b7yhpanW8c+lAplhoFPtYlB3rAGRPGtEfjLebVQeU+gz1VXuGIfl
1z0q81ZiAxO+unHsDMEKnN0yHiqfsFQ9METVeQwPI57sos6Ex+ncIeLSvrkDGjNwlr9Cun+Kf2j+
yR6yLOFFcGaWP/9h3knavmM84/JDh9UH8PwpQ4TiDLuAluY3OYc58fR/nuI4774pJHVjEHK3sAf1
PQ+MN1xuFqKdzDibKhhmbfxP1ITgxaz0nM1+7z0x18AsinFNE4P1iTH8x+GsMDBYTBGT/feqSv3b
Gbcz7KgN1sLxe0VtShRpbPOLEaFc7qrL5JD6UpdGScrJo/cYKsCbof3eKxnewkEj9zQwzYozusxB
7/6Kh0YZvDGxPM/wORkRdOPqrEZBa35/GKKb0uroHcBe1Se4Sr8+o/0T0MqUCPKf0JomOF26N8+F
BF8YOHOVv4G1/gZ/uyz57UMyvAssteNbzWAwBx0126elRzRKx8ifv8yEH1BVh/lGjQz5Sv7CxhRa
tXsUyEqbiq0p0LOkwhSS8taBPglN1Ibd4VmXMorsuIddrdbGZrH0OIfOk6gwsohq5D0dZfP+O+q5
bvdvJCwHs4MkHoKTcUZh3YiwnScUzZy1iOHQK/UqOCFkfmWLs+3dYUlWytdmYi10QNb5/XjFtu/S
6sD3P3+gsQ4HwogL+qZZUYf5e7/99/W4NiswlTEvD+XcjPCFIXPwD4RGNe/ix1qrnq0JG1yBA+9N
U4j0dlMJmVahvKvdVR9ibr2Dk9jMzS6wZNdwc6rn4D8yQrPtfZ4KbzY+9nTOQ4NMkRk/RIBcA4Jt
XsX7QP6kImH0kQiLrxiRpTAxABGwU7m8f+5FJbISh2XwjmvVylVh3PAlfkYZaOH96PsGadS9yNnY
IgniTL9wHLPT4kaKwuBMWei+FcX68kbslHlKJIHZWQYgZJT1eqPRrCe8DSeVTFaYEPCdUBkY3CGd
AoBhoJ+ZcojXSopi5j2Fx/F+bJZ7eGZA5AMLWqdCclhCicmq63vZBqEYAclCbbwJEyYMlqd/LzQc
q1vUyI5E8zubalPE3770SA6ahVq49v8jlTlzkjOYCxE+ziD5UVxQCO3seq6p/8LgUL1YCk6M7mvJ
idvjI03vmYOD+1/NWV8/dnvicspp0hq0TMsKvyRmtfillpKE5XhdR1Y9ve5Ei9G4d9TrnHsT1Erw
8F9ayD+7tZArIdHcYmHpbzV3p87DgfmnZxKKhWGjmodBp15VdQX9l2vaM7Y7mKzrZW5TVsr0IQZk
GzH7tlOyYrkQZVMJMFwiDOxuqTjY5Lox61hWXkgSxD2TkbLoHRhJQhoMyeORgw8OqOd99kb3th3q
3xWmoiRapGdqvbBtgfn73G83r+cViM4qzYvDoc7m74JLSKJh+iD8ucnUiMGd4zoeuNDDxPmts5uE
jZhOzmAl7ec8pPWB8B95rWeWvF1To5izRKQi6IK/nE5o7uEpp8KpVxjF4qYljrnBcH9byCuZSvvW
BQoF/QuEmpMAol7l/mzEVxiu+u3tVoOY1/q9/BKVZWsnx1oGmw0rzAm/B2FJwOA9saXyN5KxsqRo
GSfprCi102KEJ0duUKb5xk5U0ueDYs6xxqtMzsUABnPrfcjCpBUGKXtmXXSI5wWn3VBci32DDshD
ZR8hcoYGb3jWlUgOsiuj1cY7+68OWKWcUkCIvSK9ATbpWMUGkln5+uMRAm2XFrhHYFMmdm0bDyPL
xuPg3jz7mn4FMgEMLRlf8aqkr0X43SstNnlElTa+9kKQ1bvD6IyY2aQXLLJ+4qEfxZhVpWf9lavz
QZSBoL8rWQqDf6gy81OPjzkYP1a62R/7SEbvm3YX+bCaPJmJP2cnmg5tQkA5E+QrB0drq0GBxc/E
tc2SjFVClj1wK4VkMqByUf6cdrDnCua5duXs6UR4BuW9q4hm1APiQGm08MarS4qKCsDBhw0O09Rs
GjAjwFWA8wHlTuQpO40itJDjBgq11KoGs8vZG26ktFwgwLmPpYoptFHkVbzz1Qn2dsOtyNu97A1u
bfi5HkQPqGTariqHKpQNnFT6BVOxryM77kKL59+fJ8WwzkX7roA1VoMsn1irit8XQx9XmUPRZJl6
KPukvAEyrFobc7TcmNHGWBij+sRAV/monzFbjucF7ksxNIyLkbEw7K7hnuOYMRU2DQ82K4967EgC
LyCGt9ij3vPYO3t+Y3CeInhKH7R23MUCqy5EV1kO1Y+J8Lppnix/8CtdPMu2FGVUtuMgsHUV0Hk1
uR4hPuJvyn1fXmGksrgv3RfZ01TDUAJgNQaek8fX+johgW/+12UQOdB08JgH9tN34qvkzLcRnoEt
MNpCpXAnybfM1oF1MMVqcW1/7YItGY4pRQJH06BW//PNZA50TornmAnD47FkUOVFUzBUwPN6FnbJ
Y5jkaYrk1AbazGRepyaxAe2SZPwJO4XJxbKwIX8Ds91u0bK4v1THdRDLVARkFMEBxRQ5+qZLSXM/
5OLKGQLc8v3e2UmrH2bG5F8GC7OST1odldPuCvUuT0NPY7Fh7DnAVd21+LqxZBs/FSE1EYmEA1pw
J8P5L5ynSdDzTWOcuX+QzyUdS+iHR3+36SowI0H4H3xpTKqFjv0uv9OZzIQhffQ3bF/dsA6BnCyC
MeD4twaF/iYbINdtDMjn7dXCohySuuEphdby+YCoR49bXSgr7eH1/hEQf0rmnKH3+Nsy1hsVudCR
tkMmx+CavMFNyKkWwxQjN1OCdOdlAb1BtHQEzB8yE0UTnwdrKYxrNnRcr+NglcoAoD831UBuC7oE
MvfL2LcvhtLOyHwIrp3V69SynwoQPP2sQ0jWjMfxQ7MQTCpW1hdlT0C7XyctaKFGBlf0zd7yFg0c
eqf6+M+XMc1nmaB/HLsTRU8Xx7kYrKK9R2hXn+SxuuYDX4lfz1eI3LfqF+dQ2Vgge13NQCO+m4Hw
N9YoA3e99WpEZcQRGQF7mI5wIuN2MXZJuqzrE4ABXwLoHvVt9VtiVYj4xbKsBblQ/kL2j7Di3dug
85vUufojAjUbXvGvC1MGd+8bWz8aUvXvvjOCfdDdOE4ci+2xHcJn7QsxA7wQ32gaWAxd7LfyaeHN
DN+rCCGXOKs0zsoi0jlINZgOA8Qhlz+UoUmmvRLCLfG0MjxvrgN3Z0fR+pQM3UzIc0mQV6UCn+DI
kSDCFJWyW7IaWc0B/KmiVwhct3OhpCpUND/lIb2Twz49oDMSvcYG25Rojj/2yy2x9QALNgpmDGIU
YXi61cHcOdA9exvMj4IspZZIP73hISVzhnWHJgPpXF/5kiq3EsLoeLtXHdodPxupDRmTm6nv+p6d
Yy6WYrwxkNFLhZ/egV2C+p/KCKWRpLoqJR0Zb09/kq35hkzMPOH6QHinKKGWgQsc/Hgaifd05DWw
UJ2We3LLi3BuPoR48lNNQpYCbkIaUNPWck2jfRSsPY4YkcQyrizQLs0kFuMEgeYCc1n16j5Xu0g9
IC8xNwe31kAJnNH9iLVyjNq4/2xSJMcCFc+SNf8IzuHSBKdo1EkYAVOCLkrkqtam7j4WIF042akM
SCFQ4DxuVDbsxrWTHrd6y6+ER+wxaJeKs7Qqgpx+/JlybJBrn2ha5A98Rs7ccMnlCCyRVHuwyjVS
EqY+r/nyM2xGWRwaZmqheWUPaA7M2DrRTi2iYK23srEq0Zp8hnsWZgwubHwfUPh0ZxBIBPjYWtNr
vC568zdFKyEvl9lN52s7leZYvYIxZ1YZKJYY53tx367MiP/9W3ja7LaMcDGt82FvZIyLtFwAii8s
puLkkBLV6N/n4KlE+HnOVS0HQsDGs6FQeLHepK51KW5qYB1MTBVCqbQi/S35EGNcDP+v5BQL3hjo
C2TJa5sQ7DR6h2txtPiS0RbSJv1EqT+5jhTsbxY0LjZxHXtLzVfepKDVjQLW60wayKRV3/BxpJlG
8/j/FxDi2YdyrbG/oMr7vfO7cx7LSv+3TkwdZ3Qtzic54hhh9Q+FScNr7UYccS5B9ibaKNBAaIdq
U6TDVUVJKo292x2Ewb4L3khYdfZIWNsnaNfGBBF7n2yxPWFuPxzGxCyEiPKZ5//e3nyjPhV6Qxic
GbvZ724MxMsFoKkNaobqK0+1DfKl7Z4GdARlDhYZnn3hGhmYW1u4FmGsgkVrebC4GtViOnmPWxNF
ojgebNPjIpr0in4hU/DgUWqmaJuDRSCRbH/FCzI/kaUYeLIp26lq4muPaPEavK5pOIrxhONcIWN/
qwl/aTYSkX3VzCIZDjwHxsFVjWFaeK1D+4519Bh+QwqlZFaEsvRJZoYy8c0+I1NSLkv3PwHvkung
fv/reVpPNa6DPifBoiwm3hmWR+cUCgsXTa2KkUMqlmnpiC/Eg1Dorf5oJWuJLOOTAozmLiCumJWh
nJOX5bUw/kiNDL3I0LjLj885J9U3Cyjchx+plZSpHyM5hYOEXyHULI1qfnc3qHNNBlbDkjUHr4Ih
8X4BA14/PFWU17sGXGA6fU69tEakZxV1DyS1wjcztwvoiLsZlzgdzUxSNa7j7NU0EfVY+jcMRIb2
RktCHwDIOibpWojlncrdzmQTiKzAU35m9aHezzYvCTRX8/WbsgmJ/G6gchfKJUE3kTtbyZJnrERl
mWXhhEXKu75H7LcZSKChKMRWxZTG0MWMwBgh3zk2W7ChqeD92RPVqg/2PRhDfncLyEk9MOfLN71s
hR4pCyJfW638xKZ5yEX4TSwkrX7jF4hx5cjz2I6iDbzKEcX4kZox1Vaha94w6oANBwZT21tEzPCe
S6vEj1ivryYW6izRfFV4qeRv/AZK2HMqcKGa+boBC1O1aQMM1/SMvVagS7iMcgH40Vz13nD/T3gg
JLw5D4Cwd1ap/1eCBeQ0qqpa0rC88Yf2WbjhhVy87AY+DRR3mkdEvXA1gIkJXM6LK42m6tAe1Chh
BgFIt4HqKkb0ofOLfgieli1gpwzqlope1SHFuxtMaNUriSr+tCGh2YfCL8293fXMFskbiRxdDERp
Sm4TB54PiKXM4YgyX/bJfHVs3boLGzwJm8XwHtWlIX14ItY/GY9rgWCttFGMt4D67Tr8IxfYK9sM
e76bfw1pA3itvAGPgw50pNiXFyTBJ/ojaYhTXlV2QmNbFeLWEALnyshKk8cfKiXcrMfzioFgCyKk
rE8XoKOfMymmH96cqiI7w2ZhzdFyqzhtoymo53ZH4b8ZTiF2rWI+yWy+R5aZKJo6iCtwWtPX5WdH
kmY7li94O7nhNObU3p3VrKvoySUx4Rwa/f+/023+m42crOXz8dcBe/uQCw2bZVr9sZHjWETMsm7Y
4l8rsT0eN1IiDUCSuaoIAqeKZMySzN4HGYLzb2AXardlLfp+EzvWKE2UvRgrsdWkeCDOMHhbypKq
qykEQIMD35etxp2Qe8Etzi1RHR/WMulNuqXbBZBjaOYK+dQsH9ClusrD7rD9TIpXCnF7znzT0jpC
UdiTqI/5AZSHS80fcy8XfN1MueK5SEXbIgOhK0XqfxTukkgSBsQQZpuQ5hOJAHt4+nfADEZI6Z5U
yrfXH6vBnCqiOhCjYD8aPhK19NXNxkxycYr4ya64efE2+Trl8okKfjRZs100eLzFq9141c5/7V4U
bHRzrmM874gLratqZ8bwAE/+uPTbV+4N3mnoh3/Rz3coden/lnoLTmAdmq3hlp31FIyCbV9Q1fJa
aRzg5pn020HMl6GCn/P5hqcq8SHzOlfnHzIilEVd1TCIxb0qgAQm5bCVdfi23RAlNindadv3iba5
rrNiMZmVq2jI5mZxGg/d3jy+OprO6jv+rReb7zTtonj2FcD5o5ip83KXjj9Fl1oHCvanwtIShGZ6
BU9bXiV3Fkzz0KWQxT2MEJUNG5CITzVzv4R4GH3NvHY3bJZT7/txNyqm3nVn9NXgK2+hbb8i8Ai/
ZoQ1Iy0RIe5Sw7CF+X6XjYd14S+vDR2wz/NK0Xn6qKUqo7W+5qagDre8SYqdSw/N3lLSGk6mew5t
G3Bb3v9n4dUfQUxpfF7SfX4uCe1+VkP+sNL6L34ssjwKUT47pEexQ2RfuGcoTlK6fCopvzsWF19x
m6g4wQyTsvECRdwz4nxjVk+Nn6OevIjwbgY64jJ4bFoahTtPgLpdvJR5wq25KjDTnzd+o/7ktz49
nN/gVp3hyhIhIrrX5R+pnJx0UtTPEXbLx2Kq0WNnu5SJBHwUwZ4M4oQFOIy82cv3009AohjkwqBC
rvZ1pjKb4Pctp5XvT63PCYq4iqW68wSYDI9+OF9xdkrL4YvxSHIi9rA0usw5OVGGx9Nr6IjkTDy/
XqHwtUPLyobarsE7+b8cEVMWni/vjAGgJY4duXAHy8l1mi6ydgxwmLD+syr4IsjewzTKu/T0fi7C
aC1UK3iFFGZp2I90eEi6PiQD2vu0Kt6PBkOx1Opy94bLOhWAUy/2xKAm+vBl+jlknRg8ifqwkXH6
a4v40/9eFfm3b6Fj+sWoyqxZAtBggzU7W+EsuEQFz01F5ABpt6o/uBN9W/bTZ/PkX8Xta19hGYR2
Bi9Y5sR/9ZAuZzDn4mPyJL7+teyQw2xidADJ2i/A61RQGpeLLOiqdDwmZ/2z1fyqSwYK4arNlR10
KpXDzn5/L5aBmMsmyuvTIHsBNjTa0uLELBi2oJyHGGLIy5w+bjHUVWpYuqck6p4y//2QWSPyO1uT
7P3shaQfYULxJ6TVffFJjlf++swDe3XdbZ3zeupCaQN4VwmHCxo8CrUzFP9AATC8oRagRV9HdyDr
49Vne97wNElq34NzF/A/3SHniXc9Eg3lEVJ2lU2C0pJwE/+RAENfSMFd7xufKeM/W8xIFliFo0v+
Uaf5KfskP42fVaXOw8U4LoXuuLVglVF9KqDP0Ka8KQAlvMfDSGLvpVJJHXod8ivmiDXwMSvJ2Ktc
+Cn8E+rzSsEUAWFMc+oO9gAPr69SrpwBGLqLNMgxEjxlVGlFiOVsj663fGfEjjNsBDkQQBtJqb8b
Ug0Q2TFFY8zS1zHlNJTcLKjcaD9/9LfObLwjwQa5Jfo0gBfvg12VvnsSYM+2VobmoT1DKSL4ZNcV
TCb7QYKjcHxWUNs4BNwydTEWv0JxUtq2pnJ+fCyk9jL2oCXBV/r0w7dEFusXOQPRdSFcRd5AcN3/
vHlhF8YTqMX4YqnLML8bol0Ky8iBKXhcZWkT/2JJ5h2UtJ3hWvIBn9qSrc+fO9Kd04P/l2EWjjuF
jhCbuOIVAEoUF/ZqwxSIYaTbEIgZSZpjee8La7vRyzmXuX4T3CJRTvxAysfgEhRJXxj+lZpHndyw
oePs4N5yOcyPm7J0Lgw4sU8tLj+lYWv9OktNu7g9JUEOc3sgcfBe6F63o166XLWuVhh6nZiNBw0p
Qc8Nar8JnCj4KvkVH5TVrv+c297NNduXFSB/q+o0QN1HYprcHlC0U1+xfdSco+irhWewPkxcI9VY
nPKIqR+JZlpQN2wb4WqslBh8fxvV0ETti7snGZsuofXotv5kBrHBXNvUM5qZyrrQ8qU29rd61Wbx
r5KXckUAN0pNO8J2IzZjTS/SQaHJ9hprxq/D4UZ2SoztOmuL7KP4mHrgxR7TQ3IbewKlUKoaRqHt
AOA5xZZT9XfO9jcZE2LvMRxwfu6Lzu1JRrwcRqY01SCl1+ShiBOPdQ8/D5AgM4wiQFS/4Vd56zVy
p1BisWzrJFAQd9hZyi9X/9jsLfAKVpmzxGf7DQ3Eyx+sXukpoQl1RW3F45MZIVSe4t4MM44Lxej2
pFQDYyV6DaBhfOI8DWXG9C7BXeIuKEAoQOC1VFuaQES0VnTQGuomd2nJoF6d9g3fDhwDGuuSIbBw
j3m/fAF1Dv7f6COqWqhgtxbYhhsOl4yKZ8RF0hYdnZhTQoGTUP0eIfLXtSYqwXRWbRQPgcwLh9sM
rCvxsDD11v/81gs4g6g6PaQUQulwFkKyka5A91pE8C8rsicyZclhCoPp7dTBatZaO0OPpVlYLvWZ
6fT266U58FCfiUvKxNlGfl8ICsH1zu3H4swIXuk2Mks9X9nOkoi9K0576RHhQSHh5makC7DxUO1P
v2MfOQdNSrPDPH+CFYNwNz2EfkRLoF0dRCjTejJQHrDmn+mlgrruBLbVDo5EL+rUgKb9cEMIED3P
m0CUwMuv2W7xLT59jv4Rb0mij6LYsRgHZc3brsrhjeHJejaXQXCzoQiICHg6TNe9HiypSgk1OzsG
Nrt9uqMYl1uxsS9LJx2JlwKjBBVtoXIVoaNEVM8xc/BxCeu7Fj0HkNeugU4SRFBiJSKAa8lhp8ph
ecgLYMlI5Y5ang+kd1qGzHFHhYzgTG/MmnPM1/pdMRMPRzGVPDVstJKM9lynPGti1xFhHmHylSge
RTGBIImEs5kTnUfjIvWahTwqURaf7fg4N1Jzx9NLqaIh9HpLFrtth5kBNWsiAz9kp6rwWLfRyDta
Bo7LTlR/pBlvVmBWkUCEJA3r3Fi0GMSAY5XhDNedzzdkmEfErL0l1h6kODtEHPmn/voTNajMbsUw
jh85Jy7H8ML/dopML+gW+WM1RVd8fD3fYmVqbZxZq6NdOoW/ullTh4B4lF/iezq5Fyj71Y8uIY7v
Umkq1MW5IKp/ple0S4liFo9BnHhKJch9BXys0isQOyd5Sdq70ki9HzVr70LrNSpa3yEe5tsas6Fw
xjLlpxK1OCMNLmAOPaO0Ae90KswZ0ZsCQMoDBJCiq8AvZpmFydZCb5iAHdQBArZeoNyMj/1KCvk3
AZFNo5k4XBfukb4lucjwlsBWvr1x6g1cdvqN5eSNv32julXW2iA3vvVrAkNcVduReiDgXuzIF7Ms
kqGcSaaAal+ZDDY4y4BJUuYsDbv1pe7Y43RmYenP8wsNFFRTIrl1LjPzkHWSjKu/08J+tfWeK9Aw
jWTqKtl9HXsQMatxtbEHrvKMkYURdgqe2moDuepW3iV35JGdoEZ9qkvprv9ECqk7A+cpjKBV7zUR
MOsflrsZCxAsX41MJynw38kfVMVqZZktgQCN760tBmabH8IcQieipyZ7f5Nwc3EYEr6E85f6Zrx2
Nekydjfi4c4rig6Qr/jckch77s4SCPCi/k4SzEqc8yDzCQt24FTD6oOcNC2Hf2Q8BGzUiH1D0adv
QaIQgvmmUW1gFH0/7zIkxNu2ZBMvkeMgzpG8nziExXhj3/fvTfMSSr1hcO4ekZIgj5n1F/z3mD9+
UdijO6nMEEwm28cYh+56cIC3FL6I8ayn/z6rq8RzSGtnusKhd5KmOE2GCM9GDCNtb5yL8gBhwd8n
nVhHN4g2kEpXBDnci0NnmsAtYWbjHuEe/fVR9sinVqAhH5NRNORUfu5l338a82kCUf1Jp/2wrXlV
y+/nO9Ahv0v9JFq6rKR9T/w0Ks7WrRdR3ZxlxztnVzPMrjauKKVND15OFld0frZ6+dOWWReqYhxX
SibzxIpt6af5MAOVkUA70GOYOkt9flNi7y0stY0MtNJclvrta21JWQx1WnVxpT4qJgmWcyBYafAb
AWMpJEBfPyi5oPAUNC9iZgjF8wVNYVifexC7M7ylZnl0vhP5v2+Vc9B5vUVRxLVOpvAx8h808LHV
7TocFWy/bkrqg8C37kITtM+/rxS5x1uhq3TSqPK3X+pKnVeMWC6M52njjgFpR2xgQr+Onkkmn3dI
HoEc1a+fiEE+kwbCr+M0a3JYBa5wj0uLF+zdCiaqZSUqjISIeb6Fn6f/3u1JqNSWm4v+UCcPLbRa
6/JQVZAFZh/nwVwP5C3ocDaB8RV94pFAy5okSrDQngxERwIOypxonkNmPS1lpTZELd04zvze0WLO
N8oeYFt2PFM7lo2TFKJSvNWSCWKiodS7Cut6UGsreijv5AAVkvsqcdygfnZOcCa+NQwkmfGG1qT6
F7q/L5dHRQJorZNMfXAKhLV3DEaYLQ/EpYjrorW5vwpGBRrB6dCatWpLrqKAIaQGxdWg5JX0NkG2
7mdxxKOXFrsDl21QExY0y2DqSGOzl1O6Qqe6L6O+zJxK34y2CxpgRg1PmA4tjB7X3Dw/QVlbyfRY
U3iI45sujW5T89bYNlTYM7a4IeBLK+AOIq2Cfb78bM6od7uIHYSvlbeZz5P333U5+WomdednBxZp
AwvdW9df0VoNDsD5/RJoYpz3xpkVOjrZyBC/pH+1amlWQnLkN94TXVOt0kIH76999ZG8k7Q8fMSU
v2nQzL21POC+DDljgGTXlQYHUBxW+/kY8/1QbL8QH232imtHfvmKV5W2v6Hymu0I4ZqMHJh0rRdm
IfP6LEseb+qJZTWwsLh5zFODqTGx8tvpvP3727FBV97Ybj21eLph/kYZRnjm+4zCQXpRYWSszSnK
54AOAsaIvLFa3PAcVxyTN4SINyVVjA+OeUss5jWIv3pzWLpvYo/C7lBQ/MYy1woaR2O3upcZXV/M
5dbOZGJdoHgGL6B91pUBF6ltnny1hEu2JDVQNiOkeC7F2m8QpALBofZMLbxNMbf/MozP8euOAuyq
oTBobzDSOie0ByfN5D71LyvQNVwDe/kBHNbSjVDBSFc427wtvjCYIXoItojKECIChTDjpU39APXB
lHioTzDa/4OUokKpeH3nNLxrS9xS/EgjJbwSlqrHSgCg+fBczfX/zCqaH4euQWo27MJm7SeENmLh
4/VHuPOAs9HzrRjvp1iKNrjNOU8+m6c8Ad3uWMvPLmnzWZKgm181vooRG1xBQtHCoNeLHRByvB3L
vO44dSiYOlMGKB8zW2p9Eptq20jzqWIPrMFV73WUYNIjZGNnLdvN2QQk0aYH4GdHgZJOwOBNUi9w
yIDTbvHKmTAEyjJE5y2rVY12GmEkasT3UlAWaU1bjOyFX81ycYwTvZXKzfe2/ABhUGIqNdBP203E
RXOnPzc8t2hSxoVsj+SYlOmxlZ6ZQqTBqUfyqj9TG8OOHojDiDKI2cmrKeZN/fxTMpMwy12BV2zy
U88MbGaaC2zJMmVBDiRShogbWM9v+1qeW3eAqjwXxWnJEVzQiy4+bFjtT9SssTvdIGoTlROwJO0d
pwgOocqiOo/WR8CxPtPfQWtlnmZaLkv+fZqg+e94uC8AdojYHcZ/1Qt2eC47xo07ak/nGVWGU2zB
mlL1cOmfz6y36bMU8GDKoPYub/i/7ldrypyD1+dqZV1jbdp+cQxy47i8U1ylju5lBzDUUdHfVWxZ
Maqb7PVGjsABhbvhuccWcbSKVgcd+kpzbfVwmz5V8b86TAzkBUkJPje3kzDW/dfubpb0wY5pdJxh
ReLBi8iDb8UwNoB0cOaG55+ZkWIMzBGawt1kSFpahe1uCqfJsSHn05p0Xm1hoCpO7AdTJOnu7wV8
D2M4koXqICMv7M01FwIaXIPRqq9baXEtjugY4680a0vI6wLa+xvc/yhRY/S4cSzVBdAlNyc3Et71
5/d+ra//vvWkmRjvBpz/ONDXEwkncRD5cDuki5RXTLj06/jVMxfLacj8O04n5ufGVscjalpLN0gH
swhaRmfIPsMlsZw/DEu1MfBSoflNv+pMv2GuzvVjEgI/N3b72X0pWtL+f58Otp+KCLDmgTED03HY
aDncmSseYg5sxC100bxzRd9kPurpXIY+PBumCSyaZRuVo962zXDm1j1wt/lO6mRZf+kpl7CbcQpM
kl9C08tvH8FgNjU9K4/+4bbsuYlIyhv/7J60uqesX1fVPFt9mGikrkB3rBWglq04j3DN/4YJVC8e
CDWVI0Dek8Ice+2SqZMJPdzOptahBKE5R5k7XbHGGDH0rsqvEF+0FCgujNoKrJl0Su2Ji9vN4G2r
z8Xton6su2Sdx5RKhenEgcRTveo+s/3WVRCK6Jk8O3y1CIWtHzMKh/lTLaMEkpKc6VmYjcsbLsnl
TDYDSVGGB+L1aFVupoUALNxOTZPvhhBxl55M/56Bok6Y3VFwpS9ZCStxXXLQqX1uRLI46yzfpDVM
x44KJk4ikI0alJCyd+2BTAax77rBKLwoGPHfKQLDpS/WYh7brA7qzzX4IVUa5VrvCCTER5XC2/t5
4UYRAGnnGMwmzQElqELUPjdXKaOPB8cULrrLDWAtUnIOq9wG9nWwCD2Ve1aaAueE82x3YUtJbujZ
lhUnk+h1R+Jn7IwtupixN/hEyc8jBx4kH12C3zfqozoYOUrX4zGNEehtBK2CwFCIGOlpX/5ZAq6z
BvO6/GPJ70CKWz4FGaWj/biSsz7c/uhrqIsydH9SuLBiEngdoAC2K+ugsipxsh2EmFmYkp0WmKGl
ab8LIDIsoQ23ddg0L9n1iLOEjSPY2haG/ah24oPVJYDWDm5/Dx5yP7vYbNBkSbwdp3UjUMUhLUmL
jxvxdaEu4i1XgRdZcs/0TwILg55gcazdmoMSgcUKXZ1LW1yu9Zueg1CUltFriXNQmlyvFL46fcKa
KJlrvByQk5q8vsWqtTZmLMyxIRvfBQze7TzW4h1MymAlYRuP7h2HnyCx3F6aDsZiXQaw5G4mTZUy
30x8P8qAl6MGFXQVxrm3+eTULvv7wXSqcwnW4QgL6t9AHGh3EzNdSTgHiqxcqyOjUScprk/qY0fX
STXkGySCte6y4G5jEud91qGXWMkEBbszpUSpEn74CXfND+R5APX+qA/5bLYdqO67AeZ0TVHghMXK
MmiBdn2DNYf5/vC1GjqaP3vLt3i3f4n+md/lH8kMaT0Ve3dMyoHQfbgEO5+XFyKtck8H+KGUY+Ek
nNzSX3d01LQUUZx0rWEmHrLWeu1GAWxf6efDs6AHTdpAelhCDlCaAc//BI6+6KUxBpeWkzc6uQlM
fCy8S7oEjwSkuwZaQdc7t5mutKr+IYNlsmf3ecsSTaewKsyH6lpPyDoHzeWQ5diiMHXm6HLzQtZH
fcBDnLFli5tYwNj50gVS736uRB/kyBdzogD7yDsVaFkQk0I0OGkvBgAkHwM2JSlswgD7TeLbuer6
Ly20zroapxOhwZUSLfcSgzmWNiXEI2appKY/DBUaQeqPXlzlmC9+U5FYG2BRFSAHcma/1tLJzWtf
pAV60NHn2IJzgqAP0iElL8nj1HcXhLB7ygGUm0WRPo/1Jsk8Ockj+vfvzwZ8MQNojEPjGsBKYZIr
rQAUSRQz2X9obDbSgHoI2pPjLNFsPa2WSAPVsmoadVeZlavpglDOztZ0EETAT48G/a6GOik0yogv
2QoavZFxpwEPUOTNL2llWtxJOtu/Ejvc5UnWxEjWIVSHZnIjPo+1WnLcksGTuJqn5/7AJXSQrz/1
tHrzf8S76+vdm/YJyv1Or8E/hsvhLs9nVWjY5FZowhHw/wGmP2asEyTO3wW+zFThw0B8Xh13rnF7
w6wDS9Hyu5EfwQ68hAiZYZtGOwuY206/pwahPLnRbxBB72LDiJ035sq7t2Ln3BQ1Y5EGcgoGZeVr
Jmws85/Ml6zo6dvSGBmVtQkhwBRNRZnvHHhUPmxJMTSF/7o1i8t9zs5jdWWF1Z+OSSce25n7WLkv
8A5S3ZOBLJRD9PhBQOOfpmGjUkZlRBPRGPGWGbQ/7bNpvytheRWaXZAksFMEGAX6WSQlBSTFiwDJ
xAgWH1IdygDh6XMmXG8MxfUDVBtxtLrb0rVtBhpThrRlsuh07z38LMVrOJqMvZ/TYRqiKJfzeyVY
cDwo+PR9AqjhbCi0dJVN+6cwwDRld/FxLXXLs550Aesca0ljjuMpDICejsBDa/nvHv3pHXlNqtH1
Sr7haPH1zrVN/jwu3eGo/m/bNT9fZRWQzW45euAuwxAEs046F6/mB0dTz7Wh6UFQBVLk9htZ/Rn0
XIC3F4CP4V0dCm+W0GkyOgjmJRGf74zJp8sG5LJldAsPCWFnLxC5o0CHS7cWo0qWlD9o4DMO1LHh
0Uv2aQUvWfk8Wuo0dIYaGeAyddWgqiSGwS0UfhS6fJ8peUKiIMVtVOG2Gbb1AEeofUnJ2Dm9F7mQ
oc5oiqhAo6+HM+nwtXHTr9gIE9UftLK2+Fk/vg9ZKFPjEDkBWEFsYLplNOwlGDPObTi45N0B4mMv
+fo93bgMtuLsoR2oKB7bRxwVbeyNEL1jg9sb2WARb6eoPCOin9SHAwigISLrOOAYtMpMs7Hit+tK
+nWrdxeV552VlyVL0EUejT063eBX+NacBHxIdV2XdSQST6WQsAAQHIZEWp/jPxJ+Ouux2eMjSNYn
J1P7SHpz8vfRR8/TruPZxhk0YCW18k1qsdVnY/90QoXlCiuWxbyTk7Ob6pXw7toEns6gHk5XqGLR
qkYzlVXdxe2V9rBnC80SAIBD4w5w8/ZQ1yJEaPhlbCk9XDDSWqyhPMw05ouIxOkY1kn/Rb0vIv8j
88uMJ8pSX8bRdt3A7vJG4EJuIbIvAtdWbOZWURXPb7LQ2kSeF+eNb4tNPns8+emslIRjd2skoqeI
tG4BdzkU3qt0BRSEGM+8qM0maWGeB8ppGMKxIq1yFyY9wcRxrmIMOyvZ32RFakubIFIFAwm4tQmB
QJ2WwuuEUHLQagIi9/MN4xjD5yH8GgVMBgZNHhRPs+FNSQiLZt+u9w0qqvKw/U319DvmqvuX4IDg
yzlVbw85FeTtvN7kvOiQ0ha/PIE7FYXbR50M4eEBllZWdbPJP6hZK0gMjli9tbkrJ2q/tAhq6bSV
rA3gnAqEqO2bQ2U1vq22K2/nLGncdV+TIaEli48miFTtWyLI1wv56gZaZt3MijQAZC+GxZXPQIBR
iOvKpAh7kpaaLJwBhgrb+UMdU33F2010OeUstMmw8qCn0HTOVRr6bO27EDA+gumnZFJOch3SzZBU
b1YYSIJ/+ITCf5mR2qxApOKqh7glH1AdsBE1blSPXJFEdbYy+lOgXPVrDa3KL4M2iF8mN+P6nhFc
bQzA2AIOVWNzDquv/WsTNOGyW+KD/crdP0ZEVm3nyEqoyqkPDxO0y2yUePaQ51GdpH4boBKSic20
HZ+GYuxcUCp11T2wc1abTj84teiD0NT+JOQv0B5VtNtVVTR4oePord4UNIcPPEXxAQXrDz51ceEA
491uj7flZrbIR5+I2Wdpg7E/q/LSt7puVLbruQWiE4A39XmJjSt83bynkpo4b6N04hmkm79QpljA
NP+SNpnUxm/aLrlT7AQgZPRZFWBaYZkcc61Df3yIrDBsQb0sRWGJzPvj+y0tIT+iZYD8Xx9qw7pL
Wxq1MmxZPAAYSAULzBYS2zOR31WrwcRYvXvw9hoxBLKxuXEfJHxY5NmTrClB+ZrPB1QnbNoZNxzO
a/ySBvwcvV289sUtzrfmH5fSRQ+uQX2cj/2PtN5KlNjq3Cl8Bg+bl+vARDhAvH6BNwcMRakKLltu
/mY2WCL8btJYPyS+CYe5kvsXd9IGuN7cLID7hCApx/oGLewO2T1kt5a32DbU1T5R+E5vgjDLcr2J
ztHoojTOuTBf0Qi/b5LEsfwvj7+RvnrSoDyBdC/DFLCWI2QDuWRR+vonLAE+f+1QOtmRM/rlsr0d
aVRMu67xcW+qMwl7XccX0qG4SOMErDGFC72yG2J5/4Jg2DBQRPHPnlXl3haZRpclvgFMxr1gag8f
/SBLenCxz/u8fYAzWraGpC05Bkvjz6QWl3A4C1o8PZeT3Xmy4RwWC160MgWyRKBM76UKvpx3L31G
GRwYBngB0zbBYF6AkxKVNxoW20Lk4CXggr4vHu5AiuBRcG8rOy4VO2U7dAMsOFBktEH4eFMcjP1L
5GHxPz9lgfF1ZhMHUd2PwMKSHTLXZYa2z4/tSXYq7MB7gD5L6O2MpvW5cDnbbPz43cCaZPdq0Qiy
ZH4JMl+CNIvwjneISgAWHnhRvuA58Iq2S/wy3uDDJlB4JAY6pGtXaFHYXQJ1qx4zRRBvSesKwP2J
W/1P/izRgmN1DqPsqDFHSj7JzCOyHtef/j7cvfTQmwkOb1A0ZpPXijiIun2k7f/Et/+80moNLZvG
PaUyL6SnrF/ZDDshPGuoHLh6ry7A4p8KmevgXuM123CHPu7erJ6qs15lOiRcQoe6aGjcYOYq9u8F
eu2qvE2NFPjdEYRM14ZRosn4walCeYNjnNLW7k/nxUl3clq2sLdjt+tCpEJ9NQX0NL2wKY2a1FSS
7d38jCHU5RqWIQmyNDZ3KmBVxeFGn7N+luoM8RD8RfzYa/JS/niLayoh+Ts7ytNRidfLYJqMLRee
dZwvsxDkyVY1wBq7wXHkJL2sipLUCcttvv0m2qU1a8qKN7D3gscaKgizsmdKFE/K+TeXDWUeOP3m
3/Xjn9IODaq+TCEmN1j4UN/Y/8FJlXxOeD7dlH9Ll4yEhdj2xL9KupZoEoBb3pELEVodivR8nRyn
Q3bVgioprZuFYhXylhdIc5/oAKrrwmctG093tnA0rqBI4hYeX9m/8vmQw14ifR8UrjzqmAcvVy9q
e/bOUgvJ+O3T8Y8JVqGTb7DRFk2y6b4x0541jYq0gR+95TKIhApRoiY3EHs8pJxyQ09xBByI0RzS
cSzmTtT7OZw6HNAn2wXZXc9iGXdjCDsfZ0FVfFTJS6GfgvKafnsjpUDTBbJ6gnARERC6zg/+I2S7
OplYnop0xYJTaFz3V5vCZW9qY3+ojYoYgUU8BxQM1cYUl/AUU6cyJzynhGRnOq5BgD+n7jGt5knI
858emURyTX8FdtGKOisM5rH4YQto1KKckHCVBN/QYeXciz8l0G9ICbHjh1fFUk73nIlSxvyn/BLx
nQ6O1vSjlQ8CnBXeT6/Q83LoLnaN3+UUzWqEnfqzM5jULymHyDvTSj/YkPfffqxPawvmiRiNdQ4q
W8+58mxXXUlyr3vFmvsGdEsNVxsZ8Xdi01wfA1mfEQmkllTnObGlZmLS2/Lwrkxg04Hkl6vMl4sl
/jYuOb3C+XalflmK49phEUVaUJ9170p0iJkTJQ11lqODb+9Cj5UmqUc4qZR4DaGILhkaLosF0/U8
KC3KBtOmItrinve25yGsDJEmNhmaYr/AsjUdefSnvqsmE4UpOItK79oAX8wEOBs/BJ408/jeFLEL
z/LvTdDF/f+GPtHlAqLUuGwOK5mkQarUqsbnBLh2UdD+o/a8NYZGu1P0J/jhhP+QFyBkjRiO0CQa
jOowb30fh7AhI/6VX7qXgXT3vFzWWp2Hpyzb4JtEwL+38lSGCXCzK+zbgZUq3kKJNGAq2oYYsLdF
Xm64DksjboyWAIdD/gTOHbVoppoWl7QASdj9Rk6Nu1F/MMq9f8LewhVX+0QV2zjhAGOnvlSXXQsG
2gHOG5bcD0b9wUhprsBVQtsyohv5X+TqPpGsRO1wc0CpgAf5A8sfenYYGp/f6xcTYs5qC5imE0bv
XVu+WGzMD9ZH9+bmyvrR3TKXDaP1CjbJQwduIZaWCsLnfE402aqRfRTTzSZMWdLMbovAc7GG/MEM
0cG7HHJzWk75CJtvjrmETGT973b+SXxgBG9/1ipFwzWsL6gfxIJO6SHO6wDnA63Qp8XXsDrN0EmD
nwujgAkkU2NkNKJVuUU1uebnXHYHlUqHXd37Sndrb+u/pf2W5xXCqhU0Nk9NGU3WJ24IKPRNSrv9
cuHKGiCWKwHelKYS8TkBKlEt2wyh9NSo5NjoXBsx1feZ1t3PP3mvjXQp2uMFtWX0eTNB/spKJgUt
5v/IlJR+E67ryz69JjtMzaTkyod+folEwkTyS+G84bTyHdRwFAN/BRP4lGivin+rB3/Kq+zCdOir
dwBgjJ4w2FrJ85IBZVimqidDmz/n/ACSO8NpmPeV3yPybd/l4K+FY4rISfvBH+dq5+0M3ba9+bTq
CLivCGr1nNMMC5UiQ/uufyW1YF9wq7vHy5QJv6PgAefHoXXC7o6kiwdhe4pR9tR1JCcE62nPPNad
8tnHt5P81+QkSo6/nxNw/ipUWf0gvMP5I+8EdfuQXKrxdnAmponcLTyULWYII3hl7ekb2m1iOWNW
gqlTW4Qw9pTElu4etR+wtvElGmLsEAZqF8pecrukQsB+BxGNcBUpArrUWrHHlLIi2We38cNP02RM
3dKSCOjxf4AHlYjz4zin7DM2P3PDSFMBDopK0iGRkec5bw1k/I4WDeRGeWcGkN651H8oQY85olFa
yDuTl9WXSKCPMfnBeCtf+9OdcPsxyCeBWhfQ/RolD5CctBUoiFdoEK27fvQtR/Kq0b2r9tSuvWHN
yFt1a4vDtF8wtGSNfelHva2AUKnc5nukQVkyEvPN+sA8pH9nfqCwrVATw4n8d95SF3stCqkrP0T3
L2GPnIHSuEdzwYMSTUuMeZA7Yfdi9DPnaBCGzupSM5R5K5QtAaoDDftFE6ECGPuAO2Whv0Saj9nH
r7iXDkSpdaRSKuYXwfu/Y3zZjGHm6kRFyx91aCOWV3Ah4MF9dPHrsJv2Q3oXsfDcYgRdoIUryyAx
mKOjOLdN4GP/ojjpJ+WAMUZaqlxctzBzNuZdfa8LV47b9SR23CVzUKRkqkU2X5iVLTShsIqqjSAG
c6gomR6QKog9ClEaZMwgfQKWv4M6PBSEbrvJmbykr/nZw4jXKOTvvp3QaRpVt+eqc/1NbgM9OZXp
6yGcgrVZ+LdQb4gI7HHJS+u6yDqwd+J9yl6a44ZdSroCCLmA6sspoDWi3VZM1LnmxFum22zEPQun
i1ZYONm+48eK/uOn+FonBdv3eoAERp/xcfc00CAlAK3qapmHJpXsmaPd9VvPFuqQcJiEcIweSift
15KTIR3uaBgafKLET0jr2PGfyaBCuK2n4bywEoEUq1pUuZ04i1Z5iSIRk/4j9q2ASMYACa1rmPD7
JkHWV2m4w1z9mGgg4Vs73XDMuqhBq/JAwd57WWRC4gE328iiXLRlmz3oOJp30upHEMYni9pbEeIB
mBKVWpTBAx5TbYpmG1k6LHoHxJAVIeuevqoZp6uXay8psk9ScyDTKgURaMzxO8szWW/P6fLTQH+1
tnfRen5ZCcgNi0dIDzW2miBtPigHOZPI1KJVxhLqlDTDNW7ozYfYwb+9Jfg9jnZU0Fj/lLbEBJ9q
UbKpEz5lUQ3d8KoGveG5yKmX8kD4tjQ/K/kBD8ITtn3PyAust6guSBLnQD/VDBBvETE6z+FIYnSo
UonFDaAPVkcRJIi8KfPy6kox4NPafNQ2szIsfrYbtLcRcsTs11AxFZH9wlh9mhB4yyiN/PqWr5CF
EzxNuizSvNq++AJSK8ydl1YmvAEBEyWxClLdK5bpOwxkYULABlm3hOlTO18g4RGSrjDO9fwAVJ99
+mIGq34XVkjhg4VIkqXWl28ybKZiHNNjeHego/F9/8d4Zh7c23+NVV4nY0dqfd3YQSGELoAO9rpY
SYDwV+4LSGa7qtW7SAXg1fBN6l03JSfh6z3pBcnMOoQ3XHgLrAYAlFbB+p/C3XP3tbK1McWYwq1i
HFjP+dbD9TrRcEhVeUEREZggGSKGeGkQoZ+SHOskthOaYXgaz+kZPpHHThzLl5vV84Gd8YK2w4GN
ovP61QE1aSFxNMd7IhRjKRHZvDJGEalB0gaqmcVEuI7F9KeDUHDhrV5d8drijrnCznabGxjehiBj
os4chtD/B66dVxdGrtmU0R6jkjrp7iYDMH2KQEr2fkaDNEFSg/dGhRkMP8BGl6mGNQcNwp8LKSvb
AdPymxlLgzI+qhpBlgShMN2mCEOzRfzBfssIkkXTdf405aW2//b82fYtOlWK7CcyL+57XbYw1hk2
3g2WXMrglCWozxoxYUJLmL8gRnF7OWTr3oMLzzjaDNXp0oM4F5fvHbnHgNCArmoX8FGcb5OKQwxY
xohi6KawARi7SM6tYbRDgWCWoe061tztDiLJQCZk3i6ZHpSsLkrCeU8+nCN593VF8kT0wsDMEaCg
1ouA8x4Lovn7uEAL8913g8mfytJzsvnRbk3o2G/5x/ky46wrqQodrTUhNy/WeWIpfUlt8nGRQUS9
Y2J3K+/x/fS9tZzFFJtDPkQwoZq25xd+VtaGFBeD1XUcDN99ln2c1Ct9wLd9AnhgwD/xPfOzs2IR
GTq+kBvohUZC1HoNW2QZ5R1Wp6cPoI/rmVg39E5itA400TwnRcKjK4rs4p5RF0lann4fqoI+c2vT
UAGo5KtnjhyRwduMXE9UbZjXc3MmyYdLWBkGuUustRBJL4BqOOQEXsEYt2KY32Ej3w2qjVFAu0aE
RA1xSc2HCm1TmE8y+cJ9XI8ikL5MJqM2UI6FvKw8xJeaHBTdJ2bGNRZWYbS/n3hUKEZyXmJAo7/Q
qNHk697kTBxtyBzbHVZ/q6sJzJHhTqXA+fgpcuvQ33Cf1Zbj06BwJlWcfAW0ZVxueLuYiuKeVv/W
EMUDw9yOXBV8TBB+DeAZHiu9jQGmB9f6ueq30t5nN0GqxXIGwlh0APOfJkc0d7rLDD6p3JlEyWJg
/rGMdT/FisCAtjymt2uYH1yvGVtW7U6Blm5lUUJRzV1yMbmPAG5uGuYCKoMtPGRLkaR0dPFpd1bc
nrv7LgXoYmipBevp5O+UfUldZypPQ6xQoRelXsUIZAWWJzJHU9vlqtMRXgr6Z+A9NB1wDgq7rL9I
9+HgoLb/pGdkeNoMh9oN8m08stkek40M+0BlUSBe3yak4D+FVROLeDx3dGCxGa9pypmThZHP4im/
QPb7r+asjw6SBuIdpfkivon+ZWPI/tyHcqGYEp8lB2nUSeHrgoaG/h+W77BoRwNP/OA0CnvyJSB9
rP4IA4Y6Dffgz8a3L7WTnwRN/fUjHQD4d4RPmNVnbqbEKAefPKg9y30YjUTUAnF/NQ8YJYbp/bp4
A5Td3Jh74Hrd+j9QeT8vR8CdgWZX/EsnzJH0DWus95J0va7u9F4d6scsEzyCshRa/gKblbI5IC51
8iniOXhG8zG1TRggC7OB4o5NDugUwXc8Rl/YQiA5BhRN93Ip0FpMd31lmlRzVei4H8OfMYhhU7fL
TJgYMPUHuVSgBFKqaSksKqDBYb6xuTS38WgihwjBle+8MdtNEdJPlFUfra+s2xKMpdrOoTmyTo4L
KzNyAOabzermXa05ru0PwZ27PCmBFTJQhqq1FBIK6wDh33sE/rAILjREXkFfvl+nShuWQqNCFvUY
YvYrAGqYsx3zZ4aDs9Yp/tB6NlLcEWBEKynpimLKL7e/vGX9Nb3HBUPt0C50Cb408e2Y08cCCDbV
BAjV7hkXlRZcZFEQ3U2khDflWNA28tjZPQr1n9OCFA+1l8XuLDSWqaOWL1vmh9Mf7umDnnxNKXGk
PlIYj5JnSZoo+CeoNtDbFv01QaL6lCspu1p9uFVBi9DOZjCK4ZoFP04s41zD4CDFXT2RCdkXasa5
njp7huVWcZuVBRmZXrRSAipARCSXOHgC/6Ubo0W43jZkwcJPMCXrsSaFhQxFtnpClu8cM2cthIbv
WHR1UqDLtaucRozMFPy+Pw6ixhS+vd9GBhs0xhTCEki3i70fAgDhgotdMECHhM1EHjGuM6S8Afmo
91XdRpKuZod6Ar9JmvPCrrj5GN2++ysXHpzYhrJMuZPE9UaZvg0qUnuETZEkiTN2BVR9h+EsvafQ
Qs7eqpDUSayIuLwQof58H/Ua1flXabYO4wjH3PTKvRqHTs/J0uAVjW0CbYlA6E+tQ4Iey3eO5a/0
zegV+vFQa2VfEybclFnBWOqCp0x6tRnqYIukR7+QNqiQlpaS1CeGjYnr/FQtOF5z00lqyse3l6hp
ZumsLGEy+52jnmsq6aM4vEDKTUQrvVsT4qhI5/Hn07Vdl27GPNNwgL05++Pj1nioEcjwMSHbemmF
CWbR7sRODTdY0/i0If+AwFl7Q2H8RAzg3KHvVUj3WCouwYYnpMtTrIZWZwKeQfT0koUybXQ5oxAF
cJGkivA3JGfP7YAaCNK+r/0Q4q9kvSfC5oAiauBb+MLpZpAxN+eDxXa1vZ8yDCPsP1odoWULkLGk
5owFK4q9v2G9dXtupa+Ix4sztljnegc9y1aoN+8NarTIckJj/sPBWRlqak6NQ86ETnLZqLEjcc5N
+BLDcp3aM+F9mJ3OBif1NSh9sGfpDLLrJSZ0zTyDuFPasAKeuP5+RDLaSyoQvwbcf+hp3UVtVhaH
NNPlyjUYS3gG01REip9MkLzH6sd5ndi8qUiKyhVhcUw4MyjSHL/K/on7yvfOrvm3P0DzqDSdhF4H
euTj8o4DkT1Ffw2dKPow95aCJla/20BQAAnTPvicGx3AV+1skgcyhjoS7VHHRPtRpn/wVpU5bg4h
n6Ip2Y2TxEjYyPbhbeuQY4FFRuCpukNsDu4UT7PMjtVs7sIj3TzF0p1DxsAfZ2ed2XDPuFHfQnVU
+M+IjK1javubAl33SlwcHn3DjSVCbQJEnFdXc6VtWuqxAEL0XYo4vw9A2kz+IT2C02A5KeejIU+2
SW7XApgTfCUuxXmXCg0iCVfgusnzFmdjMQIf4ng3TSt/tt17IQH/ZcdWY9B7k69tlhMdUHK+PDmB
r0eIZr66w1ioyuvzXjEJ3IJg407i/pPFWe2185EAA01WyPix74z6TilrfJn19TqV4I40Yd1J+qAC
hlG5oJ7AwZTmOccom41Qvolmn2avLCNzHDH1b1xk1q2SzOZY9Jicxsb/3zy6ndYL2HKZq3ywFBgd
bXUdEaySn7Nd81QuV5RmHnAq+VhUVgsOYpxn5cmcTtJOP74SvS7Tn7inZELzS0/kGkanDt8XoLkX
6HEhciz9MwmXjzO0OI6IcbxydkfRkJCRuDUjgcl4V+wZHIZuJ8itDnaTqhmk0WLtFWQg54OaqUGg
PTXauwnT4koO6uNb547ZdvaYwg/F+5Ns9XTRLqzzcfJJHhN4+Q1huGOoI3tpmZkbRMJby4QwZ4w2
tbOw8hCMOHQLuIXOTuP7+5hpMyW4kl7+/5ms8X8G06gumIiuEBIhdJKfdaBCRNFkaucJ5Ruww+Sg
Vu9aKSRmpaeHUBWOa8QExz/5DDRZBA+mnuyD0yy45pgmWEedKwbz1mLb29WRrvFK4RHZDQPdIQt6
CWHejO2XX+e/MMhD8n3ctiImJ/KKv85fGZeSmJSWofZj6MdUtXQn7VmRa5eVE83WSUiXqhDHUStD
GxLjAuaukj+TFA0/ERLA/N6B1dXn9H3wt7E9/dhvksmjD8gYlxGqTmwUXqO7fGkfGkip3G4QrkJ6
iI+/2AsLsc/46Va1hlmv60e6hcBH9IyONlclx9/4VmXSHRAk7admmXfbv9pZ1cMApOjtfRCjlCgz
J/XH+wkOhLZwdy9iPfomHns33AKaQCi4RZ5t9fIU0fxRIH0huttLBr7QFimXZprFkPWUR3DB8npv
gjYbsmDkUPQk3flnkl4kQoZDLt22RIw53UVVlSo8HL0jEB05lHqiCBjkFkpQ4ewle5P+ufIwUC7s
biiKe43wOgUouVkaHbs8GY0SGPpwRdSHPd2Xoas3WNZx043X3RL9Uw2e5cH2xgwUj2sJcU1jwXmM
J7mymkb9MIb2XCpXSiPbbqVBtUdgbuin51QbXtozgFK/hxKoILCMjda84c+F1xnVsKkLJZ2/KdlY
eLR9mIuN7EXeKgD8+FBkk89gZ5pwddCFSsxzo93Wq7V/9FGpgarCwOEDP6oo5csZQ5L3N8QR7PUu
YMwm/BQAI0WebPes5BFsC08=
`pragma protect end_protected

// 
