`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
PcE5gsDZgvyoWE8AI7i1/7lVDJXEi/7qSrQHjjOc8hYHOv2VTDaG/maUPFGM69sRmOhy+rJIlJQ8
WVysV7BvzGb9UahuQTI0CTRQ4x+HRg/bSll4AiMcICzz5sZ5WMrMrONJFlh938UAoIUg75tKXdAw
THsIfPN76X/5SKjjj6bVUj6bbW058qyCwPQgWOth6PQFig/HKIOjzdtQ1yG767SP3H3Brewrgaxq
AzG0PtMOOBAz3UIxtzUsi/5AdMCIZX4Bl3pZRN1O7JKDFkZXMCPVsuy0joFjDtGGyljEqG5YQCdj
or0qVnHeBE1pP2qYYTlN5tyyXhCSpP99xeRqTA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4RIAJPEsS0n7u3OTQN9VBMTyXTcBqFM8jrPrxiFJfT8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40656)
`pragma protect data_block
rajWRfmmPc6MnJwDppJvk6t0j3u1MQGyHM2OWfegTcL+kdSm2h4uelQL4AVmF/iGcV7e9kSfgniX
g/GAlsNGvz6a/YKYmu/SFg0pt/YcyclALc7Da1jsZQSPez1xCY+/UsWNlMhhe+EuhaUyQymFCPHV
XYEb9LzGgvLHn8BhZUR8dce1arZQxsj+OaETiOgQU7Cx1bj+gO7pLhiOeZIP7MB89oOuCas/HoSt
2m+JxlYn3ljJT02r1SUyDnQSZJssv3VThbXnRpTY8Z0tLyU0MtWVKWUaVTmnzEz5FIQpx+zwlkj+
4zmVIohJh+JptJSTQyvq5p11aNkO3gTTrC1ZcyLCy/SuRkkYeQe+zeyd76n9rKE1K7FKJIXMXyai
d6tJnvfe1VGdDXrSYMi7w1Po0H9AmDCz5O9ObfWwwXJFC1RMBqQqC37E0ot0ojRb8t1sy7zLvw9t
/9pB8CcvRieus8tTB+bz6wwjDnAEME6pgjvnJ9mKpY0aBVWnicBRVBlYEntj2SiavE5KYaDH6LTn
5FlZvLv2ncxQyju4GhLLwDBN70o++Bh54PxTC+xlG2vqpABln+aCYBRXUjtAldYiWUbN80UgLCAP
t/+fsoeQ2ApRPkPK0JmauaIKCjm+L0bmAplGTbNBXqIdUvQnPq49+0KnHc874mPKkZduik7036tb
IxW0k31H94fPwTyuoPcYKi/VOyl5sByzPMv0dQTAbnlpoCAsLdiflQQr9fukzK3vg6hxS19o76Sa
PQeKpML1dV5DgT5ZKYoFuHJosXa6avJdz8HHsATvsBmw1jvKz+GzawGdEcIuxfE2xohKZ4YfAgNY
udze0/JpwAsGtIi3JEG+f9Lc7KzDtVo+7e0axUtpWWG2zchF7YBRjZ26kg5u4E7NrejsKmQn4oFZ
2qTRJZGb5SJ+gdQBQzowrZ6DlCm5Ybvng4Y+fKORBe4O+BxCB8HAkjiHJvTxpq0VwrUrB2IS9/yv
BT0mW1nWT9cr5BxcHY80c1SIh2SWvSjyo6t8HbC5zSeDNq/HCBlFXopiOaiYhaqw47uoKfrNcZxV
H0r1trD9ioKahpJlKwYaBRt+CJIqIENNh2VMLE2xWNs3B+xYwnsk/de/IOcj1iQWRoITUG33h5y1
+zkXUSFCch0fG2CfDf99ZfKPFae3/IBCbkSr3MR+cMlvRmTMWoS93L7LabWBkeZQ0yEs2Vjhq1p0
39yu13RrJCaP4ZrUCpj9h5i8+wv3y720AsSpLoy4NA43a3BAS+zCe0TSkjEMbqLU9n4TdEhxfwa+
ffSoSqza7OYtRjEqs9enDHCavm1Mbve+nPpiGcS8FpTdvkZcWffD6L9mlpP2wUPGN2WnUVrKRM/Q
TY/gCk3fFo4Qma2nCumgCMXS7awBbeUj8YaIWl7S6Q37vzsUiSu1KoM7QaoCLRiUWgkAJ/J9/8M/
Bdtlwp679jJ2BFSv2abT+GmrnxDeOeZf9MunvuEYXoEgcJcN/cuIsKxpVhbPjE6vwtcNiiLlqwVn
D75uZXixo69iV9uvHxjDatKPJ0ejY/qW+C4lRElxhuI0HkPAeQlIJM5u85bXWQ44phFbuulJFiN4
Peh/tWNZ3jrn3bUFQvJDcujr3NijU9lhll1gkJO/sOmzjIX1PRSrcqIFJQxDkwYV9NYBGiHcgSnj
pSkiyJo7kjIVF4XmGahILtXBpdUxPgp690OdaV9/jNg3AfFTTd2hR9xjIq4GR50EUeC3bgcIy9Pm
z+MVXYDmCFjsJwIazzpkV92GH0rhuGBy7libcQJM38vAeoFP1X7YTszzLda/3E46zKLf6KSvfBqU
EiuHUT9h67huXUNEzyFRSjrY7jilC4lxB9UAbR1Mtz1JtNi3mq0laantL+M02fG0Ruv0gio5YJ3c
GWEEoIXpLCWiXHMjGW6At24k3oclEG66yPTbSMuP9NFfKpoWX13wyBrPViRVdUARmxnpIzWdxVXL
4AfK4BSO4HDMMq63nGKpYFHD1vcNuMdpBWQcmC+Tck86+XQnBGq5DagaNzFfMrthl1bJxhy+rZRY
6AtgQfcQ9zUvuio61uAbBSM6BmQXBdhPPm0VeNty6ItzRbO4GRdKMS66/Tf3T+yDgo6lBhsqmr9s
tMCBzk/bJPppA90nOHEtxe4w8NgECDBuzAEZYkFaJMpbouZRhGKaNwXVnjY8RMc4hU+X87Qv1zo1
cLFwPwwgFxHI6k6VQGc0KKvvdNR9iK6YwqHJpF8ZTVSMY0oYaoeOKjjPDpAMN6RyAyLpjrRo3QSe
i4bsiUB5pxO4y0Qkovzl5f+haZG0gCw8aFE4IDkwAXlLhwzdkW8z0aqBlUOxeabL4FKPIYeRmntM
Ibz9Bo3L/xyqGzsEl+JUEdXCT+gLu3+FPrlkaZuLbhTQjPPGFyC71Yn9v2wY+CYA6ext7Sp+3Bqd
syRFhmYOsQ5pQWS/gXKTGAcj8jay/AI5LA2r1TToP+xWfGlQ5iHcNhiF1fJSOiZ8lVf2QFwOk+dY
b0pcKzlOZIB1xLVotGuOE6dLDEejIkMyQ2ODWEz7gdJBO0qwP/Be3HTwEqxQrRZeNuH/oA2QtRD3
WF/mANVkJEEp8aePN37MItwHUlRfbE/LFxeB3cHF4pk2Hf6CZZn3fAD+C0BXSl54c4loyCCd7rMO
Is4F+E0RtIQqWLfStcwvzstzr0Dref6Ktz8OhCI/Pdzs0zOyVrFtJqU87FwiOPGRWSXgKUPsmkUE
RfB4SItF4BSyvB7ngnccwkZmETdSXTm8I1GIFsJ19TIet3RNMofHHdmXfogHAFK/BvJGkn274hSs
NlIzXvER+WEdi0lspgLfzd5PuPf2P0NL15MGDfeEIvgfu9pMkNpcERvCJi0O1k380tRCug8aEq+c
zpbPT4RZWKd7gGS/dUYvsxhb2u+JBg9MMHKDmaq6N+iqoTZ8UyZofWV2uqtBD/EaHIvEQ3wz1DN4
XqfI9dHm1WWWcWA5Rn86bD0XflN/f7xwrfA3R0S9L8V5f1BA9Tv3+GfgfdcMhHEYY84d3KLHUTwI
nc+XD0EQNgGAbKRx0GzGVpVC8FWzrvuz8pRB+bWzDG8a+rGtkLyAu3oWvxJpQFzxm0MtWhO9S+M5
DjXvy5IgtNCURqdA0gKFqFrGk9FF8Nx/YNI/DK6m6fpV1OaeJGTrY/qs+1Qn0bH2Zg8nKiFspq6X
Vvv5i2Jq/77SZbr2BZAWY+95W+mL9et5vxBe1YmiJ4BdfTY+1IDeLtddpM5SvC9jz6Pp1I513hIR
L7qdrEywGLXf0VhHn7wqX7ooVajC0cqeNuPyGwAOOaNfnDmIzDf413uSTs0fzhF0gJEk6XRm4tZW
DOGUBOYtiaD9ocY69EFBDKFXWMSSVe7Z1OzCNm4yGde655NUFvk2XE4gvnbN+bEAM8YvZBnzUgjx
3QWnb+YS0Y5Rrdz3QoQVVaAOoALf6+ch6SumzE3X1ztbRqBPdaPcWBd2O3WXj6kCTUWnSM68WsG/
T5s1hdL63qkR3veyzs19uryUlClq3QvM0Z3xCERFtO3L1gcd6aLf54d6i1HIYkyrEaKrB6/3Mc9Y
oaomct6d9C4p7HwpeJpdr3wY8SVKBxuRcdff0lI6lU3S4KcYKIg2Bd4/D1+tbg4B9AYPGw5cuRre
ePeV6HleY5Ioh6MNzKhnAdV2YUM4tAnZGXvuTqPdkT2cEgP/drNGJHdN1/y1nUqyGfSnXsH+eV27
0Xay7QxKZhZ822W1gvU16IsRF90FUSgyR/yVMJ9xf7xuSk5cXy/kSQ47bs7cz/jRwsxljNaY5HIJ
4CFMXIemTPc+nqBTws4CJF1zyvMjfH1bcqjWXR+pXEoxJ1Y47RQVY/ePdMZvWZCL+IL8r+eI5FS9
nkoADtUJkeEyQONVF1aVK9PiCfDR7WyWbUPLKVeP1XGMTVv3gCzJZ3QJ09CGAjOy/4v1h/DkTn2s
smO3wJkakybuFlIyG9Fv/i6IQHvtR/o2Ul8ZABzarz/UpeJwRrJpyCeVoFp0qszXit5gnf03skZ7
kbdViXkd3h5kS7OQgbDuN3QGEH0Wk8ykBhUcRSBqPLfnd3RADLOlE0xX7pxDIA0S1BCMPxQ7hjpv
bhhJ34s82LypEIwa0KM5u2vrOcd/3IVJ+qOLWlu9AjCE0ilgPEf1+ThuKaBJZTKgKUuxrYMwqfhw
dnuV9ZI+QChWuRX+nFZnv2WiVClk1bCOnhg/sHiW3HLCR3jyS00kLHK4fknU1EaOMeN3fZmpl7Kz
20oPZzc4JhO5CxAey0Pb02klBfVcVtqjHB6VQ0dIDLMZaZtuE/bByQLNQpgPwmU7GD43hRQRiWJc
QxUWOlNiPn7AQXPPNGhDjzRugfrgLWYPu+4EuwkTMScSQxxICjgAcP9F73vGaYB106U6PgCzlSNV
jKkessGT4954wRRRG6FUR3/rMAoPFXiOUV7tJYDb0b4D8HRhrVEFcrJwHjD4kvCaJEtPQhG/NDhD
cbCLgyJa3s/idBJNRCQ4dI66vITuE2yO78UZs/G1qxVdfGJRaRPJZ7g3pRqma+159pur303eygbZ
FpqVTGONl7L4K/25JKpZ0qvbvQKKfBxYaKpucj5X+djI/UTbsgrCH34Vi4MRnUAJSmcszbddsDo2
Tdgsy3b23NFx/fKkW9MVhRce4ipRWi8OD5f1H8y5uXRPivR3stDgAFhJl+z0NZl4tTXq/kar4Afv
HTn7+/gXeV2p7Jg+kWPUefV1UTmo6swk703adWctzCnJeMc2jLmoa25TlmPR8xX2YsP8IjY9yRba
3UakXvFa6bYWy5fHptcry4RSQQVi+cKmGQhBU7PJ5vtdOLxcHqhkXUl8c3I65Opl7TJZPMSgOzw5
YQNrXVXk3jkNdEK8IYBzihDqYE0B6bjIp6gunpFlnaBMRdfrbVktxV8kMfo7N/vR+diU0Zo9nY/m
n8RIGWcaDN6lc3Yb0tEa4/xHJU1pkM6qMOxE2wMqYfV9PxmXNSLuIEoF8mFjd187L/QXG1v4ka2+
5665xnr0OWwOCbKovxDAWfJ+kmUcvXAOEGM0fhgtK1NWohC81M6n7PSBIiSvLjLzut3nKPjB8j6B
SsFrXMZ3DPv/oganOmrn9Xh9jcZQXpCptWx3hVfy/6liTxEJrv27U0AZunh9XbvjW4sPy7cYRdog
LA7p+XNXInVH/UqY/THrSFpSNuizXP6JQCGKveFCnUPilK4O0NbpMvWvc6++YM2oOuvq1fHHrYgC
ybf9d5/OSBH7Kvi8s1JMtbiq2kmTm5TUqffyeMqo2oz0Eq7GnANFWt1U/cSG30Bp3qKVjRBlMixw
WkZRrWEfZXW0Qw7+sWscfuVL3aXeGVLpnOY8gaLHeLCzOgGH+1kz3bmfgl/mUqgBMA0BvvBIpr4P
Y5gI/5BwPmqFf7Rd56JR2MuZuWmVO2+cu5vP1Qm7VONdi5Y9+fwZ3s22mtqw+cLJZUf7SE2O1T7H
m1ONbQSgCKOesqE0OYnWdrdiZ8c2TMxO1QOryFjcu0acGgvU18GazmUygT5WYNU4Duf5Wko/vWuR
BU/DwxC9uYjJCISIkN+Qezv7QlIlZORGg5E1tfpps8swiolHDU0AWWG0R3O2jn7Qn54xYz2YJseL
KyBx9hNvEB9FmoeeZzfqSjOYq1ksHKGMZZQ1aK8OmK3T2pJWWT8WGvt0LFH3C77O2uY2WPrxSZ7G
5rGGSA+IKUTu4r00Md3pRaR/KseVfmX1pyjydUSV8pZTkREPhrU2S1d0KhfNxeNp0CQ0VeQDTo3z
SrV20kU2lzbDO8QMEKRbnilrIVM4AM1BTep//SrAFdGCUwBmpUGiVxTt9VzQhdNEtTA5iyBjxKV3
RhcNz3yOds/qwyZoZD0bOFi1pn20/J+ydEAWwPRKIeMsz49tigOOaKD8FMOPmeRbLsYnUwHHnc4m
vw3ZYmjTcEpUG2/1nGEKoba4/osSrRVDWunPeLsr8bIq8V4KZD7XF3hYb+0uXNg0pBn9kaTZa5n0
MoE8X/SSald67tuKjkzKQY3m+6yOrwLcWCkne/eit+nk2BD/yCDBqn32a0FTwRTK4Cz+gn6p5+GM
hG8s3MV5zHa19nWw4f+mTUO6mTKBzhVsSh4XNiNlHSXpM8ymeLUT1f/de/FYUa8r+IcZOn1Dkm0s
1TXO605458P3o952iVIOi0/bkIGCKOAQSR17/Vw62NZpvSB03RxCjUy60mbkToeHTJmLvk1Uu2ap
EnEv6chBBbN9im6rU6yM2d/8HKZR+7ehEHsVnrHagTCAqvbWfufXEWVRZF8nc6NPGQRIRPHIpkGa
3+mEcQmi3L7pf8jbICh2nm9p2Zax8r4q53gPeHCmIYWGWIVRIq7Hc8kd1hCftLul02rSFTsAck28
x2KOEisdM0SII7uuw+ursaFhTN9BQqGsQMfWzdQE2Hb8ok1NDYtDeRgbKvAkE0zTqYUr1zxA472c
8akWNqgcJifqm/0nVbkQv+NX4sp7a3yls9aVTJBHlylMmVjYaQpYjkXGNUpT6YC3/Xlj+jEb0Q8M
X9jGJ3TRLlduK9lOE1KDym2CiD1ORqF22rIBiwaHvNe9CgWCMDghF95rRV0W2QrDMusilPf3Fdk/
nPAXlmOgHmi+7ZfFLkNlJw13CDRRtfwedDY06ZuZsvtXPjidg221MEXa0ANXuaKQ5g+16IQFNILn
b1X8CCfdJr3Zj6dprb5C0HjTL7MhtB0w7vQrCS9Wtd8cJhjc/qCNne+D4roihEtr6yyA8AnCobdm
Qj0x1VUNOj4hbfeQemuvF5tz45X+IaB4hAa78FOJFvqd/yLdBJAt+B69j/cwOx4+QfNXmFQkCrAw
IjKkorY+7nMt8D9Nmo/WMVxNPXlG1ikqq5QDC/3h5n4aVntQe0GOMGOrw8Bl8NKTzY1d1qcu1xe6
usczWzoyUUNMfJXDE9NPvlJE1J1lvCZaZeUpgJOa/JCKag3J94bYZtzqDbADLzF2hvaLJIXJhH1Z
LCrKJYlQ40lLMwLgj33A51xCozHC0WriN5XsCXo5KBQlIQ39PTGaSu5kLXFrE49ENjYWbjd6R0qS
Uvi29AHNvcFgIrUTVrdjo3C3QVR97TlbK8Wl8S0N/+n4gaRqpidPHyLivt27j/5wP27hLgcRiJW0
i9WzvHEhpwgBzyLYRsHsIi5Ujgvf18gPd3r9snkFrZ/I0tANY+Cu0ESBQqszNezfRiBPA3hwj5uT
Ebj9KNHNknfhfU+U30H+KaWb2hQjlhPy8OvitFIs2JOeopPB85Tp4oLO/NhwC3cvm8bhFNG3NLaA
CCs/9zMMAsB+Iy5vLwrQuyQsNZsU6CHEb7i+8wlRHP7JtnACCXX3ieVw0ik5SpV57/f5plrfEASu
9SGVUuwiL7GJuPt/0oTNgvOPBCyrW9RQiqatDtKleB52J4wRW0mzX2G6BaBbR65WOGfkeSlmljt5
kY6MfsbQ0tgUQehm5aqbykDEaK5rm6xUbFhYXg5L7J+CjntMYgaSDzaFuN87JC6AkRKYv4egldJf
tBzuhl+PZHaV1jw6VNnAHHl1f1VzY8EYpXuI2GWgG+O5P/jmSYQZeLkPjCa3V5y5uvLrCsSbUYu0
1bBSdmDSGOj2vJTrsVM6nkCLFJHZ/8tjv9wFn+7QPPtuIy5j+0tV8QaciOJfCFJTZanR0rfT2JOj
Mbv9oCaumr1322dMkXQRdrsjsRMttUdYygHum1P3tnBExp5NNl7GklckwKNA3jNIjvFEPqtJHTcA
Gv/7u+LaM72UWILdCnTxw1HsxY5L3IFWQVRsELFoxV9k6UTf0TsVMiFSBPlPKUbPtnOsIMoxoc++
FfGDFaG5KBo6RyyZ4aalW1lfvOUzFive2bLy81dc6WP2OSabXukBi5RNVkn+La7sk0Te7Sy929+P
0fVHzJV5j8GYNgXpyR1UeB0WDVAnYfFYVTlrtVF4guzah0O+MZLLMFmNYrMAJJ5h8zwTrF7WFByy
E4Nlcznw4OMfIS7yUne4uyycBEn+STaDhSzVnKSEShxVd+hUQZpBWJGLrShYzp7S7ZRj7ZiXUJFC
wq21rIADzzpRFrloxm/QH6/IMirkVmx3fsM0AmIb//g5rm5cMDF9OlWXfKNwf9b01L4S87gsLWxy
pIFo0CwuYFTCthksjtVBMvtR3F15YsC9DiiK19FrnRzjDEAa9oOXrJKfnPjDNTvOFvjT57kkUnxq
emCy838+FZvgRulM1PUqzinAWHn6+l0guEJ54OCo+OlmUvJsE1UVtaSDgJ6voEI1EyKBU6wH/5dy
r1RW9kURgl/d8hOr0Uux2NYuqvttpNAdL7pc+aLPCao7HK/2qb6oLUbPwRJCrROr67gvmZzlhfsD
SXfuHDTrLupIWqkdwVDxmT+L+2DqpY92RGcUyPIwsLDYz+yEYI4alY/G1vqhuFnRrzJf7YEjPUqx
YYM0E97JtAQBI8lZHe7v79uO1Pqooc0YOehwo3FxEJlrYNZDOtgWHueZrv3WF3ktCp7PjaI8ffLW
1eA6+R4c1Fs3qggjG/21jgyvIjMephgMOd6Xb+HKD5zTUoW+N9D5aGPCH7gZPgSoUv6Y92dQZGE5
2MpmtcaxUg307LRCVP2YgkUiGAC72dZJt4LP6u0W7DO71m7uwRJz9CFCO3bxfarSuBVbuo3gVA9O
8g0mZc0AEXI1Hc2y7RI8p9gr+vA01TllnsTjkvwmWUWxghWNjy8LredU6FRZ4g87cUKUvWQmHOqU
gcKX3bxBmpIaY53SvdjazDe/n+nC+iHlrYICdNg0e+j9HyBOifsJoml3IXKOUzptjKLzf1u9mPbH
/gKL0vGCIH2mqwxaXF9RWte0FNMEqPRhYAj+qRjY70IH0AVJh/x6DoqT0YQDofwlnX0jpgzxBmyU
dTtd8BFveNhWghOvgLRrtmb5nBa39zzaKTDRsTg3czKV4/Z6iysFdZpmn1wuvMdOcv1Ho2ZHFj1r
YZJ90SNcBNJVs0tMlShay/ae+iXiR67qIrK0O+anMvdNVrKh5R8YfviUv8nYoUi9Gtbav4j2oR1S
qPBZXdr71wmP2X6sNE92nGO84WYpk3NCcjyeiR5U3ThujihHYFVBQ8NQDCVM4bMnvIQGg3tvILfM
5A0rJgoXk90WPffs31xZPpijjyFWE6ph12ue12ky4M5YE++8Rbm1mloAh9NcaRDNmdCBA7w1kyKx
zMU9Sd+lpxld/wP4f62uxtYvdg5ENvkdMV37/nIWG4toNOwERDo3ZnHkMZJQdFd935PgzlOsLjc1
If1hynTr2JdcNFf1xtmXCL5osFqcQWSddtLFaDdeel4JciPnPYAWrIIIj5wDXXTP3Hi0sIlSAiHT
o1gPQuw+l6/coOz+75Q/s85feNtVrY+LfewEXPsmzzaUCHIlQXN78pgBxNnbA3wXDJsJoM8Pr5NY
AjNYZ71cpJupxgYoybPw7vB+TkR9dVyZjKrFqk/3NCHGEKxVE1qQq7fTyaWB3KbLJ3XGHUzvT8ji
TQyYt1YfG6cMrnH/SXk7peeOsQu5gcI1p8/lRlb7p+4OCUd0ycN1owaDcT5KhAfbCXPcfQ4VQr7J
rtWqal/0JbgiHxRipmcHnyk25cxZJTFcF9xVaK/Kw3OTrLf+nWrL9ETPmL20s9o7ZFBXrmjvLVq1
Xe5hdEEVYBcDmvPqT5TYw8ulHjL1tpUoF5EmgCFRaX8T7jF+FD3mYGfdX8UaD9h/324kzjq0cp9C
rC+wB/DNECXnY5gaJYfPYIdJlZuK0UZkI6sFOCmficgpUUBRg+iLSX2ShwU3XTFmej0kb75LVcyb
1o8MoFKEGmHp6nONYlecPp+HnZtuR82AoOFf7Njdlqodk/qYv1fm96hxIbcnxCSPot3zymEa6zu5
UHQIpYFfTlq5s3z+dF2JWa7i6RrkGiUER7hVomc8sTwQZPgLe/r9Dri7t+1hHk/bf0iGrseHHD9g
O0ZN4tmM6a9wqij58xF0wUqrHG9euFC7nbnJN7XpRJaFbzjRNFT1PuRsknWm/ghYCnZyBnikP62z
yA5ZDljWFqx5DbAbnjqioxQWauoQvYdbjzmJfwXfPzRX1epvU6Y17efuBhrtP4bV2aVEL+ABtubR
HsR0Z0xAzNyYtCDlbnhZ7Dv9/r/f/sh/nsUzhI+ixpZSEzPwHnJLC/oN3DXvL9LIsINoekuIO/N0
+iw67HAqTAQJEZ2qMlnaoYWG7X7vJ9co5b8DEjiOecnAZqMlG6hSwvOe9wnmIQumt8E23wo8Qp7B
PCX/i9jTfnkr6lM78H4N8gEx5Fl6lMP60qV4ywWllCpvn/glqEkG1dyWnBp6rjfPZLnzaZphGFKQ
sMbqpbHo8Ee6Q3tOwXzKKSfLbmjadBpuF/2Oz3YQ+vfysCkhaSiChFW36hU2FFvb6yMS3acG8kBR
XKXGfF3RDX0C/YOiSM6g0ArmmCMz3kUJUW/0MN6cb8B0KWeY0BHccqTQEkcuHUvz7ZBN18qBs03J
Qfam0IbiaPOwmaen8vtfSVapjRQbHEBA7yvthQvEmtZE7AgPRAuwnnlVFPO/rZhPtOET8hBXdesT
D+KlNo6HbnPYcN31T3gsW0dVpPGW3oXBqfDR3x1NFo8/41jBaR2Bsk9HmXTNj31OttwGhilipNlp
auqk0NA8lIL95sQ91L2BhNeg/op3yNhbQMJUma0EfaF0oIevU5yuswkn0HZr8lTeb2PT9sBooHD+
3+o8xhEPnM5B/oZYDxG3nY1sZg44VGGmxkLK8zpg2Zq3q+PUF2/ctV2kBGJgQLJ+gNv3y42X38tY
0j9LTeZT6Vxk+PgpTlMi/4Gjxlnz8y/0hcxy8dPG347wbhzHCAyuwHRD87UwQ+7mHG0PGVaQDbj+
Xe1mJQWqlQrvx7W7+l3VJCzuINm6NqRCR49lRG+oCpMb/GeU2PZVaGcetNweiJZStSWbf4HUOoqV
61R3qUA/iCWlClLcmgIDb9ucWCYXwgcZ1hxjnjRa7i+bXfZFrAtVT71ZxXxERyp6XTHTB/D+0Dgx
L3LaupHED9gx6llbTAGffETOsPU+WlKMSe4e2u8n7qGdMeTxQAs4l0w4PL0s3coCeYokMPdvBe4y
5amN4f16hk0C263Wa2HACBNiViXVl/KTPXODw1+XfrDUlHXhDk++uQ6Bvj0SgBFku0Vn43CMfFBS
zmcCjeRUXzXlCUq9ujRe5zyXqR/IGOejhLKBlqAHg7P4mZoJtClyK0+kuttUlkVWvDjwtIKxVwg2
kYtgKuNqJmdKwu1r1g7abs2MmZvDBM6BWEyPysLGWrq+OpsbbUs4hrnudpVS+YlfRUWeYQKl5l9k
/KW/HZMDTtha4DPdJLpX7c6a4UXPBBuRvgJQhstoy1n4jCC2MrVAnI/88h88FwsAkwf1YKE69z9N
SjPrUm5CV8gow7ULTlB4YKUJbntku543xBxcHGGp+jKSPkGfqGRFcF3SjyuKhlVGRJl+UKSOGQxC
TQHwRguqyFqZyjbpl3Ah+Jb83n7gA8wwFG+3OwDKL5WtsnsZldu0XhlkSAJP8xWfDlPcLzoKkX9/
SxhUyuax7dU7lfQ6lGKGo78nCSl1XYs5zXwUUUK+/zVydNT6Sffe5hGT3sk7DOGSBoTdXSKS3/5/
T3BtkWmgmAJDkeyAZq1NWST0HQlcDzvKX67s7KCZvdUf1KBUoPaziTATRw3hA/RQxDoHThu5kqca
1Qg0ZyGW4jh+mk/gFvZIi18Zv9om1sn/XMxRBIM0Vjp8T6g2YP2LtUXO0EO/DQpUkSfw0Xc68VJd
c6seYaUyOMfyixt2zT+PPTcM77+wybrhbDu/7t0W026sS0tKGmlJ9sF1rkrvFUyOGq7jJZKvDZV9
NhrHJ/TJ1diSTMcFiVkEOqRmmEJa2iPbphU0LIM3FUL5vGhUzbEJlSogV/KUhCMW82Sv8KzTE5SS
6hBpp7TurVqZxlW5J9qLznzdp4NhBh3YhNZv0DgBSZlr0lD4yKT2ztLw6SKwIWX6sHrXjfVFXbI0
0kHCpS8t2tF40An/ZAZEes0HCaw9LpCfOfevpo2HVT6K1VfP8WEvL8/L38Jfj+vqMHOA1q0TaNjB
Z7+d6xv68hglJY/ohfM+MLN5NbXS9i2xaYBmEB54gx2xcoodYFnAeSv8Zymfwws6Qrv2UpkXBi0K
yUexzuZKpBvB2ICoJm24n0+k9kxKJOawIzR8lIVxc/HHkTFXMoVq7ZFMgIhUwHZdZDsNeBbgMXPs
rsDmR5H9iyQ7Q9MfnljCyfMZrcGGFUTs7MNJCYsBDWwSAPAGsuNkcLT8botatjgm/GMNSsHam3AH
h7uQZMKRZHDVVKH2YNHRogoLFWKw5IAycIUedCmNGFl/iE7kticmhMreu+ShqxhSNL9TFcyzMepz
nv37ogOMMt10fd1HxT1+Z7AHhtHXqYPQQQHPZ0uxUNY2HF52cS9+5umWPCIW65UCYmyJzsdQdrPK
kpjGN1s5IiCykVYZ/rtUVbI/q0VEPTQPrUju/0XdSNlEtAeTEmvYMxOUOoOvlJTfmWYUx/BBloNC
ooqlMlqB7K2H/BYmFkh7QQtrQvFNyhrGc5994lS0p6CoD4S3/I4zLd9G3OWUUksKH1ZB9fONB0Ir
VwtjPWYjQ6hZKOC6BDPhWHLiARTp2Hz7HTn0iUtou9icoWU2hVKHp1MvKpmoBPRPeyp/mMkuPSDE
Jx9qQS2bcHETaKmhC7e6gEy34a7T9dg1fgQni1I2U9AMmOdmQoycfBUek9g0PhUSthaclIFedd6S
CotdEMHspy0fqlxg7HP/gS9Yl3rQV2l5dWa1R9ud6kD6quQxGutF0CS9mBr5ajFhL9tGiNc81ykG
6lWWqgB9GS8nnPEdjiUIQOvyZfIS2Ivzupm80e7Yt5pmreAHU5kEhQlbWf1FA7YPgl0DIsF1VHtR
k/ys6DLBIJ/g3mriEiUORUghByjKiwu4ZpqsuLWLJCxNZaQ61+SUL2b8D9KMoIExDbxMsNPv8O3Q
5xUmPQ/Woii0mckUwBmEqevp0X7FDGEiCK49OqWDLnIKGiAR9UEeTMOKizRfa8qleHybq0D12750
HEcKS6iL/JwcIjdijiDcGzcxPHAvsl3pCVpgh21G6mmVwvIIPoqZxXMrUAK46PAPoNzs22IzGbaV
pbJuZfEL/4UCJft0eVpX1TFMwg3PotDlSjhivDMv1x0njTbpl8P1MXd7SskWkbi557N9f6OW3Fax
pn3+yHTNrXGFU9VvTGQkJu8MhA20eL64y6ZBctyVS0gXx0u9WI4CrBr/YM3wsqp+YrOHm+otKG5E
dj6CFCGBDtQZDqxWK6FZoNJhoBqjw0b2NWuWMC+G+Lxia+00n/7YgCfOfT7mQ5uygglnapxdOBRp
KtDaa2ja7FyGViaYxMv7j3FBaHGBAnA49585Nl8qcgjVPY+7Dyzdz/QEgxh6C5bUkMAOPUWX3uF8
wRwTecSvKFc+w7rcgHUhdvIJVqo3NXl5DVKsJIHmf8zGd2zSQQn5rKqQocxWX68HWN5/VpMzQc+r
6wGaAgDYwBy4w+4IYcOvKH7FVO1XN1w8ntwGfC9mEa5KnmgN0ZZX9V/Uc55LQ2LO0Gf5Sj23pUWL
15QlOeDkQZks2faNzjz9X+Yc3WPVVo8kl0CCkI6MMXo5KhWRZiWDqvxIydQXQCCdkpA59INzMpcZ
HjDY1IR5LPUqk7f1TBxmHTpWBkux3JfdYIlX6KyUaCfhCGKVD3u7iAmuiGN6N5lH3jMZc5cbkRRf
mRDr6pO2XXuiwikAA6UUrl6bPw9eFf0oOYfKzN+YErZAxaUevoA9s88xclIEhc/HTXQzNFRAJ812
Cx44+7ralxC6mgpwimvKoJ8p/DRW3EgUxVverXrgGBUYWR+YlfhtRtRw65vNU2kr4HhFWaubkxn8
jdicw+w21lYJRQ9lgF2fhVbf2wI6CbSceeQ31i2UJlfmr79twnHinPPajcxWxwWPYgZnFobQhKrB
rcl8u98D1UcV2ASSLRuJ5rTV1iVOLl9mi59iaWYT4ZvS91qfVusKjckvq7mQAEz+9mkCjTCL89Tt
6y3/8239HFE76/wVqoNp04fEBEyDrzBCiv+h6PAcGdEd+OsyYiCQm/547cHulzl52FLSXsl7ZlV5
8XTDGMvJaALQtShajEmeglA7YPcN9NsdEe3HTBjx2cI0XP396anjvxYm93BAgcZJdrEdXHOCVc2U
BAe61Up2s2cq06ZgamnFK+fm83Ff425FL8ChI0mISLTwT/EWRZA+cZnUvYFhhzj5cnVTwH5LPKZy
9lDJyM3HelCQpEsApD95IaRd04qxQCnEEtkvE6sg8OucgCXSm2YUVqLk60ujOeuyyQJUKZr5g5Ox
nuF5GjE3XpQlkLsllAX1CaoZ1xpJhu29PDkS7Vu7wfj0uaCmMTSRwQeON+xeVJFL00fldB1yPBd/
rnRQ80SieIg//sV/0l/oIA1SNhg3XqTKpYoPCo+zSrNViDc8mRF1AHpzseOMHhrF35zORDrciMd9
m498rN/+ZV7lhNjTtybTxK1kQZJW+d+pEr+gYcYVbTpJopJHXzNs+VNn8q7neL/IGZbBOcTvXQQF
KXnkcVJqSk6Yn26H2tKCPFjvSh8MXbrhkV9RTVLxxOaxwBNTPHDDk06zZaq5xAGN8WVmox2wQ3A8
h7I7LfgMDqos9ePnN7ckWlb1EXTQ7PV0SDoTCgx2CmjL7LWxlpo069ue5bwc1IFyuGZFesek7kWa
E/bhyFn/28dreHjjVwixeOFBaYc5M6ItmYqh4eo+76OP7Ew12eoQvexzlKFwsaERWEwUHIVJJHq0
hO8cqUDdoGmX5nbw5TxqjA736Ry7CeagkZWWec1fl4oHjgnYWoQMMKhto5oK1rXGTzTsAJATs3hd
AeLELiZXefFRQBWL5+NmSgX/vog1NwLBPhdaqf+Q7q4rZgWFf2V7eJz/MVHCqk+8ZGiGBBSq9ctJ
pgzcDXWkQkph1NL9MCLddudE3gc4WFVdOojvNZeRGS6gW/EXQJDEsnW6/u5pcYe8K9zcCOuaeerH
ZWaZ6NT5bnTrURk0fbDkeAfvAoLKJc6lcnmmrW+Im1OnOyru+elV5rFTgr1JzgkX/2D7/OQX9Yny
RJ6Ftk/GT2E8nCIVLyNEMFvYncjL13YYeYla05wM11e2qIo4yZzBfjP7B3Ssier/1JThQ58Qfj2F
NxfR2u6qDn7tJwEaol0KiGAfz3PeJhVRbNJp2Senz9ogbXQikpeQ+UpR/9SoHxj5k9F58aZvkD9S
WKLpB7s0mSqJu3gnNDryHF427oIuuJBZX2VeTcL78QmnqLz0D5pltcq8DNJqreb+zEWG2qlXVcyG
JeGcqneforvlF7N3KFZfU3AGjc1fPTBAEWYYJW2nS64wjZEbXS5f3t0UyUyipaRM1inSaUbn4EkD
4zAtT6f5DoZHwwUzT+di8pdFeDH4GHNtNplByTRFfWkZHqZXDFaVWVX0pvA8Op93ldJ+M6jD1WP+
/CLdH8O5CYU7PjHCyIvemVmdQMEYjKsGudukQSEhXoSQ6krMXTXXmIosNQOvHxAjim5w4HmX+5aB
s3YvvWqT+JDUEIj9yahDG53J0PLTwZakWlccMseyBdsRIsnfgphdHAyutNmOfnFePKVfvKdC98JX
/AOQy9F5+ze+lUX6nAqfpiYtvIUr2Lwe2STGzQN5KjBjuugKlMelm/TAy2yThc9KRtYa6AWDDH9O
w7E/IigvOmEJXwJv32d67iqJsE101Ule6wjRyeWewsNJ6Wo1Pk/VlOpJmInQ1B8945Z9AacNoM7k
geC9mda+Me96nEiUF/bEbndGos0oZKkwEwASTrE2t4SVr4QgtV9X9Z0DqqPy8NrDQ9QZauW81Jfz
LqvDrM7o5sliiclosCktwS8kPYZA5F2kOgKg5FLWdWIsP/ApN3Nz9XVeX6jSpv2bZzAOsnj7P5aX
PyQFSHHxhYb6JabUGYKiWQDbKYAtpkznRLJqUfACPYnlXx5+n7PVCu3N1Ktc1693M9Nv0zhLmfQZ
HOJ8IhfB9DpBNIBBnJLMQ5VohyEJnOFGCtarzUoLx9TlQL8bh/8ndci2mCxJ/FFlQMh+AS955xeD
zLgjHkbaHK+O2hhSvkx4M7JXMrmh+Wb5ksBrxs7uPPwfAnUPpM9UPPwsEQyXHPe7R2qZbgUnuq89
HLRnHfraYkrxAzH2/6P5VJpp6eqp0JJXmuU3DhUw2kyNog6fK16T4zSjVSQHY1f1q3MsrGSUDDIJ
nYkcmD6FHmmO6TlEP1KZcf12D4MmeV4kLvu98AvwNGVXS4My9XDqPKeLt1k65RZ2EeHVRXggQSA8
9R0jei71dNtJCdEltLX8dhK1j008A30cQ6n21iUZj/mCxoboQmdThEMeWmVHpKoHFTZxPrT75bNz
4/VxTvWf9igPquwctalFsIuyNnACZ1i4WYhWHK+k0G7oEKzyElUPIW4gudBNLD89ApkYNTeikE/B
peZzxXWiYAGQLJpY0fSXMFotTOV0ZREIWL61N6T1U8oftPbEo+3zvZ8XpDQ/jWZXkakyLvP0fd0x
xOXh38rbyqPzM14wlGevQkv5S3B7VRmTcEbuBZ/2/9Ej80cYKEPFk8TPXAY2Cjnbx2adVI2oBOEu
5KYG9G368e+UsnqAPEUrT32kyZQggvqw7Pdnjd2rf9GL+RBxZlAup5DKLvdcgosW+jPLO+/pKowv
RC022PSmTUpWgpkldHm/NTg5Yree1aMuQuj+zZBma3eKP9ZItr6W3iowywo4pJ+Bfccqrc+cWbMZ
kqKzngTfBJSMDa535JMBZon8xvAuZuFiKJnhwhkoRNdOhIspg3aVPB+YfBL80nw8Pbic/8yfqXai
yr5ZlgfyDm2lqOCpYPRaKcjV5PJ8+f/0GhPBmMD/LsvT+gTBuzavHPgzeWpjp/U5JQqjXMxRpW74
3qtPrgQdCIII2bjEeGkMmW5Lewjq7rhC16zf0ArAjsIAJ3rhptmBqCGUg08Dbds1hqTEihp/1smu
quYoU2o/uYxjZEon6cGXJFa1ZUfqnswY3ofs2vK7SRCRO921MvlJsyaZi/R8I4hiZbgTp6VrMVNO
AYD3yQ2jmAKPhGAAGnmyyY0Vznsl0DIZre9ghw7WbqSt4vJXN/gqJzO1ouDZm6t5lwNCe2iTwJNR
x9RFyphyQR4MixC4Nb1txF+MMJnrSxKxkhxbhA2EEm6VvC6Yhnii/C0KXWZN4sOkH2oLuPfzhDpp
6PhcYXFE/8QM4S3jCtizVZEsEEFMg5iVKBx1cY63osnhvOxRZ9liFKuUqVDfoxxO/ENyV3JbK+47
nJt9kk1QjQMtXWcgGZ4ynXg+PknO4dteqHoJpmIOaPJ/0gvYBdqNOnEJ7qvOPRbmrqZU1MandP2V
hMjDcrcN/lcnCSsmObRR6ZJbuJhkw2g5k+7aXb/GhY8xZi78TWKWX3yINKQsxrtgjFnJ28rn90Vl
CUeBDlMpRWwKcT+UA2AFVjLMt3GxZq2/aOD3e5MiMXlZHJxTWqLimOMmNtGORhsnsaZSbYRrkOuk
P6iHE2/TDXe21pIZsqW9hQvc3rHPNHTGmrHjmMq/KthpqX7NpNluUARpbI+fWp1IqqX4JRg5tD3k
bcAUC1qdFLWtAOVMKpZcFII0lZkm3GW/UN3VyroTzzflwKUXb5976NYmAzrG9+L3OL6kVNf5ApVq
u3JO8AltXBJ1DAHl4ndux/NePgyfd0wnNKFYRej7pVUU/vkgGgdAhkJ1x+ksu+LLeXvpusA0Kzei
c8GscdoU3zuk45aPlH+Fajb0QKtHWwxClM3I7FfkbPe/xuSETLcz7DWUIy8Ie1Qy4LiBD8GKTyWh
LIqVAMpErAd4Qr1Lf3ihn3tWKNIZvw7fh9OWgwwWMx3wNLxT8hvsexxXzFV0Wr9iyW9K4tjC6H3Y
+QJJ5wvat7rnKPbalr6sjn8T7iuaGtXFgDVcS5fY7UkUI3L/B7cjxKaLw62M4KQYmqYmTApeOshA
YXdl/5+EYKpn8KpysmNdRHnprFfAMCMlYBpEaoY3fB+upCB1n19HAQf8wua1lZob4l1BjDeSc90a
luuRWcUIEafcC+9edxY8/qXl3fh+H+UV+F09bAlLBNrJEh43S5hh7NNZ0oIMKyfdbuv+BegEtoYB
JZYlpRmCe7nb0hHzxquuOZ1kIp7v2HB50b9ahbCxLCKv/MT7df4mSNsZl4hVAzg+z9/F9WbCKbdS
qLWEQsIY2aH4a3QXuGXuN80jX2ouIxa28BPioAXGB8mxtcZeT9E/iugKs15jxtF9IwJxrquHSRHz
ZQNf+7SHABfOcXjm7FV0HWul7uTJ4ugoqqxsfDXWk4Rf7T4vCJvkq1r5wFnJz2THcwFMnN6ia9Kf
BvFtYN+joXyfg8kyxylxn5Wuhe44lwrlr072uhU+0+eLonosGoI5A7FONv9H1r1xnPLd7LatDQaP
e+3HaYOi5i2olbpNFKkldkYJeBB+Lrlzy/s5tXVa/oUxfphv5lerZhylsVwhP1cUSe38fA1l/Bq+
Rm9CGjTYcqSGQ4Mnsyn/AGCtnE4UEMmAyNGB5QGujoa0KmUMKoRVAJH65IWkQzmh/hsml+71PjHa
9IlDtEWHjzkpIO/d7qBMkXZwsdE4vQgRfVDjyvxVVFWdh828nuWTzGRKXI0lazUTcfTmzvuK9IJ/
BlY/yTXfyhBVULVE1U5g6FrUD0aR31c8atGB0iWHOG2KVDhR2nvYWD+XR5B4Ma4mc/iuoOqCZMUj
MVzm55xk+EXnzAAxKBZ+0067SbZgw50FRNbH5BfT32FzlR81xu+x1wKF3wCAyRKdYJlLSo3SdcXo
TFACoXcKmKplBCTFuJeYqJM8/YT/fFMURzTXL8DazRICIS/MAoJoX9pIYHQjaDfDZ/kPuPQuMm7J
Xdp84dfyncpTMcWLO/A2bdxxuTPXHQUM3mAI88gi0+OO0Z7S2yr/BAKF5r/0dTY14RAIlOmSdxb8
WE5mpGe+sifecDPUanM3S8ojptWKlYej7mNeQ00/8ZjoFEnl+0sCw8O/nraPwisSzM2gUcZPo57z
cmwZ8hT2qGOV7OYEMiNfyCbRfwU0WvCj+SMtdH/b2u59nfGJ7vuzBEx19IdzmotZ0NNZ2/CNxqBs
ytoI40ne3cEQ0BIveIc3ZpVw/1tz52uXHkK37PFf2a6fbeNJoQt4eLEhM6br7ubRU4b0rLmmfiUI
P5fayO1I5zXj/+BGYyA4aQMRV8aBol2mlBjMy8Ow5MTy2K0M+MzTC2EsqZSa7bPuT8MCm3pQPg0a
k4tWHKZ7odky+tTUKcLPLBVtXEdN1S1g82HMcl08MruLsGj3RjGElXj+/TvcQ7CFYy2+Tz36PLhn
YFv5VsNylF1f0pgQCWqaZ9GyECVFWm5ymd4+egALA0OmqKmfkYYTOmoq/El6f/OE5Mq15ZvVn9sv
FvAkdjVQePUSkfw6HEEOE1stRHqeLd6Hj+XkVONTpq4N7eS93gFGHSDXSECjdigDNH8TqfGp2ufW
3RX0gNS51yAKrZEIcmJohkxWbWL8gCvDV054vt+7+ZTwTDU0vVbaw5ZGxVEMcCw43g3mtmbTq2cF
ySxj2HtvMwm90mJJoXXl8jLzqlPppoXUntjAsEHwNQDKFDLQK/lPAwvgNSMGTlBP6m6nof+mRm9U
ZTXHK71k7PvGBzhyrDitq8FqxNZudSARRks4O1sP+DeQx7BVkFW//gnCMyrz0+Ze2yMD7yxSYl7e
a31Nfrl7o/VKNeQ1pLXCThRvLpmdWoijdAAdz8VtlTGwovFb1hlVGknJeYPp43B9vIg/woJc2b7b
EFLMUkpc4KiC23vre48gNN0JFCFVkaxp6UC4gKEzUpojdFJSOUD10mJJL6I3VnADUzyHWsnKYTQb
pT3MWiysQRUvJyJEfuq4Z7Gk5LEfDwOA/A4vxVKbWFux9zuTrJRkxryO0o1Tmbyfly0cvUhRVKDi
VyhTT28J6X+HgyImVOaUjLsCywOke5ALAPt2/kSZioxcKZ+YUYoxPIi8I119soNe+ibr5DrLApGc
3BV0kljm2d7pKJfmq5KwCqJMSD4HGpOVXCiviUe6Xe2sjiNMxpX+flUjFFb8ppXEv9+lGmX2hUGD
+sQgnC3u85ZMKvo3d0myhH9VnqmhT8/Y9UmIjSypPyrPVOkwZ/wB07mf0NfWbT+jSgCi0E2iHmts
dO4JSumAq3CF6/kf+rvpbmOQO42eFeFrWrauPvZKcw7dtdMCp+ls3x3i5fLTYYiOb+nFJDMr7Vlj
P6RbNNnQkpANRjAga+wuErUIaso+9FbXIQDgAetzUkcumNLKw30RmBlSJI3ATmjerOTR/DXle1ph
FDc4M1eoZCDbzr7T5eD9oT9Y0AWdSh2G26Jhm52W96f9Qb4CyvzySAeifDFGHn4q+H5TLAFwQ0zo
XNBFxmxie27XZrgU3mIpz93R6zjMJ5uOgrze7XIVUxQaXzXfbBfG1VmMSXw8lE6L9brhQQ8nN2XS
dfs6CFMnAVRG/j+H+fZBoKwSbd8UHdNib5jqAyvkdhvxajX8RFGPWD9+QpV6rM6NeZc22qmJTxjd
cv/FlZC8u2U9DQbflM/Swk8VHKsppLOP+vHXRb2D46jq8sV1Vh+K/n1hM2jqAujbPkBlakszZBwN
UXxcqUAo9R9SlFT69qDLFsLh05/TpKDHAugmCTo636gHJ2LJp9nN2wq5E9GmpTU0NosKbyfjnH1z
2goa5ziH0lP22/cgGYC8cSR5esTST9zdDvSFm9zrxOSMMwc/8L9GXUclne4O2gmcobwmH2P6dIGo
giN0GzMSly8jndAGmI6bXg7yl8Ekvd8fzzVtEfdWPFthK39UQSX6zfBYoakfgg0ZB4qNszoIZA8K
1SnZOXPBT5s8onhtd3GAVv4NM6KRzl1sCpHadR96961agGQe5/N/fNRuGk55jnSV+cK1UUIPleu9
NhLdy1uSIpUs+knsBK25iy1xwG1PLakxDksc91kDc8l6kV7sSuy53IqQlvGtGFPAI8JA3Y9rqU1X
zVk6OMkGZbcCvSyO7Wq8jKMZmpDbUdCDEGkZkDLojfA9+KwVZSsNEH9v1X+NTFGRoDNp9yaWVs1G
+oHwO0ujgTmR/afdFiBQc4UCV/OXpeT+N7+/QamXXyL3I3NOYpOSyzlcm2Zkx3MZxWvOhwDqito0
No2LgvaSM2HuZHkF+Q/Nh6qOtfL0nZ7wGwCzYWiNFuD0oABgd7SdnWICNAqco8G9A/b/0YHz8xQ4
5LfhXTbpUlL8cgzj4y4Feyz3hgML0+KDjyoRC4G81aPfeBq8JE/nMj8AvR8aaNpsyY3rDflpkEhV
JgG+TpUZzaBXmqMNTtdEhfWnSmn7y4S45SVyLF7wpNoylzB9v165swfHMLW2sGD8xUgAJGbEZMbf
OwlA0/Ind05gcAi5+qML2bVxw+xOA3lRJWtYPwu976dBUXiR9K7d2wJ7QktLS9HPInmQdCZbXj4q
+pnBWwClsc5cHDWBzgaHhbHdOrNIIQ9jGGPhqVl1lEL80TZZ1L5zDKB1e+h7vZxf7OX3HBptmtLX
hB6rs+r1wSbVprtrtimYYo/Dg7/TRds+1F8AxRCORdLl70pQJZ6hcakc7Lmp7obTr+poASpkdssp
Q7KIYV/tj3PW/D/LipMuX4D6R2KdbKlCjYpbhPrssiB8yFI8LHMyg2Q18pZgvuRZzFujJ4xkbN80
ujSxjfnN+5sN8LNFmjFWSdmmmSwp0eupxSzKnSG3xLajGohsOwmnmGO6nLerhdwYWfSX9xAcppGa
4sJoXjRjyvUtf+vnhQH63mM73Y/vnKo64Z6pqTFBy0zNB8UMLZq1ZUJCNyrv8e1c7nrqQlwZG+f2
5d/vH1S7I1PTBv8wansY3I9vjILKWKSVpbdXffTqBYOsrxRdJY5zDY3giL8RMR+8BXY95v+Ziihr
LPQNPnnlA7bM+GhytpQurLjSOXR+RGqg7UnXMIYwdJGvkQuuso2Guk8FfqVELqorD+/PL3FwN+Gf
fME5Si05ZKndZkdPdHkXyg4FvAus7+sOfh/KBakUiWWMgF12Cd1CyFN5XueroWVVUq+c5mKgJAzF
vdw59w0EYzNRu+qaH925hJ9AsQ2kdkz4tIiAec1X1igJvhMJoTwcxv6NqoUbzv/C9g+wnlIbuBAj
LWwQPfq7E09wkkUUyjASJNJ6PCqJeJ1GytYENN5tdQZDdxCWmKN8xf+TNC4HkES4B3KhfHu/JeZi
0/wg7fc0GYG+IdJG3Ur0swR8rvY5SpzzbSZ8IpxONxI4uvDejAhigw4oruOMkXkt/vnRS6OVj/vb
ptPZG+jhzRCnX+odZQFjnNRCtLaZH62lMQA4B8vQPPO8H9CGBQIXdY2v478xSesa7eNm953GfaBy
DMKz0ogZNfd2YQfN4b+/drxqTk9fvGm2HWliJGo7hlweMsM3DH91AqQYH7pL90LiIyYitzNrHGRu
G3qs+iA0EDJuC8MCwgxOSCDaszXduGxUDetG5wXMnNgbEwQdiEN7zqevWTcdFLVZ/v0xs5gs9sS5
d4t3LsyZyUGKqxA5+zP+KOlNPDz41x3nm2dSTMOmvyR8ZZBMZap1sAxb/zmwt4F3MlzZ/M7Veh+U
G5WlxLFasbRFHE32WkEPciaiG5Qf5X7pNjzqN/EVMU6/7sABpWcJwPSy2ROdJAaUg4TIXpBMq261
e6qkL+Kgbc50vXIaj31eou4HQZPkC81hVlEPh6dqbcsVZpHkYi+90ON5mSIOa2BAaGBFUoFuLaHU
MPdWmOhAqxDHSyOiL6cWCqOZVVsISvFEd12HWzAgs9Ae9tQE7ChzZBAWuKj3Hf0Hmpnl9iEu+jFu
yxu6aZIA8PD+2swVLGSUgdtUQDTElgTps9bcQRHKjv4aWDCE1IDHrwC4TocG2H85VXuEV4X256t0
RkgUzioIQgIV8k0iGs/+wbMjbENsS16y7tbYiyWwGZcNqtlnUc+ukTYXVTMdf+pitXepuiyYWkx0
9mvaf9+q0SWSkRZ27BuNHRJY4nk5jU/oYM3DCqTTl9O7tEgVbXiqq/UzcyKPi+gQX/++sabflF+8
oaaakQ1zRo5Rr6NNvEQApvFzbGlGEoUvYShz73YDXa8C1AQU06sFPiZEQtpA3f4tZqK03+I2hL9u
PqnOL/PYfcZZRfBAWZKLUfqjCDFkeN96bXPEd6k1dWEyVMipglz4NNiIsXcpvZNNaS6ArpgTt7Na
NDOKwh2/XQfEO/oJDwRsJEdinvGHUA5DD3iAd76ozkM1hNsL6f/NHQBLeVRbr4D4fTgj8TaOdgRp
y3h3CjCkSBJvO2R75kqY4DzVMZYgf8BTmbm1DWUFfgsiFX0zzgqjU4+9nMkbZI6obOqodiG1Zb0G
550v69D674KvQ0UQ9fJZP/ydj3xESRiT9E99BxsdGVrJQYR930jCvozISBwDDsMvEQwKOzIkNzWw
GI0oMXdKV+iSj9GWaE+eHJbdzHhnFQ76hKx32oq9c828fbPxOzjBY23pIq/BQIrzMSEpFq0p0+ZF
GhjRSUqcNUchoh71GOTocWK87z7a1Lz6fZoIJvs+ejZa+FvEtDopySrFuAKb3q40u9wfDx0y64S1
akYGj6vyOe+9Mvu9I7jSP4Drv779MjwIYIjVOItcqiAGfPvdAzmiVI1iTfyBPSSiHi6+UbcOY9Q1
8yBeCEBoeiOg6YDWcvEzdPsN4qFpxg2Lxjszho6y4kU2CVXxm6+uG5Wp1ViiV9FHhZGZURcNTctX
wbPAvedlQVP8mQjkF9EcKY0AQ5S586rhG0algW7ZYGmRn3zC3GloK11gkgWngPCzdIChDVi7ocC+
KzmaClr0XNOg+s5Kgj38NbhoE6eQB5J8gngpXaVxhIZIvpuGenHKBIQePr2SYSDqwsAqxDrO2uYL
zDr6hy60CweUR3VZ11EDUJtz9coerF4HHL5TBxQGzcLJ4kHPKCwUFhofmlamoqenpAjMMXssmwy4
econ9lLnFGlwnazUB1SDIeEIPz4cS9oSFHZTwjuoi1pBDId3FxT9cQ4oDaSdz2kAaGmW7/n0YhWi
Faw/FJfCqxlSsqpjeNuHetNp5WE6+ItJ8Nw7BLNGvsGOtD89/XTKGa1ntLbsSxHaP5BIWgufdlFT
EON3o2ickYed2/gtRTuAU6SBk9NYeBa1HeWFmWycpe30VN93NdYamp6QtSmYgSYh1urCvIpOH2s2
11Hlgq/0uzuQnYWLKDRLuj1GOhpvRhdCK1tzPHhmrabZoW35f5gqOHTEhi/4azmbgoXUEsumjmoA
EocmeCgFZeLDwbfk8E3VecXTxToO+mYlHmpxFmCPFpLnXn5YZ+iLUsIybVbWa2+/1LijcUZHrsvp
WxKuLZ3eVs3TXc4TQfDn60IVYh8rg3gkko7d7GSJle38l9Vj0+e3ARFkWMFSRZgk5BNoOBDnlx6c
GSQ6518JOvnc+brf48oQ5E4876pN+LzeQIl/eW7sEWY+RIhRr/SVPtZOH8Qf/blk3Q1fflRGG5iE
LNH1kjAyBCrbxwRGXHO9nZPIoWQBuwF4FZKbv/pjojRvOEdbBU+0FLJWul3Q9ChQfLk03WLrJlV/
5O61mauIEjPpLzdakKVKFSiM0LVG/gTidqgs2SsFnZFxad2qazgNaPLspd1TRR0G6nKxc860C02j
NLJO5AdpQHag+errsTIH6hgL/HmIEppPt7axMLkMYEdnFU5t9Uplh+T1x1r02v67dWXi4LM1IYiX
HJLoygVR6bCvocvoafS4oxjpzCPup7mmd4vvsYxLWcXnl8tsLrBzIdE5kmuDsCyYwNgHTybdA3da
w1yEGGVFa0O6whuc8i7G2R577A3NDfbL37vyiJ9jrzNp5HsYSZm8TIPafNPC2SzSIkyCuHaj0hya
anMTha+l1zXDbjR43WwEzlL8ENvOetC8Zijmdg3mvRX0u0aeRi0Oi4VotR9jQ1WJDlK5iwcD6GY2
ZvzDBcx9ypZ9OC8YTU06kzUR2EY6E0/ZDDnqCZ2Y6y1uea+3ncGlZ82RDUQRD4P+JE20zCnCfrHD
28qanpHpo/suL6B7w3BPn5+UpFKKQXz5PfHgnyCSA7r10O0jxep5u5C3iZ3Uhz1K+uBpnJL/Hnek
lz8CISirnD1/xR/pMGCQX88nbf6wQOuyISqejxMBiCFgCVfO7y8QCmZxxIj4Z5nJFcrMB9I1YDlu
iwVv6d0xo/yKYdLusr64FyC118hCpFyV54XPzK4gO6EcfkwgPUkJ/oYdEFLjIWUMfUzZwaiylgK1
8EKvmoaJcaVknhxkKURsbDSRxbkWFDJRa2QR0ii5uYGnaPPzs1gJsmLf/zFSuUcYSPPMYhPTUdiN
2dH/3I2VBWrXQ0fTPqxSRTb5R4oZ8wY7zMPXVy40W7IUBe8UEDfKQBz3hXi4Y2Mb/fYKP8lmFDO2
+hWchdA4xiS5lHTN4RjNGWKlXkH2ojt802OlwYPKJfz/U4jN/1KdnMmP2RMTS0N0tGc4MzbscJMw
B2R+Z+xsBB+OGHWVHz+vGb7uM4U5Xox1sw6QalRgy8nX3Qg+PebjwLkjibOJBLVpsDUHdpxsmGBa
KSKG/oyK/JEf1JDf+eDV75BDXt9FG2YxBNuUun3C249zHy+xQJbrcH9nvAhbBX+Pp/ByhMn0Rbeg
fzjfyIrsdW1a+24ieAUPj7SXxclAKMX74cu0rsNywIv83UFf92WSz2jxWbyQZiGblsgS3EAH6dzt
VI7pShvuHnkev8CKV/IyGy0SKZ9VkG2ugKVCv0ulG5GnyrRzR9yVxWXOypWfeNSqwfHPbgMwWgN/
NLES8YgswguoM0OeoLjrcOD3bbfVoG21noC7Fsfeo+ejquROf9+pp1/Y5Wl6IxOjwD2GpdcOnER2
oX7yCnlL+WE/VuhN4PkCHWiYpLyIimv0+RE1pFcjOZHdoHXiEzt/J8mS6VD4U8xN2UF5nTDQBYZE
mtNFb9vERo9Ww1Ysd7bOcGFEZ/gn598U/ZikcfHOldkADnZKkVIfI4yv7HakvsLcUe86het9xQTd
9s945PQCqsCybqE9Ih7H5ZPp66skENIzbiGFo3X2HZrOI6+lHlPiYZIK8EpHWjAvycThoxvKmCeK
AJY3UWoIYUll2M//kC/QjoZtpHLFDZadaeqi8JfQV2uPOLOcpUCXUg9SpnB1zb+LJ1HAidE1ILMe
lvS4vDgRmuG+NNSWg0fcfNQKOtFc/SCXvhEPg++6jT/GUUc8wusSY+AGlEE03H9iLYZAoOHHYp6K
HEYh2fKD+oKIta3es9vlFygVt6ouZTrq10eJLwdAxf9qk3LOk+DLvdyVKvVei3PIAd0MIEGsbWUQ
5UtPWqruqCAM+1/qCHZQtszLDJ5hOTzv1vosPBmcDq1NH69UEeEAHZYOrieFDzCiwJVYEIT40JE9
WlB42b5ud3Uc87gqJny1n1HrZ6UF0X6KgRJYoCqsuw7hhmsii4X4Pop/GGnVGp/+PPzwJAjvnDB5
ZWQgA3Qm0FIYkAiItQaNMYWGMcmvIusck6qe8AJ9WzZZneYeb24c7Fv28i5VVv9GBOF8txYyXPgS
W9+hO4+4IopBQQlJg1lVazKrPEy/GmgprDC4OvwbN9vZDhi6yGwkwxDyAgmKHn1ojj7lnfHWTb15
vDeOjK3cFbuSsEMZSGX/nzAV8bM4cYDNACqcUJhwzZEpw0Dmy4Te/R9yleSOUaLeNm5f1PU8S+B8
jDULEutgFC421dVGT8wftLTWzGErGynG8AFp3U8b1b7SkngGOhP4/2sPy+HUL9lWklslwFFeBscI
jBdEyJNUgjtCzdbfs0vS+j7rY81L3p/PR2B8G8whDLVdP+0cC9Q+/f3TzM4jwCfdnI0G3msqKX08
vYLpSEAYrSRdwy4kflJKoHGhrL9MbaHz8D8cuEhjd9oHMPI6Q0s7eJDYk9CRts88Tls2rbZLpZPT
oyO/0EdcsY2arRx5wng5+rQMlnEX/f3tAlkbnP5kRDG6gzjYhLaW1LSQrZx+30zVT1atPMXk0P3B
JaOOX5I6/XWgufjwRVAomFQSAVEzpFj4797HBYjRQ9LI7Gm1FboVRWL4qZjlVA4uowyvy+UYyHMk
u/OjVw+QpuEwB8Bo3lBBc3HNOm10folprezb8jNC5PWwykzsgSEMxsUmPejdi9TUTNX+Kddm2al5
SxepNRcTzc/+NLKYn3dCaY5cCp/qSNTsVWYr1W+kxRyCqIgsB9FL+LD/tzi5/+WeWLGPeqnohSHx
ip0+OY0gI32zPhO+BIfWsKsaSeeiey631TV/e82B4JTwO0yMaQ9L9A4CIOvuJsRhrim/9aqZrHcT
njn8gArrZcZwkp9aOnbHYJtnxf6DrCX/vjjOk5EYiJNtgg0zDmOOZxHosZswiDRX9NdbP77fVgQw
xFLBALowWNkiQ56CCJIdbhZjEmE+M0Qg32IEb/4/ZkkMJLM2f5jk6bSlasA9w4pQBarB3yEf0kzj
k6/KPXzXshbgR8Jm62pI0nVpPKW9221GFKNPYC+rMv0KLzgQgxq8an3plbOH5uyIcnY92RXcaWU4
cEI4YH+7Ni+ExMEso8oWMU6M8+LeJtKsdZFaOgZ8nK1Rw8XTT7iI5hFSJT3uhRFrjcrhhV49FylJ
GTpieZccpMbI/QSoli0IiExtIiqRY7cZDKoH5DC/RLD+zwsNIeHSKvvjVQ6YU0VAdutcJMIVnrm2
j5VyYe1GgrRFz5Jx9B3RgiMBqp8f7BXCKlK+JXHMfZKg5+2YTgz87TEi+lbr+nzCtzLZO3mzwlWe
gtrxZLHPHi19O0r3ahCQuclUUXzO79UhocrSsqRZqtwzY7C00DVEbTCweIYKutS+LcVQVgUHRcUz
rYdiaV6W/nuacqZff1b3fHDtnT7k6bv0bNtidpnIBiLXH5CJaMZwTv+cftlD3HSpV95V5EkvRw9k
W90H8cMq5546RoyGzRQ/vCJlCn1l9ANkv5PZb4x8RcXeiDZK+b3FGBYkMPN5I9dOpWbSvgbtFLuf
w0Qj6TEnwKS3oXVz21oxMTAsrsXwUuMHO6mOcb5LpTExHt8Hrug4eBTjTbdHyJrsW8xFTaG3m2YD
6HZSqsSFQSV8jTLZlycOExuWDZT91qoUxhr16sqHBj7E/rgc5Gboiwg9eDiVwH9M1/EGzjF0sLpH
tHsBmArJb9GYeTTkPE5VwocoRImL5Vs8FLzDB8Fs28hUCbnyWmIFOskADKnNq4lqk2jW4H6sBCC4
G8nGborYqY7iOlsMCYfyiHm63O0WdA3lA9qGdVCD/g3SHiyBWMdBKrZEfk1x618gbtt+BdPaCKhe
83DlrKTGHsHK1I4bgwVT/SkZ85i4jDReW6yzwm8vZtS0kr7SLB65WbIV1TD8ZWvrM9QyC9exIq0t
oeg1HpoxO0ct32OKm+XY9wnYx0MSuZpLkm88K/qExUH7eNS79T/PMeaJx/nqp6hm7sesHBs2EHiR
KrlVC1+hBSntSPAfUyH+Ze1wi7cXfHRSSo3JVzJDAl1qQFowITF9rkbP2agcEe5blipn5702ljqs
pIKQdpSdQvc1ua2SnXkPNMYV2+EehPkAgF8PIH0xqUUK6YRpTO4V7H5XGrqWVaHEYIXPevEOZOcu
P0VWgIiITB1AQkFCg9duDdH9BmQzpG1UKtBpH60mlMoMn4AmE9uo1+n+xATuR7O0VL2CC3jm9fyQ
SbgshdplfLhwCrStk1ZsALWL4HXY0DtTV2kH4UT9Ayg43J8jSoUT41ajIVg18EA4kEH7Ed599eK3
oCbAhj4v1j50NVsvWan9F0j5oNCE0T2yC6y93JkqMoOV6Ngs5FV7DjqL+9uzmpBGFvHAdI2QQNvk
RCWnP+1AKz96zbTYIkA+qUKuPxWSULpYM8iXJuOpkiHEAR7y6IXjIdMv8xWmCUcg6vdvA3RkjhS3
KbmN42ZIbT13bqybxBbWez2E2LgY2EoR8czF8IU4JgJXX1KgwsKZxygf/owW4ARL6AWKuxZzUWoA
SnetlIKlAwgs9b4+yrfD65vscaSHNSyy0n3LDp6q+9ibyVP+n6wYGDTn3i344CX5+OveynijIBiJ
pDiPhR+VbR+8Bf7eikBFubHvzzXIXGAxuc700YI7Z30yLADrtEthCjXuSOGJMcmQRrJdQeLDFxg2
+jeu5wXH/wW+oJCCd2eSxrYRte/Jw2HhhhRa87D7EvdlxbMFewp2rRpQmzqv482dCocQ2fLeSXeE
BSm0IWvv0tdJcJTwx5ciSc5gqRsjpa1KZJPmqKAji0ESOnkiAw6rRHD+k2cmgGEqBORwTlIvTgO6
BpDl8+nAIG9Z2ENjRqtwLKE8Y14sUCAgrbVRnp+g7SrWSYlg6pPXUdujfc0JUasLDJFrTBBeS0AJ
PxqSpRjffv0Kwg2xQHEmvtFtnVf+VYaf1im9bBcj2eFAraT1D66tp0xDswYOuDH1SyMX2zVyMeMP
Yz/W/UPvJtQiqdZBoKbQG/9cjGMSOseytSlML0xiImHtMZhV0eZTvhi3IFpzEbDtZrHO4OOBh/tR
XtUeYtJnvF7raeE4Za1Bc8npVirUup9it3XgynxQnb/i910+FRktiZkU2sd7G05SiJ7YP+LM8lho
ZfSoMU3VBNCj4B8Fb72MgB0m4tKzLDNuJKCtyqQHerFvIyLjYjozONXs120iJdiwkRqWyqqNwxGX
GIFeFAA8+kBZfJKCWCQdYKqQqCTr+AlM6o1csWftXAF/zvlGbgXnsG0B2I+N/HDHacAC2LLbbpKh
/3ZLJHxOKqbC1QEs2+fFOi+LSQ85n7HHaHo4u91bMFA3De1jCErJ9qP2jjaHHW4eYmsx1amtXEki
OAxeJ/YUQXOqE5RlnJTzk1E3Qvpnp4J97TSAjhBtxRB9DO2QjSfKDZgib3maatBSLryQjLbD6dHR
niE5f5dAZgfByHTOQjjqdQR8l1/L+Ur4977zR1cIsvyv9I2TvHKXedWcHf0rXiVKh+49EMBzY1hV
6l+P+HmMQ5YQwnZ+qfHMDwIXhS6PtLHIj/lOoaNygjPgvQN2UUMw+cS59lqoLxnBhSrTmZYMbat8
KSN2ZYTghL/p7uFuiA0CHKt4Gp1d+x/iL5vmtqDObc6GKGepu3rdW6dKK3gZKXyUycJaek9hbFBF
dhxJHj30it+jeaVJQjD3SzhimU97iavKk3A3FY82DIMrE/KGN+j2B+eQHrdjpIcI/BOnGmvj1ldL
yIE2pl8ecmRL4BA39nQTzLSl6RWq7oyGUKdkpfZRg8FQCBn3SrqoOKswqLR8JF1Wi1aYhLHNrBNo
Tovrh3pjhM1+in7kyrMpylFVUv484i4B5yt7Kwkj2KUtD83byq8+OlkHj1fjz+8FRMbYBd+4mTUA
HsfJPSOSNwUZR1MVdl7yHAwX6N9h7TnxKesnLrQzzKj9mMShU7KGVZq0LYz0KJc1VmyTRe93QPvp
PY917aHBhnlnb24vUUM+DxCkonV1G0QQhvq7xWx9RN1A07sCAuosL4ZYoYM3V/GDJN47wVAOCCrk
xo+6erEs/Lmqehmr9TWS6b8m2apWbcOcDzYKw2GYw1ijc4bUK04H1WeWy+M1RjeEAP8/UKDVZAdI
2OayZMyAJLnRwqSpgVH6gP4P4dQsyN8OidHP4Vkb+jPhy16SSwU2+bID3gChuy4QAJVUy1I9bSxv
VHiQYERCnrXRTWqxXeLmvzYR3SbA/Scu2J9w1xk4/CLSAIGZ6aCA4eZXEi+og6rQyWh7gRoP1m7+
83UClBRiJWOglbJ6ROh9X5Nysqhl2PDStEshjScL8DvxLveCSeXibOHsfsaGoDotpmg2BZF0vrQG
WAFt7wWYGW2RdlgrEKu3sELQgKqflsT0lUrhbBVo85iW382btFHFh3azW352T/uMO0ZikvAXPk5N
4K4D5zTIHd+bP+GZK0nfvQJ6zgJCZmMNVT4X1uym+34n617zrXy93yVsspWl1bPRLsUA3Lk+ePzT
Z7YRJ3j0lvWGr5sKdbSNCN2KIYmF0ff28yBpaI5Qe/sZz4c4PVVQbFRasnutHh5ITbAEySWhI1k6
GPIQrUM1QKneZA8FqX0aJznMy0UJUoAiqKxoSqAOEgC4cegxTyAf4naQVcpw3gYMcBS7AxsjOwIv
lfJW5YHWCkIsD6De6gKJB9yHBSp70Oux3SBQCCx2IujbgVELQVpLjLpgA69CufNoOC1BHel1nubI
vNgTKcfjOhHkbELVshZv2zPoEeq68grMXOrK83Kaj+FCMVQmTcKtmE+7VImviutme/g2u8wtJN2X
BUTJqKPPmVImibxpTlkEYj8ddcJDzTsPm9RofqT0u2aHu0/ZokDAYpTQSo5goP/z33AKEbSeDeNd
gIhfvJk3oXpH6FHxh6LiIFmSL67Z/qs+jzpKAGdT06FqL2ZOh1q/UobShIf/WrkLmd/u/5VJJ0S6
Oe87/kMZPzvB/G2CdIg9I2vXy1QrIHZR+M/MA00XAXuI1pG37D8szjgHGRTcOB9D3rWshezFLiwY
fb8EVatJo+dcmR8crOBTswaBBvdQMSJoHLq8bAEGCcR3JQekqcsiOnR+g60jdgTcWpyhCUirsMD+
zvG1oGe4iySQk/iqLq/GWiOBi3/a6WDX2ObDwJuxkkPIlvZciVqQmhSaANPkfaKkTq2H7YbFTfch
k3I+h5DhZ9zIOW/3Q+ndJmgVRS/Xvy96rmTIcBYg1ghEdlGA9t7Ha2BybvVntKpxrBbvI/wExIiD
7VUNOJqdUibyPeeRouAhFreRGsYyYn27rsSU8qMnVTKiHv/HEKayfJt5nxScghny//bls7djpvml
709rJJ56WAaT4i3cZIkLTxoTl2QY2i40Lwdj8nQN3hPvIz+s9cR/lCCoxD1MxmSaMbzyQ8pCUz7I
leZgisN9c1YGq2k/NpJZFVfncE6CqXubwA79hmgQJAvc+vCnuBrppfg9a3UQZK0U/obP52m0EX5w
Dg/Iy0t2QOXLOUPIearJhB42RKTVXeTaKa/ITBqe3Kgr7GZqhprZR9CEicQgTyaEkxEzkgk/WUbP
wxBDaH9suKCJd9dS3l+TQekDbj4pocEC6FyVXbZZ8PDV1n2vpD4yaaoiyaITmyY1ow/BJ71w4kxf
dvjss/mpZAiPyiPybF0SaM8z1IH0MPDzoW5HOeRC8fEzfqbeKfS2PzWLBNwG56xqxigZ1MV3ueCq
xGZ9GlRy+1jetmw6IYnoEsbQ2plT7oWX+ovIZmBFPof5Rb9XVhIyfL4kfsytI0/3rnu2VHEN0Y+4
/9rXGr5qvb+OIkMfXhQsvApFGjb6uPeUdoGEEoIvJA6RwcgJmY3XO54Bpz744BIWuuZUBQ2GQDhd
qpkV4/qNDItPrEZQOUl4Qw2RfvL8Qw0FKO55JXBH2GNHbY8sbkbuqFa6dI/e8j2kiVP1tauVhXh4
20To/A7vKfQJSow3yzrsY4OsJgrAmov1z9sLh9LpWr3fp8np+GCha/BaGdOayL+N3QlgiEsbTgu3
Rx8zYo5DUVjaB7hVgAiR/dUgvhcHvnBYyUdac6xKxuR2qh48GPY5VphZ+CbhWX9Pg5TERkkPAqgf
bJhqlAAWXoiZ/xuBns+0K3aXhRe718HQkL5mMFBP0m8dRAGf6F0OmBR6C7t4o2s+6TLWsAGlWl9E
0Ll9RccuQFLOZ9L1FOHSS+YEX6R/KurvEXyzSqS/M8pr4MHcKMRgkNeQNhP9w59+mRbJzKxpb6p1
jZSo3QK97moViubnOZYoMYRSR5Za5R690IwlHFraCCeFBvTuGoEHn4rpACMKa+tZCHP9zVE6Eh/p
0i09Anv80Bcg/rry1vxi6XWjxk14ymSuZ+d9cqpRSKsoE0BKyCimZ1JNwG2mVzZ9D43xKVB5TJtD
Bu42HCWlbFzF8nJxBiQjSeDSIAItz1AYi5KzeTn6CcC9r9yXEAz/aBwioCDSvczqCuKDsNYJoYM+
phvgDQdofvg/h5UZDxYOSHxfRyTCV1sRnlspCBWLzwgyC0FbAZHOGyExrKwa1/tGNxIFQdMntB87
bk9Pcus06ZVfn87ZpgC0Yrf4l+7xDvlkPyXl6TIaZTZqDzafGS9bN/z601OyluuiW1DCHfh6Zz4b
LT/kpUT3ti0Re6E9PVo+15BUhrByegnQPY/C/oa3/Vnc7wwJm33+DQNDXT/b9HSm5TArQh1vHmkU
EXl/LSD+WvjeuvHNa1pj2pZTxqm3NaAqODLcK3z96iUCiuLr6MJNeNC8FaGDzen6hathaiKbAf87
zkvfb5G0lg7MEAPD1ZEtE92Iew6Z6ebWa68g61uruvdZ0d/wUM4/tdPW8VmIj5MWdoDeukZsLWw8
kw/bwH/DCEz4oRUpxeK6z+xhP+G5gixWG25UaPQsw/QEPmET7zLVgm5VhXmaL/qWagYYiR4y872D
s532NXWtevn6+qvftrgqwtJmjKcuhbUg1e9yi4q9sjMoE3kciQkKcrny1R9rVAktNYqH7hs9APq9
pPQWu8+tb5S/uTKAo2i6ZEPLr3KqfNBZy4SczmuXdD2DLId1m1GNWZ772EFGakCnhTxakloARYnW
Xxdpw1BupiOfDzvX80vrvmEkU1puhGPCc+VUf+VYlwd/cp+LtHOvVSqL0dPl1xny8RlSC1vCKpIP
pVhru5+OrhXLsgfa3bk9fUiDd9Ng5ZAA4Oa4bKVJOMxpC7Wv54RBSwfJ7EHe9Zb8zpV78DLffGYs
Ug+Ex2eLsyZmPEiUBh8qZeFGx8Y3XIU4pYerWBydOWQmB3ryfiDqH6nBpd+8/t1BcgbMUqaBOAUF
JrloUSuLBtDVoW3Gq9o5tHA+nifjDsfOBYa2GPplQ1bg8ztPUvHi9KJPy9tJhaMRmF9bnTGyXCVT
mWkjxasHfQOrjlXjrUwCsIZjb74O0Te0tQvFiXWR9vsM/NYoEobyEl+prJh9mCjOoIHiBdBbYfra
LlqnfqaTxqQS8yjTbVR8/XR6UdDoZrTUhU5+06PGXhR++a3IdmxJqoEgn6vP3jSBHt6omOxcyMUD
sVfL2QzUovfuAHPndz1e0oaO6McMXVnWrX9L3ul8E9w7itStxz07sSxnOCGRjiCEykJ8SOKcGI67
PGt4dvy5VlWMfy3DW6BiI53Yh5nw7slWiNrT8tpOH8GSCdpehIcdOF8SijqUqSvTwbF/YwCmRzo7
J7t6mxokVmTBfmT1/NnXl7YEC02q9AB298x/dncU4jRFQOARmW1GCkTrrM+TDEsRTiqBI71b4W7p
r2V0Je793O1Z/djIaQTiv7hqruKI3PtSFa7hGs8wI3BEg+nfpW6hExG9pH+8/ue2Ety5NxN9i0v1
bya7t7tuBDFNhY+DaKNHGwqboQsT2MpPpbfZMgYwpV96exVGGYj3uJEgrpraLh7ZfxCEnX3Ybrgd
KcilGJbwCoWuhWjxJ0He++cBRnCt8ChLcSehbLesbVnY28XdKS8p2pkH2nLl40keNTxObVtzPUBT
5iW4XF4Ad5D2z7WLMNyAh6JmL1FS4zttPgfFFI5OuBMY8KPkvzMNpfgvZQuay34S559HQyWcDHwX
eiMFWSa826Kdt9WR28BXdDrgnUXLrM8HMsbyCE5ipZO2bZbpiueZzYf8FNieXrXlwA+PhiDzw69W
uF0K9rLZDQKzFQZctOeqrOG2sUnAlY2xX3vDe4ATqRheoSAuN/nekAm9MelgbBz0JswrLZIzbjb4
PdFbaFEVrX9RomujhI6x7lKjm8ruYDsXI35Jvrqq5Ea69fhXiQ4Sfn2/FgVvHSJ1wM1WSLk5R2xy
FS16IThN/rjYl1oQJyobYUuPy+DtWxY7GgFixVHcz/XYmJdXC/mW6ON/xxNoTI1TNJGt8aFaGj/6
C7hUX+45JRRZOA6x5A7Hq4byKDIn24lEq5CQ/0EKKO+gVwUDZp/ZJhZ+xBWif9n6lH/1yS/TM8Vi
qs1AckFtPNuBeAzhTvparZiePT11jv1TGQC+DhHCKXRA+i2DYg+Jrzwln1jQETk3UVQ0infafr+F
+K4ys1Xz3ZQLyl4a/YOGuOpCRd4GCu40u2n5FJLgFwQY3VhS0MDNP04iLBTWFJa13SEUg35z9KPs
Y8p1aZgsXgT0O0Mmr8utr8GxO/sKs8EZoLFyqc0RKG55sjTLcxTigv2kmSPnAxC09ACXqsPC8jb3
LGOfp8EfqPZZ+q+9ftHWCR6E8R8dXuUg/kmqI/Npq8QKfnfIFUTgQWFQc6eD+p+4Ay5tG1jjJpsT
HWsxf//YefdbHYm2l6lXzhS3ULQXgNcPYEP7YEdbdWMsVRqqfQ58urv0qtq2pmyDiT3WtaYVjoui
uM4JJab4pcqM0v/gluyOtN0eHmi6eZn1jULpBRC/zscd3JeFs/VqzOqK4zViO0MbGlAtuXoa2fdd
3hWeydFNHr3Jd0k9pNt/mkweAcLvzl9GrUuCTFSF/lwX+a/ozL63H+PUBypRDNih7poW1+1mPdC3
TmCvzXuTuCMWQDOdls+oeCAyLqoTf9ShL7yA50GsNJ6PznNqKSBaldoZHD2KfLZC7Za05qLyc5J/
5hwN6fDXAQpKaYQVX9P7vtYxmF9P/0GmYMRe4d9BDDSpgFvsNLnVPqSleSNyPmCOVPGb7ZjkkRMK
ZE+JhXru0Nwg1ZTYJgn0hhwzHaXmY4yDmEwBT/j0oTYGfWaY+yNWmVVKrvKN1Ck9/xa+vRg2D2BC
hxJoW8iqKR6zAqceilwIarleJnFkZdRZ2GawroBJnVi6ndedxRMUcQ+Lbby7xkRSLVHEJOFJeAF3
rNIx1UWwlGgLIjhKIoR8uFv3Scf4sNjMjm/VdV3V7rtYAn5vNOqs0q221Jdr16KMwaDiYNpUj02c
7KpAE/TDtMNKA5DqfeZ9gTLA9G0COUK3WQvLr9CYi2lBlacuQVam33KcKJKOT0dXgQxeAjh4IFAf
1JjihCqjAxvOru2IY2OzoTdDOmZuJA4kp/c2yLceJPED55PBbNwGrBF9N3bqqzJtclfK4uA1o2rj
viXHwDefNoGsJv/EnENr+Vx4T/DcWRx7eSChmjPBIy5344cLB7lPdi9TtDNN8JQblFQjNmlrvklA
giLjY0yii0JervcyEb7gRtmR2B5axHiT3jgn30tgwwIUZbqVYXge+RmLVU57pSy0OYG1Vvs8Uzvr
Q3mfFpAyQ3dqNKbsKtSyYEIjIgP9m6UwtbA2+TLYN3afoKblf4gKQ1BusWfoIAvMTPzFWquEQAGs
askmERyeN2pnvJu2CBZJ5y4wb6cVebRHLd72YD77BwOGGXvsptwV56oGSRR6lx0cfKi23d5dF4/y
3sRHLB/4hf4tF1J6vRj5PmOYZ2Pcklqdi90JBTTXB+CNf3amWCT2rr0aBV2fuCClI2BT70yuCDx0
yCJSlbhjSoow2ITQ9YgNbvivzgpFMweE97cpYoo1Ysx7mkpPGI4SvZMBOSPZXBq61z6e/NcE3S08
7eAFjNSuF8m9u1s8GPIS9CJpIH1/mFboI4BzqVMiKJ2nZiXTqOr40lnJbK51Ju9wvgFnDylCB191
9jIBZHpMBJT8K0awt1+oES6PUSeSXGkxncWD877KYAl8pPFK7gzC/d5rJQRrhx71CUbrYvrDiv94
BhUojjC/5KqQDG1MjPGGmo9eYLMuPYvuTMxWc2mWCrSDVedOxD0qYMX8z4yXaXw4A2GJQncjb5w/
HgBfSxTZNj+rMei3T12ti1DZCYDnIHkZNCMK/UEvLtcTvi4rDrVkYvJDQA5XfWRyOapUekvEslxf
TLcDfnOixSs5OLqNIsnnvJpfdBSOPjh6CfbW91ziFobyT6UKUkgQvIQDK0ik+BHEpCXL9JUe6mo3
6bA6s4gWc5PRQRN2hk69r7FLckw8t4W/KkM3IdzcZFDkVw2fIUgnTExQCy6QYQh0OLpeIE23Bohv
Ti7nn7n/PUfyL9y6JS128Y/vvdxxk2Fu/IpUSnCQRlaySvmamrHsTqKZfLcC7VxIze7x3GHUSr2J
3+3UvT1n4okYK6ZxpBgmljI2iQGupufhqtppqRNG5O1v0dhuyMOMHVUQepkq990qA8kb+DyTZxQu
M8d32cD7AxmpbVZBz/2/Pz08y/ww1bR5nwCapKTwfsZAmHRxYQnCxxEyP5V1xqPKsQKbUF+SXo6J
lMiC20sPAqBxZtKLfs00sYqbQA+kEWEGiZh8Xo0Kgs52pSEQncmeCse+pempaPfq6HU/GRJ3ekHd
D5YhZDHmHDwNZlaxyHPaPMhObvJ+yriK8F4IUw5WpQkIaWzPzgQ+7+DlLeBVgQVV/sml4MKJuYVy
vtPthq09BDyusqEuqzoCb8kEPF5xMvABRvWDZRfwCvcg9YFsyHbOgdO2VoTrQwaQU9J2tPXiN4P1
1L5D0kW++pbADj/a21K95vYiWlkTW0Aq9TWiOUJamJqXodEYPDPRSnTMUU7wkQw4D2POQjeUQVcD
mI32tRCwJM0+Bf8ZkvCCnkftsO6ZMFuuicYATFODSNSx6/C5x+fkc8FRZq19U+W0S11QcvHMkmq1
VOL6KJDNH8eYx50u+rnFxQWDwVtXRH/I0wgtV9eHHv8bABkyht2uwRE6X6QqDt4QI3b30oNpYraO
0APDGNNrF4ToOdkSawDBlNeZc7P0ck4D+bpVSqzNo7KJSZDxZrCYpIVl6LT1tk1x4xDtVfVpAPA3
UXnNiGSqQntNqr0AfPpB63Fa8/TiKqpffKYqK679tfw0fSMhx4KGjA63d19Mup/G8x+yx9gpw4Kd
kFbMj0/NKHpHNtc87lDVs2VQfC/vDY9TWFcMkFGbCPnWxIpiFs/d//6uMVdNxBl5kUH5R3E4yvsC
CmyZACVHx+bCHqdoawjX0eFanTkrDoxw173O5jlB8XE3J8THkwoeIyW6fttrdagf69B4PCFADMYi
IS06K8UXSNFRnQQ1uN1OH3rHPGMHVzNrkaKBo2vSl/QsxBaa9sIYmVG78k/RJk9qSZ/RViG2ILRQ
Jz1obhyM4te7tDQmxVCqB+ysmZEaPHQV7eeXiXvQL4f2qRxIB+12MvAZqRWnxiQ2g55xNvMo56bu
XhwSNYrsuk+p0yiD2pJd2R2Lu606Nexa1W3q/XWepTLEO0ZSAqBTmETSYkzK4cxyqtvZXACkNcmt
BfNM5FnG2fzJWzBSe2TcEAXdJcRFFQrK+rs9By+HTGmzPE1pgyyGzy+LhsIV/Pq/eiEdNVKOuCbB
KtvH1dZzZaUTsTerh2WtwC/MR0vOj1I0GjQs05hJsENKuMEcSNS5hV4IDVibvbrU/w+drrALowbm
K7DDA1wU1EGVYH5UMmEWDA2fNTEfkLlmZevEoRzo14A5EMqPDxLrHJCWODPGTooHHxmDLPpuDIMT
SZD1SYsa0FRUqwexPSed0BGUuiARLTRKMdJCj+tjALzx8gsme38SpXs8g2Cj9gCr7wKAEeoUmALa
jjXFN+9IpsxlM8cj5YPjLrHlAX64W0+rYBbYa60BLaSNu6OpDYHd8ESsJZsWRygDw6jFHcOeqNJo
PqYSTaHZRvg+9HIiaGhy4vd7kDrQCA3CBA2VLCR5jeKoEXxB1WaOOtoFv1QxtzkI57znNdt2CR2o
V13CL2ykQGJKFxcoAuYIwEJhb/gYRGlRm1Pm50w7HWIwremMbZ9XCQDmhOWlZIjqneQHIpRTx7yA
4vSWQwtd7d+Cnxp8eSL7TDblWL1vA1PpmJqG3UO0FsWMeyhWJEyad6xtvTYHk12xKZASEXBELy/X
LW/V19wz8wRCkTc3DUk3xkMkevGbg6jHyH7LP4w/za6pTu8okkKmBa1fABtXCxi/ZmevyDwHyptI
iZ8jMEuCQbXljUVD7sZfrB452/MFHgs/80kMkA5L1pjs0WTtSgvx+g78Z7q1ytbWGtNvxVpxNCUl
pX2P+lqmpUxoVUOzOLC0Hjanx5W68CaBSGqF4IkN6vK2jKckdFQz83THZgMvGGBtnRTz5rLjIt3e
Zh95Zi2iooe3dk2+Sp6CPt+mVgzzwm8EuHuxmItQobfEMHLNSw47cLY/09kLxvmZkCMoFnoCjt6v
yHDoz0vvICGGJwGgYlJob3VYoyfQ8LhGuCRM542KmWpU3i5lCwRoRSyayPj1qh9iNdvkFroxgmUG
AB3V5Q43EHjG7zSyvZZMu8RezSE0zfHFwA0pKqFYaf0qIiUsSYzufe5Wnrkx5M9hAJAsoGszZaCW
7TFGI4pE97MasbQgimQdi5xe/ELYJxWvk1D75d6H2A7xfZCsiKaj5Ei8OuhqFXluxu4jE7iAkh0s
RUHDVy6ey7T8jnKG2nuEZzhMh8sL5eYCoYtPcxeAxdcgK49X5TWO3j5Y/BtcuQJl8xdyQOMHYMEC
rNkVX3Gu5vsI3s550VhC4UMS5+Oe6E7nOB9GIN+rwG0kD479YjXKUpCRHvVY8b/vsC7M62u/lVz5
WmUGU6juazbR3Uo606+NpK6H+QBlms2ihMSGelr2CC2TllneWjRHJmanC5L4tFSlLhnB/y5H5jiC
r6JD0rYV7gnNBYE9AEk8RRdy2c2tqptgHxqIMn+Lgdln97t4LGV5V7H9FSqkmro4FpgZSY9D3jsu
6OL18PNa5YndPNf2/ff7t+1+fa8LyjnqifwqhoZMxxyBTwYUldpKJWovQEdGd1gj5Vl07AttPxO3
zy3PrkLPjVTlcWUkBdIhIKtcucv/4cFhFpYK+5GrUXfYxalAg6o1wceaeFv2PVeFJLEG54f/f5KQ
mmDNDdbyJmxFT6ioBkx4QR3PakC0tNhpxLyxfm0aFQ1Dl6Nk5zkAXQW0tSCO2u3mycrgNcmdmSN2
svGO7ihOyc8uBGLMRr8pvFMqOEdY7oGA0/bw9aJKSbWPWTac74tdMl3M8JDLitfeRTy1YmURgg8p
WOYTkF/qPu9wgGHC3Kl+diG9aEemcPc+4Ew5BSbVOf6enmM2SQv+7L3i/6wvdtf2QeBrGksIXdPk
DM6w2iPzlzGVQkweLLWfW+n3yDUHPxDLw3XwqIyAtBnPubg4WG7Wc2J/0HmHHE7b5JFhibjdk2lq
KaS+k07ITALzffPNoS15EKU4GT6kIBZEsLhFjrEikjpURosCWKBk/TYFQuY9QuTJGmpUiZ8iGnqG
1wqYc5cMzwOsyZ+oXrCybGceCzy/LeBZUzHZrX3ByqCz7qlNb9goiu/RMo+zl/t+u4dvNGnN1s2W
d00I3/hXs+GlkOFPSLb9dnFl0D4fr/LYYVPbtdmMPBjmP06UQk1rtEeJ9/JF/Fu/OYWo5jKRLzLo
0vBGK+hft8UBx0GHFlOnT9Oa4pfVoi0pkzNZtIP+ar/BEAgrnS5A6FJJDrVRINKhUYmZLDHGn3PY
Y8zelnn57KJ0/BEELst37v6XeYAehMRZCVL/oHKroB7PTx4K4ZS3qqPq3X+H8uxSP8KXaqmD558b
VmP4787ONqoca1CHUrU6UQBBe5R6HOVW5jok15nlIzhMb2paBo2fmb31pKIMWTueMAb/12cWFh+w
LzJz1MtR9nav+EvcsF1Iu6HEnnNkuBzQV8fedlY8BHwQxIwPowwNF/lE+3GESyODVofP8Pwy7P/o
OFBPyRQ9+1jKNhxXIwk5OMnv6mglQi1XSLcTblWkbTEUO7ygvEZLZ/4NOrx3Z1OD2fdz9WfwgiS9
7z4zVsr/f3BuYSUHp8z9AQMPjq+Gg2LVE87bER68TzrpRnVL/JYZZJ6YRv/VO9bQinlOCjtcKNJg
gHlhLTeFQBmViYVXMuDOzniOpjx3cNPH/UwJgi0YgnXU1PLnwq+ECDroJxljWnJEaVnLseyrPf7y
3cUOfTaibGu453gjtZNzT13NbrwdOYthUYECOdtBE4kkWtQFyeqztsPMKPlEET2Y5H0QqGj7V51S
Ck3y25Uv1y4Mldrka2Qel0T5gLUqCy5loGRf47xSaWAFQysJFjFakn8FTHMHZS9+bqPkKp5lEuRr
rXu9XK/attMqJ+y5lUaPrRNn+PrrBmYbtwWqxmu9y4xeYwlpuCywOwsSWvelbJki6mIhbLaSBqyc
5diSg9ggxDYG7kq7xsjDqOxsfbgH9BhJ7XpIRPy/eKbR1XsO63+8Irc2Uzksh/WJ9z9EZzerSoxv
/oX7uD8XdMBtKKNpBISENPNvptTTC6HpGcL+LZRLU3kko/A4UH7wP7WVTxNq51ifWKs07I6++8xA
0vdiwdeQuTZfM0Mzx3y8vg6aDJ78Ay0idFS1QplUKP6P41mbBRd4B1vyDbQldastFV4QxnQf3Mup
wg4ed6ntKQN3NRzvdJuJ6sbMDMo6kPgIJ9gi55E978rJEmsZpD4CWzDOablcmNMA5NJB/2zvl0Yo
Dxo26qaSctX+YdQhj+muEzUxEoBEZG1gZa5Kg8a8t56+L7oO07G3D6zckXpfuuRfw8HRvnD4D5Pf
fF9E6QarCaF5hGhZRukkZ5pOZc8HBjQ0iaqyULK2vleivDLYKcE/jL2GBsisTmAL4jNyIpHMZEXJ
6bSb7hwxrpBT7pl9Tu89k9c5DwUNZwlFln5AgiWod2GgtVK2CTw+XA0bL6JFUreVY2FtcrqvjQKt
OLCEpQqGFe6iX4WzsV5YkCflg8qFEbCZwe91Sov9O2vhPUeVvY/4tPQhVsMMgi1tMUHSn/ChILo3
iN4n4x8JxKG1ff/J56hrc+GQp8D3kgaRwxugBEQneCLwx/b+RY9NacTvZhqPR+kVg9tHZAK+ucMX
XI3vzN9SmNZir7eajLFOCMB23q0rz2tSwrtOfJXJ+VTiRQ0UdSEyoz3ZRa+UVPZ+IMKI41hIcMJi
qhb2NKlfPmE/wyhoukSrdDhY4urllF1szF8vRZJFQRQm1wuy5sxBuKTJQs4FOrLpyCkgmd5qJxFA
FkrCUjsS72NoZvo9ILBlRtjVH9yuA27ORUUdDMwOLmQVgtPK/4ZulDawytqK3ekAN7/yVAM7qXFr
E9nIeSH1KFMbsVOJAtiDbXtd+gmt9mFhign2TBa2OtSPYEZZRayfZmvSdC7lwIOK3j0Erxxesqtx
rMlGbEeivjHgqEpBSOKKQAIea0TJtazMLlzK9DBfRlDwSxufPjU57A+ZqDW/nOCklemP7GFVKXNM
xyiDwOFA9wYdxRRek97krFYCqITzriQgAxcGb19iC/suPg8JWxcMJ3t6ymioznE2fypU54Tws80U
TwdU9aOKClNebtV3ohZ7pbqXExvdV0OQhcQODrq1++uChd4Lwu/40hjpRM/lWGUhKkdzazg0VIoe
OUKhakOpZzq9hu2Y9FboM2MjaqQD2B3XEkntON91QjEqouXvMhmOE/3gBTriP262N39d4P43ns5B
RfzdjOM2azq7UdJQNJtEeC+3Zi35jec+li0ihhg4oNfvyYD7omWHcnUcsaO1DeESEpHP3+UKkJXo
fZPPRBD7KP15I7J7+ZcvA9nj2upU4rjuFniXCS+maDp8FrqOyPS5erKxa0Fjne/XIBhlKWkCSfxG
JkTT0IkdEOVMtG9J8INdWRMgdzh7lPchZqWAPqZAxhPXveigbnj+a5IoUcufAMTspe+jYqySXGNk
OZgW4ziuDAaZ8xWsVoYRqKGACch/MzKD5qYqJRPQZs5s4taWBPHNljofP7N4QUOmztYD1EBpYtzx
4l+oFdml02asdvvJ6P0Hx1Pgmk2KCIiS7EZYqt3Mk7zBDcUURzopT0t8dgg3keqnztU+W70M8b8x
yO9IS0Mc/0+/TVVXAQPeizhvzhAC8sEQ7RxVQdn3Lx2wkBGGpigD7F7Ozsmq9c1OlvvO9SZNG2v2
2pLP0zIaxdQN7E7jiC005SVL+IkzTCXXubemvvjGfSvGfQZrGKCBKaSLhyYvxJmYflM0LJ1bTrwr
o9Z4tLglpCiwYSkN9FSxdY+nk02YDeDpbNpMkBxOXn11dbC4DdXcF6AwkMZ8m7wpqc8qV0qFlAJk
jxdjI2Dy/B6U8ZrGtOMjTnLPLSsJT3r9xpvDOlxbW8rd/eQfHrmgBNIBTbJUfYDxCd1XztvqKPPF
RjPfzYWgP4AwksiWditaw3fzPqkf3SkNGFRAeMsvlQc7LRFriV3qlW8HaZXjMKO7Lb4WvL+Plq1W
3ZWEXw3Aae7ek/PM5UnqrXkfC3D1AbLBTOq/MhaNla67eSM/abzj3Jde81HxIkKC/AzaH4eoWlrl
B+a2whsDMynnQQuucNksKBbftO+va8ccf41kMagUcEZYlAo+Rtf579vMk30lPS5uYme6p6apbFDq
vTeHoTwKDnP6heexHTmCyb5fDjMtVT5UTV1SYZAkDlIWhPMbNSDsGzGwJ4NkJUEXpdBxKjXv6w7T
6qvkfXktjlVVsezwLH/M71QJEhRnw3NrR09/+HkN9T3zz7g5V1xy0vUYsxeGENRr0/aFdcVkA7lo
qgQKtuSK+xbdyKVjV1bvqxJZrBciUZwLZmBqSaJ3xyEWdQrtb1b9FqcFoMCNxl/5ulAMw1hf6V1s
9N63a7H/ycfmi0zLBqngZN5zSkoMP4whXcsQASbBi5is1c9GMIBXnttOwuOoVxJjz+lYhQ3rP8nT
bunq+l4kG0664xLnVU+e7MPt9RGfdDaPco1vgPLyQj0oPfwn2sp508inA7eu0GuLc9+TeX1ODZzN
dvUFzsFtFsO0tMVbsBYgWU1SqtPFO82qjfQRPCPEKohxuCfbEPFiXC00Ewupw0zLtv12zOgw3LMS
18uRk2F7Vdjmt5R3pCyaIhZ6FCVA9BD5PH/d1sDx/IzzvXO63eBuGcqxqunrnm/ODmI8pfqbqjz1
1O7QRNTHTcv9uvkXKSTBHvSitmcxcuJWJic3bKW6ELSKb5IkNA/PB9Eu2wHmRBXxaamMNuZzl7S5
w2tQwIl6s/BsQjb9DyifoFHGl1IfErLxoqEEdwkfPZ1ZEysOLfRrk5H0C38MB49W1xmEKXqfbyVg
tyO3pVVBepWDeAkqnYPaBcSCUL6ks/iz7t5n5nlFHDluKF4Wf06hf9ZGfAbJhxsnQ05XvhD7fIrh
ACxhSVdxWVY7Ck47MuwptFZOT4xpagHJcGenblCvMRsMPYM0QMpN2ovr76qW9tju7Q2ORV3/uccb
N5E845AXdGY/H82cSJ86lfrimh8Co8/wWu7CAiVEe2TeZlhrEEL3kq9R+PGGJFNlGczaR90WT9aR
dqXmm2ONgB6t4Jh4kb2pl8CsOE5K5mZQfXXe/OR7WgRMiakmsW2uBEG5Dh66PjOPKnHaTjbfALLW
t0EObNm776siQLM9PjbAaUqOT4yUI9qp9sA/ijtAb43CpG5jNXLUXLN5Y9b3dFA6Q2z4fYH/Q7V4
880PWJqrHa4bbxz6UMdgwpv9P9WxogEXPddeRzxGS3bWsLQBmfeZ8uY1jaTzZLN5KBrAyxem7FPZ
zVhdLuOHd3/VctYz1AME6XCfEgh62IvyaA0Pr/FktJIWtQLxI+VgJHDxekqzcAU8TufP56Td4NZE
Nbgb9jNKqQDNOa4ND4fHVT3wJubFnMrNfSMEz2vju9EDCeMKZWtqCQot/7komSlrFHjYySSdsFk6
fXhCHvwzOEK5tiYK25O7aLQrmTHFMrzGEK+InQn9GdKtItvaL1Qp5ZpcP2pdu/EWOzx/COjk+Nkv
+Fe750JpD5TIy5hBVmk6JiQEPF515pHv+sPtv9eAQRwZQyH14J8f3NEWJMSOrhiWbhDqdF68iSWz
DzuZBSaf5Urf14OWUeyji3XQBFNDgVHhoGDzSFWaZ7+50xCHYs4wsj+96CpeNMZ6eqRvomoyJrgO
8yD7TLFsy69Ku5NkiJ2RSAfCgL5jBpNYTchLhPgV6ord144VqezJz5SPuYIa9RdShYyptjiMyW+I
X5aBWbTtn2NiGamelTbeLcPDulSEQ/z1RUM71VYyc5iN/Ag0/lSZe9cTMlUvOEgrudsbgJrZd4Cn
TWSX32XY58pAS15c/1oSkMdKCTs4ojKwLGNt6k//8EQemql7j2rYD6eq0tfqsT2CzBFL9kXoSoNx
4b+PspY5S3XA1eUkwC0nWslCOCMWH6C62PURmOsnpkw7VFaDNm72eptdYJZmLiK75eyBlfwkOmek
hf3lVsZN08LhQnK6V1k6yPvdQP2P1/x1JKD1EmQdST9G2ZRkbOx8S2kwiZgxziaK1m6S9Z4K6qHQ
2x2Vye3uzXupVLuxwstI9DDo8P/3foXXovTzWn70wQZFzK1OxgaL4qsSPcr0UcKuvv9upU+vhEA2
NrnqrMs/j2E/IJeXKg2hANY/u3uUT1wYc+svEMveiOPhNOM61ujK7pwdx3Y9mtextgWivT6otcp9
uqlX0ZFK80f6MNGffNtxFvwic+cFJSqKMLjA56v3WLJZye29UJncssTTEPA7Tb8ozXpXu0HaJPKJ
IY3EqBeBT/TY7ijfCQCOwu45F5W/zdDycJzdjW2/ugbB4j6ZrUkuNOHJh2CKOxgCerp7JwY6ozvS
1A+84LsaJTsqav+EPdOZ0JPSoFP5upiKhCrNAnwBD4A21KZVKUc0oIwtMyN++8VxUIxjitd0lAKj
769nnrISCmM5bG8PjXTHTNgvQUq75sqpASWKFON++F1Xocp5Z4Omk/b/bRyEU3euik+4yc8c0f1/
PKD7Cpe+xmClcD88aA1sgCTJ5SmeyxgyIvTyQHMKX87mZYywwkB4tiiJqi4Z1IhAQ6xHYcPeirMB
jf+nuJnb5WyGpk7Af9O88jsEeHj3GmDPLgoQQTJh+oGpJEdwhXQjSPj6/s8xk8xwYu4Js4ML/vbh
YHc8Z6V63GzwPZCyvD4so8Xn6qsbyh2m11OKBBUba4l+2ui6d0ZNPM/fV6iN+yq48AeG2Rw0gUDS
lVtmWOPdvOw6GzextaG/RM7lnE/9DC+Q271kFh/VHgKAkkZ6cHzZnL7HpxgmBmnSlQInODnD9YLF
bXnFISjLe/TX9OqxjQBSu+QLHeJxFNdVzWkoh/v1ledA8sKjiiBYCcof6FaiXyimbOkIIBKyyde7
GHVa9138TjkXHBYtktF9sds7LTausTQnropU3/R/EDzym3D4BH3jphxXwwNJSLXhssbjJi/nsuVc
imhpAcguBaw24xc9TqQjrEDAcXxk5VESIw+K9HELGApQjVOJCzpBh+uB0tqrbEoGztJ9wtIDaJfj
rz/0ceB3vMjuPdekh2S6zNXAdCu2pCjHaTKZKO351ipCqDaBJQTf11ffk+zmU0qoXW5o/yhy05qg
Vpe6079tl6/vwG5MPZjApyFOvjvlzo5oNs6eElFKh4eKx6GrCMOuy5yOROClSZGbDIxxCbK3dH5v
yZu43eU25Zd5rOsB13jFXGs3V//aXowfh2ZfMx10N+BMAh97MmSHF+vcUA99JW98OONXo02eErvV
EeAYrBjkNZz1Jw0/yAcSHibKLVPZNx6Xvqv01fP+1TiPGFe3Qr6WiGTR4nAKkNRktFEXcjOkqH/S
ETWdP+pzvhDkNWeXgIsuKK+z+NqbBNpXqDrQyTRHmdTJMJJRihggo1hYEklj00Sq4Ojve+xdiasJ
XetgOcKJUu9QqT/XeLEMsDmkriuGFcpCAwS886MkvZ/HiqpzdmtE7gFmcKX6EvI6S7m7eftLyKIV
RJbCrLsKf2u1rcK4/XJCM/INZInmjEjqz+JuoIT/cgpncLrb0o0hYa4jDMqiM3vSbMxwbLAr8IAA
Ig9H1AnJqcCTgtRjmkOwNyjf6puhbkY1+xQbnZCLC2Z3y+CGEJwr1dQt4xE699mad1yLAXeXv2Ho
rrDkKgA8yCWfD+fuo1a54YygN6dwEmUDHPQ4LWaVrUoGY0ghJFz+HX9dsT3i1+i7u+HKHQUN90KP
hBsxs+rpgPFDq03SEigr8VzJVTgXJtwTjkx0xQzhOKh+CVJW7uV0ZISLOaF60YZ5vTpVLlV/ufGh
paGVUpplSK2HTTYHh+t4GfkJosqy6vVVMQq0Jy+iDuV2q+0HnCO9f3bBYKT4WAoRwztpXeU93v6Z
W+QAV2kZWFWEps5cvJdxmiXdcHqniQhLb+qAnJU+VmRqnwb0CA4d4WIAp2IgxMYkJk96qjnbDK1l
amqTNJFLgKjXnfm7Kp5PYb9mmMCOG4MS6SjrvjSyVrIdO9P9FOQJDh/xrczRAj95ntusQI3gYlI2
jmFXT1qzinfs6hTQntYmLoWUw9ahJLutJ0HcWJPmej5gJ5txWVelLPNPoD8mMKqZw2352MGZHaQk
Yi1vW0dIEkTEd8E9IpQJZ1aS+6RajlOlL5Zck3pVEnaaIphEg8N6ZEu2aLb/HOZ1dp2h9TMFAwvs
4gAiHc6jBcDn0S2waaqGyMw2YRpfL3mWSP9IQbpwFrz0bqfuD6ETGS47aON0ddOKJBDxUGrHZd2I
L8tp9fZcywPBMa8WbM7AI/nGrKyiVlkbOFY8WOPejxujP2/2B8fb3mwzHq5OjshsguW+ipF8MmEs
iw8xojLukaQA2USynmnw4mmb6XBE5VFHCNT3Wt5tuiluS/KvhDOt0PzWtnf5Uv7hXLPtVwXoQYVv
kT4qIMs7dMBHvbRYE5wXn+u0VHN/5jIL02UjqCN10EgwxgO44vedZXTCktN1xMZYomRtsJmLb0Lg
rjnAYRJYRgHYICfn+hEDDDMJfyJl+MY83hIPMbNDc4XfTy8MdMo0axL9wCBQiwCnsMwOvfXQv1ld
dv1EKT1U9XqX86cVziYY66OkmXM0TaGTeOcsqTdkIxnjhwEkkO3gemOB9DiO5x02uy2tZU+IUVj4
eVoW9bvNAfMXOkBhKaps4Z0uf2dF0OfT0hpKkT6EIpERIYxqf0dX4rQ53tGrRbYSQAWXUUHJCeNB
4VjKTCJKiSw4P2i0XGfAxcfgEBdNr8+O3oTyrpO4MmVdgqkrcfRo5mcxYfhjb9h6OkamfEdkxScZ
AAfAYk5tmsRfAImf76F3uTQTFt4RcWYQCZllhKvUPFiG04e2Qb4WH7zB/fa2vyIvt5QW2CAx9n9O
Zc8JVEck5ugGXh70T0C0UlWBKPOR0Ys7srQoMUjugVWZ3prsmFL9JMB/5tEEnxK9jk+Kg/P4Z3jF
Pr1bej7PEBtglPT3ZtGd8RYs8EFDCOw5/sHTklef28Pls+HqdLCK4sNSsatSMaLrz3jwRefIAs0b
cwliDAWmFRXRlRK3U2PD3VV3pUnefITfzS0shX3oEDn/AUnSGQUiNF/uUdbdKLjLjmZXV8RWmY5m
QemhkBZuyjd6gTWihrKqT4hKUmChUL3JLd6GuB/uW0rcXwi0J2u/Eutn8IH1lta3eis31W9QwDqy
3iCOEiyZjzUxzZs2sPQcqpQ8ro54K2MV+NEt3LQYzD1PnSen1atfMjnNQ8qgggz+yuGomjpgXtPJ
XELrHhHbhAxP5baSWbY9R5fqs70qwsnbYSlFmlwDbN31JCpAGGu3hFqWNWH5M1vvFnoIStXQQ8AR
kkK21hDFmTedGKUl/evy+u5QQP4QhEZhLvKtg4A7plH+eiAxBMvwHQYooe92tpLf6lvlUclVA56/
/nwkJeyvoZ1pdjNw5B8CC/VC5KfdKDdKd0DWvVB6NrLz0CyZ37Pe2iQFdnpMdijWs29YQsDFMJkt
GR7H9Fu2PZcwtrI9Q5wM8XJRbFEDKKJi5CMcN+ax1G03KZ8s3HHUcFVMRXMI2mb1+WLAUdm2qTgA
QzJrVQ1cBEtgcDfRd0+JWCaX+G8Xu5ZI4/323K/wAz/9Ypys/RDVJZRYRuKIpN72Psf7BA/kMimV
Xe+b+cdzuXjPFNUVdXoRF1Laarm6GHyPPdI+XfaVOIzidLoB0MKP3k0I8JHpN4gvm1XjZ39Y6oJ6
Cm8JVA5e9hcQtEY24PvvCxoKu77xIJTnvSqLa1fuX3P1/wC8RIqdkQNnItCXEt+3hT2VRSQrICbD
9Jw3XeDY4+FrlFGGiY4I2c7bSJUMYWooFVsdlQChV7+USCFKNxJDxIYU5YU9DqIV2Vyv/HZHlY3L
mE3r038zdKhjW9SYJ8cAKp7I6Se+4fKNgR8z5iwrMHuZkQ//L9RJUrh9aGdIeBZRVPpN/tzWNfrd
qk3XxG9nIbcxZzkO3m0rqrR/eosu3nAfs11TrnDZ/Be01tF5S5QT26T2wQeEe5t3CiLHIZgFL26w
kWBbc5ObYN4I/H5gXBPx4bOx3bDc13SoLUdwS9PAGI3bEh9/JexBCen+aesy4v2Zk1iAfO3CfSBK
yBYLYsvaM00xrs+jantY/9yHDpg4Hf+KKUCW/aa/TXF6ImnpQM3zrhY45wu4cWwYuHV4XV/AoKMD
5yNus4+QUl15ghrnb/CFjczu2SZhiH94mOOyNm3GErQzwDw+RygikM8/MfDf3qHe4KQblD4Q92bD
s+lG4SPH3Xcenime56uXh9QtxeIdXCYSVyDi/hlsviA2Ic4LUZuMRoFSPVRGDBNfXtSB04D1BAuo
t7IAU8zQvAZ/lkvsYElqOSjwSHG/V4KDF0IHW1SwF6P+/fzwubB8yR6h6Cj3Lp9TYu3vl0MEKCvU
5gnmokWraBsr7PXlOSvORmOlxdBVG2QDf2HR08pAXy2520j6OiI1ybfy4EW7v3qPHmWxBt0uzErO
DFGniSxSd7FNAw9O5OxZTI+c1bfBQdfHEpEuYIEWzT8qWxkOx/WeqJfBxd0kVX+pCJYAEOxxWZRu
RefwzBK95E9rNcDHMUdZYkKYUYZkit+10mAuROZkV/KeiFL1AOymneVNu1FNOjaR1oY47qYYHsQY
zbylTA63Avb0tdGsuWEQIy4SNcWD2ebEGpTzTWhK/QqcT/Gvf5G3DdrHBrLxvk/KeJEbXnTMQSkS
7DNtM1NPZm+LWNIlXfQ6EDk9bBt8ABPzZqE9L6EiiDK/PQ8iwRdYQk56rlU6EkJqkqyVJrinG2Ic
YsytIg8AZc1RD7Vk1nrP/bH4VpVJ1YLMShPQ13edLxM9VNePQjSJE2dvY6kYqAi9+sDFj+/sCYul
UM9qVL3ooIUUFMNp7kis26g3uFACpjEZYCYyApdgEZkfXdk3YxeyyssisOwkA5s3LFAkiAjIiIfa
3/0b+4SAFqsRxiFy/HXqKn2+x2nP+gk4V15znNBBBq/iBsGgsjkXJ/wCdwyoDrSs9hT24bJbBWYt
6Q0/1bUimMvxcQ2inhtEJfmM8IaB2L5+ti+bWnHuZgK0xGR8T2oEqa6tqSP88AOfFQb558bKbh+3
5a9gDee7te62dGyAxYT2gOh3f9JIHBkzY93UlmgCW9KOLgqsUMDwINaO1tSDSMCliPE1f+AsCBZ+
ficqZ6v6RSvReWNyL5UGZx/NotOyCei0JDbRi7m4TD/1P7VUbCZ+rsTJokvM4g0PQ99DMyw9S0od
W1+jSTBbFutHs465yZdGws5AvBACBGq0BbfbHvgZMcqZRS7tP9j4g/UM0f4OsIpyNLFLPesn6LKs
mET+3DPUscxiHZn0V36E3+JSx9NkBjcxc1VfmxxH7QuliJaZurf/0SSGUrUmnTA2vFLosZNpX/Hl
+hlthR2ZawxFcXBCtlM6OXpOAUqTkKjqG18v+fTCoQHebD/ZD2/feU+2u+4RNrDfDLV1RZS03upJ
7T0LYW7D9r3wzXc6wDXXut6STkpC1pV+A6xq9f4fmqHCdwsN6DuBdLn8udmrUfsIYqNIXv91loQg
x/jxsEJY+5oHEc9R9YLWIQOu2huTzu1kf+FkEqZ9xvOgJYzwYk6t9zxR8dP1mI1BsxJPyXKWYyj2
cHLzKNFkyFgVMpyycEKGaY5oZwtsbn4x6B62HdCsccwzhQ5LUU+MxmN/QpbjATibH5mxzB3fnYa+
KEgvpLlVA6MgUKRet3+lv+S9asetb4/v0RG4k1TP69YEtjvpl2aDOs/AXwsj20r09z+QVtyQm8E8
XIqMoTrzKdmw5PlzIlsf74rvgpTV10JAdDUwdcT6JrLq8Rzvkb2YcpRgSUCKm8WuuRvDYM5rEHRV
hMvv72hLmagwVlBgL5qnGz10ix03JO8j9dGtUdUmmht0NxEstI1v3gLqBUn3elOUz2iF0kKrH3Fy
S5AocSyTlq+rkba2CtSJEiuJV4qp1MSpqdl7a5qBOzwDQnL72iv7lqS4SD7szcY/5t2JQ1gByw1e
NUPwR+E82B9qLKxzzGYXbByAwz0pqRraWYUanNG9PBtCulmd3l06zNSM//SR44JPOdMfE7L9Qw86
W1ug01klj0laDbH4Kt69fiy4/kOKo3PYUOnLBi981uOATJj2k/hN5TGog+L0VjYVkf/lKFcml02Q
eUc+YmCeHX3Fe4WVyptSfqypsLHzEGGs8e0SsCNeIacwSyz/sPb1gnNkddBcuREM4GkfNzdMu07o
52QCGbl3y93pquI3WFSOuiZBwl/V9FRYLRaMS3T1TYcZoI0QmId3ELvjQdt3kS7IIXRB0fOJT2wj
iW6pv4UMGPy99H6AryPXyvWUBZhnqDgE/zCyUqffM/F8pAdvscwUKeMJUNY3gaXW1CDNz75r5ijb
MGhVySLCC4yxc0n6jL3T0P0a/ZNJtpAUEncpcYvqXzRZyD0PfiW0terdqaIZHwWPvHN3FyNvsKgX
hrEX5NkOJ4gcG8ZXpFw1rhYsNTJXK6GAZaiC2UxzdI1erHBgYHhxbLKkexkyfzT2RPTvd7ADMLBW
x5IJwCZl5/WjtS9g2fyZbkRCT2JMCbyn4wUCrBrm3UWgUBx0hRVtdAV7SYX3cfl/kizsvbayft+z
k2rcAatBBka7IEeoaRW02Ka7q9cRVW9Yl7fMYa9sbixftEr4IgHogaSzbqNzT6YILzA1bBctcFqT
gpUAyLxfRuQ62QcftIzfFEum00lKBfxzC3Jei9LVG2YQ1H7e/nwwzzTpmpMm7kTdVpNAX2Ng6V0B
bmk7SJeFxU7hdeSMCla0D6zzOBHgcKpz+ObLt8LmK8uVxdhq4ypGJ8rbaTHSXhc33jYbtZv9oeZj
GqR6qVwdg0Mcwmzi7qaAVmw9pZpNjPgkhAqKUuDVqpEfv2zFcsSjJMnT3qAp9MyC9gRR99gWEmUE
e1WFr87ObfPaTgmDLwEYFs/xvhE17D/Dcs/LdQUZwPXByUtMevaHWze0Hg9usOddfVSo4/WrF9te
zk3Nz1HGzxqb2LVTOx0vwyxONJZatLa9WvhIdnP9Z5In/lFH1FXjPXHlIQDymQS6PfPnR7g5FkyU
/EOl9tCMZIbms8wt/eT0ZXjMv28whhMHPJgZqTDFXQ2wSq6SdkkFN90VWmq7YVmq0rxF/2C4jOrU
kQR/PlQU4MxClw/u0Cq9NlJTWNDv8ZbsBRhwH4eg7K9SJHgXk4NmS0a+5CTjrWq5ve71r4ejihpO
mqNvo33lYCplBBqFHpcHC0YXFzxLkzxpdP+uTTjkiuQa9aD/HBwyI7TX/ZFYqShC8VWE9F4kf5wZ
wGLEFoHSpnjlgueQ18jRI9RqdFtKnXqsHmDQ+qQh9ikMBFjwIpFtSsPemMytG5N7Tau05iDfcngB
W1WugrCywVmLOfbtrSGAZ7NWVBJmIiZ5wVpLJUVeNpsT9xEnLgRgdhiUgnDYvJLZtoNYCsYrkLIK
Te7IxWJda2KmsXOXS19flO967Xox8SSJa+o4jSIan3wPGvwMMC38MbIDmXqz9ljNdU597IUTTCuV
Yu9tmZ+QYwgPlYXfWFbvmFgjEkCvCwk0Y218WzTqt/Q+cAfdHco4FoKDbI/dzMad+zRuT8JhuHrZ
5bVDmFlrihMTr2iDA7G+TLFHEVm/z4VY88+6GdOh26gidqzK0ZbTlGHBmLrgBSwbPnVe86IUP8KB
XAXbqad/iP1wNmLq6fuoRZ6zMismg0ATA6r2ILR3GR+O23xwSRKoBWTQn/+EwARa8T5M8jDCMGXy
8kb3O5RZ/xQolDk2AsL/qePTO34Jj4HRy+7NIHOpRfPGTE5NAqVKNZZExjP6fUhotAaDD0b6J1bD
w+HMGfr8PkAndx7TXBomB4uKvRIKZ8fIa8P5f/bLDheefKvXv4WbhY6i7oudi+EfjRWnhJj94Cb5
mkLfQJPWT6omFKUFdF4yWhktG0WPYkNecws79TiNZgIWrcT3bddj5pNl8cVYfE+BLQUUs1Uopx05
wkhnksIu6nSPtaTbLabPByb/gdvvIUBLUXHrhHUXczbDD6rrib5nf29yAPQdQCGHEnr9QR+nTxr8
WwgeJx9PUaE/tZ0OoRn6qi1BZUxJ6YVentdgDgmD3ZLFVQWGHlSEYHdyJ96IHdHRf8Lp3YJM0Zl/
N18NzS10sCa93EhlVweBfhgmkwUr2J22dx4r3EDYa5Vztc4nOuNxHFCxuROd8QMN3ckdQ+4B7Ily
KO2MQ5PcCBYm2LLvt1cj6AzrvfgIKALU5eBMSwdTKqJ8sKYQTjzRAdogjMndkgUO2+t/0HCo/ywO
4G+Jnrdnv6jWMtkju5MceYSc4O4ROpxqVC0LqDgdDHW0klpyWuhPXuYsdNkLnz/sNFJiCccK0P87
3Wlhqe0qibqLefqeQ7eANPq/Hj8JfNuQ91Gy2rDn7auCo20YKCda88PuAr37PToarUWOnuyWU4Ag
xZROa41KUZ6LgP9ZBIGhVcwfJU4KYpECG1q3ILVlkuU5isqUP8B660uxlp7jGOUlDDOSLyFN9m3O
0i9pESrFSlHqTlOW31g79d/1ogz5ZehgdNhsfnk5mgeFK1W4tYiLEG15Y1wd9EJW/uUSSjEM44Km
+q0CuB3cGfGeXKXq6YPbcVf/8YzoTWwRALFEIUT24Xu3W0eEKKtLz/zk4pS+qkQ7pmefCJwI6Frq
XzjFTrEUHL75Gf2C8r+9eN1fDEP81s4n7AIAEvcjlXzzFClR0L/gUm7NX/ngzLsp9uFKtky4eWFv
YIlXDLY9PCaRaNiKxFVPow7OcvqmVdwy9zK1NSB25Bckr3P4AQX9Q/ZMDmN8ixlrZrp6Gk97CkK8
I3wiorCWK2tMKvcOjCyk0ftCkkylG/vRfL39QERPaZBIGuQMKFUrg3EIUQ6Kcck3cu93lVYZCCjs
OLC4MIO//KogRDCvHmckXchWUHGVg25cOzhq5Uh63gvgZ+odQ5et3Rv5N6o5iYvqTTo2JCw67AZO
Vd2EcflkmgkwqPLCdTKL3CbZfi01Gtac30e6FTlEzuvHM+hcYG3npGSSGRuUEVIqF4ENsDYAD/VG
/hDm1qneJwDtuUSAxYJPJ+Qr8klUEtBr/ABUeDL7U5KOumTumNWqhx8d5Mdt2r3rISKB6P82Xv4+
5hSWVHa5nDghqOApt2c9
`pragma protect end_protected
