`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40064)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT++8F4PPQq2cD1pLLMTjPTXpVh5mCVTmh7KwU2ZN0/MJz6GWO/3sSZzd9OCNRDnAPjQ3wg4
tI1NgRv0f47T5eD4V63LzEHwe/AKCwdjalw2LNsfIzZr61OcrkT9nR9ltb7UsGIf9tkbnkYoxOWn
WIeQ4J841QPBEaiGie+2hwjDwP13sAdkoipjCWQr8uPrSb5hm58qCukEfmVnm1HUxnUIy+waeONh
aPdsTDx84rBBk4v7nOy+ojKjkRD9q0O8WgaSIBKVLxYdo4goUSSyI/DzsVeDj2X+AiP634JG4YXU
caNSTnX5d0amtbLDEgZKJGoSQOC1ASzVtuPuB+22rXMK4yS4qGV4NKHkKN5fvcQsedFWK27AoEzk
E1wspNFBB981SfFhCIw8eB0YdkigROk5LjRXula73O1ART7kRMiBu+Vjvw8SIRctRsSwp1dgMBUK
Fl4q1N8Fyk5ziulIq7WTiEM2dO6JUkp5YYcts6nslSGyViuBkuSTMDlBY42RxSFEVBQkf+ggUKhp
uzg0jSdzncFVy77JQZHW1W7e2Dn7lL9ltz2RChEfKUl+bajAfrDFDqMplDMggFj9mL//fQPFa2ui
x+iuODh+VbA6cGQ2TQ93HBFruMdYiWx8Hf8I6Wm8MTXjvaa+/nGeeAI5jMJcToMWh3+G5rJIvgFF
315Ik/B6dqvIcvsq61HAbRi96t2blDHvr/uauyjrV7sZbrTBxX4i68J9PHmiQSHw8BU7Lj80f5Jq
UD0WxsS9qIp8bVCz0prJYUIvW+sxH7SMpdlPKzOcBuF9B70dNZbWieqxL+z+qcPEVdHLmK/kyPZ7
7ojNrkxNoTPNN9hV2JWV90p2UtGjXgEd4Px7oJ1b3u9nZjiOyIY6pSEE8IEso3f7/kiTFUKOuJG4
pnwRnsC4xRHeTYV18tqh6/IDws5tMYKL7H/TXCS9Oy8Tcf+5nnR8PBnWQX1tVQB8KzHGbRgrrQ9t
vd6W9ykijkrG/WC/rJt9AKFWnUSuGJLf78HCQEDig9QOavTcFbL7Jr1vtoMwyrZw7qr/hubSw4/Z
ocLpe5VTy3HYW6+WpymFZ2/Kp1TIPNoQtYHJTE2TbNKvn0zr38JVg3I+kEAgo1c8dtyf3yaGHTdc
h8aFDnSS3W6obL4cx73xrwV1tygequUrtF1J2Wm99NQTco+g2P/qfzkhYMx73p+vvSscYvZLP5Ne
PV9GhHV/aPZ62TJlAhFx7kWstW0ZDNOgimTiUDry4OA287KIvLQ4Ffv9WeSoGYZj+O8OeZUwVacw
1VadUey9EunxYVFxEM0CBQ2owxxRFvh5wDBakZDE/KbkTp87UAWSGB+WaH1oqFEsJ1O00EyJp6t/
0LHMsQl65vz5ccGXl2Vaqi4LtdW16UVw3BCB74Iml8aQiEBkzrQpPMxpPftPQQ4icijLNI44koRE
arYbDhs+GYoMB21rFM4U2HmzMIc+ZIsZPuyBgoURxmFTIo9kRKEURBXHQ9Fsx4jrh08WWNCtPaEN
hgnFF49lrMV5yD18uYHBuCpnzNm1Xrl69IFtvxEVCBb6fA8/utEh4aT863ddCLj7YHA8gyWrLV6U
5Nj0PnOyy89DHOCwSCQdpB6doVKJOmlc31g9TA7tQ0U5GOi6rtHv8qlkZEtmeSRi9/phKDR0iVnV
pb6WH5VNGJKFdccQMdw1JCW/RSvhsFIq07DYrCuht+dsIh1im3M2WjU7p4arCzA4o/eq+4TPRnb4
28XGM/6+d835A8F/VtRXv+PzUwWFP2iNCN/v9sTmUx5HywvumErpAHZ99ZEJ8jaEE9VJC3T7Jx4e
bukPKYPAAUgcl1Cy+onC7Y5LC+7+Wvf4rbfsdY+lDZeIUR0nQEWwtiGlSaclxOh+czgMYUnnQvMd
Egl797s3cCI7Q1uM2A0b5xHFD94xAEWo7FNddrdStVBf1qUo1kHH0rN9/InYXlaxLM/Mhb9EvCU5
tw0sDZjpeZwr4gF3cV28dvEEd5W9W4pHspYrtOm1PlvlF74gzLN8KGFMU0G8okRoN2O9n2EXxqlR
A2lPa0KaXWBjickrMrV5KqNxgmHB0nSLxm/sH4zmJdFbZ22CbP6C8c1DKGnmCt9ihtVI6EFNC6Gn
129XtMrJF7ML5i9r5ZTRAciwHr8nT9TgBDdt4PJNGBKQtBB8CEEHml6EoD7Dr72QTWgdO55PHFCQ
ybz1mRJp3+9jUgTMO4kGayrBnorESK8mI/WHzqVDK2mJ3Vf+uxuMV+i+NjXzURNQHh+LTEhQ7KhU
Hq+BTj50pCkSDQwDWDH0a8AGm/b/P9l4okhkPir+k0zFmE6rSlsByDZJGfT6AZEVHNWiOHw6XpvQ
oCcOcvJqdLd8zdbxWNJiKMPN0/kI6s7I6hV+2NKwPsKowFhzXsH8vqZ8ovOe738VOB4em6lnMTUJ
GJksf4mrn1dnp5xT4+nQPNcQVpzWuYDUEkHWY0jIh6Rv7bfGsA7pVHi1QOM5cN3QLVf0XB8HBj6/
XP2eu9fwg/dmNoASnATelFy7x+lmHAabQOfQqmuOUDuX43VZ2nTZgAhzMJnEI5PATaXPmk3wRyur
b6321d4eUUvQpdUhrH0SU8ZJDL5YlfZVnD8hBs48iLNn93PWQw7IID4rjx4ZtAU7q3JV5QNpDaPZ
JvR+wAu6xEXOSVJhtQpmyuoIdhfUwxM5qiVbdRAmUmby/OovLwoWpBSOEeU/E0PdQYY9T4D5LNZf
4zZJS8JhjGJzR7PjtLDjnfEM9dSaugVVfW+J3hp/3Z6x6JTBaa9pMb0e7nyEEWv/GOyolC64rozi
N9bh9dSgVF6OL7i0h50UCIGCFcOEtwj9qMlWzVmp8r72x22RKK76Z0zszYK4B2SUaLaWOmibWqLo
VSijC3PvenO6ngCAXZ9JX46YTRn2LNt23b6EAS1aXws553BY3wUly4IMZkl6kIEEsRpXOnSKfwb6
LfAneH1hvEkz0ACZ/5HA7m2mesJVLxX2p2a4q7N8DoAU5h0EQWxLyK7aLCD2OJNicKMiekiuhSGG
W/x0NAbA5CRjTwCPBjukyvgzG2/DprzrfaTDqsHihYp3ZS5RdXMRTYLD0hTcSMrc2b3H7Axn5zGF
2jI49oygzEoMacYpxE9uCoWc1TDv5V5VMygQh9WaGLbgIAoIAiTtfLQ0njQ283aXQIvfftYFO1c1
YfH/C04A4UAGq54mH/j9728a/4WAxXOc829crg++WdiR79Z7RSty3SsAlqAPvDdoEMnjA1ZgzDs7
OnpjA05MBjJYl7RKJleelcyla49P1mX49ZazfuZqM2OEU+nmplv8QOgfCuVj0sBW8G2qXKpQetoJ
VHBLcZn+5jOdF2CnSPd0ezCxo8knft3i3/6zPBtF72ZIpDu2vTV1ErF8ZUi4GtieLjLuMUKlZ45A
5uXMKZVlKUEqAt4Ox0hEGYZdUE3xkCZjU5yHQ61d3ip8/Hbmr81U/EXqeUjgMeDoROlz9cP0kZEO
gXRC8gP0zvZIWpWE4gmzhje4DK8aKlG/l2LLAZs/FbGw3YIHsq18pkbHhd3IMDMLALEXLVsXg1IB
SJDp0hMuvL8kZPZfZcPgJbnVSfF+VNZbO2wrdkkQDNet5SPSs7jqQ8en58do2+raXH8j2KEUYSOY
1Zik1TbvM5ZOwEQ3B/UpxvRw8hf5Gr3XB4TGpxN7CTHNEjWJGgQUc+WYBYHNpYST+UlyVYHM8efR
mrZLW2ugoabGBTyC2kIA8DYiYRtSl6ucIoMEYQ+iBRClPAInDDTLeHEq73c2vkCys9xdTJ0UTBtk
y53g+XDAiLL+51kO/BM3FwvyJX6zgpd+DwVgJzxdGm/VfY8emiizR8jCzZ1mpXnpIKmdmdpatgbr
lAMPNoMuf8M33F5maJ/7zcLG83A5adWZeLADjWVD6TMh7b8lF3n6cVCM3f0yQzb4MD//8LZS3bas
zlf/WtkLeqKhgJyEUj6dCHMY4YAvsWKFpcHUiufuoH39HOTCnWMFWrBxBOEtJ1grLE8jMVvE8CQN
spFy2n0nQ4uLKcK3DLPELlaZAreqw3HqzpHqg++wlYPzS02rx1O7gQW02btOQgoGhBcXysbbdETF
96/E+kORxNO3+5MAWXVnd8zmBy+H4DtD5MNEFwUOevwshUF1e7zgmwb+Dke6Kejm6yYZdAjGGGGQ
5J6qB5ks7R9bNe5+sEaqIiYTYIz8RfSMVJ3L0pNE0uoKBTkf+BAeJhi3ohDVp8HXVNoTi9oKNXkL
/Ao87wN4oB4XT0rEH+Qka2GrWgyriqnqmysfbKz5e99fNzf8sFeBj1wucCu+Fz+6kUmmAgW4FUQe
nKuLXRSqvlSRuDJxayfABt+pUHd5EriBU+ACAXMtGQ8JWHhG73LKuiPNSss7mo7AKOLo9X47jv2a
DG39pV0S9Nm9abNi7Yungw1W1i79UodyD2C8rNhR53l4syNUpoYR5wmF2rr+S1Lj+tGIeo4akYgt
S0VNwKNjhBSnN2DNZnENIWNNEtjxA3ccDWK02pmCFY7Sm5bGkNdvrYhQ5BMUvh2sHHJV1i9DXUaz
WDzjiJO6xJuGEDh1iZ00ANK8UhU/7OwoEdPP5KG09qZvHzPaMoAoGO3AhamPQj7XFszIMxZriorG
C/HMGGWBnvJJzSYMJm9LgY5DM2kyx6n7nRn3e/ZdzJ21cyqidhOMWoaTbQul3ueB25PGIj7En2ZY
o4sziajD1BfNLv4xBqKigH3h4Xk2bsKLKkJOIOAvttV+CYdbbw3ZZeKhgJ/aFGyFIX61nZKAfwQK
UJ6xU22LOFoFoHQ5kLfaIV//7f45dNxNSwq9YOkJK7qfZfVMQHI/CqcIiXcHuufY+V6FNepbsxis
krZHQdPv0T26ez5W8bJgEJ607DXFq+xF13hrrypUUq4LQmucB1gd0Ff96T7d2WCWZhTLVDuF4xVB
1cohZQt4yKhHqHl8CEq69yD2sBnk9QfG6SWNk5bvYmsfW79AGaCWen+PknQqEotcOb9cCT50MzGQ
x60l4F0wBSRGW4MmtZnCH7De39iE2Y4dQutCV7VPiFSG/UE+LrM6nC5m+A5AZI7JabBQU3kaT8GT
ifmcl3Wjqa6y4WwxobDv7rJLCVT7awK151veqCmZ+eoKuTZxP4vreOCyyUt8lA4H10os5g3ylNku
GS06WgJQTe8cvQqt+2pWIUdRS+YbXBYqvCOuws+n3jR21KSn/gEGJwVJYnkbjTkmaD7AFpM3s5EG
F9zeG2FTljrxQfzVGQubbQKS3LAweVIICXvdM9PBD+fJ52CjqwTkrxffjh4aYldHhTHkx+TTayid
SMvImrzlH0p5ssFBhwN0hY0wuOvMxnfgiQcGmoEXAkIZa0swkByvmM1IIkYSbm5FaTKL51VCAsfO
Oi/BuB1ll83vmz3i/suskKJ537ALbV7cxMwriWFh7RZqanPmb+Y1pbpX736ADcXFGEYbJvIywdwI
OewYmv/13QdXK7VLVUcmoE21RInNctx5JlK4ZyrtaSiy9aFXK/kbbaK9jeo6Cjm7wyfcS+ZA+And
mVcwJHon+y7lfp3zxlRSvym3s5o5ieWKYj5YLmtZ5H8CCr2d+aaTpjkLnC3VKjdARFqrXu237CuB
gw+Z+Vc7NrovEJcL/DPFUQnL/umHPAGl843vpV6wsLmPeEuunjeP3yyk3KSbbcNVxvkhzIXXoqs5
7XojWCkjWZAb5viVPuTg5bcZsnR/hF6dfeIMH7jpcDGAUhxNXks7b3UlBz/RofgTZnxrps4Yy/5m
VHHHMT8MsaNxOmRdPfuBuZTsrTJRNFjB/GPnojUFolrXJnB8KwCEhjLRd1OIhjfXkJWfpadw1f9m
S2fAdd3QaBrC3cXX/oTmFZL0SSYUHjSGppPulOSCupmf+LouW7xB/hVqI/fwIqaN6GuXEvNdGwcD
8RTF+ZWkGYDCg94ep/vgJWMZDgQdhKgk8iq2+T2N3dnlnMDPA1Nb8I1gCCWWEBohZ+FqK4EJv0tC
YBsQy2XiEfDy8juPXugHZ3jWDoA3wUTJVm89FvOeQOF9xOdCKOletn1eFXcKkDKr0P1TJPTSwlEP
xrDS5hqDQ7K+JoONiXPxsWGd939pcEKcZkVKFwcGTZ01POa8CJWk7GdtYuf4wIxqLZxP3uzCeEQ9
/6HGCIaVsUsmhdo0N3tjxyBi2A1DyeSPQWbf55GdhGO9e4yXb6dtdvcgxC62Qqrg575aH7bJcCRI
x0aV7kVeaIdwkzZ2M77RDUk7gk7mvi3LltvpKGT4nY1OmgCxYB5Kn9vmkAjte+HfPQs0O/2xXpxC
moDN1E//ryIQgWTH/RLYRqdws+26FyxjHJj6dKT38CHtAnR6CTIXR870hi8TOyZQxa0T7Vnj54TV
wx8BvNpdn+yk9QEvLu/+KVZFbDt/XiydAig8/UXLuLPXuMQTfLaqDEOZe4MLVFggsE36/r4mpVBd
yQk5OwjcwYcVhoPRqCOoy7S7hw3fXGsWlZEoMUPXbC5IMEnBJOBDjizhgS0SRk4rA0tTlkIAbSOJ
toFKM0rMjQCaoUQUp+ss+F/1sVDYHM5GCKL3EEtnyOOQm4fVRHJ4DvhX4Mx/vg8L6cSZS140C7Al
C5VqvBGG0d6OtVW/PqcQx/FH5Y+wqnTczu70fFtw4u0SSTZ3G4/atwg40oHMUvO8jahkBepIfRLi
8qB8OLxXD/b3wXtc9eowz6FOtQWaksfBOcdORKlmpOYgyFKoWP8Ed2z14FOINhdI2J8H+0fBlh7e
K/oyCP8TIbxC4nBNZYCuirx1S7FKmWZNhCltmyKNlQF7JPF5xspC0Zg+IQcQh1vOyixxF8qS3CVY
GdtO3q85zlod+FOBg31p5e8SjuI7vflRiUU6bgEGV3MH9bJJ5WwGrYPI0dBKC5UP4lJMvE5jsS6Z
VZhBI4E9V2HkGpi5KUEgjMIrT00IHkju0+mlZzj4gtWGfEAAnPZ17AD9fjcxqZL+VATcwCOYfgcd
3m6AJNZ0GljdVYYFnuf6v+wh6T0wXeX/+qMWXU/dyvVkMhltPR5zYUBvKkeR/Ekv8TzWNm3uLNXh
Rupsp3243qKtRBOH4Zzka4wpY7xB6iI5iCsUUHOs+QqC9rH1VjabErr0mRJ82/A61X9RndQbcB1J
a6dZmXoHjWgyHavQNnOXkagcfMhJm7WooFGDNBuFkuCR/KFepKYtabtYBiYQIQWJU/FO4ewDKkIr
fMXO7OEYZJuDrbLhTNMfORN3p1ZHWYmFmSMIOFSGtoMLEmAmsCRtJBY+zltvtWvag4gA6WHxGAKZ
flsxV1OIW+9Luy1+u3a3EvOXRUnN2B2uf8gi5n3cjmx4CT4BgCpJFPlFGvcsN+Awumf4nNiqcpVa
wMW+jpsU1NDKLJ394YBZgDrn74wGBjc3aYK+gfHD6IVsPcesx0lcHB5GAbshXJX9xyXWrbjhzgse
1kswOF1wDT7j/zk27NfYRSiP6poHnoP7ZLVBUgXSyM7qA4hfw25WDAVxk22/+RJBxINV5T14tmEo
1+k6OsotBEPUTPboOFBjTqJG1p3u1+ZhHTpfmAmXEgAPPfaelslKgqiWJ+z1IKWugZg1f9ieA8Fh
n5UEwhrMJB2LVrMmqTDjZIZd/zHtb7uCTZp/sR8esJtcbPMcU0T7GtRUgLrVLNO/qzJAiEdyRQpS
joQSThKGXzEnAlEsuY+Z1TNeAYoCGLEAQKtEyAe/VPX3PHyxQIcV6uIX2DshJW4KgzxCxO5h+CTZ
L77fIB0Wv7Z/8IdFGeYzHeGRaY0yjxxwpQVpQbpRi4Gsip9Wjjx1po4BsTyeQprzADOwx6wJUk9t
XOjAmysPc6MAKxXioJPbOSC3Qyx1P7/u+rqcFD287TrUbzkiTiCJKsyEEuFkGAbqjUcjcwBg/6zl
QeNk1MqlMhXAXhIIwAzDEueaPGts2matc9PAXSJxXmFxyN/KtYBHtQ9cBlSvi8N57cEqrmGj9bqO
iaNU72ZB+6Xruw7W23a63yRiih6B4cKjHn3mYu3H7I3xlIy5G42ohSwZxc6UAtic8A2B1glkxk80
RxmwxLeSvaS0wPTMzk+Q3qv0MCiL2QXqgKmge9V1ozqx5A55o2P3SJJ1Whf/5+zuLRvK/TdmIFHC
+cAAwMFSlYnoRPPYT77xwtWerJFST0IrA1m2bmHZaJeBMqvFBRWPTuHLXDtd+uaZWRV2mE88MySL
t+9pokgTAo6jDMh8FjgIWDTAdIv6LID+IZDgGR7V76rhywmjjIRQADMEct0GaTbofdgZAMp4oyC4
6YecWG5+Qs7ybtES/WLNhtS8VIXjbSF40I0SYsIXkGP39j5fcyHOoHHpqxMPBPMj7BzU+KyLgJlz
8DZFENv6U6O4szllnARFroAam2muf1tzUodZOCCWJBKXTWSqhGBefU6WqpRBAheZ4h7v2r6cFk9H
Z3VVx7CE0e/Jy5cKxh2JjmKWVwxvsjh0vEwVYDwHS3VW20dgTbCkuEKea3+RuMHoyI4/J1yS9rHm
9qtmWaIqhy560998okiZi0ZJ6cR2ncTHTSPYizijEY6dHygXhFzcjiGCcTMlck5QId6TgeVVC1/Y
pazksT+rk4lbgK95VFTqPFHRj4IstjUbvabQD3iXPZot3yFZSHabhEDZTUmBjuria+uePKyPyf+e
g2oeHmjhSAV2ETgntcIn39E4BjHmCE6HYjs/pNyPAHKh+9IuFu+dvML84QZNScOm9jwRPpZhGFQI
mha5NUc2ATl567dqwkZou+Edst/Wr9I0qu22OEH4mBVtxyLG9/h9DfM/0RYabN6o7llYrHEmkDRg
kijYkV13J3cHtGC9z7xBmkXQbWJ5iBXO5EsLORRdkluYh60ueBfTdNwWsFHf5qn0v37X7//ELYBf
sI34OtjmRf+4jVwm4rN1qWJUXh194eXs4uGtVrhcKmyQilZEPiyqBfJtyxZsXig9thM9xYcU0P3J
hKEqJ7kuf2Ddg7bV+qf+YR9UEa/yZest9QnnsFvnnPiuCYPa7dGESPAge9HqPAGvmxqswfMzvst9
YHKfooh7Rgy/nFj7NPTIVpGgNJrQLzw65IZu5qiiNYv04TGoZPg2FqLtERHIuxu4rPoCQiwX53UV
xZqiv0ragdBCLHdlZ39DjKRMOf+kRI5Yh9MHflFM25ru2giroNiQsBRcT7u35rmCuO8WbYCxIaqI
Wt32FHv2YSEDKkLPnaf9jafWyHeKDzyF8r9D9sRzEuMAz1omhNoAWRnemCqkjzf/nA4EVEGkkFj6
U+PI56QO1xPzXcFLSw90AExnmXG3f83ZWD6ifNkz82V4vuFBfqhUSj5j3GxvX1Y3vJkIqE7nP+4L
5kqtUCTiQn1VKm5bJ8gbAPXW+Gu3SUQe6PT75s/RsA3oVB3YEy9GqGavsWK50ZfjTn0G2mq44BCV
VrZe0MPXu2roVZE1FMbHbKMjMMrC2MOO54rvoFe6Fzb1+DjF+CLgmwDVGfKC/QjEoi8H+E5i880W
m0IzggQMz0Kg7t/g1M3r3B/QHC604LajRMcCGhDrwFi3Al41LX5x5EUxcPoTPwwfEe2oKBUUp08L
wC9sB1AvHaAuPy/m4v3QQgFlA/OaZB9UJMfDi33JsBprxzN4fQaG/5KfNsTH7XV6GwU5BEgP8wxq
lf9hSk3O0LRrXSjohrWX3LfPDdtp7OtEf7smskfnsLBnt4r+UvFX8hvV7OihvtC/esrFXFaX4pZf
tQKlo61LgGISaO0EmMhYSz0yz4Jp2t06JVVPV1tu5QSEsuyu4RHEX3axiJyOPQydvK+N8pRu5usm
tQ1cQ29qiFm10l5hrVrcV5W0v8q+85yKzSubhKK5Mtrv8qnt0LrqmLjQSF5dHq+APBR64C6gWKB9
mOrjl87vlbNZxmgA34O83yNnCzm+AlAFQHK5aycm8d652GRUgPrQZtCBgzCMtmtRkU7ektheQbsb
ET0dRUiQWK9qgymsAqLLQ31lQicZgsAdzbQT98PVTDn8gTFoG15fOcJ0D/F41jYeqAphVnFXSaba
fQ4jiAPd70qM+j30EilaS54l2jYAXmcpddbEONQknXnSkHet1WLjo0nUOJ8BDwpiOxb6xm6KF/cW
THNqgt/kePdMS2a+6fnHCf2fWF3xlDxQIHI+Cl4wTFJdv1uGxypjMe2vBJNmwU1MtpkJo44a9Bu+
4Jzb/Tf2mD6ZQRh+X/tvXQwbnjccTG7Kfjjb0SXbBeUjmgfxFiYnsD+JQl5xl2/TQ/ewR42IVatd
y5Vt8rOAcPP4OB6Co0eQquirLxdChA+YKLwOUx7Abc6CJznzHVYmC4Y2za4uG+k2n0XxYKpwpJWd
7/uhJowTwVe3DTbjC8PpF9ppojAFGQtF+CAGYkvlzlUqcHEUCIWPAtfzXNS4kTaaMARcSQzHWAUm
pzHmhuLRqrM+2dfNOXwZPi8UbsgrIV61xDB41JX4GeMLugKqDC9IqIXlybU7TJj/lYITejdXWdIV
hGamR4CpmjV3NFJ6ho/g6WIMqNgKvQEJ12p3xOwwcnRaM+oAUdkSyZ20FQCC+eR8SOSFTOlg0uH0
NZqT5peZtVZXTenVV85WfVrNWRrFcEpBizzyWR0lO9Z3IYfO7y5y6sihVdoyrDZET8qivze5aZrf
5P6/MAuNk2qSsqDrW4UhpiJTNK611/PoVl3HyqUMXJjoArs3v37MAM3uCvqBRArPZtZojzIAz7J4
MPp/z/+ONnKmmb0RHQSKjy3gLgUFcxHxqORkolgv9Og0F5L8/5ECPhIax8X/KaONTOW/j3tp81PA
NqvReHP+BITkBdFaWIXbUT2VXELCrqJRRBVh5q33Kr3Qp+o+Pfrz/h79gAG+yF8vjWsl2yY67SSx
rGrw/g/3eVH/d4bMIu+ZG8GfZZABhTQSQBCGdAZw8G1eRpebU8ok60pNwnLocc7XRBA86nIEy9XW
QV/brSXDRuad3pK3xwAS4Ex13x86BwfQB+65TAUKGMX2vwe1vbD355DFwF+UZG0JHp39uHzpcSlK
gSATgEPv3U7X1Fg69JFz2vzEityAEg7wJdAJxup+LYoL4n6FHdmZwT1lcB3NzchDcFuWP2KNGf8C
wk6wF1kWS8sH9CTXrqFnsnIybtylpFcd63B9f/dI2Il0dXqcNO3rmV9mJNY5/8X+HuPFrvQe0War
wdgFDBY1L97bBVVJ9g8EoijrXc34X6vSzXqTSeaseFptAmIuSzRslQCAg33u7FtMJsHXv7fe62G8
B5o2/OJBvmtw2kMuArmT/TsFwX6RGV3Tvmb2ZZOs3W/WAARMUntFQsq3UeXKslyyZCWyq67SF0zf
NLqAmz5Sf3WNtrgi4JZpZkK8MenHpI03j4OzfXVl0YAwUuLlNGmsOlYpBN7pUl9lNcQCtAksf88y
l3DevVfGd5zkEoLIHxXbiQPM8sVbzgM9TbcaC+nmHWEPFcWf5au45whcuDo/ImXjlhatj4qjZFRN
yuDHdUn9T2kHSGSwYQKGENe46k+E4P5EnaB0URkTdU3yKd9eN7ttKD2PcIxu4uHO7uYGstJANe0R
NWaMR511t4qySUdakpXMpKoTaWkmOxrcrjpnR0SjoRf1v6CLPwvjpN6qkw8GJXFK1LiM91/zjAvk
6ZdoAuQD+1HY/4TA7cD4mt2sFgy0uHiSAmK+U8/Q/AYUJM/uPWBiO2rLfj0zihtI2StxkIN3NS5f
EhKpbrAoEmh8CAnc99ub4oeaVKBUc+44S2FZ9qWAQBOSKOUl6EFVh6uYUiBMOnhXK91TFsdFvvnV
FcIZdDbyhBZaVSNSPTZW+GRyt3/6Gz22UgAO6eU6uCVDAGjUJ7MOMYBqFB5nexpRegsKUz5ZhmfO
I3m3c+DPz2bDcYxIzjnO3siCGhZZypIP5r7AWFGXglz+x56oxnmICUrcxRnUU8RbSImdBvbGbb3l
P2OjFOqXNcOcCZn2tXrZvbx9dfsdeqQrsxuir5vK5jASPW3z8SuOaPQXCmqqpn1aCTOe0yUNlZpH
z79th8Yyadia6xjbTngK/sfsnVLAlwuU44AWIwLLbHAm/kZd9lu42ZYfndWyb9JBbvHNv6uKl5eV
HX4/kzO/quDIkNzkkBf2rgio5I+oP3rP8KiG466w8qmNzKUxM6HGxCgOGYZLRSego3ZDY90g5IjW
ir9tbX0oEtflFKlRF1QIl0XxRN8l8WdJM/9AubwI3llFE5IkNE+zMqgO9LkglsRFVR2NvrdNCe4S
Tp5OsYgZ7uSqkUjRq83vHvOXuRutMDt2UXf3eO2pRmIAC5uLAl9j0cj/X86z8jXiSQiZG2CUKW9a
bnMS1Vd3f6IT/7y58jjWgAr97HZzzjhdO2RHkJNkUjTDgFr602MEDH+zYioxZww9hOp95Tw0gmJ5
mSiU4165a2r4VgMfcKvJVu3kuvRrk0bTFCf9gHvH0H8/9SH9Brdg1uAskoAhuJFOt188mgnx4RqE
Isa+X62/InxrWyuSS5QQG2LC7EbqsVOXY0LMRqkFgnSYaJyOGYlfHsEKe9Q1noR/gDJSICC+Gido
2XlzTfFF+lXlgmhlBNVZ4SQxqB8mI8N4HrAFXSrsGtapTwROdQ+HeGeHIyW97y1gYBwFAADPdXHe
c5U8/1xkpqqxZY8PjyZlb6+nHoUDAAUhYSJcd7DpxAIGSBhEpTZ2/9k8O/O/WpKOj5GyWMjLAFA9
x30LcVCEd6vWYTLYTRtZcPN0a0fY5GmkRK3G+MYhdYRHVF/UQQ2l78jcLUahtDzfN821Wq7ENkFZ
cyQImrfzLkl+Hle+Gy5WN3Swop7wgFpZx85MEmC3Ppbr5H2W2R8hx5YOpkmTw9GTzPWfk24AGE+X
gkndNnCG3UTKcdc+3894F4Le0vDGt2l2NiXTqHHh6d9mxfkevOj17hmC+zKr+yPoRXbmvzKdljxt
5aInHlK2Mfu9IaQ6vluBT5Kv5mazI8l6CayZe+56+e4aIkKbx3UIUtqeLmb2jYXoTzhW90E9VH1H
KjlO2A+0PBTzLVrr0cQqLdo9BPqvMJzmOdMZVlyjs4RnzNr7Ul1IR2gJ0g5sQIQXNgY1xFqdfN7W
snLHeVO0dxdETUfnx8mWjdw5C3MYlot0yHfAhVkGIxANphUijQVXney/hlKAS31xUpRhPAhdfZhP
fxuXl8s6eY0tNCj/dOQkGS5uwC3rreK2OtvWX3TPLRmDDc+sGfmH/rMufrQL/UA3nG/gXbZZtOyu
3yBJc6Fqty33q22KW7J5XCQy5R4Cn+rY2ZHaj3ZDg/RJMFEseOYp/kB80IrTnj6Ru46uucjUmccf
RXAXT4R1X92Z0M/9CupcKpROg08/Vp38TdvvvSDLxPqySXBKmxNxC60BrvmWgnZMjSJMdUlHmL5H
fqjhrLao0BOGUnzWsU728NEbgemOdE2upp3AV5dvPO9Ri1bRGnCzSaWu0fpoJlApk1k71XcrSacg
XHlCOj1wD/sC7vs4KoMRlZZmzagZeBD/Qq2ALP91bjErkeszkDIOwQX/kzbsxlqEue6Gnk/uWr3Y
iGlNxHeIpFwnT9I+Y6Bnzcx4YJqcSk80YOUKzSJgWhNFEingi9whkVKUQQfhRY6IrF1Z4XuPyFjq
QDHQBVC9j3Glq5DKk6vxi7Bu9eOI7lT8Obx+WIitK5ZghaWBsg0jQnwjo0jcQX3/w/tZlLBqQq+A
jwlWrhfdydz65t+dGGZwjk+h6zcqREvghbEhia8lsV10/U8dH6cgXZnAvW/yjkxKHrkENFqoMSun
y5ZWUnemFPzulJ9bsQTeStf+GO+BnGLpvHWCcMQbAZbpu2FKT2e8lNto6GFCHVrz9EJFQfXS0s4k
bwUnZpbLuwgIGwOSyXS4K4l8YIGiQNwSdUJIGOk8KnXUCyFzXhbJxN204oSSkpVWr6XGCrONF/TZ
B5qPCq6VLyM7krh1igRhwjmfFGoQlPVN4Q8guw2PhCVBX3wMYK+MqeSYj57zIAZI39AVCmIcgCff
IgPUhB1ep8J9Lbi6XXaN+x9e50G0j1/P8gBttDpUDnpoFX4Jp/W/cWMIu0GG8AVDyB2uy1aVaKWS
I03Y+oD0a/P0vkB291S3icNX6x0g5qX9vSfy9byB1n0wFy7ze41Hx9v//H0OUsh9rulgCxAEZZfj
nug02K38ZkNkJe9dmpK0U39Jvvw4OUMDOUxn3X32T3xdKzX6NDZPkzpT21mQopio35yTMMPLVisv
hmxFaTwSeEGHhrhtxy5S1WrpfBUyna4WSkXJDYu/GkZyAROY/dj0QFRk285ds6PjVPtOwdfGfEae
LMIPqwCKSGRQWd1bFE5CPMHz94Yr/PBSTXuxIDlAqINNdHM31UBmhi3CPxUtEiSHDmuApVXbAQ3I
hpUtLj6b17JDrppf1KDYu1XRSuRaBhXOb8V2kBmJQDdZfRweUin+ZIPuD7K45h67Mgo/6jpsOtI1
a6DtI5LNuNDQvA2jk79Wdgavzp8w/uODJVAxAoM/8BdcrooZ1n8Yki/rkM/n2hKbjs43TKy+PjnD
xVEPGnv+rcjhFnu2rjGG58EZGIk4yd/fpvkDODkUUSItiZRPZcHrhbPu9BDac550HtU6MoTWvXk5
0q3SkGFjY6vjELhyP0EEggiQly5P+k86uXRLTN9/orde6/FiQkjgNf1fvTqcMwxWrN44EOf6JoYy
hh0UyMjybCjcNLoeEQwzsyB0VsPlSEbbBky/PqL6tlEIpLOi59glX972eL1ZXdrTrHdVXOAc4Ttj
K1bLf3XjDcQBc/4fnLXe3l1s/Yts+jOJN0ZrUlvHEDBgmfstMcUR5MsnteVivibhdwbLmWelR9yG
le4lSpUNOcP2jaZZle2/SmchYNiLJGeXOZsBdtshmDweS/E5U9OJ1HjXrR/s9RCKO3hZ8HhdvVw2
WJdGRu/U03+gIb8MpqDocc73/ZjL5heGO8W/E8vogVTjP9wxdfDjm5RGbxz4MC2k+Y9yOWY42DEL
3TJLaE+VuA3mtZu0UnImcASSKMhObDP8Hh2xwY7JTLOg+KRlXAAnTfnvpnjh7lIM3U0GfdZTxs3g
w6AzvzpoVEvlVZV/xJSKYV3BMpfmkQyJWIxyME20ghkMHtlVdYPonoa/JCbz5ifI9daUevNnC9L7
CU4jpPZDJDSfMSbFibUHoP7oVKLGoiPtTfEc90sUgOs/YFIKkrdbU1Pq+WEJ9Mw70PSRpOFH8uJp
jhE6BNFbB7EOmtSW7bUjkjJoHy9N/Nx9O+utA1mIrkRbD5PPDwc8gQM3A/5gKQp885G9BO2rpzhb
JiOcO+KjAR616qTJVupt3BTakmkIOHkLn0a/cIRVcAd5H5EBTBrNYIgK3g0+1hl2BOM6bYFoXN4M
I0Q/gHkKWjxPgebXKj0a/8FPt+W20glV9ti6xxYgZ+jmgM6/uhEpE8fKSxGlhyDHssQo0b1qMGzB
IhRjSRB3HJu0wMYqo2e6VnYMrpm715bshEFbw2f1+EaooLAWToezhEoIHUVF10f1WFhfGo924qee
NT65qtMZemyKRk/KlL8YRn2l1JV44ziwTsodNB4KizdtNAfp6gS5EK9xbblNDmMgEYqm0Tcd0a7T
2iaIqcLtvZ9VQhWqwHbPwMV/kMnO1Car0wl58W372oCZVUPFkX3STgNbobbDhQg05H4mASPABJHd
914dPw21rdm3z3oU2nTuOJDM/YXb+tChKSYlM9T1lAJSlRzp08U8Sj3nAOAeHq5UlUHCtZ/iX1zk
7nI/d7zyU751REZxuET4rgR8FOj5BSJUl7asH7eHsRYiH2mdtkfs7WQ7diipWWLK/oMfB8/ulF7K
QluMO4NIMp4oFtb0JUNornmi0JThsGGbVgidg2rwVprQQTj+Q1yV9wDuwrD/CbUpyJ/eS3yxKsFB
RoG2psdqB2NYC94A4x4IcQ+6DnxBavSf6m/U1CUtCkxtNhkydKSgfLeHWN7a8xJknKXsMQC/6T8T
fO7fTzE63jrKuYlIAcblTfnmJMdwy9YiVUIJjmf08Ts0B0A5Rf+wbj0yLUikeEJcE9NfPrsZXjNk
rfpahJiqnego/PcJO942Em1NAZPlAJDkQW4C7smD04A+zvQOCTCC4Emki9oGn/e1vzF/VOFZKqud
HPaQyHdxGjaPf3zkmo6poT6By9MxupM9x1UZPbHugq0nfF/Y69Cr4N5g4zVFewjmK+oCjWRuQP58
hdKWaNiPb+Jz3rRLxZfIcePXfb5xXaqTYnfjh2/zLu9WOHCrnSDbtO0bqpnbT4QjDuePy+cL43IQ
3rW3Xsoevblbk0XCN4P3Gcc4wEXU+IhgaBIpVViFXvaNyE1JdoTQO7iR19muA4Jp+MLEhVSF0+F8
5cBKpwfkhGj0EKswTzy+pbpvyiwmmX7/hOXrIxNppyCNHAHDl7AyVWDrX7DMlhF+wtF/7e2wGrgs
bIjmb1/gTCYdmk6KAzlT5w0tGH+CL3wj0PwWEhrP5kW9WN6amI79450ktj7Ref0g8cIrXYEf7SXr
Epqcvu2tbu3flTP05cpfz2fink1luCAack+oR2mXYiEXHLXGiINuccmuatwHF/8FQ8iRZnany2a+
hZFrtNjHrrdpdWuegVtuQso19qs7LSqKeDeMge6Vu1uKG5cEI1Nl0DhN/jLYdHETlc4q8ODCSpW2
L6L244O55i3sG0PxYG2FCQAvI4b9Q0Ym8x2vZQkq7YZ1d352JvapjfzxxP/ywHDbhTxlcC8xhQ0p
Hd4fZqez9iHmIZusP7wpi/Xn+yD0e4HqEeXw7gmXw8BGXKoERVZPtxHDVWbTJtJsiEjf3p5X5IH4
QIxDRvZBgX7uo4mtcUkti5GGMSbgPV+WfNDKy2K+CjeuQu+6UZYzkVSbIZ1upe3ww/jkHRA4YFJp
8FQKC0RRFxrUzn+CwjmjnKCnXNdmaKgI3caiu3wY1uFPWbhEvzmaqTIbkp5OmVpkn7Wlp2W1L+se
gLK3rXnvLb8TPor1udUZGUsZZ2UXVedECnabq9UShc7r3XFDzMvgS+MG/Bj+DJRh5NyBWTFtfKAT
ipSc3Oc1VvSJ7I7VXGVM98gDMd68N7lqWrBheZxW+8WsZBbHZUSB5WUuXOfKpTNveygmDHqDC9ZP
DDjJ93H/AmgM4TiygL/BdeVFE39zwtYHEsSQwE6gNjHkSV87ARJtsESO+eTqhfHzTb3IF+QTkcJR
DYqXDMobtBWYaOPyZ/seD3KI+NaDXJD00Jrw5pWUXOO/kTLZbIvwnFb0tyDZ6I/nbcw+k9bhrnYH
Z15KsyHaCYtX0Xz9GJNEnnbrdtytzJrAEP9Mg4wqaFpL/JUFjmJk7XUn+FcXI2sQNnn9feVVrHVk
Js4fIiPl3ZlH8Ak2i53Fy55NXsndHirhueCq1E3tOd9wFy2x0ZzEchmxv4G096o6LvAtEUMqDDRh
a648TN6WKMnTseCfxE8cemZsqOGxE2cokcfIjpX4ShK+uO+pvqwUOPLyPi3JiFV9cDkD+E24zyni
xTWT4RqiCf3m0ZI9uEZdqz4IUo9sW0UgVu53aQMIHxl52oSpft0GWL0n2B9LOElVqXhhmm9gT+th
60UUfNJXy8p/W1UMidDWdadpspYjmJUtmsReOMo/dUP6xYvToEjoYtNPzBl6cp57Z7VNbPOFIQAm
lelIKzkdAh0qzvxkzmY+3xd7GKuWFhffH3kK2Y8GFV+V4ap6LMAQfdzre2KWhIeNOV+L6d7BvyL6
Ni3OB9jU1rqg4xxYnJxY9Yx94CLcLlbC1uzY1gkANILJIOCmqqoTTG3Ihb7+u1Im4v80u8Lkp+jB
NZHPO7uTgi5WGThnYREHKM0CPye9NEHQkGk9xsFS1h7/qzri3lH/rOvjdVT/mgR2ZNCKk4X3tO91
0uHpnDRqT7E2XeMCbEX76av/Lv3np+UBembcqnhtdTKONOO5/UhXIQLw8RJlP45sKjaTpvLpPtJl
CaGZoGKPyrraYIBgmausxJPBSnN6EgJTTMSbNnPusegE6SdDRVusw54GLyUDJ7hERAgqB3g0Sqmj
CQ2lvbwLwmWOXy4rMImkyRnT83eKGRaMw3T9lEY3K7PxFuswypbLvEkabVlzI7zNQG6oyIYkekL6
ADIf1FOBlWanhJddbN1n1DiA281fpilL5BQxfsfMlDGOXAiAo8NuBAepvEc7JVJiE6EmeOW4jEsa
oVVJkkd4qF+P1iDdlvJGNGKOkr6JsNnI854yNPFWO6ZEPcVycrew0xrFCzzfSPlFIru9X0ZYY2ID
Dw76b1YKixs7o4jRIBWomw6M8oBl+lyXGcMNDIu4GKyomzyyjZuAzOcOavyTUd3K7gTmi+POcUvG
2BcSjfA2LjVE/sq4stZOz1xaALCvRum6T+sYkbZlJ49lLI7xkTg+Fie616cINgbp7K/UWVnwzaLA
ONdCEgottBnpz869Ajp1ZqUKrldXt05s8oNjjkih4ct2able9eRcTimICVYRKq31KaH+OIqjIof8
9FbPonyDNVUnrmUaUgvEuVBVX9k/yeIfx6g0PN7mKl4Anv/8nNdRUMpffUSwzdBprOYk7GIKb5TE
GBQJ0UO8ZtMicSGVESiGdRwpkicptx3uG9yxoXbypf1JBBqRGdBhHIrbIvlnGLUBc5bQGoOOxgK5
z2VksHz5jxel3mc6sVf8RSFuabWRGt+uDjB3b8f1uU0pffrWsJ7LYroKjjY8aKcIt54pBdVhQJ5k
gR5EwYklCNJ0GKWzkHgy1ploKOzSis1z3kFL8zOHPPYtPdNBex4kgkKspt3gBohkhvl5YEddoU35
HDz5nn2Tl9xd6RUkqW+9VREIfII1oeW0CZx9ndpKD0EAqHztTLIt31ZslCCHQGdTPuWo1hV7AKk1
YxCGwz/buWsL6VI9Hi+YqYcH4NVHDChkgL1jKNC1hwylpv4cUIH2xeCl3Kbs4d5+Kyux0i+fjTLY
Je2qS7NDKUTsCl8YsG/F7p5SGtUxqOVm5rIj3j+ym5F3MvW8yKkxPNIO8j5HpzXS83P469eKDJp6
OvBbSiYEoh7QohwfiBPyWZkhi09DAun6sjSTvYmTQ3gXmUIGAar3aC+Be+Y8S7YCidWfQJLY1zuB
u9oqdCpSBpDyRj5bhCne1ssK1K94RPfQdQJcKgJWjjsfe3zWPiKGP6VkTVJLibLbP3zwcBCPBNgi
vgJCAzsb66TT/HsOgQLb9edkLdcxAB0QEI9rtCNiMotI0R8U9vTy6rUe/wjqeBQ3iuPhMl6TfOU3
xX0860TU9g8lbJPmkGZj/KJqdFqFqcmGc/nanceWBzt94fMTCdqKvUOMxTPTFfUrnnjiM60iro+1
jquDqzeLWzXEVRyVz/zP2yS7fVyNG1GmFAG98WKc5mlIDLY25ooGK3ZABYvwoiZ2xF9OZY7hAGaf
YGXViKHbQY9TGI+49tpie2W1AQcEsd2jZHqadM+hRAHyb45q65arktUd2VtZ0dpjr7myIA1OMraK
XIyvfPsjWbaFZQtTwFFBFW827IgfhSfeefKyl4FAwaGn1k0wkhuYF5jA1FceHFKrU/IGYCHOuY60
uKESKVWVEA/CvjIczBVunrdAxOieAOAW2a5QrLYBZYaH9FhQZetiaIAKKqLjLNORc8LQrOVJAF4o
vbureEgSwcMKWWuIF2tYHyUglVrTm7cef7am6e3DTpQo+AYjxSy0nsYZ4ZhxnlOo9iSyu0Q/nZUf
HEHdvCHymVPYZeoUc1tcAFhcV6yWLShPl9UitWtH2+q2GlAIppE+w9cKjaXs3wi79jDae0Z9i+U2
b85+/ywdh51N3/AU1O8n6QxUe3NGMOupI4+KOAdTkVbz/zrjlyU6nOLOF4+nj9JqZsCI0MNfAi1M
RgIYWqDBedJqkF+oV26PpZg5E3pxh6J76dV759Bw2gCQFLJzUgw21orp3Oc3QjKDj5ibzQGTVSHP
Ye4asUHi1nSsuQFuhlLfqiAVY5tFq574eQLp6efk5WG+waN/05fWtbJi1AoqNMYsmSxigVHlhsnj
RCiqyN46eZAI3jUPRhehhOYEuF8EUTX7ySBDpMl+Kp7yfHCeDu5ymtRiM8E3UMz6HsTdFqe6SwsF
mEO39ww+YI/EXH192dTY87NuiSBeFvVx+1nYehrRxhGd/W1Om7bKIXlZF6MaHO6OwjIPuDdb8+8w
Rjz9RRP8jc7hun0fFxpUUw2ybuVjXtGd7mLvXYnwIXelUgrYTPWhPX4pxGcACorbh1SJUaEIq2tn
rD2tqz0p0JhPsDBsqUNshgxKb2EeBdJBeApXq01yZBifK09yvEkNjFEFqqp79mNzzMOPwpR+jT3P
ONldLKoEThap83sGid5LSp74rf4TmPkjz0wPppQ4n4o7NFLGNFZ+TjEbsrLvqn6iPt00Qutu2oYg
oiBSHGu9X06W/4xcCKTPw9TcTlVBn5fDtvd9hVILh1TZDFAfKh8HkFJjIVt0BD1uf2pKqT/iYIW8
lNs8YOkxDSLOUArPHswuZb37lD0kGRbi2IsyTooM68HBL2IS5F4XIuQupJDvYBUvBWxGMSVYVag8
EQMkTOt6AbNCwj4JVeLKjw3NGCpjb0u0cbLGJbc259TJOtGnsPehPvqOeyFWY2oy/N6IgMxYQe2M
zXbQsEzLrQJ6AjMoXtlAe35TF1gdLeQGzIdphHn/96h4Z495BHd5ylsdhe9Xt87XsxY5U3AmgtT/
1TbBxNb0DkfO/ly46GE/4LsuC4JxjuzLiAHAidEdhKDHhd9DzB6z+fH1++4U2V/DjCm4Ylpx3m0M
ryKWpwS2YYXqEjPw/rv8FbW0oHm5ujj3zul/3VZj3KYB0k4ySKuHwMWiIdj5mVzTLzOd7m3eV7vf
DQ3S/r7VxSYWUsblRYP9Ff5kr4mSNkK/5RMue7mwjBhsoif24iEZdkORdus2x+j+Oe9fi7MHyqbY
rpS2LYm6YYyGqAB/L+tna42OfPzCe6nQGfnNmwsgac+Gj1KFyWhlT29YgpkHbslkH94LJWpiUXFR
LMM4wbl1qeIMq2V53HWNrQaVLQV+u5S+Hky/FvgB9Vsv2Lgl436IXGYspwHQlMgokdD0UZ+I0uEl
UeUVb/CY22n4MEaSjUEU8/JfWKz88DKPZWoDL/J5kDn/MrN3gdFNwR/QvRMUctv4TGcyCo4YDESW
S2orM0JEXTT1npsrrkJ1bDiX+crKEF/LpcDizOjaoxMd7vDcUm3yjBNfq+nL5PiVuE4j50gzOz+E
alP2gA9jVpR1ivyL+v7234Pty1ZOkndaJv8j39GedywidzY8cW2kSxz393rtvu4KdDu+4LaxkPsT
DMjEbdY219iFQfO0FEFDzoG2mFFRQg83LpMNu2G2UbG7KqyqCu4ARyVEXQ+Juq+2tI+MImp3WyG/
ocU0X74fYxuL21P3Qw2rbLaPpKQtUmSCIj/Q90nrPdkSRdNcq7matDyteqgyueB2wnmb296PsbwJ
+sFIUD2Qsmpbw1pIQNErkevK/n+2bHekT7cFrpzk15JKm3fl0iKEGcupJafUdTVfVePN/LZwdmjm
fyF8+fSDP97Y8CNi6/QzW3bx2JAyYXN/DnHPcgBSr6HtBWlyGKUG4OaL+rBifM9o1pkfOM4f+HJq
1U/XaFCLCAUGCnL03+rUDCJIQwFs+Yl0SI7TppIOAXsUfREWELTS/H1Ag0/Jv5qeZbZaAGlFTWhK
DqXHjrc9hTi+02Asx1efcpU6cNJDauSn2yKY7jN9x8DPU2uFbNLnXPDqsTHWtdUtAU4xbs5/6Qq5
MTfi5TLfqyqHVg7LWJwmOqKxjPIe6qAfFL4Kvy/xqjF2JBOVs0RWXurMMdQU8Gl9Rl4iE3yT+d+X
1XSeaviAPjm67h/3GW4f7lAXKn7wl1lBEvo420t284eDp/si7yaaP7WvLjwQc7z09YIiGFMqmta3
oWXfbR1QCEOQziCFOkAxbWVK2v723NBIo3LzpzWyrVFg3p6P8CV6fM+TDp9GptkfTkxxhrD4pZKN
fVO7C6RVEHSZaA+2nDJiQQetgwiZ3pENMeMqSDQJ4gkkjOiytNghxD41h094n6KB1gAA75FQ1o0R
u7jUWw0cUBKhG9pehw+LPpxQCRGV88tMPWB+KDAcn7PfkgLvMGPfmKPzfS154rN3SIgMnSMRT4KL
lsmBQ4ysxoq5hOU60btbuarbQnyQyRFVlJtxvL9wOlaFpoltGCdwXLxu15HJD3PR+6PCCyj/NPsL
WIKzbvgsuypC2cwyKIhC3vdngFr0ZCdKK+DedfZRvndWK4/JKmfpHkWPkk3/G4aNPd/HKVx5VYO3
Y60vlx+mTaQ5G5Uj77NAtJzCp9xX0iSZ2thxH3urHwIhqdKHBCPcRdhSlMl7bkwpUsgYz9d7mk8z
BCj+MpGY6kVRIA13V57ANAv7xVqOsK2JWqgdhnWC45pJo7EyKz9YPF+plmhwvhRIFTSSXSFAsDAi
r9gNMSSpZ15Um2gRxaJL2/8JxZdutY3df8qa86yhVV8bRucIM3zvERrveK1jZb1NlffiKSJxzxkE
Jgx2PcLxwvLXwkB2baUcjS5E202BR+jerXR9fjU8fc6oVBhxthWJwlzXDhpAOjzPV52wszUTCmQT
C799wZrDXEJAxl6O3rMbDIu4Rf5hmXior4TYeVMhDt+nI86LuH/tgJGOdXOJStbGSDi24+SoTHux
CBHFJ2AXGDjAOI25GDY3IBVV4rzHzuTF0/ySLwcNePXGPRqsky+4fqbsIQ+Savm9th28AoJmXI4o
8xpy9zCxQQwxcFmgXIaKUz7jKiIzXCgR/j0NXMZ/jmxwmrVg6lkWTOde6CeCpkBFcUOtRT4qF0TJ
uQ1gMu2g1tk90EhQKKSYRFDioPzLFMg0N7RKF3CnNJ28inX0u7DFADhJzZR3Eers4F47utvmaNoh
J/wNsNPyGCSW7NZRzYJnN8ZPXtsUoLlkj2E9/xIco/enasFaCGVNSFfUroVyz35ZPFvIXWVV7p+l
SybCTtmZsSV4gRJMDEl8A4is2A5An+RpDBH3fpV7Wza/CFPBJGUtby/NsjAkJGAJ+qLUvcJ27zDP
pkt6Z8eQpw9N0lexG/wiLd/oBe+cO1mghiFNOy+3UbLRDucl1vO5i7aMCD01/Xpb0uA59Yv2ouqf
g3x+OXdaPG1UT0f//x2xW0BRs+Mo2qNxUliHBSzI+adIU86OAB6o2DxiNPnmOH1Y+3nzd3D49c1E
dI2cy49dcu373LEND3AtVD7ExXQnkPWcyBoHNVbAufqY4qeUYcTwIzn2WhEmhadPoE1KUzuOvJsF
3Ysp2rwryHcPUkKg2wWso8CY//diEvwIBKXbA4200G5+WMiipjKzD70p3n3Fo1V0tzKloiGG9pzh
K7FO/4lrZv/OMoVw6weCZEmbelGWkDCSk0drgpvrr8ImWmPjsm0ngFna/zPRcmEPviZGkYqdkjDf
7U+B6nU0xPKx/6n+9mn7UZsUyfOz6coMof9OrhK4W00RkSFWDja/k8Hq3bL4B5Pc7yKStfYmb9sx
JZKSGlWlX+pgETVqn7Xrf/EANLtiltH73k4fyAqy3tC0aQnnj0Wogmas0h3dwwPMKiO8bg92PSxD
iMKJ168zs8xpCPsbdmBwoRg+FmutWT/pTd5JwGnOXzB/ndr5bg0mIRAUTMcDxMIxfWHPfCSjfMrA
+KFA/j4ZceLv84YKfREH+wgglncyR21R81sYq0odvqjL7Z3VUGDvagkjvejbcyYAF5CHKU3TCMkp
YbjewlkD9V5ZxFq+rYxZ4KWST1eSx9Ht/BczcomzwWC4xK8nZNVwRRjZkfD6hVtq5TmiX8l2RIWp
uLNDTMbB5/2POjscvMJrDEkwfJiNAPUd8IbpufL3xf76NXS9hUv5WUC0OjPpM25F6XueU9SGYttg
2fZjddHxyT7rYuD4FcIYTE3te82Gyz1HKhsz6p53kVkCoB7T59siyTwFnt/2Wl3Ofy7uVVukT/vl
pFcxKIvy+5aQ/fRcOC7GzSIJ42f82dQMSTiAg5LZ54jQ5g5gzN+T/0xD+7n3CCdbmD3HcSMEwoC1
jEZLuYgVqa4MPIqPA186BJLr+B/Mw43o5NUhRj0EwTwCwqWsggr08GvXb2DRtLUOdhNxOmxCpVc5
OYOWB4YqToEfQamYkg/w9tljxHm5gQcuQ5d5pflHtZxhmeBdgG6bT4OUF2tTJz2nvP/Mi7OvuYRV
UmeKFHCzwFnOla0tQx/oZniLdJoeffXqvKE6ZVbCbVZ2gbjwPJLM6NQDmoBk2YNqE6bTIh8p3ZmB
yq6E2ip8Gaa+L+MSpsGgTCR5w0kIU/NVfTeDgqdENVb/GAWwSladUQ3AM+YyxABXxJfGpxHnE398
99qaA0M5IAup81U6txAmgSHSTyExAL7NbRTkyGP7KFkurA5SQuMzEgWJQ2ma7cLTKLqApqzYc+gx
/RxCgnT0DVxi7VO4c79GAu0j1kkm0yksHCmphRU5YxIqp1xJurNgtcGJQ0fWTwU6utorBNMmdtVe
Q+a3W4DO0DiZh8Ti1Mpw8egicgyUoDE7qDaF2cav499k0jTYwCar0MWy4+5Szj9aPu3iwdi7c4pU
AaN7JXaUP24wKF9IpHBOorWCBZhvA+PR5PeULhRxMB3qEFpr6H4h/2N4KTwCXaCjNHNmK5X3PWKj
0jshXwczYQ0H2aXdyMP4IsV7hCQz2Z3+xoANqVSdBlgzK3dVxrbOV+cR0PediFVhMq6NERE4Pygh
3C8kYubPLPIlU/C9EmoGtNuzQKyhCSvB010hZvS257jUI40h2ChmWD/xzIrXnJ/kPWsHh0o7Qcuw
Uki+lng+6H9yRl2HZ+fsx7nPE0sYRMLyByulIie3cVeKu5w6mbbQB6heDcF1ksCz1zNOxs0gw2Z7
I02kYOZvR+KNNB+nvuu+2jfpU82J8IGsnvrPpxWXCiHGf/ics0s8x0JkDJGwu1fx5BKuFY5lA9H8
od362BRm+NWOjaSTVKIEGa5AWO8v/h89j1OkX8xSrDgJ0fwqmo/RMtaV8HGkOxFk7lWYvBhaPfO5
GNBuXGsC7LnDaqArl1NxgsbknC4YfkZUGCq+h1Y8Xbt3VuNbKZ4pMhHz8hAceY3B+wUTNIflxN8Z
xncpZgH30SRrJVoMyT/Zl0dannI0hydOeRFNXN2O4g/igqOOUERFXfcqgGiWm5JMcTNTLh5CSwue
d7OKZ+HmKo+S2N/XHMF6j1LKydPJjWR04L5Eh0uebWwjRUahGyyjzQ0e/gLmhpHyUM6oJFVLgBq8
0FAQRQ1Wq3xRJIjptj7Viri0dGgbXb2VuJbdw1JMB8RXanq4i/aDt5vNHYLGMvrLhkGGMr3X/wtG
f39IV5vkuYTsHivYn2p/Rr4KbbZ4O0ZDioRQRW1KAkc6asZq0VnvUMDQAMdjRoQgKwAI9vfaDwpm
3EXa2r4UZfR+TwtzJiRhDGhJAflXTGLLgFMRo0Fml6BLXIUTSeuLTNV8WC4f81vfkAXq0Bc6OH3t
5gRMht4+wQLsJm/zd48FviqJTk9neeyZSlb7qdkW4eS/irwuRUXC/1byavYl/OUKyzGBRDqNhm2o
XUPDT/v9CosTgNd9NJtCX+KCglEup2NvzOw0o9u55b7OmQYL/FZz5Dcxxlf0ddjugWERHwHSCfv+
ik8mtdoB9RI4V5bQXlK1iU3BGQLVYKiOpXIrCpntBPhDgVmfKvXRW0gtg8gyt4trv91grHrCWu1S
QzH/ookkjMo+NmmcJomDN35GOSTPcqv6BjFVRj0DqPgt2/gZ6FjpKq/h9mg71GFjGIsE1h5eqLlh
/EV2lj036KCeTYdcvl/s392S4hpKY7aTz1roWNrEHI25c+CRhs+8ed0sZ2vo1RIUNFJ7l1LiDDgS
TGt1lX05e0tnFH5MeR5PVpk5ktQOlo2R3TslI3QR2XkryGOsS3/GvUcQBDIVPhywbzLbV1GkUZqJ
lGqWzU7KTDtlC+TV4eWUoZKdrw/qUO7DZDVZ472cUiPVkFAW6Lo/mUdxU5LI3/T805L6XVqK/sYJ
C3k7nTIzTIu0MkKgNB7Q4YbQMdHILmcPZpyqlflsuJzZJP4p4CfsiAaMMqpaNjdFXTZsbj30Qf6Q
iSOqHRk1FMNu2vydEUEiMI0TqM0Tn5JfxfJP9rhwAMBne92OH91ioSvqjRjyLOYe8Z2VhEr7kaFy
mkBtZ2y9MIrM3m7ZhL9Ykle+IDrW/kzROYwcXfA11nIknz59RHp54K37maycaJQ4oFYiRDxSSTOG
4zNpoOdH+Xg4p31rD15Dcn+3oJ+yKYm4GN6RC3dq3MS6NeiqTlOQzQieTPyGG6yGYHBNAtRSdM5H
79x5ebsF9cOH7fy9RL+/xXnabeDCaTSmUonjy5jR8X0B1CKfiex5qsexIsJ8tUZ9PTPNyeKIN62d
pbMkyTT3kBXf66rkPubmOLqd8mOfnBLkIxb3DGkbIJLNgmjJe8bX78unBa8X6BxSUoZfA6zZX5R3
yD3wxcwNdM8cdLn6fznjtPCPg96kuvPo5gLd9tJ1HA1h+rXbJDbdqXtrK6U90D9QSkhw+OBB7xHY
T3A0gkIgfdPchTxgSz6RzJpq/luxyIUDUziFStbOsGIgWppOAacLHUgw1MGpW29/CtaoYIYYNHrc
DkKHnB/ewjBpFqhjDWeTgQBMiq+7SFf4srnnCGKBwGzs5cUqLOvzqwfRmMgHNjs7weSeGw7JAla2
lOo7dltZRmIydBCFGPwbZQBgBrjCmmI1+qsmOjlSkyCxQy4DEAfBj802JfDelkaNL/DFeYhkcpmQ
+FOedj4NRaTcwfnmQRjiQNoKbqKxGnuVcvOA3c2CTbuOD+GjklH4wnXkeCWcJiGGKSds0uj7JlyS
nYbhOonT+1T7f2hhVXqKwu2skyiyNSCbWsU6LPp5/DgO4JKODc/7YslXyYfkzhh+U3gTAXqGozxw
FPJp8ewzxvs3Qa/NyyObq47Vm+f+F6w28VQITDTXe12majXtglxin9aE1Gy2wnqvRlPQpdBB0vYD
o8tjDKb2fcZYnNKVDY6opzdhgyPz5BwVagwoUGtTAS5MlwQpGfJVeBBEyZOHW0lFSpCdBckIZZjm
eGGGy5Rh9hyH2ov0l38VoFC6L4FxQ/N1t1+xuB1z9tIxruYSoBIrkowQ66S0E8MK81ZpUV7SVm4x
x9Z9P3ca9s+RzHwKhcu7yVihaDorcTaplorlo5s7vzkF/P8wqiVbuxC91MZw2wFn/BRMFjj+WnSb
WZdw67TIgLyHfZeXR8fUmEgmP3lGLECJihEGUFnZIJi8/Yp2ipSm35RxQb3rzA6saba+5BbcnTIe
V6vMZFS2QRPqY7tRhE6ivMm1Yw4PAZxiKgqb9fsdfoETY5CRnFbKWrvbO0rZl1UTGpmdLaOw9OUD
2N0jf77+mApKTUaHps7pfJNl96AE+Ph5r0mpvyKb8tDcqgSfq/Ael+JA/+p135XrL2UShBTY0IwN
IvR5HFvaFoX1j8Pzg77DTHN1LM9bJpoCYZFxB87rT+nM201nHtaf8EG8uRSTmCso6xijU1DLM7zB
s2HY0O+7aSYpaXFBMNXUAZr6XJbjKqzXsgNaVRcDi3IClh4E6xSk8aaC5uPBKuRnGVazl26wt5HJ
G6DbGXgQjGa1f77J5wDEUMtKbZBeJrqJ1fm8Mm7bq1Z6lP6brp+48LTlF6fjEU2Di7fF0PT6ehGw
aTWpW3h4tSx6Z1+aT7S2bplwK/cvwCbzcKLzWU47u7gVIAbowEqCwnfaox71cMUeyx6omuDTge8t
kJVfUjVD6F0exQoiF56Z/0pfPwN+qhXVaRcJrC3nMS+f1ubVGcoeMNPkzqIIKA9SqgWB0rit8K1D
IFAF3r3F8J+jXK8veWCpza8SxlZ7q31yAgVa4cEYWFGLGPNHkaKTwXeiXCLpglDXa3YkOnaabrSS
nfg0bmq5mhfCLUoS8SeBcCgaq2pxWswONPiQS9mu2Z1l3unDXySDt4xaGBlYtDMUa+cEKHvzULEn
kJT6XXE3EACUT84TNif0OIQsgMvMNuU9cg5BJW2+HvSi7ZkumGqmsRiHQbrdw/NP/QF5ReZ/odCw
p7eN9gMM+QnnbXqNf0XnuKHSAxSfGpNh6o/H69joiGpS6u91UPq4/Kk13wlZC569rC0Dw0fSv8CQ
vke8QBkMrtaxPXcFvFOZG/77HIyNWpFz9Fu4LNaIdM/h7M9x3gg+kt8ZNHTTPk8FDn9wO3/ljMK9
QD1B4KOufimNwx36drkasmhbeWDxwsO7LiA9atSGJl/gl1+ODj7vkEkNZLqc473Y9WM+MWe7KBag
ZKB9qVkRL3SEkStzlGV/GG/36b1JzPtIoHJWbU6CYD1XrSv9vNv+XIWfZ6ZvEhEBMgHXrpqpqUOd
dvY8ywhzhf6//OW7UlWUfmDdB72uSVKbF4myn6qhZKoCtpfMSNxKgu+tO1gelRiSSds9W23knfv1
ltENO6xLxYyQhiYGC5iaMLcin3lH1VhGUslGFxCxGCFKhSUISp0M30CUhBrH+s/SqZHipT33+AmC
28r9vGrhPEYC2pQW3vPu13/yhcWrzBpJrr9/gfz40gGsSM45f5/BwUBhZf9DDhRzpUVPiRE2JBKV
Qd6Ln9pQ6571jbOU5k4202y3XCcYT4fKzPby5qp0TE+Qb43rhn9CEvBVvHbEBcoDH9PZ3PhBFEtC
rFsMEum4xJ1DcPysslHsjgIuR7Pm06pMb9wJOpDtFXkt9TVsRaG/euexlz87MkI/eNNseF6soK5r
Ct+jJSgnF3PzVEe9uGLlPXAMGFZeYJGPnYzOjZ4FiR6tBQONl5Jd31GaYj3G27phC2nv/wUxh41w
q/Ox2OgA2RArzCKCF7RHYAJYjVpNgsrJd/1Y/m8ku0VLgvvNun4JU/8N9s2ZmdkqSHe8PmchYYDD
HranJsPQ1cnmJRg7tyOKr3pQMh4Zs/F9+/3izFazD0XeaBsTpiShRl3fUqW2Fk32pSNJ8CUWDa06
Kp+9oVGrvHTGXO/EbnCqAALCVbs/indg4jT/kDAAi3PL8WvLiUymJpsSfXJdtsA959opINhMro1J
C6UiZzMuqAxDhSNvhizIMOJoJhW5kekTiDzZ16uslCMl0c8cHX99i3xLwxJazqkjv7qC7f7B7V2k
y7LzvnQ7jMrc74y37U2KD1wntqjtMtrxCnwCifOdZ/pe+ptxdL4b0BNaloCnzY7aflDXfbPv//Q2
Qhx9FdBGNZiK36Q1PaR+y882o+IpcbnGDi7T9qMxEfg09sgjIRV5Pl5Lvau0UjBIOB2+3hUjCiA4
EuMwFNgkLR4CIBnKY4a99QFm+1HSsPxRA/KooTU1jkC9+FAc0TD+uW11Gw7HySYoq8u4ijXN5J8E
XiSF5TBDIhCFR9J0CBS9ODooa0UjOj+VCQjcoE3v59YTiH+ClvKO1T+3Fvb0PBpyXfGrZBK1qM55
kcRDgB9d7lRIOTDyrHTT81BmzGGFWFX2ym53h+njqSBG4VnkfnLe7/pSU6vetMoKFt5L3TywsMXa
NbTapxEqFlyYHo9xOVjASTW/WscwdbzamlqsMpXfl0BUYXYd8SP4bbt3FXnsr7tAwpJAerJHQ2pv
HgIw0nFAEEool2V7NIoNc86DlcuXfgqX93YLT4xZgZ9BXBn82u8uCaQpPBjn86pI7mJNGY+gxJIP
wsc5paBeDRRkGOYrsYiD/+WT6QDx1vQGZmD5Mt+Qb/dX6po+dg7rznnY27PZsm7lNHKpAm96oyrU
4KUITNXxsdvW+x/1IbhEv6ig5EKerP6KBR4b4sbsR8QHzca5IyzzXmyGAQcFueUO/3fPY/ADfNYB
pdsyS/+4RKfxDuRP9UhCocfOvoT0Jb5iB9vGs6yh68wn5wTIN7wkmNgHKuewAsCtef8cdqbUGcu8
O+xcgD7u9ZujOot9gBRMif1rxZbFcZfrSeZgk9i7XbXom6GZHys6eoevTF6q+t71AApWqUHqhlGC
HjJQ/cfTzytdPfgeDNf8o6A/TutkN1CMJAyAPiGN43r0L5hitFOr0U9sf+y2JnOKegNnaD9mJ6Em
pOSegKnITrScRGjHwwUXP4wIMANk91uXIXUk5PH1q/aMuO+KErcMSFCOqPPUmzb5oGC2KUu2Gi7l
zJpsvses8TevB6eukB6gGQKNV9xTX3YwqYK46TwFLNJ+94S0TuqjvUXJ1Ib2S8QUpNowo8sMS4gY
By3PWhm4hYiracQJbqnwcGpnW/DrZk6WeFuNsxZhf6jMQQXMTGzAH3k08iBQ6atXbVqGyyrvz3pr
LBW/fdgT0QQrL3+Vx1WoUzSBTAWInmVm2NKrBwNdtygnfS/X72Jnhy0YJlGf3uPh82X2xu2/gBuT
n0+1MWoKSa0jTF0bQd/LSTjSaFlZ8PgqVh8ptfwm9twG55TXTc3kRj5Sae32qyDad1GzalCDKRRv
SNiYhI92sa6ye4cPxqXqwXe9PLBIqoziUE/TebteLdW6/LZ8pVrrS5LHfF4S9+0nIqOMfHKvNSyy
U3lzgiMSzi0o5QD9xO51Fn/99guispO5ug5SxjfWfSNCF1hFGulp1ELJYd79fF95exKZR5u8pZN2
KqlxKOF46r4nJ1tGp8Rn7sWmW7GnPkPx+j/OtWQOBHhCzS9wSL/TkFN2eBm0t6ktYjEgPDmn3O6h
PJrjGCLcrazruu3Pqt1ir4kPfnHEBsxXlsQbviyhaYIZ5+wwQc+OKxCm+HC29+lQkH+GiwcI6ISQ
Mptly43hoSxCtc097WgP7VOOg8W1mCKKjPPcEsz+E2K7sF/4QKMPnhvclnFk9FYu1c5EmTqsUlgs
4wKsdsry4KcyolbUxOHyiORqfh035o6uUuXVxbeAEsUuMOc4L2cH7iuAUolXpFq++0kWeuFDp0Dh
6Ts2pRYTE4Fx/D6PBBm9P49rSGQ5wXYXCs5mFh/2urE3TIrCYydet7IN/t/Eo71KocRIgzPyyiNU
UzZCyQQY+SSZk2ZsJQ/QPQqjg8SId61e1uZcQ8gXRA6oYbl/EybZlcf9Jw2k/cmrza7YR6i4WVab
9W4KKl80rBmC1guluWO4sBfiwkaPpDllUq4SZAECyWUHElsezorrxuYzMpRUfdpqndOKcuRHQoFY
JY7xkGPJbBTlufPfw1CqvrlynsPivzT3AeqbEnyXf3jCIMeSVgmA6Aze/e35MH95BNviN9ujz2bP
I2KPzB17f/WwcnUXF70R53XtUds0j2wugXQs4p2lNczzXNndCcanmADiQDuNXN7JenQpnThugCtS
vvLhxyDK6n6+hb6gRGrlqrZ4Xd35CTVcvSgN9U6N3zeZo61oQz20BD+RZprCZqAeIpRBIdjlka0F
r18cOK3dQ/YC8Ba40vZ4D2LHrkdzAtw3EzcpdYr0n+Y0IxLT3ME1c2Yw6bvPCcRovoNtvMfeV2KQ
/EFBNkRkwjQ/28UkQFiv60EF8Xdtyfe0tK3ezq5k5v6zl9eWsAe8TKQqxENRZi4pPJU4L1HYhdLK
7Afudv6FT3gjTrcffS1ifoYj0Eg/lEgrLmyt4vRLSEHKMegGUNoINuXTElG61WuIlTImJx7Rb20n
rn1FKGBSe2B9xwuH8dwKPsaRvWnrYA48bdDWHQN0d2G7Hv2ppbcyJdAwLtBzh/vcygQiPcfpg46X
L/TiJ3gRrfkrLzJeMTH/ENfwTHOMC1D9XybstBnf/0dSIvrRUMHVncJBLEQcmghMeliMMpsY+WpZ
i0K2DLhlTdg5C1fM5BDjWWU/yH1M9/1n6vnkPZ6ns9djoWnYWYcr4MnWlwFv1tANbjk/M8GFZrUh
B/BtnJ4lGfNDqdPOk4/tbu7lDrwT4W96a+QfI5qqDq1AH1I87G0R5vbhHrR+1eEX3pruocfzI5Md
rdPXGIX+ySS5ti5vPSxXDxlXe0LI1/uT35a5tyMAVI3O6FraRJX1spgKgcCLxjdiJRMn86kXLSp6
lBlP5D+sxnP7B4znoma3gmBXTCZ81yX2qE5d8iWzX0q2usaD4Sm4RB06Eed7wtUX8R0c0yvbhZmH
zHQNN4/x4TM0hGfbx6iCZNNaL/Md8J2y5TfgTQT/Rkd68UGagAkH2dyX0j23CXm3HU0N/SHP0qAh
Yuf4Yno5uSR9c56ZWzQpJh8WwLG6EzO1Wpsx4dOQOGc4FimP6WJjUaVl+fNDMHqEf6lq+zIcxtc1
+FtQcq08X40dJlcOUo9cp8qaPoESRExw/cyScsSCQpUoNFi3fm3otTt4+2K3Ub8Qfh3Ghl+8ERPF
Ox1b1cBokeQSY1tMYMFIMlRq9+0X8b6F1eXvrNstDezzCBqzj0AcOJiRrT/i7xjgQUXiYVmy8NC/
Sip3QbV47eArO+VaUzXlLfySmNpAMJVI5NCop2fGpcjuywUplveSILlxSDa6gDGmS7X91RmEfQ0v
d0SwKFVpiqxuY4gdwjTdfZlAn8mJ73sXsiglukkbWSu01lq9fMDP9E1RgxbIwf7cHrNYrWx5OPFb
HD1Psco9YOIlkz1Alig+LJScSS2QukLUXE8Ax3KDcYmmjwo9KshXo9JR4kNMaIxWaPIhfrHSB99L
KpxCN0PPOm8XVnLv3X3saBhk3XRS3yyqxOQQ7hqeIjKBWATliZDlzaSjsgqOsB4l/R091T8vhayN
x+5Xc3pba2SRI+PT5BaHQEshQqP9I2FCxj9KFzeMjHWdxYD6Fh1/RVDae8oO2/GdnL8ry5CNB70Z
cSeqYLiEL8/ZNiXm0rp6bc+Dei3t7HIXub+gJvgtIVOANqMdt1nftWVgZ8fKTwwwZpPm+Gasv/R5
dxB6h9jvbs8/mKra1HA4YJ0PKZW0h00NzKpXHJNAC2Sw/hm3OBlEaG8ym61yJ9IFEGJ/b3/trsqm
z6PfZWNSSA00m7/0L5ASPdRXLtydXJBNen770PUzGozHkpqBVx/0gj7Sy6Px9ucVEmdvpeg2jAyD
gtxrDBOOTylHkWG+7THAJuIthqFRi9TWG37+i/RNkSyPkOLIN/34w7K/zOSAcdhsDXnMb27UWypJ
rUTDldTnaRvwZmlUmFO4UrNhjfUnlsGn42zfV5jsgsTe1vrXmQCZtBFpHSWaIYNx00X/E/TKa2cr
4ZfECAdH/oxZ5LGgSoJ+SwxSW4VHNVEch5rFt/2xNoEGsBoPZbnNzK56K4JKkWaGiiLCQFnZlroU
r4DOlUCahaxA3EGgKw/md8D8S2Ntls4AOhhN2QYpOifo746oCYym8KZ1jC15d5atBJkP4Rjp1OUs
TGETmZ/41iwgeaqEYctLwVdCZFyI3qyRN8bNmgll7D128Viu2hx6I/gxyvHuiA3W4sU3dqZB5EtS
v4qTFjs3yKjdUMTyqJBkj/vZ98PFGeLai/+1lkgZ1Lc3k2Aq90lDsXwlcA/38Agt4oXKnbhOS9YR
x5lBK554nd2X9qSckQMPXp5TURzKlSlz4m7lwMFcdDT4xQ0Xq073rfU3dfyiq8dHu0XNWmW7Bxpj
owf/OURwKwJrbbAvenD+asgPULb45++08ekgcVlbGHCUaQmTaZbVC9ZTHHxsT8lBu3J1v0yU9CzJ
IMzR+ciRxDXBKtm7n3IJO7FLTxrkk6URseiJ6WyK56ZHSn5gCMWTLUiANuT427XFCbbKteADGL+R
Vu0lCm+TdT67YoLiCA0Fv1t08LLjuGLWZ8ATm7mK89UGXqbsnVeBaTzIhAjylwlJ7obQp19EqtIY
cwuJ7pDXOsGhO1Z5SOPT+voq6mAZGybgWbJArfpG1abGC8XNnOc/HBHEMY8vWRHYWVHr9M3HsjOc
4Q7DjYHPOvbm7IPFMN8YWOWs3RMOLICaU1I5BKXDAGPUNP1o4E1LUx3lczkqAVZi2q6sTIHuZwqk
iVZXAZ7ONFBl9C02iMg6iYkH1yyHPo1olL05QTSBhU4PPC0DlpmDljbji/9/RinFGaFp0euffEkG
hNYwfs2kK8nfGHdD2nBYeopOWsnyepYX157Z3/CUkXkNps5bqO/0phlEdD2iJmfhYAtXefHrRqBh
grdNujWi11+7wTEXKo48AHXSHCXQecuMejkD+kGk34qOFWXCZS+LbYuoQTc90alrusFZmm1FnXzN
IFLpQFRcqKaW/y1pPYRoOgkJkQpaR4mc7zjYO/igoZPkyDtXIO/Tb5uaLhAgkgnldAGQv9Gbj81x
RwBGWx/BSFYCFOArDsWbLs2i8ltxE+EPhGQKhZBcDv29W+68mLcPJ3lS5zgxAD6X7IbWYkDETqtu
HQGhLTtViGOpxJCLi+3NFZv4mkFvSDgQPob18Ghwjn6Mjj+nXUReLEPdwIcPT12h1tMHjqHAPfJm
wEDlNHCVeJp/Uer2iC2GA3+y3YRP/7dIAhbQ1SiEiH/OVIS0a3ze1qdCPerP5fI8igwEt14w6y++
M/lGKl/sJaQ8PVmcbHDQsvWsHODpkgMHFFNw/phx1S8WWSsTUfXGtvzH85m9r39W+iQAXESX/Lrp
QjounrPhbTY3/g23T/zuURbuS52x8LzoRgkJpdMO/T1j6xNd8mpR4zbC9VSB1Lpd2V/z9hxfVCdB
L8V9ZR1wWwmAZnK1jsQSQnU1L3MRWj/Cz+PdNQv9HmuJoid4hCF2dXKiKZBCdVLwImaamuxlWiEb
hlBFKiSe584yvNREoOAXPU6pMFOEhaGDbvSZjXNgoj+0Fse5ryr/r2Kv0Hp1BfUW/1tBqVJoAdM6
U6xKIVgTkOno4Nt1Nz1VnvqGhyk9iS/afIMwL7r6bD2OaiE4F3Elg1sIDVGKKvWTEhT91sJzIL7S
F26W8Uc6Ap2PuASzfNc6dvn+6/DWWjA/N5eCA1B9g7XTuPaUL467/bXwK32KFczwooQcoUrTFVP+
DEr/bhcBJE2e2tEO3iolUIZDtayPk17/BVsEiWuZ6RRfI1k1d/gJnliL3buBbmRHfhRCSIJ2wSju
RlygBzin7c7YMVASFh758LCUWC7gtYf453m7ZkB6h0aRGK+cQbRMlPxKGt4dex5GYZj4W1snDSg0
dAtMtfHEHr6VEYs2Z2NVxF+61szaL7OFpwsvT8JPuzssoNF27qveu7HSnj3+p69m/R3jXWq8xA0q
l0KHac8ZOViYC9JhoO7uaa2M9UxvPbUEWJzO1axQXsHPoBxIj17E2mAbj+5YlUVjb3XZ30NBxbt3
Dsth4js93M4wOJELXjR+2zB4oYA+HPbIwtKVI9jrSeBwdnEhdWaZZRIGeSOwaxbnbtPJnmhdys2F
EnLc7mXtnCUmwwZnHg3lgz8T+sewXmqjaBSzTHHJFLU+dSXXAqVIrtpo/7PE7Ply1AzrE9DX+nT9
86o1WU4rjVjoBJ//tUucHEoTuLqff0LmB22GxH869JFwndzwBZuPl+sS+MShP66IdGnaNAP+DQsO
nHyA9s+iMbYAg17iYdVYGwLf4UeDpQ/lbYzW9JOtGGS13wE6RIjzdA9trGQ7vIBsZqgFQnzixu0k
3GqOMEmW+NRaJ4sSY5JrdyTVO5KzReVIy/b6S+BISKoJvOurU8KOmYL2ZT4TWeAj3lSHN8ptLGm0
CDhTSEr7xwEmCoTxLMOs1y7QDKY25Q3Y09+gZTiiRw4P1jyEDu+svvL+YvzQ/Fu6ZRzgcTy2cmNz
krr1l0xhmSj9XjBU19/nsSacD6U9IExnZlYziQDYDAmse4RuvQYgDHxCB7+B2OTBKeUoWGzSeFSV
CNFKI0e4iyhL/uG2ITx1qxCpYLxUWXblgnYZiPCi/FHKT96BbdLUd6abz03MrhQWyXbIYbVuV7fK
pm0V/Q3SyQqNzD6rBDX5F3McSn3leYz3B4XB7QtDIgIlwlpf6e9YXIj2Rmw7TMdGu5s/LPfNGRQ9
UfipHWyY6P12VdjND98sg73p54/mZP/OuCtmte618Gt/B2kS8Qpe/sw1NFPX9zoLWCp5EzJPX1uo
QLE3saPzQqL5Q6KqnpO8KmB/GfgzWfUrXHops332oAAV4KqTYXiiEWcmU8BFfMM+KsoP26Le8MF2
pefg4LXVfADMaJtK+qrIZHhkE/V/TjJQy5LaO64o+g+6yTm9lhxkzVnIMX4wdUJc3VXKM3vZuQzv
Ds17vI7yAcSxzuoUMI9pgEuZxSdOH14X1kS1LJ4g/cezyjpIc9wUGFpI2GOqbg2n7aMuMPjFH35g
9T5qbIJlkXbGEqlVUzv2L+IYiB9ckUJDhqwBx4TUlaePygk7voG9y38C3HDCzzhwHiMHea3Wahlz
9+jjBNcSYHpiKRMi/q43ATP7uJXCmvmeOCnWT8RNXLpyYclgRQZtDyLx5je8wU6iG4yRQYO5taii
s647io1vSScHg86zZgHlRKETEUk0tEJGJ6rUrIqURCzk1gJIQ7CHlCehrF82LVWWBWTv30ZvDC86
B4IX3SeHpprj0uXJhONaX3qsUcIEySE36BNIC5DQIGhRCIHmWL8h90GldUg9nzxtz7bxHB9zRct5
hL1EKHiV2taMXMl+iJjEdRGHebnl+LYGYo3CATx4p9gF2LP0JWY+zS82lV+eHJotv7bag+7iguzm
rRYJwhlxaSntEMUcKKE0zyJ80y1N0FMnT7U5iu+tPMAE0IlkeXMJ+HcIYohVLILB+flA4ojc/j0g
ENzu9J0YsjSQ5uqaqu9v/IFr4bBQe2J2hNT4XVgNIZpWEA1oBjg6J7b02+R5OnKbPGER9urgj2Cm
w00D5DGxU0V7D5aJ3YZzrkwEbginf9yWjIQ+aMyG8dLvucAK6UxCbWNmvs+rBzUON+Q1Um0btKCF
csNDtMQ9ciAEzxJ0PaKZwfeRqrzBv5PFFvH9GMSEbgdH9IJukNELb2no1HcpyGQK8CJrkpqa3Zc0
NbL7ZKUxKTSS5w/DxdpPy/jkLG5NHb66k/yAPNp4yqjCR5tkf4sIlIY64pXz91araxF9teLG7V30
Sqdpcpgq5vlzsSAlftAAHFnanZT6tpAtB+lbk2HfOnCVvZm2tQ07jtfx0qOUnpn79k2RX2x5AL6C
RZyufBkBTgydZMg9T+wW1nQHnO7Uzhct70fqLEt5yDtxK1t/luYsYJ9opMejzp+wKQBmWLprNInW
btncrQzDP8MG4gHLYpUkPO0xgiv3ewnBWkbl29hHTFRj9VJs6gELuNwfrmft4b25eaA/7fZTYH5S
igQXXzpF/HjWpREK+JC3l0d4WNHenkdL/0TmfHldfLHwMLCgHS3QaCj/SnVYIzuGrElD+0tPzHbr
RjhkHdoqwsUiuUO/NBZz62auc0OxPGlR0xvmrU00B7/v3oneg6e9xPB0eE0XpyEQfgunSy+51rgB
n4DEEcR2tnTdsoRpJMbiK9QhxZ/X3KnMVRVtctKHcM9lOs7Qm+7rcT3Jpap2xLr9asi3HjGyE5AO
pUir+lvgZZ/Eh2Kj6K/ot4ANqEdIqdBtOPRHSPUDXERq1DKnBRSrPc+Crg8a+3PTWpgwSu72PUjx
1S7/gS8rln+SEkhPDkD1Zsf8pVbbjEu74F3K0Sf61ZzeNWX4ATyV6ee2Mn+E4ViS0+MhZ2nbxzu7
Fd2UW+a4QAxFXMweM8x+tLIy4EXIvMRC9lye1O3sXen2cdH4m4ic7wRvpW7Gc4TxGpF8dj7hG9aw
WvTwut13tH8ZJ60YxJVnIfTLsbaQ5ZT2lO+tugZ/ZvDnN8VU6JYGYPVnUWIJuEFGIQ+WjcwZjfC4
voijvWZK5RmPxl5m20IR+cR2hQJ/N3aq0HeJcLnHOGamrBJG8yRXvpnjeeuk5CNiIfDGoMDj7NVJ
W1IfWtnI9LrYi5XzYNIwePJSWV9Mhnh7L1pNwUvjNHgTqVmPe4EoOGJmhbVvZGFdosmwP5olfDxJ
FAGGTmDXTruAtRkKvN9q5j3V0Gn80nyq4QiBDTT/PmtHWDFyGGhbegYy0PlOOtX4btkO3+RunxfL
M5DsCcK+jWw3nP7fOoWRvTGyu9dELzGkbwI6JFZ8CAZ6TxdUJjuSQ/w7xREmR/mF/8roHxQ49Yvf
FEikMacUvJ8T6LG9l18wVaDT0OXtgufm8/9p8cT0PX1t/Oaj+JNmWZm7cz9owhb88bByN4IUYsRK
qdGXgWu5auvZC0TSFQjTPW5axeiGB3FAe5r4dK/FI2UzUuw324J8gW1ZtRRSasLyBUuV9w76YRAy
XfPMU/790LGQJFyNoC5RmuAyJim7z9tbCCWTyQpJ8nzTIwtsJ1u5IMH3dQBM/h2hFQCcvEniCc6w
KYN4zNxJBTXaJU4hdc/VOvN/eSI5eALdd1A1uf73mic+QtegFhyf6XBcFrcpv9CBwILB1U/6zfLw
TkUKXL8l3IYn11OKLTzwr0/aUZURRV/YNC86zZV1CYFWZgdByVKpQ74rZJsgM42RcFYszNBISiZF
yAw3BUhGsrkK4h20MN/jrCLbf1eyl7M14ZwLje8ktop0Mj44y04KuipiV1FzoEOxpSOu4R819tjV
WMnpGKTZAryT7AlblZJEtcMnUsCW2vdsaEgwW62AleJBaCNIdpL1I8YEdeOUV53tegD162wxC5z9
IqxAhaxAIzI5+Bgv12vIOjRWSofMfDr+OUq0c0AcpXQTeFvsTit8FRcgZrc1VZE8qdm8GsFRqW15
Y3k+JPsJ0qXP9UPEpIVmeC3GX9IGndiUad5/HN2vA/F6To0URLHXF+FfruN20Kj92tVlWM/7AyMq
gDVfoYPr/tcWPOQkZ+CdcRISjgTbcvLTNQMuxZpo+ug3ySR1tev3i9hwhH6jIW7wZBqCQroJAuNK
77rAfVpaHdNxZSmf9SCR3AurfMAjrtLyNG8+EaGpA4mdarwwkp6ujH23RFIw7mKe5UrMDR5yCr6k
MkxiSkMBAGeoO3TcHzMwLet0FO5srGfJmej8OMWJLpX/pOwZRf3e68sYs+1z3C3+PdfthDUD0z9v
cYMElbrEj00t/AA3AUN/sjerLrJ6P07oiA9TKkiyDEBuvKuI9hOhgThQw3svXdjv8cEuDxFgJJ9+
FbdvnnE6XvWj57ppEkwVFAaPKMcLrq4by0Vnr/JrfvWskz2Re8WM+N7x3vSEjF8z9AUq8PROF7q9
19ILSnn2VAwEnl0Po7t3eh92Bcfi8OAQ479PXB7kQITlpzkjT3vlwRoDeYNbhanIp9eYikZuG9ou
hPyF3e8A2XLkxM1vqvZXm0gPX+3NHZZuPv9G5Fq9f+gxKXTHoaUabueIEWWIq4KrQ6wPmRqHuS+g
Tk3EwJaT7qyN0IJ8PkYsWoDe27T1krSiEYGOWHpEwJvzjwvDf/Z17X1xjcwlBvHshakkMETDsWqj
ezOpav8JN9dUOUKsWBJArxWMSHzFJEZqs/vHL3OzXduSoglWqk2A/tfv7pbeIkY1G/PjcU8ztntV
x1MaBntCJRy1JelFH6O0cZXbo8+eCds0j5LRXpExND9A+3UL6davuJuAUj0xeVDkQCUvw6KLdfCt
58u+C25oIkozYA5jJHlvTy/aCNAZDtm4ZAXA1i2cbMNIQhgilzaEy6I66i4MxoC53FwyN1fjxj91
/GIkELMUSBbKK+s/yGWK5Os4IqRQ75bI3cAp/te6jMSYtZDHbDXze5qr0ZMfswDIOqiIjWoacml3
nDGUG+5NJKd3cqkoBIL4yqWetm/+ZqNSvdjfoJ0jyp+3oHby4E1kSOubasuSvijszVv6SmvdMUX0
0r7JZgutUxGOlKr+XayBxZAcEYH9z/oo2u+7gXUyBMPo7w+sORJkdR0+QkoysLZ7gCNPnzL259M8
xXdssjsi0fjuK51wJrq0KdgWyen7C2u4iBS+z3OX0LVrCxi5ShQuQlP/jlW8NeiaPQGmt8lysLCd
hrY2bpnPXVN8SAb6gD9kRGITIxNEec0SFPxUjiMdXFHJjGXCqFl7enaJ5v2nNHJMtnPSaAjI3Zhk
r71OfAD9/uTZnwtlNy/vqH9f18P/q/b5Rky6+LS3EIwmpHwVnQMT85beNs+t1Fgrl1OvVrC9A3Hr
Iaus0E+Ip2crUGtrQ78337TG22wqGLc4K1erv7YrjRLUHIw2qTdQj/juxk/riX3nbdx8MxcN9ljn
4UICqmYZkTycrqIMXZm+XmiMaszLYCyD16K6o3vo12nJy16qS4eNtEx17l/A1t8BCvDc4NyoRCnL
CTWwc7c2fHk5nqVw2qH87oSyjloN7CxeXCpGN0mSIQaklIG9s9TWQZrWiWprOe7nMOOnIC9+jgeR
mtRNOUm/DbbUnrZqgDNVKzTH614EwUHQVRJdcxFuYfnL7TMcESgdpDmCobrefCvLwbI2lwFRleE7
82nZnjOXtE2mXlUIGbEqEHC5F9yXNuo5ofqMJGED7/mLKoNhHxmXvRrIU6H9mP9UQWuZN4pNKSBN
o6F+8en6soNZ78AVEfdR84M9UoPlF8dBYCrX4f1kBrypgMhhB6BZgka9u0dtmCDXswgPi/yBBPyN
B1HxHsuaTnU3r9LDDl1OEgOwbI/ru2TzElmwmD7ucFjAD8+mmAwoLOztrqyJ+Lpx2pyKaHKXwXbL
1fp5qc8RF9RPI8VPHti5GTOcdy/Oac7BXGeJeNMshuVFYIJU236pRocf07AanFh6FPA4OskKbACU
iZbfrQJXrHyx/7L/mb3QuXzkujg+66rh9xqqIea8nnWB9x/OKdKDTT+Neb/N++uA/Ge46NRH8IAj
sChyLH/H4qIdLSu/wemogEBLiHfPHwcQA8czShBBpy7Sqmp0Sc4JYqCdec48FjFfqoTVH8oAPhj+
azCITmXvdoUWw+PuvcVfwcaAA53XkT/urcKr/6FGMFGPBckFMHjuqTXxcJSPVFXGtIgfelwwYNf3
bGWYe6gqVCm2slZRbuMyCcSJ9xNU3cIN2eoQ3Uz/va2pjYAnsCGJQSF4Ud0hhkE4Jj5jVo5iQ/gJ
yvUAyybKmyytEGnuQdKcTzDcqVhSm+sjOtAUB2+JeT57wocO51uqRt8DEDrMSJtUqmb7HWRwzf6Q
86Yy2PNAYo2sjRRTrCUKrHpR0uR3ZNe3M7gEMeX87wCKkjQtPDR8F8KQXu/l3ICVkpG9gqKAg/1q
H/AQ/SVvcniWnq9i5HKvZlsMjYgjHprCZs7rLFDCWrO4D2vRgCYVsM5pZPXQ1UVS+nwijRMx549b
CaVrfHSvAeRdTbBTSV+JoJP8a/SQeYBAnUKs2mEhC8iZRP25ZULvoPm0Emk7k2JnNNOhFVzxAmDy
C2DMIp5j05/83zUe/eGrVmwxjLG27S9GmU5y2WCCMuj2o9zAenfGpA+Kuw8R+OsMhFGMSDSlNQAU
hwok9a4q/TCSbL+t50R3j9mz9t64UJe218CO3QjKa3RrZ4OdcGvMTeEj5ZNWGLpCyUHENTeNup+p
t0ykdcIz3JnA+5nblh2tzGzlxzEa7vDfqtAXaGJvZyy3EeryCuBF1rO+iAW4JRyYVxSKsLWPbLiG
oDunTkF0HPTL3w4SL9ROkQfCX9/fz3ZScRw+XIRVC7S3CURxGuMcMrwWa7sAlSMSg+QHeBBEIgPA
Z7lV6M4SUJt8/O22LcRaNPsBbnmv2KAvZcaZ4kxcTzT2px6UMlouGupVTHPPxL0i4aPTy69bVVS4
tzjrtvcE8w4kLlu2bz4DHYud066fPkM/jXdkikDmMdXLW2mHub3ntzTx5rrJiZodFAUoKZ4hrpWK
NyeVob+G7phF08RLkCXq/EHsslqhTNKztXbOEzUWn+ZLdhVuaDuBcM2kmV5qrVPLUrUIkP6mrRWw
KH8fDeO1Hh+jO5Xw68c8yoA+oUg5W2DwuNelSMhLGP/ycRycN0ikpPCJ5s4n6QpQh/Zpd5naBHYe
QtMz3G3Y6j9MofAxAcqeuIgcsUgc7aoWN/khG6mOHTu2snCzlpP5lHBIDhmjE+1ihfY18DE8ODY7
ILWDpiyi4TpboXAS3+V0HsvBCcfMuXX3dkUFtWrtdwihCYVtpwQ8MYmJeE19PTlWOcOxjvBmjNR0
xrvFnGnMZo9t61/jI15s7EHy3/UNzMfvItztEkGJPswOMnvyJyQ6qvDCmyfbdiXPTZVtMsP05j47
zNgp2veGGWzq6n1Sr6uryeECJlQsuJJpsC/EZ352ygCYJAYxd/YTVQRW0lK6ePCLj6fmkjZSBMpl
B1a+n6MnPbywJQ8pAGP9Fpdq2xMDEvnnFgBpdqcOlwnMyAQo2tGv9yrOrMjLIelPJCveDU8jCbc1
GOrKmsQn9Q0cnNpZpnV+noxpPYjI/HpKYfy45uGnpbjsM5zIJX36yvEigNpUZlpsK2NXYKaa/Peb
pqBtkaqVK8ZwPXuG3Fn7HBd9JvtGmA7YcKDwZ5FJeAVX6UKGyM9RGrHyuJx/xdt24NTmtx4IIL2C
BF4+Kw4xZzFRCv00+WUtfm3rV9Ml8ceQ/kdJiWPSDzszjwevh8lVex4yg0G0h1f8AaNzA960PCGs
densnEy1Qnf4ks6HjabVjoTD4EFgALufhM6dLoRzjbJChlL1V0CO4SdpCZVp3jHcYHFzabH4XzZK
zCQ0k3mvCAlz8G3iuBZs7S5lIr0uzxJW1nDjxt6P5TTsi6YgWWi8i7cgdRYS9Rge5ot/9xJpIg+B
IJg2VZeUdu09PD3xamG2dhU9Bd1IZI5SzbBpHywwtGOnx+5ezBNjHhBX9MLgnYPhBbUXG3bAnxV8
3pRhkDEd4szaE6EkHC4jgd6YK6ONFzKHX39obfU1zsI+Uz2pH7Xe9IMw71yfb3r0FVdqkCgmDDEF
3PsxNlWMJb3AJ3cIAbqmJ/Dtsl0kGCU0ShHDLOXsIR1/J1g5qUJVo9il4OYH9KKWniaQdu8A24g3
wuSam07qbdelux695NhuvTFwYqOaIdcJOG7yg3c5QaOGnHr79NTeO01vxAFKrBpXPMNuN6Bj36bU
2nw8rRK3a9AD0BFUo3HrXnv/pBz4yVksKfQPYvfi2P8ueogQCvrCmLLU4HrCYrMcIJO1H35yp1LP
vtOoTriWmC8hs3jPPZkNU+aIfNam5U+adK08xpneHsQIb6ncpHS1g/+sD1vxohEdwbleTz93y94J
iJGys+cgjFcD8xWcjxJjMy2tpCZiVVKE3SIr8FYmD4Y4iKNtbzCuYajJbIBq5JqqeNupAB3+tpH0
BhErftz8zecSBmPOY93ytgn6a/85IMc2vqZFuPW+P2Qms7dBIwY/SKuXE6KJfWzM8KBz4KI4HJUV
D2FXbalcg7Vmx85inS7s/86lEKVRyye7NxZfZa3x9B1VJegZp+ZuigwNDWikvsWgPkno4L14JhTx
+pMD21ts7ntrpXRl0IC1BAjiulP+5l1atV8pG8CibmSi5yAia3Zgfe3izm/3cFzaiDS47WIrIiP2
8/Go32VlZavBoDo38T1H2WU684FK0dbvo7IYiNOH3inUbjC5yFHc8EYM3ETp0A/xOd5ZAAseFt14
T7RmnWtkKdU2QYR8Ljr9jl4hQu7PO6WedtO4Wnn6prk1HmmhIxa29kw7MWTy75bMWCW2d9gLXHSo
OpX+TKZuATvQSv83ppD/zHsWej9+3ZBIfb/C9Bw8vD/veYZxKUiGYyowS4evUFDWQjSB041BcNpo
CQEO4ZaDOm10zHT1bB4l6xH9Fz7IDPBISRmpYvR4Fvs1uDyIq2cd5fHqmHPZmdkC7SFgFPg8XU3J
k7VSvw3Lnkt4cCw99XT2GxlHAyUER+S5cYYZOFs5p+r5JXKsALKkVuGUKqZt4NO9EtRbkkm5lNCD
uPq1eBnJmHefGVdjNsWx2Nisb3EFoFdmmmyhqLdoP0CvKFLZhRsnUmK7b+YLrFWOLvI+78MX5CVb
ZYT7j945TQ079P93ewmvzmognlTWwIcB0gODdKVc48FrlDy854RG52nk47TZR/B8oQGAWxHB0nr7
R85pIsJcDjkZeRSRkNYzaLHVEwL9d9W+3LxDVZqHYroEwGHoE2Wf+0ZVz1Ck7t1WzE4dGAJCg4sk
Wjo+CjMYncfef0dfx1YKmFPZd2IHA52STk4Q8SDRrSLFux2uz3qb1gLhXaZMrf3KiwJfcW6p0gpn
nIY0/FtQMGdKMklt+KWWLjdWLfjpWUY7djz6t7WJx2ZhMNt6zMFZn5/ZdpFn/aEoOUDT1Sdp56M0
cnx94X0HMtCL7Y3P1sJsomXJMUCBm57Uy9zp4YJiy6NBOKAnUalNbrY/t4j5zNUNyVSylXirbFsb
6tj4pYGys242U36SUV4qpOcKBg5DJVC4GG9c+KvFEesS04RgjVOUnFC2XcnmIVPU/oHQeTNWj0KN
yuSeooRi4F8gJ+gM/1kupOx55EqBAPJBfcphP8TISGTe2yf3TxuZ139Jo2teQ4hVehWFJd6JLad3
TPHOjtjYFwYrsG3FqSekRj/cAAWGqiCIvDVRI8NN/2YE3U2CKEMZ7bosrlkSVXR+aPsw00F5aNxZ
Z11aKTv5qeVEgppRrMFepwVZIN9VhKG14apV6KU+YH8Qmv6HdcE2moLsVwrNoTt68+ieRyhyQ0yU
RRmAMBvjVYIgCXd6xo6hgEEbR3WF4hZWLuWRh+MxpRyhld+5z8gH12dyjh5jpAYQhNmNTMDbi7vW
PP05IkHeh2AKqISJifxrtc9+nzXNgxdT6VDQtHh3dn8+FsTyi5/Zfunb3vOdI1qZtAo1gndy/8ZJ
vaVUUybt9lq9giXn1kAneMKSjosP0J2ftMo7TrZXQ0t7Dvu606ce13126MqhXaSgJ+zMSdJmuyHF
hSlJShZhRTbd2oa9ldWPRXcMUGRi8SjodjxheM4O2zMgqnrkpgeSNioNhciJxEy8NZS8hfFtl8U9
HYfoBHSWhy51pQAJm1nASdKNmqxrOCPREMBjE72ELQZZKtIEHbw4M8vOPuGqpI6QOF2eylZbE2C9
9JgRvBgFXJ7GOJnvpON9sGpOwMjcpYI65ilamrMZWTEHFZZYwg+HxGZ4WQoaynJYKHzCxEaIXipI
WL8wks2WjkeQsf59ugdWUe5MdmqLdFvJ3YKoV7uC0InY7t3rExSwdW5htgeMM/WdbTWZvOfhbUf5
dqlrXhsFQN8OG3C+eUm9URZ8NVS9F+KibAlmkJJD+aLuo/BlagdCnTPs6uCnEw1HsyKeg8a8+3SK
n2h89J/C2TjST+yDZPQRp3e8+32f41vQGgcfsUuH1Vn4GivO2OUkr45nvPzrnVA4WPtkAPLAgDn1
XrvTi3AxCQ9ksTIqd5dgh/I7OO/9kzPnQd185S6NL2tuGpllZPYX9SISwaGZPvfvVy8Ek4CGCnSF
nM0bl+1Cnl9l8hHmRHTl7JKrabs41KjNIS/un8AIwS+PknAzmOiPYcyGLvO2qr1AuTy3KY7wIh+W
+1/Bm6DwZPfddiKBWvYfcuDn6Frcc6+sA0gp+IRq53eIEoycAFR9aQrRDXMWK3uN47JuBVX7PVDk
7Iq3bA8BzfY3lPPD/aZy11lne637u3Tol/pdfiYY0rco/eVBf5TgsV66pBwdfbfrXOUn9C0ezUmL
Y53lvUjuiwR5pakKkM4Y8aCa9tiCnSoX8JQTUWPfjhW9G6c47nC7m5KyLObtZll37LkQsWZcSBNe
AJOlB9kN58OvZuuimSBRcvxzQjAoly0LoJgiJ6ffmMfl/f+XTdkGoz8Vo7Ijg+FmFS3PgzWe8lz3
phRCAzimAqIRVcI6mz57pmZJ7KUJ665MCwRoQ95LCduS1W3+kPROwKnDYibMHdwiqQTmct+l08OI
5ikkcFvJ/qGkSGyW3XPUyQt6HRB934wQt4J2KxxEcJFnZvD0/7HZjgkakRLQf+nyQh9ZNw0CzJ6j
LmyVjgTYNs622RYzyQtgXz8sgvqzboY4YRummKeC8Jt2WlrO5QjO8+1qchZcuraD45cpbVE7hZhu
8QIJD+PbHNTXdIUh5HPMSI6Z/qLaexUme7YsAv65/01cID7JQ+YyVjz2khi8BQnhCxE7mtc5RMxd
8kXm3POt9A7mqqKKhpnaPeIJFZ/4Nrus8sv1zLEDXeTSH27iVnfrbdI/90AFj7j4koVkTi+oM+Ub
C0Bomxn2MEQUH8Vdejz4+pa283ZVOyPY24wt5w32ZqYipyrKQOS0R/+cwm3WrgbV/gHbZRgayS8J
0zjmCZdQKDE1kXu0nJZtDHzFuo9ewQLEBjaNVO3yFvcyGmwUk17mxjPy6RFM7+EFukPOtGfrHD8e
Ykc7eQ1zPsjMJ/Zm2zISR1pLat7SUqS1tjmPrgCRUSyQ9NtuSZIKMOMfGqXB2NaEGyGDzaIyVDxk
B2BhyaZ9f06xX9bry19jePMUq7LsuV0oX0AOaf3yXn3vKOi+aRwcys4ldLtqd92js0xoAIxX/MQr
kPxKyUZcrypoU+i4pAVuMA/0DUq1kNy+NbDQgDj26EMv865WEj3LN6cczcyMvtIp5PA7mIB4pYTA
Z/6L8jXYWrX+Y4JRPYhXtTV68Jihkd6qYybUjuqVbXhE1/x/1wdJ5kxxzTFs34csodpLz8zf2zCF
tkOYGhj79EJeO68mYb/RqqqUsaRgmCsQO01SrcEiOAH1KdhsF7+SAlFx2JD+Se5fgxEdnPMOsaKo
1eLFOSrLYWC9PPM6flnSFQhAp/Rgt/yrN20MmxCGHhbAtVNe+eNKKr8v3BdVnptnH0b81sgFAhPT
7jkbmtEMpbjs8xEUKGyK8r8qGUp4EVlOTKJUMacRy+rL4RuwsdtQBs/NTNT5xcj3hpkXdEg18ZXN
jcMjyGRCinftR7jqFvqxK4126YccxMYZZJf25TC8TFlGgTMPArgIuZqsxq93wWBpNBSmx6QumiH2
TvF+szuc6e4NKaKhVTfUpj3jsJ1hKhn1fzCEiAI5i8mz1bPgRJPu97DAJOiZQ3C/DvxlqtCQVVej
npZF1Ts30LHEg1y5HidBwdduZbA+KkD6CBB3Q/rqG7Ec+y98Y/Kqc1cup9wR5SzLhu2NZRPOkPxP
iVWu8pTgZ/7ySHdF2ald4XpI/jwClhxCDabMe1Byo+VH7o9t3eKBYgtc7R6rl7LbBSVGjWU42zMY
FUxyfMFMQU9Grp1LY/wL7yknX1W4CvZu2t2PTmEvYUE/fmvUSgNH4sJOTFo7a/+g5s1eBPo0uDOF
YTXEjny/IU59DKwB5Ur9ujOTdMALVBmr70qCz+bPdCBz7i+zj9Wvq9ykO0WnLGWvqo5UKy3Oeqs0
DOdRU+IspVrEkymKyGjbNSqV8LWN/H5wl9PjeGwb5vxQ7DN7BYEk+e164qDyF0TsH6LkJnDZh4aX
nWPJzu/46VamiaXIKfcvZx7ld7z2g5QEy6kk+dZoYvjsqyCr+tcuYEITgAofTZh569QwLrhOWbtW
7mg8QG5LUy+VJ3ALTnsQNX5uKn2O1/YsU4kC3W0L6QgcccAA69Pkv9h2iPVkg3rMlPilaYuAvcKa
n/9CDmaPz1ZikPysPYwcniE6r/jklAb9dQbHfEa0D2s2XlYMOYMhOxPip+5HV4DzP17phqRkGD57
whAqjbFrRdWN6bo8kHcsyn9WrlRWXkePNzpvo+8KPad3HCfKPUWP2O/Mbgngtpq3F2qBMMraux0z
I1BqXawJk9nQ/08sBjii0XrAIqoqS2CzchdszAYNAYAtmvZ6SNJXQvn4NV/erwpxS31RipBpapXY
wD4J9A7TV+Cp2PsuIFqNAxOUChkoFA+So9Fje+GnTwLc/yv3Ypk1rAwy3pxLuiFZU2TBjB9qpllb
6J//3LNbWeHkxwYei0Nr/OnDx3avIfCu4FDzhKyAPCp4/I47MV9P0UaOBhcpsUjIz3zX2/Tklix/
L5XM7k8Dv8ZI3oDqI2mCkTkL20uSEiVSu4TG8aOyXDOwTPWGPD1Yiz2y0VzsGvuH0y9F3MfR7tl3
gdYV7RR4eyzr/QgKRYw9vZuS1jiQC68D8w+ZWhK3cZr3pXqJMMVLLCPGJPIQ7hWCUebCAKAEj53D
BU6uvoBpRjt6kJwA5QvM/saHweptXH2V0ElD6qUP/6BxxEccinonfm3nHqrXLIeDFV3SOolL8Cp6
v1spddPCqQExn+gNwRYDACSlFvj7qjbdNHcQR87YmtRZ0orWzSnZupOceqEDuuutFGofCLi/hxlF
r7vaP9i1GuplXVgJw3guzQ+GU3Kobqeoutuclz4pmm07VanbZP88+/G8gQ6EReLdBo4Kj5YPaKzQ
xd5KEX72+GuTlZAO08iSX6Ba9TxQBLxJ/JxZ/gs/RhLvpb7XkQJW2AalYuaTudjVsCrDCzJhxetz
c2qEPa6/nLn8s1l0RSFvoPveWhO3h/OabO5wPb5TnhEiD37xvh1z/2DvvzY9gBXkegmidoqqomWo
J04sK5PX/NCt735Q64vmfuXO23KD7jNfVUksFpMIQn342ML1wrZfAgMvmV0dnT3jU0gbLdAwD64C
ipdN83ZJK3N3pQvXJsCamSdXQ0S40vFy+FLTUwramPyAOmg/QY5Je18roR1hsyGGpw8ETjhc0x4K
VJ6kZ0n/pgqAim4KUJV3WwMKUauBM3ZTACVxA+Act7mlG0/1Ssf9PExPwEdgW6EGvN7es39j5E5I
OxJdlTMdOSzeA3HYhs1tCvjA/3QlwXlZLfU8KL0w6BMcqutUaSilnxjw6LUqgdX5B/qVaqn1BYkT
6i78QIBRjiiPNaw7c6IO89Vigz/8wqNggVQsRmfoBONgo/enHPx/KJvIsCHfISzwp9lUJvPdjJS1
X7BQrbuXo0Ohfhujr1UDj+SjZa6rqbYfdiQ/TTkQQasV26Iohy0gBjZlj9LJjMm58TbzDFUtlLob
W0wd6osKoHz7WDu9O2udBdB/goPvDYYNRtlebF3MuD88OrPk3xScuLyTcH9r69Qd1iPfTvg1OObD
wU73qH1iDI265GjuLXPM4xaNGjXvYU1O5qG88p+72yQToZxSlBDSkKxgkLjx1RkzqWg3gFfnbXPh
s7CVEx7NMEVBKle+0z9a/gNjj2ioQjNnAO3y27lRzlt2fXtLol6yJ84dtFzLllXUU6tIe0KhoJyb
Rzqi2p1gOM7tNO1gcIiHB3thwsRouy8e+2EIwtaUsmv1GTXt45ZuVSHH0NA8/puEGWvCtkpcuaTg
qBtKcu0Y6K0kpHJo9heH1njm878SeZ0XevJNdRhW9exWiP5vECQy6gt6wohQDHJ38rGZAEjeM7t1
wZUJpUvA5DAUrZv30tSCJ5eY7/axKqNeQcqUNfYk/ZkXc5uJMPqxSdYjE5PgUuUMqi/wAOC5ntWY
mknC+b+0wwy0jHtwfKSB9+8bNY6E+drJEWDRv06tknkmS9ZzUrchCOXZBvF6Cn7CIrKZNP8fazDO
TPoCUtalMdR/lNarSF4Xp7w4lMuFHC58BPJUAxXKS7I9GVtysUMdrmDPGYjRS46PLvJGAA77Kt9p
auUWIij3e/q1JXsN47StyLXMml4K6KRiRJsL0MU9OtqgQPFV5usSAD3AQuv/ETJkXfePmtM67lZv
Vrohb3/oFBN6oWwlT/tNEzJUGxUkzdTQIaoZWFGcW/bkBQ+06TsD9DSOoHVTpooinwo/+s4LC5yS
fqnHCGP8qzmgEIELdOZWAD1nKFv+SZat2NoXbqzcvbfOpBJusanod0r/KOuQyN4aTtCsr7fyLuAj
i7uLG/R3mjzPtEISXFDLeMRgpL6C+2dHyczTFcOx6wADOMRz6MEm4ddbiYobnxx/ckuWOP0SKrt0
nWCOL/ErOOcRXHwv4bjcPw35BfJrd2P1z3GhM82nxPe2CC2tuLdEvlWbWEMQWqqZsK8XM3OUadbb
YFaEJENVW7LBPfNycW1whV7AUX3xPYZSMAMhgmQLRMPlSXPzyR8IXLpurKzdODwdOpZWcG4r/e/z
9XK/82B91dprkHXKIUChyn9mrSJdcgYH1upES+LAc3eaH45yy4WhNHfMn2Fyqv2X59OAMivTGIhv
oz3ufypzUTc9eLr+kTs5X1okNmjZLcoNzBsmdAFP+1FDwXNkKesoaH8kgeH54PmfKeJ6BKyT2D5g
3LPlbIdL9CY9jm19LGsPwo/AG6mtXtT8EP8noH/SCOfXbe3kmZIioNjpGVgPl7KkBfrfpbi4MhE4
VvHrcWGg2ihypSSDJgmFGdrBdmd05WYiMuRLTL9GNBmW7/DUiFkDV10aPRcHqkF0pCKdGFTAEz83
GHJy8hAJyji2Nztf/ACC0VydHz6ldP72QCnGAr7oTqpkPGBKHPfd9R8kz1FtU3HA1VoesDlvWkrd
X/NfJdJ9wv4mJqS1MJs5KBetg5gxFYE/SeEF/TkQP4OAUwVmJGvcBkSkiF/SihKXT79xup6rJpES
+5FQs3jdpG4KlwPB7aRQXKV77I1NVw7xGU7lzrVDKwNnz39FcRGMHnG6PthiB4AdrDqoGwk8JOc6
uRuaOVOBZzAncAuBb7f/sllx//pYMOssRBzvE959yJNePST3fwfqQ4idVjtjEg+o1tIR7vCJ2nnP
0tHtYlj8F0F1ebFyRmhr5TkUTiOrlraKEwG/gwEs4wo1vTKgLIQ1Lrg9Ot0k90UEQbVN9lfvbmPs
3EPxOIT6zxqHmVVUNuK0VuqpKEhfz+Ey+moMU6lnv2bBMl9FOxVSeEhx6LnKEjeWqHB1InqsXtIh
5Zr0bOAVZ3K1mtlZnz89NS9iXfz88cbENLloTXRMJemV5jry04BCpEP2pg79V0WLWOmrN3JxRlQ8
1ECb8cRBANGpHxvTGipmOhbuo6ZWxcaQmMjOddgBrX4MMvyOg9/AJZwCuzT7mxuh2df/fCGZ5cEK
QpRX1DE/lvejAA3dhXgS+iGcput1fZbL2JVKZe7+OHol30oiAXHrdomXZjoCGBc4lv0YXevqC4Sc
/dIdYIl0HlXMBQZwAbj9iIxGHzkPG3uxBF+vSxVLoVxRAMbRDWmlJ0HOND/bn0z4nhJVQP/3YY9F
NNkWzYFfLDdWLgICAplTCRJBHMyHzrrZz+I1TUXYHe///a+vCcF1dCDBDxBpUTp5Ve67e5OuX7yF
MX8T8n3U6zQJtUoHsmhV8ScLzX9YZT+sb6/L40jEuesdVYJmtca8K4jwNoywbOOTLcBsrsquAIRo
AsqQ8nbveHXQMrBMJN6l8RgbFg1fs+Ju2ng+mhSHCGB+RrYQI+c6h/fh6mlnKFTbYbUJu+AvIBr5
URtf6sOQBYZvSUrniaDlVnj7tkXhbb5opLpZeYXEFZk7th+CxQWVzqX491Q4GBTuyjdisNDd/tOW
nvK+oa5HUI6fN5SWhmgAnsHgc1nYzGdM7gQy3d2QlSJITs7dB3y8OSlP69qXb3vcLpzUvUfZDirx
PVMV3ffL/ZG78bm5d6AUQ3ftSgRvbBBkNmJeJhflWIvppq5AtlG0+whRIpNu03zN6xr7go/zjKT1
VqnzStYDjAXW1mL9KCJQhDcIsuDNjunor/4Pmi9hgUwumDk8HqJ6Vhmh/0TOYk6ioDlt5yXTTAbY
tFSio901q5WP64oHQ6xLUioNOu9P5WW9ZTGJqHrc3FvJBgBxO/jCpxa2Mw+4uG5SPEcq2100URvl
oG6aulSlusS/UTfyBwrbWgqVaK+sPQQz5Vck/ksv1mfdeOLwr55yrMARNePrfARXuRRZrDPmccOO
nNWf0vd93/t5OfzGOz4mx/40VlP7SL8zmkQ++QmaVMJ0i+hxeaKHKREON4hkVAQpmgRKVTbPE3A8
W2RBSFC3MeRC0+craUL2jR1POexX/G5gvBrA6Jy9dJDF/Wjpiz//rqQrrPYzTsBY6GBAVe+3st0H
a+iGAOggEnfjNK61Dasoynj0OeezFSS8WAPbbi+a12t6N0bC76eIuKM17Sm0qATAJkF6dKM0ESiW
GTqTPhxn+GQu+kWYI5gnFiP/L9pnnkZw/yLLy2BzA2oaD5f5vSGjQJL1RFipviFQuzJb6nVtLS0x
NNssgNqHyc1tEeZvraAKJ1NYhxwcU0tYfF1nuoRAKwKmG3P8c6NTIf/HZtrZ+3/OMYP9Bc7lUrMT
Og5Xs06rMIXLH9Uyi3oyujc8EuJyAaPB9Pxg1Oz/KevALFjtwx3KyS9VZd7tAvQcNH49b6O983wq
WtZef6fxjv7p2iKdoAoYvUKS+l+348tslmEK0Mplf0/9rA3HU7DCtUAFndZtGlhPhepvPY5QTG6g
ronxpalEMtYUeKypG/z5Kw+W+VHv4GTXB4lFG7DYwCKoa1YXmwhfGc9Fkh6ULXp/elKHuQL3zv04
85GeCjmbA9XQBXCLUYdmcXCFeZ8qx043GU+sLhQhJx4J9buW9EyGQ0duD8CUvEEYzAIsxq2GB9NO
Jahv+WbHwJHN2Jzha+8ZlcgCxGX5trCFb5Ns2ascRp1ceFynBVf5XDJu5nSeaInUCk65UCccfDgC
bN248uIKQtsSotirpj8P2jqL2hSZ3JXrkyg+2K5R6CqyMX4r6tsa4DuO05qNlLyoqwSzh7K8pNSh
oNMoEG+j/HopmVHi2O+1iF01zrezn8yn1pLL2RzbLEtU4QtB1uHUsrLOsk58RwJRwul8k1o1sF2T
olouOmXJoZ6geIh1Y+ponIIXttPDR1YTBmHUvTbil6hXivucpNrB72hrvNVNTGmeGLXa9pQ5smM3
EBruRyFlBeiuBIHfgxfWKEBbuTi/a+A8/tg5UnsIMr481EBG8xAJNmswF7D6SsT4S8d7Yuc3Y2ic
2ZTGx0q47fDnopL659UGL9h8LejfpvIixTAWuuBeKnjbaknCJdOp1Nn8Pbe31L5533xnmhEwA/TN
1WoF8j9Xwjml46/RemlyCEmt/+wmH/VLqeb+hTk4p6XIGvJnqh3RwcyL8gv4IZ032XHQ7KLllGH1
Bfkj145ge9Rd4/dhboEhy3lP9hoXLg6k+Q8w/llGDpKqr4JWWrTBcF+RAKfC2QNJGvzCJxfPXiwL
VBdur6hs93i62yIxiAyoV1OdmtHvsYHFxZFuVqkhzfvfEEB7nIrRPtMwlEn4iuUIhS3Xq3s7KUlV
zyE0vh1vFoenrssqLXp/jA+ZibdO+hAtaQCvSIMKrUl0AmLlzzKXq97wPUuBclhIem2aPZIkW2GG
rUdrWpBxNiLPperf4TtMhMSPu76etwj1k2vlxCl64wfQX1EuaE+Ev19lwGh6JuCUcXFeOeUB7HiO
MW8Mn8QcIIv93hwE0KyAKAbFxZD4LVgDtkJs1c00ctMq7PyCuFvdIeL8diHCV+tVavcMs8Vyfz2f
CTJH8opfHiAWWeUeDGKsO0L8V0VeJ10pnk8lYM4mS5ufnSc9KdfM9hDL5i30QrKMA0D1aowgeahC
LedBXpSuUTVaix1qa+tZCQLSrVu8CbhXK3SAtUfFCwcNvZ3jrp48YvCnv1yqwtmD7YE=
`pragma protect end_protected
