`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 24688)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQElds9yIbLvJzi52IPmE3e+JRN2
1dGI+PWA25fjnwovZmrXRUliArqhyqn95sw2xPQSD8kSkLXpEy1HEI9BvKxRDtQMgdBCaLMHKBU8
HdFeakF721+RBzKOZKA8M1kHcRv/mK5eZQW/YC7pOlOLBNE22I2Fh57uLeiu47OQ5fiN8ItYwmEq
r7FQeS+Q4+OkmhHymM/5Ecnj7bzoTJXHGUWM2MQe2vqGW3WwP5D+R09QLKb7eCOi9yXRaHYjnUyX
hbCj58Xsyf7GQxu9rvy9s0WVJFaLYd3/Rmrpb1CCXkEYp+YltADXj3TA3MYZ4/jgykUp7Kaeq04Q
VpOPskJlxTD6cwXLmyv0yrVcYTwy/NVkOJM1HmYYIpW9UtHiwAIBQM4XNJWvTgLaE6mEbDnrm5pg
y7oTbtQQAyXYD0EOulBtISYKtkodNkXWww3wGTFTAaaLBZTGzodhCfr22wlK+DLFn0WjAfLosB3p
ShdTtjH2mvwAO2dw9ZGKyb8tPpYAk7dW0iRbDd2FcLGmGW4f2odLx3H3Fi1K1XoCHk2oBAeMCrKA
0U/LJYL5Xv/z/tCb5/XOKguudYC5JN75r8OjgxTO9XGR9olsNwWn0M7iFxjvAtRE2ygHr+kfQoIE
1+lasISoGq/zb5uNEoN2J+tCYlT0jnrfoiMEM1Qe/q2kwXoacx8UgGOKnjs98HC6f4ZoQCI5n6ZA
CqVqRbpfrsQwCHYVCMnh9HW7DrVWEJpZ4tJ+pXKzNRP3ffB2Dui/w7BFkyKemX6RFaDxnt76L1Dx
YOhCnCfffnX2aEjD6fba5PT0K68poAazgBkj8puic5jhPWSZVWHjAZoZPsGAYhsI0Ds9yqMRaxaT
nfc9Z44wuA/TDS96CKAPA58BXxOc59qmPdeBGtZCjgKP3f6alHutbOG0Vsx4FhT2RZH2E8hMGswM
ODXJTPzpCIFUM8hbf5Qi7LtJiWJI3iVGFBZvHKqxdH3J+R1+ej4i7JCoqJtxJfrUZvXa8sIW9de/
OpT2HX02cJdt0/Bqu0VIosOAFo37th4gBC9Mso7f7MZmBK/X6MuAb6V+Zu6IpI4Lystziys8/ATL
9TNYqi9yB3usQe9Npry/tA87sCrIWfypCYhfhI4V9hyh40NOzYMVSTrIatK32/PjdmtjcIgNDqmu
ew7Si3wy4Wlgeth/xgdFJ2YJ2JCmfhrsj1RxlNIBuYuvZpjRlRUVGAmSg+lqolP7BsO51U1r8Nw0
ZYBS4eFro31SXOhFBg6Vjky9z9RiWAqgtznrRD5Sde6+S3O942XySBRJN/Et9nw3MttAWi1h76nw
TAJUC2Blj87g/h82JA4wAy37WZ67zfXtzl1RAJnUCq5q4t6NzPF1nOmGJkm1LpdgCzQRchpFmfqE
pfnR8vNOk+l/D808tdS39F3Js0rOF/WXLGFCKylHAmTtAwc6lqDQZwrD8/46vT2Zkjz8V2JGLggR
dVGq0HCdWjYCl8Ish4ARJrKCHG8yurWJw4G/f3LMgTy9DdWvfeQ+ZjtXMaCFVQdblKP50KnczZxf
9JEa1on6QWrniigosZVxIe9yfvP6qWEhUTuVJ8eYFbMR9ndW1rtSls76Hb78pl283akK7lmApK2t
HCGmZE5e0/5V/VI87cWRme82+VtknORAvL+wcaX3Q5QDQnp3VVdcrmw0Ml+LB16JmzUXG3RgmwPl
oZZ2AK6iTwGoPOqX6Ghoxk49lxNBS7JK8o0ScoNzC97MyNi7BzzF/d3eDreOkaLan+l/nefoVEj/
DMoVjuTl3DwH1LO10ETvuCB1mhGirIMgYRS4DJuLmLAmCpNJQSA+VyhNYb4RxvObwDBZbT/0pChU
clJeDeWMN8Y1uGV4mE57AlTbpPVj3BMWDtuuOyCxQdkYMoG1jxYJUbcJeBWtCRXl+VuEuBvCViVt
WQ4mte+fUUe3ef46ybvWtZykwNen9ALGUVTZLApFkZva68Ap5vnBAXLAHPkaA809h40B65ZaaSfT
diLioJOJQiRynNMraC5NCoxuUJsfxNjXyRCNwZ0SWTFuW3J2K39WawmSAvT7fUFinmVwPHSy1k0D
C3LGG1xF/jekcnosKk2PA1wdfhPGbuoX8jdrEnTqKVIWP3G9J/mcHvaLaFL8nTFgVxuTFzanGs/r
lpgne7WG+ZIf9R7Y86oyPC+s+zBIPRkvN63M3ifhfHdzeK7JuROpNHyR0tlTn+qoE318ODUIJkT0
Ga+OUwQ8h9l0G8EACkSacrIcE+GCJUf1BFe8pBLCouzJ6aNHSzUd3il/sfmP3AkNZrkCIGsmD4fT
ViKZ9kRDdaW4TNc5lPE/z2eUywdJDWthmKaNTwxk0lURhfq/aF4Lb6R7jzqh7lFX3Pc0G6NXzXGe
WJb2AZSTzdnZOcJWqL1R6u30vLsUzD32JCMxn7UH96TKv/rbc7+dRsxvKrJalUhbWnhzkngttQp2
NK1jy5EwR+qtyGOKEp/sJ9rVPnNh7ekOex6ADMQ2BqseCxwcl6uprNlXsGmIJ/yAmDgrUZWUZ9Tq
hNfPjcaK6bWa8fDXL+YSfDBZgx26gyryTOxGODq6cVxLRSz5yEutcKNWYfD5/i2mh8C5cY0tEivv
WoYIPQsmWdtMkm8ibNhTzaOdgJJNUyRR7GxiEvqXbmxUQ2HwEK2tW/G7k9lHVauH4Ky5tGXzVr/7
scoceFKc0ykqU/Z8z2pKZSfD/u0tjM3SyvyGej05lOmWhjxr1m2f3Cj5hqjPzRV506D01eLWHDNG
C2OS/okiNLzqTZGEHBVRQQ+1I6auOje5ulZ/xwLUnFTOXGWgzIXesWA3NQyW7OMILzSIpL0RaEBY
lhfoDZxXDPvg9h8FRHyNEXOFAKXDzhSfhVzLsiumIh2uX1jhS5NWE4XEMkY9aQ6Zrxd74bKNKTEK
6sK/NEBR92cegxIy0lLBLRzbm6saM1VSfdfs9joCCKIt37sR4T2SdHxMDTsTxN5NYTZGKlqk3i5X
ozb8cJDf80Tf4maHBQj2F/VKk/atEm0tcvd0z3EFdA1jt6SkrtrxWgFpzsBLfecBB4JNs9nLanI1
YEuNrR25LO9dxeIi31Qx1WkJbhp9MMIrZvtatwLaaHvWl6aG903u+qHh4a4Oz0GqzbgwnAiq8vsn
Lni3NrlQiepzhs84p5/74tngvqbhj6Z5Mzx4WYllZk28wC4MM/i7WpFLUd9dEYPmenRKnktUTLnP
mN3/vpes/PHQH2DVb1vyeoLFVCa6L+kvrady8jNqg2MSRGZflv9b0yKi9zAk2GMZ2iW2qNdys9X7
LoJI0slx3+kBed+1Ax3RODUtTbtp6OpdkZeUgxnsImLV72Yli4Bpz0waL2eRLkxLl6RWEFOCDMqR
l4DkdjPreyx0MVm42+pWrV3zUsHuzOZQ6wp09xSCvXqygGw3BObSMIN+mWEMtDddQO71FExp48o1
pKJF9FuLrI2Lwqdgt8hxVEO3JeCzgoJU7WZpVwkG/7/7v/Llod8AjjalM9kjlmx4FFm4mGoZQSha
RQ8nl/s8ilUALUOy5krL+dmBA1yR3EX6bz5LnYd7ZKynXiihA676ulVS2vKrzC5ht3/qqkExiIZB
kXZnoNISYrjFXi5kYGZYCy5k5ifvNVBjPHrLsYpDw943NONAVTPAKu8txWoq40WyFfd4tywDdKR7
x/9lHFfQU4JkJwqiLcE1OGx08hY/XQzKjXV1RBvcUm3+AkcwZ7B1FYRqCMKfanPFe8O+xYiIJC13
zFlX4jPub5T3eGRqD4NSQSFoT7WYyVmiWGShlVbBz52wpqfrqbEqM+6KgUvmI3uPsyJn8mg3Q76G
nRRR203gdvit+jOPeLNb/VeP1oba0jthE/zVLCawv3dTxBgqJiuWMr3VgDAu8XRJMs/CuLotYHoF
VPxDO1arGwXq+CGLNq2fRqVZJSY11XEP3FGJJ/kD4zu+NCCkHKy+2bqagEWs90bJokwvbWGNFk8D
3mjMevzdVAhBWmSh4R1AelQzrVkv4aWZKkD76zia1wAF04GTkoHl/lE9Q83dSolKFFNOKost8MjL
5DQSNuwt2+2MCVbtSxg4WFGkgOGunxe4+YcF8JrzwbD2Ss3G84qIjytF3zKDBX38advHX2PsRT9z
GlT4IJRULu6j/aJYOAJ/vrSBJzsAPG/YedLfX82I4syfRWd4iUR2JUmPYf5gP8+HYtCIJibpMtHk
wvMMwnuPneliRuYRCvPpTFDwDgdXTYRIxkJXn1oa0vOff4lnPssm8w+3jbbfY8k42QbQeeXZmVfv
WECYQa+EBk29e4GlMITJOgNimBqj0tQd3QkceLlZgaTSZ9u1s6l2gAnW7+elM3xsXMmInx+8+DkR
0gLHXuQasnazZIMGflDlvFxchz3RftFLGGvKUnu75PwzqZyiRly6wC6AGZQ7fgRlsg9TdAGBjf0O
UaKp06tMaA3DgimGR++dhZVunTNxCRXprIZfe1cbCEydPOrk/WL5TKEb+VL/tGcP9f6gW8qirdrE
0/w2R4ML+0WpO42dlXIvXziVMy1dnyNhUOmrLx9h/+7c2pNqyh/CkZUR3TyZyVG0ffJUJ7N0Z6ev
qBjtko7Uf0jsnP1aFysJC1wL93pDFQvSGzn43wKbEQ/Li5BmTcDFmqTbrhhDZDMG0Ri7j9/PYhT4
jS3m2FjDQh59VgYx5AMxtFVc9kJgQP7VPiviau+ibJhSgXMLEs/J+hlGVuUddUKM5Sm76UKvxiKw
NTfojRu4vI9u9Q3B1AZgNz2aS1/usz1zupGj88UX4EZc1Yr6pUINX86IXh0ixWcmLsRh4enj/7Kr
CSyfXMVnGql42RXzdTQnEIC0ruOvXIqDsWmOytEAKZ3XRpE6GSspu44c6WavqkQAEtUqvcHJ0UGC
Pj8d6K20Ijtf1uiTzo6ARlO8bvA1StaGqvFcUOzW6X9zz1lGnIZMrZz/HjhmRPL08ROSUf7g7dEs
tWyaNqYL18qaWWh/tQ6kJ3er3bNAr5lCHYHsI2zEXppreHYfhS1gyWN9yUJyaOriwCk2GhC7Gj0m
Vgno5JudiqreQGZFt/wgD+feEPpCchpGhXekXZNpyf3/pIfXAzph/VbeVQS4bUNAT1hmFUkHTMdM
z9cz0XR+R+bQYFP9W7Tz60f1JajUFPDh54Gqae6dVSkG3F3cN93ojOxTRpwHxgt0sMB8/DrpF9Tl
g9Nl0FVy+rdDUVB76PAZcSOs/xHaBazvUvLZXKIdsFnJmp+1amfiWNMc5DoduxWJ6uBjZo8x8DP+
Yo0DbUMKIWHc36l7wIAFpHgs7/gTb+cLENIlUoj0qkqrWQoEUPcVNoqh/HHrAHQ8Vdv8ABuAd5Ud
uqQNOVoCPtEAE7FzQvq6yD1o+e4wMPa4PaiQaLI8yeWVCapv4XPUoy2m8SoNjr/tTLo7FefNaxJn
/PY71HGpesPYmH86xgGYhBj06g5SimYckTCKcNgRW3TtuZ0ylgVsATJC1cqAMoD/wngsNH2qMFn4
vnavo5/BXkXcKawDlgWYM5xAz+xm/2x+1EYv0qlIxqOpG9OdVEE+lhpgW6+DD8K+qCBRWDX6VP4b
538HcYQq3yWWLBBQGga1351YV53qr8o9cLFFx6QXfdcwKi7Z1wXy9UQgzeII2TTvfQBf01VeSMkk
mMXWhUaWYnG7q4PL69QS6+TMJ1d29rDRVNBEDzPHznVaJfiPp97MDxlEh+ycEW/8KrxzCU736i99
/iPUksRzkFmeBKg0goe1Wrz7laiseGJ3eBF/Dm2JseAFrs1nTFwt07LRI+XUM1Xe8oMH48fBPIR0
ibNh3H78NeU8qIgJFolAcLNegHV2/P6WetBWJd190ajljsfVJKVGRIwnBxWOmSxf1DlGUsQDbmlq
i7po19dA5ypAddb83MsaIUAqVFglKYUif5rx+GUipx48ZSz+SdhHBQkZn8zL9pgBF0DjtDS4lb+2
zxeV6kbjV9Ck/ifBNmxdpVLKzxHTvORxbzqE9tWHRlz5TCiiuf/b8JmsAFaFC3l84dxeG2wWYHe3
LOH4bArC8KKT8wGNJUdbIO5Ay8hDuPn3bFwkV/SF1Bxgh+yqs2ZGTt0uoEaOkzTsr/JLNA/F9/3S
fyrrpasp2wmYtJtiQMPptboPWDSrCuF1ei3GYBuA9NtIqpKLysOLUhIL5XL3IFe6o8vRv2TdQniE
xXqPR9cTJ0aBkog7IC68E8GA4w9SXfSxAYgetU6pMMNrQyptt3QyK39JZm1YorxjtpvOaDxWv6W3
07gJfR5g/R49VxBf2VH7UE54XIqUDGaTDdvt9YvmNQCeazlYwM9Eme/garsvPuoDbrmvHV0Eyq2Z
i8CzvOli4LZ5WqvzD54ovd0TtDUGfTHW/0oxFOqnTBbja9tPCtdXstFA2xF7ACfhWE1IQfo9QFp5
Y+7UnRjkBHFiq9NFdLxgOjHs8ER7hZrNFM3lQq25Nmq1Ttiryowb7OU6jdH5M5hFigbwmJRU8h7C
4KKGMlCdfYc2j8AHRRokUWMiTdJu0PIgWBDwcB0AlPORwVgy/QoPlRZ7RqRZTDS05x78GMJ+QA4q
poDrWKBzVW+FZXhFo56d+rurJoDVaWOKb38hTxz3m1nMGrFhETfpbWjoABPi+74R6Z3wSlsfLv4U
apZRfyY5iKAmF0ts9l/LrnqYLIYYX08mgwWduxu1gj6GIvTaK4DNg+AoMh8HzhH0WRnybxkiGGfl
bL8/0nC3R8ypfGGhxvXS6aSvEKsmRFl+AthA7HxyouH7CKQsFfQiWto7xvIijXkHBC9OXhRMHia1
iWTQRS0h2cL5s4f75a5NArkYcC4tH52hKF7qcY9aiT0tqCfygW1ietQwxLm6mSoz3FTJ+6Xvx+7N
PELQpovTlQ30ZuKtFUo+kN6o5QmyV/2A+irrILn2cM8mO6/MMwrx/jcN2kGYOV74966u1PpjS9cb
FKmhSPWuZDU18k7ghML10cGnmU683di+ICYhJ/Lbgm9HMQVjeMUJheE59CjFscGvoEQlB6oTfUJo
3n1egG1JW359Sf9xdrlV77AfSfM1j/RSqi+LtaRmHCm7XMCJ/rFLi7QxdnAdMPiVpRdKoiF/+drt
TP52FMNROn1Mq94wDSoRBZ/q0bevJB7L6gLXoUAKC1Gx5Z5mr4xrX/u8BUvXQpmBGzP72TtFMksY
RluzIHfh85WRz70oVUhtjWqVTB6SIGriHynro1ipQ8bhol4p9bdERITaBavTT6haWSXB4SGIUSEQ
GbamicOlNykqZVVfd8pv80/x1H8RoEGf5dl/GgFRNsJviEFepTCkksqTEe6ssJVE2pLL/crkkzmT
3kmsFIpfJUoI+8u/S4eIwOrzLaGemJerOr0JhJgD39+IncKnnapesX0fxyJYsZBwRIXSXY5vNVLv
G5inTp2zxhb0J08szPfruDa0hgMzn0N1zlEQb5e8+G+nY3Rg3L6lBe/7vFOIrHszHE38cq0s9jt8
C8yijeLW//oOhw50wWuzxOWrSv3sbKhvQBFvi3uGh5o0K1Y9oqJ9eB1UEdM+Bb25zf5H/ahrDi3V
ar/nmcsG3SI6Pi6GV1Lptm75oErIYuRkfNlL/p28IThuRI1ahNuenf5e4NBbL4s4Zr+BiN6WDSk9
G+ueoAVmDBn8+LyiVlOMpDrzvjBbfHkRwqwlii0BPV8RZOhy5YcNqhe6dvsmmw5b2c1cB/GuPxWy
Vn8zGikC42NqkLy+jfGlyQq7c6Uh9t9RC0/pWIC9eNLu+mBAnQ6Hazvz4vcnnU0ZQLlBrgAMe73J
5xNQ7DxSruaY6qEmdYkEZO8t4IPL7uEFon9LglQzxUVI1b+utbFWVYU96hp9uTLd7Af6b2MqQgfj
vqMMhmyt44qE/ik04D8qLdn09Jc7h6p4USzsCwGv5A5JpTblCmw6oAWsT5nP/Xb8y5ZLionGbsm1
phOggF2xmm92trH4I9/zDZTNMv9a9aE6oUeXcltkNFszJ+yCyk1o4iovsVq+ayOMPKh/dvTK1It8
mGSwIAJDssAVSOMWGXWkKipLyWyOKF+RJEy7Raq1nlzulg4UDeibEzz4V6vB9DEUes4/g/RlfUof
ZHnsimYcjwIJNiXFzXRD8MwgcNHZcLByH498Q0VSePLKlDaYmZTcOwzq3GWwOVravPb3SO/otEJb
aBnPDiAUFN6z3mwyg1jfQoSqGEG++2SO5hl1h4TREtvx+FChrp4UUaLlWLee8Rspi3h5MKnVIOO0
ewXzFX+B/ARz2liIr4DjMATg9ftXQJxdSJaoCc7lqCzOumZY6tkR5kMQO13aS52ZgFsaUwgeKQyM
pvFMapbXNU6GWk2ufJBwCEJVIu0p8a+PTGVEFU6ocK8OATQe0c9jnN27llSKOR7IATDRmdCu5I4g
s2R+AAfDpN2gkp/nDp02boTMZ8dBzdeNgZ+aB6LrLQC4IakyslaSB1mYhKuFt5iCqwPShnOzAz0z
QmB0bD0/gNbhNbSxRWgRHc1bVE0VMcjwPc/UVLJ61WX/O6+lv4a3kW5rRPtWrnZYF3EdQ9R71gyi
I8ZTlLfk5BF1t291NNaDz9t96P3uOP4kXif2seY1/7bVlCSndOj3hynOtHL/eGESxieQnhRrsPzs
VK4INz7w4evDnqj+3WY4SWJT50xAK8YrQtkMe8+zsiexgi73CI2QMASFJ4oWFnChDZvKHJSrQ23z
jKOV3jR0ijJtMP7lsCKh0kLGCLeicyD3i7y8HIur52jZXr1JCmlmSFJLRwLzLSpX2B+uhsXXM/5R
TofFz5g4Hg8pkiZ36uWGimfPtvMxuSrknX37mkAHX6wNJyRODjSmvjqXC3cAn77y12iKjFtvH/jz
bRjC52JWO8qjrWWgOKt4zokqCvC/zrXw+HiYD3giYzIzKiwT+BUftblZ9/iQxrdlL8swa7V16Jpo
PfdWEwVsyhrK8AnKTse0tb/HAfxyxj5hzJ1P3HJEBnviGrEWNhDbOXm+SXAXDqNRw9+iy6mtTqmO
BAUllvyHY7irfUGuh8vpNo8/R/F1KfMQMfdE5xT3STlkPXwl++q+VuGyP45pqv9Q0S+Iiwz+sV11
sIIwQy0/IlsKG51zucxSEXplFOjstgcpNEMwLrc7qHI24zUc5psLPDioV/ZQBvJPytk3wYuo+v1c
iFaVbtJGpyuyIKyWVfUworsx6MXNylE+K+gCnSnHS+M/cMSjXQsrWystl5g4H+c8VbFfDQfsy3xP
kHYWiC+/7yEqN2u+FeRkL05Jj7WBJ+PNP+Xmgq5QApwox9JeG3jDqL1SzQ9GNgEoBU/ssodzz0ub
GSAloTej35SYaenZ6apkC1FfCGD0AWA6wXBaTW6XIFueJWC5PznOGI6AvfKBC5TZElazU+5XGlFB
Gzb+agSAAwnpAswFI/w1NSdO/ercg/jItEc8FBCxe4BBMn89VK8CE541TwBwD3WjxM8uGp5Y9TZV
XRZXQl6pDH/3rULr4SJ97zNP/NcpGEcLeUG+cXG0PIvKoC6lQR2Ckn9HvGzpRsIlp+7+DJsuvv4y
om/CvYpfwttfncVbuqdLN34bE67MHNvkhGSXP/Br5Hg55eESy0tA+zNNcITSeUJg52k1OyoXRUjk
5zNIatcwm4UF3AD8YPkH4nsBF9WhBD2tWzmrIuXPmVd0JN9+sG0sASaDhz/wFiOXLuHBAK+mTr0f
0SOW2CRRD2q6hAg+9St5RXmwXtwX42CKzc6KKCYTeR4jT6DxBesrUgZsRxW1rqQLcW83XDS1k022
ccp9b13Ex765zXdFsETb3+Cz07OItyPFAjifTVyt0D5gOQheTuFANLrCYo7DZquyYoTieyi1y8Mz
sbr+73ywJPubx9gHLgNe/6u5XdVmVFHlZCDTRgltagK2tpNzAkM2riClCef3gk1LH+BUyJ2hWi1c
mSlUTbu+02JsB01SNbtvuw5I9lY1lEd5lFh1BbvH4wK0sU8X1yc4A54Px8a9HHUWLSbAkFLS/Cuy
888/vpncGW4jsmvHjJCAR9DHf0ZWiayzn6WJBA6dzA7O2WJP5wW6NIQ4ZEj1GbIXNyrm5xswVq+j
IY+7D7I0bDj1j0IiVvP1s1tC9XL49d+4z5/PaTSRcSBlpR69Yv/lEwkUL83t5ZQyxBNyz15mlP7q
mWLejVA9v6wa+hljGA8LyAJv+vukMPOMod5Go5kMJjmBvLw1sNQp3KEkp/6cE+ZnxyWjr6TZbJTk
kq2sowJVYWHzIO7Tm2Q44geO+CXd2DHwB0a/NSrarSM4BoDEvtdxuxm9xvUuZPNHFWs3tDz9sS7t
rHHOOf0JAIsGP3iQEu3VpGQQR7WdpdJWMrYrvE2tvI8Pv6RQj4aPUDZsf61oELZbYohZLorI5eEN
HW/XENSFG3ANPpd5dg2XtnVaLqH6MdhHTLjgtCiGOx/ICuHVeoSPjs4Kl6Wuvbh0GUOAVZv7IiE9
9Ec78kWcSWxC8Qi5YotUhATSrLiLlcn+9gNDQHZk4A82AWJ9/FG3czfmQsqGBUlVfXbb5ZmLgQHL
G6CUFT2iSTZUCDDLGxCB1i1tjlGaIU4N3BHV//7PjKU4mcUsvvUMJtdpX6KagdR5j+JSyWqPLeBN
hQFkztpiGcs0b9Y3JAM/t5feIWYqvTNvMYIWQ4heqSCJlDvNbBvhJkmELwKhz5ZZaUcg8MkcgJ3N
zdzgClNBHZFdktYFzyW3CQd2KFNB4a7sEtejTCwPf+/JqbpoeGHRt4Ks8tcjpog54oDSD2xWBD7q
iTTvfwoFGRvxgap5KG8ESi05L7xgtQ1alVcdYB7sRylCuP0oH4r9285UJ4XtG1pA1Y1miyYPDY8p
LSNPHRaNegXMUx7jhTbvmWDqQBuR1bTfFZoXXsPs7jUh/tH0bZXn/9qc7Iw/znd3A9qbmYp6fGUH
PoK5FvtS4MJK01dwdKjFB3hCzr3Jv/su3OpF9FU4GKCGb81Dyb1KBwcVy42umdF1PBS6tCyZwxRM
Qa8o94CQ+9oaL/9UqTzxodayKRqdX6eblx9SXwdQatjC3qKQxOta13ENLCSvfhgFHdE7Bm7FHK6w
LhuFZOB6jLGPl9hA7oHscAyIXaP4hukAsJnHNxLkfNUUlJolXD3WJR+rtpx7EgoP9HebzIo8OBR+
OogSeD0mNM8JdQA+Q6gK6R8acZMXyUtBjjZY9A3wPXa/H+9+gS4drP7IBg6w6QjlepjoYRi+Yty2
UIvU1IuLZnZjA3yPHGv6Nbcgz4bH1K5IhwZw/NIwRtJnwPpHEHxdjS0IWAsGMoBM8aS5DoxFJ5sz
dHSp/8bJi7G/fc8wGoSyx91sxJ5tbnIiTGGiI1AUsUzAJN/2IhPtS6Kvp98uJhfKuSsNHgGtbrd9
gja8gC+ueVx1XyHIE0q8IJcTlcTUVI2qU6EW8/aYbm0kBKJ/s+p+jgkNWm+Bgv37OP+aOJE0ZlM5
f/gWtgD/l/sRI38YFoyhSzyBV3KDfE3tDp1S1FEpOrMKa9aKWj1WKPujDBl9lPqrsDRyDt0hAG+8
QkgO3948Jd6tIzmf7x5otSmIjGL6GdwXrII2GLpsASrueTzvJiU1Gxx7Z81N3fRmYkGJ+fx3Lujs
KvADc/8lj4TYz9Hi2jqyZZica9aJNSI4i5debuYcX+whWKpMfD14BvOnaO1+jlIK2kcTTpNkI0NW
RSF+KLnRmK61LYdWc+7ujGtke3o8ftdvOcwuNUZuMIp8duBfAm8FEzJfvspxylCSfUU2s4QGkwo/
lCIJyJ3xQ07KDkF/nhusmBZkrF7SpulKkAGb85zDebaddhChidRwNOz7Y6M77JJwWAHpSwAAETsN
eK4WI4nBIVynODrsiDccvhs/7AdIJJLMlb8ReHTUodK7+o329hW81p9zYESv5vGP31dFdDzduqwT
8nvNXOCWxldZlesT9SwRlCJkZblFc0IWuHuK2PzngnM38hF1xwn3LmAJs/PCyWo4X7HrD8j2hb1A
8gUKvylSn3PNHOYMtSq9AledEhwyMnFtLZTrVcfF/NkTZUKj98/W90GGeadeUYMB8IM2Bp5Y9TFL
aVeJPJg4F4iok5Mf6ABzt/Q3R3859ioZ6jWF71W/jZVETyS0ChOcj8aqyR2b9DbU5qyDop9e2Hth
Y3fhSOfZeMbPz+j3yQXbyiEEJ5Es8PvbLko4zjoS5ULKTkKMabYh7JaOjubUmAq5zk9QkHgOW5Yw
4IXrqnj7rqRvkXtTMkOnoD0R7wuVrW9Jqj3/Hwq3HaC05jJKooMndUM4RhMEtX4JuJHEZ9wWLkh2
oiQuQF0Zxgivwzm3K4jBjTaIH3OEc38bHsxLguZ+vRhCg2Suvp2x7NwMJOSsWPtpmF9HJcdOx0a8
oO9Alg73SwQpYKsnQ9t9oTNqyf8/7J3DVqO8HH3FvPgsCmlO/LOx/FeUHZXkNo8wderkFU40zRaK
aPa6hnofyy+mGBpnwjxSYddY/Az2vfPMUIO088fgwiBEqLJxB3GY9WjyXTtSVb9wpQQo6s2Oi0ta
YDExd56pyiLkxXIA8hOE6IMFRWIMHtCepStvw8qd4r62/QQYs6w4kdnUE0vGJMPgZXz6oaC+fONG
HD6GYq/mPTnSU1QTMVZTpLXgwjiylOVZd8X4XmeS7ja0CZ9RyFvMbBTxDuvFuEbb4K7ocecNY6RG
cv/PWOp6x0GEppx7ZskMhtSbkNWr0cxtCaKE/UWyHfJ5sS5IaD1GDRZHufLZfcj/PYm90WoZH9k0
sEVBE+yCzlp+stqBy5dX2ZUC5efH0bK2LjrD2PazkCobsVJ14lGUDoKYH3P7VATThYHd6Hg0Aw/G
o99/8ueNPBwbNDCzLgS8X60gj/K7NZlSaWpdI9jZ9cIQxzRWBtsDAbcMkOdHKuSbVZADHeen4gX4
wZRPvT19+SEQAKhZk+7iTJU/Mw/oQrOut7F1RbHh/G60mIiN8upPiKXLx7SV0KXPMxQeZOkmBEdg
xcmxgIEry7mbaYY2WLCS1UaFS2xo/9nWdrgjk821GIDr5zX7xE4l2MRbewxfxlgzPZNFaPm5t6qw
RawCkFxfzp0b3y3xDNhtj7FmOhGPsPYnpHlFSGyAd/S0mGANqWK46KXUtUlTA+7oPLuA8fzS1SxP
MLiyv/bjQ42htMgzX1/yHjCqH5TogZ5zedqm4cv0JgLiz/b3kdKeSeXSQ2remobJ6UBpNo4YK+ax
U0FwGsEGMtR1GinhC4LRLxBIw1Ul2frIql0kP0dNkHgPxuedlyySiOYQOO6kOZJt3rNP9XDx904w
apxNu+ONjKJVDMDeyFFy+/geelMzx7xzM/uGBsAuK/8eIzMinlYVHs0IW1focg/8XP5WqHQRpofm
EoAaJrFkV6g5YFaD4vI+Ts3StqfFXxRlrnJNsalxydi9xTuq8rJC6dMXSbEudz2P3nUgorRvxJFx
Zp5rQtIivLJc4NpvtZG1etqyzuHOqA7gwkbpN1p0ZRuw3/Vu2KZ8NDlDbeRHgZmXhHrVnk45pryq
7WZ5QG203oYeb1y+wqTu5FvHkjXnZa6V/sosshlOPUDcwGzbH7QZo3qWbwZtpAtFhQAVbNgK3Pzz
K29/avO1jul7YPlSbIQhmkBpm+poHWFcp8Zw7OL2qF2vs2lVbeWBVzbAOtoOTUONRrm8z/RPuNrV
v41MgI0pkqm0ioJWyKrhoUgGZYNuOtmE/j2x2Fedfvy7gGAfmSKhAb7SnJyd6p5RBTT+aPhg4pdw
MfOpL7cZlnsnHucpW1kAaFZOXFQMJKxU2BeL1Ywoc3YEkDFD9gFZdI3o2zCg0mcvPGAqAajLTwVI
Ik9ZJvEWz6mepaAMqdF5BZ/c8yRO/npsDOiXfaxWSxSG0Ugy1v3iCLRRZoETYyVapplBOPR0SO6A
HZvD2O0riej7zROzOOylpsiTlAXOrp/G1/8FUu13WW4X7vKiF1iAufEftUYaTjTs62//sqpam0sl
ALWi65V+jqhc5191vTFfxkuNtJAl9lN2o8nvls/dYhsgEZ/T2lQ8d4ZoiVT/2u+Js8g2SZTrrQFV
0VvOtecD9V0294g3fAxR5a457rA4Za18TaaGolRrlONN5C6ujedgiiIi8bJ/x52bXCj0BTxp0DcL
LEwc3RCWEoFsJcy8uvegvH9TQbpM8VuT4E6nnnEyAQW/5heE2KSv7t6vB/sefyqcOjRI0C49sUjr
q+JdQjXf+x2jzitdTouh9S9WfzpIJHg7bOp3808CIS1BCk0qq8OJaHxYj0/l1FpxJ81/YLbvxm+v
HhPyRQHaFA2NKzd0OpYMss1iNgHaQfb2wcY32ICmK+5tvXd+9UgUbXraEa6CLG8GL2XDw2fZr/+X
1/8yMwd+DyQHC2Y53rAoPR+p9zmDDT3ElrjDClk6s4RGl/TzPmi5qljb2ts/xVZcaDob+5AhPtsc
Ku9BGMwKaKZO++2+OkUJe7t3zh1k5K2oPrdxGjmHSSTKxhCPHg661+WY/8+QS9JpsahC/YP1t02o
FKDG+KdDmqMYZZjOzayppY3RLhV658EA5n2mmnz9IYee/+IXeHZ4G72CeZt7hGALVTwt4dkgkrgZ
EbDAc+T/vKP/7WQo6uj54cvIIDO/0jAM9rbpELi2q6RQYnVmVWhimHQ7XoZfFaFo+6IOFeXtl+Wg
Q0196ietPOd/nkw4DkAbc4MeTd9h9tue/zHtE8mqmuuqBUAPygjLso3ZcudcqTtM6uKGBaXE/ZOA
Uy9Kr2VxDZ+3KduM4eD4tYHutb3JNeCkyZ4X1rYIUlZrmvSUOXbauThVwbdbHls0zQhBvxBpcC3I
1QXfIMSWq4S0tMt3yujgxLBMS37HYifDGvzGIt6BbX2K7gdzB/6/GMzEZKU94cnWXzDyWqtfP7Id
LGeNiWVGnZG9fp0r5J6Kio1eWLIwd0NvTZ03hsV0O7M6j9Ke1DqKOsNPTKHSduRf2uq929VhAfY0
CtXWZB//0jhhW4XpIutgZa8ZFXBVDVxNMvdIdDLuqUTsXkIf4C54yEiiYtr9ClLUkwLcI054rPO6
4W3IEpFZoR1I0ba21LTCJ/bjepDMb38ltjHPwuRYGNLhW2bTUljIuCaZwVCi8iyoQaS+tzbIJHav
mtjjWEVdBSubsamSaXL7l/WAsn5f2jzJ5P/Enn57vAqwg1ZxpUws8XU5PsTRmvEQgwFQAMEJUcWs
TYjDez+RsluXzj6sgMphBj8HdWO+GJZ2Bjp2ndmGa0NIUluDDUg1dMjOmyzZzLmLV2oWalwt2Q1R
okqtP4Z2OlNYNQBtudPA0l7kKotC/veiPfnGc9coO4aip83EVY6mH+0UfJobOERy0eDmjxx25krk
+Uk9/AVuIScu4IYvlXswSazd+O7ML9W9qA9C2fDfvTLK7F2TGKQSvcAbEdMzgDDVvrf/XLjKPFWs
uTZZbOiBe8SRCtbCKfHKtan+o1Z8rFbqaagVJlrHfF9ox5Au/WU/G5LGToYSwxv90oxnktyP3jx/
Tx3Zr+v8/ShMzFasLgrLb4Tyv9YbU49yFYNxnlkNuJze8HxAH+AIrC2qTWcV6vLvpEpHqrhAsT1W
m4ko1QEm9cV8OTG3tvR0+HqE4oe//hdDuKvVPq+9oGXNbm8yGcxp08nG2LFNK0JP0xcCkIZLdXo2
XXjePMcvM1EpLnVsDcm2EI7QgetNa0jzRDL09O7cHsMZfqDVWQEMUdRMcUbr36Pc21EBhu3y1Y3Z
iU4AgWeb3D6bwNbmTucd3T5aaFhVwl7NjO502i4FFBYzy7xzJdzeoQIl3foe36GViQo2V1v15LFC
zvUaLYMjfmI+Ajjb0CtYARUCoQqhuWDXSr1ZgmkZ9s9S8futRYkhTqbp+SrsbzuCMMB4MuKSqQcD
NKdaYXVrNs4fcG8mXf2ZXR0M6uZnHec+4fk6sZKbIIF1Qh8l+xOE5qlGhT1443mMYYSVhcpqLXdT
0bizy85KOxX+MPUHm8GEW0JFfXf/llAngu34EUxnpOnxCmSa238l43foqh15iZtPfGSx9JkKFkn7
w9+7uyHyQYRvIkbpTCa4+t9YMKbN5W76QhaE7WXRaA5Nn8XuKd9tU7y5oADfvuzGRBJeyGFSRRKE
cMnl2f25zUBYGLKpdI/6yMCuOIRnyJ9zijduEvbLs8e//Y3N62ji4p4O8P0V0ccWUxhxlSM78JCx
JmoPbFR2RV7g3uBBSTraUzTXE8l7QYdI6ZIYNgcyDkOZubRHdc0VhtzNUiI22Bclabx7sU8wenLb
20M9TBy5fa67kflYda8ehyimOcmsrBuqFYPFwYu0HCuwP/djQ8HcNIkHhd9exwHMRigrzXNenUql
0hAdITcSucD2AbYL2gHF72nCElSMA7s2JZswMMn3VUaP80XKtrMEfaAWdVVVz04y7hpEva80SrtF
Qg9W54ekZkFj8gDQhAuYw6K4C9I72ry1rz1+i9IAPdDVoL8VyFg1Zhm55/SOwecw6izVLeTWWa7K
awpGzSGTIDn6RQh0h2XGtPez6AEz17jrCDQhgf9Z5ReYLMuaS1cNuyE7eFv431I+BfpwzoAAkydX
1BhjBOYyJ3Mp2mZSK7jr0e1IOAkqSOL7D3R58huhNK09bxBqkFtaOqtONSL0dgPpzrr+xISIMFVh
W5S7kAzeAKb59F+yvCOfjBFSJYArubZMUmGKzvXmmd3EaIDWPfl90LoM5LG/p42I1nOsOFel2AfQ
692gea2FTHuWv/lUR6s/KrI4/LIPBJ4GOp+pHEM/rd6T13SnGs42Uka9TQ7uMjZxXsMvxwtbRSu/
qBdyTDpfeSrA/JttRvDTcBF976TBVI4brbLIABb0ITFJePc40JNpPqq0VKPSrnQA+vv5jAKac03d
LqvI4VVLjRIX9rfj49aPVMpDyEr8/QYvQIlrY4DBU+2uH2HIwoYFv2nruLfCgQUBlI3YqJValv1v
DEQkqNCdqpE/TSV3I8AFtC4BZe3azNDLtH/pUGIggFJSUThilC7kSruudKlq9yQz18Wxckg3ci8x
KiuOzuxBZkLu3RV4URibq+hHewXP+dgsW1LGunOCtl91Fgg2sy1gHH5JQzNoScYbTUgwKxM+ZfHM
7m7p96eK/BA5nS7JN96qFmCG00Se0enLn57fMeIuC4fByDIGLmCfKB/fqyZA5cWFJ1BtO8S7W3U4
vkXYqqyydAsx3le0WYm1e1xyYGj+9UWDwKonIDtnEuTlpoBPdiIghGQNHPb4OzjEjeOr/MGW6K6R
3Ln3cRY91SVV989Ibexr49xsXuOvI5khsiMfiQd4HK9q/2Qj8KoPK3KMDeJwThXWQT7tEef1EVFg
NGbhQ6JXRkl6ufjHVNBKz1nzbtHOaiqGMpuDJuv8exPUXU/eEjGTH/JKg4GoFOLam9G44owGIZhZ
nwCCsXX6iQMrgt33EeSwBVA4tTtubgPu9NUuWfCS76oP6QDzcadZJmBWJKhcLH08f+nJaRrjb/gh
pGm/hPQsGtLifnb6p6kKLQ29eDaI+P6iv/8lYqij3F+woPfke5qcBvTAhUzqw5Jd0nuFD9drbIxO
0AdnRlbXo2OBgTIJ2nioZM9kKCtgpDF8xF9hfcpjMYjCDXcPX8y/YMBYSLunALGa/RyVlJVFXkmY
zUbHlvIHu+WuUozlaaZHEjxilE5tPuhTJLdeiJKAkDR/wQgPXGdUtoHZ9Nw9WwI0CjMFGl4aAH+g
uEbtf7ia2tcjliLphY++0hsB2wqSqaBdIvrKT7+dYKc6rH/KIqs9SXEv350I+SQyFO5Y18qemlK0
VeAZq1/GeW3CK6RQL23GAk5jqmkOVRboazvQ06oaEpdk3tEeliGVsqIqQBLT9ydDlrHHp8HTrgMe
7az25IaumJ+kj+FHE76N++aimY/w/itWir8Wc60aOpJasx/nml4MWN7RakJgb5SoBRytdFfnye4/
x9JX4yNmim6UGqCJo2dk7nBWO7ZXz12tBOQzKR0NZr1Tx1vaUDsNhbjS5ytbh8L8nh/A9lFR5qTh
oXMxU9xYB9a8T2TQHgN2VtzUwIRGiIBbcqx/wGsINfdJUnNFIxbtwDqM8AA/xmN/FkatdSJ2SIp6
0ZcCfgjcNsBw4Fmv5h0lNQLPqCpciztitzbQ1w15QzJQhmIsEtKBTxtSrRlgt2BP1aGA8Xi5wwzY
LiBMA3kkZTLiiTecIgZE6CeWvQUIxG4Q8dpwFXr4AUaTQR/CupLkoc03y461H0I1fd7f1aD6F3K6
nDerxW98j1hf7I4fRO4hZbuAe2BoOvp18vQYEFE9PY6RNGomD7aZJ/arufjUWSzRhOK9GvwZJQ9m
nOTCEF0VZCtoqJJrfyKMht6NcVVbJvWMaACpzZ2XkcHxmeEKG6rSYA2Eij87c8u6vDKD8a2HrIpK
vjfTjWg6gHeqBlQe4kPz/pvY/nfcqz4ZcGVFKvwzJoiybPHo4sSrlm9F5NZh/tM/uJiUOtzYf9ID
uKMIYRltQ0P6vb/rgS02sy1xb/xgVUxY7SNZG6h1IQDRViO2swlvTUT7s6JEsCp5pNYebDuMdTDM
uzrNXnPmtBw4DCkse25IpHgfNEyxpuX8OpvPeu3/OTZbVr2uXg5lapkwExM6rhdBPn4y6T4/9avW
LMocct0H3z5WOtXBRFEhNKFPpHEWHuCLKai28UUZJEjZhNPJpUaxCi3oj9BqFk4VtyqNsQ7cfcgf
XoPbB3U6cOhG1T3WbkE97+y6lJvXWtvPXrWz839O4/UxBsnw7ScbuvZGuUGjlcr7zgT3H+b9/YfS
uzdufSbc3hgHGGMExdDrK7ffCmXQ08AMulzSpistFzmgRxXgGjz1pjJOWrf5NcLGMJoZIFsaCFqy
0ryr8G4gAj/hbCRbdYt8CCkTHENnjHjL1hw0p/Z67UzSEIUHF3p3S5m4B3z1A++T+9C9KuS2JR/S
m2pAf+Mbf1tFpUal6kxd04pdIU2QzfGTurs1o9bY9hmKOW0yKX9MSMB0iCWqT5auRM3Tp+pUjhv+
4wxXO97aler3rwsAQttO9RVGjeFdZg//z57cZKKTA+4D3gk9+/LggYFeqHQmRRNqhO6z0rFy+cPu
bLJbxssNTvAlmHF7A1AqAd5ILJjPVxgALwaEtCWat630ZSkNh5TpA3kTj+qFhAkWlMl9MH8WOqEg
GfO7HwH7Ffbrr3Z4dH0u8GU8c0B+qU0hBXYK3N27XNfx6m07oKfpt2HxshkXaTvQqVM1mON4qV+P
S6YYRM8PN+/ALKDAtr3ebQSSbojHERDkS6hR8gDgMjAC4TuyWaWa5+2gPUC19FVtI+672vjOqL+J
5ywrw0GJ5291x9PGScxcUTVq0fAnX2N9vSu93WVh7zA3JiXca8D3n3kjzSvrg+kthMs4xEPgmKR4
x/RDELk4T8E9DWRE72+d36WrdYWuZFyJ1iSB/BGHAwLFGieWfb6X7wZqDSGB+7O0vBhE/b6Gmx69
+3A7vlHtDyqLOR8Bs6dIO8uYUMGUtVeZOTKf87tFz5EHxrQ03GQaC736RetGYAvO0DCkFX5kGeBb
SRqCRpFXbrls2q8EBbhTdHtsgXI6t7b4c6Qa/jGyBkBVQV9FYLqyYMregKeHMIqdaNHDg6IJesE1
snUL8RlgEEqb2Y4A1Suoek/Uqq7tDOoVDQpuW63B0nJjO/3DJ/Hc9KVN3aha/MHSB8VdPydrviF8
uGHYW3Bdq98TQdcsfSCd2wPXSeCtLpscO9yBBVOPHOJYVg45+R15er5O1oQogZRFI1QhZds6tn/b
uoDamAGKbtMLEl6tr7RX371QGQNsrJr7Bsm47UKwnQgc2BHzMiSGRZaP/0RD9bOW182WbRQAfM1C
VDJ7hqCmBhxc8PtmOQv+nd6NOLSjbnlffsOxsKQhgeX7TXnWc3MMnz1K6JH0Ymxb0uphWTD7mXsE
NHS4Axx4oe/kaHYVV4pc2L+/bwXux2sMIfG0gB7QM0pgN0Ambbgg2+8uuG0y9dL77PrR4QlLvIdW
q97GH85lqJIlrVxBHtU3By5zGPDoOXpXGP0b57qYJHls+6btaHJwPcaa7yGXHKkOmdmEjAixIGq1
HiOaJxFTCjpjzRR3xOQJu24HbXCUL4wV4Es592ZIgbfrLSGsnbEcB/CCrf6++qYgqZTe1jhAO2p+
idOO8BOylZS3FlbaSwIjhT1zFgowP/AxXNfwT5yqeU2GDr5X8Bwu1XLb/vb+e4YCDBpNSCYFP/Ee
hJ4yLte+vs2j20g39SbsDCxpz++W9O9B7ilWRepX0DqV280uGla3b30Y1XGItPlz2/kJHvSA51tC
GdyydeE5Tq34kAMT+eoSnarnHYAaHCVQy12KawKxRhEWKPaqi0UpqJiiyMnObEJwqDog+PI3Sbwc
aR7L9cf6r/MGwaijBd/iY+B1RbShtrucxS3Zyvw7JsNCZ6BujkA4fMFZK4KmT2S39RhnJtgndyzq
guybWMs5JEmdaguBv/dNdJgpHlmeXdRESXtR55e1Jk+ciApjKI1nbq+E+ttqYICfMPei0jcQv/OX
Kiqw9G+Loov/14a3hsNsVlAm4r+r9JguZzVDCpHfSwRHLciLfTDT/RIu/s8wJQLLk6YCAHQuJbdi
yhbw0bsyzgdts3YPZ0GFHd5SGU189UU0PfJ9pSXtO0i8jgHFOW1mj1d1smJXGDfPG9wtJF7CK+Iq
O3K5SWPtHCOJcpuX2zy2awdWQ7karHfW2b6WoHrV2ECtUQh0eoiixgdD6UBtYo/zOW3LjWzzk/Wq
RdiMX/9IiyE6MKXZjXJXRitzE8s1obj2U079oqYCFfsFQRZyvR/uZOyN0FG6QyayIr1JALrk6oWM
RVRVbtlht7QuoSxJENikxALtbwdh0bkZWWSxuMQ4x6DApjqj2eLMD4iL+Dzz3/5wKhgIueGr6JEm
FCpGosJrsCFJFDqb9wbyrXdEyMd7BcmRrP0cfpiOSk8g2oWHobQKxFtamEQ6SndGMuwQA/ZEqFZ8
b/IDZUA6Wa2sx1qzdAFu0Dr9Mv7z8eQ+97rTfIvXEwA9Ju1jIi+6XJzWlG0MwVWIANbUSNGf7clO
dknxSPiMceYO8PslDkZpPKUSt83tEeMxDHvJudpdzxlu6Mo2cUc0NW00cpJXfBcnPxJ2uF2IWLJ+
h8VTm38hoUOqw6snDUV+6u39QdiEU2TPiSU/+AtKvcVPuhLHdc5y6UHHvlK/ttbXMj2hcLU6z5aF
BWzMoFFv23lTM20yLK1Chn2XrcMdeD6DgGvwJoowOHjmln9WamoZj6VqUgRMSwhbDvXhwv1z1n/y
f3CQe60jK8h4rxZSot4LFPNhqwNM0u68sdVUUR5xUxr7PJ4B9rPL6xv82GrOQ2DXZwKaQWMDXD1p
kqm5UOVjDdGsihUt80TL4ATw0d4SnGH9pD3k1gDA3WWVTWbCgHFLTY13M6HZX5NDQRo1PqL/pWrg
nU4WyGEAbwDjalWx7GmaFw8nWyHWItPkgFW1FIj2NNq3sTFFAq2OKU1QuVNoPSjbcBnJzaDnyjua
Q7FlOhwPuPlX83beo06+lDz8rc/txdDYFz72HjbnEatH3ZYgEjlosOgsQ/eHJFqZHMqCVJTwl88R
W7uzLc5reccBjVJufe9Yo9QAhXxAumd2tsm2/2YA1jD5aPA6JxwVpjkwX+TrAMqDmjDfStsaKvwV
CgSpRrdRU19yalqtSgvyWwZiHLpQsTLFtICO6DTA+dNxbjUN578UTSvRNrKw7T5+V64P205/5kjC
UQ+LCwSCD50EHjK9AAsoOP7OSo1wGXrcEh9MB0y+cFrinwBytaWV6oIH+fncKAlWkiaNX0X+tlSp
4ClWfrN4FMcCPR7Kw/GGwgxg5QRp9N5fJ/qFBDLs/evGxQik11b79jS/j02J6+NdiHg/ki6TprEV
V5BP6+nkCPOt5ZHNxvqWfZhDCZeA8gefAuoDFvurgBBMJxJA3aD2TOXFpArdxzjq3Aegt878bnhF
VWJR/aa3uhFN9iTIzWbpqTvUJ+vMpOTV4T9sOSaD8aCrBJmlRQm0U2LZ+/4Lm5tZJSOFgG5CcWsG
JgmG1isN68tABijgfYirirLns93mWZZBXrj4AOp17QxSn0FOOlpl9XMoxHOYO8LuNdZEbgPeAo4o
6I9d+Hd/TAWQGnTUExTKrsF1iEAhV9QRiP8Qu50WIRpCPwxT/j9BHcJylCBm8mRovQOqqbwZs5Pq
cCh+6a1NyMCGq0TcactCEmSMoYM5eT2Ur1YBTKHkzulOqcyw3+/4SAGq+SI3jPhAacI0GPCQeDpa
C1mV53mgL+D7YHeSSQ6sZK4UDdSlXfUWQIgQa3bH2/bdwCXG0dXHdUkgo/jvsQhdEzTiZJUd2WrJ
FWDGysFfJdut8hpT+Y91koGL7PkaP3a/fIH6ObWRjrYgyPAakDuzHxkF1Wt31roWGF0vNgtObb53
LKAx8m4QYBqIN8tbn0MW3b3IOe10JwyOKVw0iM5PgxW+ZaCSkZZ1BmgMeMORfJqomysa339i55Fv
4+F7TysM+bjlTNewmv8b479FId8KJN+qFR6MISPo5xi+DGO5KdrRyjylMC7RNFeqci9a8sg7PpTv
bPVOWxGDUvUFIbtRG0b/4vACguf3G34CUV/Xs0u4c6g+jXFKWZKsht3w8kq6kEGfpgDqGB4eGFTq
9QKimT6LkqUfXLSk6vzGtc5zuXz6AFIrpgp/wk7s+A5rBfpDGSc5DhgWmJpagIBJtme3YUBb79ft
u4i2L1mhEUdij9KqTekyguP1LELi41p8lChsvRWECBIfrYvQ/4I6xP9NSEJH97PWoWnDDD6BOTgZ
EWnaBxj3Cm56A8iLpmhYG0YQGeOvQMgIg1tsRuZpU78/32UhFZGCL09CbOF9SEBe5i8ltvBWi7EQ
gJUtzdTm/od1qvVL7ZPgPPG8Hi0Z/wZyRMgxiXF+94W6rB+otiLxI9Dzd4gbIQfMLvtVq5qoB3Jo
2hkUreKniYmGmpG4i1QGOnSoZvtdXal1/tjrPRLPM6dW0BCh1x6TzPMbpMxFtIvcuEP7Iyh6XsVZ
t8RMUs+ndH1gDH3v2ulAgJ8Eb5L6hylNTqy0aj3BU52PTJEA0aows+TLFPJm1KEC1W17mz+mVFSU
Ksh78U4HFAN1ykPlUDxbhfwbzNntT8NTIjET1/iyg6WJoo7QVKUB4M2CpcRsWRKkG0vPejiemWFR
zAJowT01vrjHJu1JKudfk4dzFHcJ6XDX7+iP6fSPXf74xZ3w6h5V8Rhtm7T6B8Xl593isB19OT5X
6rS4A/rrugyQ5YYAIe+k9YDXtzDZTKUjIsAgdqi7U7mmXxfa3b7esGI+JT9AZ4nrNbHTv0Wdr8Uu
MbMQyGHQBfVW1a/vRF2jXk8eOA4cYt9EAXjKpDVOeb6z1pTt9ilgLQM+CcT3Et3XYToL4FX/HD7K
0v7orMfmt9/u5Mh+5Rdp/oluJxGetTuMPRRgFlXymhVa0PG5XmogtY67704B9gh/UlIZ8iyNuaRa
b0asGr11n679GQVaZWqrUDRCzdttj10a7FeH07n+0NvUsB1dlEQChFRe5nVbH0qRtL3FD6oWXgkr
1SuhUBMIcIpamjIFLRIBpsc6+s0l1lqE89X1Gl77vJOVIa0JcHPtAsfstS6MEZo6OaRpoflaOpZJ
HsDtzB0Sfxp+Uln5Ny+Y8Ka+uGHYkHJ4t3DULxAvDMn09TeV0aL0VB2hfRJAlrT93BU2J1ZnbCjI
HSL4PB/bnK4TFq+Hr5D/svuGxSVusRQDPn4GhG7sv5UHUPf40h/JOZPnxsgTYDj5jQhw80rO8/+6
CadYygR7zWxsHhpra3f6+7lTG6lDI9wLsphD4Vix4FSDBL0XItvDiE4WZ+W4pOq9Sa1F3QuIfU+n
iUp9x2NDGzIThrbyBRM74L7tPGjZ9yKH42saFJ3fv0kwsVI88AmF/EqCtP9tWzAG0i6h8YoQbE9J
QHYUiHCM8ikyHvta5MACkql8UdmYMJXZsmuu0LTWDra6sU3XpJmsT9MP0CgRhllspPWi7qxsui9W
ZAD5TC66d4oxA7URBq/fLg4p41FK11Z02tSSDYGw3o9JPlFLahwzU8jP5y6DLhNXLsVmGbWjyTIP
9PXpojVsz7cc0IQqBZp9txkHYkMxt+wiTcFaWQ09n2ahSyPXfNJDg3Yiw32KL4YVHBIvhEblrB6V
VUsBm1oe13Ggh5Jy2oqHRtnxMsBsLIfM764zZXZBt8beVrGw7JUtmc8Tml5jNotI2/BnMTo8QwTb
vkEQnN4GKp9n4c6F1j3Uw0FF4MVJc9jgbq8aIBejn1rUawtGyFTG5nQ5K3ry7c4qrVNP/htSQrqG
9dBQT1M2nAdMki936OEodGxdPhxPcXjdGB28I1Y9Qn2LZyE1r6GRrhXmkFCd3zFo+YXqC+hS5IQR
XssNFFfIovWpDub9fMeaCre7KKHQtz3Bj7XbHy9DIJsidjPS7+5mR7ZexWgvlrSHpouLrXOE9wop
qZzMNMq+Azkkik7rqARHVHkAaGXEIyTwi4swOxuJFL1L51UvMYEfTpY8nRz5xDfnZ7C9TvN99UQn
CEhb+kpx427PhOPw4TbL5h13GqVaHv1S29iT87WvZmT0XJ4GJZ4sXy7XZZSPNBBiuA1KwLQfWec6
tyv5jOWQUOBB4HlzwxPtBbD6kOjGEs8iHWWZrNvolTYEJJSBKDqzEkkj2Vy6A8tapJfvrwhweeTl
XlDSDYmDF4/S8oLCgB+TXTun7HNqnHejDABqBIF0VjAEPjsG5ZFShR/jfiKZQDihVcy7Jaq50yMd
nCTWF9LYsZJ3mk35+fPqDn+i0RwCkjjU7/YiD8FGRwxWEr+f9ZZFYwhvclPdde/kSKIcCgkW5j5W
K4Ltf+Nv2MxLSLR9AE5B7MH9iibl9fjVvcqLemn8JxcsQGzoX4jR2/nj62F9xqCltn6ZF13BWgHf
IgQaZ5XHdBaAqgKQY0N8Ui5Jb7OgPTwJ0a3Z4JaZpihMI2ZsI7h0AJ4xGo/+80tSJFdlxyqGGVPM
EtwMcJpm8TVuaGNsbgDVGJo/q5aw4aM0mOX6P/dDqbcZU11sY6HlrbaBbzcqOYfQ31tCekQq43UF
DBzZbcX69j+skt0z8ImCxi4tPW1UPrccXa8RNErlT5odtRfDxW2c6pI+TViQKSCyTaUythqoKnvK
NHyx6H68vSgEMkCl6lxjilQ2T8SiOCiiABxpC1E9w1fyA5Dw+3XXv+6wa3XwPMhJzYaXRO+jX66w
MyRd3qZMnU+EWE3uUWBiWMxrff4ya8GRrv++HXQR1dBzRNovg+if3RHCAnQiBdmQYZDMh3Rp3sUv
XopsrYIWGm++loCrViSkid9NZHiGLA383ppNaTSRS/rWHa1gSJe1ZOalAwbaBLE4tryswgfEBe+d
eXABeuv3lDfmgLLKiUCmzguJ6YQRPNj6Mq+c/0IXbvfGR/S96bxTIbUdYaL34mRUZKB8dkAEmV3p
j9/uJOL1nhRT76Wtw2qRzLskIQU0bnPfCkW10JfoNmPtlEXIWtvPsJTV+ryjAoFv5h7ix3MOcmTZ
cqBUvZ4zwKpFr0Vw9fChkuwceT93oz+hseFfzVOP/9WXivCp7jnV3OghV0uzhDHEykMhdGSbmYZb
DPiCHmwlOIPwp/4u/852arAXTeVvnD55ms99VptaiHi4azfrUnwgr+riunTIRQMmYYvFmedcGZJr
SvWzAk2Nys0TpTOz/Y9/0kkhPBjmzAQaWNGr9AeU+f6QiFRMKUkciTbLNno9zLHQKY9zug3Kbk/v
Llp6txRVVUwfJNSfXap55AhaDLKsPeAdJv2JaVQNRpJYFVwCdx0HI13iBAZEGy2h4lTgDUc2UW9j
INpHnZv1wKC60vSZHQyPhWWqgNQDnm7RfctaLc0QR6x13IDO1mA/W71kq0/iO4qiRQBpNvvw5azh
Eyf2y9DxgtCBiWp8eL9/F1Rnod/TfTVjObAlJbDanQuckQpifBTlyvTIs/3cYM6Nwr85iCMRamgX
w6m7Hix3V1EYMhLB73rSDmCoYNlD32BTdfMGm2sT3rxbD9c7pQy5LZNb6ldcTgDpccK9EgLjCGIG
in9y9INbizdDpnWKCuLka8UzayvGz642URIWjz/2ARqbQ/z8I/ByDGy/7WIRxmmogj1172/lnMsP
nnWqqnzVJQBFk2d9n3UfeMwki6/iRv8AJQGrfFOZxmbfWWaj57wYywlTC2Puw2XKCEGRATs6iAHH
7xqzpdhs+i7Bg2tbI5Og14WYIi/qAMPHPM9rO6/dUcIZCcmvdsP3OHHqVLqGUhWEAVpfTg1SR/AL
hJIqCBFo9ajDhaOvRowIRJukD04AUYrjuEO+Z+zge7ihzGnIbkNq6gX6gRNpL79Uz3gOMUj5qZBp
zrjltejw0gt0I6ELwYGV+Im19F5ggtmjYaMfmuTgOfw8cAbRk2IEQ0zSqWKDc75pyUEyB6AswKVq
EuleKlydNQX5GZC6p9SdTUYbqPWJd2ESthD/1r68tAwerHRj8WOH8Czzipnna4v/Qba9mwd/rC81
Qjw5jdrJ/hqCHTVIOuqwpaTEQ8G2F826t2tn63e2V/TBhnC3DB+rAd9Lp2ds0uQaAMruh3ui8vXf
tD7WhWt5bIMLikGtb/KycIgJZWF55zKYbo6CO56VAfUooiIzu1yaSJyn4r3PckjTsVsH1fUgkXRr
Hf2ohH2Bwp7J307DPy+sQrsJJJ/nPrnquVJBjEE3z6uvtLTriD+OIDTurJ4EbzvnYHF8O74TCCKf
p/LbFjACD3N+E0rCTR5NURwdOXT6hxx47gAHksplVJ848+L8hyUe2vxbfCWGZ3GsU01Kc06YJDX9
AmTwyBhtXJVFQLYJDakDC9/ezYDq3TxTO57nV58CCrYITewOL1ThoLdJ5SOAeBFGOMJQmkDEASk0
NUPYnTzIlA7bpyKtO5Z6jQBwvZ6VgHFui8/BZk0jB+psT7IX7o/7AOr2LSN4vvTS1BbYabbZrGkE
ND6Fkt8DEdJQsnJ0Jdx3niOzzTEh0itzjk6WX5XVDxLFm5pcDPFNts43vfKMVfxi+tNTp/TZ5G0O
9iWqCD1QBSjM4PdyRVKB1/gG/+rq2+42fVYyFlljLIR8REn4PI7BIXD3qo+MuYljbcNpvJdsmwie
gj+JZuENGBJq7HVnpFvoPbVawYGmF45nmwOLRPofQ1nZNctwaaJ3xLlH99qJB6ao9fynIrx6VOAu
kb1SDwbnSDwT1uaLZvskD+dHNT7GcbtrKajdUbuJcbgIGX6cXGZmBFRLc85MeDDAmgovV+sAomFt
O7aMxC8eD5H54jvzfegb9C6f0QTFEhh7Jsiruvtk/1XCK7yD3dFheRrdpDOUiqlM4IEeVs7DZW17
+7HvPyTPBqYlpwBye0DdFPcVf9ZnC9OJpnB184uEDN/g+5njKQXicg2c7CkCUDtZHR680WvfSPtj
9s0jc/P3tAqS9bOQg4hoQIE+6g/9C3a6pTk4JfgBev+TbO+7qEGb50dSDMXI+MDHIdhKFWmu5pz+
kUEOSS95vbfWCViPQ1GSd53DzvvndEmbX2rZIhmCLVI3H2yJA5Co6tzTifJ4jPSKETnRE86BVarg
S93ru3RuLljpUaKmVKykRA+yAE7XiJT9zguf3/GD5EwzcQjleKmx9BtlKRXWX9k8+Wf8eV3Uzrra
cshLFz2Dq49rY9LLeunm3emKNL9QwJBy5U+52JgANDkmdmrkiITF1ttfVReCYoEY+cRnkhie2Pe2
+VJTEkg7PV4PIdzErcVlkWUJ7NWV8dGNBvmFVWF3ZdGnjhv2CEfUNM/UNFFO9i9isKMD7bZpUjTg
XTQUqip0HGOi+WxEvaRZZEqj6d105rfxZ3XnGu5iaXW1y0vug0FDgyKgSLS1rspzZj3VFJx/CSi4
dk+7TWFM6RH2Rd5L45bQaKdXHGZr+WGXcM7+k0RVqkAfholluvVl6x4YnalLWALbedgtx52aH+nq
d5HpdB0eapzGv3GmdwVCN/tAxQpMJfN15uDMIQsmco6WHrmnA1CvQzGaw2yNiQuGiu8glt+up9Ce
+p13VER48TAYEGXsrewsO8GnWjOMSJFyQVpf6uN0IkMg1xTuLoybmVpO/iSs5TG2oet4eV3XAV00
kfOLLFPZroQcS8UXjsY4/tSy6txsPjB/CMHiATK2Jm5S6aZJ1BLVIn/oma/ErYsrGhNDDblol9WH
79TnuzVfK6Hudd6ahYY4Ed3VIXS6T90ny2TxUkt+KVfpmcF0f3NChlWZ3U+x4n1IU50zYyLZnkrd
LrgLhHHtlsLtjyQ8PaMiLgNteoPxbN8BCtgwc0D1+taTtANZbX7vQCPwIuc6oH3Fa3Wi+T/xAaet
5uCm1h/cAPhmWdz73teVRtRnuDJThsaLGVn5PeSy4LNyPBpGHUNJehJUsnqNab9N3roqKIxFMxF6
xt0m5CcnO9foDulWPtYMaKnOozO3XX0CgGt8cMiTb/dxymCFBqVJD3wFsCakERv/7LgeGqTGM544
FmBw3UD4KINiBEphACZzzb5qkZqunINDNalRKu76T1BhAGM2RQvYeCFhiz1dwagnFanIWJ5ZiACG
Ddwt8NlQFo3yc6vvSH6Et7W4ixS8YjHYkM9xnF/40BRAV6iOBKN+X6UNrv5NanUrI8Wc6En7NC0U
ufrQFs92DqMjBmyD9nptj4hcuzIdIAAOKWEg3uNB21FjX/CyxdmBGWvJOM+1L30kMPpedjDwc762
FoUR+w4/4DBMQnLSoTNjQLo8bfdsJBmEVElAI6y2W+IJqm+zJwUUhra+6HfXZUcvwzke78vNpCv4
hhIeMsY8pdnkKWdKV3cTPW03aYvsEUqFNDb6XAY9uUkC9UmaxE2ndtORnapt+zEVqV1Vx6KoOfNK
PdtYsyZvQJtemhqMuitv2r7Y/MRVzcku035ACJ/5vaLQv236CGdR30wI5cGDf+Z/kPc13jPwtHiY
DiXYQZaQIKAusCzMt7Wdxwjb1Oi++rK+drXa+Ol1Zhuzo3jGqICrywyeuh92cSITwUk+WBuYkNvY
sqTVeaBLp6sZCOl/10lmJnZqyIeHqxIq9W0YN/4d1G6OLBjNevT14YQg9ONLXfG+v45gxo5rTLEb
ilP//s5fyPIb39uRGxZ9/qLtjJYqfnQbNtggEy2/QiIIfa/rup7CFnDD6RRXYxcvf0FRjSNYRXpB
QUaXNGVKhPhvsoxB39Tm5a+6l1sIdDm9uL4qPmdJIn3oAOMJb4D9fzfSG+OTsqqqrbtSpmHeJBZt
6rU9HdWsHc1lQoXRj4U8oprE/NpoZ0HBbf45/OoIwr3f+EsZcXYozLD7Bf75RyG+ccaHZps63B8X
q9e8cKW8gnf7nu0x0EFxm94r3NRHfSbi9j4tBIyFrGOSsol0npVxQEwzhbsYo/j7WQRJptZF0dts
hiWy3ov5wg111UkJyLcq7KMcxKARz5oZ1Kx/toyCmNbMjBdSJKIt0zfLGPNMKvSvx3ZW+t0AaXHr
R6eNhEYwI0pVdenMQFoXtedxl7UBUibL1mcePv7D2pogtb1Dr1DUiWImns0E9yY0A//SagaWvYJH
4HnUhcOEFhNVtiNcooceFSCrPKwF1NSOZQOuYULovJn34ySszIqoaGOlj2lqiR2Z9M7Itkm13J68
DRCCETZAGPErOhtdofX9fB2v/YYDHYt7PUT+0Pbyi+mnQBHMETWkjtpqPjBIIOAFqYi2dgbob9hx
AuIPAvXz3mQESoh09d/EVVxLo8tWeuT4EoZcS2Vtm/d/B/OXRSFJoRDGOhDjB/Q23x3ta4Z3+z94
bUv8qZA6ZfrmMfJ1iqD74qeaW1g560Yve3tf/Jbn1GFwDYRMjJq2PCW73YcGL0iFBbZN8vjqtYjb
x6TGxf4Nfds8pA6xi8VNgK3mDEt53n2Qk41QzxyEvTFJaDpNURnZ/Y1huCkD/YxDvrGBu90ktzAa
gR9+n6ku7rHCa/DAdk8lVel/uUlZdVAEBdPwzPMpc2DKYfQEhMnttNbN8TwcktMSlP03dL2dGptG
i5PVRQXnnZFAnzS7SDvFeKjmZKdbVRkgGGiMixqD9+yvsfIR1CSOshVvvgSa5I+PQVb2GzMci4oa
abxJnrtdoqLSwIih+izU1bVw6PevekYpfzgT6LetPWfWGFYAeWa+r7ya+/BftX8FWIRBb23hGIdS
Kg8ptPcRT8vnBz5lORDjckcaHCkLN1eo4sWNqAvoQAvpe2i4zLfVn/LtZuJNxpkhMtT9RQd8kb01
2rqUFMXGo9InQ8QM9IPBATIY+rz07R7z05vvxcKR3Kdv3oWZClJtrBpd2csqfNrLC6/q2k6D7Ocg
+5dsHzFEK+lqMUCPJ6da+tnmhsR532Lkq8VK6cLiJLZk/iaq6Z408uVKxfTS4FmcJlKh6WS04Y0A
30u2mn0zhxsc1ZiU0EdiuuMmK6fLwvwbKzWmTSM20oUj/zl2BN47X949KbcVXnbF8lE9CDKb8+9L
HhrRHjHBPUD//qe8pqkmYLOdaU2eHoX1RpSXbW8vIeGgkW1ueCAXkPcBI2yhVZeNhzTW6RFMydR0
PyUQPsFKmTKXJMPnNUT9K/9kGUN5vbg34QHgT8/DuKERj9czDhi/5pPMUfQsnCSsjkqORUM055OK
dwufOlDWImbRtFsWgAtvV0oH21Ach73utMG/mDcyDKbQudKOd+EZ7HMQSQn/c6FSxAktH+cPON4F
EbfVnLTvyyabPYvJic+DEt9r3plQyo4hpzbH1++Z0+S+6h775N1OkIq2awiEisiCX+5eOL0sjw++
UIkzQvfSxmpH87YytnB2ZBQ6+Nz33q0HL8nH73t3qhKu5t3kR6axaN2/9h8dT/zAvWEYN7Cgu4PD
R+g+aimK0n/mn8bh/84UTdsfK3ZVgLktkCJH+jpZJ40oTyJoohDOGVCRpB/WB0KrFG8WDHwkUvby
rmo9dXQTulGH8V/Q96DRlc/+El+Hs3AqNV/Z6o6ZvNnx4lTZ/0sTDH/4hYif7n3a9H7g3sXwuffL
Styl1hmVQHSppwcXitb75vPI1nSyBEafvqeYgJgwFyZ6IPkGEyCH1lKh6rKOKSGqnNqbeotVsWqu
qYoGmegb9ROnvdHB70ovAGe/DKpK9S9LcC5TRFsRqgLYVTzlDgkRuIchuEKR+BK+e3xK5SQbh1/s
2vA+coaHkUEH4uGbIUNGVBKSfLo/71lO8S0lwOeX56vFkuPqQ6CEhi1ppvsxBes3MjjK6RMurSwT
pi/nmGiKumzm7yDlwlUtmikqdooBUNoglICI0EqvOB4zt0r3lQ+2oo7e5ig4x3bMnLHJE2B8l73q
ypQ1zp+Ai63MUqC4qiI7BOuSSpcokJ84fMfLbC3jlCFJhc0hMKc/uR6rit1nEMUOYyGP96mm85co
3ogZzER/4ZZYT/oRG5bJQaDlNdy3jH4f/vJxWsvbWEvFMNZ0X3+O7Qto9VGqFhW7tqRbP/RKnQ+4
0F59+dd+HZkaVWVU3lXiDdQWaJLomDvIhuI56HECg/iPaG0FYVt5tYyMGGsM/5mmnwSkbasUOtFv
LxNfjwao5ds221k8G97ZOg8P0OLLCseM0O/tbrQ2yrOwmW4wjyNtld3taESomzXpIi69bXszztmm
r2n2ZqwEpTtWbSv8Cnmen4aBS8uXpomgM+RzTJ8hvJQ2zgVyXLTr03zWsF6nSdWR6OT+zabejqJB
Gg3zjPUByfzUAmLoO08QBoRM/m3mPEQf/f5xWSze4GXzceG8w+LJkY6ijJKiedxL95u/yWtv3jDV
YZxztjXWaXriMpFB67Zwzr3O26WKU7XwzuE/gdiXAmpXlFhh8eJklKVAn9p0I7wxxrNH3VUNqtRb
1D0Iq6m200Wp0ul7tChK/J+zcrM01YMeWCd1pT81GxadeokQZhFrNdcDdftCIwtq6zZxpmu8KQW2
UeOXlmbvFXbypGGMS9Jmsst7mMLTaEFt0s54Iz2zuEvKZ5eXhxiAM076BkXZwC4c2b8yt69fNVvH
9tWiMCq0I1WkOnjVwAoIdvw5N67Rds5OBxu4Uxq/OCi+PmGTgeMv0O3JVdXcWlPWF4qltgSbPJ0T
RqOac2blFUWKdJTdqURRY8HqGwO49FbHv9+L0PO19oXFHz9/DxE8wDMHP0424FXmQTBY/QwlGDPx
Ky2mUMxQNA==
`pragma protect end_protected
