/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 303392)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B60UGYywDetHFadc3GMQ/M71wx/dqyn3Ra5zg1ThIp1GKmBHD6CZkI1/z
/+2HDeyH43b/WF/JJZNAAWBfyUlBhEw4tIVfJJtn/Y/VonJpyHA0qy5vOzfsQ925ZMtCzod7jBm1
jc7Hc41YYchmkX7sww/Ux4KrQ55rlfv7Q7WwT/CeWETpnTxuGohrKXI+KUKd9yEdpEEdyPfi8YqL
z5MMNEUSeOH3Y3UJx8ULaWTwQh8n/pgylhRETUa7hlQRX4Vs3Dqyslrp7xrXq6zOGQO0cAcnnGeR
dM38n8Zj4u6d/DW+/Fs3pPEEqmVc9pOmva1MpM1d1UysXcXbm8Sh7qWZMLDUYxwAqzHW6WjkcZnX
YBi+ppISua4HxfLJCzYlixRp1vkaa2xyKhsQ5GSzjm0eB8ULUxBLYEBW4uhO8uvm/Hg1G8dJGcTa
eAbz0Q6k2peIti3JLsA0UqvQ5j+CR4G8UgtdHmzfQ0d83bcHQ7sw4LUV9+rzzrNfEgdGXbaAQeRh
Kb5Z0wCAHqXM8SELO/6lj6wJpMPIAVoT/kcrlfeM1xwuAHLFojOFXm4GhE0u2svjweHJmJmOAU/U
IZ7Y3X12d5Av1MFZmTXiNDdfvJg+r8aieAs1kTGVX2ehubarsABSoi951amkwXGCL9eZJsbr2U6M
JGU0LdjBJnwgX20w4C/PgiknZ6Q0FcGUXxcw6duRMOrDprq3OVgeIXLJeDPh395NJV+9W/NLet2k
m2JYfmGh07nxkvQxuDJu7Z4BJLS2c9uIVN8yy1bvlD1eBXfrkboslrnMTDYmek4G/+WqNd3rtNzs
OW68dhNRYsqgILqfTNqJfVg7ZF01/ZvPzYCKZoPvwXdCmKQD1zdedVp+6YdPlkdy6YibBIWCWm5H
fYDLnxje4glTwjkpncLZhefurprnC+n5aErlOW2SNpg320/IskGPwic7EHO7GgVprBAOIPJiiV87
3VT9kzrpuFvYwL0m5P3Lv05kbhtfzKN3FIWeFQAEAe9cfdTZBdkr41V9xE86rQnvAy6FpsUm0pBL
gJ2BJ6wV/aBCx06GYpKtXYJthaTK7wzUr3m8xKNdyUDtrKY5r+IMuuA4XHBxdc8cI9vSt/du88Ug
usLYIfP1Xwven2c5dGFDiSHKNtb/siVA4AYFhuCi8nHevA9kVSWNxjictjzA+hnqSmORNDGd71Uc
HrLIa/k0sXEbn+ugvxn9wJWDRBIsUTBtSVhMfFRTrdO59p8ZM2a+K2K1W01KnDVU/QLqj4CO6Z8p
RPEatIqma+h8Zo9QRkZ1MT6ZGkg2JtrkO2UyoSkrrDTQcD6GumRAzWGkpyebvxXf6eRJXGp2Uv71
85PGBskbEWJMtm83b7+6avAGdXIDxylHmCoSuDTBNaYU44ijGt17NORr6LfRUQdDWRcGbztfDC0I
fL67Z8MhoTxk6zDWrun0mOuXYzueHtbf0/METWrWarX/Em6reiPM4EMuDSgk2oGUhnuURCoVo8St
eCCNpSyuxf1Xs+gjYLosIkcjpHzVk07cDu4B40qxnENC0eeiSXBCoYqokLDey+YO79/rMSzaZTXV
jelf9F5gw74h8n1/TjK3jetGp91/XYd0GmUMit+hg4BtCguGuWAVeyHT3OvNdfCDU6uiU5aVguwF
Xs4MdM8dhAD+u0IJ0HHVzx/+COipdRaRn+6wdScX+I0gguOjGlm4P8of/6ChkhcCy5alxb1x55sk
+4rBFETeI701ILWm9ltzXAvUS0ilGE6Knh7StHlu1vMSY4SNP46NvTkIe2xSpJVjjok+63GYzLOc
7vgJOlwXpTCbDFcC/Rf0xOe9LJGw8P58ny1H//EUjXfUT3rPcjzvgwMgz0VkxrSKSUjYSI4v0c3t
yXqwXC99BqpcT9sG90+FS6HSahkCh1zVHbD+UBqmythG4SvrmMqCe+4WODLYaGkOFUDLiMWnC1xt
N3AXNgxBYY3j8BkLsbna9Jl8DflfN9FIj7SGz+IDfvNEWWf3YcdnwZgK8bdi5embOcVCfrtrjJb2
8gPY9xT6k68ZpWLJmDzzTR3AXUy+KGMOF+kj8M7LM07NYNBY5WYALOG9Ewe8F8HpVdfkwLrq174R
bLMdgq7tvi5SSoPvYG0GXABXi6HDuZxVb38Qyc02Pxx1MNUCtL4i0tMsXqzpFBrsgXyxkDRlopHQ
byG1vfB8Ct13FglqfqWzJcTta62oeIZU1waM7u9LcMN+UHpzIGQ69qsglrlq/NQRzAZ0uanoUMxu
15Y6EkVD22VsuykwmeqSOnx3WuZBCQ6QhTLMieCTKv3p5FUBO83F/eucuQ8nTh6jIVSe3ybhmEIF
5mL5k7UmOWnFzwjaxl1hwNr/7uoicAabwOrK+gAi2yZL34kpS2Gyl788C8F1trvtCYCOmOxfO5rx
tpzfS3eFc0x+Ni3We8y5mFJd7+e+jMELZviSgJ1jr5uKPizTV7wR8pS3KkCpHBew3+A/otYeGYSn
Iv2PB7FPd56Jc1ARxm+tEhUj/FhcequYx0A+KneevdZF1YUbNSKbEDJV4cUMzTnPFJGOgSky0ysV
Uiz/EPwnUqZipCteU+61Mlr38d3tr8RSRKkL6zQpSK/FEyh1qJkRvKCiAA/nV77v+3AA9iIYp94f
NbCWyZ/fKEMjfwmR0NMHtgTjnsL4sxJIvlzYcgVx51tdxFXB4I6ajyBl0klCqbDioSL7okK6mgGu
6rNbrkKqOx2zSXa1c3vFQ2pu+diHBRtAkWlm/WRcDa/73RD/a+ImBMem0yvs/Udopwl4Wx/+Xlhv
miCbDGowrhR3KcCXUYxT/fSMRBZKUgg/qn9NQIphiLCF87Z1ifx/O5sPCzYEeqACHOmzRGS7C53v
VYd8SlBeOzroUkNByzS7hbNBdMb9tsnQ8Z1XmAKC4R/JQUdukBRMlSbG5IkvtpIdKga5iMXCJ0FD
GV/8CsX3KkWZ+MGeXXBZkyTAn84FR6ZQl6e9CuG36Xz+VenSU0m+mc6rUTJWz/uXMH+6gI10D2x2
SlQcIl3Sgo3TxU0ArdKaqmt67Pk6p3TCz7jLILHG7Wb61dqPv76XtxOxkbF1S3rdkr0BvLEmVlIe
NbRJCJ6kwnLKNaNM/OL8pwLEt6e3XwOL5WoCcA1Ooa9KJS3M/6i7B5kUf3C0/drz/vwFJRachzQv
Cg85Vrao7cwxMuzLI+mZUQIZOL1lt9pFvxd0PG0Hh8KmGP2ZJ9iN48DRUYKmmRkKgBeZmauvX0Ea
FdHy/bqj1uj69Vh/TV0qyHhqfsru2e2COleHAE6VeEAoBPDSF74r2f/Zvy+1xTg3Rdd+wAzhcF+q
PIR+2bA/f7PpcrNKAzCG3GACznAWMvjVZ20fKGGipaMwZSk5PvyUdrBQnA7jNvEq2/jdSOxxEdKG
pr9aDiySG/gSGn07QtG2q69a00iDYbeHPxJntWxBXEEuy9Bk7yfCbNiM3fU483apnmwsiGuzKxEl
USxcqMa7OiuOprElTDbQN3Ty1K8S1iuA4YnpCWI9ulXLoZMz+unFybWx0kclYSqho5U1w+mhAGFw
6T4rQjqOnXFVrHIXtF5Wyz83KG55sJ4iDPtvQqRDN8r22meVAXyIwAcbahn4xxFQR31vxNGBVyTI
Clj2kFn4GaWprCBSFSa2KIn5solwXqmPFJKN5TqVIEdL9tUYWart7HJt+kaHTGVHgP9eYJZ8OaBd
78gJJRgHj54Pjs8AnOCXtoOTnxQtCtZWF6cJL8tdFijCS//3xLnMFljOuh36wksCJgw4TvhoOCNU
p/uvkqN83bdK2JJlkPH0ISSP5bhbLHW1+XxWFCAiVJgPkyL7P9iHwvW4j946egUBnNzWBC4liKPD
xA3/8HRvqlBZY5a+fxKR+4TVx5WR8Ge4htP7hQP8BKNmE5NNvW8f4xBUzGw7CM5nApbpFSazmOGD
2AhakxP5ntJhoS/+XnJ4uzm9k0ykbZ+kUs3yZWhxayVAsXVhquOdE2W8LVberwt3g5CHEwac9BtN
6t9t4qHpxNHHOvroGuuMYdktbt10sCtSv/7WZRb3oJ50GFVxe4GSTuyEwhhl4tilqk2rGdhlWBZu
0xir8KrSNH4ThWz+z4WKSd8wL/ymMaD4k4Id6l/C6vO6LpSR6wujxPIc1vhC5gSBbogsIZmeCJCV
5E4oSS7mPc7jgQ0Jig4FCWZJmd2zPFo3uq+ZGEzK8FaAp92CCtOdqxxoqjHd3sQ9vB+yTLNvxed6
sMo49p82xPjQ37RdNDDgn2ifJ4/E/VaZPy9xotm9k9NGSCwk7zGR/VqNPHhqUoOvnybvFt53g1ln
DpwF4fnxmXcQmX++GImr/4dA3mIGUL0dT2s2bvQ1orEj+Rl184CYMCGks7sGtIrMZwDR+HelwkFK
zw2lANrtzzNbH5T7nThZBfMTOyi3RJoGq+Zv+OVnE5JbT1bCcPW/A+3S99sapzx5FqADo40Pruwv
+4hWWB1uUeETuBC4xrdksMDNmKWNLbRpxqYgrD4nIeZojIeGYskag68WwayoESTOcNUE6Xc1bXZL
MBs468dwkuQkaHtaH5Y4Zcidn3OBPl55aRcTDMkfI7+k/cHWIvMUaMov4sK62H7zVFcc+pRooUHR
zsN+9bg2RN1WpmEI94EbQPMkbMBG0m+eDNrHnlRiktk13k2tSh0wa+xkySGzXWeiX0NYgEZw90NS
zyj12LIjJDGSr8Oi0WYMhqjZM0nqlhRoPBHAbpRUielhp+b8bYUPlnoj/B/JB3yOly41ETU1c2B3
LNsQEQdWJjkDM/D/9CW3W6v7Cgz5sQbzuldgUu16cL4/VU6rAAvxESyGozGIsfjJdzG1h6Ry04t9
1NClYLcXgj0pUbW22McGAsRNRkiC3QFpnisZfSz1upLcvtWIZOxqA5E3Q30P5onw3ixuXP5cWQKW
MjeReWA7MvHiwapa4j5XP4FGnLk9KRt9TZPcdrp5I9AfrBP8rBY7OwhgrEgctvfWV/29vbz8nZOj
0/MoOOusjjXWgB8T8+rc4wdb99R+6d1O0Go+mW1CgM5mGUsOk/wu3K+7pLUBwdPwO7SLp94KVssc
jkDOM1pjy76U8Gjeg2GSDICl4t7ijh4HhBTWEvLVRN+E0oUwti3AI7fNaWl5DOehIgk7croYANfa
ilAe4DICuvivW/iwKBmdnfMICvkcSIEMuwfT/b24cOqaBs3RFHeijNzlygxMvFugGwabvaM+5xgv
pQRQV1YomOgHS0rii4ulW6jK/pTOTna70sHHJR7CBIZOVEl1SY/mWEmVrrOGsyNcTNBsV0QVXt6r
SwNH6MsGaAvOmHCvt5r+g6hEmemNR6OitGy4/O1LIJ/1E/4hRZchGODeupFM4A9//hS1Iv6AE6sG
6bCDOstlL2tjAqYSvFgvFzhLWBQ4BwqTBTpkqSQW9cOS6I2YuZZn4JN37+tYVYJ6DggcpmPJjd6g
SgNRNve4QhhTfEP/HmqpWp+prpR/3JtPuKcogJhhms8KhTwH4e4ojMA9+oY/TnLiwoL7+58h7obh
cWpVfA9JeXT2zt4OL+Bo2PG53BhCsOC+PjZJtuAsWdVzBz8eub7QPfuX/tc6NL4A2UIkqxHJDYy+
hRuOBXZmH3c+mMpnHRnAq4ArbzJWBXODGi0y/fbayNgxTCcm7B6p/Jbmsm0R3IF4WJ9Ry5GlFHvJ
sd8ayV3Mv97NqDH588Mt4KUv8suL8b8P8QPleIRzNp4ctTEguY+IRUdigWJjOn74Vu3ICzHolE4y
B6UER8fXvUDJ6lXcXwhS1BsofyUpYkIU4iMPC0rc7x+BeFX5ey1oTvyW8SV4Wvnf0tbuBz1KQIDP
+awnKtSsmRBMk3IwBf8ygQOP6zyBhVcn3pVgrv2qfCvfzWtDY2g5twRx8SmhcWSmwLtmJukTfXVD
p10JgG1950wbp4G8KbJ13/zTrb/I0qYcdylnw/V+1PHdhOkS1pA9ZYj8e/im2S64R4r9fMytetHx
Eeo74M9qxIMZANknJauakTkabvLX+s7EglIQ1Urria19B9LM1Q+zqL9moUshcfLCxqkcAqxzCRDS
3T4+xgEz8KpMXGX8r8CE7f9GdQhjYvypH1J08uXJCXUMUC2Tyuyv58M9RXhjbrYMaclyvukn5nX4
Uo/mQS7bjR/QZEiXiOq6osaPct1bd63AVMms+SG4xRcQKiJUNk2sdMb0gdo3uyBbpO7OZJU/F9mK
1rUR4dWJy6WsspZsUpuSoXk7PbHIKxurmX3fl+cq1KOIyrKgOUN7YNWz5W/vPSC4i0WNGuYjEPCI
/IEb40X9EReL+/SeY24b0SBk98geYp7mFEPaNWwwBs/OFu4qqpYcXLCYrXfQQAcaH8T8hhUhcDpZ
hL6pIN8l86tseDKEkjIp7vPhEa8N1lUMzf6XD52oIGS+7ePV8j06b+pBQJcRG/t38Ch8BREqX2DU
shLyrMUUm+8wGzVQXajMsghJGPLJ4oUoAzyEoPBSqK1KLpESyoKBu1uoUTKyAAw1opHWi6U9kcBg
6wJoLnSbKvqAPx3tP1MJotUg/bUReeT0Ip3YwCGM8/ptdaLVReUXjeJHr5cTIR0T6VKee54TjZSY
xVF1PnaO+P7hKAo522ut9sXxIaqGU30DSQrVMp+A1CxibJBcQdVXpJ2cA3Xk8o18x1qL5kaYr3Ek
a6f1XJfJw5znx3MRAVjhSrf3ULYAY9RpBpvraD8/+Mp2YQMosN8VWHk0unBIBEXrTAP48d6TG6Iz
zvNECQoLMrr0FUJlAJNXZj0mBXb3vPjOWfKYd55rpBSJ5qwc5ORBTfo9pRPGf7WQRfKX5uRa9HRs
2V1iRbZWmptoP3UaitFBPLssdgE/O90xsky4bPZC2GGtM8RAQjAkyLdfEPS7O9pqzB4ayNpxIv+c
QpNkhuZobchrJW4qW/h63kSlQ3dGN+SvA+w7Yyz1XuH21x83Vr+1uWCqfvfSGqOwMrjhmgpNApIP
rSVjSVlp62SCAFbC392i9JF7SMY+UIUOHYxzElA52vEbwzyLrn2s5MdGtfZoM3gTuTvl9NHdYT0C
QHAotGPq+XxWv1QhHQCI7zNQJW6ZUfaikuqBl84bu4qyt1SvKf13bKuI+pXOWy06nwS28cK/Em8f
PENiRlAd2ic7Knd78hzj0cWBD1U1P6mEWluoa/4KUfYKD6/N0UY2NX/f+icHKbvNrM/gII9QzJ7K
oGqayibX5nxounZn3dRINXjAKVLQFW8HxAksc7QAlpwoy9/hUrIpLB0Y3UJgebjqcG6X8Ouw/8xA
n9uUYK4KH+FV4mVykn5/1DlU43pRiYmEImDbOhwvspW6ZfqCrUphwJtzCb170Ppan4T5YrFQ93S3
kwQbH0DG5LgllzHU7RcxwrznWjcQch4lRc6c4qIsOlWLvumdFAhnmLj8CmP3gWqLpdOqAfpY7nTB
3dHy7WnrImUx3o4WaoLH/Sxh4pE6OLhJHQskkAbnQ3H8tTZ5PPPee3MEqIYZzH7Wfpj3ctXdYpjj
4ob2VQDPq7F8vaY7TTRirXZmmUKzt94ejOrrMlY5H9fYNJQPJVPbQbRQUQMiDa6OecwN9xYkuhxJ
ODOj7hpTytIAnjgOMGi/8y5lZ5SPUmlZLnQSHZ/RUhC0ViQwGlrY+fG7z8DdMAHJnwxwORlIZYT6
56Fsws6o+f7L0XBzJvRC39gf0Kwpo5FekTJDWKaC+/8h1fzXtV91cboP8gqmIhNBXmozr40iOC8F
4z58Nz9IKBpt4YKf6YMJJAc/6xwPWuM1aox9WGkwE0Bq/K9N53x9Auqlw4iZSKMf6z6P0GH4oswR
qHRgluMCNqqivJau01+U+YeD5W4Cefva+S1vY0k2jhf5u6Of8Fb1OjH3b1TpvfJ/XYglaSN15QRv
ihABrf769W6hKwlSy9wLkBnq1J4Un00AKrOZVqlhGxdiAniIMbQLl3ZVKEIxbSwwwTZIDqOsKEhb
iVpp3mQZL8I6p1DjwG6vf2hDsamjHCWlXeNgnbvfVgWZRNpuxht6XFobTQ4TIZTFR/8aGZ4Af7ql
/YdQP4ILKETP0uPbEKaxN/lST4f0IrGppWss0ysi5rKg0txizc06dEXGX7iIfdchPNCrd6NqXcHK
cCYjMBQuE9DqBkE1I445EYCIjlkruhyo2A/sRFQnsViNtCojsiftz76wWZExcihwVHK7zQiavLXo
yCetqc5YAFoGHdlN0kU0o/XksndbX6bsMEJO/n2vuPYGBcf9mA5wdIZgmtOfyxWXkbNP4cSAbj3C
XTjvmZkRngtPfiSDRpQcAW0qBCH5wNuYgDTLx7uFpEIkc1altne5pIBZDGly6GrdcIQ9IWKPITd9
4Ex4bh2mKWrdHYL+PWLtAEaIN6cSWQsfAsVLnQ1kanWqPdOdU9srCwIfK2MAFYNV/kF9dF6Ib75H
Q1u0voUn7g2QnYJT+FWsPEMmaWjDmmQC33Hex6bODJlhCdbctSLcxQECmiT9Nx4+RQ/IIoO0UiA+
t4AynLHkBD3GGqMYQATcQtD1xpoJbZ15oH3aEUMz8hJ3qu0BFtF8XgVzTExnXC4XSF688aoPiBmZ
vVhR/rOEA8uXtESV2WWcML7o2H3yTu/LQjEh0DxZ3iqjn9P2f+OO6oNd39cjOblWRF2oZrlK0GVK
BLJk9ffO03HaCpC9RYVyXOb5YADNBLt/C/JZdnzNlBjytvYUqi48WGDWqs8MSfBF8wfEg2l+W6z5
OUPmRFwnBdQL2e/4rq26ZHmuFFLH9+v4kOvMDYlWZTnIItK4lBojCbFlNUKwQVKoDc93Az1nm+Qt
UtDR0obkX1pUvaJ4Je24f1eB9zG9NqXBrMmRL8oWekXC6DUYoxpde49UKhop7OnczlXzbvgr8wkQ
ldYSMr3YUU0FamtrwoopKXuciB+kqMeBkA4L1y7N0c/jvkPizRgySAClJLpUpMLKpxcwjXbI8YwJ
s3uUEHDYdVH+06/Nkq1+LtTRh64uNzOYJ7JgYe5SCYxCO2j+VfHnO2v48AzFk2SfLRtgOcVAAzcr
jzzXWsNQ92i55j8jK8j4jfgolOPiEhIcSzQJgwNbZXrRPD6jLJXxKlVxY4fz/l7EXLfc6uag8RM7
tb6z2BHXb2isrCG0ATPe97GhLoGp9eW5Vda6E/f+fJe8tHAds3TyN9sdVfG+kALAk4c0kB6Xd7xO
kLHwyBLXSxSehG1Sj6VYhdpBeZODj7V/Fr0+tsd+igxh4CNaWJvIxlIBISfw5GFC17aJB29VEoXW
GzqhHD5Z1/TMHhAwLbaVIk6UPOJNayoxBFGc2SNFTlU8+dLPnyVUCDtpHJ3pK+Gpcj4z8AUO4nsa
Xb8FgVxGl48v/XisiH3eOsXcWlj4pAWnURGnvKst1or1DlnnMzilghacY84QoAfE4sbbSPgVveyc
xw+lQkNrlsldP0xWMXXu1gjCLzhW9T7EgOpUcaK3I37wBVO7edKHvP74QQuQI2SdS5xC2ZKDQhVv
BQBjmm8wSeHhFLl1QOV7+XqZQ2484922vZUGTb9HN1nAdYM8MjuPl189D4p13eETFBYe0hJ99lAE
dlPxVzkJ2TPGiV2Zc3S+cFtWhv5J96TZDqP++Klfhv9J2bPa1WXdrPOAsyuUVagpPxsckS3g74HT
irE+R57ODn0ZowE8HoI8oc5cAon0KRRr43wOQhsEHu4Z544mRz2OKE01FsUZhqdnLCde4YmZ7Kb3
N57eFVk1ZY5uJF+VglakZP2JEey94LLyHHiMTfYWyIldKQoWw0s1QIITxIMeXbeUjdTLEwsUuY+A
ZvTWu67wjl0RAQzHWRKd4MrM1DUVrSP5y+4e6sat85PS+9M+Vx7mGNawwitSGyp36oian08TRPj+
R06bRMWiCHQQ+BxF4WKoWuPxY52FUyV7/CeGD+q7/WwK0HyM8YroigOueuYLJoSKILpuqXLiT73D
GZPQlxhmQrfRuD9iDkZaW7OoERvMeVKVXceiA0huJluOZs1CGAdWYPeVr/xSRQqLWmV/S4u9FkSR
x75v74Ar3PJMYjBal8atXvY/ccHHHxIR46S6rr+j/NHHOuDRkrqD0wFRF01Rf1CDVFXU0kLhVui7
KDaouDKl1R6IVnMO0x7inCJW9AAiC0iNcXJs5p+9lUPsXDMCuIib5Ov9cKJEJKwk5pt7jrzP4n35
gK/aTcXr3qH8Ko9XjmTEYD2Fc6DQQqPayZ/Z4woO06hxaj5EOlJS4WPKoBNUz0Na/iJh6LKaJior
m+WQu+gQhQnO7gKt4STeotB/uyd3Uc7/BSA2j6xXjfdA5ST7yENHcDGYKKeXhHmDTJruBAkrzgER
NSgc6OBql5ZMnzFsHon1qF3kJNrVZ6PiLa832YrkPjqS77quhrpYlBbX2TUfrZLvRnl9wwsnowhE
Fv0sX+IoWvoS5Cn5ERZNRnIxbxT4O57e1EuVtjDLQ2AZNZOzTVvdJCW/TJg/IH118OJIG1V+OIe5
57O9lrdAlNRs9HbiYM1tsr86USOIw5gYuHqDXTjdMYRhMF8pCkcHC98McikZxXfvsOAdEKQYkSad
CrxD/hPQWMAZNJc1Dgju1lhADR94T2eciLlxsUskSqljSXFavZE6tLD0CtPDkQFSQDa41miP0hiA
3TGMWVW0CZhgKg8C0H7ZDdOewrQAd5VUn/wbDsv03Bvpy2hAGBYeNHLqThJgCV+tE4X3Tt/RsEGU
VD16clLhEheENvkdDeVvWXeaH3gJGotblwYUxaktABrLI2BbA+bAHZRRZ2/iDw3Y5+e2YktlK7Qr
SlE6bx9PU8yyUFvN1GbpZuf+zMATWHaHKFbdwUapz9fUqB5E7ijOJf5tU8GMCZNL/g8kE1qS4CD7
Vedj15mufA29Ken5VzbTB3rKqlsnoSR9ieq3z6g8V7X788UA9xjDImTxs0qxJ0TWmCuk6OOfDqGE
s25Jnga12m2mWPunNjc/WLbchPy8MUKS5FwVTL4+gHKKF+4EJgXkV1iWljhx6hwBbHanxhce14kc
K179v1JTB0exg8eBC59/hpR1JUcP7eZ1rhAg9+FMZ3niFsI5oWS502ri24X5GT8OeWDi5+hkuWV/
q2e4NiG9VTpmGF1uwDsa0olKS0Tg+eMlxh7+XH04mf2LCRSuJSuMZMTXUHIibZq/kFzU0cv5bzmd
nODKz53vvR8uo0pa2vC/6Bbq1hGcLbcR5nsWXSIh09A+4JDsJqjFbHYUpI+u3tZQqmS4lEYc+SZB
tLmHTvoW0khFaQDtG18NKO/9PBsqzsN+MLTnNd7flyXF8PD+IPNsKAFHHpbZMt2PGzuwa5fwbZgl
8HCzfEcCWXBkyV2VDnPpnH2nOPB3FewUucSsvdYOqDoKkjIhrIa5YWX5mmZ9ZtO2P4930LkdK9uJ
CCOlms/o6Gb4NnJdA7VQp0/1GEBQZcBoFBTbIIu/uuAeaPUze9sL0sflb5pJBXck15Lg/uKyVmEZ
hAvtRbAHupZBOJnKBZWaqqrjHiaA2XlF5SahvkRfkdB8BIYg1+HuAu1dtxbjwEmW7rmvZAInIh4c
8tZCRStdV8tmzN6KV+fCWTVqQir8UNDc+n3A4uHZn9j3u89ownwnfmpBQCnemywUfqaHrKvWMxgi
CmXJYOcRAmRqpcCvYM8crOwi2X6oUykcPjBCJOQJhTOilzYxRJ3BGs4Bqd2kYkricLt+rdKRhALU
K5hF0cV5k9WxgrKH6IhBcbgN4RIqiTrbxfqkAtBezWSyde5jK7MFX3kIvXeWvvBNpGzcdbX2Nrrt
mf+OhxJJdzFJbJ+q73eyWn8tY7zRe/kob4D15EbO2wSe4Ht0AkCEEoG0LxeWSQEWkfav8WgfXfvw
HSdNwW2if1Ah7l/d3vxub6c62RussmSshYQDiuc12Nsl1PwpCX2rTVmfNXgXpJ5FrlmlLzBPUlPu
CrLj9dEFPIKZqE2oVrJ3uIiHDqNOToLIHlO5vsFyOQF0+m4Y6j3EcsOQP/Vkm7iIGQ5AZwwft34n
keml3LG/4S1HrtkkLNaWA64GqCBJIP0pcmleZ48e1mde4ndDLfXvNiZwzXB4TF9zBas3Ln4mr0dL
3GLrEGI2iF01VK+8kYv6iKJAPpfPkEZUMvrUXG1S8EG5PrmEHqX23uS3994okSZdKDTbsTyoaWv+
UI3GuoDsrpNLEFT533C/FOAjC+7qqyVL54Apw9dbBO/DgniW9VXyxxdLlG9G6qIZHf2MJC0ICqL1
dY1Pvkki4ITMAap5mmzS75Wti+88qjR2IOxNfj7bB8oMEf6LwzKyZwG85oz1Q7NFvFBp7OlpRmv7
RKaCK9cBS7RIAHHfYohfdqMPA9TaLewhZ8PNzP71L/PPbJdBZOCEyyIkajuJAYeoLZMD0DMGthYP
zAhffrFWCpiijyJqpZyVUqgnpD4T52VOZpX//ibKkmu7MGCwWYP75eSnyoLv2EaJnS6dE+8ST/5b
hHZ9hOabL6xCppPm1wlCl+ZNcY+haiiKn1BhMJ1OQJr82D/E2fMYk+vVFSxzJvoE8wniW5fo8aIl
zrCkXgBCTBb4/3ir3KeLWbwEibBg/G2IL7aLTLllY+iQFghyqWAcUlBK9BDkvXoDqifm7t6wg6QR
4XK2UIvadrEVtai3gmLta8h81xrxEeuW8wMqb5IAqLusBRPwEFTzvqYpduDBB2MRBxeb3qoH+NaS
w+HNHowIi8xXACGDFdUh8AYT/65vsIE6pesQRSGpzWGcOeXOUNrkPHZDsLWctkWWBjY2rLtARNbS
+JcEc62OkvBy++T2eRs169Sg47GEE0Lk6O+1nSlaO5UtHEQPaApJq4C2a0IfWQRAHo9K8GmXmbbY
NYzF3iB68xwysVGHYQN8WzOPz1a0km+mLpD/PfGklHru9SnKvT7uqePD7Ze7xHoAAMyJIfIFpWK8
U5JpnV7EiFraibJi17Mv59j1tFdsuNL09J+AILiQXU5YfSNOrGvlzUGdOoZHsoNOhs9/VT9MFgwe
tBoY76SvQZtQ+3of6Xm9PjidfENgyEEp1y1ebdnzfOo7ojfbpKEm2DphEi6PizciRerw+GRLGx0G
D0f50YHxMbk8BHCnhN3miz0GYOeInKqWmqTshHneIG13dDPo8zxETbtSlNFIwJaUF89AGt12ebDR
XfPEJ2DKr0SiqgqNoTdk634gV4VusY3mOKgSs2Rpvw9lpwavQCOztYkWj62qG3SuV2y/Tn50nwzt
4fc4HL67TlN75gX6an3FZ1xaH8/rBQRbDMcuDQes9MGNtQKCM8NHIUxC4szN/Klc3XhfOU/VKnPw
/jSJPKc6+7e4bgh6HXK0gHSanI4ceVD3CtWiZYcr1DbawBK9Dy54Xjgap0lUtFdxmEtyvQVCsPlg
w1RhrilzEf2Fg1kWcIXN5PsX0h842iREu6DawUqheR4bPPqvgxuoj/sfLPooYjR9g2cMm1ECLFEC
SROLfAz/exLeOSgQ+/Wk4l8ctSH2n9L9Ig4KGJghCCn/Scc/r+NN2O1XkdYTvxX6+pZX5PCxK4Mx
SNGypaDoabh2dSaipC5LVdI6t8u4BK1bILdzoRZU85gKdD9GP4ZYYKwLZgrRWUAeyXDg+AI6pb5R
HQPDgLeQf3FYMsu/eoM7vjh2cPsCQnSI/EWnyMG/98CEtsVKO+i7chwSWkjShM1NyTsS+B2I8Oda
fAcz0R/jSk6auejk2HtZkjUEBfps7l7dppsgb8qTLap4+dOB7pxmK9lYanW1gtUCHUlRcc97qolx
eI3BEnhCNXYH1ZY9etNuQAo4pe7W8pNQ61wePh1aVpGXrPTVleEV+R651j1qzbRBMyBkjxLMLGpK
Tag3L2JLT5dP2y+zHwydUGwwYwXx4u5dLELF9o+3iNs1XC64OZh90ObusKTBjI+C5jwwZ/izdwnK
Po1JJy8RnFb+QlnXSslZJhmMrvXLk3aqUkJUAKVqbgNgaJXTmV+D377kpAUf0fDaa7a1kwB2oUF8
Rd5d2KqSqnM/QPGCIwovGIrYCKfYNQ9mNwZ0Es4RGKeBDdb8KHg3HCkskEYJLb3NsXgZQOonbjy1
SONkfbRi58VTtNJzRQrTShWSvg2jpFVh3QnQAHZWhHwE0dc0/Zcytxi2rRfYowCVhANqjpax9I3b
+Nfsk0E0JmTS/No5JL3WqIJgBLMD6AsEMb5g8qimbGdyusvbiHk2Zk83/bHm2rxLS95zW1+Vj1IF
g9LigWWrPpgYPK4b7TnjGKb5sauTMmD6ssVsVxFUTeeXeiTApmLKC6p5svoig2Wkmp8XjsEkirQj
e8Ll/YeZ4DL3u3VW/dF8lU2kWJibD8nleirLEywHbKlmHExmpCqkkGGagnBS6IuOIAmwJUU/kY2l
3MbPevSdlZlYPx7zynTDrg1EHhWYCuYcLTxKXegr/LHygHOlYhy7oLC6Cwf7PFXVAqr745Ld6kWB
/7/HGcR+xPRUgFW+sm+6ARgT7nYrBk452xC5cYByqskD/niG2RIOVK8oGcvHNZrQbisppYQWpEKZ
3qPhnIk8K+3NhiJg57l4noUdTF++Ofyfpb/jGw2GUX9xOyBzF9CMWTJMmm3zWw2E6ftMywhsZcIT
8ukbJ5rm26I5359d8S3nDubX4PqrlKckFTKdNBekVB+eXYDq65h5BkPyr1CQkyLfq65kj13IpPxC
M4GhYpqXAZ1JGzELLk3/41KzGFLilPeapj6J7/wbtWYdY6/DWLN3KS/AhIhjuOnFPs3+bRbxkxbw
8qCbsxsZr1AyXW+y9ikyIfilhZSxbFvrQeoGQIR9fQQED7TISSMspl5ZcEupQmV9o86eV0xWv3IG
GKO/b2rgpYtcUXDyVbUWvFRcUFo87mZvJwSn38NH5+SRJzhiJGdcSCWW5WijxQYHd6DYb/zjXKO7
TGTKanEH3eieWl8eYJ0OCVIa6WJcqmw2qmchQUa2w/MmVB+t3jCAXczK7vrkaVPSU5HdqPfI+z66
9S6chp6B6UMz0j4Us09QdiZKMNmai0U7/VpQRFJK6w943OQcYSt4wcQpRQJ8X08qk/cMnna2bk0B
hcWnF+0qDRLzDMaC8n2NZc4FhqSG3h8G6OUmzHeH9N/RzdaYF6/hDe6UHQJClxaGXG902wuRp1OW
kvf/YJdPcPdE0GhQ+35K6JjpF6BHsAfWv2UTFmVxglWAiCuoNWqiM9UNwLKd/0AgNv6aSc180Hbp
2xzMYPCehLDeVkZhrIqAKulPBQlWgFsnQOou/UXIaObKP6boHcS+PmMPMO3iw8irWgzVPsQOZwoF
W9sl3ZZPr/3F5YDVs3KmQabgvS9id8tvf1f6JWfDOE717qB6rjf4CO/erDCnqcaxSzhIKBQotYFL
AhButgi5P68MF+pSVJyK0Qk2+ZGmTfP8F5vizbg2j4G3IbHr6tx0TOX+7b6UwB8uYSJ6DW+Mppu4
I2kPllBhBBaAFjQXvKuOpaa954zD3hLk060DnqPJ8Ss32jrebC88/XCXYVGhwHKk/+LdWIQZspXu
o4pufLDGiRU91wbB4IDUvpGgKUdDO/PLaWxdyTWVO76L2nKpSkqxT8c/n1I97bzFvrRQoNnXHOfj
VD4P2vcygLFiMmcWTsUS//6f47vU0cReIicgLGeLQPZeeikIeZitXUQNsZnhiTB0d0nS1C0TsykL
IBItNkR7V4HCvup/fNafqNsDQ0Oz2TzdrYZaSvt2S0Ah1FURwzkq3EwU2HHcNZnXSZgMMkKzriR2
uSamXjM9uWtUvNSd122ksZvp0xGbaQa6mZ0F00S2QzypfhdHbTD7CX+V3Ig1uvFwuZ/xHr02d4+H
ZvMM17y4PTLEpo0zZ+i8WHWJqz3D83rmw2UoDm1jCeW8ymJ25aE1/u2QaBvZJwzt3yXW9OCuFEdC
MwS33Hn6vrd34sYQ8QBvDjptvltcQoIBzXmw5P6873ymN6IoFR8AhpagGobPL7UVhseSyHnHUmAb
/TySfOWWbKL9R33RGVFkg/+J5OAMYIIN8356z0heB9BeUiqAbN6s2JkZAT2bM7/8Sec2BwaUXyeT
p+mh0xyAgK7Ucu8Hok6WyvgJPfRGQ0c9cGghDIe3thacAcLd81jSB0V20IAHmXHcwVCFx/VCxl/s
KeQSYa8Lzufy9pfShQHX8tjYcqm1WZSxC0TVAIei0kEklXtAJ4+R19mSWwWAOC8vOcda7cP+YiHQ
vEFnkZKuyfoRnLwVnxGwgGuVW9v0DQt7DSz+PLtGnsz2IyNNSMMHsKnhXSTT+6CTbraGAcknn+r/
y1hTDBebeAc3i5E2dZoEMLUadEa3gNjK4W2iBdyxmwTx0pJnse1jRG+SnKNtecGdr7bibN1l2uPf
8Jb7xO1uESI7tKCtzvlHFYoAJuT4kDwJhQ5Cc+xNeL0kEtAre/fiep3lpaqRG3eC1kpAI0H7jmtr
6aOgY7Xkn0ciOTZfZIRxYnRw5/Dq8EkQXnUIJr/En7yRzB9ys2dKwpyT/lO0g5oSDLxSYGsSpaDL
YLRo9yDUnBXQ1cev1rx5dF70WBsqLXBkCAyzUdK7f2tFUONtnRK2uWSSpOnpbKJam6EsB9phGLmv
yFTehWtgpr+dLgw7cE5yy4CutQZUNixRY8gtYoni1eF1HsEq9V//xn9RmKG/IEeuOOEIqryTnqt2
wMsGGIBov19Kyfzh/sQQ4Ovis82YDFqOP+ydONy7QmyPtr4hwvVN58fnYQ8XTsew116TGAkFkiI+
3YXXlKbtWM+aiMVm1oKE365DBIisq+S2v/w5n9Es0xyT8XtsrAvdn4fnijkfhMWDkY6tf5PqsWjR
XOru2vyFIBjBHf7A6ym8p45zBqfOdidcl+G+Zp1FNfmxd3cghRx8ObvK39q7OdNHL6BWO7qTpM5c
kTOXSUH0oE+dhulI+UnrC7f53NA/efZvLiAOztn04sY9vKJ/Gg+qcSvtOuvEaXEOZl3RSKclIE8M
tWKz5npYRlbZL++60S0Vh+geBPs3eYv9qEapuau1AQ/c9Zc0M99ekQZayVNS30aprzMPdiBbh5Jd
nH1yLh80dAgitnefQc49G4C9jvMk4iVOyZ/Vu8iODUv9ffVp7SZ1PHCglRLxyiR67csiLVQALRnd
4wwiE6P9lF2E2S5llQtbfNu0tBjsm3qTX73nHJfbLvKoIqTOEfwObm41AxhCYtT1eonKRa3bTaz3
QUuX2xyNh/s659oRTazcOn2zKYn32XLbSoljSLxGNzOFUR8m1ALIBdH2TrX7DQk4mIMhXCAsSwF8
3pVfXIs7PvWLP/SKOj0+GxpqJ5peITyjsC1KTgLblJ7gaTcRJXUmc7oGwXhIwZuYyMhgWu4BWsn9
90A3o1k0xTBayZxjaFFy3DSIYOAiFVRblqoYnH3sZN2yTY5a/liIB7WcdnDBd7cKyENvGsErw+j1
1BeAsR8a8sVeqtMydS+WwUgD4r0TFzga/EBmx46D+hwysApyKULM5Z2S0Fhg2ecOIoVMvNLXA4dK
CA3RAkXm6G/soSzwgD4uYqYEYpqPiMFTpP2CdXwunasnn3CtZvqydJZxV/GOu6EfSWAW3zX2Rm7U
kl5r6gHpRBfA+1xRucUX/6hFECO3zKqsUkyCySdUsUmZwzRmMOylmmc8JI+YEA6vtTRfnJfItv+r
/mQZw4Gc+kj+sJRgAKPqwH9cv4tan65AHJR8QuUeAK94Q7u3qm2rwmZfoEUtB2vMwj7DoG6c8T8j
dcn41QMcXDhe46uO9KTmyH0lHILS3yl1gux64XvA4uSvQ+h8UMFmGMCMuuvDK/LJr5tEBf6JrDQ/
GiKNDbhXM3tagdl4uqoN3XxdfXiKaoXQpdgaBBSSk6HWZuVE3NmNi4TBao6eXzadpUkUvk4xXsYC
iEBZRlR9lrkZ7DmGvPv6AUNoOB93WiHz3rLclP/NQSOdtpiTTtXJF/1yPlOt8AOdrxbRXAuIVsSZ
7aiWYOEQZwa+OGC+T6ZaB3qhaXiVgc33RV6/ppEK6mJP0YoyumY6Utozr0LLPYuYZ8JmynMSZ9nW
DE/EF9Z50M4ZKb7DKIoScl7woNWlMhrDfAsrPNHOjz84OpMCozqSsOrituYC64Bi2rcvE5nLaOaI
nriBrBQ3db/RQO0mht0LlhoPoesC0lhLL2U6bzzruEiHTVJuOSH/Q/hN4V2DPh4Q43Q462iB68ck
rdz6LQfytIPzMpL8jvIDTZz6uzP4pdh06+ZnmxuhEU+70pR5t3MZE38rrmC7y655kmRnLEcbOScR
+Tan4HVp28eeiqXnTfc+Ip7Uq8JeK+DK0U39tQfEZNQT71HMy4cY//niXPtTl9/w4Z+RVZGNeQ1z
Dgg2wLSCJ37PMX6nUCmysnO2IqQLZwYOgMJ8bDdWevUPLR/8HXYkObO81mLa3B+w9F2H5xgLi5zi
o3zuJt9rqJ90yqF1C6XRH0M45XSs4iYFs8CHfxDpBty8uh9A/InKOcgofauA9HH1YDmlmSK03ZNU
NBkxgYJvLvONQlklwc8jbC2GQtJi4AMERuY2C+QGAsCtDWeEE+Dh8l8wlpZCxci/AJZbWYw2KOMK
Gy68VjaxIQvlimjaVGOMkzqsaqZ5LJsyRJGYgPhW4HtdxMk0GRtOFvjS2Y0f8gsl8WKvkUGMboll
/K+VD+aCiczys5vofW2XeSQl8U+5cViUNGLepefp5SNUXCdEQg+p909jxlzrdSBq1gNFQ5vZbPlh
IXEpVAVIpBzacyN2MEZp6yP9cuMO7Lqiba6dljWOZ7M75+tWZay7Z+3n5XUhqFkP+g0nnmv1isOG
/fcXQrFi1vKjIXuQX5GOkFPWvoPv6PEcnm+n8Ic8hO9P6eG7835EpgdtdC+RwawkNrgD/mgEmLgx
bx9LqmzO9KHcER+6Chha00CqYnhqEobeoxRp4jv4mzymX3xAvoS2Iz9OsFuCaZHEpwq4DphIGDyI
SMc5Jj5NKTeEIymXwFzBFmymwi3dv0cXNGroJL7Mmq3FzlxDfEIzxNWhYCEplgz6Pz+kRtgsEFv6
jvUFOZfj1RR1811lcfdq7h9fsig79xZSkH2Sncon98m5jmb7DJupgCWhDzh0EQjtBGtyNaBDWjOk
6QU3kJL2qIlHZFl/yG07xfPJk/krdt02jqm7doM+pJZFPWUqQCmFmtRSBhBEmmGKtiytG+ZZa0W4
wZ3xpsLnqnNcCcOVnoprZsUMW42yrankQ6mNYYcIQVtIWbAqxi7aMgqba+yZpB+kiD1A13pHRxcF
BI1nJA1ZKf0usrrTu12QrKXqatt3QG8AYx/qyIXQSmJt7+jlSq1K5lvieWPsXVds1OLJjw402OmM
K3QLcybdu/3YEv5LWHdLx8AXOIJNbXxXZtrz3qKi4k6LgpXOPnZ2ba/SjStgDsDA5w2MCtibP/4P
2+AEqmLEWghs1OBA5lAnsvC5vJmps66Cykl78P6ze4r/KY2FIz9Y2Cg3BoJi5KlkxBlMc6FCR+Wl
ec2d9+TN9jIMudkzs/2FjqPzX/rMEjm7QUwZgzZJMLsK8f1jW88Lfkh2n92i5H+F1Nbu+GfmJu1g
yoTlIBdmVDdXUCdxSi1O4pDfxd94QFnPst1m/kSnLMpWDlsztrx2eVzP7q/O1bmoTXJXQQZ7O/GM
jiRd0uVTeEUOVoEQOfFsuabw5QUnQgaFHCNxM8OFARy2OinoHmerdYxFFPMkArw6XLmuZZpABHe5
+YoToNi15gaSJgGVzCF9gFmpfuw6oKL52HZ0//Qs7YuPaEF0qVBWbQmPh8iamGnKDol4r48vjIUC
VaH/gJO+pDwnQ0PKRf+kCi7jI0XqDmv15dAqdfDn3E/ZqJfoNFprVS0JgqQcaTXo1FdPb36u6/fz
hbLnVsPR8hf5gCx7DxwAQsUREoqJoWpN6ds2NlPdCXjuuRSyY5kkzErK8y9nqyqr/haOkKdyDr2d
jrCA1xod6/L+MXJmSb4CWn/FImUQPhPg2MmGnfvFVx2Oo4TDABvGFX5hZVr9YVvGJePQxfsQBimP
Mp3Oh5w5/AwstHymDiCXgXzuF47nOwS71yfoEb1Qm/7QXG7zR8ZMYGB9s8ilCivoX7VMUItAyZs4
6SgVJskYiHsvA7XNNAamtcnyRYDYzI7IeTen4XaUkVALnJzYVbNtHpnyz57lgbrwdt00bS9745Yg
Y/JfUiU6VCKEHAd7ifnyVN6DnV4eo5gyJReQNKyx28bfDAtn7iIPlhHxMkwzYcW0sG/tAQP+m/Og
VQLs5tSeHCpoLnY5A2wqPh3Fsjw6JUsc/HC2tqkutky5HxC0YAhAE8YZ4fuzxzkx31ofLneEWpvV
ziqZ7e0UB6bIzwokygLO3HgBnED9cl3kAU6/njsKY0CmDr6EyLiNFrjRe5lB+P+gL3tDWcNMzsk/
yAEBiH354MXERKkpXeFvnMOq0AhoAqVdA/pEQjKip03DGOGYx7nophFmHzJXqn9N8UGsEP8qTRmo
vAWCMPXaRoy+Y3OFKKboUH8rTaV0/W5yGNd/1LtePLpPE2QJh5j8oku6hScB4uiW5A62qFIqm2Gy
iuYTeNe7xolFaCgZ3kltdvJP5g5ZnZxin2aF+JGkLg7ECHX8+tvFJnnWVAaSnNFF9ii5NmpbEeWY
DRE9vrqLxLFo/SzGLHKPQkl67bh/dtgtR+3qHwcRB8l6QFVC71eymPyycNkMS7s6qpa2C3WBLmjh
FA3rScyRLnvWCHHpduPl1HI8wfLDjCBo+vmDBmmFRKZ7SvFzdRyvOlwC8zDNzGYRgXy1nXhTAKuh
IqvnVBUg1Aw5TscZFX8Oj8AaPollnFARcWvZvxXFLkEVCqFfNgUtUwq8UHYbzgnhzwcsVpQ/4btm
H+Z7+WV2xgdnH8O3mhhuzNnKhvJkIHP7xX4a6IK7mT/bnDtz28KH1Sueb5EZ47qbi/6rOUYiHG6U
Zwu+nrpRE/x9VTO+zxwBTa/SJNrJOdW3DIwzZH9r9gk/XhQil/myo+W4Fden6FcZAwWkmYcxElTc
3y7UkC1zGnTtiGKPAet3ukAz1Y97esN78TsYnS4Ufrk/SS6/30LPlRC08NLRxfpWeiUJwEHjsYIY
+M00luQbQpol9+jU0FpzWK/0sLCKwD1IvN0MULZwdd5sVE5KKLREeXinwpRonCsYjTjt5Ze8v+dS
ji8VNhdz58Q+VN6pJIFGR0ywLr2XM2uOocHAillsqrEXISFIsrhftMgUbcGb3eyYVg5E0QEki7ZU
nEecmBtJq0w5bQw4HtpVpo7LwVQ6cCQHQRZwA1fQG9UsTJQ3QhrvYPBQq98vpK0XvyTwkp4Sx4fb
ekWqjsgCtW9PB4Wy7PBmu+fb4GJnmbbQIHHTCxg77oycgH+1QyYkz9whbKr22hRkSg2x3TgmY0ys
49/XrXiu0VaPph3uhD2NSAPFRmkC2dRSIhM86uzvqi8WAB+Wa+xXfavzs4GePK9s02utbvxcn0C/
JyQmMFoeNMXYOEt3uIXeTm8XLGrO6Z8Fay6LNPmzIlm1UZS6s20nxJ7rWuLFc2/IwojbZj6oQAAd
ylnMtBv9l1o8am6IHkT92jhDOweJvzhVZT/n9qBqX0UDqP+Zdvw8TzwtcpFGCmHByK+ohxgIpi7N
OH1bvS+Rt/JFn2dgsOjfkL90AcQ1JQMHVAutgFlwHAYs5PTnu3Lf2iMI0HM3WpxqnfamL7e8PL9R
SIZLMWY6Ud4tSMu+R95wTAhgkNxSUtJnFLZfQ/atMHVkPLyr714q0eKQmvZ+Q+sdYQDuSUExaQWn
HOX88Kjy2/pUIjwY04W/+ZlTeVxbTI/7PTiMKNSzS/MvWVuuU4fa0K4EW7cEmCmbm5Po98h8GQXV
sVx7thw4ZE5WxbITgshChjqeFoHlNgpqHebIltx5Ys1VgWPx+dw0ncO0ppgSkM357ZVgzisAOTQg
FSWlkGgOOOzqaGqwQI5ZtqkTVeDvbUmDufM5xii1Sxcdt6fkzwlJj2GfkqpCkLPHrbeQzV2CCWHF
NG1hBTA9dE8jP5ebGI/K2A4uSBrQzNcg/SJ9DICqxGoDENS1D7e2az67whfoyVDV9uD73s64u36H
c6JxKiSDz3/SjcOisLfMmUTgnmUfAln2a4ZT3AooHYyTk8TwwmEPo+1Hgpq88+PQcTaLwX8FzIS9
AMdCeSwYs5HI8+lrzNMhG9Wgxyqt0SHdFbbs2c9Kk5b6mSyw6kGIRlxVCOqsuASf774eBu1AtAWG
sFbMTNaiNkc5jifrUMiHs1zPT80z4SivJydXifGztyA27GZdyKBzauAUaUmDu9Fv3O53SDegrQGu
nILKLPYEMRVPCDGdWOMQ1KUVwLf+S5rD8Ru5jVbGCUh0eb5eWS20c8z4w5vB7sS/8WDlXa/sBZoR
/NcetOTSb/2GFGxL145EiSZ/vvMmdN3cau42+0Blb2zJy6yv9yPaDuCb5Wt12o9WgntGOecr2mgo
PTCPcJ/8cKc6OQJZRNxBiPGXtVaJaMZlSF3nBl1r6D7qcUEoTy2ZW+QFdq91UzrnZC8nCpQ4FHa+
14Ih5Q9FdbmGE+h5AxyhNOlKyZYdXz5zYhui4aPGvUw6vEwhf7SWH+8vPVMSFIQZ+4rtGPs2AADR
00fFOjLHdrFq3HZQVgpFagntz2Q+b7CfsScPaKqHTCBzuKue0NDNHag4nVmOhBtWLmMpXJ9E2dej
Px/L9baUM78GDgYJ/9vBnY1+tdtGRNLt3kXzOx2yf2tzKQbP+z7IBbvHRGa7FkZco/HO9vrOCTiu
siqkVyMKWb6xRQrIgguxcIPskV8RwtEykpVwXfa8Bzb7egA4B0pT+x0/Az+EZjKN0ibJZ85u+UB5
Cv9pdXjdqUtRmcdC14ygxHLmRqVLYgE34w0Qd2Fx0kQpKo2vdSUN3NBNm6FJ8HjHbE27edAeQpKN
pm5TdtRRXaGEzhaROTnF5B3zgoGA0e3nCmcPZZ1rAu7sl2GEOriQXFOv/7skpwkIyCyirzTKWvp4
aYU5en1TLkNul0rc+8zDXpryMwedMMuxvcWrzX6jX2qtcgFA0zcnGsXY+VbsGs6dh2F1JbsaSRKO
GFm3E0mlXNutaqNZ6bJVM2cINhKafqKgNilo3GWD6bOT1y9F41VdC4k6MGUQPRnGhSJ8g69u9AMO
3aukzUmkBNXDpPmKnJMiSAa8ofISbAA9nokbm4es/dL79Cchh0v1DgUUUMZ/HKCIk++Nmr/0crcp
pga21VjBADirnDptBIHDi/XxYsi5TQFDHDCZxwrAf8FczXwW69W+Wd3sVk75n3o5ZHqIbYDUrJ4D
ogpoUOGExuLED3hYIr2flDMvxdislfo+K1Zi24fcwDBlcbJTf3WpDWUCaFtCXQmomZm9faSjkoK/
QR40Ld+QY3L7HFWKH9KlIPrcYT9ztvUWnbACARgBWXRR8I4OxgI5N6U4fjVOFKyiYXOd+zxQydPd
oX7mAEpZIhgUBlkh6xHt4hvWq+vQf27hnfpNOCOzZvFrekZpQBZTgk8557iMlIb3QlqQs/fWdfJD
fN3Ym9CnqHfsJmyVXm0xIXAup5r1ejcPql122B+xmJ7YXirCPRPbXXcryl04VYxsyg3TYiwDzVVM
SA6cRW2zPGN3w784ZD6+acn9aIz98P+Pz8SZ06f9zLaa3K53Af7351Hq10mDvfHFDkojm2cg3KKc
U5YrNdCXcLYNcph7JOKhbO/YNOTqUDpj7IWZMarm2Nl3MJOCu+lm5eBtnJWnt2neUrEh8ynkNQJe
P5xbG8aO6hSoX+y55Q0Hk6+4NvGf8bVEr4vPO5y7qDntk/XCWRzdvDMfYslj6SSwt2QoqvQeljr4
Gi1cQPEV/L5sUnDZ96zHrszXNfxdRmAR72JLD2FtNn2HOUQombQ2nU9oZY1TvCqWvqwy+A0z6HjA
7HRe5CSlfndxeH+sOGsKBR4IVgXJWgsy0Pq7P4B4da2gJvUdrIgL6+7sSlPYglpSwBen8qsQr/i4
Kyf5daAo6SBDEyOo8HUSf638UKrpmP2j4l/6yH5+JBGlDix3DNAUMJv5DYFqExZHlGaitkj5tXV6
OW0GoNK9ZeUp/2jmtbpxKAPfPJucCu0qjZoDh6sxUfx+gpm1aMaeVtIqvkaLCHr/+f/2Cpizxye8
tjAvQUwupU1ehfk8fMa1Y+Wd4ZRe+aWG95NDUgpUtYHByvS8BhHtip/Ilacs98TWEqRzSY/v0zw2
NoWnt0ULw4elc35uvaw5DmBR1Qva5DyJN5wk+0t9/2ArJZoYyE0cbGPctjCpIx2nVl7hjtaw+Wch
qgRFZxrCKzZf04nL/8b1nV7SXJMQfoU32KmFm3JpmSs+np1bpnAEolew1piPo5yUVxRPFLxZGsfP
uTZdpZrzhnFJqU//5IAfr8aTHZQwIltyltEsKPmaLzq/dsh1kwpvOJohg59znp18FA0WLtNGQgkd
Ry7vCWkvqxufU/PKOpRbEzJD8+so4ikoYm42IOul14wl1Z3TdimAfjZ+gGAgKAl9cGFCzMkyz9hu
gs5Ib2hVGRnk5FN1OY4HhPvfRK/5Gg7lSD1jaDw0WivUso4CY60VsebDtP43jHn/vTO1pkoWVZvw
+REvghCP7v7yuWIGVCsuAnbKRGbq6WaWh3aMV0XQ1CYeDaVkE8FoRhe+Dvty9T50QV8G03+SsnaD
8OyX9IcVksHGMHtzqOmtDwuybUsXhh0rOr74Qc61M/MIh4v9GAPwTOIqbFct2WDCh2/EUQtzRELM
9NiWnS7KU8OB48w6Ow/vW/VkIo9aMF4+gl260Q9P65v67khaHEh292owyiPY/g8Rn3bWU2RMpIv0
Oc3O7g56Y4CVnUSOO/HB4pQ17xWf0xyD3Tr3ucALyD3wDCys4DN7NECHlx4pdz2bKUsUy7cRqOjx
ro5l1CdGz1RbbeNtXTrymDKWHHBhl9O3CkQQoDTDb9msH7DznSVq0mGSiHmzejaj/pevKiHpOqFa
V5FpsGDXtAWKHFnlnZuZuFJ8Cg0zT1jJrWZwp0wQReJyqTtu5DeKkWlMvORBfktE5QZ7FP/Sh8J9
d5Sw3LkvEi2Z/44+wifmfpQgmsfQq0dPoxH3LsDGQMzGhy5vDDPnizgedQPgBVuEEMzaG0GYRLIo
vgN2mgr1LpyvzE5nI0pL19ZNUchDouJloQmzYgH43SOphgmzDkkizxkBoBacASSr0MHQDcV/DLDu
N/MuYK63WG/spNyMnPs5NEi5G7sRVHZV/rQgo0pjTz4IS0KOszDHMDfIiUTcKiYfpzogHv9tDknf
kZJ6BYUaSx9V5T6WnZWCtRLU4xn6ndCn3xb1dQAlGBIZXj6FVg4diNPPXClE02DO19MyRBnGWK39
RdCQNXGAYtvYMJFQtzj12CQbe7O9eMTNaM4Cs2JZK6RTXEynFxSBJKIfbrCO7ov9NDQ+ZgoGwAAo
o03KQzXdb6/rLXOrUByspc0yRPHZLAgIzN5NZPRkNONr9rO1PuY48klTEqx2vAs9up1GSKtAqkGC
rsDHSafqduoXjoVIZ0c6u3JSJ3k7QPSIYcnOqoIAksADheXDXjmCPLCCZjoVC7XBnUuEJYiQbFOT
5cI9KOgw6OqQiF3jB5ccUkEP2YLWiWsq1UAu0midX9X7QYWNvgTcjazhAMppUy5XtewQ4Eb/htBa
cpAXtlS0FvsD+wqy53Z6HZLwsNBOdxu1PJo7Vj4Kw8RGak2XlXuKYw6CiocPDgNyWKucZs4Wr1YM
MbS2YFeSiSCR994F5TTD3JVDNgcjwze5BzXsOnaqb41h4jDlcCnAwrRxFI2WuRqgUW+Ls6xrRyT8
3aUNYw6cLRNDvra6Wj3z9XyHGTspEKM1WlTeh5i8Q7qwgwM9lz0VKJDqzS0WZH8DqQd8n6mDPxVY
oojlPxTUIOLwSekvtO2x7ye/yev8fLHbwCdvXy3WOBqs8oxXARHYFq3eyspHxA0UlOSs6wl6AwaD
gosIEqK6qf1Pg9++GM7PIQ1OyOcVN1uX4+1LQw7ErkufL37/2YzMPMzXLMVNZJPQ5Og0BTXXJyxq
2VWhuf9/osCduwQeah6g2iIM1ieaYNgsqBtRZrfACOC1EoV4BNofuWMHHPLLYkMk/M1FTtpD5R0X
Cv8VHTyxvBDLG42r95NJKrBlEt5wr3z/j3GvbUgDSk1dNpys8JFXGKFL77k1Zc58glG55SKm20pe
7hRTTN7fUFnTQl1AhIb5wKbme1+RFZ9mE5qQgAAQDvRje7FvFTK0X+SyJ7AnXy7cshe+GQt0rWSV
WbMEnCqMaWp1MA/k1Mr9Fo4kwgEq0IJuEd4VGy1YvlgAk6QSrS5KVd8Zgw9KkNaPjF23axqrLYRM
psT/6KJUl74gn0DhO2h0fuiHIVhb/2FDwX5qWuVj8waCFocFJy8ILPquGRKBR8iiQaImAcc6nZuP
01OZB1Ujo24/0wScxpvevAqJ7sEer1nrkWeSVQRsycshcM6i7tWUKmDwUs6KOLsvcntu+8tvXUSX
ctVAKDJsk+M22xL0MW3Diyguhq0u11FXOcA9LxJtoaD9vxkJAIkRpKtRMh5hwKTrbEy0lslSngtK
7oB3rgReH+sAPpnMRB0o8mI2Kb4nu3N0Y9ABjpDO+C/nFWxgCtPORGKe/Z/5tfmXggNgfrLB+Rb6
yDIOp3BUm6ajHkxUuhV0SZLyy3B19n8g2z/szi9H0zZO7liETlsn3WBQ2BaTsu4JXkzX+7yS6xZf
BodpGaHPJr7519SHlxZhG4B3eXkAVdExgr8h4z8heDCPS2nB/sjqrwayt8BbRNKAmDMbDEGSd9cr
1rLsV0IJtlnyCusArGlbBiG1vGDs/Y+JFeAbyD2FN+CM3LpvSgxrRfxVOT5cqV0DokoAj0lwsUE3
ogOo73MRf2hk2eNTpd4KdIBrQS9h/2Df9Eb2e5vZklrPXLE0mHXeGVPLRa56VdyMklOkPg1Vwt9E
XUg+U8BAw0dd2pRU2yGL6vzg3L4dE/t3zfHGkMdSgIqDpu6meOYxfdjj+ZmtIEFn3f8vwYbHRfvt
9WSj2hHMaxiQvfz9KEwAx85f5MqQc/oFoGQX2mgaPhVdYVXmGencguGy+MYPu5+zM1DGl0TIWHsj
6EaLPRx2GG+/XGmQq8IANOUZd+CjT2KK9JMAz7yB2D5lDIN7qAQ/U10Iw25FdI6BH56jznesQvnK
ak0yxgkx054f47rHt9Ye1vEQ7Y/GEf3jBzEbDDMkwDm7dlm/sJsZnGDqfwNRCVfPHXbSdhdrg8Wf
f3t5NmYf/9cwwRH/c2R5trx3n8hnnfHsrZtcrWMOWS6HJ+Arz8KAlXzE1m4wig52JDkXQYUaClE4
TS6dKz2JXbh/llYYNcH12IIXQJw3bcve9zqlZnJfVZuED6NHL2HFTgtPKmHB4rHtVv8rNUsbmqNv
WosNc7SSgDtXW0DijU2oEqn1e/6ShnRGnjbdCJVo4nb5Ue2k0I6+fNXjG/n0Rm5ulb7oKqBsynl/
sj5Nq4q8QTcsdc56HE1JhlT3X7UmeQv3DgjMok7MX7VzvsqxrsehuCKdNNijyTu/PgxN00xNtuQE
z70Zq+NdIbE1mbjTE9asLe2W5p94E6+UNtuHc90ZRIk3ruluKDeS8q0CdetASdwDxre3mVjBrGfd
O6Aq8Dbvs24aH7mCuMhIutZ//6dM/5uR7+JK/yQzjcpTydvwz5tEgc9bLPW93LLisMLwdF8LdyPt
OK6ZmnPa1hjJE3InAT7mTq2nfniVmVsE5devosEYfI5EyoSw7EuWo4C97XMhYpghV0f4OaYyF+yL
ZvnglxQwvuI1AcBML8AjmwUbZ0zvprULoD58ZSCfNKuQ4CRg1O4GNRwhLxW0G02overbGduZ762M
e9t/2USOIRAYMnBGcW7nzHprdKgWIG87nRiIt2o1kQZyisSjfyqbtdb2G9dGTqpDLR8YnKbUzo/t
q34bmqrFMmi1ZqZvA+gHLHr1yNEKQrDGu2iBdT7QGUv0i9KlqmNomPCExKhFzpUSTHXzdB5lC+ue
kWMOVrQUt9PiJejWaB3jLf8ukvWqKc04EKHYDC7krlmLmtcnMr93atvjO6p+H5Qagh39tUnpQJdQ
cyp7OpO+siVJxKDmP70zXdGRf03t1yTOlZLxbqOEPDhmbtZvfJ4xwB6uvkOssG5zo43sVh22Jn3R
nG5COpVDS3ko87CME/S7Xm/4SZu0EPMMwvdx8pgQuioM05hanOpJpYrMqi0RqVs7RkXaYpaok+jX
1+so8rH/DHEr7qoSn55Ca0aNsjdEaLROoIFXqkMryUDWOnOaka5tXVSkBiyLik7QJ4Ar2mzNCjiX
R8yTqmRuBdZ+cwqnOqfzu4LDL9PVgWDE/YRcZN5EzS8ZXqGeblRl0CIDHEEROOxLqEWGYQpOIKG1
DFfUCCMAlJKOa4BPT4jQqTvo2CkyCPo3E7O4WZArzzJx/Boig09/J2LHcGGsMW1fCAdGlyeR9kEl
4ScZf/AKUZgY883s2bAZtKVqHmneXAmNlU7t5m1O9SfWYFCFQ54HIVcLwp/1ecTmH/QZDZZtaYRh
C3U6mcSk/sF8X8ESheNduPxcaOmzMq3IL6DfrXGEcXJhOf3gKRgGEHf1wy/Bzd4CzkgcbWONTcei
/Yn7Q5FEb0Fze2vvuOhoIfpYBKte7mlvalaozMyhm+vDAPQ8rrpxWLDCNKwoMKW3gj5nURF21RN/
H/wO1H8TrnKit5WQTeyVi+Vbve1Vdm6Xn7KwE85p+JjecV1+zIrAWglClThQTG9zb7qvOLDFumS+
ZANbJKb9dKbEio5cGZOia0+ktRdKJBodVnomTnNBkmlY+uYwMi4F7JKer1TpG78W7pRtJkxqnl94
EV2Nvgh3CJpMkdi2lbEoiYW6dBPtOht0g1CHcPfiSBhfweh0LqIaSYGc3d5EJ1JD5tuIR8My+GPa
dGd4xdd2TfxdkwkoK3SQNmZKAJTQlcXV3qTydQ+ebWTM86fLdwifltXFU53zKhbjcU6guD0zJYV1
2z2qEdrSnTwY/9ciOUMpQDiiKAUaKoh/aIX46miMkSx+dTreN0pviyoLMk4Jfoa3E1E7eqT09Gyf
05egUHE7iNQ5405spt5E8HP9Icux6ow7cjQdkcIL/ASRa3laidjJG1OL8Ea0V02FslfYzGcg/Tuk
lKFuF+wgxK8GvTkk3Ux9JOW41n8pIOZr9LBfH84yW3M1Q1CcXw9FX+f7wPHjWamp5m/uUveMB5ku
Y1Q/RTtzdaoQA69O5htjfFRusVsMrsVKfgsDECSZ3FKZcurGpprWQEhUCtTd/qliwv0Mefljae+4
IdGGX/yWleXiC7FRuVpjiDynfhZ/pz+j0kuzSkdJ5P+4PxiWW8YlNMH0QusMUIaR6AQGtvbLJ2i+
shmpOxD7cUISk4JTSAMOf+/D/vtuRaNsUA6h4xmH/pIJhqLTPfWjUjC8WEHsUqynY/V0lrUJIwFF
bisyIlxz8rH/N6UEQCP1YuAsF2d2Ur8lZ159SpjCJBof6i5QbrhdZjHhlaoXbAi30nHaRGNauu2j
nAeSpnAb1PhtGs0YXUkJv0ufbhUOJ1RiWFBJ0vvSEPgV8E+YOGTxesQYZ5MsK6e0I7rGscaBfgRF
2349kZRzu5XbgQdZHuafvex0SG9EEmQzp2+zERjdRIIhPeicQqLLjqTJ3CSb44uWrHhCb0xe/Nc9
AycHdtbSMZC2mbI187aiNZx0OsfdVYwGme6g3XWNEX60DaBFTH0bFdZTqlCOOaR3qMbeo9HeNW1L
Cm+Y5POw3M8nuZFnMikp4RAnHXeln7GavsAaAYMXYIboGFj+cu4jS6G8rZdSJRciI9Mo4DYO6CqO
slowczqoYT7M5Qw5ZtFOQfduYD7Vj+GYCocr1cnonsbQoArJTUeA02oeaMYggJVbuviie64efVZI
6l6fgNgAxS8COYwSPuCdbUokhhOyo9jTnzx2H1p30GIr8HOpuZ+pUohOlqwWPDYcd4yyGqj5BY/X
OwSkoR19LK1R2z+QFc5y7oAMALVBXDYjlswd+m0dJsvl6Ow8PNhdENgO/p4ztqRevI7uYAnAvDin
BWB9myygf4/SwD1J+Owks71o39eh+aOySUU7Rzz0fHgj4LVDSem50BYxNdEZYv/49WFbtMfuqJvU
LYQRyZjEkcFEHz9WcJgp75ohZvLKR0TICW1xO9epO7W4pGaiU+G6eNgSAgN2tEIWWXo5C0wSq1S9
dHUxebclElMDGYVTTOMYBYoOVTkPtXQa6ZXgRl8QU4aGIrHIISzOPAV0eTHPSH4L4Tj5AtYGeObj
OOWjP7Kh/1Pk87MF6ZuK3U6LQev3h4xj9/ko6iHFeciWM2G6fh57naMKpQp10J5azXhIx3SM1GTl
Vko00aNCOvNnWJH4/KB/c/VhXA1hAMR4Uj7Bw5hMHi8h4qTShpZj8O/NoaV/ko6LnSQs9Wn8oPys
SXTI0/W/8FggKnn+vKY9uFrhyVrOZ44/WzDZLkK3wJGIcSwvx/7iWbGRUfl8aRSKpTkmI0b5kTrB
xCZ38YxX4hJgnTyqfKoDTfPoy/6VAA/fXsBDlw64NiAp+b53wZ64SkgckG+y+FEDiGpWK/vywJBf
JBDfKDL86Vyuhy93mM9SC1t4itAnSlZyThmOPJWb4rqZ1vOaQ/pTg1L4RYEmQpfB4chRwGUYh9Hh
+eVwT9htQ+nS8oWBNc/oBFva0CXnD6X9pB6O2JS7VBu/27WJp6jC8sPzNBZeUWmGuz5Rn808ECkD
YPIwvzjuoX++j6OPOL9qd6KokBEmSB5aUxzrvDo67zf5tBlMXDTUr/OcDCvFSHJwZ1rFNMgQbobC
PCClldzQffJrnoLdYxQ3rdY5RQAPuKtihZNTYnk1iNpoEG2/dtOtfFNlrMML9dyx4pxDonFyoddL
2X+iUL1+q6JmtzUeTjjeb7I+FlyB7tncWo7KHQchiWifenM1t98g4BUCUggGlMWHpfL2wQUAxRaZ
8MpjqwK+cuG6HcfxOsXrrhrDvrT6HZICWRoLVR9hY3CJ19OjRa5QqxNS4HUFBqSy4Cho6CNlaei5
KXZfMf1xa/YZyYrvPgxIm+uH6OLMX29E8N5tyIUoowCSrPeNno+aiNr/8Jw+giZYjNAxSEXBvFbo
vLXfXbDi4CgfX83sX1iq5Cs5jJbCQQ5StTeO2OYujZRM8vuyrmoACg0y3hOPLjake8JpSQ8R6MQZ
O022LvgJJoYbiKgvFoUQA8eHxAOMd4n++AB+qH+Oy2fVp7uQ+SHWQpqDBIdfhSioHI3xImx6M1Ef
ZzcUqFbtX+TXLHUILq72croUy1oTTDtfa1xcWNBzwydS+wrVYkJc+TGRoox1V14DuTyKQgKztjIW
6WWp2JUTtxg5JALlXcdeQ3oR0r5XXZ5Sx/LoYVayHyFpjoXVWfNB/TKmXG0zWEkTNdBmmw94HKoY
jMMOus008mH/pQUcJh5x9hM1qFWOezRGA0gvcKxL12m0Fqw47/jFfMB3CZ2LHDT6xs4AHiicuU6w
EK+5uSgLQyn01DsCeZv1hSp6ffSvUQgfRgaXJ0lBIJnr9Le9aWII/JiOKFvfSZtgzeeH493fLQuO
Cf+SMcylLcxVhlpVU5iCXbZQIpXNgaUqkfovFLSS/rQTyIAqVgxwSXdnYEwja/qWIMdToMQEW2eJ
tf5ZhdbBd2T7ntHDtp615VWwdqreVpr5nNUWv29uekM65z+1gSBvJXLpA2vLwltUUEZHD3btzRtx
kH96u5cSqRMSXA5ngqx1Tg0LCcMfuD5aR2WAYPTpNhuZLNZrHAhMZcqm6+Pyxn//yK4QtRyJTjt2
Z+MIO0ddY8d+yob0Wp9F85eaFNCbxlEVXZMc5PiOEPUgf+mX2slk2ngh8m8Ce1eR//QF7nde62r3
S5BWSGOft48XaeG2rhu+Ti6sLZKIhbqNnv/+23Kssu9hgtl1ykYs41TsHI563gv3iFSyuZTrgf5b
kjs/vJRXzIeWeQaQSeEB7o6x5LvQk/0DIM1G5bOhlGJd5QGkY/GHworWJYLRJ8XHtfwD+ldaFBBf
mEFjtsK0AzxDosPRo8hvh0xe4Q/atZOW28f/mf3ggDuMLnA/L2nP/lAVZTVHivXv6osJix1syu98
pS7wCIVrSmWo78rwIGNNgT7OODZLYKxlfSsqUcIBk/D1r44XLT82Q2KCy613KlH0SlQ3a22IvDT9
5xhs6ZII+jO5Ovvz2hLBLrsRXszWQAoZrLsx7+uxponB/83nmhsU38DSRf0QmJAyB9T5ZIO/392G
1lXJnkccUeiB49aIzl8LimV3UGuu7sj6NNp/KjaDh9XCr/5hm997q0jSn0LmfGvdhUJHwLxB3qyX
It4EdjXdK6SILH02D1WXtNTOBXHuKesUSjxEt9Y9UzXQx8Sw4C2yf6qkS9Apbn/nHnYrNHi3T+mj
vfFsF+fPEu/0LZhXqwMkPvQeFINE+ZDapykY1CmSbUI62XIhatFIgQ75mR38/jffmWyQd7tLU9A1
5eX/zXhXxRQ8S9InjGLeV2dFV1XtoMzpbkcTtCQoxCS00r77AKeKZe+yFeSt06uorwuQ8HI9pY06
BZEPdynsjjqLQqflB+avna/P1xCUWXVnolhkIP/BX/2KU95IBxQ51PypqTVh3h0nZ99di2vLdBfq
nCLKiIuwG7xc5j3OHpXTtKKWcK54ACS3yFN99FEZnlmTPBTQcMAJOdeiRFzX2MLXJKycOpfQIha7
v/gIgPznsQ3mJ/vE0SLXqqe20bLs2NZHoVvdmHrTlFIcKTco0WBcltMm0336cSsomYsSupf5WyQm
0bLgZdQh+eZ5XNm/g07TmlJnMblMhxJsusqNPYx04AAupsFSBFl10bCtiTJwkUTMuM5m2TiV7tZz
AtPeBozjijIe8IfH+o0lE6mOLG0AwG7P0txcAK+UBzn8LM0wHLLaQFOnh/2CdYQCY7xqbamdOOl0
IJ0PW7YiOQVaxen4YBGZhycP7ZssGy4qh4WRqrpU0AFZPHQ3+cxg5oOHvDsnjLJg5+/Pc+5/0Anv
I3X+hXsATCaEzmKjFRI8LorYuD7Th+dVaTAd0Nk90opdgQseBoui3zeOqlqGciM/XiCXH9pRiPnr
5X1ucjoxdpI0L/ZJokNhngkj9mZFanM+BrzbKyI4H1yhbtmlkL/uNX55m2Rbmo/eaavKRu2fR/be
MrHSPtzyQVdeqB+ZmCT5o9HZHTozTQZKaQSIUikfVAKsqousThr3s7X4MjcdgW8oDWcSfKu3wt2K
zNC1y92jixl/QO4hzYLc7drFdseZmLQXPMA7SYo8VmeHaL8XakrrWHvnP26LfqMbSG+41MxPP44l
oMobYzahwJ2OlhOL3dNPpQmlFNPtO6uJlcbeOTvIZHDR/x/fx+nT4Dju9AzzGMUICBPYZLrjmVVp
oBAw22bZdh7TH7AHp6dgjLc/Hf44Gvy3okH4ZrsRuztvvnzphkxf2c1VdxbH48rb1mL3MlQDQaXQ
mmXkSSo2xfKr0ELwt0rxUIEDdFw7KqEEZ1whqvP1fPNXO80KXYbQUSjkyj+l2LR9QsWwruO/RP3v
Ndv8ANe6r1AlvNPNFfHgH2hBf1YMyWwku5DqjVQANpwLgGd6NriuKHN732ygDstb0Op0l/QdG6/Z
AmnSPdI6hSm2TPfnQyWVTyl2yUxCLZADo3kc911cBwkHEU++Ygzusw9wPo65zgbQUm00VgbzEe6q
Fb3vl0wC4yVIrCjGKlsw4gsuH7PRslIPjTrIi+WQ9JBuJkPF5RJra/d6R+ENzs+Jx15VWFZXMLbB
R84Jzm6OiSXK8xx8jFFbu7EEp6rw/hyZGJgdgYGD4BcsXdghW3kBLIYmEvLC+z9jvY5K0Vi0Byi1
Dpdc1cnw1nfh2X3Tf1xzEhJQmheC2aH1RxA+dQXZa5o3ccV4hYeCnd4OCaq5bOmfFv9mHx2okWQU
Vg7J6N7z5jBlaRLXiBWmfjObl4VApWb0pTysCqwZkd5K6hATArzEEjXUeTpRiINmidaMtMGZmisJ
uqd0HO6/9SjPz8gwSYpcbBsFuLqoNGwUKFNiZndHT12s0MwGBVpFYimBdqFVjxPLaHJkz/om1diT
c8A5hz8LWSGDlzt0OjULgiqqLY1v8Hsh2POdxNg2MxnVT91av2UZTqskNguf32jnlNKNvF8srynr
6GR2VLHR3SdF+sskvAukfTGl0RoXgcwP+7LB1GDeOAh2T6noiAOGRfqGTVznIehC0To35YlF04Ay
tEAIIaqTLXvvdnQiBiJmWbIuYkclamBdOIry9G1Ck6Z7HxciMZ49dm62w+Klqb7dQr8fLwNh8WYL
Xwmjla505pe6gxGzdeCapu3Gz+QcFDgSgCJidBSt0ZY3kjz0ZIM5DoxQx8kzON6gn359KcK7vNXa
tcUzPz7zJavftWWEBXWJtCWPYTpwLia5JnSnL1YIf+1HI/Nl0e0SxwJEroF3VwlzW03MlDIFSNhE
EheAGyqWHIUAr7YufzyLjmxnYaFtxTfo2oNC2oy9sZIWy9PzX/M168XJ22ZzPorm5tUCkNYiwUAX
sr7skXVoQJhVEw8lGMIZj3nsqDAuuWhWMlmWH53YOtzseONyhUX9LJGHbOF97oasq/tco1HqAmoi
cFCpijHBok6cuWnmr9LSotkGfX5MftnW/+YOns/ShpolAUwLXjSv68oy+EGuJebcuSi4syJYhcbU
oUBd/IpcfK0JMvlzJRCYxHzPxDnPV8mI8Fi1eRtht2/UdjKaUbrfvWip69wGDFfCcLFUeXrDZGci
Oc4MCvEpzEeqWPKmVHV+U8yvX38yhk/n27H+NiHXZ0N7SCUFLwd6zhq9KtQQ1LtGPnjzsa4gq3co
itrZLE+gk700gNgFF1gr3yVWqtl0BHtFfNFGnimAlL6p8vFK9pBekDmOuESJ3hHHid/KctXDJllt
YGmqDVTBUTqQGo509UrtJOJsV/7NFBorZX3GXS6BTK+MB/0tCEQ9z78pBtHfsyXC0rk/oAalDv07
r8ziRB0Rdzuz4PUZIa7IzTptfdZb/foWMbQ8PTy3Jxku/7wH2Id8ojpP+kOY/sUuRRJZ6tIG1niR
hj7ucxRw1IWZ/Xd1fdjhzXNYDS9Qo7k4hszDAyOqpQUP1H+p8132l8/lrAcs1h3uKu0fobXrpqQ1
SVcQEC9Ia36/1uWkNqHrB8ift9oxTJlr3v+LdBMSGBDwBzaiGu9gDfDO/fBLL7SfsrJSbaRjJJk2
1neTRFdO4cgnB/MVkhgEylyz85fMXS6xcnoar6EORN1AZstIMDdnMEW1QxQULvLB1Od8rx/Zf/NS
EkOXTCM9aYDYmbFyVSgcwi44tgeV9SacSmDLVqlIHxgPhLznhOe4iuDDH+Hie5+A/CvUqtB9d/qz
XjilHGqKy4zlBPWnmI7pYMFrit6ec3hKIaaVFtC5NDnM21sxv9VBZxk8RyLj2w+RDSlL4kr36pp1
9MQREIsL1Z42FDnQ+Im66CSqpwIuAxBynMnurYpeFaLn5luZ869Y6MJu0SREBLWY/cdzkTOD/sr2
Arx+wtv1MGYzcI9PTQqQCyOpmUxTjavFpBw7hP2uaHZGuFsuWKHJgGhlnlwk9+/7tVone2m0z3Vc
WrfZRi+go3NtPDXW3S7u9E6tpwZIdWFZCMWoCW5p0+pjb0lx1kXctP+u+kPlvp0PDnP8oB0JIZcy
iq0enVQ/ZpD0ydSsxjVWnYZowaEJzjLnVdcTwHbisTJB4qB8qWVreh8MDpPGXAqpLi6JSzQefAdg
pPtyiukC/oJCHYEIY6QfIjsWGPUjg6K40aTLrrbCc5QYG/42FGmNfXkQx2+vmHWlYeHb1q6ec0pd
a3syJ7a8zzHPflPOEGbOiqmsxDIxMspD0Yp4y1A98PwanMx5xELDr5QJl87EeAdn1W5WX0fC9Gy1
J6R6BofGkwGG0Rijb8QRYzGgAWpq5+UOFkb0OPnKv01lRtW7eqaobvvTE/oWAjeH7nZFYKjbZaNJ
DB7414uxuKYT7087T4hrrDui1yLAyZTnmUyZvtzTO/3X05h388eTeCX16ip2Tf/DckxyKzk2B5OA
39/c61oIdiPxOr3LutB5JYD2FX8CamDh7brsnoun+tpV4ouRnPH9odftD4QGbkkwt7HiffqrbU8Z
kCBNAcq1047b3abUsVWg3+8rpr04CsID8gBZL4U13uIx3YX42L7OLhKpUU52+1OlCbK9NsNEuYH0
64wHRtqNl/xYksLY5mA9O32g0D/xOyhq7sXULHCopoP2mYcCJ/1UiX5M0/YS+bNBa0SR8VhR1ZDn
UmgDbs0Mnb6bCaCi9WK5n4xHdjLmlTiHJ2c0ic4sYfcjdhKt+7xB0R37H3lUJXZTBoHgodjngg/C
D7ZJ7JV++6UcbND1uFJjk/80bSxUZXsO294/g4DeE1Wv09fcpueMEJybncipT/jzAwqZGxkLwzu5
Uk63QKEwMIdjhdMfOQ1xeCRWEatQL9aN05G791GXwIaIxnI5KJXXzGUFF1xwJmTNIfBjSZsjTFSH
RyQ+Kh1yzmnn7HofpqeGiXSAnXly2Drt1b0HM3h+9Jzc2VE3XBHkeSPacfqMPVmHrrUE3nAsdweZ
FJ9GpW4AKakgrVXof4tWOeHEZWo9xbQ8GVuzSqD2ETiFWat+LdzH4ivMB/lTJ0Hy9zwGTODqJHfX
KHvWfYF0TrnN7HRbfOgP4xnyuewdWVoVtrkyKiu/DPqqUQf5aPIwzXLGbg6t/asp7CGxrX4v5vET
0TB9NaD73vm4PYFHmBbPnXsYwiKyRIdtdxFuYmbOIDZZhoBOeiM7oO0YmRjZ9iS1100NEAUQNqGE
iiT0ST6jwyw5Ipftr4mxHAVQtfHcQWNuIfalRjSyAl/SEwufuPD+h2qBo+buDadD8pRvGzStlKes
KtHA4P9eyylZi9C+MEx2795UuGl8Yk9kPtBVnL0KR27LwcnpkDifWCCL6XU/Jt74XncqtDaZ2+7I
IvDSmrxJqcgGPVggpG6Ww6RKqGsN527UzGT3SCmJ3Zl684zmZD7peAQ/f2lHjPeMwbq44RPZHU4y
qp0pKX4iGAVE/wbRAecUWDpXFMmU6CyIWZOghQZ1Z2HTycNGl/eN/Y8rzsLj7EY/w9QyO8yQBjSz
/gjHB8WY067tiQH1vB1fcQy4FFMVkLBHgjh3FW6AS9sYs1qIwem7nBFWw2tOCY7LeZ5cO0vTKM81
oFwBhWOqrux9KIRkvyJq9iDM3J6G3ofL65eg7XMYsGBs8g7nzKNFvO38+aOGhjFYAJ9UlGBg0XwY
naOoTuQApJI+5xKXwxAprHTa77tvzV45ED/1LjORH50vgGWuSgre6pwHNRk5LxF0kUbsKXEhPVJc
Y/ZgEeVekNAmpBooUGIktCz3WkHP7cVTQlG8UOx/mgfRDzfRpyAYW5wpej6sbJp8dZkSMsi+4Bnf
WcLXdEDO4ChVAwpvlyrIrRzQoOQLrLb3Q+3EiyJLFJXW6kIUeNMEMC9FWKu3CHWPkTCQSv/39vdQ
Ypp61CRQkLQSovekkbrTCUZfD1wSjYKI5RyS4ck5h5H/RY5rr1AvA3fT45ZDxe1i9atwrfKbsmsR
2r3oP7Kf9jot2Y+RABu5XB7Eq0AZ2hwWloa7zH2S0NxPVVSZEzUXi0EiZmN1kRwV4tF2YEXoGNEq
50USU2ALxs54zRb8UdMJPshWgmV43PvYlr/o099lBQ9waogZmoYSfxVCnnMbxIbCj5HJwM/y6eAn
on4jIvQF/13PF4KsZCFLo/tRRNK5age4Tnti6lTLFPoEMTrRn0/C2aqduZPRoiy/hxVX7eskFUUR
tHB1B3GYORi846+AW/fVJChn6M8ThLpe0VrqOpSKfOtB2LumcduANrTydc7evc6Q04+Cy8wVnW7u
q4dyroHo20bLPnLxwfgJ7eqQ5aopqhJ8mwSOycddwDPHBfqzfSF8uUySGJoJV7jTuDId/ZPfelTZ
/sEtd+wIBFiOaThWIpTVhFdYM2ISnEcxZuCouYBIr2KcCPLnunqhOsZ4ARvrj2xSG1MRMggYXkri
XO0Qe53dvwQa7TAsuZQbxaPG10gxfpFyWoqzv7aIvcUfQvtP49W7DXXbiZ/lF7u5K8q+bDkoA1Pi
WOLcI6KsvxKgqbH0yAzaPCj+hSeAh3igKZSllKV2Sof153HVGFU4MU1wiAdMpl5lKHcNyZcwIbBD
FqMTDAJx8T1hIuRB5okB5kok/NFmxWL5Pe9CDAHTMw9/XHSBEV+nhLu3/os/OVA+wdZMBIPqqMy3
Nv7wHPC3i8g5lvX1ZzRbrP5O72wDPJMxn7gfnQPUHJBT4ivpsaXgDOTU3/dUw4uec2PLUcwCiwdy
Cw5B3Zr37YogZlwC2jbZAB7D9bbb/S6F7Of2VTkIPSKFzLalMGyZdVp/6SgfysbSdD1t0E5lbh+7
deaQtn7n89Mzfa2JWdOlVQEiHZkAetn8zXGBVm5jQKvMrPUpmEIHvEYO7g+BmtvWHpe/5QZ63MWT
O8kRyMSxCG7e0m5HEt17uur4GjgNFMx48eVvhjk1N+cmIYixGrC/JFaWtWKD7rRQveyhvtNlzkmP
nb2MwzdhPg8O/yRMLobxmGCNbBhnY/B7tTbc9F5Ua2w6ur6+twSqoyyb+igNQeDmosPKzfRdpF1U
lrpD4ceflFrL9OPAJQJvg2O8JFtyWl/BRMZ9HFA/0D35mREjy6a6+c1eCi/QFNLJZq4XyrY9nz+I
cvaYoTCvP3O3T/gnGD8e2YFRhakzJ7I0VxNl7Pg9LUsCJd1nlxzudXtnktcuisK9F2pRDB61mQwD
igDJz6z6gKwoch2BNBSB4G2zShCIwYXyIq69D+eWbk/ZIA8ZwPnvPZXnkl5esWA/65Pk+UOeQQd5
48oQnBY7sR4zXkAWuOnMZxL+fCyZdKj4LIQDIqPXMskaWpI/sUykMXaN12ouPNrOsmIZVrf0c70k
jwfCHXCo4wOl4mzQCkKroLloSjUvbPtHYpKuCpbGA7g5CEBo4B5rMKcttpZBGP1E96723Do6oWdH
7VlRC+GRvInrTeD18BF9P4xw2rHguHohAkRadrPawkvXl19MCTdMrlFk21RUQ8fD/QgP+XIfXRbE
yHeH0VgVZ54W/bx/QyMJkgS7qlv9r5X7YF15t0G89diTo/W/0RaI4Jk1f8TS649+gMBmXDmpBwqk
Y7tMfpczUZJxTn1tmMgdmDB0wRHK0Q2n60pGRJM0UDPrsNlxX4hjTLDlXc2MG7HLKy/gWF0GxYEm
idFlUPWc1ER6F3z7GM5RgYaEd7DTFu8HldKHHdOtMuIynmY1QUO8YU4BpoFpuh0opuW+OAyHQAIS
nu1hhM/nOzWUZco6D9UO/aCtrzfZ12zXB1jGgj18nA1BJCWb/aqogOPAVQK1pajLrNHCWvCAPVGT
+6ldri/xm2hhin75RmIm6DqGW2Je5GOdSg1ar2qyfUTpZctb9a1v+uZYZ75MxjOMJJBv996rajcd
MXRFR9c1leWla9Y4OsuKitrNXaka2JQ3SbrSXHl15HanYGtbLizD+MVenXTEg3UPI9ytPg6BsIby
XFbBmfSNBJ4sfXHe6bIUu1nKfPuye63kaYz9GtAz2NjILY/EdyjS4ric0CkUGL2JIj5wZn/kSIeY
wUUFQGIQwfjsLGSdgPDJCCWopfrWkfNzPqarhGTIa4tPepxOsvGCkgqjnfhG21XUaoCrVwND7v8b
e6xkr8pjXXSsEOpDuTL5cHzxnbGDjsMAHmxwIynPXfm8o1czx+X+/YcO5MdRmzhWU8dDoJZL9wWL
g9GbGHAwxZpbdyi97Ty/HysfmgNnWeaJxagRt/mIuZILgktEbXvqvs93NrHwtd5k1HDH2uTQ0BYx
k5lPXyBG3R/GLSYddBUwk01sYBbr23JpWgLWuNW+XiBgUcoP04PZEt5pZ3SpqVp1I0P4d/y9BHRM
U7LmOq7/1Wx7Pg3jnaruHHJueNSsms1iy0gkFnmoMf82l8Guzfd/eK5WOQ11RpkDw2lVn4RS0F62
OojKuokUUw8v4+RnhIWFnXg5I2V7Iy/G6bPal4K1/NGOrfJGCakEsl6oPUzj0nDm2lHGhSql9J08
hkoqsguDLHBEM9XJz/6r8W4170cTPP/lXq/mpeicl0iP3buXgQQpdlI92cTJnraKQdNaaxsvpefY
DsAqjXkb7gB0h0JAoPL0E2ggXo48/dR/B1xcwXTdhMfB20tcKHPkLJzQZ7BaZUrkxwdiioeVWxhx
6Z0LEFzoOSPkUchMtAMPQ4/cyFyo7l5vOe837QBtQM0lobQEmXRUFPIOU4Zp3/djwsGAEEJhD4Cy
WLY9OdT6QM8D2BDeuVSS3MzO9+7zu+dwKYaSQo4jgSzxUTkdXUmzawkq8rlggOXswRAlzJQIuFPX
UvU3S+VTG9sXsFAIv8/hN2UUPBzUy9+lAjXON24KOIYd/2GEpQRtpBlmKFxouoK01EAGkflZ5PbB
4v4ulTvxvMVsEBsiCbSRJddWeMFc0dOHtcIdn1Zgy7i4pmPcirFyVzIPcXeR7ABJVNaCiVFfxrpk
To/tYgSG/PI4cEgkYykVJI2qFOZuL8Q2Xnr3QUxAoqJu+20RUu6VjjT3Zp2mBafOImNOcdOMca7z
18QPnrMiRk9RnWR+IYRdJ7lyubftsWhjABa67JH8/DhLoZfUHu0jawwaCpcwGUmFKmQr0St+cSb/
UfpvN/9rTDH1w26i75XYpKLOSNfQv8nOGEN+96nLpNK8Ikqm1GelFlcDdNzuDbQEPfUN00hhSiNo
S7tlWHLOcRdLAZGg+y0UGAAL96jwDAX04FPB7TvxmKleBadqXZNcXGSbbiqI5f18fQWTbuvGaHHn
PIbtauQo90Bu4++KYbe/VxeqVEs3gia+5DNWgiNfqOEh/ScOvhgXzMyUDUFOIttMasXQ9UFjydJH
3Kkj8NO2wW9AQbM1Cm6SinX2i2g+I109ofHKp10sCOgrToFhkGApPL6MGV2fIGXQ4lmYfG/V8iSE
NfvSmAgP8y8VxxiGlRP/y8K1QxQJCc7BugztSDSYfoyy2kvuVKgESS4CWrJwr6XMkTuSOSD0ZprS
6SvrcoWdGoo/vyWYFyX64hmxnICFyvM2a6x7al7abVYla9XF9ROXnihV7lTvBdwXg0T/czF65KZN
5y1PrrH5s37nwHqhSAnZxYPrYW9gKr17Vo8Ee5kwRvvguqP513V+qk3H2P19RIWK4cV0zSdm7nHi
/X7WEpn/CySDH7HB46lYiHmkUMvyw8lX5TwuOt2sEB1j1oIe0aQXCWIdPKqjsXy11naNYOJ++J8T
7sBcVFeZRiOHUjY6QNxxipgtLjIl+ssuUsT1ySQDPNrcRkbMr8eMrVNBaIMEQ34bhtCHIIGwHVK4
Dv3nXI3tcvBgHRaH2h2QYgG4sFJQ9N86xo9lZ58seMScnmqPye7AmjrJKk/EsEOkZh0dICMVsghl
uRVL/nbm8Kpk6N73MJNgPZkz13VJCaIkpt6hnWtrZrjXCGkXP27pqfmeBzEylQrOhFWKOuCiHOIl
+aR67u7vuhRbLoV9XiKehtiAb1ZGxY1id8tTEDjNT84L6nCpkyDGRFfSl05yCHHBnhLTEluLt2wp
7G2NEt8hizPmNRgEGBtOdT0dtf2EJuaZb8yAD0vNkmD3M7mZ/q717Ocx17TC3hwt0osU88CpLbC4
8lnIvEuMT4pE/cg+AacMnYRRplLsIcQKOvz91zF+Hjgm5mN2DIQphBpD1n8hj7usA3diRqsLc31z
SHIy4szMdmKhHmDQHrU8JlUu/BjUOOTKNkzwidOd+4KL/9J0taxxDPHqFm8C4mJV9CtMsnav1soO
1lg0Apk6A18ZzjAmV4RfYn+kknlXGPSIlsZ8FSPJGULwExShWQXhUsQKuqOEaBFOfEbS7wRfUtN2
+ryUDuYdbiFD9AGzL+ZqnxxLUwhp+S3+Q36ON7S7iBLCm5yX1YZqfLecCA5EtolRcOthFgLo5f62
aktUGj2hD2MqRypsAlt59dke3RDPe9dlx3sj5FkGA15TfZR6TJrmFWv64xjslDOJjDPdlGvydXcm
2Ai5yfR2ZBo8iK9ZSbjEbisgxBQGlPMIzWjZciAuROAjSmmQ2JIJqS4PHnup0EI4yt57lPTQBs6Q
bMjuy88y9kbxcYWe+ARFqi993TpoHKBDNhtqypge2SCGIq3SSwKoquG+gpU7tcRVCHnkpeXCwvOU
LvOu54/sxlZCaMLamMcpA2dd8RL8gJCE7VcIjVvP/eLOJ9Kd5yyzxo2XFde3XmKbfXIk8e4jLrx/
3Gje089DzSVBRfZ6dPjixXRbx2aoBXozy3ZrI2eqr13wQWXQnPPAkR/v+CPo/P7BZYhoNW73Mi5P
czroHBfAUtIDify6FhwuCRHhVzEFvtvaWnATEa24djKE08cgf05ml0tpazjWOtaLjv0Yp17BP4H6
SinvF+J+vtWw+R7cCrKo25ecN9s7HQO6LXlbrheIDzCqJlcVMVSwBY1KXX9IN8Vq+NYyM1sW+HFn
E68/KvVuVOgD+PVIzC8FPS1x1T4xeIeqLdA/lCUqzHPrS7sweqQpHPvK8Mc/jdQiwBeaL7vOqSFU
Kc9nyUutCBw0Vy/ddfgQ1q/H9WpZ+V8IzTKlJ1Yb712wtxK6dPRHqTqzN6JZpLRjv/rpIMZtm00Q
BMd96BgE1n2o9Q5BrmwwHZT0CcEZ8uCeFDCOWOmUfpMMsqtRQJ+KeZPYm+9dxhpD7GAJdzST94+K
Nup0ffSUgrvM4HEo92JLkhvgqOeTIIwQtPABtwyionjoRtppkRufojlmCKfBHqHoOy8H4k9eL4wS
UtxGe1DmjHOd2u4HuJgqiPOOCnhWtJd99zPYHNEREjzGvQgE2yRJ+1l+uyOObqojde/ddiWXaoJb
M80/U8ghy+w6XmMV3hbuRNFNMmlHHR9Q6YcYMN0dihSTjwNPxTzHi49q+m2xm5OQuxCiL5QzrTKC
3LF4vNguDpjA5kOQqptjMALq77OXfvuUwwUl8dkMLGHCapqkJMjBBQXgzeeDRSlvtfD/W9VtAmNA
0a1moHoVB7+MgzpLoU9X62bIvRjCyMfLSzY9vE5uv6pI7lTY2IWzO+IODeNTqXtH/blz7whLbzPV
IB+0rWm8wsRqAW07Bx5Zr2bQ8dKAChHQXh8n0/9vLMM9z35R32I/KBvDTEd24g2JDSvT4yD81MFO
TO5PO4F64GDVlJqD2yRUHtI4AYA3ANuzSNI4G4s02M1FggeASD+ToiuyM8CxB5mzAgvsbiACEoBV
HUkn9TK9NIJqHC2bvR3MvBRybc8fC2Uw4JzCFnCmZLv1FQWJn60L81LqeHKsJ1ZtyhVWt6wKbN5B
mbj8Ium37NYowOyOFX01OQvIRIYlGZhi78qXUL+erJ/x3MlhhodvlgLRFDHk1JEZZfjHIEc2ISj2
PdgVJnlsX8H+M7X7/zf3CG0266q7/m07SaOPHhVAaKcin0rvD22lfWteBVPOZbKaSzOGImSZhfbr
sxXRvQ9r4Qja/Bs3xNylinpbMxukMwaoSwz5aMxEgD8pRh5iheDFwSCzAvZwt+poU3v//mVwHutO
lSQAuZq4deCCl1aoCmMWyHAQ4i6lHGtJZ37SdBwzeTRUOtWC8KiCw5OkK47KzUyWJrmzbcl0gsnm
Z2xJEHrF5fwCxIWqX+WiO9fig8UQPhiKCgoO3jdkI/7gIsKvjFxozx9z2FK+HmEGMYP8Motbwv4E
cnNtzDxjRdfZQTUHXHkFUBEpteO8PkJ2EsySCdzZcDr9aU6UxFQdQa2qot4MgjA8mkRiLdYws5LM
RUrROd+YkgFT/1URG6BcYo6r8n8xWVk+3P2Dh2P0qpTzx+N2f5dwQqtWux9mhse4pAszouEtwRRZ
IUZ/dORBcsmV1qh8c9pXg1SO42rb2h2xtWw/oHrrjqXUxSl07vx3sR4nwcLhV4AfM2V4fy6+ZDI1
On2reCmhHz0AGdA2t6i0s1pUjAtxpGwjABslxx8MSjEN3YrwWAYpeB6MDCpyYCqVSinQy0ih8199
oLPYAPyqwA+wycVbPMbmLcSE1CsWePN5JUlYTFQtqKsc6vNJ3rgcI3rK8RovyUYgAFU2ZQeReb6R
SXnqn/z+Ie4huobtcympddpVv6vavRTmnAV8T9ngFgqAqHbF0RnqlvO6b0blfS8AB27d+nY56OEu
oL4pRjN/Nm1GGiRLStZh1k5e7gaRJ/6LJZhuXo1F8N6nEnUS84o433k5te9oGhgutSRjYiYl2QSR
gUiszD08YyO5JefSNl9VH9dqmG548PyHFrQPNhbHYxxQyYDTDIowHeEd+U8r+eqEZ8WWVnZGC9Wy
xSd7h/XVAwfdZOXu9DP93T9Rli9QKn6BYrhgQOLqHcDMTCSCC0/bdMEbDu3gJcxhHnUAop7/BGo2
LqdgPLyolap3GcG6fSRtMD2y4n6OL6osfxrB5BS0aNA5oruF5eITbmVICETvnRQMhj36JqCyuEOx
XKq5SQL4PymaEoY0hX++D+CIBdA4WJRsSdQx5317z6b18LuU6oZPCvHDWR4CJkMgql+qLbItfH5e
j3F4eDo0oRKwhJR+7AQ09BAVpyUY/0kQyvpvaAyaU2r3P40R7wYO528aiLSDTqVadbQEjV6Iwkjm
KvSKiLicrAF7/y1AO3q4R8MxM9kG+nr6RG51ptI6SYNjeeUOcZdohV9pIXg9eg7blINi3Xm/5pFG
8zSPMu+F3NPm+22aW1pfhDDWoluwOP6Co8IYBN2pIwcY/zCeGkNlYsEhfRGK+OdnhNhhS1tUUDq0
PDafhjLjuwu8YNr14+j8wrKv1JdU1PYWe8aMtYj0XM8NhjgKZUCy0tm8hypSoXK6JB2P2yngvNS4
60Zhd1jxKGvIwXI1NylLLqLwHpLTPbSRSycBcwiNGx6pXqC2cZnxwAWO+MvDeZmM2d6G1TDRdirG
eZgWbILZeIPDvlkPZqT/LXR7GeI8PuytujyBF1Xmm+mhpT+1x6OpzXVa+yZmf09npAZi9MOGO3TB
XxM6ePH7zXRpLSQSfyxJAHJnknUrQ+gNc69/3h2KQnZCaE0hSDeWVjrqZMDCQu6zCsGOOdMnFlww
b6vatokbxlXHZTPR4jliz/BtcSU+oLN6Ssw/vgiOLm7qmM1cQBTuVZDAuSCHIATFjJoPD53ZbYws
SJiVqJYz9tcKl5AKW+88hnLH/AlJpa9Qn3AbB0NT8g2piCA22aIjqMU8/qZAoV/6vKqzyJGZRviJ
jzsm0hvAUfYYDAXmU6HZSCUGDEM+WbvgN72FiYzGySCyo2WCOKZshcXS/1XaM+EpgHB1W4Jw2LT+
ctQlp0Wgl6m1il71bth6zFkfEEBJWmtMmEWID4ufqg32byZXC+szttiDSICoD/ykyreiZdegijG5
3EcAVzZ2aQ1iBYMREnwGQ2lkbQsNzBqdITw3lBriaeXHiEZHbS+gqmCzMKwn+D4VeWVpROqr0i7Z
vmOw7S7QQPhZCrGmBeS4RLz/HaIjrBabG+tjtvJ1k63L0c9zHqYZW7Zdw6ifZTmJCxYIFd+1+8q9
OBB2eezLiEjoy/Vtgs5r9iARC3IrbHUVmxyoZmNYmexvK3SOYBCEVH6got543MPtp2Zw+q59rAe3
NLs+1Dbo7Z7RuSTjOIZUc2rSdd92XKcJviKo0N2eohq/soXYBZIOC6Q+P2kJtBAFLig9K8Sw0kwN
xrBdyOVxvm9PwOgtfdnYFBsFsSld908BBXS27+ljr26B6VgoRIJndMqXK0uq0nNU9/CGx041g8rT
5ztIao1wKndMYgaf3n4sqQptNpcOj2upmht6ixXNzdZmeRCuCOf4/AecN3i9jj/kXELta6rTMaUM
GSHrOch/grVrd5t4zUlklc9n8V/Lrk71iY/oXwN/oI6S0fr5nceJYtA1ZOiykv4rHZeuQgvU6Tz1
evoybYTfBEwGoLPJHWm2hXFbfGZ/BsMoCztn7iZMDePm7WCIKqs1Qyi4lOHq/qrlwa9qsUQiDa92
hSbaTXUefXo4FIgratv7+OPc5CC2nlrbuCDz4s755WWExzQS5MLguYl92UNmJMk1j8x/nCrNl7CH
eBEisQccgvHuEEmO/F7qqIaWxINK6RGux5a3vQT9Prqtu/X6hOXwK/yjy/mCjQphqC8v864r5Pol
8S47wqsCOcWXD27KwEJqRvENpUoSisRViWP0Ff9Q8tNftoYGerivT2s8nuDfZJP7XundQECMp3Gu
eVAZlMgwB/4i29KTFbPpe+5i39xrNHUUIS4KAVdpH7nnkx3ZxruDysLQsHB0eOqHzSKUnm4/Tmri
sNmqp37Gel6ISVAG7ZR716Ftfipz4DDfBTZiaZj3/am9U3ToaCDvKCC0NuRyphFxX0BwNuuOvWXw
z1vrPlc8u+en1voLBPoti47jTTm1ltEQP/7lI6bv8m2udOz5RUlUmdAJHLkbsVtp0Mqhpau7prAU
Gc0z/0TwgfhZMKSe8JkhX5fBCnMuh8vle5SpxB6uaYrgPtXpk1L81zXRXX/78mv2Fvh5dp+7ebVQ
ljTrf+Zuz6TVMXX3+hkpjwQe59ouDQLO9HZPvWh4N7PUIMW4vasFdpKi3j6cB9+PdrQ/CuZF3SpO
c6P+5pmRrrFRc+erqzcODN+FSvznccIfhq5A/UZrH7T9edPHp/GHEgjtXs5gg2HT/wzirB7Ehn8U
E66DrVWglF1BChDuVeIREJLHCP/WqsiqZSIUHZnuqtrTrb6vLKkHs/aMRTO8t9fuo+mwXRWmeEhX
pf15NtIIX2MMxW86A+LFTlYS5gn+AoKYIOfKzSfsi4mWBBvig5NAi+uS1mUjH28yaYGs/lAG1CYs
MGgW7oEqFHUfuHhsyXAfGVKhEXmbZmMEHeHs3X33A1N5IlaPmujGJymRaZQENIwhfx5sIAaPuPOf
c8DlthLkqFnGc60Vh53IbLjJl8HE4fVJ22WJayO8GcJSMmgN4uVepNwi9dQlOXecKxotIqck+zVZ
7KtAMoxJJc2005xmj+t9JDNzamJ76SizpyMAH6spMpndn2+D9DM44vPdJ4i+sIzwDpzON/aB5Uqv
ESNEmROEwPce0kDHeaOuUQDcgNtiTVu6qZlG0onqZYb5bYoUIFPHy8S3fxFI98mwtp5YiRSnHjJl
tgemtjulqTqH6yccZReQFc99hD13FndqfVWSiEUe4M84/roogs1xZg0FsAcFlkA5Iy18FX1oFX9p
pdsnfJsS+taKfJ1cHyQTxA3+gYdVPKeat9YnFJ7X1zsoTQIedUYaz0PRtEMfWg61skTu1brpZcZs
z3FkNsHPWDN3Vn8FWWeLVsAcOfZjJ+S48Nw+nrVnEo/hROzT8BNVxHC6mY2NIVMG+PGhGCnRCKME
l7zwd7ESMJaO0Kqe7GCRY0kPA9HxVBg0CmGl0DzInjksiJEuueWMS8mQ0ycQEdRa1Y9m9atId5/s
MZjo2i0mNg4x9wXX/FvxYKy0S1F9+9EW5S9CkD8ktloc11XdSTkwEZS0QNL06Xs+1DKsIw7Q4xyd
jqIadRnDOjfrfooopZLzMLKtg0DDKxaAdwEQcayQZTa9IZZrAVH8v+7fQ3VbshN+POW+nQVakmnA
V0hVRE1oZ2oNl4L+JY27rY2vZv01m2shZXoBcHIa14X+JR9X5INzWGZcU53ff88TeL/Tjdk8Ny2U
XCl3Yg/EIWT+H1eVWQwAM9kBdqQPxH6cOPqr9u+6ww4fKnOkPe7MskR8OUPVYRKi247lUVSXP9w8
TXEWVb5JfwvO8yFCChbDU/xuug5mMhcBG8WBmf6yIXgAEbmj3soGgXWjOXRolVt5XD5iA257YXXJ
MhY0VH3b5bWxaf0Yar6lKyf4NwPFBZNYwbRhxMFSf4ycMKZrIoYHgLSVr9oFDv0QDOJ9M0ktSXJj
FJlE7xqyBj3oAhLnuErFuwmzQ7iTNmt/UThSejg1lhHUhoMsQdVwZhTJthU6DHcCCU4YUhzZkVn4
IeYZn3qTXIN6OVidjrppgQYlbd2h92/5I+vJlDJmbNiBdmcfIJgNClyt6KeHR/LZbTNTf7s+ULrA
jsr7dYWlvq1MXKElgNg3zgo4h7eLE438fiGmg6SDiR2DMqkPPxEzGOs5CuD9a3YroRD2awjY4jNL
cafieWTTDnbGdBHlIq4QpiaOepVjj94pZEJU8eGzaO8XiSVOO3pkvNO7SGH8V+DRcqbdJHk/cy/n
CmAhFHv4EWGUqH4pn2A40FoKgCxIoBqgb7NGEOD2VYaPFXYZ0cGmPwqLEDufbS+YJqgQyoofiBCE
3a13IVFAgXwL04uNHW0L0MMimUmZQ4jEdwKoXVWOgkDdVSPGFNoRjYXu3zxWltDPba3bedXc2riH
B+dOV1m9KmfzNgruC+a2ymK0cGsGpGRqu96itgqOChM6UrQqp6gR1Y4TU4oVj2w7wTDNW22r5n9R
VFuIPUHPNG8vdTICrx9CYSb/hmP5NcfUE+l34uJIB8+hf2LPX4jb+rHNoWqral0E2j2tkDRmQ9v1
Pvv/2IT2TCNOBLzeErHAflHgjtE/97MttkcTfup0udXCt4vatlqp9bgRbFtJeGVmkZnNIGno/vmx
N3QWh//iyv3JoO1HUJZ6PdTvLzoV7fLcxf0Q/xX0zkC3hyWEjVsb1m6TeJ1wkPHFAoat4Zrf7a+9
kyqKoT3UBGwHjo2EeyaR5a2L9DVEtgxNpwS1BvGzAbCADU+CJYlkWtYpewo+AVOLe74P/99OaQWK
lcamc4JeBaH1X5q7z9g87qNy3zhrMB/GF4tB4MwgIGcLw5NWaHioc3egyHGWDi1cW3nAFX3s6gqo
GkvEe2wa2eYW5zjOqthITm2CjG2fU35YaYypIU6hO1wZ4Qkm9Ml4wrtv+lL+iookufaJcUaK1SkY
6hUJEe8rw7Q6tjeeY3qJohQKOkHXrzAhH0OF5DHg8QzVvCAtYTyHFkYqP60N2R8XmN5GWTLBRWVE
HbFIdwpLV0az3pvLbxdCnNCJZrZlCF3YMhTHhT2aOzN0tH7uP5tEmmNjCnTSBEKyGnhe6pfXKrKJ
NBBjdSF3/I6oxH5B4h0MUFYwPs6tdDi6uQsgtsxZVqQibOlS80FtHi8CHBh9lEdc6NkAGorYbniw
jFgEd46r63qhs8FOm9pqJchHYNAP+qtBqA01CqnUJj23Pms5tEY0pW8xKvMPgwQMKdTgZ3NEZf4x
2GRKkHd/23GjzYgq7gOJJJnZHooan6r/Ar4Q1veByYKjAMn82rDfmzxRNUntYzyzszdWJsQXMyna
2osLVGW4RWK4grQQHv+ZiMYqhqAlkSTYK6vMtNYL1IxmeD5qOspIcqmxFD9Rmhbmkb1QYonQ+nOy
mtdVf5DpZATyS4YJr93tw5poZX7sv2fcbKo+x93O8FGwt036dB/r1yNCCdfBzlajzT3WyaMML4qg
OKoN6WTi+sxR8q0RJXEwrb8TPoIrxkHow1g/DjOEOHloUSwagh3PvmgVOzv6WMj9w+iudXbY0DRb
g1jnEOlhGhHvXZA/LzTpTJ41/8FeztdUEKk4JO6TyuymAIOHyVn28VtwllOZ7bJZixVzZpCIZMWk
6LWUI/TZUJRuc/5nd4Toxeihl7ZHpNELBAqLtOqPmeY649EzGk60f9SrUaKyOFaDf4dD6bRpReiR
8ZXEafbQt+mQxb0kVpvIuaDgPiUHLBnA/4vNlR5WJdtY9MYvRkmIEV1LChi6bi74EBPqfpiy30ry
NSBxj7BWkE5piGtNW6eWasoNAs2qLClWNTQs7KZu4wz01oneB4INhw7qqsuSmSeryxEqBtbRc8AB
t1JFvE8xcrcPSvpZob8fM55jQY9zCrpe+dPqAG8kRbMBlOvg5+sqC1PzNq5a/Wjtc710Nu0zrGH4
kxj101Fhlw8P6uX6H4xR8z8cYCDwpHSmGXNBrKn/QOwn12AXIq0+pcV5Z0RVtg0Vp8cbXlP/j//r
bRmriKAhy+8lh4ioiIIDisZmLGwishVtO1ZJxeKx8ScjaU+8NiMVii0sKe85NAgkss7Wtv8TM4tW
2hGJo5VgoRkJbN/AkDarjZrLRz0oKAH+jvtwzJaAauHnTlmz818enlCB31lVfZ2LTnAGgBouW8dq
8ybeoC/Tt/lhUpPjLOxhAlwhP5gytQheEkvNCRJkOvouWgL8uPK9hCRPh4nHn6P0ghDJ0J9d1rDf
WQ+6s1a+wV1vAIDfwihsdubspivY9TVrFO3/W4LMPcr7mHRuqb/RLUEzTlh0JASCufLB/AOVx0qk
VWrmA2ueT8w42kCKQiIOTLHmNb88dDpsp7SxhHkL0HwJciH+xhHyYsme5KSr7lnJ+TRyfOJBhNJn
9YV+1lYKlA5jAd5mkG0oSuBEzlgbD9TAWeqjw6fFNAGGjiOeK4eplVK0ToNI03SKQ0OhLWV4Kvm0
HxEr1x0Nf1voezwSdh4zBkmIBWoXbWb3+HjGQ2YC57EWBQ0HMxtpSqGFzb9UnorUBQlUbKf1csuK
wDNSYcBKU1umqtYans+qWJVI3xRa3TP1uX4A+5yCLivZRlHKKc7uKHNsGSYUblV9IKHiO+U6NN/f
vLWoKbipQOl82Y07vJizzaEsZTdrS+1PgycQBgl8JAXazGGIjvB9pcEpZWXG/CSh3vUMLttVJ+qX
4ub5WlECt5ca/YrSVtSYnPbR1AeIiodpjPCi1PqEqUbmMBiEFkMaP9QL1qpY+tJGhtgx+s/uEVyb
j4d5v0zqFXi6EwVEaIu5VZxWGKgEMyWk0HqQnd8iQox3Lf3IYHFszjiTjVonFAQsBhatD8oc+kZS
LgsVQ3pbP0VpzkOKvFZ5Bg+Df3kWSnFsGvk9PLWxlBJjQTM0Qp3X1nSPqFgCcWA2zOUaGR142psQ
yxN9Axil4eZmPA5ym2gyPv2RdGA03K+VUxcodOaxFrKt6ZprNcQpo28BRa1WR3qwQN3OtBd/esNO
hapH4psE13TpZ0o/QqNRS75ZJ5IA094HMs0G9K63vQXPicm9C+95VZGqs9hoyAqzAXYhO1E5u1yI
2vhrmSMX4k6SQR9UdUevSdF/qj/n0VHFXCKnlcPHb3ucofF7k69KufKpScRFV9ruKPVb/YxNqmkZ
j/N7igwFbSJStThwd5MCcFs4Pbl8o3/RP/fsGjd8iVAACIyz2LzIHYDCfnl/qMqhEO9iVXSg7Tg+
pZmXO6qgFQWiHu09LIjIw0LL82HxpqRJJ6g07cnI+vpMc0J9GxZowNRys+tAGyfA9uSvwaye2oKr
RCZ/6G1wb4OA2YZpT/w2zXn0FHupefIfVcW5xQI9ta5jQb+bvEmJDR7zxPs4kgp5F6Qd8CWJn9JE
GeYa087v/VN+CZ94AUz5CTgdX+afM9YSjVUB9Ms6pJQQHQm9c/h++ZxMwSTx9z9BtwBLoTYOkHCt
RN1MS10ni7JAYOWPyoSpRsmzvA/PZE0eFBxHiOY5X3UgMuCWFI8QIX42wJY1do6jbfWPUVQtUfJd
dkoxTNI9M9NydvM+PuKEya0UaheFaxt2e9nhPyiVdGNP/FMzJorr08XE78NRRRJXUj6mf1+RxQ+r
znIfUspxXOUbnQV+V92Pt3hf9aQduq2d00vi2LGI/n57fV9yN3RjtUgPZdrNZosGfhJ7eudg1Ppv
h8yd6kayioPLsfaR7Zp73ZbDAyy54xyvUG4PLlvz8WAwXv4Jxq875vnqT/TVN7M4V3lxjQZofdfu
2p7t0pSbLyXYVxDJWl91PFHWJQRbDFfXRG26GWKyx2nCG2aF3ohqQG6HwKs6wZaYgNTwX/pAoaqx
826HNSjedcmxxeN3lUiRJbC/f3TEVfDP4C9qGRDIAuxgxE9V/QAncNlZgVFd/JWFHjhyALJp8LNX
Jw2kfuFxsRF0dPt0QJMG57xDjnvgMVkQv6TIa+V5WHI81z5mlJWt3mXGyXgCZcvAKE5Jw5jeZ2fy
V/Xf+ag+FR0i7LguYny/+l67kkQrjNNONSSTIHOEzrqS23+McvDqyReh/5L7EVmPiUlVBI0ONrKz
OoWslQJtvjwrnH+4kgMbjHUG44gkSk4V7lXSpyt3pnRTHW/0Xb8gqsYVjQw2M2nqefmUY5Htnqp4
+PaQteybiD1YEB/fdXBELgqh+VOAXGOZuaWwcCHu3ybyBnIFsDCk+VOEehR9ezziGXGZgCtVdFgl
h90OkjYV3F3XanvQp0sX7pdwAKG12oxK0GoWYQx5I66GnuTYVJo34gKupYIqMllJx49dyrb1Uyen
zWdx6Tb3o4HWj2vmjklHFq8MEBmGfkAMcC1UsMUokHFM3jy7XXjsyXxxBMptn6lBzCA1ndoXXl/s
G4gkVwZ60woRsDq4lq2TW+rfM+1t8Ac3rUlIbCVwSVe0RaWJPegPDLsFvTk/JDaASX8i1a3eJw/0
1tTSofGM1ohMe/g5NC6CxVEqiIqUeNxuSK8ilrttrQ3SqY7/J9bMlb/s3zcTOmCXQjE2O4Geq8Gt
9EhFS+RzGwCHvz+yxLhMcz6WE3pZtj2MlkRK5VIxL+cqBXmXeZatstrQ0QcxYdpbwSf8gNY9/+73
wX82PHtPFvCmuEfJsOmG+JYjPN8dUg4PCxRgS7DMRVwR4CckIX7dsBXLsAqILWM8k/cB6WGTaRgv
jddnexcPG0ppsI/a0dKadPZ8a+QudSgH9vYXwfsypgRFbB1wUgmLcRLW4/pWoxAW2bobTiyaXGw7
iGCdKTW2dqlX4C/PRjgJyrGAPS7St/tS2/xm2i0euYF820wvX7RqU5vWpALF6XavZB18rcxyFfiM
DMCo+4pdXYTn9joayntSPuiQ3I9L2V6WExLQAFIFJFuP7LzOJQgtb/UOuesnrtng1wvQVs+SKQsz
skGpVE43F8y0cg793b4w4CnQD0b6r9Tdn28Hr8rwlx1Fvf68U6E3zGczaQ63eS188t7bK1Z3c5ql
M9oTWdPgVd0eiC6maon0TH6aNS0iV3CXceXl8LArDvV+WtiqahY6JhRQHYbpVQa9hxlzPFYqXj5b
jZ24IIQXWlWnVyvFPueSXamUROd7k3ZcOrMaQbSIdCpfu4fsgwZAEWCV1WV0ANb8DRsL+Vx1H3oc
mBHkz502hksIJ+s1faqxgtvLYeeKx7TQQdRV/jnKJj/3PDyemf+Cb7Gp0X71KP+IJfsZheFyFYxh
m4aUaYhGr4HTQJeelZeQv8j0+x9QWf48P7YZ56V3Z/f57lliM2sVdNNYGG6SQsnI73CXGrB7teB9
sUIXUj0aoro/NE2uxQY1QSVrG4XmmL9/fWDHp9xWJeSZ9zm+9+hmqn58qYyqDHlIzd1CqySCEvCT
7QHIz9+MIAnh7ujxVQFSMbYhMzy6ZiYkNo98pmWGzqkKaN/59WRqVZhr5LomeBPtDGR7eRZFOYG9
5c+WY97gpLxWNnFLBWlC503u1Ragf+Q2cf6poWYZiCFtUU7Jivt7H4lc9fWX5CqxO+DsqWUUEmLi
o5q3W4ZF6AchENdPYqO3ZFGwOuX7Cx8yHGzD1RiewUsD2DDKWWsMJEF2RdpHw4cB6KvnyXb2MgNv
iyX6+jdU9cjyMe4rgmh1W906gpc9BLG2DvnX64p1OykMj4J2pF2p9IRAkR4t500Fk9/yMR7ofHGz
fblUWNhEGAM0pH2HKLfODChQzQWbp83lOqXTQ2FrP45ldC4ocDvqxsDsPmFh9mEMaqVTqL/k8CEh
rUdI5mJEt3r/44MUJgdvLk9S4kD2Wx21vrL4IIQR5lk3h2AoP1F/Pz3OnW9cYp1C7XbcAo3JWPtO
yEvxxgODzrOszZnS6i6fh1hf14HUdPEhYgfN2jhxOY4Fh79ERX1pLNjKypRXIwmBwetA6fnCw5ja
xpVpqKZq4T+Q1Prxc2kg5g+5UhPcXWgUf0C27xLtpk4vTrUuoCckUHcpN7S3bgE06dRe3mBJegho
AsX3thwt7QndurU+tmHdYWfHAQYyJDnivszqKJugk7sXPVe5iPAT/TNf6dRh/da1SX+tmjb+jy7h
yJj5qsI+D69C1P6gfDOd2rp0lMrxkn4E0HHh2IwnKFJk4OlwpIPWi+VQol6e0/ctOUnXwvZA20zt
MJ7qMUXTV+jl2vZXDNocW/7fblzqkBLZy8uKLpaFxwl/OvjXOxNebQK4xinaPsT7wNz+5ep3Z1jP
qyiaMcb0YehWOLw/YBLExv2bp/IIfCpb69WS/QVNFg7D/O46bu2TgGINl9cxdKjzIaYUuyDtP4rQ
tIzniRyiYb6evfcofX0Um3G6xOJIpMlYpVc6+M2EcazVyEY7ez57mnSiaiZHCu9mWAbEnPVzJSDS
41WOvMMMZvbZt8aO1lF/j+t0aufwGzVD7p5BMh98E+6R8uW5bukbu7gSO+8/tzo6ulQ4RpaQ2S5w
6cBb79HFaxwFmRFSNvE2jq/olUYcUNU8ZbKzaYZvz63Zz4WmvcyYErDRyDFbQyxrcMCirpY+g1D7
p5Zz/g+quYWupzITZwQ+z1DQXiDtWiafRV5xtflYvlF3gp+inA5yy370DybtEVRztrk2BHXw1Izj
MZabBWVuYvz1+lmb4kkc8RywELLQ7+ZCwPfehZx/8aDF8mR8VlsiHNFiDbfI0P0izgxIlW8u9Qdq
NzOvcvFFGVznHcxgiJZZft7Ekmm5I/L/XrwJNFsmCvCzmC7phLRoIIlYOI7j1NJH1A7fQC+7wTb3
QtfcWMnCrVLKv0rZpENWtJbETczCxpLAD/FTQqATZ0GemkBVNnzjm3SC5e0i+GgZzFOc+OKgbKFR
IA5/Ssw9gzFuDBmS2O/iJBLlwWYaAPQvCxrQSKS6moN8MkKuvydZ8vIumL66N/FcX3rwloxh2yyy
zZOEzWMXRHZnflkzTMKzpq1P5q+Yx1o72nJ0/f+HWZ/T0ikwLACh22RM/DcgK5lKFI19wGhmWJ5w
cUAofCwYHz1dsKl2lW/r5PFCTUXSgYND9m/SgLFA1yEMskNJGaaTkrpMXOKvfcu4KTX+HNWZgfP9
/C5q3KV0gPpZjrOxvSfEXd+KpqCfyzpXrb187H358RiYhAJKLJNBWsHZxik/FOQQalNY0+JHHx1t
nVLnrj4J4hlh+QquyU8ayJJ2fcLCpfMpxnQ8wUIu5vMLDzWQEJl7kK41sd6m7JqJFoOVa/UrVg1V
HhQeU7rY8F8EO1HIBaq6vaKaiIiy+D1eOmrkA/T90DIUC9waQZBv10RSUArpsQd0xyVaO/XMsrbk
ERC77bvlQ6ZIJEdosZa1sz79T/9ztQICGRhd1HAxoBrVTh0eEO0+xD6A6K+ySvG/dme0AtcvPnSm
9lnZv3F4Rh7hNfij4oKe3zRLVkGiAn/jxMz8TsA9BMuJ9gGdJx1DuTH4+tb8x6S0lpbS+oOQiw/I
QSIYnZOqVCDuarolZZOsvMQXcbPR1A77d18kilpqpWQi00y4AW0pkMNe9UI6yjGVNv8jtNytJ5nn
x3IVViDGcA7kXy2xWOidrceOvs05UQ+IcDACOjOIuJJnMg7yeiZjO1A9gByKymYZWfpkJST7L9g4
sdX5nNxaCEovg5ZGfCOFK7fvVZV/1WG2kSsJWC/PBM7ixtOk7/Kx/9MkDwO05Sq6TcrilKF6nEZ+
ZsydEK8MEcbRalbfFqcrSWxyKa6QY4L7WkUwnYCDBYx+XzBpDT3PHjXuDvNB6aCuVErWFzjtHs7G
nnwWlJT+5qDARf2SHIyq+LFhAUOIxNAYtYhyB7w+gAZYwC206RUW82FI/rMZFNtRwyUzy/TT1tYZ
S5r9bfVxUd/RDMggFGDHX3Z3twq3DjGsCQ5AIbeJHbzJcwlUA/Xb1SCezhOH0d05oVRyVUBBBffF
goJWAQBI15wCmrRPcA6cnH92BPGrUC5MRgo9+KPYobfWCK3aOd2dUZNZtg4hL6P8OgRbiSKwc7mY
01qvB+203Oz/GQuK8fwzw/iJ+nWg5wYCtLkR57agppdLkMtlM3Ix9QQKapp62RRWPiKRg9mwpiKv
p3a5aax3GePmC1sp1nY29Y5T8T5Eq2tgGjHFK4A9X0KEw/GCCVJNKvnCQXvucF60581kOeZ9Gg+l
1xxBjk8bq3mTCraCsRw4X9Xyl6xtRc1e8EGscZpXTMvs6tGOW6cWVDKWN6Sg5Z9tHKTe8IJXmujB
y418tfETT9wMR4pphIPncSGHh3jj/21OCeLl958Dg5iAPJoyrdcLfHjbw3bDSqvktW8EIkZ6C8Ln
tTyRR3KV/U3Y1pB0tobG6VRLIXX7uGRusP2PsQsL5zLxPr600zz/pent4vX8zQID0Q6t+fu9Zv0q
pYQBpEGQoPQpUsKJZHE2ygtM9PrJ2bN2aPbGmWVjRJzIgpOky9EFHigyLsWa1zbsFr9ftcOiYifi
oW4RxHkjAF/76S4LPRVDHSUDr9vy3G1Nv0+J3z1P04A0EJWXvpBVP8pG3afWBhcgkfMLF74vj6Hc
+/pkrl5FemZJdWrgHYhj2Uy74yaRXYohqQ/QPdM4eru/bZb8JEiQ9Z0jpoEbDlnUOSmoU1gW9k7R
f0GlQ7WbfeopJzjXHCNeb+mdbC1FdnHH1ffdX3sV3wGscViubeZdAvO91zlKYhd3hRRHtk+DOH6O
CbBakvsoV7ZTrF9+y6KFgo4X1Urm0OYqL4hQYxC4WkFIdXNArj1uy/9XFZsrvhJLzPYHd392sg0R
RWIpNoNljwt0MksqeMgzpCn/znqxfu+JeFyeailwXjGXp2EERqNzctprBnEzx8ZSfx8+sf53HZ7v
/ah6ruZ/KMs5D6ki8nfjQTSaILEInHtrI35IPLMR+r2yp46x01KG3WVOJLyGSEb6xm+SGWTUggmA
YX4jY/vELWGhCjQzMhjA1naL0q5XSaVpCEqQtGOXFXLhx57ws/ZKg1qOAJZZDWFWIJUvtzMXBULq
hwnlVqq+cMiAlrdvtJwhPSHmWHAumV7GLpdkW2wKvB6wULIyKhxjcjyO1teOSRLSuq78bFz/QSqN
KGzTPbgNEKM4AK637ggZwNLx2z+YbS0VItJIxeRMFahoshwosVAD0zfEmd71q8Z9mww40RYwg0Sa
5N2/Dfr+5fdcLZ35y/XS+42jYqu72E8d2TWUlqQqly85KhdYEUDVNebRXz/36L7IuCXdMneD0o8t
aRwdYM4NWeAxyQVPuvV8AcBK3+NsQz+WvITkm6JBKVz7vDKsaaMNWLFucocQKNcdzR/PSpr5lqh9
Qv5nEptKuO5pPUxvJlcr1i2zTQWo7ponAPn4wj+BHQeJ0XLA/qWky/VyA0wSsi49fpZShS5mYYz4
UMU3xUkVY22Qn45lMM+2zBTJYjGdv20kPkKAwBNnT+2YN7vfVGskg0e/WxeFGCta8i4bAgnV6ksw
ZXA9PqeN+r2acMZPcYgEseya0+c9qiBwpOW2pFOG2lBWWQ3HEE0RsC3iaLq6E4K3RH+yHXPFv0wo
8M3jsvYstjlFxjEvipEF/E1d+LLLDt57B+npdnMA47D5+s71hjqUjXdPzi5fQqvHGlK6iy4bsHd6
nlghMSWaKiZ6td61R7kiuEE9MViKcPkky2zkbuX6CkJ01tGC6boz3GeNPcgeJET0xmTNd19bphxn
qpv0zy0Pf8FaYgrSV3WyhiA1jTeo3hzt3rRHTMeqk+iaah7Et42XqiwFPxv6zLrvGNcv8NiYo9N0
GXtvqCOXvQg77pewcjj6iA5X2+W3dNeFi9zIQXQHFt5bjTqqD2Pbhb0BfcMlzwRioEKHQBFyLoZs
AnXPKCafiNzLBFqVwMhj5fWxAa6n+snXq7ct7E28gkIv8NXXazuehOzWFQ3s5P9gD4Q88QFbkmKU
NSqtRN2qlAK/qopIu2kZ7uattRXjR1xYObJ3g+pA7zbJ6gjw7JJ2uV8Dhz+W20o4TZg/oMgik/s/
ta1WSC7MkElEL7tlSHH8sxndVsTNDrnlcbEzTFoEPYm0JsYWaRY3U3KyKKFsDZFCGA47+w1UH/0h
46lCJCKHQVkmPTsQRjO3NEraHXO33OWUIFq4jKAEYSTkzVDggiMJQ9GZcrjWhr4lpeLBVNO1FMjd
3k72oD9f2s7JbU4lrMsj/GCfPlX8qbu2oq5GiVbbjk5ujBmwAHYKMywCrrGO8WvXS1Jzo9VCkKFL
daTm/RaFK5cbbC5yhHXwPMGzj1dD+dBMI7Rv3CyyNHbrx334v/G91MAGMOSYb6gIK16fwenLIWFG
kiXx2LQjPYLuBMnMAsWBoFstuyWgj3AQHS0llwuBerAko8Dhaog/IUkAvaDMY+1WJnt2Bfn3aYD1
iPWQwgOKiGGo/zzQ1EE6vamzQyV5Ia7BuBzOr242moMF92Pa+6JKnzzD1wN7G7M3hcAcmtcGsYgY
Tg9YwedGXvKFygURwzpT/HyDb4d26GwSly313xuABcvBHSF9FksTWwj90mN7sWYYBy8uNg6ltTfJ
/eT6VOEJ8m8DweeZ7z5zpD2dics/1ubxYJn+LfndK4i36G/Qj2dm/RQ+kzvrwYpklyKfazKSPUPW
r0Lx21+i2PZjgaqoB2zryJi4623xHVwCOc5EiKZmmYE4OpeZoFgjhakpWrVSDOrDAN46Xb2S1fVU
eIi5r2kWq+XXX/TSl+7mc7+YVwZX0ZzUsvdFRL39AAvI3gfh+3jtrPaRgCvZ9QTVW7Tk9/NON6qU
9i32CVi71E8cgURdcw28kAza2Cnr9WHO+YZQtYxycqU4HFD1UOt51pdyWLpH2UyWFHdFrxSvJOYl
V4YTKLMgDi6LUirVBcW6JOWNaCX1uJAs5vWE3Fnz3bGhV1b9tgIHe73xFfOisz9+iWdV+TccvXdP
BOgLnWuLER5q5saZmN3FFNG+wPV+T2zS+gw5rZVWpnj6GE/BmVR4zMp3Eg0pnFwEDz6UaZNgzist
QZiZ0vTzjprqsWRFvIcEB6xPEzUb+ADvaARksOec364gV7YRMPvQfDuN5BngS3LQd0YVGwrkee8I
cb4z+VBxybWm347RVIGl7luI4ha+v5HGcqQvMRps9GKXVWPXuPYgsZ7+cGre/C2Wc9hq158UMxaO
t+JlniwdqITi4UKELdw33QRK/8DyJF955JSyOm4qGA9TRtFGbVqb5zMNm3Duh5SyWu0i98e1UIwu
Wc+wJQpfW37+Lf1Bi/3NtzSscx81nxL1/MtA7/dbXFYZWU7BnhplYpM5U1n1ueLFYtLuTLQrSNCI
CgveZITCSeL27zejyRHp8+foAhgY6K5UkYRHccnf96tDjlh7MTT5dCgk35NA5LP5F9BZ81CaAzXi
wKIzAUF+xxcYueDGtQC7g6WQgO8YU1gkAshLxfJg9NBEevsiy/XLg0OmU2Zq9xXupZaWfDwegMFo
9TCCbEwBJpU3IbIQyUKWuzNlsZ83EuVJQ4g6ctkx2PhM+KxEmK+VIZxFszV6LuVZsY0MDhi28Ndo
RuwvP9u3dSOb3mJwkotMxv1JApY84vmFj42+RLvOORXo6GFCVmSGMj1HJZoVt6+YkXFpxccOg/f0
7MHH48kdmRwsVrvIs6u7tvHeCRWoDdl6k1wNmL0Nj6bwZlQ/wET1Zm8mQejiyOfmi+5MS2ZmGXdy
RBwY1mDsYSgzfaGzdNJl8NCGM/8AALG/yhHofbW+xj+FLGwMRXLN7+ZGSRIwsyotCkcy3oAOa4BZ
dlBY+iDbaD5akwU8eYY6i1zPrcpobOMekywvW0GeqM7NzU3362C6oSrVRYVuh76agekDHA9cAUMM
T04PgE96lNN/CuGjWeQYGh3w+rgqM3rJjs/QEzghn95ybmum3lBHMqQolYcaWVlgg473gPAwIKP8
tWHcasDWhXShkaPOkZnMrl2hUelfNzU9lD5vFHSHzVpTDCyKh5cb80ppI8PuQ4K7tT8i0gR/8idc
tukBXpLP1jiaV8/HZJarwU6tAytrLCiF1mLgA49tUn2C+A7vbBIFNnPvL/9uxAXeG0j1rYJfPJq4
n3TKxScIPGoT3Ihi3avii2IJpEZ3Gtnv+RX0vw83ItpVqVXWmRyNYl/sv68GRT7BPTNzfPEtcLDK
sy0yxuszvapey8jktzL8aoDDr0ho1h8LGmaD2awupbJ1lXbU423iG2M/OBQAmB3BOD4Kt4UQjH6Z
krTjDxNqI1Ez3rBk4zeuIX0O496N6QPnpynAuz7QIyoj0QJwyfexZoSuKmE/dxWJdwn/wflFy+D/
tI/eE4qvb+VqW9qQ3iQB4jgcPHA7nEeRnYyniyiEEW9sC7cPXq6p+9Zr9lj5qfP4NPfd1pUcQE3L
vXfkPwnUWw/E9kUL16E1SMvxmr/pStWbVriSd8As3X0/x3koBwH650eTNoPMBeaKcOrD6cDatlP1
tfPu53GdP7Dvo6UuPvo6I4BW+dsz0o+HYu3K95O4tfSSLMlt4llyVjDPaO+KXBHElja/kBXF+fG+
jaVg1a8afQ9uPy6F3+nFN3VP6QpQK0k1k044G+Dt846O7ytRqFWSVfgN6JnAtW7nSfULvnIzafQH
ML4nOXqYbUVHS/IE6HWz9ePIzk5HrE3wEwYCEyKy4v9BcNPhGtR8HhMvCiG5ken+ot00c0bROIUx
pnqA3/JoTJB/05kq0diXCs+q79MUe4/FBTFtP4oSIxinQKJYwUuY30GlLxXoNnUUvP2drE60zrZs
uz6PmVy4Kaf6fz2cZfQEjFsS86azdEaJkZa+WLCyV7LXPsCqucZ7UFnl2S7fhHD1JaqiVSZkrJBD
AJil8kC2wdAFcxCdQH8z4JhLpeQJgQJv8iebHPgO2Rpcx7vUAfs4K3r4US11gTVQwyTS0IXa7tuu
FdGom9KJk7ec9lXqi4+PgG1weO+hT6nw3ct4SHdsSmL/Xs+3r6uaJj/D9aTQtkdj1I6MQXsh8NiG
NUxOeLvOoE2ORlcxSGBPYDiBX3ZHc8cPkDhMp9L6hhUOLLyc9zZPqRwrlVDOt++iD9oBCH6J7qFx
FdN0HUwF3IuKgd+/aGU7lFWfrS65r2jdJFAb3hhp95H3g6sDkayixhIgpbuBNSMKKU6Kww7HjpOt
6cpLq2rg2mc9PPCyRlT8Sb1jSVNfB0snpqSZ4umfQJ0uzwPuOgjINiCV8Ba3LemN/bYP93NPAeVt
ZYulOwHWhdv5kKczRArDAt/azeSxnHTb+xBMuhotImC0hQOSIyapzJEUV3ER5ab/7r9lYLlQXpI5
D0ULLAoem4X/Mg9z6qOCmtAv/pQxyPZ47EGk1vbA4s7gbVIjFomwRTUwonRLyYvRDkOHfUeVzZod
0j9SZY8BX4Lxk24FJ0V9mJi61UJz53O6Fpa0tuMx3nqvdYowATPFORxzZ5DRtQzofGjvv1VrVLqa
a0l4N1UpNH3c4k5n4rTA7veqty3LaohoZ75HvqssF43qPEbPI0Ud5S6k1D1B6nQer768bmtrxIXE
OyhpLdYfEb5O291p4rPaObTkcECHQAeNh6FGOCHHOmZoaIu/VmkcJtbvKMlofGzf+F2AH9avghSw
xHGdlYwdgOMHyo5cgwLbctn4+OAtN6VS47Zi4XJwNNMJWCwSwTH80rY8LFYoMCMVY173RxBUcJjJ
yYA7rHel+Yi6p8yQPd/aLTfwyjfSRFER9UwSS/Klq4IjOTzqNjFRp0s4AnB1hPhxgJnIc491oyp8
NVKWBa4zylzd3H1mSKR/vjEDrihLsh4osOEHBsy6A7Q/6pkcMONpA7Xftwg6axPpcT9vGFYaBBHH
kjY7OjymsRTZ7w0a9nVxeBfpTJDqT29r8i7pqjQEx5cPIw8hDJnBYSHzu0u7OUmS3quIQYieT46K
x/uRG40WTWESTYFkTJGiZkJmcXkprV9MbJoPCg9feC1aEK4gTq/3xDrBa2U2rGkiGr9utkTOr66d
jtFVlxfVOlstV5Majd7tolGTWhHYbds2rWdBonLzKkrxZnCunW9WFGvhRCpiZysvsqq6jwgCNvj+
fx/Egx0vb/LdVoRIGw5IFLucb/3gL2PPxcyJt9O5IIbegkvXE9lM8qysfXVQHc/ioGlZmuhQbG/z
83vDuT55KNXzEN2IuVtTHeuh3/rVDlg0OHDONN1lUa4I6r4JugAM7u3uiRa9kPcODrmbcbnLGGB3
D8ZPIUlb3Rb01T+qPkjTcOBzb8V9czqdro9AhALpO3nAHdnfwqCAkQ3eeBNdx/Rk/GNZKLM2xALF
zRyB+N1OxRTd6dknqEeTFG3pV9hWL67/qi7fTyaXpJa0m/OdBr9jaPS+Q7tuIQ6RPAP9tA4thJv5
GTkQsHLb5s8R/birg1I7K4uVU2DkGZWuh2Vcim++IlV3ieRBBBJnqQV1xm011gHHZfbf0vax3pBf
6b6cFhe371uVI24yxMAk5ppDUe46xwstnBBG/a8Z7aRxipdqCGAtjUdJoqZGwNzDMZdsYiF3uGG0
Evs/vjc15D1fQe5/CfOlvS2jl0RWDV2lQqYKd6HI4RPdGzTxRHV8ORmVp0iide8skkFRsJ5w5cNs
6zWsJ2CK7yOoIAP8S63fChxHfv4m/YfjI2YqhGogkm/R3WSq7bHD1Z0xgFu4vm74qg2S2FBgC8Me
JYSvr08BBSOCEQHuOTEPwvePmF0ExlNhtJsghytnd+Zkh0Uu/jvlH0zpD/38vEFEGPX6ISHBDC/C
2tyFZPjrE+I126ZCFFLK3wBTmNW7gvDISkKuLaAUEABX+Jq5J6L+sFaZY42aDNGR/hSMRw5pMW/l
XMg0wB1wP+ry84MvN07IPRFnkzz7W1+9g/guF3HYc6O2EURmux5niRqAIhCO5dbNY/cqUDxGGBqz
9+2Egbda0b3eZxq31skUKG/pnP/LCBkbyGxlvyI8bh/5D6tEf4HBFQ4VNAhZNLJjb5ezXPX4eDzo
O+kXobY/9ET+Rg7W4FI4FxiNy7aHUz0F8/qtWnsXlphUo9NgOoLgMKMZkQaq+bz6vvIcBhk8pjj/
WJlcAWTsj4d6+oaHtRQ2O1e4aeXSgvVAkEk9jEZh7/FHtW8pPJcE7DZmbZn0DtULtpz6P4M/GO23
+31Uj9gNsQ/bW0IRRJ9jiSYBYGOz1jN0bOVF13HXkQS6o8LAyzShd2tPitigsftrkZBOOEMkai/p
8E6vP1JKxBRo8eW7JlgZdv93Q1SlRLZufFi0GY7kI8sHsycnQHlsnA5rNsqCaIb0UKCDrOvagAr1
/6OU23JnWpFzQR7T7J02qATSNVQr0jBrzqEItx2ZCuuP/0FTl5U6FCgqqs2Bkzx2tPc7cddhcjM+
SNUoSKnaWwu/Dv7WkJbz0DqQ5ZrPjtdo0VC8Gf3FaesM5yXHixsfpA3XL3ogCqy3eK+RiUa2qdhL
TgzvhIIovbdkfnDa//gbDoUsy7ZKULaSzQfx4z+aTbVecj48YdFLGv2v/tq32CAlvdCynamRB/w9
V27DuLN7z6g5KlHsg1e5DRhz2YpHb1Vk30elK/5fx+CPc1DI+p9uZT12TpjGBESDqokc+IbgS1nb
tnO+QV7lDFpa2+WTvj68Ix2omN8WNKxwBtV3CaM1WSbUJ+9WM/n7cUfu8ANevGPyW9EqwD1+LcFt
nZFxmxw1E4sh7zpD0O4O9LVJUDYhIDNu/cH/GgWgRh/lXCB1EZrzoWwty62a6WLn5VY0JjG3xagO
EHrJruCBoTiLefy+hU7pANyPVtZNabSdVyzRfUe47J1tiAgBJWNRGYQwVp+IuSUCvaEYJvREnn5i
ScxkQlowxU4zmZlt1aEtDhEcRwbI3nx4QAgrjOJns+KnyEWYYoqi2PW7OQ2hjZG1rWUqqShFeW7H
ApFCzEE30yal1OyPOMPIPwCp9vyojUFOj75ubD3nvzt+dEJ1yc/5kciDsUr/FZZonTVE0HeRgWPL
/jSw4F+0tO3MqTgI3CLr5YNNkmA77fH26m5pRHLePklN7PtjjEJVA1tIWLziQBEHxXWYNK1Ym5pB
PKHY2JzIbn/OypVP2EbkGuMG2gk0p2AMpxwL/llQ6GhiscDK0pflC9VkZ1WEnn7dnPNHAGsYstqx
eUAyMLEPHRgrstBFOOX1b5gA8GA+X8lDjs1zd0uMMOH8NTIuFD/rw4R50K0/HxA7L06IuceSA8qz
J0bRoDkfyG3J37c3w1n1uRmevAmx3B1LNVkfOq4U6XhucaG12lPmPkwKAIc7imrphME5ZlYYej6A
Hx9Tqt4zfx6ZeXZWTrbCBBTXNgQ6u7T7AHaPOgIQvLOQbViO2L+Qmt5RmKobYLi5mnoakqqWRZpX
9GaS41rOhs5dwVj+fk+So9Ls9S5XQbPt03j7z/LMpkz4fsfav8/NDnwLU/a0o/3uUtj1uNs+e68D
3XYE0bDF7PtFYIcolUxs5cH8mc3ixvxUx5/5jUCn8dA40NaeUjLUay1Nu50AbTfT38hQB8rkGdmc
ecHMnaNmkfKkguTRCFCdmj5zAGDtwcso09rfbP2c8lojfOMQSP9gogKLWYEeHbqdiwAytwpHmW45
yxD2vzSmLxfblOvhzWtBXNPSSWQNocHnb8YvOjSaErHK85PD2zi9TZsagMosKXyL3NSSpsDHZRWM
JvJEUbDyffIq33xlgsk2I0psIaJJ4U8vszTS16i03loeTVGti59Qnf2bxsn/q+JUrEFEtA7Iw8zw
e7BDbruzWg7utM6gHSqjz4qv2O3EWMYtMBK1aoX+Ub0sUYk7wGVVy6WgbxXE8RnlOLG8q4tvcdvu
yjgZEOGCgvPMSt9FajwQ/h6BZ1zdVlCEsw7RNS4UT5VKueJU11Udt2FTuJsLAG1eu57Jur21B/gd
FZpc8ZZPFNt+yEXHow83KDe02a0JHCYz949m4YmbtR4AimjAie122QucbcUHtGMzzw2wh2d5asNk
/+YyGaA/kt1Tk97X0ldPjeOEkrrcT1rFTme/N0aFGs/uomxkKQqiZke2VqCZQepkxoYhlq9JcdLg
VHvGz5KEWFM3cuJKT7cqUT2r+wD3kR1j5Ep8CAKKCZUVA+1+m77orI4uBy+Yyzf40TaHI4+TgFDi
mFAosxvUlAJ4KW9bn0Pgo8g0nYU+CGza+jerUtWjL9N+i6OquRpEMFBuz25kS9Rg5rJYiSnaN2zG
u2XhD5Lm5Kftwc9FrdpO7cdbcGp1iT+4uxKjjI/IrZba6FKgEDImd+mCcRl3Jw2wwQHiVueAqmGD
y0n8pI9vkLdKwamx6PyE+CNEHN+f/BL1T6lLPGNeS743QpqZAp5VMhhXAye5r9gjAaS3oXKxbogH
f4cpsmAOvcHc3C9Gj4Z587sF25b2uGRd0hnNeI8XgUdaMAvXxuk/XEARkyVf9c5Jkn/YakG5j+f8
nAPSYsjY0kyrJgpabwcpnbUJD7cN8v8jaODLnbtUd+7A6uqqd1+tte8Af26S2CM7zYd3Ax7OGoa9
0G0GrAcxOfRuqKRg4r9pN4vY3hxuFGKxX8T+/n9ppUxZ6sNDdNi459e0WZu0y4pArg+pRzXvhW0O
Av+9OPx2Zfl0YzxBu5/uLtj4WNB3GviqPmRotF5aK6B/qJRTcHlgcuvOLDD/0dVGUr7JWrjOjZgG
lxYfNV6UR5sgCBdigtXfkKp5IwReLuYqxiItbOSeKP9AFgSmSuy7OAQe7ckSmIxSO8+oF4QLUwZn
XUjSsDkr8+fL5fDtoq8XscRzORofOr7WRJ18xZZXLL6YlsxFjQqhScASMPj+jrq3fncSDRsgvUfQ
/ih9ofC13xPIQ2F9q5Qe/TI/rRsFgZLsZJ2e4aewz5js1Sty+O/SQsRG3oThvKLMDvkWB3RPf4Im
GhcGo7OYjihjPlJvcfaL4Hq7IJRmfO9GsDJqaUxOXmu9LAio/4aApVAUuC1i6IbOlLKHXx8eWFXI
snB4W9pdHpINShqj7UnDCKivlLU3d0k0uFGas8AqcawxrjFmH/Do+p+zBLyBGestCGreyClJBfVg
aWfT0XrLvqMJbiSBdy84xZzLmH2jl9e/V33qIZ2RNb7dlfWBrXkoIIK8AkkcMEKIT8mxMkIOoEfF
YNrsC7HllXFp+FxcgjPCQmv+driQbVRPpSznTG8mFDiAm/C5o7nE/DxhPxYqmeBmHmfNgc1SBzAQ
JcsxktpUtmdn8yg8AF103fq3Hy9vaNCBIq68sZYgwyavW+H7O++S9tAMWjR4JmNUneP6HtsWvWfp
i4EAW0iBZYSS63RsQhYFiCsYMuDRH5IEt31sB3bynP9JAL9m0Tiy1lt8nBIc5cllwr0EW+PoEa4U
XZv4UQRovq6IuqBtrTGjXrW6n+LsxXds8mi2MVcS/nqFFQDoVWyStXewOv0B/MweszHTjUIZYtp/
9vzdOkm8IsoQr1t/jUjt9l9zGWKERRpSom+UjEX2wwsMLlMXhWfdOmBHYWYX+/CNeKEF9CLR3O+q
ol9TRkf6hG8NU0FqlxiA1Raxk8XEN4iohW1i/OSmLm16gaHeoMpwgX/dCJMA3lZZBJVh31DrojiN
graoOfiJOi6CbI9/o59KZ5DOcwrzhQOtkypLN0YAgG7c4kRAh6bUatAO81sCO19KGF41FhkFYeCV
tJzY4LL2tB7pA48251ag0my/pyqnUj+yP6qpSuRvjmyFh/+qFEPHQrPPwh5gze3Ymf/Dvtfohz6P
FjAFrROdPZHLdzLAz4eDVCwK98swjnZ2R769gAqQhmDeunznC17Hh4JdMdS7/6kSa5tKw1PXtSZI
8RFQo4CsESmCSW4RYFhxyrr4UdLHPUNt4+e3M6dxziYYtFu0Nwr0fbZxCbnRmQTazB50qtBaocur
YacyihZxIp9GHm+PXeKV3/STcXTgnkDVV2MOPo9e+RsTVQubNJCo2Wg1i/0IDTvt7Tn3c8xbIkR3
wqMJ3suwpEgS351/OqIQ6geguSx4QgcF1C15+UdjJRENUAEQGhsI5vRMj6AaP0wPI5VWFJhnoEym
50vYzT99bolTUO8Hol8Zky8v8xJgWmfX3eIUaA4sklb8k4bnfk1DCPX2qRcNslx2O7HQxk7c50fQ
3EB7R85eCTxuHZSUhgziy8FbQD/0ozVdTOKGBfQTijOCCpKGelm5SGJFuva87FL7Ywwwx8MzeI+2
VRE7a9T2YuB6cUzeqN3lCy8Cw5cHClXXbLgDBCGN9oNqImUbtrdc9h6Q2PfTHeqV76Vcj+sKsEqB
vrorB0GVDa8iC0AbVozraefAdgJCv7uGRcdvB8/OFEIqT177mnt0q7VmnWzftYdZiDl+XY7uSywq
uw0uwrJvjfY6zm8Izg/EI9N3l4u9Oyp+8Q79uxLEm22QexiijNIIQR3PqijZCqLpGbU+S2GkqIWX
tqB99l8N92oSYt78Jf0Kyg0YuqvqbRed/alMmbD5XxN/U1cXzUIcnNsySqMNdyZkGRJLEnw91PeF
6mKtjj7CuM2O7815NSuVDYZYmzw8A0M8CjJwTN+ORTZS4N3Qg0Z/+Df7mhWjQRworF4Uv9YtLatW
U25NFYAjIKdw2Oe78wDO2upivF72n0Y690s/cstZah53pPVhrpBKDMw8kIduNLbLwuh8WgGMVn4Y
1KLxe997lDX3jq7DVMn4R2ySepXEhSXYa3zA7x0c1NydQTk2eq6dP0x6Hu3kgcYZncDJ+aRNBDaK
OFicArl5io6pTAu+t5wa4jp3EjfBKdM6NsqUqNrQuMH74WyUmU/d+8fbZyl0j8Vb2pzv8vdouxfb
Fkbnj5Tave4hQYLipbTHitBOXJiVvHh8IaQ47u0JbCfc57WLmcJzbuSdJRaeP1MEvqecCpDp+zMt
6Zhvm4Jki4bbHS7/p0tsjEsI93Pb179aINZ7bLcevPN2uVRm9oBkhw7T7/FUxgAs/62DKMiuDD7O
5GcNbmxGmtaSrOkcs1MWHYsISd6IpiaqC4xXMFoOnc8TuhLPnSRoVxMHbqtEYb4E9nGLDK9UxcTq
ESHZiEQIBveaIFvY0fgZByEKjg07DXQGNSrzkjuer8rpA62pOiOVwDPViTexPehDAuQgtQoucLK9
5Z/e+FRVlloWFkcx58DiNlCyM8iy4MFvE2LhzAQ2UdA4tk8mHLKX5mvwayjttAU7/oZG1EUlp4ec
rN4kRRM/j22RFdAbOZuKArCrsyHqRvmHinAPtS8LPkVBf1vtn8uXl5FbGOV9Vq1B9DCdRUDAJ3j5
pjATu0HG1N5SO+OMqka5if6/d54/xJ7bXM2sJkt+U/rnLZJPJ7cdUfR88UMzh1jSB0ICtb/Hw148
IAgP/wbR5sqTeoNjUs/tOcETDX8SRnm56xPTsiG+C3yTgNF5timjr1hDy4Rhri6Oj3ce/iAEtssS
+ipsjqmtX7RE+mYcAt0UBQu4moUeiDMV5nS0AuqENYg34qZ72dthmCXBHkYZS8Sbu7+KMJHBfpBU
+4t4FbxbFwuAPQGzNblJDdk0EFv/BDtDzByc6N2HDpIUBcTeHqQ6eYuKHOMTWPJa5Iqdl2GksN9Z
QSYpozF9cr5ZOW56mZol8FNLs4S6Zqyj0zAznUPB9je0lgB1d+yFBs3dZOA+BhaVnWIBLoFmA9MT
4qfuggY2F21Ufjx53cQ+enAYKi32BTfloZy7KODod3ovfDpp8BhwLxW7v/lWD1bIjNlf587ZeSfS
hD6I9zSpmMywLIlMSyvCPCotuyghynGXUP/V+9SxoXbCOQzYADvYA3GmZTRNNMLvPKxldaV8GRBe
gvm9mMKonfxJfOE1HNEkPzjApQpztT/prY5AAeCLU1vY0tLaqWvxyoKGOVmpc0n2vSTcQUIlMUgP
Xa2PuU5uEMLY5xIAGWYkgdl5cuXZvorgOrk5lVhbsSV229t1m4dRZJrTgU8tzXdfgxHEgU7aOmSd
1U4NuKHuluXeilJ/qQd5IxN5fhOQvSYWSLhudoD0GNOVme1vQhd32ALcxWYwxxRj/wxmwmXC4qGq
pU6VTsizIzRtY9OJtPKJYkRa3zZR7P6U9iG8jeqZmlPoR7UVRfLIs8C+kw6UgomW2TBK6Dp0b/+e
7Teb2gYLZeu4ESKwQkcSbJgia0zk+K1x+SrR5yTBDxVEHvMJRgW40P0SbwvSE7RtuxkV8tJRnBpC
T9ej8+2Nq0abvNqgx80TQWN6s5LHAWYmO6epOxhRfTlxb+m0imCyd9K41ng71jQd7k9pYtcIDXFw
qdyGr2Pj0PYbBK1V6ITxMG/es67ITZbtIWRu9Ly0PTZ9q7MGJNYudYWHMn7wVqWlrOqVpP1PFlir
Hzly/0E0JoDBL3g4wZIBiGQE17PXXMX8i//5nsbQOAf5BD0fVnyr6CYuL09As87m9BjWZPvrZBUC
wovrhmLWTooL0SyfhMQNkwdgcQDeI2g2UFVNtaqLHDiwy76pqq8wJe0Cqa48XMCd8xJ9gB21AMkA
NlV2gDtX6slPSSlzUugNMBeVoLVoZr2sXvLROPoox09NPTXVBqcPiHLPWWsaRik7cJEx6m9JvCBD
20ofGEDJwzRpq19PBvZKIXJsgA6QruchYaxoPsMs8BrzmFK/6vXEI8oCEIUz1hy1PGQnwixyTAlK
r90W92DOrqSVSZApfF/n1ovTiGnDZRZR7MIFO1okeNGnRaX88jly6rv1vRNNGp6wFXNpHYG8SQkz
kXD1jRD0dwrl536jVnowxE25WAL9+bkQ+aKADWePeX02xQOCWs8WTwQ7iRyIb5he6kyOIgJIn221
NKEsZAi87D6oy/zxQmRgDGhi+69jP2LG/m4BEM3LNkDSvRpAWl+5Pew2bR/yLfGgp9zhl0j94Xo6
rMjOL0xxnRBft8JMcx1mmEnxzOjz6YUbru3619ct0O4tUo95J9HI7Z1HPlhXA81gtnsQvAxTx/o+
Nix9DQyq+VSHpLpN5i3Qs1aQX6ulx+lGwPkT9E7D0VO1Wufn2m9+2Nuut6Uw4BJ4WPSlOkmvAD+i
ur9cDjRMoFbMKdKEfrN/Ivkzj7H3LcXReYaAfq13j6K7J+8L+JThCRWHWb0Lu9Tl5wO+AWypKzxh
+WLYLo94/JrS2URtPA5FHPHfrNYPWQQug/ZgVdwjZ/CzkUMhJlB8VpY5wzgZW4MWQDsHH5bGrk7e
/LK6KotluFBd9+dOZehp+0otRx+QNF0l4LjElnCxTDaeUoVadg+zH6KzdQ2e1FEa9uOFC+fkk7cE
Zv2tdRrhSl7OWGcahl4dEXCpgkCqEdq7iUL2oCSV5M5X6Nu+oz9uh0MWdqUXw/T885wdarnwRpc4
VDYQFd2yW4jbpsSCWVhJBO+6++KsHEBiqiFifWyznSvPa1fMLYKJ8VjDkh8EAFwOhCYk+k5PetKv
lGFY7RO6CshSSkcWqPZ3Wg9xZ6s4S4kOtCtI74TafrbqFe0vwNKLzt9+7szmnaTepVJNMS8SVUyc
R7UhoY1Jel0adFtihP7+xyZU/PiqCk58+W+FRqFvr6GDascr/0BX/yOkUC0Y6twANPYLcCKtFOaS
HDJBbNNJuWx3YXdhUr+O8f28K4Tn6+7zQTKsuryU/O9vHeSxArKu+Jur16j3KFCRjjhZTXUbZUpL
Apa/WCVU4i35hIhG1v0pCEIU09oSWv8sBdzSaXEo28//Up8FOiv6lwnNkp65ERJcc9US8GnLgbsC
f4K5j8lCx2SpoZlp0PGtE/Z+THuLavM8mVTy9oJGOoLNXpSespzC0PNiFHPW3qqV4+fNUDuGqljO
6KApDvk8WFkhBxNe4Ho+U99vqksphThoco948++O8VxqMm1i+A6wDRd1/H7ravGEYizancI/kqFa
gAPOHvStn/uUPJMtsSDZzdT0cr4SJN1BBD5cRg4f4PLwBX2pzkmKy8/67jcOLJSv6vYxYVvvPGS3
aF3m1LeUFItj4I6kPOjP/+PsNBwo9tS+kIJcohpfemN7RaNPVFoZHwvuZKoWPPU8jmAtp/OJX2VT
caqO/yaPjJHpEsE7kpIMUf9agDu+QGWnX2OzYygKB7OMz37NOlQczh+1fWVmsMhKDdoEgvkZc5Jq
Bs47Lu9I53IoNfnVTMnMOpgb/cXrAjAuRUcxzmo0jhqCfHVVChzFLDmPILkadAKEkPSnmAVae8Dr
Y09tyoHdXon7vwoNrROPwg/+IbqRhUvIqAARRguzhU84t+KEhbvFhzK1Mc+7GBJBlbvjD+dxX24/
WyEiA2awqJiMJ3waIRKYKkT2zJEiFUsgYBQY3S8Ky8kjH23ZnWWVB5B9mbcyHV7tv9W4Ntv0WeeJ
lfzQ6RiJc0pWXTx+siXFmC6NgPoSkdHpNx3PDcXvw8IpVLZOJyMc0baGzoAs2y6FodF1eGzhHRt3
+HTonwfgHp3uImWmpmeBEyi73/31UtHbrrlhyNrD7GqJXs0smH/bLrjsUQKdeFF/UqZ+gt2tKXl3
OSw/GfTAqSiyInEAvsjK7D0qXw3B4rkVRfKiviYCzF8sI+U/Km6HogOMYFuBY8Vvu5F2PTKxHWYS
5WjQ8OmgylQ/T88GwRCzbfhOKtozH0807a7kCIoD1M1WINHoXBuovTQgFAc7Or/IWCk5PEJJFW+I
08q5HzY7UZ0uNVaoK5CQqfN58d4o1RdQbtXWSsBUhUr6Wf5N6xzVzTD3yoejvIuamwQfu58P0nSV
XVEJT3pIXFUBghgEZt8zRgNFaCVTBRYy6mGmM14/3UdF4vOXiYpAxQV0L9+CQD0hNAFhbLHkd79j
ye/QqSHZNrcqHSohE7xa4ekJ+tf4EpN+Hb5v0RgG451AiHpAlwaa7UOE971ZOxVDzvj+JhR47rke
0MYVCdPuyK7aWs3aolc3OjLbHkxqhOKweIWvdxhu0++KCR5qDlp6tVyZ8LMTW9qaMENTTgw5xF7p
XadDYa1jBxAGLyv7euQWECQqd2NmnD/+0wmqud92QSA16Nt/FSoVIelSAETilQgmPHPY3I0+Q6VU
SdKnwR1WFcQe6LHFDwTUdRjRjxjMSTKUt9IEnt2rIgc1eJ2ibSCAyVaW8/f6m8sYYY1YSd3iClI0
PJcs6lhB0WvVqKTmKhEELZTXTqnzWwCOq3uIPDT6MMcDMstJqS+fYVSGIiVTlHCSvHdz5nzTfnjD
mxLB+s4yzccm7I02CbYMvlA0jn9GofGFJR+u66uuTKUs7jD2ohApfIXJ0ugcKVc5TEgYR6QlrNm/
NlbltpuqgvKiPT8bkvAoAuy8O3dpgPrs+ZZhdqzNzEP4NFS+aGRZhiLue0IKqLqbT7ocG7WQ/ECz
/bhRhTQSrtcPvdM657v0jHtolbKsCPbXc/hGFCROjMqZHWXWjhQ7pqPOCo6SjNQ2Ocz8vIRoVNys
6VTfA/GorAINfdoTia5XFTxKHx4yP5VN4LsbLOEzieoCXo7XKO94AcRa5EJ2avrtoQUaLxnaT4d7
7C5bkA8AExGLrR64turp3YMwlJzg/oinl32BBgoTrN+yc02kHXYChki9bl6QijVhDATd2os3f9y5
q9LhX2Fw8y7xYpDaH/yr+BpbvY3X06ukzXUR9GmsmC3qlCCJg0dEkTFgMHSMGeMm3/z9+czwDjIL
BF248BAbJEYk7xldHAc+GFNQNNVJyLHewxESZx1r9JXyEIdP+A4n1kFy+acYpuimPDcp8tnEXbhj
N3xlTvDW5848iFqyemkknBe10zihCDeOYjMknbhFx3leF1s1cUszs/hI2JeDOoftXaNaOKlwqk7X
PaByMJY1iLggglvjc6Pim4i+zL/e1I8Ttw0ekcdycrkJuwCNTIVgV5M+z3qdq41I7ZAPGnLlLK5h
42/478UxbE2QTPkdXPAkdNtt2TD4PnvfW9IbTO/pv0yJbPNRJulfpxR8oojLoV8R/URglh+yunK6
Y0r3+gAUsJcBJ+hGUuCGVBzN58wg3wFsiIYr8Sbvs2PoWeSMCR3bLSjlioEnhqQEQ67972HjLMK4
Nd5T8oTCNtO2kJYVSg0uQfmZEQLm+MnraiyTBrgTEDYVYdIafBT4HPSXZwBZt/cxuSY/3AZjJnl9
GsiYg24NL0GB5HsC34GAj5ZhYJsYMrPeIUF04ZKFQFWeKL8XoOnF5muRkxcfafR0SNwz1PFitqYS
MczcBYUyQonI9HEoajNgp5EU47FmcYtSRSiewHeN8e5qWGP6SQTrjb89kGc4xOhL0nlaWflNAoDm
qEgA6ramVw7GMGgXpPeJRfBcYr1VcPN/iBObmQCkJwXRv7mtIhzN1TqWpd4LatmcWmimTdFc+NL3
PymIbmnlLSCaeaOG8mrRV0npejSZdA9cou2iTp8D3sb+sTXNknzMf/Crhi9AKvfOcmiZWf0Dru7m
3b2/yZW0s5ekFvavhUMnyQs/NsnJMIoDx1l0AR27XlsU1avFAj9BfyGjuDNCK83MgOGspoth0aKK
QkD9iImBbvZF6Qm1uJPvi9MCmcpr2CJOkwJe4BI4Soffk52+Rgq+OnzPpsfUTBId0ggOr+XlQvtF
kzwnr2IDWDg650KTFBRQdXvka3SAbbkFN30C3t7JU9tADp0WTYOWJpC6w4NvNdT4nZjiOolle13/
tNQgZr7s/qi+bcaLIS76ujfF+xEs7EmYBpuyr/ONMSrokSR0IL3oHch0MiYMTGUaQeACTyHe5VWj
vxZgkTUzKb773mOM47dzzIpanoEkS3/eWG3kg52V0qq9nyHcIsHLBU9bIjZPu0W2Ld3zS+AOTD4W
zMCkhgNpMAOzDPhUBwBQBVrULKddgaqCxLOkKA0Q+eot3H3vB7Ib2T3wKjnyMyRa0bvRZnZWwuZS
S0mkHQS99xuryoaha4rfhTPlr/NwonstFy0VogOvhbgCUizXBzJ4WdEFnefrWIPjHPrqEjWYby1F
G5dz8SmOeHXvUu5ftuyjZxTiD/rsYn3Ukd6XKHxNE3DnIxaD4BIKbh77PRWdNf/+mMg3Ujo2mqDZ
kPXthwFIiz4Nv+IutJIS3AUBVlgqJqB59nYBs/z11LqFL+oQksOxHdpjKtNC5tkMnCdGk/fsf0oW
u3tuJ1YY76G8Cx7FnZifyXKZKP2pNLxPotnNGlt2Ovuy4hFmBOpO0/rJzommTMq0X0+m1Rz4f2iV
0bufJQLwq18H24xq/1q4hipTmIsVn5T/1PIbCIdz/UIGYFJWcIN9m7afKSiFDmzdOr71Zb+DMho8
GYbsa+ShgEjvNBpsBUp2vlnufH5e7hbnGXV90yAejlzrSGgaUQFXImyY6RdJpJByf7vYIqduYcZ2
MMUU4nlYYG+46TM4rKEfwfXZxH+DkyPy3bzJ/0Q+qocKRfOhEY43793UhZLOzALhn8MZajQhWcK3
F6jc87gwY3L5F5H18oxKVDP81cYXOnPTLVIExWdRR2qz8FlSS7uoe9ghmMPXWCLTncsADK7czomt
C6gfMxxdvpaQmZhi84FdVmqUxlS+1jvvL1CggLEmsxbi/HTy+QcyMNV19usdePA3DwtPN70HkQby
+YUum17RPAVSxn4Uqz5Oso3VHVIniN+/vG2uErUHRSb0u8eMehv2jZWl//KX6vyCFyw64NNSqMFv
1Z6i6YpHHIH3e8Rk7B/DQjuheCX2Ar7s/Zepvyjwd9WAiYQ0A/YL31yBDY4cO2A+TDAm53n8P9Zn
G1cBGiGpvyAlYk3TPCoa+GVc+PYMWUO3Dvmk21FIrFr58zBcNYnMY/D3zhAoNrIJ3J1jQ7qrY+A0
/u4bhJp7W+djutKjjs5wwaNCBSCIHDePIUcimPBhKW/12wngeL2E9hbqkshNhLXjsUO/OHjf1zbV
pAtXBD4Gw+SgWb2OWUVT+Raxy/6tgbLKOciHJu9lBYFcb7NMiQr64x/Ld9o1r6emCiH4U/TjwGnm
+bwwASIeVqo9d2+b9DIh+rvwE+lago3nOItNnCeLE0HsXk4mdc9H+Q2fhUKyvwgnYCPHvkSD42/Z
rOiBVItoAf8hP3rjaWWS0qwp3ji2mI0dQiKWWqdKoyvjhIZsOPAuX1OuVgMWUuAa5SnPueuFySM8
TcFLCjroOZSSi/QMGRQZT7YEfrWflwolinlHoSTJNuh+aqM9itCTF75CdbDqkjQ1BaoZvZ+ZMyrB
2fFgfwpFz5omDY3SFu6VCj7UgUov6BJ/w/E+bK3DQp4a4u7XGYn2Ea56sgZMMBhvfo4AIpd2ugQk
mKWIlYCwDVb5lO31br0f4WFeBKVfSf9Td+X+S9OYAofpuK5WVL9KYArVKumBqKqgT8gGk83JnJRH
4dPaIL2VrC0B1r2GfXNH89IF0KIqqeoFoUtl96QR4fxTg4j+fqNxDLlywErt4M4kV9ABDmelIb2s
ImLK5IbDDp8+cVovMRU6a+73UYeFy7/aqq0nlQXepjFCLnmFIyFmlbr3+EQiQPzuaoKMEkClOwoD
akN/YPhzt/qjC1SBra7fCeWmRF05Pg5z3R+sZEYxndMsjV3VBR7W9QPk89JdSaoBhy8qwX3V3d1S
hI8NUMRSh2sBzSxr7zrZe1kodLYbYpFUcm1iArodiEiQJhq934+jikOWyfmfGersKURPE9HfU/xf
xaqmVzmFpzTbrG9Q7Bymn2FLuMLi7obx21j+X4U5qHIbHnhippjNY83QTyR45p6k4yn/8oTRTCpr
gaGEUQTxRfh9XvC/YYU4IuZ75pxbUmilVo5UM11nt75ONT/iYesROLueNSIs9HY/ZQfMNEIDSRMy
jOYObrJRo/zZlA+cMhAKdJBiioSIkotuvbO1j5TyjJo+LuOWk7aKle4Wq9M7BgDb2baBSJiDWPNJ
MXfsfC0Sqf97J1G10jjwk+F8o/yRHLZMniIufSCVzZPZh2tgUaybYjJ213JqE+JALP2dKHOhkvct
CID3tPlR8wYfWT6hfWFQpaQ/1DfBDvBJ5dPHLM+i48U2wfL+m5ZkLWXXh01LMLtDGSvPZBhTIb8v
/DmkvwWJgc1hL8zB9tExWczBnFCs48rCb763u8OZTVymK7fhWlu+OdhFYOR0pmpljKAtx8BCcGc1
CEYdDhWB8smajvXxn8RuIfd42QHYfEPbh+26zGXZHoxssAFO6M9BqihOvA3WqAYQ4FqTyKYsMvSb
lpqGp93ybz2TpwQAl/tWrRQV1j2vXTI8wVeiJ8cz11ckBXLkvKxLsGEkmYoeKGlSJisp9J6GgoyR
+RJDEb300aa7LR3vUUK0mWZH8LUtslz9GTo6YXFq/K4+A5gKdfWh0apH2IWWqjBkaytzpiok4mIk
ilrxSXh4cVAFZ9chalkhYT1FU67BqMUMTNw/3XzN+tqpx0GgrQ8nDgO4HkjRXLguTxrlqb7lIw6a
/sUysiqaweWpoQk38tcZxNLecbIMtZqPK4lw01DGQCZiypaExwPaKryaNYbiNrkkYXWd14qkrw63
OWanl+hSQZWZrxku9NG5FObwjavgbHsrgWFPc5wzGxJCeliLMz/3H2hbbTf2cFnZgNp7xN/i42P/
G6prq4sT/qDBTwy5XuUHIaByHDjuGC1MoAa8Hh2AJNb4bdTFHsKbrUhDW5EM9O+gRgUX/9NgS5tE
D2+dTaQFCroedgcqTFMWgRw456IUegvlvST6piFSnW5ATwM9JqA8tUBgtR39T2R/WIMqgUlbOiWd
Ge/5lT+8R1j0/axzgctE0854JAWubTzXtKdxNiwqD5/dd3kKWEBn76wO7tAzhDRpBHc36gpefzMx
s/S9xlb3yZ2DWlJBqJHF6ANuYF0KPtaNnyn66bvnQaYvcoIx5QX5rYcOwdwTjT2UQPSunCdQcIcq
4DCqhFZd6iacK0zAic73h3x7mkMVrV06GvHUCv15Z4dxV1Xp+G6joumVID4/u1GmGxG75MN3mkEQ
x6JRmTrxLVyF/8FebhoIC27gQq9HzK+I1Iu4dYk7HNInq/z7EjGb8b3IrowBEG6llYCSg3uxaPbW
T5PXFZAD10ZuRI1tGZtStIbnUgASkZZoL88pwumQvtkLI4qP+eBE5lJdWNicsnibpQaoHIXWwA8E
EU/TTRp9jika2Dx6kw6leyat6YwRojvTyWTiE9BHKtNecAtS/rTO2GiqWaI+0pJF8SL/2sfcZQke
U8VEcgF34deGq3Ycppj3+lkspkGznnvSnYGG0KocYgDTwFHNQurEixNmiUyfrZRkmMTdAPqMwhGz
FbuNyNBfJ6ts6g3s1vR3B+sTwXYBJIVHOcw5rN+GyjSaFECaqQ+yU0b44Y/0c01lZg5ICHzh/YXM
pFER5GHzq6BE5vtmii/slE+DPMjRbfsQm/tLKiXZBb2MSI/HF+2sMaM7bHdvYFnlXDKOniZhtHwo
5Cc8luqHT2Y2miyR7Yroef0xeL9Hhr9GhfTNUU6WSvn1txi1jmWiwI5a69oD2faotH8VUdJdo3yK
KDxTJ3nQQiPUkmwSRA0mN+BYRD0Bw9uHZ2STTIhjAAVpSBbmgt3O78cGUFo6b1PTh25RktK3yy4O
1AOpA+tUOM9CBiWxURN2FsYNScHstFMXqWSj2HStft65vglb9x/3pBywEb9T3heL50S6J430vLR6
84erEcE78VWIQFAq/FwrRWrUOvBMq2O0jf5ta+xfj/3OT+zbuKU8YDWvxjyzwRS/Ve89KF/ET5r4
5PVnMkEo1kemYWDsjjxP5zs1J2XPaNE0mzEW/7fTsKpMjshYCp+J2mYQDW1t3MB46CVaQH8+Wvun
1bLzqWf845aOQgXxG31L53XlSf6leDBqiYBFmdr6sZpCxMUJZmuF9pUFbqCCgmM3IADYHiUx/vl5
BlzYhi+HF9UF0k3960pi8BTWn5B0dI57IZ4Mz1VAHhexMd0Csqwdf6ptrFYlMvlhgwJCqYW4HjTE
AMrGbIgzBKtkvYnRKb3/kz2eF5w+BXelIW2eqP4XbABEpB5ZqRtCLF6D5d3dcXZc8SoRJ2tllgdw
BZhCLMf3keYQkNFb6iUetma54qJL1I7jpWBUVgdJoCzDMVXl5yrFRudIk2PzfYd1lALP3c8OfK5h
k5quzyjed7cx0D6K7DDtHxK7VN9jPTZYwyy3nH7ux84Hhx3+Pt+Jsbb5Lsph4/49CbVU2bgD9jwZ
2CWhLBXdqsdER6skDVEYG8B4/SPvtcRGjbm1ZslC3/CotcgAz2y2E6UJXJoKb2sDtjdAW+Qa3BLR
wssrJzChS8AnJPzY2VXOOHrLzqbrCHgn+mL8KA0iYQy/sJsvdZG6xDnfr+jaXCBnpgGYBK78kw0j
y1WVtesoPQ9KqGpbcbtwOf8sgNXiGJ8TM1+w1jiPg9Ad3Jmv7IIW8PHiJkctky9sk5NupYwVU2kq
CzXxjUDuq/Ym/p2fYo8ASs8p+OVwzDehKMzX7w7jlNMRhjJ0+ld8ygKHpNyIREYLGgN9bw0+YE6r
1yvIKjVn59kDyl/GOCghmiGrvGtE/wk7bRJJQr3QK5YucGVK8BwENmzHcm20SXrWzTSsmkxOvOqS
3e7xzgQgOYC+hNptMJH1/D98EYToL1ZdCIZSBB6oQYCKG92urPBkGbVMHRnx763IP6vCkipYYH3e
8DAh8sY3Jr915YImdTnCIYDvqKbDf91D5WWnUwf6VJ0YRb5qav4Vc2fnuLUG4a34dFj2gpN8ejzN
/VrXeLhkN6zWlBAlsgrueWHoZtj71p//bQ0YPclPVBjfb+Pn5S6CJU7HUL5hnPzrzO0TJP3wqqsT
fvEu5ANBFYBzHYj1mRJL0jFw25KPCStCE+N5b6xPt1YQZtoMLudJ2V6Xp3xZsoVExN9JJdo5fieR
CxsxS9jw5OWpDvv7WexNysE+Mp4QeCDT7y/N7QNQBVLQJAsuzSUY2LPc1QiykgbyrtArgQ24HWS4
b2hb+QSB9ecxC4Qq9S4x/LcaGnuLGbHsWt2wzDYQ4kbKaKfHHuq7zsyUK4RQ+rcB5KWATe/8C+ch
zEaO/mQzqw481I5JT9sUjRF0Rsf5IFZQ7DDf3gpwocQxvcGSS8MO6P5MBq/ZXCUPJJAktf1Au5Hk
MHzwS0y/PbP9kqxXkIbmVERXU1mwkt5XomvnZ8ZbT4NzpYQqQdlSVqVgIhfzIe+E42Hx8ypClAlH
GLIF7AzVfNVwpowtU0UkIuk2k7ZEFyOcyp62JfUz74HXSyKJeW58p4nH6TujQUC9PXDN5qPhiZF1
9WIo06SNsWZ5+nukL7wNQ9i422V4vwDtd/kDSwUX4sFqwiCkVGwinRbXAJcs+oshgxGMMDo6fNrJ
TCnTFvWhHIpgrNSVhNnbBnfw2bXnUt3bkSUwIH5FyNxtC81e6CdJpa5pTqAKPxrfIUpvWFS8Etg/
H9Wf/eiEi6g4toY3NwdyiSNhKQze2Sva1fatPC52ft5aXQbWUfrnLSW6Oa9gy+Yf0t+APZbs7FI8
kIMi7N1zcyhfwAwQ+/ylSgV5rns/kShGXTy1i3YbbF5IM0IrvFTnHDYOEGBArJxcl0QlAmhuJyC2
HmesuvyLq9DoWCF+X67RVsZV6FRDjw4R5LT8kZE8Bs9mEJNiRDPBlCIPqjyRUnrlkLh9u0iBHi+4
IVFzpFFypoqQFJ4NJSZno0c9dMOZ/IdHQYZYaAqhjNM20zvZG6PBm7T4YerLs6q7TKm1BwegOMXf
4/FvuhcmLbNifj9ZLiOcB52ssqWoFP9vj/e4zu0IH12rbaRB8D2Gwqfu584GY8ZyLmT9IKU7MUEI
PYXErUmfHlI2tmHluky3dvXqofNNLbX9m5DWn3zxCzD8dgv2T4vP/grOJ2wgU7MkCa/cidcNnYsD
tVQbzY9X2ITIwlfCleKyvS9MbX7/B53Cwtx8FLeQ2poeba3dEbE2OkHFkOn6tWUZ9lbN1oZeu0wV
0nEI37etU7ZqjzvfqYF+78eKMQq2/SnpG9909UdIq7YFsf56rX9NYRiAdWqSt0VlOh8M+qlB1CTL
1R8tvg3/hC0uTFEFwpi+J4YaKvrDndUlvx4wqhmzFnOZ7BLtc2rMbig3IoNoUJOXxMm9ztxRUMgB
7p2cwc5Hd19lQcNK6GPGjfVC29vyRZfAGGhV1s7x1amxfra+DebnxQXVRC2C2umL58XQOBmbKXLQ
pyUQgh1Un3P/Fmt8AGlhjod/0FaOAFRlClot4VoktbTfcuYxDfrHTgcOwAJFEVNyV2nwwfW4EJrn
jN3DBlFxh0laNtRmtjj//YmjnNKhuz3mP1VNjsBQzC8YSwjmpJ1pVQq8laVLnUeokXsat7zfVFX+
36od1zNZDtvhgeOmEDDWD+g754QUAZaCDsQrFt2lfhnXkyq9WPXaE4dwFBlEOxbL+oJdCoRLp1BG
z8wInPb//DB6CnFHjeCXbbZT9cb4YgryENqgQxwq2lajViXYlEGhPdWxyhN1p3nF0pT+m6d0Xyz2
sjT0Kz8OVOtapeFxXluKwle4aDsA0VSAjAD3Y8xQL77ZDbV4UPc4MYCkhFkg/vXcmXnLz7B85Vss
yRUyZEOeGw0FuCcHai/FNArJq3tqSK/XC/RGww0xECK3YFfFXxu1U8by9bkJe2p/DMD2c9q3uAum
PVdYGQOu8Vywi+w/Xnv5SsOtJWTCnET35lvHslUGHORanmN/3Od+rOcfRsJtuvi9qDw6qVa3uOUR
rUAYYW7FuCe9UouDrmCxvW/db4RzlvALcpBN9QWsnwXzlsmsAaUo2OsOFeYRRdjvQN3A0CsvpIW9
QlYDvWqbqYMJT8O0Jn5OU0DsU8auhsFylcQXwXDXkmzu8u/D24wX7o/3thPkuAPKd7c2fWM7zw82
y8PQ82bnHBMeg3lpiUQ/HjO4bLNy5bZOP1EkVTjJ+wlyNtIUbcqT8PitGaT2+8bKp5Kgy875Y/ux
KTXg2UL7Cuc+LwP3q3q8G8ukBNluJjMjML5idT7VR4xE37mKBJdUBCltB8Io32bQ3oYfAgaFgTKt
hjLiXCoEXME2HoLD5JMbSQIsmat1XKjxcO82KTvhNt+ZIG7xoPZ1iynFXsE8ca14S7Dw26gVQ8M8
hAB5NwlsOlYXhzRtXVWxkAhuOFcRONWhbyultu7lB/I8PD+IAt+LuY6q7LIeWDGydOpt7kH3D5OT
Xj1N0l1j+vVFP0fX7Wi1Zl+X7+KzfVqebmEncm3yWUQfbxNWCC8cvEo4dgxIWBFTqu6ZpUs0W2G8
TzE4G25zsGWZwyjpOOd5hqVdhRxmooQ0nDlbG+FwF83bGu2D6VXXFdzh47s+OmlCoUlKXnw/a5a0
ETtHuP2C8GXIt3Xsy2HYSOfvAirveJMI/tDUAhjCdt2cSv6CpC8tO8tRuw2p9ATCXhjuh3T2Y4pF
BEaaE9z7wP/RJovWV7q8LFB99n9xP1mG9ekL/eejuxIecYin8ua1zh+A8jh48eSniGrNCFLUOnks
QPlqTPkj95VA8oT7aVX8jLa4SO2CB6mhhX51kaPEwxY1MohzybAS64m1CTbYo0r5kPGOX0hlNzGO
DudwPyZpV/OmxEmz22gdS4ELWJWpK8na9eHyco1ZOVc6Den2hhVy6gILShF7Mj5fzpmV1ZHXOQ64
3uSHJQrMYGpi52pHHmPl/LRQXEf+WsjVxGubGy0kXf2mNUvIhW/ZV9Awt75LUpTrY1mIz1HMZgBa
bFw5CSq3t1zoPsDVLblAztpQda5kCOlt85F1qq/Q175zrfv7oRbhzxyHNr8K4i3srp3GIIuFliCh
Vio4VehPy9rOWNd97RKPSZQDBxjTexMXf+ZiBBThZoDc/6xkZEStmqKJbBqUQOs4x9Tf8L8oqU9K
7MBqqZNc+Akkuq7Br/XKAoVgvxxDH1t4l5G78TmQ5A+fl2kTyRjaZw57TY8xHl3N3vQL9YoVKYPa
xGWKA+I8RNyOieZKNgRY+ZEIA2+g04fc+qx68nKtvxDwk8+iT6or+r8wc36BmWMEJdYnRgNxT9f2
Y/rNuNBBoT2xc6ShbGKg+wCpd7+b2O5Vc4kNAZA15gf5kYl6A2MAo40iyZk6w2Z5XZhYqEwT+gPQ
bdBtHy3fQVR/VU0YFmzidGGv3zgnKwsuAJAtnZ9WQHlgbmnS1ivwctjVFwP31QldmDHaEgaZUiiV
2ZAmXW6sNqY4iwPTQ05wezynIotkh8GxiCakpzSJjarbEuSznCBZi7pRq16mbseheeAt0HB01X9/
GDPQ2zk8yuG9Nzfq4tC+1dF5FHsrgDOchkut7ft3mvQqUJ6o1E7jBJcXn2EFvuNgEqHbkp4hpj1M
dMp3oCRaEmx2ACt81W0WdpxgPTHgsSQSrt6mMuFZoGoFUT6VpHAS3YOz4/KjXhIh6GEGnVYPVP82
tTtfDxOQf6iN+xm9UuPbJzxGr4yy2OagRa6HSg2NFfvTiXsja1ioCO7zbVnZgwUgOLjJH5Wr7aWl
QVn+iyvFHt0Vbo12oYwBe16ltAgcAzDilnFOMAyDtSKBuNT6/l2dMkfXEAbGglEF3hJWzAQ1joYE
PfNxIQaTIpumGEwcmOEXSXZwOqrG6Fb1JP6wu5zDALwY4N1g25InH9m2CC9bDTROM2Yz5gzVqr0K
QfuHN2An+lszaDvdTg0MiGsnIFnugoW4OPZeeZRppqfRSVh95WqBV0DusxG0BDzB73OAQEjJDLz4
AnT3LpMkGtsAatJQA5JNupu2TNAk27VjBfrvMts3+NNw6uERr6yknKljlEj2xHOtFxQR8mc7GZQ6
Gk+b3ywVqOhcVOJuLXxVwfU1Ylapf4zAmb2xPIs/lsdmGL3l8qg5Vf6P/kBqCpKDb5rOapnZBjAC
e43Igb/VmWVVFTnYLZgonh71q5zThCLY+0/i/2AwxSQ3U+Xjm//fkGW9Z3E7dVh4YdDCFaDb6u0L
C14NCrN5YFjWJKSkmqvTskGd85qhPJUVwDK+4liurUp+Q/QfakZdXTFeyZqXj443ToKYyZ3QKu2Y
Pt3tgrhQJ57zdCv89uXZpeu5FTFEWinBVctOt8fNaIA6OXy29ESU9F620aK2yfl6E7rFJ5fRXIuT
8aahpMVr4x3mKbUtpgjVgL3ReMdLBvc9yCwfETrto3NIih0vAbAqdONiGYTliC11OUVajvJ1Fzhw
1nFNunND5lu7NsVx7cWTb1R4u8Opc4QNSKBHZf4oa4a21zO2udL4k3TvE0L2AnD0k2yskkGWZQvT
Vqm7v+aMOsG3T7rzfHnsQ+dlbtkKko3FCH5twETBY48v3fLQzUdeUR6pIF33pE/VXdx26qKX1Dms
A/jazRoFSafbhvcv/KBZb42yjGCx/r3meAI2+NCC5E/x5vKX4fZ/T5+E3Z+esmyTLQNqC5+efXaf
MEjklVcCYbv8Dczorwx2yrRbwgTkMunCI2eYfEUQ31cYJ1lKiribhpxiZvMnHoQHo1/hHfVlpsNo
iQm4WMgW86kVwPUNXukD31Qe62iHDXFyWN/4n1t1hyyGDUbM+xGOEC/99ydb2y69XtGWqY9Sho1i
EDDXEhkVZ+zuOhJFQ/tjZ0HvN4KW32W4J2rrmQ0BpI6c3/sJs9gBm8d9A6D8B7e6DmDNy3mJk7dc
vRDIOifBiC4iNcOwavnjlO8uGPSUNEKWHy98a88Wx5CkCDdegwZe7Gif/upHa8lPYAXMni68llJT
bigR69vP6gxpRk2GhLn4DwOnnhtceI00ifJzwkaGswZ9YIP2n5tkCBSljl7M4zmLKyI5y35d8jEF
7+VjXmtXtR5RjtH8sIQldO0gEGiKrx8PNu/Eukf+EQCg3ehiVnbBVZCpUNFFBefwGyv+hXVyeG0T
ZwL8aew0VmRsXNgLc9OcGU8xmlwS2HrvFer6dgBymFn5TJ4i/pQCQgqXnA6TiBp0sGoGFxeTofB+
mK9PDQyVvWwsIvDTk0SOXLYxXm+bk5UXcC8lxgDB19eJ2LXi5t2IOSKWIOAR43QZJ7SPg33U1wwG
PZgFoi0D9I2AA/n1hK3OaVLE5zRn7V2njVWJsoa1vwTsAU120mn6nETBTefDswKVSgrdPcSg+bPJ
UakfA0JtdQNxXMNkzSE60xgXZ80oXqLj4/6W1dO7pV91PX/Z5Tnj6vbTjTYCwVNavlTQyUl0NP6x
uDa6/Pd9rS7Xd0kxf9KXUbS0EidzbLdYpe+L9iRdf5JM970PpCyvRG4Ko/eeHz8bFyTLGs/K1Vl0
3H+x3PuyI7j9z1MAGs4PbBl+ep5sqauiMry+pJMFkxGVxP/QNhZzyV4A0yHn6ovwKewDvW02RCzP
BsGqmw63xcJXTInpQJK4LCBC/xWJvm8RgjDX//fAunRtaZsk9el5oGTUvuPGQ21CjgArysO0PCB/
Dok5OAmg3BFip+2Ky6IDj0FQPRd/WFCf28X7mHxcqS+QqCrKkduK8XD0ncnJgpF+A9zoi6hhaysj
u3CcD9c2+D1WLiNQeQXrzSR8tybmojY6/neL9t2WVmLe2EqRjzuGAclk9dtMuFAu4koK8EQR9IeE
YoOOldKj6XJ9eSfejZjP0iq3F/U+hElWIkyRcF/ASIT/y+XEg8ks7ZXS78DoE+ACYaF5tZtmoIcX
ZKBSyTIXegeYp6/xoWNK+KOOBA961sedA5jMI8SFjZo0aZH7n3Pos3fsz4KobYsj5HRlqfj0/vsp
gcn7Tmzz+vy+0u6/XLs3a1Fp3ILr8HidnaSUmP9Z7T1xaUO2huT1b68c5W4lZ23H3Opj4Qr9/KtY
qlvcCRp+QsOEmLbMKmsMh7X/ovNHgwfZ5PlW96QvdLUBZ/as+FzlLl5NENCr4694Z6bCs0rb9UkA
mAGcgSCY4TA9Xtpm/XSUA37GIwA4R8brjTpg0KDXg3egQBIIWvgKKobms9gk80FKxYinyh4g3Tn3
xHpcqxf3GfDuO4yBYjX/57ATUK4UzDwMv2zog12G5/shdrPgKUPzbCObA8ih/C/YFnylI16Ghsr1
mUfukVsi/4Z3eZy5eLy4JcxPR83wfNGnAb3nAYDZUDZBqgMraNTfcHD+ZR+WarPIS19gFzSB2+dA
8tcvgz3/UhdH4tzVkpciMTwiEKiopSdXaQQQSpsV1wH5c7bGHCsiglGJOMn0dljtuYyPHFLktF45
DhovLlxE/ufC6SyVFwgtvmoxab8K5oFAPNOmSpknWrWRKmMpiGQeNfJuNncggeX4gHiD4GpZDoz6
KyedZTsvDII7gS3i0scWgCyCSQwTxjN4PMgx6GIGppFJk6/6sna2MnfxENnT1AbRGbo9Q2W/HJVH
uuCh7adyy5Re6W7P5va+HGSPuGeH+HzpVo+ePlS6psw5ZR3LfunXJpuUVsOymrRwz8aB+TrJ2pJP
zfZre2+br5F9+yaKi+rN6VOjkeLhmU1b9A/wP3Z6WxcCuIeM1j90RIVIt2dePuXEsV6IE2e9bBqL
tpbG0/9ux9faGk4fbF2glH/fgoVhVzhjqvhw1lNwh1ulPJ5X9+qeF1iXNjV1ychAznMq8P+QS4YV
DPjPmRSP+pGvT2lXcZfAlDkMRrOqqKzCh8xejHrf01eUtFt6LBDB3B/wl64FsxCsmJRQD1TMnsoU
ycmUTss+/i9kIzsZOMvgTti+k5eU3MyIrFv2CHQ3Efo+0v3M/fpv7Pdmg7o0oe6sD1+3YkPJomdl
4DEM4xIePNLVYX5UNySC9eGY9toR7fX2iwBuZV/JHNTKOlPpmllRO0JLFQGo5XZYqLijcMB/x4//
IPL1dmtVRaxYarmDfh6pC/AhTGj8dpM2Vgpc7pnmAHV6lu1ktQRwGTgsdQUZII0tsiF6TAVSBQ0V
eKL8/mLBOA3vagzP59lMYKemCGQTvoihZLQWy8KHifM760nZ4Bf4gZg2vIR966HI/DclmfspVeyQ
mlpJtoFY93q6Il+nU4w2zKUrizlWOQjNk5S7Skx9TRmFPEpQCxyjhSvdSMtt3cfCODsmTTJvL4DH
ZVHkv6+FBXzcCX4mDefAF+iF1VnLIUYq8CQwDZ3g63BzzzCnImTDH5h9D/CCqzCyjLywEq8a6eU6
VM7JlsXkQQeVWmBlVPgKk1HXstvikqMuHAEuaqrluYqKdFX7qIX7EbEeKI/3i+qKtrGiK+WH4qKw
Ja9St3p/RNXLC8YAxmxeG39cb1aYaHDaLfZ8yuyTcoq4Z1MfeecvPT0x+mKmf/Zi05iX+iRVnDPt
eAD+cpp0Z4/jN+Cquz0iKPSY+JBXMW9X9iRj53KJdTfynnf0nCU3IXVZCbGX+h8/WhF5E/LLqa9X
cwmplAdKEQM3O20CodUpehNxQNT8fs/TSmf5q842PjhRIUlQP+AZDy5iuHztiwDD+rMWM858z4es
mb3ZIdRaPp13CK7uPjY1BVST2jXCrVqLtG6XpDk5ok9Oc59nvaY2NjPynvli5dcsiqJ/xM4tQYuw
GFLIpeBGuaykFgl85VjNPOzm5YYD18NfGqlg+89Gz4AjDDi34LYXbzb7g/6mMp2165cMeeOWwzeq
Gh9hoxVft0YTkPVa2pvYZNOyvaLE8d0algFiCFhw0j/C2SnjuiZVWMcokRl9VZHqMb0Dxzv8zdoK
Pj2OOi2Uv6xkTl13WRWsGCra+976Ql6BMlozp8sXdw30AImACpAYG8uOMsDvZ5QBWgeiJZOeGPZn
80yZlJJCyU7J7uBt5GCgXxAWkPvfe3N/kB2XUTvlqL77x59x5ywsgRuxCMYJTx+c1CGo6cQCWxyY
7clqNAbi2lF0FYTEQMIPotqE3yVYnxZds16z57r/Yu7OswNmNGIYqCzWNrdXhMD8uTHIiMWFDFST
Nxh1ilDu2LnAxBqN3PM/ZeF5sRUu+K1KlQFRSIBgT6anjtsdlsTi0nqXwXoBCCm0Rryxsuy41AjX
++oY1DuL5wGhjCfeuvYIHZZUlAspMadUY2l33nazSc88spPXhiI8/wRVdc2AFmfustZql8BKELkV
KlmCVJIAiqHUIfzIrN6IsIIisGIq0mmqN2bOGq01U5JCrmgCoYvmpEHTjxOeHVA50wqF0o8HbTh+
and/V5JmftmFsuQ6E32Mcc7cGEatW7ZKsudHe2nHXhBfpjdm4RKj2rqeSgc84XkcM713qkbfDk8W
5d1pblsKgfURdMp4+tMerwhCCmX+YcZucVgWLxtXhJbAN2Yt935BxiHd+R90vDG73jZwn7GhEJlV
kEyTHZLgb5949rpStce7fv7SiSabsrsbo4pEw5FnLrFdawu1GYOtMWxN2hNfajzwgzNccA8jdXl1
cBwlGTlIwvfBYnFVHh3Ej5FT0bMXSYRUbkrn0DNi/ub+u5SMwlOShuEZgiM6q3omfMV6yBiNdd2E
LIrDXEY43uNDVll3DY273x9cbAFKtDbO4LxjIP6RDhPwegnYnHnbJLC7Zm7m6fSIX84Cx65wmhd/
pGJmCe5TMYlY5gHec8goZaAsGg5MZC223c+e6ux4hElkwLJnwvAuz5x/ZYkbx7xJ3ECq3OFLeQy2
RAMuRdPYjH4rvF8kVAp0PnfhCBIhNAJXBsRusb86KjW0cRBk42xl23raeIzMPqcn+8HIH1T6SSnY
x6QvgZkhRtJu9eDPQu6sWYLHG52RG40iMTxdxDFvznR4+Dtge7q1NzC8zcbOH1ZzLGZVj8PdzLR+
2BlLqEen0KTrsAbOhVcnZSgjqTYg6Cd9pouvIfzqX3Ou6+y5Ba4RpPFuO4aBOxkPIN9P1jQ6H5ut
WYK8E8L/hMciKsKfU6QwkJwcVUp4d/BWxzQULeWhxbmI9ZMsr8ZO4VEf0a9iEWFwyfwAbX5dS/br
Wn8EOFh4rmsndEc+lIGaTkAPGFAUzJ0YX6G7ymeWQCywjPk9YKWbX3bzZUlzrF+JAzBM7PVumHqR
rWfrFf9zdxIhN4652Cd2GoTATc2rQV01PnfF3Ma3sDvcLl1perPJRloos4rJWuPyj9tYuz8fmVML
nt1arIqjIz314yboel0p8+HC4QCAPvWAnIcCg+SDuTFAeQnsDOgAnV+VSzsrekMu8uKx3kffv0RF
xRVH0kpcAghy5eoKeXx+837VUgeE3AEJfO1+vEsfF1b3oaKCAansHU7MfjQZUNQICP6k6OHoEQP5
6jd2QMn37fohjUBOghrnWnq4HJ945amrvObRpv8ZfVmKL2jW2mTvyAjK7s2Gp6EwkOPZI2NfgcaS
SxyXJXIWN7ou0bQlJQBTclIDBZM6CoeHiEHujvJwWLnfZCNNxCkoCSeOCl6kQJYE/OevXUESrWOl
SjwM4nAG3reB9vHRx23JuxqsyqL5GnPofR/ad/UyATvGVJNNtn4F9TzRNHfKd1Csn92gj8cSQSfk
6U5OITUpZZ7CaTsj9EIsMjbjWuMMH2ztTRNOeNmwBKlC7p96ft0DGtJtrNvd+KSUe9I0cOxp4SpJ
UmNbBTyvdGoyfvnqqAyZQSeCB2POlbfE08zqiSzt9q1vP9NnMbnG26qL+ghhC/fM+yilZHNROzfj
d+ooZPWQtBek20RGTv1iss2H55wcoc2UWm+QcQ3QGeD5cezR5CGlMm/SczpRwLnymfzon1qBPAM2
9qaacInaKnuJR09YsmOjDjmdm9S1jCI6M/XzirBhPprcgdXazPsSWb1iu7aB/5gAHDiHIhQ/rktl
JAetSr2vxjf377JoPjK7i8YwQLOUfLXi+hFJtXa8RBgR02n+3JRU0Q8lR3JDK8gWnmnfFv64bWme
d+JFixkevD486+5SGGvXLZtPiqPZq7nJgcU8bQ5EY/Q+qUs+lIypyEY2M2YbyzegwSeEm8rbXs/N
icA4xyMvynx9fvSBAInBQ2Cc6K5E5mJ67+jZWV0VabLT7HpncR5htUtKseNeAVfM44AeGLLdZfgE
375skQikfkh2OmiRBOSHCy+RJ5Vd2ci5/ak5C677IiMEV9lUf6zwRLgC8g3KZcerphVjzC9F8C61
YEbrpn19qRq6q1kzqfngmiLKTX7CdpJTV8v4ab4WyGbg+i/PYxes8SgFa0VeuIdZu1iXIVbM8Bhy
/jsp6moOYzK3i70STaF3c63EvzyGsEngPOyWsKeQ/QUhByIKrTEssfjD+gbAzJupKVSdFH9J6hRO
bLUlJ220eTLsVAk9PqJ8+sPailA/HFvZlBDVfwo8U1mK/RFA7UalpT8sBTE4x7ksN+szhG6OUVY1
qajuDihqJjiQupIo4l7OR4e9gesOF3PjzTlYrmKnV+FFZlW9ciCGFGCnnhMMSe3YGCyLia8p0ZYY
0b3u5EgrRrxX7qmysw7HtQgJPmek+onbjE3XiOfWb4u7inwPiTATD4prrWd7V4ZSkPXrU18FlfIG
4IJ/O7EeVzHplS56fn7WabTmN7tC3FqUciNM5GDNTGDEN9IYXfOf4jCuz0kXiSpEN/GKgs8uYV2+
ZYhI225+R/lgPx4pvrDZuCOm8JhgNwvgB2lQxZCKC/dth7PZwvnYzDzKsXAjZpHNtg4+1o8P8yCG
NnHkdZm+Mn4QzmxVCEjitzR8vN6oTAh+kkglVYnV5s6E61ZTB+x9KOhQsl2StRZRkiRsZC1TD8jM
u+FYqVqetEajWbl7t645+seyBpCb3FvRrvwBIbahEiozOsAiODMouI66VjtpMijnAH0SB20sSBMh
6VtA43MWd+FfeDN2cTeeno43Pks/JS4TbUBn5/oMIwKmYGPfSEFGt6SZPYgLuPEj1JokIOceaiRd
B8vLbGs3JYmJCBq2m6EALKCqFEqQ62WZO0git6BKCvKiz53I2srUeuo1DALFGcX7Q4wzuq+Gn8Dw
buZtdfFA60VF8JGB95JiVQ9V2EfHwGadibZLZTCz/TPdefhgcagMPjOubLjd+yMsLQApiR3Xm+cp
wCYKvply3fra5aP4GHX/iOGUNx9UKknT7xY2AMl/gp2MtSeFlpbxUvaQXwsXbdIxlHByWmxpXIBR
1CE9YfAW8YFlyFjnsGsmgjOcTgCa+ydNl3xE13vA1xWWZ04Raj+bmU3CCxJMYwtvy2xhX3T+4fwH
xqgISgUeg4be3OXH4BJ5cAVTtu7E1KkrwomTiNyBM7rYZIzVuHY0E3iL71Rg+eadwdw+J7J3XGuG
k8kogp+tNxcEoX2BQjwdMwba/achFpq8zImjdxmBxk7nzV3zSbqlCHM5oOIOW4g7KCLfStHCIYjU
L43KOyEGkspnzfuUYKkVARRaMrCbY8JEiB8XXhK+S2NdIksh7mgXExTXxBZZrdyBMFjMSDqTmBRx
3JC5vzRqhDMMzIpXLnm5vlJpxwx3rCt5OVgGC9017O5pxVbHBDFlxLpY/oH3Q3/v81NHlr2xmpve
MsXL6qJbukRDtAb8gnodC+BKtQwLksFhkz1/ox4W3isoltafDckXt/uQq4+0bUSCsCxOsnvDykVJ
JSXdOaleLFD6ZWg8zN2eJx1V5K51TXkBXf632x2a3MIIUBWCsPSi9DH1hYKyTbs3hwyvAOLCU4kT
0Vbkj1NdyT6xebAIEAuBCXPYMOhpjOnFq0Lm1s8YgfqEK4fROKsEXe2lMULxUjIADft+qNxsy7pP
tfzCz5IAZf78ccUD3FoaaBEUGhP5CzHw2ijaEkpfUuR7EgxV097ufsP1dIUxPa2jQMxoFouKHqRd
aVh5HYW2kwgmJuspLvmi1yffEJrMg+/5/ytIo5s6dLOCHzz0jnt8R8ysAqaLgBcKLCh0E+wgOLNv
0Qd1Er+ouZUxZclTt/9pecbIc31Cnhwa5BfDjFBjx/wvFox7iaOeqThytQTN4F6tXY4dSgx0ODrl
MQH86myd7QSwKLu36v/wauVVcRgRKlhePc7NUXsudE5KRZBzCq+w+alXqO6IjqiHtHg2b9i0vIMC
gSCofR/f65HJE3sOqIKaXkFf0E3YbPt7kzrlHH1L5gZQOw2X333mEoBF8EkPJfGbQ4Lg+jtNNglj
Akm+Tz21oYPXMYcsahIeaVarDiA7uFg7LfWqrOMvO5Ifs44LfNyARzvJN1Ct/uR049hW8zsO9fP4
pGUzP4e+RGUSWqs68ocPPfwLIjwgYTMU+ec7thrXV/yAyFaoZWnMytLQRxW2ajvKuEsL46uxdJDN
/h9lDGWUxMxgaZ3wie1LOHz4+8qLPtxnro3b5lX8iaVbVD1ueFgTlCeLhWFYysGkBiqGdUpYqj1R
XQS5HCIytbO1OJThaO1NVZqF9MFU1NxeFzmHE/Uu7KsnIyAZrkWHIJ3D+oz1Hgz5awL3XkLp2uK7
9+Id0yHiDbSUxmU7UAHQB4ttYH3hKJ8SdDgIuRMZOUnGVxTGpNl5VDCDpvBDrvZCwncHck/T3/GI
aCRzGUTOUw+SAiaEkGsAqUX9/pJp1CM2pF18oZh+6cq2rWR8x6QsHqpvp6GWIOMe+FTm5bPxQfZr
ZJHb4N4ZglIKszWF0er7U+byMmYwR0HkblYrhn0g6csDxDwcOsJ2dNVUn8kofVsPpS6tTspq4JWN
KLqo5J52Y16bv3CtpSBx/c1ZnCahLWyJiukc8VIXHvFkSdKE0jyHjsKiRCnYOjEDnffUFmPen6JT
A4EHQ1feCj4VPw6E9P5Q0ThG8OxbkPSBkgTReI+KuCn9ITAnlH020kNboZJrKtSE9SV6C8pfYSOr
1k0plnGTd++vzNtp9RQovH9i66EBIJonF4aRa29KR/O4H1HalcrZVnM5QtKjDQVh6ru3nlK2OBLh
eLzqScQev4Bhn2fiduFwyr6I65SWA5tlrFiz869l2R1A1nMWJ02NQI40uo8Dh22TozMPyVgCzHWf
60x2KlX8UQ2brakCu+YVBwEnoHEKFe6Yg14p/i20980+kCQbQzX9E50KxxH9NPQyDS6Rx+pX4OQo
leUWLJi8Nd0cCBHGx4H1um/QJNP0ga5DlLIL1PiqMn0MO8S8609cqSQbW0pacg6mBbMyl21PXQPo
Ui9LbjMkPeQQ1K5mp9mih+m7T1iHes3QHDluIqaXOLFwIrIvaGtAq4K+17WV9Cf7mxCXNM7a2Dce
Qy1SjFW/etNHpQ6nY0Lo1Iyw4OUYKd4Yx/Ew018W+FfCO2xIz7g5yoPe7tE2+eu0UgqMUiTxytrg
jnymnIHF0cXzK7mZRIAGCA7Fx2P17kzXuKgxTKoQbV/tUlrJhLq/VL+mj7Yaw/2wYcnk/cYkXWnc
/Fdl1R7frCqzKGyuOlW7Ej+2ZmXYnE/ahQairC6HW9ZPpi+hGpSiv10ko6YQUtt1QeQ+nuf6FG60
TlOMQSyVH6Wts7zFCX4xOHwC/I5DlYFiHa51qmoD2YYI0TXoNm492K1CwToDPDWYhfsWBpSV5b0i
T/AYqU4brKZvMp5tGF64FO2LXRwlwKItQ3FOc0J7AbRfogWs+Vt2VfRGR17aUoF4bSpZIwR5J6UQ
+h0SAGNYRbDn5tLrsE7xBgn9mpFPwytPK6Z92UfzQ28oWFB3t3FR5fC6N2UCtNzRAwiiFEsqD3Cg
5UCyrw0t59CjwVi7xTdlLKx8ZYERKSLCyI39FzIXss9+2/U6xL6QTfNyM3UUvIEbyp8O+vAMKXuQ
7cUargyXICwsY7nnIUQhOsSPktlRyfmDaduX3YzojoVY3wOVTcCA4rbjcl+AXuvHLIKSZn5NQwRd
/BKPENgAPRFsY9yzLYfO7mod3bvDhIg3iooIjJL2xBv36CbAe1RYtHZOvxBCyYLHqbdAFqKnFD/f
HulO16EXB+pk7Gn3huMn+h3F3TCPyucucHT3EcCkku+plvcpSxhtPhlU5Txe19XnV7gEKe07SBdr
svwgMAP4+EegHQv36KqRys/s0ojZRds9AWbXScIXiF5b/wiBVrFm3lMnBVaBP/3mIYisOnkamVHD
b3WcZBV47K8QT/6C2Re6tFohZFS+TuwExZzvs8oN+zRqdXRKGyEc3ZPh0oURmpLmd12Y6cNh48tY
cngknGmFS6msJhFQ7G67j8bsUXmpl/fgrDZbR/zsDgwDpmFA+mPsOi4RUexO8G4S1fSvnhbZYSm5
cqcWqL1hx18fSA7y1/iA+ZhJ70X/qqDxkXmLXXWb2wGbVqNobJEu5Pf66olQyPPQSTvtc4Ogz3be
ToOJwMVlXCjr4XLzIixbys+zNkuuNOnt4Ag0WGhobf6yt5UYEyuGlDtfhEZ90CRPLP3yhh8T1Xif
7zt2cQJ+mo4WLTDEei0+nmuGH1NOiaLadizUTYLY6JW4gIxAa+RUeR32nIzk7e4zCdoQOQEjU+cL
hCsQh19aT75nw6jzb5DkvAtCBPEXnu0hs3mg9JHzFSwd4jV8QNDhahaU0xC4wDne6JhKgBDyAI8o
5VtOtvl8V8rdDvIoqZs/XtoWVLvGiwF7AAy80CfqKSyO6DOaJLc5F1fHmtOWrJWmORItH5hpO9Zz
6sSvBp9MXW+zX3GrnBCcSJt9fDymxJeLryKa3KPu4ckMu7MByBJ5H2qDf2u2jLeykOoNb+xlXS8G
rfQ4FH2ouhwq04DnZVYs/YoqSna6+9upfw4eO4y5wxhDcXyHeOG8SaBAu36NkSEnTPbCJfRc2PvW
Az6/iu7fOXKG4yoM67EQsrCTgQKNOhmUJdgVJLNCUnk/TTqFv3hjoUrlnj2VdGJkiBx770J/un92
gpQR5c9GEX3uAOfrnYzM1FvRCBzg4G+sGKDU8DFyf+gc0Cj7NW1o+9CzBEOXF9jZWaz/ISFRyMo9
f5K25tzWoy4EBNOG0jMUkgt7Yz+j2+aUOOd9Cc4hrzGb5ezLORklRRfhLs9GvuzmpBCvZNy8xY6E
UOmnH6o8tUa0Bh35oIGPzsP8Vqgsra8Tylnp3O9WzX08mrh9OtauIRK3Yw55PQKeYVrB6KzxNKA8
Ge1l4PIteWjejI4vUvoqAP4+mgjkMKsMq8ieTS2Cy+HDSHWbdd226ImySo2EAOBQ0eJEnouTRGnR
jChX7b980+BEMkC2y9iszibYMMhlEygzUcLbfSSk7mFqyNT7ef5eILt9DOm1lijxtSTxNBn419Ii
0mJ9fV2F3UpUUFLyfLxxgVOF9FMlvtLuOa1kB5N+H22q1cLUkVAwPd0waj7O3KzsZ6q8KdnqNS0z
FBiCrNP8s+zqmS+AD5QsuYZFbX/jCJijo5mulBt3hzb9VS9gZdY44FnO/atXhcivhhLoxKhDcxQp
XN1uuzStRYJdrI99JUWRMK5qAE/K79ANP2Dua5Q/k+ATFXPJjVLmJQim983ozWSZiJbzi9ovquNx
UTbRtYrqKhQMn5/ZFBZvPeoHNcTsatXDBj4BnZccmvOkOGbgPMjT7lwo48pVnIrmqmOibKb7ZCol
/uOIJ0s0N1q52wgbwnqK6wwLVjyl0OvS0LtRliuGRZKrCl9NTb3FmaLwH0WJy2/hl7nUrAk1IXKU
sxbeahx06/RWd2glYKppDGYpyZC3o+uL8v+YrK3MSQIO2wWa8bZkT3p+xYh2Je8eJaPTGik2j+uk
EAJf7FxOPV6Yv8FjNZBM9zeus7pAeo5dFZemkcxi8MLQT2h6UhYXJONeUNSEOAd+8+JAjOVSztJB
SLbhf7UUYMvjfJ+UyMpD52OVhWwt/ae02ElU8WwniP1445rQOXmqCF4YnzOfxh87qJPHKlTEsLB0
/GJt6WTRDlKdzoVNnzy+Gd+b7j95xj+zN7+LUM+G1zgVz7H9tY6z4LBJGE2P8cV4Z/8wlwDmtLwF
I5lyN84bpBzIBoHaljSaaSkEPuEt0bBZcaQ8O76aI196zTyQM/DowrQhF+wJEk4BfBuVaI/kARMd
6STf5FxVvOBIx+dtXJ6/NKAwJFXVXabOKUpam0TgAUlkZEWS4/RNvo4524J/Zkbqd7dzD/2MU429
aKxoSJip0YDHCFDcK2KqNhR7nm9Zp4Css2HoSoDcziVsqUBa18rhdlRQJpmu/fql1PHgeaD6RQ2Z
me7Qh7T50nup9uZ00hxxMUgnQ73rfaHhyv1JHSUsJNfgCdEgYGTOmlvPD6PoEm0OHJcRXI7bGSNt
Znnq4H/+rw3XCKBtaFNX7R/F+VErmv7dsOdnPHzXnUXGNdUbhJzThy+V5sRaS2XnY6O2Dx4x0PQE
c+HKK+k+MnN+CdRDen4ygOXkTFHS6QllR4QipGhBUW77b6F/oBPnePF6geiNf4mPLKRiiq46BCYi
eA/lSFS95ok0iPRWW3XCc5D5TULGxL3Fr/D8HhDBNeIBZLuJQ7o/FMlh4Wn0E5hHcGZ2BxgIjTMj
wPSaD8XHVfjtGtXvoZj+/UDztJzk8z+9M1eNJyVy343+2vOqd0H2x6o6q9Fi1osqYjkwlhuFpqey
mgnDFj6pk8diAyhT7rTSUFPDusz+T1m94KuMC7mtNcm+eXwxS4gLmOAkOYhzOQHDTChM/v4TFJ6S
sBKehFvzxcPen5PXLU8w9f3pX+x3GsXC8vLaD2Ln10sAvi+phRh0dPDg0/eoV/c1YbF0RCCi96Nu
RxupU0Vop3fb9Dk8XgJ0SbX4wqyc8IPQHQJxItAPv/dNAqEshHPuv5wXyDKxpJSCmMKrOZJ5XLF5
AX8HFsNivNxk9LN0aFYgYcZZFXI6U2qYAJM9y2OmSXZEtx6QeXeSMZEZArc5NFp3DIf8GpH8U7jS
ljoE3iLZG2ooaZLBLpWiaW5WjueBYNHGF+6G4zYxqddwFK+WMoyWEa8VMY21A3P8uE78zvaRCEPS
xz0lUOT/N5vMOwFlZXPOG0KFMHD2tqzNhNl4/5UB/opSkWOAZzBZeVszUgKrPpnOeOQ3Rr1NzhVD
Ic+xZUWWycDzvA84So0YLJCJCov22X24NZN8bIT8i1UrdEWU+ge6IMCVMP795Oh6RL+5V8DOKdsA
MYzPxujOyM5p/uFDXPVLdhzaWklLwFux0HNiigIzYC13SHmlWLDaOi1Xq63lB5T3tXstk0DWsBkM
ZACRU3SYoISYrqg3m+MB9m0pr2bgNNKEuuINARqQsMMKnro4J5BOvIQWEStCWkTFhbeQ29YlZDsW
IiFnBYfdZbF6Bl7Ovr2E6mOLwecX91SLqlzVu3RiJbbaTZp+GXCDTb17E8bk+YZhXtbqdB2pGenR
tyNqcOpqaFi5HTKPwgm/KvRH+FH1k/zxFbg+iMXQordWRhg4sN9QIP+gftUrXFhciIerGA3OAs5+
RK4GTLdIiy7YkaOtTtg1lNmXrd5b/clrnChkZkx/StLL62QXUS7uHzirv6KxpTXUwqY5KnosYTH8
LhHO5dRgu0B2a8jwrWFH0CDtfpejSjReIv91711vny/PZCk9OOoqyq7u/PJxNVlxBU3k3c0FT8gp
dLLzz4zVhyx9hBQAcuhd7ULMCuRmp+VZEly3X2OTI4LRObiELZqdf7yVbxPWdB4qwKn3tN7/34/B
FZBH6S4zV6d6dKsCZW7e3cH1iUbWF7fvHsB+BE7wA1+eMxA8YaXUsUdOS/L03uY4hlguYRG4FAz5
kcr1dRDhKn7kc/cSRKyHQmLCTcxZXFCr6+4ZGTewUI3Xzw7Eyr5MIeTCP4FOYuTYcz05uMEY2Rrd
+ximufhPW3o7AijJ7zlAiczpmSa1mZNptYsVjT/2EOT2CpiapDQMMfe7Gv1rKgxPhQ8sODKJjKXz
olqgAexdExYHO2fLibwKvkscgck/NEXHMNnwNmhXzHKXv50BSXk2ccRdCR0kv0Ab2dnUaycVtj3G
KIkkmb+IsukIj0Gln3bYBE4c9YjoAh5p9VeEu70L8S2kGHbQzoeoPCgj/jDpRvaYLinWTFJ1H8p+
9WfGU9S8a/wNPIpmqiWwgcJwa/OBsO5G/hB21Vxbkiwt97xn4hkzvP8AffcexkihCWHb+Rv89vX9
XyIe5IjJHCH1WU159H3ALlAeCEpPDG5tj2u2A+zF4bvgROkEnAF46k9wToOBfhJNZUSWOxMrNWwB
iEKEvfopLZm0ReH+Yi2aEdgggCKUl/FChXPs0igj0S/fxKof2WhZNTGZl4tf81gcm7NidIDEimXS
ZUKSCavlYsxNeJg8ncuVgAkkwLfZrt9XmUzhHU5BWnq7J/1mGrFXurmRzbw7yJ7i2t977uXv9kS2
DR1b5ztPvUcs10sNilA26Sa1/FBvs53ducwRNVmPH7fIF4AGa8/CKgvlCaDiCIpVkKuzBKtktX2J
oss8/zWLASxg04pDWEA0boON5nAwjrmhkBO2mvJpvmj2qkb88KlZN1jllo47QWbZxKng2L/cn6uU
mq7NVl34/vEIEPXYZYsD7y6/ZbTO4Y79p7CQXRWTttBIhRVxw9ECpgHeYevhdnAG5BdswfRSSlTp
xt7AsNYfMt3vbHvCpFKaJdRJBeZQtSicYxiI5wl0iJb0N/7H5WAgndJ21WKJr9BQ6siHRfg3AiO0
SCqQ2lJ2NfE1lkFwP9YDtGRj14vDVeKytslO3WLYnf/5QLgcjyRwR0EwM6A4v22CF7T19En066UT
3PuSeC9Vcx/Lzm+bu0Tq2rOajcZf36AhHIGyQ+zwgr9Sm42tWS9krWqddJaPr2KG04NvYpJuIOUE
c2BnoMKkqoVUtaeFC+Kvn26nS5QkwWkajqmluwTCAz3dH9AOC4ns3kQIs6KnqwZK3Li56aN1PMjg
2vhSz+hBc3cYfxxgS0SbxWDKTmEbE/a2yThiGJ/p7X6TaDJpdvF9WBOslP0uC0FK9sIw2nrnWosE
EWITfVu2kNCoCjzxP4fPG4gNqWDfTpUbc2K7AGPn+lk6UWpMvXK0CkQa1C3u/fMVF9RnPItljzMW
2a7S3Thujm5qdf67LJ9ohQKwOI7K5xcTK4CF40VR3dDcUglGn4k9YxaeQ4Ll124ciPP5F0InWW3J
7qfpoVFw0MuPkiGFWD46m4r1NE9Cl4EDQBIz9kOqn2sB7vjBKVgsuOK0ChPQTwfOYGqJlgYQKdpA
rjcLPvUf+MUBoKiGe/DJcPyxkIso4Nd8GK5Q0/U4HBqU2spTjrWlboRbb5UZXrAQK7O2acYZ54b3
g77pPxTthUOs6iw5D014yv0R7buG5/X6VogVBZ30pA1RKRZp0q+SC8/IhP9xVyY25fVs3ZRZxcck
D/RvzhHaYb0wX4RCnc8qsmBqr4D6ljmwObaUcBNOYNNJzia51qCIDxLuoKCZPlXZzJjg+N4hHRG2
Fq4Wu89J2qN886ITVHgWOisAFKaZGhXNb2Im4L1FpMi7kGQNiEJpiGUvc5wuc2VSE3U74B4iqZOP
kjCkNa07iLMHCt+/htWm+lphJe9JF2VfdK2gbiP67s9+wfySAx/gYDFqXdHOWfMYsVM1m5yply+1
X0Ba2NHcYnksJnOcBpON/822CPwLrwYbl3xIXu3+PvMtOqWhtBjLHtxYZnokk3Fx+oH5ied7JGaI
DJKmPJOiu2IZ8bajrmzQDWZHfZaUsdnPN6bNaGF+J0lDTfZPO5Fl9kLG9umLfyEtaFxTSt3HKkfk
kE79cKF+uT+JxDPqe26GHL8qZuy+1MUDDDW4qjR1rX9M/DJNLbDIrSfq+Utig1bLF8V+UvnopKE1
9My1lZf8yG1wO7siCEh3335cHBGvS7etIJVhY+dX6CzpzIptIlF0P46mUy3fnUBfEh1fNeJQTQg3
u7OPKdAD7CxP0lJr7UyKZPh+fchQtFYBHo0aUnvuOmLSr4pb0JoFKhbyKMbwYY6ecXKuA//yXOMO
QkeVo2hZQgixRZtC+a3KvRaCL3Zf1gewwG2k66dMnNeT2le8yI3bEFcx7o19wm76Qi+s3Psl+qFN
Ld+282ArByO00WqQD7ew/TMDA8pMREpMPf3iBsi7kCRocu3iPuJEol/y+8qLpD8+h+ohDQIqcZz+
ArIfakAl7K7kCIyGZG+ZrdXUTWw8KGGzSFwN6pOcUhA0foSXqdoMxr5YAZRS791nTuNPyNvMSCDi
skc2s9GAcOl4GOQ6CbfSK0PqgcRJLDcnq6bBbFwMHVSvh5Y9atwYGwf3fOSqQvXBT3/i4lMbe0TU
mQRONzMAoSbHSBg1AZM+YBvKUtutGHlge12tEhpxG/nfHBO0qlgl/pYg0up587Hg0RsPCkMgYvXM
VCpHKRfQX7zeul37z8khmvlSoekxxg5JJzIM9sdiEevt6wl82HYN6CjVSFobD1obITVo2kXbtIic
CVt5vSPVjbGDFVBLFJxtrm0KJEVV/pd+UF/UlNdfSN/UU1HwnoqmTsSfFkXHU0Ltd0M+sesDukUB
egmiR+3JqTOn4eIp7O021EdZTv64CosJOYYQbrMx+ISXqIrOxh7Pqq7/DSxnpSHTvSKNyqq2+fr3
A/qJFKmqD7cogN0dYGMAktAhZxuEaxisp0vV/rBzD0suPA+GNDatDReRUexmaSKLTdLrjvIJXIdK
FKmTQ0BKwVGgGDWin6KY3FCc95+psJvpmjVFTu7aACP9qQp+PuxHYEmUxENRNyGb7Oj1QGIY4eM3
gjdvqoJewXJSBRWw0zz14LgHdfc4h0awPdnYkCSC4z3ImJgvuLbcRSnjktLfdF1kLPv43f6ivCLQ
A3jHP3Yr2ao4qaPbJozHR81VwCafhRceBDeUf2qSBS3rH0JjQ41qAzGEFP+bJ70Ocz39ho7nVAJm
E2FlnFpiPUSWJUoY6nOy+psZ4SJy8uvwGYUdJ+wv09uXMe6tv1EwVbxnxRy6Rx/GEIg0ev8ZR1Xe
SgEkg3vgikT1BPiD+VlHloFco9yDgfaYVos9KHmOEswTXy3BvnjScmiBpzeZMxdixsr9K/9UQIpc
9Qvm+jPei+9Ul1M+xo3H2qpLn3hQlegfjlf/ru4DEKghlwgo8ZPR1CbWXCtHTWAq2/sB7S+5nk49
iinDBP9G2GKQP/HZpudv5PZWOTITD3ex2TJ4h1IkJntTx0jmlf/CFPOnnt+3ENOY/0GlTwI3YXLC
gGAj8JOY5YlpKSfJAObSx9SussLc0R8RNOnf28IQgs+A+UOxLalwhP7E7KwaV2xPHTQoDAGVPM11
SLmWj2uatMsJgu3hv7DI0HjUMB8J7Ri2PETzJsQiACgPUBNiIOOXU5flX69U6QZaPm0yWcH4Qsb3
bZRnVx+cjoHwiRCrWMMDK46vuF4psucTkm8cz6qxSibqK8wKZRExNw81iXqCarYHMOQy4hKaVr16
UVPN2UWZe0S+cOqug2/PFzcjypir1u2HzdNylf/j0+tIXacRKFdB+XJD8elmqCsb98ljRBKgxTW/
B4WmAFswsEG4wGlIHm90da84B3tQBPpPysXFresJK7xt7LpDM46INOkShrZpkEbwUuQM7gBp8V+w
RMXOJ3WkrjyJW6MZkarH7L8NosS+EgiP/WgGKs2b01xB5tG6EGU2Qm1lI427EIc5cye1RNjdnWVW
yB2LKOZyV2IG/XEvmXXOWcyhCTXxucl+TKLPGVcwSHnTzTcTM37xnGw1CpH6q7LTgi0yOvBS18DN
fIiu85VrcLcIHKkE74OaVyLIg8sRk6H/hhScz+7RvyhO1d+SqKnluHSKY1zXVCLMyz8PFhjsJ2dc
F+qY13U1GOMMNxhUkxY56gHUTfrJiue2KmFAgWAR4BabwaFfKB1FAIC/krL1M8sEC+WU1cOjRnPc
BTyriNJenx+5XLlfpOyENwd/PpBJ4/leekLGxw3QZyTLmYBplQ5mZVDAZ7i2ac6sHyNlxGFzXUnU
TdB0KsYovWdDaaeVTSJxjTRcB5w26Ryw8KOwX8+ThY+IiHiEnhlWJsLd+ONDZnS92yOQ1CBeJlEG
aesdcwiODMaqwpdg/3BcaiQz5CIhwyKtVKd2lYzVrBn4qnv7vz2sUISqfJpIrss/aBPrYIfmqZ9d
V7nRlhDocvQ0dz8JiPLF/ZlRo1ILeusCsD5CTvgwLWNmSAg/uUCGDRA/eWysWK/RPkyW5NUmLl+c
hhN1IAXTTr6geOY0PDrjeNYkfqzK21g2WZyY0MH4KZtniTMnmd9sGyjSsqhDpJUnDkMzudzQgknd
UPiCACPTlfwWlKUzBk7eFKkMgsaio+JxyA0JEParg+tpmol0BWkLj2iWv2A6DCbiU11ahXwPg/lM
EHJ+VYy1iP9eSro/8POz45jR1n4fZtfwn+AW1Fb3/dplqe1y5Xr55IYwcaJyVB+s5Ntf7R8h9wuu
0FQ6MqXdion4nh5vFs1ChTt4Rnmd9G9RhSCc7IMrnSfpbASX59chg1L7wYSJhHh365j3+SRaVFIP
n+t4hw3pM+JqblyZj0lThHOSV0QF3ZWAmMyYpkxPfCNlYMMtKuMdJv8BjYgn9RfoHEwXuuUwH4ET
vkRQw9OKNJdpjYEJyBi5XP3fUkrVLPo/x9Xu2VfTkRPiQm/VFD0mn0ITB4lF9O+dV9+Rnk3uZ+Ej
nRO3IVHQUL24O4kdQSED7k7HdTmmfmQhvGvwv5CK+xSrhEAgqs/B6mIV3ksTB5SPhSIXgG9ZIxq0
HyxL/AvvBux9fzJdiYITtA8KW/pvohGFHEsp3y5QMFsVHWkT1vNfVnN/ol2YjSjw+8BPyosvpUSw
JxyuCcM0cTTloFKRWNXnzA2jhJTuqXHGqWYgCOrsD3IBytBx7ORW+UEL4aOepTvuITKmnflZdEJM
Q3RlxmWz8jr74vRE2J6uhCCPS42+5HSOXmAvysQmVB6N7UOnCXImF8PNHOIoXavXFYS1XfjeFjZD
8kAEJrk675GKV+4Lo7bCWFFL3JdE0jgMIWljiPOrA8Vlmdmpniy/R/jeaMU5MDWyPCEw8qvybU+z
8TWEFi6i5gJXDYlNHVRKBEVA0V17Pnl1uRLZtt3VqfQtO6T00RMpX79ObstYWvgsF4rJimlb0BiY
ZTnuECwE6z3ryt2nym47W81zugrku4CLXrXArTUyFq5hEIo01cjv0YPMR/cU70avZ3JuCo4iOqPb
5iKY8Xy5be/S/0HpNuX6LPlygx72CcK8X6jrVD5/PGn6xvf1QcvPuoyCYYGS17nYN0uEcBqQNM+w
c87zzHmosNc3vR+aSR2GacREquN/pvdSt+iZIFKzwbLBSVA/jgEo98gGEoFmLeGwl4xIbY+jWfLO
7bFaPCckuHo4839KqsASnMg3QeLPmMcSigA229ETWMjPEwVoL0fGDlEztz5sYkn6q45q1ttgQgLx
9hcX7KeDfSC6nBDfoE6I2UsGNqKGSN3m8spsRIpA4gh2VJD+nxsYIDrFDbSeFOdi2T64nUWS993V
HMAt9vASiItZ8JnZYU8Ulc/fIg9Iqu/lOBA3d4vkbERIrvr5FMVlYVD/CoHtLQTCTZwOZ4JEr07j
WCT4/4PJhrK061ps2MIQvg9Yc6+Wspbllftv/WihQ6bSEOL0AlXW1csC8BXIFQs7xqqqncHrY01I
Mwx9dP1Vv33h/51MfUweqaKUm6AF5IN1EOQjfagwS3w2aBAM0bY7KP/WbRNtrMwi2C0k4ChgkEY8
PR7U+Sz+dz6FN2dx1Pd0ymP4EWh06laNLiCZDrb0VMmxt8B97CXSqlRVYX0PS07+qSIkachMlqL+
2XjYyYgDJA/ABHOGsHVTYQw0YZPzuVfgnh5wbAXK68uV4u7XAEDYMY3Xb3iq0WxmV0etgMl3EpAR
7SJfy4XWXEV9xKc5K7BhlR2NAfChRWOojqiYPQH0nQT5Af0CoBcS4pDuWddarLgGOiThc68WK/De
NP2HahhQDtteqB+eqkLxE97RdIhWxdXMWWnQnD+lGZyn1JX6vxg740iKDr/LqR6TbjZf6BDqtEwh
B7e2GQO/gyu88wSewnSxodZ1+wbVO1WgroMHV9VCBO/V+8Shy6yrTfHH8D9RpY1J71ykWjI3IJmE
JunLx66Ikzuhrs0GTya/1DbxzxfviJOMTFvEvZoWlOlan/Y9RI9U8ITZRPElLRHksKt7kIC1hhXK
nptABIhAw55O1tEReT6LsLc4W1Qta9vKfSq7jB6hfmylYi2pNoCzMBQ3rJaP7aton8letRPTegVi
KOrmFOIQ5QoPndgMRFRhvXaB8R3QcFEekuTWdzJ5ESByn+BMrYkeeXP4iJX74jKT6rzdCSxgZ02j
VgafvilOobv4SfajH9KoNDxsmvpqh3c7P/gF305h6rbw1D2fWe09zxit6ixPklU6aI/vCk4Z/G5u
0WPGEUKpZ7R9345QBakJHjZSQ42qwboGqNpCvDVFX1wYN/ICY5U6f/ANxb+1JZintlu2LM5lh6N2
nbFMZM9KXjXTIlOb8t1LmcYuu8XfZezoKs3wL3sLxq1Mqh4tnq3syYYv5g17g36S2SxGqJ2OfcI3
ie2j0z/7uYc12WpyXbQn27ltPf25fblJweeneLapzvNhpycL6SSYjz7WnHGykkgQZLuKO6rRnS7H
Y99e//6litRNgomHu9Yihn7vvtnkUbfyN2/wdWCA204jlpeXUQsYtGHPiE5RSVH36SnPNU6/NvWR
UeoHgrXaBizV7pxvm3f6MYVb9Y4IQu5i3KEHYSbR2E/0l86sKZHDmCBNkrOz6JxCgr4o8eTWnyHC
2CqVpXJgnyBXgI+qjhu/ub30SuD9VG4UvhGgzM6jLs0wc44RHTEmLO3WheQeu0YQeEO+Ckxv+CjU
IKvNw6O8Tvu+lX7qAQaeBg+4y3JF+u337nqfXLywC9ivp4EpIyTVyYiSiLGQw/FoTfkfTieoBKYk
rqofmOyfCmIrTQOBqdNMvk14oemq2ThIRoSRT9JVL8WgR8TesUn2X7TgYTsEFbSUh/3nZ8invEUw
Wg4IqG7+USTp6dbJaqOyi4CdwtHKU3Yc9w1uhhQciecF9aU1X4wwH5EfJGJzQAcdJZN0SCH/ywjW
dA9BFu/lVXpkBNnVI0UxOtqEhkUbtdcSogh+jrZP7AonyWYLyaemDZR5ILvi1Fwfn+hM57HZcWkQ
TD3R0Ie//xz698nSymm9bSMFHF8KvGhVh70JVsQGD7VqLjdOE/rZleGoVxqehrS/kSUscQSrxIYM
+4cWz/I1gTq55O8PbN/J0g33C08SOu0piSfH9HzqQKhNyN/x2Li6fPJ/Rit9SXdHiShd0QepirHC
iRbux2tZS+RmoXp6E32IefEeq+up5XUWuw49a+75GBUMb57zDJq2D8MU17+44HFm6hx0QDYkg1Rq
VE7vU9AOadF0GftvTjF2i6goO9wMxVGoSNejcAQylEXfMYmPd3Bh7RUYHBdMeg5EyV79B8HY/FgS
jC6f+LLm+l6jFU5TfTwOYH8JhedpZw3LcBlrhaiD5tO1FMueVW3H0SCS1mvvP/eDkf1H3c6VLRT1
BqEYW7nNERBuiDvhx7o2KxvuSUrVXXkkg5BQ9BnMTrWRndCV1da7iEmmVp/6UN/f80DOj2pTJFUX
/utCADNcm09pomCSpcUu7Va2gF0vU9gfp8dIb9ZktDUSPUrLs0yNvW4AEBBfPIKe8m9OE6Xm8q5f
yZ7nRHopuxsCiLSbehWz+pbxnxJZgZVzEKFPUCd92NzgSA2YCtB5/HKY2juW1SACKO76tYKOW9Vy
010IyxsoacbOBeBsJxcB8vLwtNQO+ZsoE6BTSnTSuPbzun9uMbvtN53377y0HOrcXt+/Bh3L5sSF
d5OQH4R8jtR0C5jv1R6EBZ6YAZNeMfUgtu+G0uTAPySaiwfxMzWYsvPEpKOEgaBjFMelq8huH6v3
QNit3Il6V+z1kOmFOIHkPJyvm8hdtbHbpTOTgG8A00aFJxaZm1P/T6bem//XC3RaYNnslg5vcdQV
IVCiIHXqtGGJOe5zKvk9GBDL6mZEMv1j7bKyzedwQqAcztbC1iI5gghbODvdwUYYfm7VrhtT/O+E
phM46pOQ/4ig8L5XlYVlbJf+lXTLVPxLLWISpsD5KpoJvyEv/BLSOaawRwkHYO/nB6AYNA1ZTpEX
rKNeFB6MbRhJ12rQ7eVrQXy8IsRX+ha/sTrx4YpnRlUSPzSEJ600QPCKQITZGnsi1gw4jaI7ORHE
RTQ9PmUt3BEaEKCrsCG0CqjXNRVy45Qh8QejbYTll3FqDfbE7L/wCbPYtZr1TpH+meVUqzT//vSv
la6Ai3WZrHqmXH38BBnynOwecNOYLjMD4W5VINHsbIwUNOBpR+xke3ixjl3NDQlS+HpeTE2XFJ1m
16zYAXd5WHI8mg/jHHE081LbJx5uWjl/GUpQG90t/mH4n6Xx7WI+evvZeBZH+FXAm+Wc8sa2eul9
xI+xhxFUw097SMtShglEj2tS1YMPkjpWBRLOJkFdrhrS67yF+wF5leOV+yLe/Nw7Nxf13gJjhZn9
ZCOYlUAT30wu0DBKiogMVvbD90EINQRD6IgaXqnygfGXA8SUipHILORu/PyZRQxrKH2bgm/s+gSC
FM6LMj+QYxdvT2Gnk6SQWWczUF0YRmm/yh8sOq399WHjr4Sfd9lnKuIxGBcw58hg9UxMi7XV9YzC
hhZ/FScaWBJt6MczYGRMDa8MyuDNYArSvckoMAkf1/9Qhzebx4Fb2nLHdAKoFLmrVSHq5h5JYgXZ
YmrkD8tzuTJZY5JmUbYkF7i68RWCCdSOWMqdFb0LiITIOTpVNkWAgwO5k+ys4PvBdY8YxMXc6Jny
egryBaA66hqsm/FD9q/J+trwIKui6Ls0mJx3jcrT4n45yf9jMoccmPG0GajTbwbcLdv6fs5KXFGl
ilmPzzQ1LIjvCMsmvQj1TW0JS58lioKWjnH43gqN5974VI9lQ112NCzFiycNlua+zK5qCa3Ri+05
N8XJC98z2YHBV4DzLfbcBZV9Mur6P8Y56F83gVh9qdW3cWu0q8HX8qmXrLPlZFKec6NdAbaeDQ2q
eA75LgIguDVP5fs2X17hU9H7PlXgSWHbo1bTEsJt/yHv7BTTT71RvcY7HoZJcx7hzP4S6W69gMP6
5Jit3eza/dGUFktGHgnSfRy3JEtdQpV8xUZI8WA7ALkkTmZkLYjbSSyaAIQWJtJcDOsJYwDgJwFF
dmB6c1+rq+8mC5D1aYkXfxSbhr7QmDfqz1LI74nQT0SqQiKB5P8831SIrfLILOopfvsD8d7aIwl+
2fhNtN9m//UbDBXNsX0hGQACsWsWJ0GbgG/IsLcI0P7M9z4ibtGIhdcn4MOeycrUpIDTeeVtfv3a
LKb5JdpYQKtLgpWBd01IJbH/JvfV49ZiNaX2SfGaZAG5lpIttSJLYaVpkh7OcmViLQm3MoiYDfyO
nErzd7qWZ9xIPE5db2q0p4ZVkE7BMtmvB2l0cjgH7vR/jSlPrORKq8vJUB97SXy7QZocXv/aNsRz
baO9CEqTxBUzp3qYlpHoLXjSZZbJax6DntFzthMLo91zNLHNHo0v++2I11WnKHb3GZXA1Jkk3m6o
4pLS5rwXIlKtH7T+7yIstcH6WfDbvHSSutaqesXeGy6vHG81EZnXotKpGU8X0POO2IXOBRnGEQTR
r3XTT1QAAVOgmtMpSnvWXmH+/SOys+aOnuYgip2/YVgId5nvR/ONZO4+kZt/nPPOnPF09Q+VGOLo
qH7SGcMD6VDr3Z78UZSVVslazNK8aTAZlNPpP5VfA8NHMezqwm5PIJ5GgeR8wzxUQhAvATKf6kqQ
urOJo2ftVxTkF7D9/j59XyGQ9NkUKLsGdnNRiTc72X+3ufcXFJOEdvvnDa3HE4w/Qzm5+SR0wxqE
uM9+fYHl5ISJvMvI7b2rKy3MKlPpUBXL/dxMGoEgHfkkW6efHvbjysf7BfJSBbXMGrpLbjkIJ1ac
EcihOi3Eky+XWwobB0e5egL8IipB/lHwNODm3FBcLDVj+aW9mWxbCAH19w53NQR5k/OUaeBgcPeg
wiiN5Y+kQ+2G7E8uPALr75A5Krf7ht741GYg6BHhJCZ9GHVoosNMZFacLppGcOElzIpgfbrBbgPK
dFsaEdtFsLdZcDVN/xDg1aAFcuzo33098hLPVjXJCZNGLe5crUd/qg+MVgbxK41u4i5jv99POcg4
39rpUBB1B/fZrvTFqYEXOd+MrzdI5aSZ8cQ67dsbfyFfSIwLutO9EfLQI5KIaDnwFzVOT5iYdadk
dvOOHIn2K7JPi9+AKeenP6bjz9lEA+/NgcF68jOECTbw22zDrYn4y4tSZhCAIS61+tM55QrdAF7d
skIDnovQmdaxPpVNbpNrJYhXGvtzOb/WnSZQNjEz5BN8JU7+Y44XO/ukUhF8xdrM7V5BHQ4J3uHZ
EO2IIiO/oSMtbtF+TEUd5M4rspifjOcbfasRE4+fJHdl9ixgx6RTGhLjvQFRpKEcCH082ahbGzLG
lqjnF1BjG5ApaElseSUtvimxkPEmRhz08jXnRE0AHMV8V0TB40KtpwptI9pKClEFx4i1AIK4CjuH
RNbzm+wQDLj51FU7P4DnfWq+RLiHBnzFZ8uj7A2wFBxCa+yZkHA9IOK0tem6mFKUGTwCE90+b4NQ
xl3ekF51QdR1Oi8d3ogQSBjxs4FUddXSQ4Sioiyw6SbAR6g4QseqHRpPiayw1F2bhiU+B2gDvAk6
PRn8dkBj1qBOB0RQNUlo5ZPA/OvGbzTqCrxIdhUR74mZoPJn+Jfz4+DpfWTRFHV7SpsPXozzm13G
7siu+aP6uubnpUQGwuIl3nSvQvpsjP3z0zXmVjGi1OCeI8ORRYjtltkFE8I2TFAwlz477afyJoDj
rah/Mku8hwrTZZFhk06oipny3Nrlp9FhfALfq4e2rChI6EfGtCLExCVmsI4K0wHEaR7ZQ0bTbrpN
jNThkGXHMYSDkzNg4dIBofBLZBcnZ+3dvvOZ8A7Swn+nBFAaIjZHZQ6rk5iLmQIR7kc1qY7D92qs
/EY/fVXSOPggBcGkHdYg/kWuggFAUkG4hNYRCFVz9JBalWj6nbhVeJbjBSsqa/P9Qx+ufKe4dXnL
3zpKPdsPJSF0PW/u3vKKN2fjodjTf7Vf9rzufaZDTIPwoMHVI5bZx1TsgKVEF1YuLcpf6m30AQQN
MCmAyIqboDI2O95/ll+EJvxUnWNnXVCOzalsPmcnGY/75HEvoy8lfSNTPfV6bNIpjUql1P0um+Zd
Nze+ZAB+1sYImuikqAFuVNqlvQ54mYhE6Y2gL1BOR/HNSkTorbV6VWgqvZv9twaOe+iakQN+IKQd
l5N9wRzOs2HhUhGtsXJENtP+BXBHpAi3r5+Wtq13jdc5zaNWSGNNdjVrzCiRnledYVglLn75XWhc
LH7S8ywvn8Vi8VRVbBcEoOZl8bN/GZ0uNurKvZv3/VNsM6G1d8gdXihziA9pmCjhxJ8Ffm2WSu6y
NNJkOFSvIUk7CQcfuzZ6nvgJrZnDSiKaazl0vm9f+4r/VNCv7axuwn51RBwOpr/VUPjlYcO6i7Uy
3Ew9qWclQpzNjLt7Asfk8J0171zI6/1dwQ7KlmNOXqTA5sS+Gt0SXmZmxIvWSpAwB6ScXViENuN7
8lnfcMqL52gGrFFVpdHUaKEgCrpjQtf8LYMYsbwscXZVV8CaF6i9EytlfDkQiMLS6nZLjE+bajrp
dm5x7UqjgFikjSy0i61W6FDYYn9R8NV1tRb5bEX0XZsmhHaea/S6ewXfD/ZZlkkUCUf+0R6Zo1y0
dXHcOgKSPrJzhslMZKevwOiJGa1Rqs7qEC4WsDWVA7f1ZynRu/mt2Uo5oqGg0ebmx6wXp3hWqgQw
BbzCNLmFbHKTTYTLXJgA2gnYuj5FRyhxQq8BCIX3M5b5om9mlcID7WPlrpJTcjbtprZIHW5tknVq
laGT9upiAJLENuRvLV7yJQ9pHnwfbLP+7QQgDFVzWZ7zdMmO/IoK01o5+gZ11kiNhuOYXYTzbpWm
EFDs86GAws0zNoIi0wf33Jrw8axpUztGKE/mE40i/BwNFFJdRdFpygy7pRgOPWG13nh6CpE7AtCT
zMUNR9hB9R88F/4pUdsXuFKN+dZwCeGD6HZvjR0+Kddh4VnVT1dxizDTZEyOC42MLRgtiAx3OFhp
Z/P6jSciw0q49jH9i0g3uFFQArIiJJnKfql3gf7+roo8iX2eXTyKKFNb484gku4peF3rQ61YcwTX
LKrGC9y8blw99NcYu4Bi7KYgscl4DrlPq4lRM+RMPyIfGZLosBI4SwDkD/AtZMsWhNeGEiH3tBd0
M5FE9f1p927oZmUL/Z0U/9LQTV/XZW8Ig9+jmX4lY9Sw2rxpvqQE5eNGbx18gVz6UzCsUJml/ttF
IN6SkKy8l0g+Ebtwct0tTKVnurkhAj2M5AQl7X9kKpw28sxPm917TU1LtMLYHu6K7W3RtF+oBHAN
mkJ1vBWBtzSLkmCFZ71ePT5WeRv7YjAHDEkvtjU4EJCBk2AE4HrA819GrB2Zd0DfD9DpV3RljWXj
I0eHxpdqkCJlxo2LCAptptbKBzPspDucAPLua+XoTIohRRrna2BkyMhumGZhZTBXTtmEglIAmcJ0
j70BM7C4+Sjtad/4xKTqVgt9n0E0gIndy+j7V6G/47uFiG2SxiPiZYQqqUIMsUJZERJox6lskC0r
SnIbhYgXgmY9EW/WU4Us/OsDD/vZFxxpxeN+eOnelE7QOwBo6Wb1fBt6cSLOcsvLxcITibITtjoQ
/loqF22C8ZZLFpc456H1jdVTuql80kYbYYLyc25yR/kbyzijx4wYCuYS/dpylSPkv6Re7ZevhZ6u
wg1aZxxa5gLSHdAe08EWBbJcO81mCgvt87DwnwcMvBzvYctoVZIb+ANG+NAYWOlHvQGR+cZ1BRPV
UhZU3+JWG7xpkBsixvBrH5KUx0X2zK6lgzBZUYUZkyJX/uqFLB2vZOU48el3mu0NTUKb7JZ9wKoH
zTeTqSy7vX0E/wcFxb10wXjzyk5he1jkDuh2nHp1WQ92EMDxlA7pHP7LxfQGpHm70lkxrStIILzc
iqTUQv9RwXVEzlboxpTmxKmiDcpH3gcns9F2OaBqzcy/yBjgZur+BiAbMcZL2jPjSJb9aP3v0FcW
JC7rUWj0UDfolsmxnsOL9nea0GJx2HupLRLFx4htICHqhYiM1EbPczBskTbcNsrQYHHwfkxqmdtE
E6Rm0MAL1w2vHBjeT44IjBWvq8hkYCfiSGSzFFwhFAXbzZUD8KxvaXtFmXJXhmejTvaD2+MsB9hM
o3Td1q351hEYWYdD7i8Ud/2FsQCNgfZkGWoUX2K1V0Sm5YVVyeUoZYBwR2Ip1pFBGo8zI1DiVifm
rOv68XFd0bc4GIHnreCmt4GVPgBGIqHGRXs8w5TjELthc0MqXd64LOZFRtAyydPSYNkdwG6dtZeh
kmOVBV1jQXk1AsC2CIYxuaRsbVqms+hZMCKBInhoJKz6vVaG6drsQpAG907xLX2/rHxBmFyy/F19
VWdJugW2VxJglZaMKpRUPfIYJekePLbVitBRRhF+uC42I2Ij2Kbd8ECyqQMrfaXh3blISviVqNXp
3oGnUMppSz0/M5MD6837/4W6oCK/8uBsK4kG2R+HBKfn3RXYreYEd4rrqeDoQzLUPhCbU/IOZi0s
e2q1UZE/7Bm+YM+ugMY+OOmYvNinUhk+iX8+RvFL5ACkPZ8hcgiI7nSxnTo+MLawHDK09oUVf3s3
kQOXIq5G8to4W3D9Yf103Y/hq3VIhKi4F7abcAM6Pux4vgrn+QaAYmfh6Ak3riUTtZ0fkiNzmLq3
P8j92QbS6o69+77HXYqgp/owzLJh47+lmSeceesv9J46JV7HEEnwVNMyEgtju8VmsmBZXhTMKGZI
je8hJhc1MEKrhnYGqRyGzl5PCp+ld4WwXloPfUh1RfdSna/N5M0yiUxyIfcSH6BToSpqGkHzQO/A
P1IUfRTFsyS+3WZzNxv77zfn6YCkY9UqZEnenGJzmrwLGzqjHtTjwqfBKuJizXiynIDYd3hnWWJ3
kSvZczy8xJa8vU5UDlAgmyyu3jF16cEmkZkFrHn7unryNWMH6S8oEDmJDCG4RBH2Xx1bQnQMsrmk
CUH02TdpCFIlDxEZ0sKcOUxoNuBJ6SQMIFd/09Z9hEBV+0nGqMYYZAY18bR8QB5lMRED9hTvcVXI
gIfymieadKcgG7EzaxbEP0BTdbd1W3p1AjFp9ojadDqHLk6854FkhVdabY/F5+Or6zZQx0bXuigg
veKW1q7vYazqxwVYT9dsb12tIFCqfQL+r8eJwI3rpHrHzoSW01VFcUWzQfsaxDSnp4RN8BdK+M0R
iXHJ/oRu1YvRXGOzNSyyfmVyFyKAMz14CtELtZJ951AL1XGkYC/lireNFMTDmsYXD38uCmnJiRV5
fbQyC7YVDgDINtIFR3j4ppOUrx7+cALchVjGjDjJIwYuqxNtk1SffD9I7b9jbrTMBED06L47Dexo
TQFP2Vz4o7Lel4HDJHThUZzwVcB4c9VUJoj5oTxqi7BuiA0KrLpnqz6wpXESGam0Rd5m0yzJwIuT
2l42nYCg7BA0zc+I8tIdjAE7cHwV5NmbOMkoQhy2EWpbedDAZnjRr4bfPEoEuxrilC9d8EMIhnTC
f6/V4WW3RQyZVl+ta9xbNR70PnS30dQPWLDxBeojHAyIQ1I2aOTe3oPQor/0l5j6DY28QiKweyit
QmOihTPF+Lmeo3vuPraBl93laGzm9htmeoD8fqOnXxd9SN7kjavj2mRntowwVhdLOjR3s8RLNHWN
LMyRA5zwUSgouD6uMytYBZyAXE6mwlPYX1KWQhWOCCer82Y0TPmGZ8BhI2g/tLgYehAbe85YA5MS
ngx6ebyWiap8CdZB59Sab7OYAhYQcZVIYS+qj4oWTVHWHOFX48yRv0fkgheSRHMs6mqAtpC81qMA
s/NwxvdnTxCmScm9RrEEyONJmCu6VGbZFpd4e9QZaFxQmYy7SuZj5QDhhV4Fv4xf5CxwXflweExj
/r+n70Io3+KMJoaH1ypbcKTNY2eHUXcv9gv0Ee1WMKZk6O1JgODnJX8X0ScPWQAknFeYiz0pjIml
MLlAWgtksGEzMVkqyw3a36/8fmm8c99bXit/tMcnl49zJZRQt9VruFfIvmCJkNqZPBpdJ5JlR7X9
FEZByj9QU2fBRHEOiTjzVt1TP/e9zMon2rTEvuUqBrRIijNSdiBai0uKkms5304wY0YiSNfS6T6T
cQJopMm5rkZZqAJ4k4zmGpjS2E9Dque3H21OtilZ7Wex4ZDy+imKZFX9tktwPhB7xiUsIz3xeDyA
gZzhfKJUKRWUw2rpQLClnp04BdonmWLCQ0ZlBRxmBbzBrBsIXhT7uxjYciTUtg8dO7Xz3J2ILT+P
gWil0VyA4MIeQz5uObun/dM3KGQ8dbXGrj45CQYQU5499ZJhunjU+bYVDXE4kHWHADfSr9+g8Iu9
aYNBFvbEykj2FfH3fvBmENC4fDgFYmMeoKNTBmsFcKNN19n3eJtJA1usAlbHHNzi2UTPFp70RYv9
90n1xQa27y9iiITNHhKaRbK0onMAOd0I+ySyDAipYwy7KKBa+4n4CB9iWmBwr8SiGuLtrIIoBiNk
vG/c1hmXYftbL4wWnN7XnJD9KyzIJ2pyLTS4dg4c9K87pbfBEy8yPg2vRjgQOISkm325AQI1at8g
DxJVoOteE85gFpMpduul5+xrVq5+DVFgpCIFwfEsCkBsUuprR6H5RQ1SAyJY7uLrD3pMl4mXN3rJ
4+UMUgWGjcfIvBZre7tvviB9zMqvUESZicGh+jk3YtA2D1VmiOeBjWQOxhufMRVo1qno2zjo+GZ9
hPM1PcJsPHJ7FCRr/H4vK8t643acdhGTXOzSXsdYhzBvKcCtADAfG5kiN2q6zNrs/qfCbyyYx6m3
wyhuLB01cElgcfX/0GoHTwELh2iCzhH9EcbvWizRz88ZlDxZnvtG2sG8w2IcGTPd+Ac47njFaxrQ
OMSmm1fZGAwxQuHFrs2Qvg75HH67TPCgbvXftGIVGR8jjVrFp32NIusqy7cTQpARj0YDS13TAWzu
iKIm429bGZ5V8F04WNqKC8yZNpzHcOjxL8nTo1qlr72cqffTFz0dWCLU5cy0lYLxf4B8x5Nbol7Y
grT56wMvXm0tRzHgbcVddmnLPq/NRppuR1/d2tbx9SOQGQ9R607gmsecUOe8tBx8zGWAR3CTrjjo
6q4Z3HL8jNy9G19LCDWqk/hF3qiHnm1Xhc4zml0dtam/7o6CEgnGfPku7c4lvtAL6/QLWj7IAZdy
m0AgP6Hc89VsQkBg4E3UJ3peUjDjPbC4PiDO7aNQhC+qo3GXZY5kyqg2jsn5NXhRa9tAWUXG52TA
loF0BMb6nKkPmMa6H69eLLD67dMO9+V+BM2sP4fzLeCIJcIQFt+8BTIBLjkyvOPKj/NVukVLmlsC
H2O4JhWy+a+4AIJjWCNS6Qhc9Ll/E0A23FA35iTgX/Bf2WTeHukYiygqfW2Tg7ct36h5kV4vqitL
rOU7t+whOlw5JEhSVKGObn9nOniLIkxvtrz5K1xEKqrUSQ5MB3/rASiWdyT6z+IZfOl3TUGRE8cv
8hY+SYzifg/GfwiVBNyY4LBcXeRS1X3qK3KxecmPxYZrFiw1VCMHvj7NvkfeBM3C90m7O8k8oXoq
tWXybK481XwVTOEBYtzpr4aSZEkt/ZbU8iS/DUEhGW1MqSZFFXK2aZcrj2O+kkBzbfk0jfo1Wdo6
kTplOp12uxeSRktCitWHlMWEpU6j13QF+S/yR6UF4Cu56uvauKvUbzlKqgur4Yot39pwwh99yr5B
8jnnKtOsWmvnS1QIz4MXvZNLPOfYoVZDKDd60QRWcJZa/0b8MuAY6Th3IIj2DA8tgMsNm3Hr+QT/
3sy+nEBC8/AvKSmD4HO1AGYwA3PBLIT9PcHTk47BLKCC1gulcuFKEKiRiq5r0H6x+artDpmZLjdY
ZxwJIejV7OXSfczD8l1wVSBFzi4H0Ls0KCy/ty4vmRQIeX02OA4InRFmoE9hfQvFXzt9+w/8sxYl
B+gCNn4J8WQR3SwIuZQPHUvAKEY0X1hJNECJ5cq1AsiUTthMExHozybZJcHyD8F604Q23y75/PvS
+enALlYsiMGM+V2FTyMxwbU9pApd2lNkyOCZSbw9qEQ9qUT/kd2ahbUN375F5ZVap5fJWmqcQzxW
qL+1I2c7tM5XC+ZYzHK/3TsA+3yk96hqYbahpvYJAiZVpI0kmjJHSUsTYBIARiK06CuSA+yz0v6p
gfmOCDooRmx/V9xsYFJAHXkSc3+gyn2v2aO47MvndVsMU9MJ90qQFSMuicVnBCXt+R+GOS+o9lub
cCqk4+aP2L4hGgSEsBBynAc2Tp21bSTsbp/CeypyDVPAExZYbGFoY29MQopjTwpSYu7WZZN1XyMY
UQM2OyQkungvWOSA7vpYNaf8od81dLaG91Gpg8sDgm/VpqlyEPMUGsRgvi5wD6hWfWoVx8WvvBG6
+iLaEb7QiShHeEbvor3zehigQlKSYAKLRFM4TtBfPULbjD7dyOj6R6SuQEtTZSiowoM7eh92hAAf
hocF67VTDaS9bVls1WFT5/0iearVvHrpcTSijSzf36Eqb3X0XT0Es0qORGmdkxX8kCUtNGfgvwqo
LHu8U6QG1TCVlg72DvVrpoEgqnaVPH9RZdRvqXodUYN59cA9dxX8hGOxCMEYeJJ+damCOyDzywO2
hTZJamIiRfSps/2CgFBUe7vjRQ0EyERUyFAwzo4uiZ3M525TVZn9akF0kL6J9EAUc5nN02q00Hi3
KsGJlmfTezjS+OzezQEDwUsQdllqDONBhHJDfyOwDkM2gzjuhpgVURuFXTolHAX5JBkW/elQ+5Zk
n5aS5oy+H/xNhIWJ2JURbQ4fdiB3pLK1ErvjSZoVp71aJeiq/ZF8H5EaM54T/0aZkXcuqECAY4QH
DKuLcWIEYTZZJFVLpIHZmA3WMEhqFv1Y4v54lto2Nb0HbX/wAYpVgw1JtOkD1/ocOETvTUCHR6E2
8zBoTR5FRZIzAyd6yhAxSUN07EUhT3GfE1PmNAsApXNKFALIOU8CLRZATL1KFGdvM+kXMlJH31zo
jrWs1+8k0isE4eM0EP8EIdh3FpMzTBDvmz2U878ItmRr8hW80yf4hdcH+VWRYlDhMPZe6Lh2x/N/
5K8wmcje9zeJNfX0zugziVV61BbAaPXjZo6FwIeWz56jQePeUdiDjSzRZRXr7hrRLD+eXg1zTut5
yqx/D5Rm5swHdXXTbfajhnzzPJE/8LKcXfH5STme908WH3Xip+PJsSQcZwIuSe0Ng0tpKHq8tbia
oeQ2e3cGvtYMlLGkRrTCvbAqQ/nDq83Lwe0bX5vT0M/i/p4HkwDlfLvhh1GhLEPcqqsD9HG1mwO6
DPjt4XifRH7YQY2rbKC2J0iXNeorlrXT7LhsizOk64ccfIMpAxiTMtHPMr9D1BFeEDvZpIB2IG8V
E7b1MbcSNYWvKgq2QFDYCGeiG+0CAtxXUs0fH2o6Z9lOdOnFynckGxCRcakZlFPNWJ9NH8C1ykhf
axYL8Oe+WojsVRL++ubAUT0AjROHOMnsmgdOFhIsQy7gvzbZi3tczNyjP3zVQIezocjnUDf3aj6m
riaxniwleXyBEzRspxWHOBguZSMJmCkYyoel73Mkk0csbQswLYhTcvodMi92cyxfhbEwKOLp9j2x
gx0tYf6W3g6sVd5BDkuF/EhcUUpmleMUn7O719hYrpsKurMaO43fsdz24PXX9dazihhuFOv4IOal
9K+FxUr7vnJwd+Y1byOzfYb7r+JLDwXmMsCg7YBj1dIFbKNN34u+wOH/NWjNFa1huZE7B6MMmXto
pBvKCsSDjXcnoF14pESLgJs2CCCUeyigOGshw6k5IbS5i4h+2eTXuKaFuKu1zxVUdYLjRpqnHd5z
+CQ3HCjojcX4ivPdsufdrRA4ED66U9HlFGz0rAG0U5ABt7tjZpgnOG+qYHWyMw2b2MTyx2AsBczD
nwswjZ7hLxK+jyhYQNnaqHY8X+sBCFx/chERelKZBZ23Jm6ck8/S865buhBIWJNxdvsqjeV42QQx
3DWgXYrVyWEzqntS4+UubjlqQMcbEPCpAenFIiJD+aYLu8zua9bn7ijM5j3kW0cAG3o0lzx9ANSL
sYdeUVvF1Fk3H+t3AiKfcfjXGW+hPWHwrBgPeCIP0Cf7zBcoJDTMm+XfhqVpX3UV2lBOl2bg1rtn
trRzBjFuewdMFItlQjIyV6Q4uOHMYyG4zfOaBKEnFLWoTotKxtHkLQRRbWk+Q9nySDWi3w+Yo6oq
upokSRILsvzK9ntFrE88LQHV3oclrTe5aYObyWxjPIGQFQ6lxXOcuVBQ7W1r/0DXsEkjmB8sOJ4k
BD+unUdGGzTKf1mM7mToLmN6PZiiFp/XNaFo677zhHap3Ns0CDywtfOqcCPusQVZ42BII/Jj0Hnw
VMjPnaofBL9kIvHWAl+2WVRchXxd4Iq0LW+mQulHs9+WXrH5plbAuiprOawiKnfHm2t6kt8X6yq5
avHvOnmNKbwJZpmw24Hk4ODgDaVexfm3GPxj4dCfdJvwa+DKqfDcTovJECAjHDIoIZRwvI4eVvt8
JkhH+OxESo/7kR3I15dZuZfiFdJVbNmbci7SPtOzFWbRHG5Hv5xNcGu7ksI1LCvbaLmF2hffD3hx
JQw719347sCEhuM9xtkE75g9gA8a+fLXHm5Nh4T8ufFwE/QqXBzHrIC8RV61H+RCFsAp8jwun7nc
vfgpcVqP7/ORxIXoU2yaSNfC/zo+48OJTZ6lhv9NLZsvG1mTF/TGUJUZLtrQYkvxMmUYAi7knYxF
KtnM6X40jRJue/ryztBamZx0NtUVcCBLa77et3lFhMKvbAHfnYC22qksE0+o9sYNPR+laDhSoj4r
ZsgqNnuFhE4gAAtz7amkEJDe6RlVvkFidzKa7Rz1tbgMNg3JjsnogJfOVii8ob+1SZw2oHY8rJs/
Hkh1vcEcMH51Z0eu9hfEg0r0wdZgrqJMfKzEovDal4UkuHfR0Ao7GuK2JIzCqRu+zjWisBtWqVkI
4kyxpB1yksdLYPBbFbFOVX9RAJG5jOD02C9J5PhnWrqDPPWWP9LZNg2l4JlWijgVbRR2O8+1Tjik
MBXOD07uQx7eeIt3qBea/n9QTkpbMFbi738No55nRbNQkt1itb1tU+B21wWKbRAXjAtQB7ardykc
3+9+yt/qY+4aNIaSrNEqPICJiXm3WMp/dpJ1kiMAdFiyid0FvzZ0TrndX68gtjrCxy7Qj3yNCSnt
cD/nG+LKQow4xe/P2DoefS/wY+cZuevwukfvF9MxLrA1OW50o/JrrY3R3fGlaeeNWk+kQcn8ZE77
33WGrD32bCEHhXQ/6dP0Ojp8thFGm0I/rVKSAgMIqfbkytcv/XErZd8Z+wSo1Kt2c5z4OOkjFPGs
31E7MQ52k2ab6R6Rfy896OQMmDSCuOubtdg4wIDJ72biJBPogJgkLXDIZ+QC2IJrVb3YApsA+iP4
61Y5VSrt7trjIfsyejzJ/plyUSCRnUdUH/04hDoGrXwpIrk6w/74YGmCloo2JYqXUSzKUXoyrxwk
qYxnQCnW96qLLuFK9Eg1Uk/pEX+ye/FS4Gxe1CUNY94TtQfCFxhqLa4nrzynyuxEaz0sbkmF14ZG
d3/DwStSHW8HOyutcFgP3dxMDkqyWYj1eaEc6YLT3rCzf6EHVVGFDpvyp6IVKyorZy24X+rhbj7Q
BNM1AEkH+9UWDVdKrOCQ9W0WC+85TxOjugPuw4cOTV4IF9Jmk3NLWmav+JQxBjfou5AQTN/NlLpE
lzpGBI2h/NrB7GQSFkSyZxeQ20CtoHtKjuLibhDIVcBcv2vj5tkk4pkrnkYXMuN8ia6OWBfq97I7
EeU16iysD7T7Oq6tmqg8Bbf3at/2+vzNrnULS+MIQZpoEtIIhr/ENQzB6cyM5XvHgW6eQUWQovRu
vd7+i8Gqm2R8MQon2FJ4/1hwgZDgvGtTVRgNnXLEQ1ovQsPetDWulLEvZBcgzU16fambUW1aOe1Q
N6T+qKAd4BrkY3A8393nc3Alw3it/n4TxXyNoV7DmuwG4kU8fDMMGYKI5z7rAH92g60s8QqQl9EE
hDAKeBh7PZda+NwmRj18vJVbKwSGUwjNur6rSgiB9TOpl1pwqdNv4aW8FwY207saYU3+42s/Mwno
U4lxHqPYQVPELP5OnvCi1BoARsNEyqzNQfScwlzcYwPjXwNGgchaYEOsAKPbkkEIJVY2sbHp2aRO
9cNUQw1n1917sWKiimpD1aS24BCfyCxFvhWAZDYGlh/YfSTSDRJ1dC+ig943gPD6slEVVynL/z93
snw4xjQ14p62Pvyofs3AgjwRsjF2y2fGqTKfebEuYfgwuy8skn8HM/IEZ/i5uPYVKGAlxOSVRbjQ
MBUQi69C0U/CqvdWjG1zWiXAmaBA8DKFAsEXmG2wi1SGOcX5qPtVf1vq4e5lFCIGQX9ydFPdnLjz
H7yViFjMvs9UIrTibJKIRH+n6HKbjrnugpnOjieRG3Kcu8vl+VQtew3R9ucpTbyCnE88z2S75bve
adjfr/w/FfEJdfvjJR4C6P/OWvm3O9uc6CE/JysL/4ZA2+OLofZXPcM9g+h4Q3AEMTEdG/xcOULn
47J8mTrtHSztyUEJ7P/00guCT+xdsamzkX/nVT0bKv2k0XaF4uQOAcfslEaDj4HUxA/pXtopH8Fr
fBQoUJS9QgHuCfwOAcEY9FjoeunQqAReLoqgpDQB7O2+v2axgNCo4xXFBsgeIanSzq+7kDbbeC4q
egc3qA89h8DXwLjFoI2PTMu2AqKVPpRMmsXxLKEWV9joDIyxgJXYZNZvdpUbkejVNvKAIgh43vvK
vEgkaennQJy0m3Qj5OAPRDdYE0RukSDlJ6BDjrcIKlpxbY6W64370PeaZpUoV5VW5Chtrk7UPNLF
E0fT47isyz9IYvXD1SgkKD/+1CsdnLqkg367jkIhTimoDCj7JOVgicYfyo+qJCrSiJHtOz+idLJV
SwylYk07Sq2LAu55dWf3H2Uj1GTHUkNmT8JoCHhv5QNL5pJJwdNHi9Bj2ZXVAhb7BcpiP8k+4//6
mTI3tIMi42uDktnGMOTv3H2+i/hmcqJSurM2MGwmomCh0scISZxf5u3qZxVRcko58VENzNR0ahtK
uDmvLKChTCRSp3NnbhSJEMOXXoND1bVkW7fC17D51Yegv5qSEDaZYPtBKKyrnFV9X6ntCLeUlBnY
GpHmqs5kqVRzufxavXBFl72lRFx3Np+IgBRWxXArjSO5bYdgw/rhK3sdDZ+uwL6NEyGeWpJGmZDo
L/o1/Bfs7ndy8EieXg7GJF4nGCNfE0rEFkQ6uxR0PFyqbcgXgIX9CTcYyhgjuNYGfx42BD5JHeSC
j/jDh0DNvLbswaA9sSIrPgJVZPYYZWfH59Lvy+Jq/28HUv1cgngkYCbsG/3C0qlSKG+Ge2urYQq4
Gn7SPwHrMauySPurYQVXx9cWdvIY9mgHvpBkOsYfXqV2jOsFF9wgMTRImHBKdwbGwuW4UWLnhkMA
HYfsMPXW5y2+wnbXEb3k6nmiJNkCV61cqpNWVZ/4oS4EN74lH2fZ4at+uOTNOHldGnTzym6xmwKO
yDN7E80FA+i8kYiwR6LnGfBhO7qYqzPPmwwWG6McJoJbmv1uyw/Vwa5hKRGI9PXxD8VGkFi9TpDj
IUsCTbt+ziDvn972qjJUrXNK+EvUEvkUOzb6KxiZDonVb357LJBCevdsW1maU/po8HDkQ7jnbLZ3
XJb6SeAmwHUmZVTksfmz+6YJ86uNjADERA61+6qVQBfSEDbnMRUuUOuQBY4BHMbr2iRSM4+GvJ2y
GfM1jcoq2BcFIvXwUG/pXAnMTluggJgQP6bLnIV3b23k1B85qmiPmaoDURFjvapyiAP3Zw2J/6zN
e7XpvA2E+gSlVOwnmGifXbko2Ln7WjtkVtMM8bzfP//nYweno0c93V9fNLTLM27FHEX2DYEo7142
ac4TnL5WXPsAuRBY6fSRspeJK4A7/Uo2dcqEo9Rh6NIQeKhIdIRnxbyDdAXFnf6ARelv04vFWitd
z0haZKbV/djYoiPkmkRmRB0xDAfi2JJ/aRPYnK8ZVQ/OTf/AW1zNErsmzF+K717CaqRW4MWPHHxb
vscZtzQwL1aBSgnrAaRlBfhg+jMlGOO+CcG2rr7N35p7FYzBI0ZJfO2cqW6F3Oar4FwLELVcJdDJ
OuxUHjkipn1d1swn4Jz4Fgv0xljNx2hBuhVtF9N4SemXEhE65JMSnW4+2J2wC1RIw0Pw6mSxxYH4
8lL0oZwkFuSNxc1afqcLNFO87wRPL7kPwtrZClXI3BR/dJIaf5BVrJVYoUxYuJoA/ETpj0VXsjiF
heqsXPtraOezD/u1q2wi1F8lQPkVz/ACb8o+6zMuZQHHReFlaYxt6d7/r41oirBoOqLlaB3LXU+f
n3S0enpC/f30yw8hrsis5CEMfz9f731S5MauQpyPy983H8LP1ybK/2Tq82hL78y/MBqYrdSALUjq
HJTSQSW1Nb14lFEScc4TLOdNWSDdx9z+JwtYE6LTltebIE9gLh2wfUd2t3PGmDVT8Ic0Cw4kHeqZ
fagpQ1IVN74bxaWdsAC4FjGrmWjwPj8c73+ebV6NzAbP8G2+6si1yxfdYjfR7Z7mLH5CAPzpWVBe
p3Amk3zsDb4uGU99Wn/XdZHp+BLISQPv9CUU8u/YETC6kxmZQ7SEKdeuqcjZSmQnXDsoUPkj6Il6
aLEPWDMS7jldBD8f+9qCVD2sQKw7UFf41udlKe0GbG8NUrAN21I2KIFdalN/Jm3PcyxwMabSgbpb
OQWYDEplhVlz7MQbnhjmhN5aIo8qyULNAMV8kn2gS68px7LHk/b6/gI3up9KqUu9bOZrjKVLctz3
vBYbdjHVv6ZkYQKFGkBc+mzyAUFdJeB+Gle0Mv1mab+gT7VOSiCRmh9O5jfrCTaX1uPL2ZjwUkGH
7AfMVGcvMeYAEwwOVLrfznk2EhCcgq/NgaOgi/ZAYYMg4ddhhrpZ1p7wxCXx4myXRsUcXUVocflF
GJTn3cYVIcLh6ZS25eKyiFwTbWKrym0NsLsoXfDbQlaZuSqe+6temEyJp0GlaLjSl/hX5omDaJAv
p+icPGPBretNMVoS9g/xoeGDoQnYX2ScYXrad0CD3RyeaW4jCR5+7zTzSLUoCBoN8XXuJ0hhdsMI
9Lp0r6YF5qqz+yXiTWTyuTzXcWNE+8z8ONWE+NmyGdsAnJvLfrKuCAjCkn/g9irCfoe4+aNdCB0e
UL9RPhEdubCADyX9qR7LPHNmj6eJcsl/u1WRI9ejnQdqB4FQ0NJ0Omq+JlQ2y+y/RHXokJMeVEyw
D3PjDqKIKc8TAnnPyNnAzFWGxOpzQW2R6++HyE+3gtYUPfXJcqRJimMDeDPoZB/gJvyvwupN9c+u
7t2pDHkO1eVC33xc2mifMiVprhseHUbXImwfIgtdC9Msko6Udi6aB56LoO0bz0Em+kr4pn16QUYo
Y/iucsnZ8Xdcn1qljU3AgiEpzA19d9ueY8l/IZP+qA5xA4WKObaJuIhuBqB2RHiw+qBk5f+u7eZ0
BsuHsB5K+sU52EV0xdlusT03czCIHBPvIKh+bhCU6silnumiW/3uSiYmFNxR5CD6Wf4AHT42PTp4
QVA9qHSt9mlD0zANxLjBwiFM6oiycWbyf8Buy9aRmIbpND0ouwlmVEcWbjD7C3aMVmB0xZ9tP63u
kng/SYccMx+n9dMdFkS/X3NtSw9ez/OC0KsOGNmlUO7o6R2l7Qe4v6RxGjinTIF0SoAFNsCWpHLu
i9kRW4+In/1kZDMvZaSbGdAkLkgd0sIdjvdIpfvQgaWCEuVB9rJE1q+J2Q+VCmEhqclZzaHyYSZj
adCIMYNQPnijALI/u4JJLubLXwdkYkBxO8ext7vi+e2ILgY2KZ0CFWkdD5Iwf/H4vchg2mvGnrRT
K18yZA4AW2LLdFeILa5nMU3gdAmufIcQgJeUt9QOYtzuREQ8r2gHwvmAMeYmJEzil+8sFeO5DnpN
QHT0FmRVYGGBHuso3nKQ5k2OBcqYysvprNvkMkNfoYTH/J7mAAxJQR9gO9DfakrdPiOZrohKKHNq
6oofjlLVFFF23hHRcAfS+ovx9wo2wtFRebagmiFts5p48FhgF9Jv1MQJLCc8SsRxEpOvHsC7dv4h
7bDEbcJ5V8cRQRomKiDcxdyS7CU6uzdfDCOBQMMO7r83RKOvFJYzOfQkbmwHtHFjcfimO8hFV7yN
nUftBUHOKmMuFjtXqD8sMHhnFbfTaEH0+BZoObyI6KfqTxR5NDsqZVZaKkMrgLW9XLCoIL55yLAj
/B1fTBcUSSHFwm/phetK19UG3YsiM9NUHta2i1HIePaT2K00AOgxewe9+JSN65Dgfs85UdLGpAWj
5DT7c1AJlv5OBZiAGSAOCfg4mgHE51rEcCtQGkviVWyHa2hHr+cmisoxaC/sG+Q46HJHLQCo5Gxk
lLoFmyheiZJ8EsYJn5f5YDrkrvXRoR2Ei7+7Rj8iWbbCTlAI1l9p5kroT0pWG5oFSnwnB5fltIyM
tYK3tXxyKXbBzXzua4+ImjHgduLBjeLLPgzyeFJkvKJnY/u5ovznEn3xJpEAfiD2U3NFMN5QAAGm
6ZHOaLu/gt4CbvjW6j1BTxy6SR5khYNJvR9Y1Mr/GlXVRy6J89YOQ4YvvtVmihXUATdDeB9CqLxr
5P4hFEgP52rxEZoz+4AVO85GH/YtgZXau4NefYsVSASv8OOfvJS9ujXbHj7LbyAwh2A7w3EKj+6L
19j0S99TOW48/Tuvag/IfscnsDUByKYGMHA1plH2HKFRhNMkyjKhUqzcmuR+slpPJO8UDZcTu6FI
Ce6qY1RwArKiBYD7JOm11QIVbUtDGFUkue7RAbVGLMjZ9wb55FAz7XvGUDE44Hsmb8xa64D5vt/x
Feol2WBNCQ8Ja9Fjilfdg3NJmOeAlGEGU+GDrJnQmKnQjVY58UwwFdq/jub81C6PfhkQJYWfAo2R
1fkxQXES3/1BxaOX/AH8xDx+X39+qEGcfWIXdhEOATAcMYg3q/MpNgOQV51s6gAW9m+Alc68wB7I
D1hvTAH8B9gfEZ9LEUsO6el4i7KLsmDNgTWQJrGHndN2Irj7EWvzCWVruQ+HaGXJ5j0LoGn7lX16
2YVk6ZET0z2A3IuLEqjdJzuzyIuhLphxLaxA8C5sa9R5PcNphX2Qa3f4fMH1ekp3IFB7DtdRjGEx
akOZLVxVv6GToJh7BEeTOfj1l2PL2fL4tc5a31ZQigUkbZFhP8mNPiBZM7YA1QFfDth6gy7Cr+4Y
PGiNjYJd+P4E0T3Gp6SNJt4tWPDGOZvUyNr72l0t+KgtLev+IhIWFZWtr31DTY7td3zqezGAR8DU
OeomFCT98dgVenicmyNf1M0uVI7iWNbZs4AXXP7UIf+uu8iO2VnwkKss7Kek1hEPPTLE3YTiLPu/
aRDaDRpbBHpQ8BIpLiMqCrxCWQfBvuA50LAwOnLT2zrs3O1VjO2hjefloBvdKk1sLk8h8EoXWr4l
0Kv3huCiL+hMb/0O70T3UAdIGfN0BYt7VQc/waS0Pz3tq1rz2BgtpDje/S7iSZlfou7O/9nG6Cfm
d/BLr7TGsD2z9uLiaA6G5KAL/S8mQrMJkw0WG+0/QEws29i68YnHAqj+WkH2xN+diRwHqDWDJvBA
506c0sYMYJflwwteQRyxau5QcANmCVESUuhFLpsHGJerxyvjEPwGbZV/4H2Eh0aRTlLQzAZ8gMnZ
XqGZmXAqeJMTrog3JV1Xkyuplhy7rG+Q6Q0hTllJYjN9kr+9WtnVScaIWmNEhu8fAJV7hjTzAb6z
H8efnfC+qLH7BqFcOBtRGMphf+dqz8bjq5oghd+8OovAN4VZLWKw5KkrQDDMjzb34bdqCsM8mKuz
PkJXVIJEmzLvfaGZmuO4ZHhQtsJCcbtmfB/2MCkTlhOqD8IlpWuO4KGFUqahmKixBlKTNIAt2Ucx
2wZ+ikcLRqCSizGQYfjbJCiZFzVrNGOizcUoact5m/0Gd60qTeEsmaobFTPGSyqVOwAlzYxa3F4/
z+ZxXuHz27KqrNyEQwo90uaw9aGWiMmJ54yuUHIcM1FXQhZCVPIiPMLndTznFzCiJbF/yAP08kEO
phntA+LpqGoRFPIX4ySNInw7fnLx2ETOYSmDqeo6f3oinlc/G43YC/Q1q3MUt/zORKe3hZi0IuQv
5Tpg7Pp8ORAXsO2qpJGTSAUX+DcDZ49WIhEU3o18OC1kT4ata1X/GXnIJhsou+3vVODgoVkSjNk8
mOHk9fqBa9dKjP+YxRBWpX2GolO8RmnfE9vDiSPAE7AiQtIJWyDgNSmeQy+AZ/W1oE8uGESvOY22
Et/wbvbfMHGVh0FU3ZtstNcv7crl0ajEXO0KD4bcrw338V0NbZ8k3W4YWSMvgGaobGSCq5ge1s3+
CXw1/B6NYxj6Twbz15HLiaUZ4Jpb3GaE5Txq94KIjCGENLj67shV6+qOoO7VmKqxYDzEv5mgtdyx
f56wD5UkmWOxkIwKwrPk3C7kZ1FcSTjwAopNhOgoYq6efpkpg9R5l5rodDyVZdzFYQotL/w+6hOU
L77xn8RLs/2e2Juf+H0VEcBMuhLJVjMsm1N2WQn3bmH4QUs0OToBgylgfhhNYMKYZEOZw3XjJ80w
z5G8jonktfRE7irw3vjc1QUC26n/wSuB9QvqvJ1EEDWE1tOtJaOGf8uhXf4sSKNNZFjJWdgNdhSn
eQbVzdN9us2OOjyt3myZBAOh8sZgQGodYkH9OgNbBPUtveQMgWTeRsJyBCJc5DBjLw9YbHmSnSt0
uPRdXTf4fytM/Hrvi7gq1V6GnLS3cpKAq8N+3zZMj7LoO4TcWbkdW8ZPuxci8Q/3rexT1AmX/Duu
ClF3mGFQt5Q1OQxbXGc0LbgDotdgOWk0GuP3+WGBLJ9s9dZn2RDUkPtlVY+Y34hYuRj/KS+9eAMu
qoh3HlipMmdj1d6d96OQVk/QUxVKGkUWepRnbyaLcY7xhoR8t0P7ClEtgxq5rtjXs0jI6aq3YgTO
GAUv36ZEEue+hC80DEZPkobthEh9vW6+GVWuu6AFKdS2xrpxboIbXmSMhexVCmVbBPqr/m5W7B5Z
K6+MEp3+CM4B7zp3geE2CqK0QLif4SDiNQtrtweIWXK8o6/V3DhNZSexlzdFJR/iV/p1vsHSx52E
BdEmTD8E2TclL9QeUbQoEbwWGLaIiY2H9XJGbY0S9zsIh2jQTdloaaCOFO0PyLlQaxwQ2vVm1lNB
z887H7j9YKcaEbdPeAQjbbi5z066poEJ5QSHu6DGQKWhRzZFQz/Mf8skIXEztT9yQX9rKtRl58aM
xWbaVUyUbEAtBsnytNFjqCXj69bzINZBIg/9K4WC1l3sEVl45ljRkuykTDFs5uMQez0cHfx45Hwv
D4KRvUeB7JC3CE0/XhaTyqQFN5DDrGl1HvZSJN1G/3GZcaTIIxra6pcMi9kr7nNPztH6nj4DSkfS
78HZt4RVQKRw2a+hEba32vMvcVKqmvvM3GWE22CWy8IyF2GdWcjBPEmqeM2AiC3lGaq1c3ZiwWcI
cSH+sMxcvubE6PAv470uN55N/kKe9pshYT1R7ejlfv//d4H7jB22tbKf6hm5NW3uR0ce9iRZbHl3
zKqD0OzojzmBBLfsLGGuCDwBpVMAX7bbrNWLPayBT9ALFH9F/sD19KLBUv/XN9dHNHcwyyuZ6SaA
2C1MMlmAqrgL2MkU8m4kSTOzUk2jqBLKL1pVm7jnzz80Cpl7OfkjbuKTb/FJmGSzjRIJ3N88wnCT
f+LWC/GHgbLMCav8FAKKR/Fgi323mA+fnC6kvMe9UouOx8hu/SllZpRI2IrUoVFACVvRiTZC2qfb
jkuv9ZkN9aEenHGHwugY2XeB9rSqkoyvzqV0ZsAr4JY/U6xoruAYOdkyIFnEsDp1/8hNJaqGKFWm
66NVd3OtD1d8ExxptNHazstnjQV5Ax9iDN8DnEbGpbwX9St+HBZQWVEuiGjia8i/KpnPptrAVM4r
T3p/DMztUJRJ6GaidsvmTzSps39jhmyl+eLy4kazN9BY/NWhKMvGVMjG/LkcBIEH7lPbCkwDuwGY
HW1loSrGP1cT8xuTMgAfD4dTS6aysTt8O6AesfaJ+PHDKRstqJuLC1Uwq0DQXP39kK09hj8sW3S3
M1RxHmb7ZhIsPWVCpRf3NxVXgMGLLNIzB1Fc/8cBjTDaoDoaji6KDrZdbOuJnFO1TxKw6SkWKWUG
METJ4vU7HubZ855KEbsS5sMYN+bNswhfaAn0kIu4+U+dGrLv9oxNpkhIytk3gZKIwr0yXiGf7fsE
s6db93qzg2fCWH5pdncTpg2X0/KToTnP4Ud/uuGfqWnAd4jRUnAbTGdclUtBDQW+jwdmaeAqzYJ5
7oQiAhO/bzbJDBLrvDuP1SDBsK1TAY8JQx/Oc4mcBxUru0zdM3K06+s9MGSutfBgRAxxJ8ruEdLD
KixSNB2jVwyuTgwqUmK2DzdMbe4mlYcMEVoz3rNyrPOudGcGZiY8MyZM3gWRYN12Qli1/1h3jAVU
1hWBs2Y5Di8Rz8VgusmG5uldf3Os3ImGpfCgZ7OpHP1OLuP6DD6MVcAAJRKkYevPn80WZqvvjSM8
2dfcgpskI9eG2y//7xKHtpL/H0ICUOLlXQJeyZUjB8pihRPIdJoMEmc3pP3PLUOZ52Zb5ihrjagB
s+RFuJJYJd50cIUbIgzPk7dYxnwjD1BqP4M/jkB8A+vx2HWdrSNPKuje7a0GfJiEz3EK+RLBZPWp
ivCRB2ttHQOG6Or+So+KxZZ+xTs/Z88bZJpuUF6tuROSaC2eiH7RXiIppBQiwh6oQb/ly51KmnAY
XzrUggZpC4nHct57chGjj2ztu4GCKmJYw6Yjco82gIYEiEzq1SEJxXNwZkkn+Eua6xnF4XT1LJ0n
bBNOU0Cqyr3XHDwagwlHI1ZMVDvtTcDKsZmQEGu7QBSvbGU/dK/2capEIL6c0yZEe/XKMWFJSzgb
Afwe614dWhW0RqPO0a0XCK9TXhVAjDKUL5erhKdcaBLklgZDLtSBh7lLoFjKZSAZ7RIUtIdGJKIZ
WoDzxaaVtPhbBi3Qzx+jQc0U2yPlK29K/GYV3J2WYB9iKDpYvr5vTtPcvaonzz6QsLk9VCi+Nm+S
+6MGDEZtvABItQE1p4vGFCKk9CORb+L5f8rHPIvz0uN2EYS6PLc80qMnbV7XigMHUmvwwyCPT3pV
xGKnqTQpDEVwmcY39ns6NCm1BfQ43ERu/ZJ1/6A44ie/vGWPO+oflx8v7itUdHkTrA/qwBGBn7c6
omGa3/yQrqv1McYOc19XhNxMCPwVi8VnMnh8uHd+DN+Uf0KZ56iK4lCovjcdTRswa/jAkHw/ZC7c
iy1RnGU2J/rvQ+7pIacWXexvInIUQDtHOO1JhlXMIog45MWgczoE0nOC3ASdLk8va/AQE0kQ4z3W
CYes2WF61FxmlR0oM8aXpW6xQjcT6nHUssCLr1pORDFkdgDl1HU+AjZNjyT66hmSRtKf5DQFDNRy
XeeLDV6jzOXE8F+0SAVQPggZSBHOmmperUNWBA+mu4Md0bXrmBbvSfg4dZz+b2fFUjxHsj/owlkg
PJtly/b8z3Eoa7CqSAGt6lq02mPXR9Vmcp7DzRemkwqkH/8Gh0j0dNg+eob2qEFYk9MlfztnctwY
M6fGsjH5ZGuzDE9Ll+T1l0V38sFivLrgZLubqaaEmcpsvmDd8jQlJfIfM5p6ZyvGLGjLlEslGhjv
a74JWJFrMRwK31nY617Xk8Scy4S0ftcm/tEvFr1iWUy4pMGlBuI2e13WWabMZo8Z493Kd8BI5SYo
qC3pDLUlhBfA8cgDVGaSxc8iopTs2LcHviVYgO6oPhCVdUlxWG2PmNk1EnsEO8jUN8IFywPD61ey
0gbeKgTkY5XAqgItfJZiSH5HCPJU2hzLX2gh4zmiTV1wF5vuElFxqXd/+LoC/N+BG7uIBxmXmhdM
S8P4m1fl4Oot8lMId1NTx4dmgsR3+NiU/+CnzLUeQaAjTdJWm2n1j0GPvIRY19gfi66GtCN6vMx6
xh8pV8nucoVcRi4QCsn8C2bv+4fN6NPEna3EOz/QchOEdFI6qPdhP77wHCIaiN/Llg2iKJDvUmz/
3lbz0yxcmxsTBwRLKAoIPOAH0zLzF5lU5jDeW5fFgKfl54cczGwWQLxgY6KiE1vPmkKv/pd0PMZC
rK13t8euPt/kQtlEKu8kEOqnUyTbhTesjljddt0C/YGen7U6j58tP2Wcb9nY5Wc1I/r56ZvGJ+Td
AnVwNvNuCdIK8NUMDlWuaKeoqlv6tA6AHQuLvWV5XgZB3kPinhQt5CsOSERm8dwK2cRHa8UQJdr1
jeL294G3KSJgQh4oa4go3olPTYFaTG4U1T0MG/f42qceNsNer7yr8AUpZsDtj3nQGEwGuGriT3no
B10yX9UHnQ8Pv2MObhjdYUpOHfUvERCWwgufMOJdV3XAN2o1FRfTNtWDQh5EKDQVGmhX4KIZvdt1
/vDkSqzKjRTOLpLgpPMm0xNe/v7FfIFe2/wXRn4ZKgjhkRIax8H4Oes7Cf1k9W2Wftq3hoh7qnPS
Cl9HBSoLIRIAIQSXsWYfm1vD2zuJWfSgGSvvPSc/jvuAI/iv6BSD78LiGe2Z7XzVyTqcs0JxBUaB
2L2ZaYrZnHpC7GO/y//6AQvVQhpuepf+ijMDNvBYRxMGKKUAlYKYLYKAKlSyQgPI/4xeucHAWvgL
RezyD2YQkELkX3pNe64E3ZzAJT1fEsfFFWmPNI23DT+3DEoK8PST5ObnBNcik60P1mvEDZThC03M
dK4IWNGnJF8T0kzam5t65kbHhQ5CTWlrvXLH78tgQjqy4n0Z61GDUIZgUxA95WFv+xZJLPsoDpN4
IQ/0dRKamW1sUJ8jOUhuDBO429cVd4Z0Sq0gZ41WfDTMnS1xptCUKESc5gumuk7DrgOctYShoafj
D4ozNJ48ym0W1zxRi6S7YOuRdXmdAwZPLLMik3IKzKvDk+OnAisXxbJoFCkfI/FkBJql6VtT9QxB
g/P/+oqH5cw2ICIC31LTtqQOr1z9VfpYp/NF1OzXYxpFKo4gwOawmdV3k2DJgAAyxxsut2X5WZjz
qrll+sQL85PmeF5KzH+KrNXF1L79+f4g0ngbAkZyQmVl8HdLfTEFLxPHggv6EM2nXU+s/Y4qaWM9
6Ck5wvDZtvSfHI6pXFBo/mq+sny6jmaMVvgWvDJvTNeVh7ApQeox58fdm2ym9ziupNCd9mpUVXXh
MG19Ur7IHNZ0nmYJwoWzC1QzyKneS4is9ca8a13CDp6LP8/jhDZiq3ZPLbgOaBUzW0hppZPv+x2o
wUNjJszMwIm2xXflnNh/dk9EvSeap5YvRVkHZ3Chke9RVinizMSkYIMovAlrbGrqfc4cm2eZNaYA
YT8F2eFWlEIv/3l7M1vLQauoskgJGuHoZ18rbsf25foel4XFA+o08kNMgq2KuB7Do78P+9IU1M5I
vduL3gvoycYe4fXu79VzjdC4KaVc6tObWolH2d4heS2xr85a8000jivXD24XMUPa/rXA1xqhfCnT
FSgSYDB62VdQIQAsGOorUVlISYYoEKjVqrcuIN4lu7Ce2sm73FQkcFDp+hlQSQD44dxeAo/d5fKW
8iTK4zLL1XvPQkWDo1TAEUqFNM1Sc2KbxI/C7Dx6Ts822Xq1trK0uOv84XtW6dNrl7OlrVqAGEee
GRhri5ZitA2TwG2AT7JNdkSv2XDQbO1+NE1KPQk2EoEz563tTQriWPj6IJdT5wyzrUg9ukt15zb7
DQJwvv1rivIsg1cD0v2P4sLb3dWZpSICZHKEMNb/d+GEuv/Q5bYaeL2fGokM6QFr9hRz2GMyxksw
k4hgPF7MAPbviYy2OcTQuN3ERULwU8Jjxg3gf+d+WiXktVfH3EpteliI0Q2uSRR6lWBkSnv9vXcH
xeJK0iIVf8PIZuogn28siSDxFdh7xXUGDd6SJGfOS7kL/4pAFJxlM6594zeydznm0I14/V8PCh9P
zw6o0F+8znY+xMh0DP8gY3jAtZ6JgmkokzWkIX5bM9DbVemhImnN9tbOvt5+TX0wZvpkCt1DLTFc
3z68gFAA6jYdP8WJG3DLzbD++yruRqxEdSroa5NL5x9G0hjD2psAbfiorWC4ePzTExSDvPejcUBb
2SpMWhUVQ0on6QXMwxu+/WYGjA0zChEyXqFg5hlpMLZ7GLJ4/OTXkq/1sDmKVtiRnL5SvkJC+Fiu
8M9JA2q2SY1r9/VrzRlNHIyEUmcp69FgM1+nNS9jl1nsyUDtJACrYmrF7AYI/rT7N4ANA8ntbrHC
9MCgkEBtwPt7jY9r3k+CK7A2c83wZ2uHlMIL333Nswo7NlX3+JjCT5jrzCuNARffsm3KrYlE82sU
XsE5SdfZLaJcNavJZ5LVxFlBi8rvh/DjhTtj8xGqeyyG6v+I/mqATCOMg5bFVbOPr9QlQnZoLlqD
IHumeX+iS40W3zHwq1kOPbgjJ9b2x8uzVNfrFcY0OwcGouJ2rzpLfuQwr2VuB5iLh2Jg/a28P6vq
3tKQW/E1ENBWpgdiP1CqeBzHymy6ub942fE7Q6hHyrpXxVGLePA3k/U3/PHlzwbTptgJKv578NRQ
4bXd74rHMlYyPbHnCQD9IM1tymZ2rjDZarHaUKYHwJTR3YAb+DzHsp4jzCInuunObxBqZ6nvfVrs
el/fxP0mvE87cNeQK7liwoXx3JuS6Xhj7xi+lyxHO783s/x5lEP6tj37SJjD8ppxdlEHIFSSL8JD
sjiCPMC2FRhdG/lfxjPVD10nNGWCSXnjCh7Ki5SPu1Vp0lYUEMBN1Oxj6/Ghx1KUfu+mMvsPO/fH
j3vXo+arw0GOWzkmoarkEazj5f/G6X227Bk90Hsbhg25oLypQczB5LEdWa4FgV3qpX1sxt1ARscP
WGFImxWLt0I8rpUhpu6rAr+jBRLyzWJJnd6OsxFGOl+S+csZLghWs1WnXppsRKG3VTK+4l5GO1uy
tw3MuN7MEBqx4WloKemUXcDDMY/uomzpFXEUzJ/byOy0ewpohudgz49WflRBtU6379DdN5FbKw3g
37HhX8xfXHvB7GKxDiZPZqEoxa1zNN+rl0AzfvQ56kbbdu8IGBEouzo/mvxhJhl2rpTqbufWRCZv
D90CIw8fhs+ayCqolKyXkukx+khe0gc35XZM42kPDngawcNWG+Ax/tXTgFLP0/WhYNOoeN82X4rB
BXEQQU2nVSv9Et1MtonHE/B/5GPtRE9PVtMJ4+pkmTJ3g+ugxrrFHRJ5nokeOy9fpCww4OvEaTki
zUhmdAb6LRzr39R4IYrhjE3wXd3GxEI98Bv7K9e2l2zhrn64RSjzS0KUu00V5yIAoFF6lpwFIM43
Hz+8vpsG9XXUcu4LtihLWVfAfhFiDJ0GAphnxW/UonGmzIVVQUT9TSPSVpoySfR1HPjV0jPE85/X
hAA9d0N5JM5Ecd3LxQ+20p9MEdeUqRd0FLuU0zzto3QgDGq9toUMOlJd62BF00/D/qVIM1Qhx2GM
HnE3rgeDLQE2+A9RgiejG3b2MXcibROzk1hGLQnfMx9f+0kXSKmqSB2gMvxrTd4ifc/hnQmwCCKl
qg7601qQ7biTI6o/c1itFFHgDmfyNnIhMDmmGBfl2TeWzWazCOtk+Ob5sF+s3ZCu0bb8WUFODNTo
DL1knGpuuUKO/CfB8YOgrPg3IEKNkMXZpVlyTgVywZpdXQ83iC2f6nUWpc3CRiwcLyp50/On7kaS
VFETwRVjRtDfUUmIpM8iAPlYJu2wAiI8CPCnVnbyaeOrxeedqDc2P5oZ9SsJN+UO4iZmLJt6p11g
+Gdcu6gbTFen3TJKT9dkw/xdJKI8P4MdoNJjsyeglssv7Q57PMHuo6PZQ9IPlFtrSB8MN7y0pNxO
FaAcXB8j2e/BAtBdxkSuNsMNEOV6uHQpDpS3ofwhEqF7vOfaH5jMRMh8NTS+vhWZQRxpyfNHj/mI
DZIsZHNjrNhG2E60ptFSe7ycvhWtepE9woTEe7UmYjkRUPHzta4dkxDu+8HeNtUX7nHTHtdMHIQk
+XmDnsmLoN18uzE5kvGYtgMDdN1rvL+67A28M0CfIMDv6bPWjWjmaL0XWG3j9bntTYYbS+psPbao
pCsjOooGl+JsYMVID9LUjdvlCiruq3LhRy466++/gusCz2Z4IXaPqJz5n+e6o3oXIqdko58snG34
IHvAllSus9AIC4LSzEKwuxbwd7iGhl0XAQb4bpLtlnbS1Pt9tawRIn+x1UdNyn/oSVS1VsmitE87
9lZU5na0vc2rtv0KKsbOGg13i43yP7oPWhvvsTB4f4ZIda/YAb9SM9YswWt3QlS+TVF4qfpn6XkD
0GxZlqQwRWCamjf/tg01TWw0hLpcSETG+We0aC4F6pggg6GJhOmNzvHTF3ZEkwQN/YCH5XCMJuuC
KKVF4XyJOoK5rc6oR2LqcJs8+0fkSQNXbm3PAe+6zoXozT3aygFoHI+hYG1Zv0FWIJPqHug5cSrW
QqQ/vxMVBQYib+f8Ndg0Xd5+fBrH04Y1xRbndyevzvk6UJ/+SRjatuE8vVm8VG3OFeEPGKJXC2Ci
m5R/9NDPzMn8Khs3bUHwiVGImqMK7PBgS0QZno1+jp4m8LtZwlHEiePy0Vv3PssYUSYDglZh3vtR
MOX/vbQK6S+V7jBtivUjMpB4sKO/8Vg7tda+/78ruPix+tztIrCN2vmDqmr7pgLQAFjQ2QfTVR9S
pwzl+yGiJ7eD5BMQjRYbIBgeo01ZOC4e3fPn5C1Cql39mduQ74WDVk5PyxNP9WnIEU66iREaHZPt
UAbRrSl3G6I2h4zkkzga3S1DMStY/gNwhrHgyvMvzQ8rkuHbxgG28pg1vzfFoyoUd5lY6kiPQMCJ
ZGishlfy0i17awzo1tFG6fUt0dig4bJmbZLTdjvikW1JXiVxuihgQ5o+yX5/kzpu+KPD+HxTYhDf
5d7iotdrR6sfRNWAK39VmOOEIyOMRB1jZ+09xFD3XrtUPBK1rtQYJl1AueRmCI6abxfWXd9dFfYE
jK4sLbAVCNwxlGxE2oTOn2hbbzoj4clz4W8W0jcM41E8+DJQRcER3sIawKu8Rpw+8R5/V8o/Godi
gyJ/RefJ2gSms5UVqjNL7koAJ6GXNYGxKdtas0+7XfYEbMz4nI8zqD5qrjKAw+hAIQfX0vDFoYTY
BSL3moDYKOqs94Q7bzCy+UoKDUZktEJ2m6QJGHVHOXBkujIRfYeq88xVkIgJf207H/xZ8Fdyh/Rj
DEJE9MR+ooRqgcuP5QLTWVt6adM0pdGjrOQEKzm+hXHSNCnjN1KM1kIk4DYp48ZXNkkAjxKI2mfn
H7rWeE10/9qhJevz9KzFe3xbH14/TppkDWl1eqP3zINRio5aZjFgQbl/UKQPUCxd8+UEplZr76bR
bgHyDOJkayLxOdALhKyY/EV0Hsida3h6Tyidqoyn6gw2yz3mrc958vSzj0YGWfpx0tuoAjolShaZ
vGKplPKzLxIAP2LrQpwz4aYs9Qvw0eRn8hC5gKqpYuMMwCqehehU/ofRuns4fqKz6QNrXKNTd7IM
b706RKCmJDfpoi0DXTzHIA3QYjElFwpekpzdgYyCtXDeWKPjdMcU2jMhMdwA2a8pnhSeOMr0ttYX
RL+PxXLCE0GI2GCmfWMxfct+nQuxHJf6uthiPV9YCnenr/Zg6vaiwBIuiFZxbprW7mo3QxVmTt/D
3MAfhEY2vOEDAsibRryeMPgAZMCVdGbrteGLxcFavafihwcgZCUrYLSP3+6NJW0OR0pzlZdut4mu
y8HDlk44ncC5NpyI8IENwjzyjF8F6Y+SUIkgFx8hEg2LdlFgPqqAgr77v7qimQQlQnED/tARL5+s
jPXaSRiPl+qYuyDe1nCWnJ2dwn0VCw/Y8PKwqBU8ykt7ITMLSeCmwMvlJR0/vgGWULzjko8OjP4N
ZYp/MjelSR4lQtjMb6yKcSh9NPxgB59mAsP07IGy/UHst4KarfPDMMhTq9HclPDziz+YYeehtps5
HTLbpLADdRwTqZypk2TW/26L1zXv9FQYwLS/MraHf25V5eSHOpXgbGmV4nOKVZltYbJeJ0Jfazmb
xAdivO/WseGjRD/DYAkK0Gp2rMnH5Ru3Lj8v93Bm2hg0BVUi7f9Xu9nGY2JMtvkY+SV9BePd9UK0
QBBwYDKhbjFVPO+4n1ePaIRUmSEndwf61easjdlb8Kyg4Z84pw3YTOcS1NqIgVTR79zmcgv0gKe8
vp7oDRG4qtSYTZclNK7yJhivTeqsgmkRPmRkkgP9z5xV5Ktwpp3B8omvbwbwAviaaK5OM5EV5Xul
AxK6GjTb/RqJObHS7m6hJmTtihGKnQzNUrtEGmVTWum1VfxWw4zR6PtFXoRbvItVUGc4vCF6Iahk
k5nSAX+ftFH8/C5Kk7Oht7r8j7MBlcmrsgSWd6ORkvAKCrLiJa8gaWmhfHiEjgRHUN0C7faFtj94
k9B7lbsApv3EL+6pW5lkcoR9F31b5R3jgEX0zyRGC8ZhX11YTUzCh4lxcXpSTAHgqGR9J9Fbx3M3
JF8xCJymARc88HCOuWGJTWJDzmHrqeVyapA8CAb2W5SAi+sUr8HfEKS0LEyvBu6uBmLZVRCWKEw5
6p+GNlAePK2X2UZK+OpCy/dqwtL6NTXgEAfQN7Fs3gEIHqu9NLqUpa1QZPLI326Q0coQLIDFOBcz
0NgqxmTGubaoiA8bbJaSHwlOQAqr1BqHWdajfmsK2ysksa0JKweSumSr5Cdg61QwhCqYoB2TFOWf
QpHxSyelBjUBtIydebDeNt0oJxOlLHcoXsmiQnIpSEVQW54WOmqiWjOSZU9qQn+2DypZGVl0ML22
6L8BQMdhNuqWtfNOcHtn4j9yEZn8aRC/8ffsUR/0w6oo2R1ipIx4njOtWWjN4cOQMAkWXtd+pyRa
eItoOspqnowutpD96QZ9zVgpwDEzWXuQYw+umu8sm3IOmtCBiZLwEftFvUimZ6hukYB3w73Wb22n
ps7x95A63OogSJuxxgY3Z7+WEO55db/MhGBOOtAsUcE/xTSiJH9GMOQJsznj9CmWPrq9CoOh9t+c
+eDTxxY8YYD4p4OSDkOkOliVNQsfcn+xg6RSzvVMCkFw7pfex/V6gZorK4yLpnv3zHZd035n2UgA
GJtcHeRQfyKFogRpxf0O59oe08XaCT0bVff9co7XqwV0pGSt/fz4JinogEvZR8vUd31/VGNjQ7Vo
WiSEOx2NPOC9NLBhEQL5Z9Oa4ZZn7iK6xotIER0QWr/AhkxjVlqpmChFjH9Zfv1+B3D99yrVnYvA
AouVgYvTcOZzE7Sop2fnonFoJAE1LtULYYaDTAZ8bYK3KAqJZqoH77G/OYeyrtc++C7lCNx8nXH5
rKEuankMw//jkavSZb4CrOFEaayrUhWiuY3eEOfzI5SD/xLxGuomcvkJ/ZdIuJ/xlWAfWcX+yB/3
B+v6F/79AJAqYs3tIxlW+zDtxxQuUUuR74PMl5Xa9aZr5YIPTqTdfRZJykwy3pOqZC2bm8Gv+TaX
/6UtJIL9XN0SJvpQqjyuqYcxxf+zrAyJf9IFNsRqAvvMSlsh3jAdFpcIt9259pLnmEtgTUHtDBX2
7ozty2TVV4k15YJxu7PcG42OW/4JSgp9Z8BS1lcDd0wS2JP3YO8St8BSiBhDb3m4zFy+1XgML4fh
nyt2AWxYSXOiQ0d0dXUsV6S8thnBeEu7ClN0XTXZApd0tQ3xFSgcelehqjjQIYKlwXxIc2+bFAMB
lOybuAztDdMEmgZ1928+FVCpMhG9dWCyT7PlTzMZgH0uJ/VUuS5YiZ5FTPzP1tSLdSy6ocyOPF73
9l/AKZ7XNF75aNtaETf9kl/Ma8aOjqOIv4U/4gV6y8OFyL6AkUdfBgOJ/MXWYSAvSnCP4rwPjiCj
wvIMOn+Gqgpra8Mhs0FNPxwVev+jA1FdYyxRJJr9ExylgqkMbiAXZr3VEErQG3+CA1HAmaz0PUYJ
d64i/29US0fmwa+K50K9kKoIx5mznUyn1+m7DAeOxHiF1kKQl1v/jKzJHSmrmIn0O453zlI9DiKN
yD4k+GdAqM9S/BtShGWmdk93b8eVIbJkFlgFeprP8u177dkzhE1YhwIo4TH2MoeZ12YFBAsCYKNZ
zYu2NIll97kj6LPPpQNzJyC+UabsEfEfyV9JhfODwlO70ut6GR2Nvpl42gimyJDV9Nvoh+aeahWn
CtgUONq2L1pi5UZNamZyOFx5ygQjty4Fr58CUJ7jMx/HrVy+TsCoTY6MpVyTEi3IAr1MoChn37Id
LvlEICt30wIE+Q5u1zP2Vp+CQHDR+aOBm1gM9BPO6ATHaHg+IkP/YpdsCVSkanXmVijgjjMLzFjf
cOOzJDlX02fevrgjWckaGiqlHsZFKc1JtgATGjAmVtOklmRSzN4shEPF135fEscyZZjoqv+lmlAT
bR1akuQzByH1TOsTyAjuBiYLf0NxjRJ4RLAV4w2LJ9jIbNCShTVufX2vgmXTgleu05A0zMlKtlyg
Fja2jFpj7A6VlwuOYlKkZx9WVt+6bymyJPlu2ro5rIDi0mwlcLlcftLf0dp8irHCEwYPgZEsb6hN
pg1gVQIO10pc6Litm2iIjSe4UNpy1BudHblAlzrSFkJpnbZjY8AL+PFYjGytQH8uDsLoR3LejgI3
8rNiMGQuNgLfwRXXmM2c2khdvyaBM0Bxh+PoPERgpbw9fA7e+b/SN+w+5UWH2Ss6LhP5vhcd5ho/
8ASHbD/WjQnaJ8HsEgg1sdrJ9MzwMLw7QpuaH9sS+H/PnbxzbWlrqgT2oRTElxxV3wHz0V03Tcjr
881q2gC4xsGS6gsYGpFqPisFLvdVLbz8GoSGIH9GHEhhtf2tj5glM6whRuTQtUtCsHXrwMic5bW5
hpDZFKmw1KuDLuDPln0S/HZFNAkkIf5+HZElhddwApY5XraaPvtC2st9558N4DZPufcv+scItGRC
ko2m88O8/Gb/452Y5Arvbtr1ghQin5NkyAbjsi8c1fcBonJTGix4tX9y5/UWXtME7lv2NS5kqmzn
Gb3LBZPr4V7yf51vJPd/MK/xUYCEuruEc6jC7dO4e9FCWdGnvtISPp5zEurjtUC1dj/8kOq4JwnA
qSAnGIMqN0aqHErI9ydn70l5lQACNcjOrxVrA+8haegS3c4TD5FyDmrgFnwr6P7bpLqrkmtTMIqD
BwRtz32HwmN/oXfbRAbTt4yShhy3CEHMnPWvVaRI1nDMzM+f5bIBkaKz+LXzNxABEPeamz58vxcR
T6g5v3ANbPuKs0WbUtPeg+AJEleD8/bSI4gPoW7q3v1OxxynEQ9YMP2h67X7JYMQkL7qlBYmH/95
EGN5fKCNlNQZLnzQYhcLGYf9JsA7+xxk63QJh98PY4wOOeFrgwiJN5vpqc50cc/Mp2C0U3MtDw9B
ci7gc04po5IQg8lQP7D4WxiOOEf75QSpKuAXAH6HZjOJ5K2GgY81MEsDTySXpV58Wi6RNkt7xW4c
NidoMF1nQz2/x8vwuHs2kfdpbJKTX2qRlNGP4BwTbx4BvSYYthku3eAnuDlAmR0hcvcoYcx0rQww
ulHcRs1Cahimb56M4uTyLZKTgn+xXWlczsbzDqBsZTpVGuv1ENSMqqJAv1C6sXIIWtJ+xKxSIffl
qEJOAz485LNYO79waQu4lbRk+nfNCjIZz+S70VZfE4+j3Svo+KLY14w4/sgJn5ZnPlrLGZFtm9gg
j2ClMePhr+iiAlD0VDDaM0EeepDzURcRiBh7ycNLKOXCiLp/beEoxfv8pjRuLvzMe7kJmYsB6ASj
ojKxNEdk0dRXBQWH8VPKmw0hDfTIFd1xAiTq78zac3sI+XvFes4vq2/K1q/Y9w2mxgzji7+fKmJj
L+HEV6BMAuJoLakZlT3cIqRWcm3uULkOkZZyYpCiibgtySDmvZjLZ+mnIYUOj5AoRNwYJYBBFScq
SS5kkk0qRc5HDZNR4BQHfBqtV3ffFTZYwCO1XX79TSIqG9H8VphyM/ZxAJGVI81TGQAX9d+eHvoO
1qmF9+5KRjgXYOk05t8V4riuvM1PMBYTWDuIB78F/NKbYvZTxtdyrLCWsU6XfLGL5HhgmWNuiXN1
gUmH08lvf3UqZ7SpXidaN59F/m23WGKrnY6CuwrlSeSf2KFL9INtm9sifH8wCG8wmuWFsV4BRKHQ
7/PvttukVHYqrBiR5guBpw8K4QeY59cPHvROjVkaRDT/JjV+hMHGCHN/ZcfJ44Vb+63N5cTvFPNG
vbluF2+ceb+hYCLOCsW5BHy6ZZkvLOuwMBzZduU0uSKucy0wTRZcP590xKuEOfeA8RGyr25vJrAF
ybx5SR/KURdr2+ZIEBBP9wWlBIUnoGjQ4q3QU8BwpxJW7AfSbCZanMIeHksTAuJt76A7xg0e28/v
gHCdCROwyJLaAscaJYeTlWbcQhefC5icKmVW+Hk/HMh21ZnHUvf+CUYTua9WOOKgezM9JmKP8xVs
UKEgHQ2dBPXAjgOGLVrCUNiKcrvDCWufGWQkY+sReK+AiEHJVJjqPgalkuqi+imNZVFixBrqWv06
A0oLxSi0g1BNzxGAkfcCMgwHqkU/UxcMjFHv1Wwkq2E44tXm8/vKCtYI4SK9IQ5X72nZeC155d28
IEnzu6JkCiXF/o0hovYqOFxkbfY144QRUbF1GCdmr1z1aQpmeM47TM6UyYVH2QRQZJj4dTmDDjV3
nQNfljyVwIwIMOCxS+vnQdtqy/E20QBAGcdc+ehmsjAJhLIm9zI9vo9YjvPw+seS6V1OTc6mV9yl
0EZqVq9TNI1Ux7F1ibmJH/eBtGzi5Cvr6fj/hMB3SWYWqxD5T2drdFY2kjApSKAnpcBSxRPvsLgW
yNtjfNC217zOou31wLofrG264fi9RxOiihTaxEmmGfxPUcLXO9S6K59Qklp6qFurQFxx4Gan2jnZ
kmi5c8o7VuTjNuXiOq/yoAGqIIZSiFny0oEJsd0Y4ySfwFYrhwL8rTVQFfcrKKYJM/j2a3rnDfkx
ZqSxIWS72juXilK0u32AyxofLvdAoXRfkkx6SZDYrRUUGwZifGfLmW1OIpNu+Qw8CSPb4FPEIvS1
+WznbtXMoTStLrD3dSyCj0x8vbuqubvicMcLjeZ2wWumsE37G/g8vth64ObLZLJPlafGahNCvfoY
4Tyv/g8Yn9E6U8Db4+aWVE+Oei5gKFvuMSwSPqmKcXR6YA1y7QuANUMJHySzufUZL3sYsaDNTrLN
TQaxgbTqMI+APu4lkco5CyJU/Ahf1djvxMDHGDmwGbQkMYRNTN8ECp7mEPxU2PT5wIydoYTsiqRY
Bh7teIZklpCyhGq3Naqz7nhTIlTpYl71bjPJwTTsyrZz1KRmxHIH4bp162aHElwKPEEfC517WDty
t5jed6793q1WTe+GYtcDd9O0LI2rfn9scMstiU4VV4ct3n1lhJydAmRD+7xfeXKBtR016S2sw/8E
2iYN0I6bLZsD0XoiaVSrF9taHa18gujQgLVFUR6LY4Y0PLDtRzGTx5GbyMVo/fI41v6+x/n0hPgH
mZizvzA6zhp8tV7/2HGKjljx8GDRxTvT3pYozo2RH+F2DtwbL/Wk3lHdV1sYtFMJLbV7bGj2Iqi7
zFbC6AypX3lqPpQlZbNR02ARdyjxrLYS6W7eCEs3H0ihWvjnOI5W0hf01OBbXGpYRXEsGvA4EvwD
J1tGfsZeP76GHtpTvxaPOl0eQDcPDAiXIr0CnJVcM/cBlBQEzIogORx2uFnLb4wp73k+xQLy++8y
6iJqVfxjwt0E6A1fbJD02uhb6bVOGDij7Xd2TJZQ0shYM5rM36sbpBm68unnjCez6gk6AtFTozQ9
Dd4XWUmV9LQ6trNwrbkNmfEjDT/IUOGNUfiy5x79yDLJUV6AGazrM9cKr+ZxIz8l3HsuScaoEZFe
mUgWpbLex1k3r9GU31vLeGylrO5TQMQ9/I6cjeErE/ahYY0gLC6vWfuc8AHFCG+KNsDoW2JLOPO+
+rllUgmZgvVvQc238+fPcU/zpQqYNdqw6rVlQ4eXyvhGu7OaaVD8EjDPJbzcSRsnsjBQPccVBGFp
jDpzl5MxBdmqmBudW93/LSXx2BUBQ1dWK4MxSrV+3GlS1iZ/cswOBYDxBUwrQ4NNlI6clVDKA1qC
JB0DEru0We9ickwK/xWCIhrOddjTpWWnQlbdxd1iAaxvq086Q+GuNs9uep+E6/s0gWrER2aClGUr
l5ZNbkU7s/69Vvn5lss6BKOXWbNYTMElgTVSNgveosQB6xSbamFpjt6O0pd5zUkVt1Tvhz7K6ik6
ZziAXbW7sAHMu28ek+AY/aMkdlmKSsM+3GkJV8P693eBj4pDmHDpF4B1sPzjxmdM7ULSfVpMqWkc
KuESFxEtQl2P4D6DsPJt/EBkDBiZ7+Lr0+QVczHg4m1smlVTrIYrlAoomftIStjHuk6W0iZdd+6a
Am92nCmxvRYe4ZwFIXU+vFttRNw5x/JK9WQyuOdkZFr7GhU8u0lm20mRHBqsWM+8U3rnFaQb2yPA
9vu5AWVW+Jv/4C6hsF5VnctLiybOEUJth6uja/wH3uvSI8g+ZH8GCzhpcNVj3wH5j59wamTYmC1f
9UiITnUJ+7WJQmbjqpEnfOY/px/xouaseuIt+umYqvILFf5LYbCe4R2fdyBw0f0mS5Emo7pNCP09
NIv9AuT9kciDtpwbH5tE92yH7dYesEiJmw71wnc/gfM/ku1c7ZmNfy4Aq0vyh+x5iBOFRLhCarQR
4qiHR4XnoRx4eFAq3YStLHrjK1C/UwzSL46FPfKUO/VGo2l5xyOTnF5nhwT6jdOSgZsmSy+kIqPi
6T7IzxpdOVMXtPeTrwspWbhd1RTjICkE2tSNTAj03mG+E/wt5Oeeb15GvQ1AVDjsyWUHT9cZ+NEB
edhzxcjQ+478J31tXkeAPLg9y3yDVhqjJlWhQMDnsRRbzjN9AXCrlapk+e1NB5cbB/TN9ZSoko9x
21KRF09u+PAiN2FbPiVsEHeYYfw00EFLSd8iMK7Jn5Ea+EAB/jQZj86bnaY6t+IOrQXgz00aX/uk
2EM1cwXSbAZmAI73CvjDIWYxNJ6At0K395bxzmatXahFD6ZFq6eCwjPSAhuTJWY7U43uTmutsNx8
eT/J4WfdgbHGsjiwgR88dVx66dZAiRXqd+dHYssNSHjUuXde+7htPRpxsB3YFL5W+zaCv68CQPXD
OzhCHi+L3ZPZolNmTCZHQ4RFQjqzZudU9wFlwO+l1/SaDvT7W00Oz4UU0saAmNLIQcJ4EVcJIf/z
ixTPcn6SNSSAX4Ujk3PXbknfdRc1FJI8t9DI4Usgd0eOnVO+MsuUXgsBYxPkrraUQUuMAHFIoF80
qPw0++J8/E4KlK32pcJJV/rGcqZnS9sr5p0tm4dKZH2/bOWJ9zaxG7ORMhFJrL4ULWW2ggDM/RCQ
8DQjqJbV8rpR5CHX/50raUNXi4Izp8tjY5sgdAk2g2PtJqTmRNQigQ0J4/jGyIenDhCnbzljCHn4
qrWFUHlDB/uLhAEJj8QmIv//71rgij7ViUiEmei0jzYRJ2Nkffv0zseRItbUvBzA65ph9ytuMTzT
Kxnrr7ZOi59fXtXHc2GDKmRtR0yQN2WobNwLz9Q2GgyfSR3SxWsByWnKxvfdMAfL776WPyXiZWMa
cQuFmZTcERAWTQtIfepKYonk8rDC5VMzE+sR3RzPcz9HNlmj23r9xd15Bc8Z0sJwOGY7CM54OEhx
xlAuMRCV61IVLsDmNfXDC5JmgRpFyLHyyj5rFMyAiegwaAvUd//yMkMeHvmFhTAnJMwAP6l7a9Cg
N7GDbilt87y73VU9hB+w2DuY1wQK0skoBdpeuYV8FRU2qtUjxmiV+VzcSrSDn7SvhXpzvZXgUu2E
RNoPTI9L3btIxHrsa1mohuRcV8FCcyF3EQBwnBACWoqrCzpTeh7FcZX+JV0Q3QeUN8edbV6LyJ+M
8nUlAEp1QlF4RoYxlQhGSefl1GMSih1YlIxHtTW+5r4xuHrPfQPiAzDFplQA/ry9c2+pBA9ryNBe
2bYFZtEN+JbuKoqBUZrnqC9Rv/uJE4tJMYlHm/L2YmZiGp4YtwfkG5t8LhO2xU3+bXkt6PTmoewT
rrQqHxLae4gHHTTw4tcPU3Rjrfy66HbXCu06LS6EVkrbxwe1F34ak2UFFL9pSD436TrpGrH/rolm
EUPZfDWa7yr+S0Q/rcDqwwFii6SPEYxKMFHwMQmy7t24A3XuxKvavIO5etlrDfaCgwwww/meGYRT
AQ8Q0XbxORUN+mh3v1DTCczo+mGhZxn6VGTvbx9dl2EKHs5rBXdqv50fm85eXEF4jrsYOWAS7ePl
Y63uqdbiRpQqQsF65xtLOt++KaDrZwiLK23lv+G8olNBE4TZ40xwrjnDQaiT9U2taH+qxZfjImmj
yWKdybg3+Ny1GjgVsktYzRNBYD67CaF2VaFfMBjOVAUiYaqGxmB9l9ncub0Sx8VMZMpJeEUCneti
JO1udYrkhXO0DhjPLhICGnE39BB3wNRVtjYXekr96MtAKJ1UzuWsmQ4EEeN1eOpaACRuLot3Ta3G
2zb1DeUiwF+AQ7iS8wNbQuQ20+8TISEpRutNt0ebQKzvZHDmGE9KxseAer7LuVVmSyEaVaXA4Lqq
xppugBVvOYKARZ9PoSKDYX8r6NU6Jz2kqI8txVzQnsjzx05sTC3zvPzo+qHb8ajlWvxUEdU0/T23
Sa6+KeVp9HGLlQEpkIVQRCDvbs60Y3K/kw4r/CGz8TeWlefb+8fjmTggjfyydhwkxTxbMia+8kgp
+O8X///jRuJL70qddTEymSUYUtCDDwU2dNfFkV1ATGvpB3Z2Z70hQ+P+9bp35i6cZmhTH7KVCphX
H/j6ShO9DhcCjbaxQ3GuAl9/r7aMogO2CtyI06rdzrQ+0iWPerfaA4GsZC2xydBuTisDK9zUwfwJ
N/T87VeUTtk5C9/ot4FWFA1Kd2IBdv8U6qoNdNujnkPgEoEmr2khb1fP/ztEIjmzAnufFJMURN5+
7FayqrMes6mK0/+qg5ayTFgRuSGPS2CopSXXrSamkevZFIyY5SOuyPE/UhqvOVv246V1ClICFoz6
Dmejk7a2s76OmxDAHlipIC+8ses3ImVc2/ynuDZPqkRNJVze6FkZvs/T+9Gt/VWt4COUvXMBZo9X
kWnPbyE9gcmSY6mgFLb+zetLJzs510sFVDd7c0ITcoHFd8MORWgvNtpIRZI7i7X7BMrG6DZ4hSAp
mD1ZnktQVM5HM1G58Vms2Mnuw75BJTDvHNN2w8VmGBOyzn3ICmHyXWfQ3ckMflpHCvnBE0UL67H1
ON6VRD7DU9im2vQsDBHfWj2jh3xuo7WRSJjauQg7QdnIcJ5ALS9HumFb/x0dwDOzE3PDf7IP/vGb
KFIVJb6ZrFdKlF4ySrGNeOc/4/zTlaUzsDa9br5Sjba6leILxVBJd9juTx+4bvxdGNCHq229L7kg
KUHm75eLCQ3dwIXerIbEChu/XhkymAAiFtSiic4mbBWqlpcJ+SEI5dP23cMgkwZukZykj/G2zR0b
xxQprErskFtkykTx6aPf9/G5bOm49CMI9flqUqiVXx5e5Lzql8u1MgLoKrmKWXWGTJeex+asqx1H
33IqnXVLeip8qhQZzAEFQw3s9lbKfSItZf2w6b2hKsgaw04Pe/YRb2fKr/G2C61k1EKaB7zopmtV
bpmtScja4fjF7JFTOdYP1St3RMJNUQ8HRTJzKUh1MKgC9KlAwsDfs0mPWtpDb08b93htX0US8Va8
UmhftlkoAh66/6lJF6J3r77/8IXFpZmsdq3MDcarLQORvNY3FJ3XDgEYEABGtBdD0wUKI/LIqrM+
eBSS5s+Obo9uXgeQ9TIcNmSDBgFXf0r9art4vSCektesgWIvD2J5LabMfk5gdXxEvfsx/ayFxYJB
B8gn9BnZW/Dh4tiDE/2duF+3fJWe1TUVW9+bCWL/7qi5oA25dQXlv/42RxkYb2qNqmfdfULMQaDi
BLIqs4ZTU29lSZp2/9E8A0i9sJshI0atWBgsEgpRIaF+nv9OJyzXfljKt1nHZ5/wxFyhWyymT78p
TNkgCDAP4lgMt3VCej0zV/17wN25QeliWWxHfX9ZJUkyeJVE6mmJ59dU1vb1fMRiwCJe5pwNjjFB
FZYwIfw2l7u1RBsQT79r41QsUEG7UGC+DEuIEE/wVepjchTsFiNkAkcR/izI8KGDTDZF2QzQMGSa
7osF61IQDXRstur/S1PM5Oe6bg/ZV9mNXGMClJnIpCCvuk77ckagNYpiNweQjQIpgPvW1T8MOTBl
qOrTiNij+H350dxlQegXYWd4uAqeP6Dtwo7z2Ti9dc0coWdGMWMlLOWmPmXQ77UIkO+Hacj4Hqzd
IyLolHuGq8oftRWQZ3cLZu0koOjlhZSySZwcUAXjEztcVQmPj7dASvGcYm10k6mJq2kl5e+kJAaZ
z5zGCBo8Ji6pCokXM2mLkIzgDcg9kUTj0cT2KKg/zTjGboVZ9ylBR/upS6WkSB5AU4q84ifPWZUm
xbODtd3XphMmS6klE7bW16SSbyToZaN0JPVClTiCmcU5Aq+BbcOB7vfIXq2T2ddCmPjqqZo2CDvd
3feTSrhOF0sECs8sbbbx14u+bbodFwpKsv/KX1r6nA52aJzmowTBFfaA04rFBGltGmYjWR+zB3a+
RkQjhbDLLnmTOAU52YzwI+L6RJzAKcw7DOuTUIxJa7DmC/z0bH/yf2mrv8yhYXMgXoFI4/ZWM5eO
++q3eA6itks8Sn2SPj5C6N9ycpCu85Dy/5TMj023v8R6YoboAUrjnY+DK0ld6DD3TMGCFLyC1w+L
sUunSXNe/W3TXv3iDjeg8Pw4MAjzYtj1g/sf9iI3I9m6m9QBczPcM5OkatXMzhINKICiZVkyEQsH
NjvacvxJcoSaVoufOKiEM4GA02QTn3LOLcFzC/bWEh+Pra27BOU1Z8WmmZdZAIt8l/bleupmGjQ2
tuIgyxCBDGdiMx6h9OyC2GIZ9wQCTm1r8k+9M1F9Ke6Jy4u9yXROYWAkpw2s4C1ZKnDN96lu9jX4
TcyBFnXUIghnBDVzmNLeLyN5qbYWxICk30KmNyMNGnnrjZvSrqBS6dnPSkTFsNDW4h6gUpGfe/aY
osDUydKFSc+8pmCp9lDQ/DcIgimgzxwrXUmg21CJtTI2I7icBgxoc0rAkNu1evipmit05xJ6aYEP
KuqhB19ZCY9mdkH4FJcW966Y9kzmW0ffOcbq/FfI6SToBm0HTUXlYOZAv0JFU2VcjVpEnzjt52x1
4gonODKQCF0XZ/QoOt+j03nu99twuXNi1nryZwVmdRXrmI2cVVlwKPnNrdLN+X303ajNF7qCwul7
epaQaMer1QrGehLydygGB0MN9+JZRuP9CIqBrFPLdIAHySXwZXEbTgH75xvdYHzIoSha2q1zZ7XS
4ITl7cpZf0xoLxJdJPmja0yr364y7ldcmu3DGYzk5YhGjTKt2n36Eyuas57lZ3QSzhVUROWcf6hP
o29zPwo97mss5vhib8UQ3SazHE7o3Ej4/2Bb4DorqbQ7s1eH/4QP4sBuKb44I58qB0b3bPjoiYsp
JtrFAV/SkmmRstNCpJp0TFvBTreyqyBLAWNkqs1dFkx88ACzK6mOgoIv39d5Oi/q0Su+Su9oM7Kn
uiId6No615OVYbZf0ksjMgLm1NarGbi3A0iVVPzb88e3Zd9gDGGBDuS37LwaPHQoeO8ypVeNpokY
FAsH4NXoV5YrKzIpZkLDeBaHzY9NNjDmF92LXW88Lb4v0oSWzL+2WfOQ5qdMKc1NhaKhcjAK3Fv1
Ti1dZCVITHHWR6i9DjQC+fP0VN0HSh4Lx/ZNieztfBvUJ1sNM0ahunjc/xo4bvaMANJHcSkX3gMP
hlJzaq0dtQyN0qMmkEJo0GZfGBENs9RqXCR5fkRkt+0KcBqcLvs9TxFToP6hDElz95t8ANZtrnNM
CQBcOodd4fQe7tqwrsf8U5k3CpEN5Fz7WlCwzD2fiSnciE5YvN373ADYfcLM9xcvkoizHwe925Nx
LbyzkVcbrxJ/GJlFaW0Qg0sPZXJus81Ct66eilceHLhHodYuju+B9fAP2hCvwUv0e/Mc+A+T1dOi
vlxcSIP2ZxDkVqRS+5JE26cCJdWxEOK73X2GkPSYPXMur/2XwZMprnlFpBmZqKkVsPIF42Dh7nS/
qqHxO84imtOKhE92YYKEGIEXHHeGQvWQ4qjW80umGV7QB7MQN82n+pLKJ0FAG89yCuoo0yr+Dkb2
xl00L1PwUvS+cJ/xFc7u13X3tzxpFmNRk5vxEmPDPX0hrsPrI9g3nbVLp6dAKRDs2ppJzJ5U/6de
f8D4vHBVtkBh22NFvqdTcJUAHdf28SW++RsblCtFpPpGnuIP1u78EBR1aBVX2fSPJPp/dfaSltNV
7Q9JExLAPxeeyu88G/TbeuRP7Oc4thRBCo6zmS22hCModleuy6GLUF9MmHoxlC273Lz5EzJjlxf4
b/4R5sfVTdV5FnVcHySrnZPpu5XClpiZ4Yqo6Zkv8DD7yYYvmD7uKl7cQTv6MStT0DQFBIVeDZpQ
FRCkNdN06dD1AkPi0X1eTPdcKy6iT9AKckBrXbw0TUtB22xrsQOEnmOeCL4biJdGB92RSSxuV4Rk
yt+zdTU6C5Og/fWdTaRz3E4EH2EcRcmiLTy/0ZEabIMOWxeul4eseMD6nTDiNo55GPrKCvcuDIDE
HCOk4zgLnkkEUg62UtoTLS2BLyjMqGLTOUmWVvS5qOc5rXq013AiQJKAeaGD7T6uesk7Jxv70phv
mRETZS9oTcOrm29ZzSn+RIGC8Abe/L/xCcYRM+mRDkr8vX7SEcL8qlH+M8wfzxWUot9h8YmCtGgD
WvjwNb/V6pEt0zT9H0ri79c/ro4pN/pFSe+0f3m+/TDgWwlvNTCK8jF1dZGWQvLnT/0IAeAO2TZQ
G7JgJIfnlMzNFFgCymecwk82vvwXTlmyJQrujPrHWFPRuLCjBImYdLdhxuNuDlS8de6qXBLZAlvH
MdD1VQkh5C1E0A/do5+u+iAgwY+0c5MYnT6iRSi5I1dfzv2rta94NTZtcJFL1Ecj85ZkfcRbc2p8
RfS2V6GyRgPpIjDC3Tz+4ez0oX5YW+DPIKXsKMUr7djWLG0Ec83F/Uh4SyPl960t8K8lsoVWXys5
sI3edM5fGrGQAhA7iOK5AUA4gHy7nGtk9K/HyJotKA5i7VZOTJSWOEw5m4JJoxN3PD1sMopL1Qxa
P0WHEbXriPvSp+jLnvYo4VrUFqHC2SSPty1/lTCV42MX+YPuJvtDLsSAGTAE4pdJ0ITRs8C5E2q4
P7U0XzV8yASBFoiQ4WFjm4FFlMq5pCjgorurPuag1Nn4LknLqMGqiKKi6L3d4ia8rPQCAmbO+/gz
h+hAz0jQXuIpI9cUaRsOpIQEnv0gxXbWgX9nvu8q8q2e8L7xfJt30lbTAtgu1/uUro+iSUEa1vBN
a58OqGxdoL0vFEkAlpxZX+Nhh1q7AOa4V2zKPUPK28MKDrxSs1fS0P3HBejiQIqexY7wd5VrHQmc
LSDbbfkl/uumC0G2K4TLkfc4thnPE9LO3iFu1gdLrAfF79LiY/5zNMdU9o5SK8nRYd5kGy/+pS2T
tvt2c8qrP0JXUGmzDzIJ2912HYyiMOAQ2YUsZX8nVk1OpelFl3SpoP9pqMYFnaiJRfUhSP85aRKk
+RjHYKjIAvBINMXXlZU6Fju0zMQsk8ZbbvuReyOdebjQlKHi2a4WrHzOqivxbRLB7bIc89RpbQmA
ACii09bWi96n26RsCFKQa5NyBAcNapDukoi/1YwW4+ZNtKS61pkTcx6svGJYaeYkZVJAsHoGRJRs
Ti0CnLxeMUBRd2/XgODbULHfiBVDJc5S6dKxxXqqLYQlnEPc2y0cQmloSKo23NrjsKER/9qnnjkH
gK9t4ydqnJeL0B7CnvfFxH3vzf2woTB9bVBTDB/PzG9PLcnGpr3kEG3DYg1ChH4uKVx1FcGG3czY
knZVwfMX/3lDdfLBn733a6FPMBpT8Fqey3mhj6AOTV6lE4w6ggG2vFgBmyUhi1eUFgDCTPdLys4C
E/qUIQbpXfPgSJ27IQXExMXk/ixmQMxxZ2hlq8SMlkmRKcJMcYpajn2Aei27V+Q5gFpGmodGu0BL
mnYlh97yvbxwBowbV99c7SNRhbYw4OXkP5v8ath8W9lDxKjffGrJl/RyQ/osf7y/tUk/VT4+EEiy
KR8wwIISmiDpXXnfT+XmL+8ETt3hVfGMPOHTxR5iUkScOqOU1tlznlaACPof70fINaqknnFWkgvX
iuTREkQR7DnhdjbOzWyMSUT572ZBsQffLQx3V17WaTTdfVA/go5+eBkv+wYNeNTrSvfdklq48VYi
igJUjNRp7/4E7HOt3T/8hRYvV7S9j+a45d2qq2+b7Nk301myIB5we35QkShZrRdbuAMD8q81hL96
Lmecv9aW0hnLgc//iZyIazWTV2N1h802E8qkHcFd+A7tPYzsNmL06eTT1nmkRVyjNnR/kj5J++D5
t44QPNRULSlj6lznFt9+yE9aT1o/lqHDK428mRjoFhKkJ/0h5iRI4GKS6B45TK6o4T38xYkkHj8E
/gJj+XfUw5a2Az/wt4qyr/bxKWCGUlkUMickbxmTSvr7LzSwRkey/fYjCpitxRswJ+yFdlqDOYj5
HWqYRkATIOmgmdMkAeVJaMk99vCRYHCYaKZ2HxOn3yjFK4u8XzQiK4BjPPKA6HlpSwmDO/tw2Zwa
AuWR62DOduK3uaP9rozSRHht9ZYbum4YRmo31uYP/Lon041c10JlxOHz2W8QwFpPL7a0hBjrWw3m
PEfybjVNEYgX5LM2O1eSjyNAehO5rC2NwO+Ag7nWY0m6Q6rwdXBv7S02O8dUygArrvPsHqrz7qIr
KX6wDdPtRdakWgPvEwv0ThJ1k4OtzGDpA0PfCt+uHKWRiIpMORbUAM/ptHQEKydy5wY6AhTvK3ex
D43Yp25DCTyBkPgpOQwahGYezIWpPoBrkKxaDGFmfAjL+0SAXGrokbwZ/7A2EjtAMn2/RGXT9u0/
vqHzUQkQa2mdZUucUrTTfoutBxmV7NcPSO/LhQIQkZIpadINHXuqyKCBrJacCGsemnfj+5EaQozT
4C1wzkh3TulzrI66NOigMShWUR7NmwdVf/Rp6JSztGdThrm7SWlfhpRZP3cpkvJlVg2XP0fhwGCx
HDsTWEwYeM5oUnEUO9Yt0/07TVonJJA4QZ4PcGwZtBAqohQTwqnKF+5EJ64o74030Jq7FamhHffY
X7mSjVQ/ATGrixlu4Gb4NBr7du6Cy/8D7KmI0QjLrqcSyl15SZ9K3JBZMHrRheK8BBgSdzyRpbzv
jjkxB3C7PjZn1r5uxIbRtANLybtw71Jb5uP9UwIF6MyNDxg5f08zVjif+fMJ77T52RpGw8EpEkqk
WVCe3j+uNTfbqsyYEAuTAnUuOZxIqly89P5COmKHax80OXDlPyotQAZrz2tzWnhxU0b0rfZ9bVmh
O/Ch9Mm8K7Cgva+x143OWz8emGYexfFqSYmkkkI8QWlFA4mBioTglbJpbiivgsbiJT/wNxOHpZ/a
+FIKv/Np6GB/vGtMKrXHWLh8agoQEYdKO3IxoH/5O0fW5zX7ymH8R06u/4356FccyoffUfYN7zuS
ZaU98LlgdsYMxzayb+W1ARc61Kzqo0W4VWIvtI6SXFoqLjhDVnKF9d2uCAT+1WTtWtliDt+DuF0I
cGGCOT+Kn2UZL9KjjxDah8sSlGy7OTlrO25rE5ZLT5Mh3SAM//dzgPsuWnlS3vJz8Nqxm1SBQpiJ
j4qdb/9NXVFSnzMMogz1/W8eljonCGvTzdxms5GUEahRL9t8ZR8y1rqkNk3qo/itJoNQiWBKBCYM
/o2K49hbAJp0TIYSK3q/uYuqjL1qKyHcWovdLaAFGahVwJ5bcTjDo4OptvmdUhTQYQP76Yd3lAR4
e6Z3NsfZye+44pPDb9rWmwXdgmwLyLRDLfkzVBPyy3JmSkNuyQcKIeOrwmJOjyv5EkAjgQgbk0ZG
BOVxb9mVcVCrshKBwtvd8tfGLnDUqy6k5pjk1T40dZSnbIRggKTUoDoCpouT9wycyXzTkjAXgJI8
5QX2z9TZbBOYlrGGfkx91rL56otIzACDP3L8xlhPHYHLAUrTofxYSdAtEoCrRP5m39E6OrNbdWqJ
bNq4saRNl99j0wtFGiikHE+OdIOxK53cJhO8EWZwLkz+n8en4Y5qhvQQ8HBXtDhnM7rzaZ92qvWd
cXFJ/i2XIrODs3JxuzzZmx8tP827B2bqIhoKCs5G37ZJQqllFsWEKhvdO3JYqVNMhSZ9d7S+r6cm
skzSX7an6H4A2PdkHK8VNKF02jsDPUE5WNyk03XURjRr3BlrT8ZwunkJviCAh3RRl/7Mhn5fxFAK
qFhzU+x8q2Y8W3BZl5GZsKS+q16k7BvnXDQUPgkkj0cnpdMbhR8C81T2uxSYb1d+8z7bwSwt7o8s
XRaL9Lb+SN2HITvIcqWPc3fJVp37ZveW+FvQFnBfiz4Kep+vO8tJoyZawUE1QskD8RysQVHD9GCg
tfyyC7Vh3asA4Ct8Dd/mkuyIT7LMs4dl6dVH+GYvOfjPhZlyorPPOiBDNacaPobSWmC+4WvCB0iX
j17t++Zi4VtIzfry32+xFqSgdYnpm24rRG10OvSzn3DQ1YmIbeSiVLy7BJBY4xxu6naRGbjS1qHD
d3yO58yv5VfS0OUmdwsjqhG6F6QDMr3eMjVOMIrsiEBTwMVWuok5vp2ZfykfHmpEL2Z3MlieEg9+
K/2RIKP2iMwI0vfHIzmdNQe79XebqJnifFCMgc4lDe8ap1tUOEDUxbS18+mFNSwYggQ3GRV4LbZn
yB+ZB1ADcgRx5MnLGPwk2o1z4YkMq/qUsbh9DecwV486I9Bf/2Of6kfHGtUOxhdLpfJ5sdb98rIM
eHWVcJLS/zXhZHT2+eZwCOuzpWpBbqXt4cnTZuwiRuprALwY244gmoqbFRy2GyYcKiII5MytecUk
xgmSiORYICHgWZlyDoXpN4z0asVQe4q0f14f7uwUzX7rZyqjLFITOs2YgS+N8YLGzruxTLd+NIJQ
KekV93HzGkGlUfh5sGgDrFjaSH2soiChPOLJ6oQTabq5JWMDF17CZ8xBZKTblYQaMT8hW2+DPelF
f7yPSzuKPplNpV7n0yiHxGrufKGvgXkJn+Gq/EJxhyxcf0eZmKOAk/KChNOlFRh8pK9htsqNwL8g
Da2/EHpONOszHFX3h58YDWgGkM+8MlrlClEnai2j+DFLwiPeUvRGh52esUucjKmMDD3bS5IXcmRi
lwqFbR8MvIF6zVPtLQhpIzju+ZSCPkKpm9C6e4rrJdaIGnszXdDc3jkbqJ3etfvcVBi46txjQush
gHeej3KC1cvZape9hU+7C+1qR4h+r2N1WAdZ69FkDB5NiGWunYfH+p+LWBCpYDlewTbh69lJO4yl
HmLw4UEjVvpm1bEw0sw4RWDQDq79iYH0biwWczwHeoMtdehmMjzMZ+up0yOnvGPPTm3TlyUspL/e
Lbtsey44iRA29csKy5O5iLqw/gv2qJH1XcOgsIJcgMsuWrTnLXMtDRqfNeeaa3bFHujrm8zgrJrC
HMVKfbs3FrL8TfA81ZDZ3RHGSKfqQBd4CueC17PRvxpDt/Fv51M5RRmaj3GKjJ1W4mH1sSFBfaai
sPw00YKkVAB74qbIdJg1aa4t0yJiSVxyfIx0tyI4WTsN7W2NRj5RIya6xl1NfMUMBsqnJEfKc1Na
sUJPpcS0UvrHJ0jp0PJilkuMeEVx2nwl1sW1Z1uUMhKhlANJd4xcfQ35Fqr1M/YYNGO36ISb2auh
EZJ8SBFvXpxXoh6HSy35Y4UJCwDOlyojSGJICi2fjOR8dKB/gR0/IEoenXZIyIuQEGg/aAl62Z5t
yFvk+jrv7ExCGQnz1GzK/pIm1eCi61UFF3WDcpXU/vuIbT/sZBl7WhaaELQ/BvFjp5NaYglEkq4b
WzHRd4ot8Z8Qvr7rTNSV4GwowwporAJq1okUC2NZsMtFpY9XukQeyUsJKuYrRki04LADdekHmbAC
GqOfKL7te3p8SaVEkekAKZ7U2AeYKWLmRpWGIrxklHJdBDa1ZdeVWNloFtOGDTQxgS/3FE/EpD2E
Lvv755TJb1OKn+jtkl+AvV9HKUWoy8+y9n0k/H04rbDgaSw/lHpUfYuuaTEQ9/K2b7tTJQHq6XOs
4z6BWF7prYxkZ0C+QVcNSKOlcTaS7xRnW6rjO1dh4jVz07XMJvdsvO/PmkJO0A7D+f8pUW7tENOZ
5ZR3+uDyDJmcXpduux/Hn/MKRSO+C9zQg5dGpf8BRtCjSWasWD4z3ebp/Uz38c5Pa2Of9wLHK2w+
J0pWXNSRJ++B3AnZ2zTSUljXWYdJ4+X5M35tA4GbYabS3GNo49uwO9xXZHDk5GTDxgFG+iVP7zPV
Iz/3YjE2OV46ghr9g4pvDrWK2I22+djvJD4X9wkE8WYcfe3b2GU4fxCV2usIO401lZrJyioPiF27
/NSfXFVI3BVOXmXTs1fsf4kB4cdwhfkNOH6YMXzB66PvBQ9FegF9/9kDMfgw6yTw2249MMNEMUq8
sS3XiAe+CQ+w9oDRvj4t13Kcvy2QDwLoeEkQaMYd8FKDpjBHfmUb+hDmEvFq7yS/anbOSWdRK8v0
s9dKQ3KARhaCzuXIUBbBfOxMWB9xISpS1LfLo6oH7S6sn1PR0H4WYBz3SsoFF+sHR4OoyTCPe5g9
1kzUIjx8p3PqUnWXchSlJ/SgV2eA2stQBp2S+v/Y2ZSnu67nbE6YBVvv3kUscjagf/2p7k6uRIXI
bEB9FSW3dXWYCjN7zLwD9jP5iwJZU/YP8CD1C5bGVegYarznvvOJnu5tVmY5wFEpCMW+i/vuHNR4
MyOVWJquBk6MX0SUrewpFVsOcFZoWSWqYXi2EKzoAv9wYwT44U9P2NWKo8Aynduth21EraU9hM2D
ttL8n0uynvAIBQIAGTyG9a5RG1WO+GGzvRvJFA5FJgLAXumnVKr0OOv2ZQ/PK/y/UZ7xMaYVQ++k
rSeuZNPTW0LTI56C0JTofoZCLO1c3pp2b+r/c7vNBd3IamDTYNztT8+uLKtqNuzPUpEpvSXWPU5I
aPS76XVmmO6mkpL1UeWgdcJnbeBC1G3P7cajvzf/TtnXPf6UsxzxgnmywVxiklt1+VPbPYGkkXaj
yefFA+dqaqdIUxJHI/iZgisGllX3F4cuBwITVxczi3fLFQlBNf2gzX41ogtMSn6ICOIkOtztP82K
DM68SR1ah/iOerNCDlLfPnKidW7ukHnLZWQ3vPNg3o/K7yJNXapaoDHcbirRCpieq7xVxviC/VA7
AC5MxjYhWOmRWgX7QRQf+GKc+4NTxdKDi/tZb1gE1X7fKpozxVZ2pm4V5hNRx+HnkZKjVe0SUZln
nSSigTl3LdcNlELtq3G0fURfQTQa7cQbN8aEHc1Zs8LnVFV7QsRy4ifXBprTdeVRIu0dM3qKPOnC
HnfE2LJNqrK8fv1UWGaYfVpCWhTnvOC7gkXow2MOejop9deGDxBL2qymn6rGkGi3HOcLCKiGHiDQ
SI0rsreZaPwVvZHxbaSEVjySJMN/gVYY4yKjzKbXGwGAZ0BiWVF7N3YHtdDIwCDQOrTEvdXQzmpA
2wIpWygM8/D8noTi1j0qGQUBEC0lHF5q82iWcgcEV7Pi33uuH9jGcs60QDb4NRVMv8zBCQijaXuY
M+uTB3T1u4L4zbHBe2cUtEwMFxv6uX2m4wMtqyfNGS12k7CmpaBgch+dm8q4enJ0bzOEA+8h3YOQ
uL7rXh88/nrnff8iJG8rXmsye9Cn81qclTazw/QmLOQfKZxJgQfBPF6n+u8R+pVgXuT5m7ARynlo
FUsypIHryax+MC/IiedCOSuUXBxLwpbQJNRtsOv/SHPgstIl2uZo8/q2s37cEC7eA2GNt5LJZ3QF
Wp0sf0zzCNk3isKP3IwEoQqRa20AKW9FtmC0M+R3YNjZ8xFTFpUuus0LyipfNRFnqqN1IfU2C2OO
DsDyMn9IVzlCS/S80K8s2fDowTyWaWIXDIAX1ZgLZxi8OWXII05utjrWDWP8IC8cJzPjbP76Qb36
ofT1L8YqI1rQAMbp1xN2Qw2oOB9wRKU+9jf+u6RA6ALfJ1cbafnYaKpZX03iJeBfc0WDzJ78aiJG
RwM9mW4N5CDo6I09XFl7d8xPrYHxqwGUemj3qfoSWz3YzyCMKGD4XD6ZOW+w+snjhM1N8fTQwH+4
k2RBgZpim75KZgLWMp/OUpwGpC3ad1JuJ604E7lEpov4+Ac+vInkqWIrgHI3EzH9gjV8nDUyC4Bc
G9ridk0pUzU/AkKIx9mNBbak0u+irY4noC+g9t//FAYsYjKEsgNZ6QJp06SfxNb33VRRYQJdNlMu
TrYq9dceN8UPBbeWyNE4aIFwkOQKmgri40sLlY72KThW5+jSwMFbEMihpfiEpi9Hidx8DCyHNb4y
zhfdG8hy+XkpZeohVnKqGv02Wy9nRwlcfrzp6h5jALaBDFg0DoIAs6N6krY24QHKPffh6u5vNUrm
paDpzVDlQ7uy5q3dwWn6RLsfWcOX+iMASK0qSwcc9xvevHNFGmCUt/IcOwPsJcialMqx7DWt/GHS
zfSPJB2zgTbi2MzJ19s8K3yzauA1N2HSwZHSJuJ4KEXoOSA20chjiAQcZHJ7Roujo6I9eeLmXthz
9QuesLjgPwuvDweCKQLI80S9JvQA+M0DbT0DpywC1cAZbio1L6h9+tK9MwUH9/+XVbz05/7qpNXm
AzWnDzpZ7Nl2zduYpDtmjFX7ZCryOf8CrZrVjFbdTt8xEqNy6yH83dlqokjzkG2LTWhmzTQuTaUt
ex7yzuv+Uw/Mbar9gLFQAJioLUl2bvec5XdyP532LHR9xggBl/cma6GZeckg2NYkiqG5rI0mUil0
hvyHfsmiL6FiodFeieNBH+ju4fckcYll/Nox6RVDko8rRQXYOdZFUkRzWEgnxt3Se100A0MdeIbm
A/T9HpWQUjP19x7y6UZkgpnopizIGzfMv61y2dhsRsM3Kqsp7t5cLS85DTHt8d1dRFu2j4pKLRbW
M9068KdIqRYiHVuqBt2AavQimg725wHVQGbY2elevL4oVTB6eq9u6NqZjfkfesYfdZIFrh3oWZhG
72KLXu89hwd1J+anKlGuggEGaVOKmRAIcHp49eJrTcJEKf1dIJ2v3S4VVWlGmgqJ4h2+WYhh5Q/0
JdLJhQnqphj+k5ADFhwLtGG//3DtTAYAXR439SV6yWhS7xQu5SR+c8IigLhFlECYAQbvOe+bPlxY
uhilSVM9jGnCqLHaM4KOBl2tz366lbSIbxC4IbdF5F0EGkc5XPMKITKNSx9Y1/Im+yxDQVEgrxjS
aptK+lt55kEP8zn06odsl9744tfWjXf3XlS9aIy/7eY7WJ9NHwfoH9WpJU9pIWw1b4fopPRv81mi
4M1AcTVZK+uYTWSAkqGczUkJk5m2L2wrED1gyVqdZ0PicEg/RbKMsE2Tphy/NlcaqSAAw72yhlsG
0QltOwXO1+jy6pMLVG+EEVimWPTOYOT+NCubTG05OL1qaz1CvPhJdTauDD9Fc8hJmkutpQhufxgj
9zscTUQ/PUawVC/b3KbFAhAqB5v5JrECV9MEm/n7n1LbDBE64/3mMdBReNqJI/Tj00XNWx4C/1hK
xiDQOMPx3OAXeSww6p22JGgjQwiiGjjbGcjGb5bD5o/qtWvkCX1aYiHU1FdzSI5hSJxCYAB3t/av
vzXVn5o0rRx8hZJNhDTm54QCe7O0NHjnvut1YIMCLSNB0xEDiLfVVcH7Ma2xIq0jD/9A1aYLoHpu
fGMBvPYvCgzgX3UEJQG3y4IwF8yU7x4jlVozNrf8SEL+C/yJI7EY0dJGjv/xUW/oR87RH3bQFvHP
y+Ja6rMd/RVxwtZw5iHqeqj3plGjAvBeUdYsWq+ShhqHJGghvjg+IwGSDQToHlAYksc1wFPq1lbb
j/xDuSTDH+MmsCB4v5vi6312w0CRtmsbpE9fwnXpPFrzHLuVIz8466tjw8CmsUY5ZFZ+zfvdSlAt
UZkFu6r8Qum+q8uUVqypRugr3NCB+qvpWo71IQw+adkGTEwg3BlVxWMVtBWxpemsc3Cz3yCphmJb
DSbK2Vs5zE79+sumCWubZRfPwVWLvtS+15ptPgbYSxAxOUwWbgt5RIPX5n6Nd5NGwdMCG6u+vSaF
9KmpTwR2/QmWphkz5la8IX74eMbixWaT+vNhF7cZerhebLVz8cu4DmQdwdBCAnUit7fR9Mw9yg+d
kIudA2x0uBez06QoELR8d+Cv/wL2u6X4NhYRuW+5ZM9UiB5B3HUu8aIhYNmigkLOvVZWBrNPqm9r
EXK91KumpMDOhlcpQkua5zAa9YR3BvvjQKrb3Yc2r41m9j24FIswaYJaA+MQimLNvpQlasRTz1ID
3oyJ4oMah0GHoAvqNvmHi1H8VIyCCgpBc+9/SIcPbfwl0+HubdQQjqbmaFs8YkmvB2sS0B4MpsJf
HXXpeZ4xV1uCnsX2Dhj7DPeOlF32qbu/YejmHMUjOr6PnqrRph797maHFJ521b/qf8+Uhw4GYl2r
y0xGoz2pxGTCGOROIA3V4D2h0K/ut/Kg7cS4GjNpmLCwK4Q3yXURoztpzQw7it7qveShcpeO57y6
KsMdbK4uoFG19xWFes+7D6jLNM6vJ5O5a1fSyWAlhMJIAYz7uJ3CVu6USQoor8FaNaq0h7vW1BcM
xTeyInlikeewIdsKhayxUWe59jWrXwBbNkZ5rokPdaZ8fr98B4/msAdu4pcXq9ABtnRPfwaGb0xz
yLGwk3Qk1quOYevYtvWoazWb3m3sL51GG8O2IJhazNG5G3ZZfrEEb55UESiQs5/E4onjk8c2QTE/
PjJwE2u0vZbZWj4zc/f0myfrl3aBSXsIulkTt6UQzC561CFjlRMKVPGMRggc9D2/fq6TGzeM0CA8
FDhprpRic1twMmEJytBlmMhzkv8sOO3kU+c1NR6HqoYn7+p/qJb9gbgzRqbCyGxW2WV+fpiYIMgw
oNMfV0p0Ruj0n6ACenbmbUm8hOlrY7Dpn+pkx578ElemZunx0bnloBrN3MeMlTv58e103tu6eLBE
5s5FD2/MmLCegcnmTd790wTF+IdlHGpLFICx4LA7lLulmxag/gCpLjiLvdHVT7IEfJVQ7a/jFWVN
sZz+wymkmZA6lar/4edx0wixR84LQZcnMJgWU2zQRk63mkNPn8PzOFYIBZN7yqe97lbgkdfBtZm2
bDXmL2bKGWflceufyGRak5eFrQx4xxx3oTCyeMJH99C8jrW2yxQXKOZBEP22lG/ud22tfIwqXPsA
XsohUMJdC03fOtx593a5OXDMJi72IVQCBgmS5hJwAPL5XcRmbLVD/9yCq68UU1ZkSNWitYMq8XuW
oWiIjtjUSGAIxLkZDv+a70qPRSXpbDELZvwFNjAvDBQHHy6sUKFdefeuPv5ks7Gi0zfhx7OPN8mU
LeEax+c5tCccUSVUBK4wVg10ph6nBA1uKKyvqB1wDwaDpMgEhTwFveHbfRUrjHPN5EKtB+H8AEQZ
V1AiroI47rxpFZTry4Qf+shPjZ2jTMziZxWt7Klli6J8nCzHuN5LassiMwsgO2Nzr4pZQG0T4YG3
RNbGRRiogzXt6zT/ERSQjJCciSs+VW/zD+GT5Hxt6craouj7h0+O6assoD229eyU+o15LePyZU/Z
eMGe58YG6FirQoRHHUB0tvEItKgPayJ6dsTcLO8e0ClUvpejXI2mZu0wzcYWAo568WqBB04rVTE6
4Krl5B8K5c0rbCwhCX3YeYN7CgTYcFdE8Pi77jbGvwjPJe2ayxVFxidR/t1Mbb3z892Es5DdvAiK
iVdSd2Ubf1fh4hZhFZT2RWDzBanV+Tc8PC49VdbdFxyTch0xsCK+PpkdZiEY72oYrNu8LvgKujz5
CHV9RNoG6p3h3mnM/En6707BbirdQVx/rg/XyvtwEzmD9gj0yj3NdGbuSpNGHaHWUlKBdLn02WA1
LRbmBhVhNhc++eoDmWUD8gOGXSaDg8LoWds9SBGP0b8nwERVwlRYgYniIXaarApMfDgizS1QKFTm
LFKaWBtKTZmFbH46CTjUe9NL3iQWr2+sHeuWEyrHbtXO1Zz5Ed5aK+TFSZKZk1QnO/VOQ3N/ez5g
1OOOo+hhYaQBLwnUiXlXLxlWggNFxjKxr+gGbDYspTqv6U+dcbmf5aW0kl4hNS5nC1A8/y0BUPhv
/mUioIhFCUDYgXZIfn7RSdFQ8X9A85zkw6LteFHGD1e2tknplNxhF9tp7Nd92VrPimb4o4qdL/Th
tiX84iS56yawQ9bw4qd550IQXLf384o0ya5JrHrBvoVEMcOF4suC0EUgSjWHA9U0/QUR0kHlaQqx
BrXjiS6XzXbhO4mtNM1Znzv5bGs5dOqeBEI1B/AAlpdpVas7HAsWP9vmYCjAd9X1dmQYdy1gT2b8
o0CcaQad85o6UVVuRF24VGoRPI/f5E756GTh9mISOVbeIH3rIAjhfPNus6GbZ1Dinql4W6tPipdt
apI/7cH1rhxueBGll6O0P2jIo13LR0BQRlNsWsuh74Lm52LsZ/fFi3jEXH5+Hy060Dxy4XSNQ8Tw
77cYNIwtnGoMO8Zunoexa6OmibKIc45ruNZDGoAWNFr7CALaQfk9d+kN7fBy21KhathfV82zxm5M
MVdq4IxKNyMFKwXCfBVWi7R03VHhKBQP34dWibHO98CPUtOT0Pl4uBTz98SX+xH8EeB2NG1MiCZb
KMIaTk9R8JXtG32B7cjVSjR+WOWmYgPNJdbor34GNbg7GhVFQI3F2TGpH9z5HKJZIAvQOBr8an8r
X4km/v+Pw+ITEKw/6Invj1SUHrUCHAIe6u9I0icP/FncUGBW70w12JlRSF3Fzk+K7Y2xtO1NYfZN
XuiNGzxsNZD0x+KxO5qkl65md4bIDX3NtVYBUKl4dr50qT9Js9udxwOMdj0xhIDwmiwkIeXpwgt4
DRumhv7rd+SUaUVjYjscojIG6w7bbzlc6LeJmgE87e598k4QYPc9AXM/BsEbJyY66KMxiVv+oDbW
yeyaSQP/wB9Zc5qqNJCJR9gIpfPMtg+7tcl0hjvPdrIttJyErAEjAcI8Q2hp/acFKp83UbDCHkD1
ChfiJmRe9iffCyJmBquzXzLnphYJG4z8/XgL+7X8O7buxMYmqdQxkIz/dXFEYyuoxOxHVGig/+lr
/p7LPj0AXZzCv8oBJy9IO9GaHCaUSU2jKoXXgfI7Byv/Z/hHwQSd+ZZhKZNiCvtItlVHg+XsYmk/
kdY0y5QSq5O1BsSIB8OSRqEuabydaiMOlWomH7PIyLgpAKjQ/PdWaVCWG8W0iq79RJWG6GFxj13O
n7C9qyFhqKOgTRKnOQkRP9OxQhy0MH7UZXFCd5IWtiha/25moE26Sfvz+BAdrbFtFgYCw8AdjXHC
XGVy4BWDO0gSVSMKUHiCSF88lskxNn9YckXmjQp3/5795N257SkO3jQqqzZAv/6Du2pPINmBY/g/
2gn0wd5Dq44mgxY4oe2b1Pg4gHYpfatbkHpBGVifb/1UlemaUHyBk0GAVj7IlSmyJCDqAoNtLaBG
EyE/nyL1TaeRt5JfaLe2P/7qnF2aSqCRLc9aqIt8ih9OKVPi6z7tRHlJaqWadvCN189+EZTrQE27
oy8ZPzAI+/4l/WfGF0enNHwgiblJRTVUQB4vksUUY0izWdo5p+bLycYu3uzyCOwvTGzCaKHPjmZW
L3jKoFjydiAXKXZzrOIF2vjNG4+bc4eWm160JEOd4SjDfOol9uIgmx3INrzBltN6HYfZTXB0agHy
/yBEuySaRgEx4MZoTkR/DS5bus8f2JpW/rqTGjQMF9u6heNwHXiRK+lrOn+hAJwhhVbAFbAYnaod
OWT5Gbpppkex3RENgGWQ9R8DSNtPW7n9eKeH2rxOJ7Bx47lGqnfHzjhfdoMdvoIZcfUVDQXVscXO
nL1cRJluQQkoaG+O4e9yloWg02p5G66XiLdU8ufgcrHSB3A7smGRHJC2qz4SRl2Na+FLLpiXmlAk
8Dva1h+SV4ki9C6S2ddTYXlxKNS69gOp2QP+IDsnDG2peVGC7bQRmlaS0ko1DQfJ8+9MjeuN3Qfx
DMsMx5Zr7fZ3m6+AotAaveY3Q2EBd5vYcqoQnyWuyLmw3tKwcwR+X2cEqdzvBq8NngYrefdiv8D5
fUChgx37CxtpauoogJAJqm/d7KGmTt204QOGqaNucSxfpOWrkoFHkn7SfmnvKYhHKsLEuMYBWJql
mEI4vilOpFSMeijPbGRWXSmj9EaGOh7rO0kqM89598rW6WvHRM4hRRA4RrqkbBwRdnlYhUlvvzbQ
p31d4JBuYaDLDu7We8Y7gM08JLCldYf54apt3GlDjflUyVAWs8JyltK2Hgez/OmnQgFAWtyxwx/z
ZmHnRHgggifMUbJo13dLXWAdnNFvkshIam6fAeeZpENQb+ZV5cp+RvEUzZAsKPA0pBPhCzMvuhZH
eMagosWlXhZu8Ub/Bh10YSUKGAQn+RYfQ5dOd+YXQozAgowujCCegKFBRl825SRA6NhN8hjfCA0G
0lBfyjlmHKyMee967O7B3BBT42ICWF6JExv4GWbXLUczkERM2PYms3yXCM0uAacb77dT2nAE81fe
n49nAy4+f1Xn0nCK+GTc8eZ0O3e0zhD1V2NngR6EZGq4u2aIz9Gm2DgcArBonYmFZFLISd/uZkZr
qnbBIYnKc13OPg9+hbzlV/x1jjmCa5rWb8Dpg+FklXIZMgNJjALGCpAc8152BGv/goZ8vQJildCq
cAAR9rVt2i0Emqa8iw/Xv6NgH27kx91YzBDAz6qKFiynXcuwYAvuldg249n2P56tGlbBcEAkC5uw
OsZRKiIR2q/jbVEka8NsJMwzoSpbS6OiywFBEznY0iPujZbb0sJn6TDfx6VCNpZJmLiaoIFfjjwo
SCQ6ipJqcSxnsS4wxXiuAhgwGWOjcTDryT4cDlcIV5VF8D5CsIEPOypcLEn3OBqeZEsWrY4Xryf9
Yvi0mDj4ckwIch7Fh/+cymUUeqaKz2Ozq6D9ZGyG39n5qmFtx1Iw/Mxu2uHC4H2uEQf3vnYk9lFH
ZqqyUNsdErnOwSBWAGB5yQMfGybid0S1+nCTLfreaHjKCr9l0MyttcgSWMy7+qpX11Y2nb2eUIJQ
8cf7fUGW4FE0fS5TwavBnluIJVvNDviko0zgrtNNW/Ba2B7ysGEX+4QK1EeK60iiLyO88O5ztd+s
SigktTa/N/3DobyKsuZSA57aKd3VCpy5cbc9B6YUqnZ2DSObD7mfOrgUG0/1oM468YM2qR+6izb1
bZx1xdqse7wbYebztbGGvlbzFtwvFvgtvUAhmTDmf2hmTJM5popexxToWbAnGOlalKi+Ptew1TjV
XSwyV7B8LroWy2jvHxJJUyhGn5VAtSdA+J8st2Fl0xEE+6uP8UA4tTeHR8999waXqDF8FC7kZ1/2
s4KGIzLuuRvvDPXTlBJ0z4hAw/Z979xD5tMXrxOFFXFD8Bn1U8LjIzE9RBcuQM9koL6whw8FmdZU
CaHgNDcbKpHb1vQLy5RtdqMhkkS3cpQOP8kiWgc7ZI7ZUAtOkj/x/EmHEiCBNfNlaN6d0Fm5rc1f
zQBjbLOpZzouGieSk2FGNLuO24HgmhjhQWI6DzNhIrcb/6j7r8SrjX96ceyXzXRcTWJEG1ZBDrZx
xqmQBmQLRJls+WxHBeTE3pTs7eNLKrtfOjf1XTlMh7wihGvs+Jngt5yyX+oMztHU6/KuA08njpuk
FzYHAxlluy4kofH18RX4KEihk+Z14jeGV/uOWpwoQXrFF7FtaU50nk7roGGELxJHDCaaefuwjs6a
65j8TQruul3vnEwqcbDQe4SBhElOZ+D9gSbWB5vrJNVpr3wDWGKtcKxrOWlTtr9EO/xUcWn2RSwl
h2DMDFi0DJm+i1eLAZ4tYUB7dpifxqjKQCgvRbf5wOYvoKqfnHIhkM193P6apeAEu8310Z6KSnXe
BFyj+0KUmkVC6EqW3KcMh62ICinh2HpqCB0shwjntOkxiLCkL1beYpNRNPMfNR2r/cWIdGrEbFi7
KT3V+s0fBC4k7XrZv5N+8MjUAJa1+cshrzJ9fRAO0krd3o+srfXyjPH10KWN68UDHRVPaRQWTGFK
b0g5xdlbaSBY5psTVDbx/KPhfWmxADjLP95vzN3wJZaeZRRnAX6sJ/nf5RfGGrzlYrkV1mqyir3H
OltKk50oK4oni7DnXLBf9XSd7jlFzz1K3bN8ZCsQNmqJMDepipTkG3PVGAoLU1tUp0PwgQ6XkXPC
zDf79D4P4BsrhZZ4GYhM1df/y9jqka6qSDbVfJC9omg6SyKZ9wgRryScpv62MZSXmyHZJDDtY1JW
PQfc9wd5zY+N5eOUJvx+ElJnPw+Nilg5PJaCXy2CpRsMgEv8IU/sj6YWIY7pHTIu+1opwE/C0iwc
bvPGWzejWXgvJD0FBG9pMTFrshA0oofmcycOL4S0Vieo+wVyivS0yMCjBT7jyBWjTlP8kVcHcbJD
33PUnjAlfYo+t1oGYrRx8D7lcs/46lmbYaX1HCo7x9oQedoakgA1nzJ6MKk/m15A0gTTgnxchBVO
z/G3QdGeKSFBr/lwPVwpdMVaDzHfmFN7e0BFGQ5BtMM41Tbg4P/QJqKbL8MPR3pWhELdhKwgU0rc
ZOmTMI6FdQzCu7jJEn+OSXFmJQfUzNeTOUdxq7V7YBrUD4wRgXMsySgSoWt34t91mtWYMhlgW2Rk
undBIG3QjgFRJYbrNOPKjq0QHaoVVgAo/DZ+jKDyMQt6YSYKQ4msiQX0TNR2PjHj1N2UBcQN5/Ek
tbSu+6PC4aUJOskHC1b9m6B4wangEXZDTD3IesdYIJ1kSGw6denAh0wGPb0uEchpjO7nU8LUc0+/
dEBXEUh5iGv65Vcyy3v7BRNxwSKDOF/b4ZW3mOK5kDSn0re57rN9nmMdHdOhrLYECi4P8fQ2/geg
xWZroImpj0XVPy1lCcZBS2/m9EIxzZtunZWrI9dWhO2XCFpApzRmYDBXzp9Kb9Cvo2m68/Qub8S8
UZhpQQveziw520wV6Vzi9gptgUA+cM4KEEDM5SFqssYs6AP3stfnHPFkFuJ3RcfzSkbdmJ6aUOLR
CjDG7/EL0SpwfxxImA/VP0TaC5xK0dK69HL45CCkHAxIpnK6hSZPRv6fskLdKUH6uh+MWYTzbaz1
c6dTxUJJXQCHzjdsnO13T80JUQK+QPVzFBjkuPaqinitj05BnE75eZKdqZTkk/hPeqmfmYJQaIs6
SbEx/dmooRSm3XzQb7bjxeYWzNWA4dpIEmti1Ln8xXCRwC+gqEzVzKvthURaq/rxbQ0HBVGihggZ
gTYaaS3aWxrOgvj6+kOH8T+upUX/ljZNW5XX109aqyh/Sy2k44pHJzznhdSvdIJRRsDEqVj0hbag
OmH8LWlxNXjeGWG16PxcZDYhpeNaLlgEK0N5vtTcFoZpQeI/r3ZmHF38BMazdok1bB20fosb55zh
bYLcgMUP3MI6H7O5yJ9Qd3A2Hf+ch2l/xl33Bly2wMo1loAoRhEDk94JmHge4xSlFp0PVLaj87Fh
mSrhTVtvH8oCKfmjKksQcfcNEJIlcZ+UgtZ9m3Dm4oWTcX2bw6bYoneO00txMLd0nUBlvTDr9WBn
jc94WUZNFuth6TgZG5w4JJAJRHQnfALnpQPvW5MWjVsN3xIeynemNIBylH7TBrs+fCi65xNOBOAW
Gr7uOcBR2rxXkriLsqO0eG3iLtL6nhOqUQW44AkbP03VNIW1y1Bia4/Jzq1r6V8uR7oynq8yqe9i
QPQfPUZ0OkrHmPeACrZTdDTCszgEtj7xBcFByPvGoFWYjvIWy3U7MoTqwoea/UwT0Xv9QPwcg0mZ
HOk/gQLVkcfEZAM+NDg9f7n5z90bSis2tH9S//cQRv7L7SyYFWnItOwEhxcdTSmfBJigk4kI/7px
vc6AQarmDBodyJVCSy27pdPFhAhLkadF6vIGxX8WS85ECMfgdzer98fN5l9QomgLgKEQBLDX0Qey
fKFlyD9Cojz8FRt8ngR/UbeaIAhlvH9qZCmQZpbcD+MpkWQfn1GwdK1yPUo1dgZl1HKkgJ0Wr1ZS
V/VuvRNUZcbwINcjllxXZRhZYvZ99B/tbZWw+xfZAomVflTxASUxaLaxnlpscd5ttaTT7Af9y4Lm
UTgn8mCrbDD1wa7OWrEmwgXqA6GP0Erd7oLMGJuRO+IyOmHgvQFQG8+V+Jw6KWiHdh2Jay+GJY0c
wBUQ/GRmLX0bkAeOm3No2HTxY+b0iCYm1k9BJfPfIkISbjiQ1zyR7l6lCFQUPOMLCTs/U9akzW7C
PVt1jt4N9Ig75+OY9B0WycMjNH6vSibkD8KQH8MNP7pYhT6eg3qlPJqNAnSPEpiDnGOq3lZFjpbv
AKw9hfudd+vPVXW6A9ZRhQPmMnTJvcEdLNmsjQLd+2zvHaRywhvKY8VI66Z5edDTIquUd/bsnHF8
mJJ+U7OwTqUsDKt3Ivb7RqIT1hcoY7lgSHsSNB5WH5aEGZAqUUk/JDAoi5s+S+1V2uCz8/NSO6d/
m8BuFr2gBcc/4ztFtoY5Tvww2eq2178p4mBFAVBRzy/PSEZ3RZAw+dHdFCBUDiAwAj63cwu4mmYJ
sd9QeApPgApFkc1AJghgh7GLYIRmB7wmKXDhH5tRewGFnj5EpBX2Mn5TAA1fKQG226pL2S0uYJNg
0Udfv/WgBK5fmRIGaSu0fyBeRCr6UlduvumbfzcBzlYQ6w5sUj/ez5l+wL+Kfp6g7fYDrUlkgOWU
9QNJuoaKrgijWVpbU+6hkz0JQ3m8nB/D0j9JH9tikIEkdM31lXWVcQp7c3E8NiVQIoFN2r9u6z6h
AZPk4EGmgGw6GRH7cqmDl/MdMJfSz51vJWIxp4U7ZMSWDqiviCMAEUur+6PmfS9VppfuInkoii8Z
pvKz1GNB5+eXg1CQh5mkhDdS3VcXewkHOGzGMFvxDIx8/IWU4XulRbOo/LD9XbktqRzWeHBAf5ya
ZCCPPM5LIstfXpYNH6zb+OfI0DoBDj/OaLpKcXrMCjSQkMpaBhvNE/Le+bvsPyhUq60czO8KgaRZ
1BVQX8Cl/XO8XH4HNxfmEMbuDcSAH8J1As4zUT+pHUzTAREh5NwvX4/zbzk7zse92NPu0RPJhWCs
pGKvekU7a3PKQQBsxZoKbNGH0cTZJ+5sKX5yiaMiMXIYp8o+6eJ+QJAuNznV/QR2bRlBZQH4xlyQ
ncsZEFOM3AyY+fpjSpLmWHJBX3Kf77N2saDQKmoTegBL3vOIY7gS7yKkAx+DuKbAWcefZbxiWBW5
cI+AwYuI0bgcbKn7OBOBsNe71RANOeIYjx1rUw8aUXvPgC2tHbrf92/Lrnmw9UE7Ade7FvAQJezE
zYY2fqvcnzaJQ8FE8MmwKp/VSyzspg2IZZvKhXNeZ1NkH8M8qWyYXOEq9LGSsXJV6PiG1UACn/xM
TQT4GaaOFjTaoMLEEtGxChBnAhePcTU/9Sk25hb/zGLf0en6iA0HewW7wRF7KLlQ+W30WxEBWk9i
hlzy07JTRA6942ld+ErQ+dVbc8GGpiZ3+VSfR9tCF+tJ33A+/8GZBZmdl1oPGw9XTXhMTu1NUMng
MLct5e5RJsA1wFcJsO1EVVe+6JqWKudRcYbqvWYFeEymx2kTpovINx2Zbd3YCbvXifdSWjxG5gsl
QHxuRLW+UDi+NQasbfegUwzZ0ThdBbwUfqqz+jeeM93DUAJshDxaXMnKQVShsdSj/6FrrbjdRCQs
QCGUIuKwPOS1/8lLgpBuvl8Zm22aA86HSsG3L4B6bxvkyq82DA4dZg/Ff41JhP6fTvQbJA2p8aaK
f3IlCLcuWFtmGBQIOdwswlzkH0L/lu6O8Hxilq58dL6PXhvqU7C1QGl+5XPeHEvvVO4TA5icdxn6
Xl2sU/9JGYhQAK6dYOTZ//eIMjYrv4wpxBN8urw/yem2IyVAy9iaA6rDqwG3Nxtq5cw2TzA1c9Pw
aSotJ8++LCLNMhWsEaUuiFI5i5fwKlHkCiS7zIfuJ0M/a+e0mVm3uBuIe9rzd31LrVI2PiSVuN/R
rRxqgPpbQzWscWcfS6Ye52ANxPx/IaQW8cSvBK0Dgd4nLC39hu3qWNTi/fP3kXrTZhO2j2HxOfPJ
b136jjyleA9RZeEeSArshUJcMMD0URMMjgWNdT+MHKbYMVi4V9D7+qRLiapeU/EXK6aY2BDC2piF
qif+yJqqcoBOdbR2ivePsA17vm1cFaUSn4STVLAkQqdo9Y230XzxOF2Hasb0+V60AFvafkXVfwDx
xhJyfmby9WJ+hnch6sdZ/SeT1jdxJeyz7zU70uqa4lnw2nJbVH5LUFNkm4sWocqlqZJbfJYARUju
llaxiWN8HPp7Ekbr5N0F8tqNu3jY2M//z7mbu5QYj+MELVpbJqCQX8RUmJKIiuZHh6H2ameplt0X
KVtiZKMU5l+htYqL/yn0oWoqHollCxiuMVudF7KERJAgNzwwM49kpKYbKoeZyls0CAvAH/Dn9neC
8wibPhOs0bXihQCPS/wyB626ufyDZ7OUJzrsWTqqu9oTcSADsLwK+zX6fisfFdRP8b0P1jRxzWAI
rVMtzAmQuBHm4I4RBlaVcRkbzT7bzWQlO2ocEh3np9C+eBSBgk5pX5DmlwIb1yPqOUAznYAIs1C8
5f239qoDEk5xbtdxio5WWzoC/n2sp/uO3P2oFvB6dU2bqIA6lfvoez357zKnQu2m1uW1Ea2wMUci
sxBPh0R/CbpByIOtW+MCDBbIVMVq7zlKnAq7SHPIfF8xeurHz27S9X6WhvQevjmUtgcL1oeDRc7L
13mtuPjsyBaXsKsHhpaKK/rbMuyQ9R62BYmsdMH1J5rkyLRHVgciFW6NCTri6sbOqZ7uba2Ng2rW
2ne9e8EmumDV5wMIB/WLQ7i9Hjjo8E8Zw9SzBC35WmSTNuBEfB61WwUFawNiFhgngyBotv0+AZyV
o2OxTodwmbs0N6IoRegrVaSXmKJK2i2mWQ2lyFdug59fN72Lu6EhxsH4vydysUY1Afbb9w0Za9Fe
DU/IEdBgXhy/wxf8s/DxOm/fZzwPC5+VgE3AmyU0mxGia9x3slrFKNEJEnclUR8kia7H/ewxznOZ
xAKH8z69fFbSK7YcUlAn8ccRaVZLBeaG/qwb0gtgLV2aKciDph6+hkp5XZquibmWq9KGJ2uI1zIS
JQRG6ZS4hM5oXbnmcLz3PAQzvc9rubeOfjTzRaoO+YcaHTZdVTF59xDOVgzJJEMTSxMf9s2zcQKZ
RxqYFlWfKiVMA8mlb67Md09qWiKaJe53rqPJpD+QuvFVUgZXDhg8/4nb+MBXl0MBBLN6BNgCbDsd
kico8lcxlAklOBTdJM6xUuSJGl3OiTIU1SsRSpeEjgVUllvmnVOuBnxKJa5QTjTmRo/cRAN9TfVv
cF+r85ln5kWVWW2gELjH/MhYBcC/yU1RR0MmETtDMztDhj1TC95ByoOHWkSY4yvMW5oYyYGIx1It
MfTevrhmM5Q2GorDW/ak9U+DTbs+nu56byQUAAvbbr0MFTPyGXVYiO/YDD8//OuaTT7vouT5Cgck
FjEqsYWQzgzd9S5HvgesuMSM6K7OTU2EjAMXVFc3tWBpa4Co2Y71SHDiS9ZUtU2dKVn7n4R+7AGF
5LM/YJmSMPmRQy+XHwz7YmVQ5e0s8pW88sSbKAzo2f41hsd8sK3kbryXCz8Eze4J5vN4BCYbniO+
y2pXFD5YnvV3L59NZ0BZCf0Ng/idG4lntIaMsN8aotigIPAoE4Rd2s5Kwj1wfzD3yLwHQ5NTBDCP
EoP3Lu0qtkW9j9TZeDFihGbz1Evw8wWECfSgGbu/KfPqQDnsCRDUSsxl51kACPC3QVR60mUKzUHY
TiXILTjDLMuG4e+KOZ41gIYPsQkyOTzCaU30aR2cmceV2D/tZeltKTM4FKU7gobmZdxx850BV+12
KB8oCudoS2pwBJtMnmDUKUvIBv55KVDSTdVSkUId1N7WN8awV+0aQzkivucM3FpxW8auLI9qH+0i
ztOD4iQEA1ljxNaIKmL34TTtYH27IB8T6aU68jU/GA5ZfoxivuC8QzRljjqAvnnb3FoXg/9v7nlf
k5OI9nCeTpw2ToMmv2J9+JUZRq3fb5mGx6UD+jItPG4TOn32XZm2PwoUnoT/McqxCPJDKGSBqZQs
OeASRHSG30iFr+qk5utofTcC93fZXysKpOW5TdRLtUjyLkA8Ss30wJ5feu0q8TcU1Fennah1IYu5
rhLiTWVST9mifd0xewa03f85+uk72Oopry1ejm5Jcye56IVc8Mjy8J58LxYPMBQt3GoUFpzQ5Bld
5dnDHoVuIjPlpIyI73ZIFVxU6W9DMAg/3E9VjC78x7Isp5rGiC9+LNWyWjrbQzey8zyScqtS2zJq
h1qoRiboJuN7ZXBLd3xjnBsaVQLwb+S2m9VoCutHVKEsPY7sCJ3TnECTm46aRONLIGNYgVAOlfNV
1R2CemhQAZVE/USbCotpFD5IIoJP2JxhT+iz0FlROoeHIIq27QC/eN8IKYYe8+COCU/TkDArLsMw
lph083Q5sZPDY8yvBGv7Fxd1XESPX7jn5TJo64DSnzvJ3i0mdnqRuBkYw6Kh0ia7uxqvjiCymHHU
pjigcIybg/2JqAH4h5nFUx0eq1pg7EPUqIgCcpUfD5Ap3sfmLPN4KvreuQiHEwUgflP+p4yO/sHZ
DlY12BAwapoEtj/m+deG5z7ciku7JzQUSuMWnps4oRrNWESiM+C9R7WWAnyytptHzd4C24Bn+hjD
/ybvfNj6HJ6yrZVMQMyq+0nfrbAD25Z4+TqWoVFxbpGQtEaeErv6hhEyXEj/z1XvG2wtLjwcMVLt
5TW8ve0V4gLD4Ks/jMy/1N7foI5E633hYf5D1IArtp7Ynpah4D5QR9NH1td4wGC0oWKHrqAx3/aW
M7CpjgFMrz3GI30tpCcMupFlVTEK2/6fDs5RrpNG1N4Sxir70Bo98aJRqw8S2e5SvgW77iElDybQ
jwav600ZeT9CGjaYW7nJL1kKV6mGYHQVneTbX7M4leKIhTCl9PMZQjTYaL032lQhM5ZZVe0UWzRN
cxoyoN+QX9SsI/uyYuFQiZsKvrU5MWZ1yKz8W+W7luJTHLZyPRD1nz+wCbw+3SrMtK5yJbFza8HD
++vrGmTFVQl8zrVd2tmGJJycrvWfUwWIX/4YkRjMVbZ7C9bStXaCv/gZf/Gb6kDQm7eAVETA06dN
mrXMet5R3vTh1ibyWiSPCO1bYLHSM5qlU5+DXOpbMVZsTRw0PxPW3rijCdab7eOTUvhM8Xmpc/fs
MUVWz0GCriRObkllcUPOepUV+ACcD1mHMSx4LerlTrUH2GVjSGJKFsAtWOFOTdq0T/PBmT5SDWpt
PM/13vgddt/eS3cIiIO+KkrYkO3OsLeCWkUJusrsvM9QeXJK30WWVTQ4K2XIMSOUaEQGc4j61gx2
EklTh0cDNhStDODKIbhfNQ+UrN7BRfTS1yt5X0OVDbWGR7xHbqzHQvCMEd5Yt5pyw5NILwVAMGUd
Kh6aqs8988MRtW1km1X+55d53cKlagPfVzw04wYsD25ZLzz49pJM+RQaud+B696DX3JgugC1UVuF
l35rmeH4KQRzvG3FOTbjrZUEcCneQU1QfraM9fqJnBmGz6wwr35A9K21neYguqYvG2kYy8AwmsiV
Vo1w+hvw0z4qLChnyWMzan96CARA5G/VhuG9OklpsTNbs6vcW/sWimVbI05nskaHqH3HV+LCD97P
mbgZjODSCR3U+cDEW6jehT/7p7lgi7NQF2uP0+zHLlyivpwWaLWvYAt509mWjo+RyGNtWZZS7b0V
UHgwEEBCaPI7RM6y7G8hWfHFUpycMyyt2rXf2TzSGgusGOX/XrxO4HEJad+BFeEQrjz2ms4vNVVD
iLmsf5yqJD+YnFJeFe6txOApLW29t2XswtCDEzfH3aB/mmHWfU834cRuQZmfnBViBb88sX0dMmcc
XVg05+5YgUjgWGvr6zvi2Rx+LPxkJFiGvsyw/lh6w+q+9kWQ0BX6PQxJrMMerbFxepiIc9osUZIL
fFzkhSMg8ctpx7Y2FHFzKoLcH3Uf4HBp9D8qLRNUWQz3lsyKlspk6A/CYxuRBJz9rfm53wiOcp4P
HmAIu68xUTKhyxISzXwBD2s7RmfO3h5TReI2H+KbIi3V1BOkSD1W6XxKn03EBIQbSEsp9rANyO/f
+eEbQkVc/bOlUVuLMI0ZRK45RMDJV6Z+WRIEV8uDEKtnS36JyYNrP1ijyH+vWjikSdc2XIolImwY
nHugvPm7HqDJ1MnWW/IzT0BZq+Q5EMdXnXg0dRoelZx8kJnTu4neKCD3QKEJmgYym2vGLWPRY/8C
TqYPGa9ZSj5aCLdYHPtrZM+fISAZEoda98KjjgGjRL9x3zrwHBGQMTsyOWwnIysWhjfWMoCZiXWn
QLXsyvSs8IJ/ktn18Fp1ei8/4DBt1PrZU36H9dhyJ/TZEFk2+tTDvR1iZbiEUAkUYjxpbFcxXh9N
Tt29YVOFTFV5iaUuAe15BbqcbP4dlTEH82Y4bj0bYVfSbyngfSDyZNm0pF6U6/+9FGwTbHKQmOqL
BsEOJ2jdKFFZmvGym08T+xTvUTBNnR3u+ByGhDjKQdAcRpdNlkbbbssYci7mPGpBq6r44i7+PXMD
8bkKAXdMd8d2GuZGWIM5A4qIZxfhAGWm1472AnVoIbJiJWUN3qh9fduHrRfkzgUpZb5nxn+qTHvc
9t/WUw3lSAme0a2wheCTioC8XRZA/MKhUQXjsEf5jRAflqqo3QQhvF+T6yXwDnRxGuPc3c9UlGXO
NuE6XygDSxZ9LzToSLqDIK7dmJmZODRwP/TMGHpLz7FBVXYTR0NoqWVUwKO5PricmxoCPpsA/+mD
kui3X+AbIJGyJs2wFrQmg0jnwUr6Bx+R19aj+f7M9bfkHh7YdNh7qEjgUWHgIOQWV2AmXzL3z4Ed
cs+IeFDw+8CSHf+P4Q3ZCG+uN3guyO5Fhni0PgLRn+aOXV3ofY/0KZD8EJf2WgsFDv2uTQykmTFa
s3wM1GpudyJdJRDvVzD0Yq6Sn8viNSuaB7LfpTNjC/nV2RC/4j2BjISLSMASxK0e2w0ZSGdPIpQ8
PpAnifCZZCu6SOSG5bCPpD1F5AIiizWY3HtmhBn844SXCNki03h7l7j8JOc+f8GepSKINaXp1WMw
Zh1e9orKzxjrFRLk0vw/SySM2soRK9XrCUj4yVqDcz50c909KozMhGtfNqHE40OgGJU0/fW+XSc6
tPGdCPxSrUcHkwsYw9DqWP6jILAbaTMjMfafzG2vZoOIloJA2/F8t/GM2QTE0MwVPb3sLJgfr0XK
1zp6G+zTJlmASO6zHFvwzwv5Rzd83vwIWfO/tupfUF0PRzQV6a4q5kwWdoan7/ekG+xfyCL1AfBB
oMG0oJ2KLxYBJ6HscDz9hYVfpHQ6jAi9WYeG4GCXtv5vxov9o2K5ZOThxpnTFX7lJC9aWEa1AKUr
+cEAH+qmf4Z3XWGlv+2hMLkRcn0SulLTakquFwCmxUqpPWofPA89EDi2+aRQtwz1y+tsKmJsDUzu
GPtSMu+uoeHX3+L23VX/4xA2u2fMUkl3BI77e4NlVdnVxEhu64w/NpzKFGmIQm9iyzM5dEOEWs5j
7SfUX4wlEnzX0X9Tg4KOrDX26wcAUiUpHCu7DHrg6KGvD56tMvkhsCyvrNcvpT3tllyrJwE7jA93
2jsBBxreZAJ0gCtw59RK4T9bNQ+RUQhmA4jPIjkro7xPxPYlXESZG05ZelFZSrPRXA4zOqx4M1FJ
qWnDG7JFQIXjPVuFNwEE381WYchmwC9wIbhjcGIcmT8ETDMdO/XBMFpszMU2ni9AOrBZOqSShS/3
z5USmoO+rpTHKQ/eSK/IatI78mOpyv9/0w6eteM7ZEV6eHQu9XzeGEAqzA7WjgX+1/4ni+zB3nxR
Gb9Vofor0yEvBxomdc02/NDUoKT8MkxtCrU35e1qpSrW9dt9UMkopqu28xI1/a6YbVo15jgpuZgM
vXbDmGTn9dNNQABj95keVCZXWLGwzSOzqgz9IFITaFZRw075hlv4IqGkLEfqgwIqaKjPNhDEXXDI
vrUnhc95mq+k/zS2+gEKmLRDagRUR7EIszm1pFNIvlLucD/zMAAsLLu1aM/r/o/9fIYJgfarCR+h
lEQhgjmijcGkoBU2pfEZNedoH9XorY++rrG6JmyPWnKlgBTTfrvf5Ug3RKOpV7fty4qtHDYv6btG
CPthGBUafNxEl2gzO4w88ZlaqMvXhltJGPhHwhwtKn0MkodHE4SO1tA2qmRkFqECjKFCiaJ5Dt3L
JC0jL7KsVrMcgx7Van2EKGQKQPbqZBflHIiUwG1Nmzyl94le5ptWDJ7icsZb42jDSR3HRL3cBwtd
SB4ZeEAJeeaq7BftbauM4V+y/LOH8TcjQwApAGHUp68MMaSN4Ux+8SmDCv3KXtwlT2xXoFmHEc7R
LrkHNvmYN3fUr2Fy2bj5oPwazacs1yHKPFdFLftQQzpuwOazgskNM+Spg6MVYZtq2Qs8ByOvpYES
43U09cykm+cyrmxIgE9GwsaP2elXJQHgej4B3T1IkjcdbonDg2f9Vl8/rFwchvdMAnD3W+kvOtWC
hjBbt2VLlLem4lMsiml56/h8N2OwnEMuZaLTW5/jh9eytY4dki2tClHc9Q7ffzvRYksVh6gHspzo
ekwKBPRvaSAFXXIuSDJu6MnzNAw77Y8+jgGCe4oN2KL35W2/iqFZ/zr8DxQKoIdgK/rQv5fnO2Lz
cUIHARfq5EUxUa1b84c4UdhE9J+xOmrg9lhXHJwfnyWxCP7KZsIrjONHxvxfy7uKYJ7H0UcUX42N
aOpKjhbZubOTAXaL9zZKR/wlVTyG4zby6OHThM6i3npBYH1XCI8PUmjuew6gcR/AlAvWHHkPhu6x
SOO1NQIyMHczSYSUFunIxNAH6F5BqXtrF1ZuLGTJGJIZRZjbVIKqpJ9SBZJ2jY4Jo1bjyk5x3JGs
3AUGr+/5FSOxrCKz8mZoM5SUL+bNEzFIWJy+ZxN8uBDWHe3RiKqjIPjymQmpAEVsXe0xapfqr5Kj
EPcow968JIXovs40iwDNj7XYsqnY+i0GWdjJql+U6cX8bklmDDgzf/q7sWKQtTyXdvUjZZHhqRzS
xsxgL3A+0BpWU89QHzZ4W0LsVa5QdtP7dX2X2gnAffYGCPG2MB+rV+tgGpeB1k/eVSdguWLhoybT
GZ7Lv6Tmdr6wHyY1kW3x0Jv1QwISUzXQIAkggUUpHoaKyRiUaySvWEe4/MMR30DQxj6kE+mgPI5M
GH+O24XFBWYBsiCAyLqrDofLsWShY41yhLGHyTOMqUEi/fE291wIJfdyT+b5lQkfUGctgTrHnhbg
l8hMxKCZ78ukgwx3Oegc2Ivde12s+RClT1ny/OoEpkGtF+u/LuGChu6aTzRMi3SmxSqskZ0WhHks
WoadDIoD+9TrLShS0Y6PXQLSYilQ+ZjGUmhumpjb2JR/fXP5WGb6YaSCFuoezMPpG59U5UWKaJDh
HRO9NG5bQX2og+OLn0nK7ZP7aj/APsUyt5Id/hcv3myYxgefuDqTI2NL5GkU59nFnFdlhwrpcuUH
OSeFXl/s3+Gvh0YRlLm4yZ3v16KMzFpw1ZOHO1jJVGryf9q7n4z1LsRi5sglk9QU4l7UBAaQEciU
ffeUAZnfJ++D+ADjPzXV9UWhXU8vuQJB8deR8h7ZqsnVxUQEj3sZZrnb1zGHNbO91HvoPuSblGKt
P3cCfOBbBvfgGjlA2CQD732eZFszD9OcU5U0QjVtHtO1ex+3m+7WxcWVU/s7QnRy9cx4tUOxlNY5
HnJABTwesACRp142ROVQukGQRbi6QSRxtxoGl6IxqXlP+k43bZt5M/Y8smR/x5Wy9oOxd4AZgPYg
J5XPsf+k68bflO2s0arKiHwFqf89EH0Q2/iXTQj3K2awVPX3M9O3TG2FW5L20U9+OR+rdUM1J/iy
QRl1Ri1b6t3hAeyNIHVlTy06elbN5/7aFN6sxtt7Gs4xuuD2tB8z2krvKqZUcp9SOxzJ8fYlUZ41
VUai23uJs2UeBCWu1KTKTiozlkqm8WBcfZP77un1QtEF7Kl68QttCHfXIlKAWs+IlMLzZ2QVNPv3
xv+MIDl5L+KZ5BElBN7EuT1ykv4HAKGU1DSEd9mPLQwiVbkKxS0ujv3+lyAkpMhHE00RD4PTOR3w
DxqFTwRmLNsaA03xyE6Q0UhUoheJ9mntM/Gu07pZAkFLzBfWO0+eO5BW4ZUFNm9elnXH11P612CH
SGwLYLcdF8YcxfJzzmahfvA4BhoEySqclvKyQln/64ATxs75HOgLXg3/UWTPpdxoXmuMQH1N0ufm
7shaibkWporw/c8S0mf/CuuYAJzlDQ6RhnRGw/+GEMGoWolhkNrIVHCfSp3L1b1b4DPA22EHpnTR
9MOK4QHOD2spUkWCOZDNhrOraLYmtHnnt0cUmiI5qDROjViRPHtVB5sjov0/45FwC41sk0HBqCtw
LBam0DSFx+SnBmEL775WaHsdBvnMgm37wqJOeo8FgtBoBrV8Ltj+CHaOBvpaeWzR4EGoHiV1ZxWV
Jw9qtKAR3eGypTcgNFEEyM88PTbbNkXPwgekChlp+5pFGFWOUF1kRae8tEoVAArZDfsAgxMycJnj
OX0qhsaJubj2wn/IwjKhIMj5hsWWonBVybIvOf1mfYh7vIJXRns4I5wnhmkvFQvag7w4DAeVlchS
WotfYyRkDoskbYO9LN6nq7Thtpe8IeIgRsMImd9Yw+hSrYgle25V8M5iRxhbIZ84qUquy19rhRmG
g1rW78XZK4gBYiRX0hkfn0UBRl+b5AkZ0VixBKiV0yTYzByPw+ik3FUd0sxre3zh2ykYlIkkZ+Yy
fSrJI0NU9BuPyki2fIVW4qGtF4YSvqZL+Yv7KzyX/AGbATuIFsg5fknGe6Upc4Mv5kwCllpPBsOp
aSbXLJkjrGwTb8Ld57mCv8pxUcmR7vFsNoXuj8yuTIQxq0U3O4K8u0GPn3thscBaqZnZ4rlCQ33k
Gmnd/8LIbuWKjV1F8O/lkDVjd52ToLA6lme1hEA7wMaXSf7vjXvJM1X14krNS3447hQY/dsEkExr
5E9WLCBhWR2q6Pk5rzlPgUkbIAGYWB2b07QTDzSyRQryYoTFyDoqZls8oXpHnsE2tojx34zSgh2Y
ZLeOarNzRuvr1Sj0vxTAvavFZvW3qVtweCUAdivri+kVP72/WdwOwGH9TF+QeqhwM3d+E/aqqw8+
grXtZUzzYRN8ZZiZSpgGjCw9VM6A9xVE4D5x6pTcCLXy2IkCKdoN1BHqbiwZwnjj0rq0TaC4v0ZF
pKtC0NH2utHvwVQ2u1zheJt1camR2V0VtVT0PB+92oUg5Y45c7UJbb+ywQzTrFuPWN5nICw+u8wY
pZAbHcYJr6NlM6IVspCgr44AElkSX1hLqIGDaavtGW1KghK2CdXmz/mTBWdSQjD1Auzl9iCHYmWT
W0CWaNGGdvWzfNwpSGrHnOfaPhRSGmnalmzOs5BYPhPFAFNn2Ul3LavFRA21lI99B/GEb/ftZdez
GFAGYt9kzRoyfzIjzfosTs5IGZib+ChFa4b5UFdlP9NnDeqCKLh53w2xFrljBesCSikIn4zACOaN
CR3iKR06UxtUxLdv4F2qartZZx+MOt0VjLdaBKnHg4hzBdRaSqBdq8itn2O68erXAIXOyKBJ8XLz
GmqE+9fV7VNwp/pqzhLuk7uEtzzCHydyNn1ye8+X8i1pjMKNp45dj5EylEMPQwAjjKGwOfYcPVk+
v/MxsL62mmFGZPbCdhEWpSy3WqkDftZZKTobsT0y1tyakJwfaeN1Qxs6jwj1EiQVL5mrxBxL9QKs
aM0A3gAkZuBp5idsIu1JnA+Z5PbA4B2D3UrqCJ5sUbhug/gQ2JoetE9ayT4TSDDTQy6etdSIhcK7
E3sp2aIjpxHAh5vx5yuVSzgHFODw2P6qpcMqZ/ocQmUQLKZbQ1tLpwiafccz3/CZge7NPqy3Riaj
l50oWlAQJBsb8/gn+2kPoUwTjNPgtN9Sc+ABE4kvYBcx+vwBU0RTsy5hoDYe2UXHaejpzIp5UqIZ
G+Oc8nydGf7S7TZ9XVpRmy1WkULsTWm2BvPszFaxHOqSRMTQNtzjvTWHb+i1EmG8BQ4UARjzLR3k
WLGZzS3cBiDBF4SZeWWWH5kpuQMmUdM5cMnlb7ZFasv1mVcjDtHWXY3RcQ5wv6ceuLDO2jNPZNjc
j8QDNfPQi5ckAaZWjbrq8oelMlvH81mt92lgIjAGjqnUHuFpFgBi1XQ9HYDumiZL7UL5RLx33on/
uUwJ0/SmNOsFkMtoJyikK9VOwKYrAzBQqG8H0s4toxuGZDraQNCvK2oTXRwYI9gJI0B9WCrDj64d
uWXlMiVfcWxpB4clTxFOZvMo4tLTDKsvDL3X2OYp3zR4cpHIDq4RsklrR3dSEh9lkgUA6yCBqHXb
waxjcfoLXzWKrRJddrbZDUAgpai4gZiiVBeV1eM5w0TEkhYZSK4w3ZYBG61LLJ2pFUYwHVhRd/q9
S8D86ZMFNLqM6m++X2KqXvBfK8y5baqkx+VBrakWudsCRnAZ0W53MLU4A+nAP3Nav5/wE5jc35Hl
CKSeHKdSj6bVL7RGQ0FFrVamdcDhVbo479pVyuR/NLus3eIoaD/r1NPBM0uppfCljTWzh704ZbPU
SeNw6u4ZwPA8ONkwLD3S8CWNOA3nrsA1MR8TJ3596vRCj4YhMhgoqY7INlOMiI3Hc0pNsa+Y4TIs
avetLbktf984FBz5UxcGTTwR7HEUN/UwJrb+q1mc6tycdKYOG6D9qtO+ETQBZRlQGFDVRNnCzNB8
mqwb+ppltD8BxTcqAD6/DScRDFy5xZVFm1mVG3uuXs6F9C8UqWRYgASSD9nAnLpcDRw7D0QGUEzy
ow9I80kp96BOdFaz7Y/xHQgUD0y/CtdGrwXN1BHyCxy+0gG1fowY+M1Yti862RzgE/yUUufVOJEV
Ms5Fl/cEeZjhD83lHMNRPcppfG9tiRM2SLKyMjXW2u85V9qtZhJDdSH8upE0PVz/r3I6wqwywcwZ
mPszAcybYZsYVwHU3zF2ji2Cm1BAep5Zw/2O4MyhzL76IcFzlYTYpjwAhEEbIjLaxB1MzcIQZ/rk
JS6KutAb3eDwicjuTLWGcP9QYEf/3j5my7siU8N35ZxG3Kx8I/z6SVpSliDWIXXxEieM+pKSvx9S
uR8Qox5WItTCy6nR/CWPFIhuFn9+I/TsQTzgjwCEkAu5owand2OFf893mj95Qnb37ea9Lgale/zK
4G7drXTLEKP+nzthvqe7TgSP7tsgjDVEKJ3a9v/BkgCjjwUfT6UQZV3rd9CEBAbGn1DycoTHfuZq
eGiSM0oqgVYH8jtyrK58OOoZBnbJe7Ubpj60Gs3Zlnj3dw4SkiJO97+mDzKSkal79aFfBxArDwHv
MeIdo6xbr4ONuUlLqmV0EWaz+NWrecx/VhWuiAP4Sl5WzzQ8tjuDL1SV6MNihoirkwnNl7anfkbl
cWK7jI36t5c1b/9RwyVy4waGrR3ZF7sWvadV5DY16F2e++IbZhy8hir2ERhMnCaS/LLKgtw/yjSJ
kgvJmKdkwPCidluv58Uqe6r4AV81meSE9LIsateFm2vCFx7USnCEuJ+vKjZIntGvQ1Ml5CVN7/eu
vXDAxjS5fkDfClw8/KmwVmAgsb3H3PK6t3SvvEYPe80mPLhUwFOBzNEv/jyWnzQvnNLD3yr0J7dj
o9oIaZW4kCOv2iyN2R4ZlNlRY9a5cvN23ioFkqG1rIgpj2x3jj2l1vUbQg8vfj5t7zTBKpDNWg6X
eHB3HrABKHdgohLY9SJF6zOyLFqycnkuNElHHOD3TCV4sKgYw02ugIAodsqpyOmK9IhoewzWrilT
YEZEWaM6hD52UftB52VyV5Er4kwyG5/Kq1Ttc+5MDPrDtoDxJJO4xWKp5YO4Xy6ONUOJBoECYnqv
s3LivZKGKBYm29WfyRegi73rjHoWpB3UC+bkg94l5+VgRLMiL4QKVe1IG9Lz/VLV900Hi22b87g4
1VMrpUpASFTrUVDY4ZrNstgDHlzsIIagXfgpDJvI6zonUIPDAhZ47xVOWnwMMnLRbJ304Ih5DDIV
e374pabNQOYfAhMzSE/SMRCILCMTfr8zplA92k3XvFKbCto9iue7910Ogsq5YU1WoKfD5PAxnBdd
bCSv2xcmqGBVZLpngE4fssRzvvYCNp7lv/gu3vWkh7vYC9cKm+ptNC/DL+4Vmjp2ynEN72Xt+NNW
Ky2LAbMdkuwQNzEb7T6Z+5v41/GQ9pWsWUeb0JcU5+LRaWvNA5Lg7apGaq3JXjg67EtLTirgXTgn
mRlKsOnmmr0c/ksnE/OdRyuWU51LbwZ8b94fRR8hb6oqL0a+9Ky5/TXF9BqV2yCbwhtcUifpp/mi
M5mu42+cBJWldNfW7ZoBtQVfguxDmWyUsJV+whwGNY+/Axagj3CGSscx6NwI+bnh/3QOgnlmcZRP
72wbKhnBqh1Z+ZcJNL+80o5sizt0SCDZZQZ9kf/L8jiZTGjeFOkHSKNrJfydDvzMK4s+W01Lkh7M
SsRmzfKKGIAKkALuWYurngdZ0MzjmpI6ZvEctsbO7Bzod/EAGmvrJafwpqkqkvcFk818q+5AobCq
syvuV/jLYTecO8F3iN7japQP46NFrLp07v+IH4GEYZjsz+qkY3ku+0rcbJhi4o9Rmkm1QJz1UHcV
gjg+SpUoCY7UwGGfv/6gMhTu0O86DrDFmDOWwU01JIWTumFWep2YRTMKCB+JESUm8KAggB3AwI5W
N9fWvbW1xs66H7RfmgFXsY9pr5zsUabK61D0h1A/p6kaz3bU6bYGqwsem/tymSoNDzy0lE5kuUCP
BEABJJETDCzVY70STW3dX4dwIbtyusLaDsdeKLQcs5OJnlUjbfNNc7Vpv9QwVyDz/3+RM5ms5TG5
3aPnwJU1KATIXzimIYXz3v6swVF8ekJzdyxQlFv0+9AyRzVI/4iW1GM/lkCkZNSrF1A0OsEBPYmf
YUNokqOtpxe6monm1k09QsVxYqSdHQfziFEwWpxmPgKY0cXPQGhG2hKRVXaX5loFA5xVIWdYybwj
5vAFcQvCizjD6+1kpZd9B0v2tk8nX2J2/TUFztVHDIWUx+L2XHwSzeNeQV3b/g468pyhsUjMHq2z
+QGSlaQ3PQ7MOYjvin5LUX6qv/iP2/8VF88Baem/zoadsc03UVmzMa3MgzdO8XoAbEnkxfiVGNkD
qSAoF2ufo5/r/Hdsfc3CaLsWE7PXpg2tQin2S/Kyq55gdKws902wqbM2axd1uF7Cxxpa/H57qS7q
0epKnh15zICsqWGz3K+nMW7RxWjpWg7EQanflOMIIfJXH14FlGaoKJkTCzxdPgUUnu78WJ1iVAAN
Cqh3jC9xzvssXO6XDE1Z1ZO1VE9VsDFlF/IaclxsPO4RsOZN3ZAK7CkBKkq06R1iYB7furK23Bzo
7Q9Zr7ZmjN7qMshBpqgVi1u2AGTMMVg90EqWq59LuC9ngSLx7mBrt5L5/zrz6qiJSde+E7JpaF77
l6KD9Lwe6WOO6onVxdkWVOKWUipX676LZLqzyucXojTc40RlzQHBuMO2GNJvKdH9YVE+uaVmJ3Zt
c4j41gIWXegcDuI7yILGZeIDIzSs4Mpq/Iy/JE7qJSiCVGTTN3m28GKMQ5bbZF1QTh/yrNSdawsv
rKlq0tXxqJ10VlfPKI/Fty9b8MxWjBRCwGlcCaniA6lXJK0tjBdZOgVYgMplM6b035q0NXMy1qK2
jwRD7r8ZcoXifUGNjT1r21zGSc6lSPyoevpnbaFD7wBHPX/2slfyq3/4Upoze4+QQR4qWIl1HxiK
EyHObPg2D1b8QZYUTGzEsldcgCRIpLe/IQfV2Y0Lt313sNo4QsQrviM5aN9GCLwQPYTD8VEqMwiA
5SBiVgiSVeAaROVXPUGW5HrEvV87FppbCgoO5TOReiCm7cbmFUSI3ql6AhR0IjQKBRhZ1sTYONu0
o115vgx8MO+oZ9yZXw+8fCskKTi2FoN1jiwYATobh9CATqsVyFxw/qeMQaXgNcLWmqURmQVEtrc9
q4m0Ge2cKCkhAGOr0CVWImcEIXiT1GPshSVQBAwg/R9VLM7latLugUW0RWY6Kz3fpcYDyDl06kCB
UN9sDoMPxvwo281fH2uhBI5cpX6AmsHJoJ2dypaLxF4uiQoyHuxpXQrOnDxKhBOm74tGt1Oc03Kt
Z1W9wA+JeKxPmpe0HmvaYUqoEDQL0wN3A/FqaK1E09USJQx3drT6hECNv72rI3XjmCdhqKDBq/Co
+nRdDxTdlOERnB5aC5oz/qWb8swwT3VTdL5P9tiDZQljGuSxSR4w+MAhB1s/ZWVV696VzTzVpPKg
jg28Aq4BlKXt2dPjkh4C5ZSzGvZ/1EvP1TjvaPNzzTJiXT2HOCujIGVIZl7ZA/S281OvpTyBgNao
g7OtvV5BK9kl3ExwMw12rw6/6HROqE23Femi0RlmSEfnqm2s2E+o5puhQVOoIQvaaYQIF8wuOtv3
y/KPh759F9mS0iIFxcHtai0vYvK/ktfHODfn+1zZwZq9znc4vDAPa0PdEkNqc6DOUpYCba91xOEx
2PxPBLZm6JQaGLwGfnHHixH8Sjk7cyOiVRgU6yvtW/pqTT6fJcQ8w4L16VXcOVBYnVwDeEyw8wb6
djU5E5Kqr9HPuxvYLGUEpuhgX1NfHboYmQTSabrZj4SyNjbMXjpKM0z16ZzkHBUzG/tZNL/eruey
4kdT87Ps9/CiHYWuNKf1okKYUn63kIJa1zca8aUS3MrzFQDGMjOL147QWNZb7Q8ZVArFYxu60RAN
UkSXdMa79Jp8uK/RRCm2phGey8DrU/m8UBOvX62nQSoypF3ma2Sz5rnKERTCBE+zvrqhakRPEFnV
dW0ERmiui8rbaC0OhallFHHdjjp+2nshv8W9Dqvbd7QToD6ja0TM3fFM0GGfEqB/5lWLA+1cptsc
enUBmsfjHKBVoa+CzW3usobgsv4+ks3rv6wFIni1Lp2LdLBVTCcUVoxkbegdFhzHeYrFDa+J5pLZ
ejd1K28Od1Ve0IfQpWr2xrPhAWTskiUITiR6dogdCSPhknWn18OumZzD2OAs7//gMNH9m20bNdMu
vjdj+S/HjGRMRGTrxrILSO93/iLTn/fBAhpS+a55C5wagqggGddwiml7IUBk5J3CDrWkx3YXucjE
1o1qYNlsEU8JvIdy3E0MmGli7BIE+y/UOJCcdcP8qdR0+9MYpJtz/uI4bo7cRKVRyRnML+BkuNV7
6Wp4xvrpHbpVnbMH31P47HsPscwl4MAuIgzOsc7J81DDlK5MRtjRCLSgvd7zQPu2sNaQhVrJuErc
cs/3W1EHg9uoSDHuH787V4RGX4TQxlyC58KyDfR/UzObM2IHO8mlkFduslk+uu312yMYFShf7ZgM
uyCTptQAvM7hyHB9aiD8h6DiBZW5nlGkb3mY4/oALQY0r0gTSFR2PmEUfAhi7uunx4Ln18XvVXgk
XvV/MNzszBOxuuehGPUcSW9/WRb0q1yudbVxzEKSFJWuzZ8/yq8qwi/21XQA/bX8h9Si1rwU3+H7
l2fgMxnmU5+IazFjXbVXMd4Gf4hJFmBvOuQOkX+kFbU+Q1YVtpfdN8mHwAv5Av7XnHil+TKQTUHc
Hahe6jWeK7xAGG17fkPMoPFwGlQ9OhqwRtzATb7ivbj28t6GjW/mVU0LAxTtlD+TDIAabktX/7m9
ZTys9p/OnyUcun3PyCQpV6pe0Oji/PVML0/rLNvr2tS5CnNakOxhwxWB7Js6qM87VDZOTcICfCDO
inmDwsLzhMjl4i6NxwdzdIg/FUEbmyVaKKqiPrLgHVhEs8P/EBsJDd+M3l5F4DDXWDsYxGgNtM9N
BBNYI7orbXUrjBere4I0Vn0OX6KaGPwvtlGo4BdVTGB6fN8bkQqEhKhQCDV6LgfhJ2k3LqS2OXL6
RwXw+j8x46zF0usmuAp+1SJXKnUX+5IPeZpJclG0ozxfAFOj2GDJly8kvyK1rwfOKpaRU7u2+POn
VxvWEQ5Hp6FSGPwYi6DYf5jqTxXxvjeToyD3th2Wq5NlnXG/7x+8dh47mUFH9zTetl+WlhQQHeXb
e5dfMzyxcAiteWbT/NT1hCiF8gCWsi8dN4rkkRrrdwcN7ec7L7gzmBEiK48mWXO7Lb6gIdlJSCSz
l7ik/VHqErf4ZnMNriJ5bvkByvNqaP6ZNQxYJzP5Bja6ndMIPV3IdCxexGDp/wn0oI7ypj6pYjv8
v6p6/yENDBnoHwGGCzKoMARKz6by7jq0TWqj44AacdDE/A/giMqwwJ0Y45W9t11RDpz10dqRd4SU
qb07FbEYbbQHc0ltOb2PKhKYzy9Hb5qoBGJnOMvfvQmurZUfQoAp07I3HGi1Jdwd9S9OEWh46hs7
PICiLK7jfUk88KOrcKWBKgWxHHA8zDp6tMS/GE+voUKLzwe/W/ID0apObUolc8pT5TypL1CYudAZ
xOwquIhH/aIKCAwVbU9MGh30XvgJlGGFy1xeWfPciQjTcSjNNZyFWb5VsAtw6PaVAi3ygc1LbN5u
39RKY9aU3tAnaU377+iSTbw/V31ZcIrS21Q/c4KqljXp9ZGLUzJypGXfXXdKLUrhe1OU/AMhJq6Y
tX7/S1idvqj8o9VjRx3pVyA5xcFsOvVo2GC53d1oTPIs+vkSGqqCye5gQbkY2hCoVBQZ11ocXpee
mP5nZzn8lYiFOLQaZCHo1YAaahilUwBWq6k9xcF0WChWMnxjvRiin5NBbmlTZrrvA4U7BPt8YD7q
64k5C2SonGTcxVZuUeRDOlRvcL5UPBeJJA9oWXoWK5iPRb7J7VgMq3dOFTemPxZRb+wlSC6bdO2Y
cw52v4AjqqEGMQ5T4AIVwt/LPk+hdNy637kwqQqmVsO7biL35Z7cVLd8bNx3e4ip+BG/Ca78wvvR
sZGovzBtSCaDEBLc4nZ8eurvRX/QCNUcNNmtNXqk0Iw1K5MLCwVOIfNNIPo9fX7gGihx/sVMQuEF
QS+1GgX+/8FDPvRjFk7oXjZzffb+q43+OnSCs0XF7azYx/of9TPAJZGdVQvoRsgy3WpSzAHv6WmE
O9jF+erQD4e0XvElqBMpibrL3+TPt6tzHTKqPnvcS7Hy/HGXwwDAy/xsjvclcB0/MEOMoS+5dnZt
+F7T2ElMCQYMYztpdKQRxfIBgg9Lyo+49YKg9JKfn85ZYolOrZ1JQISgga4+d3X/glUdIUz5GDiB
vfABy5sGCedHWqVwbQ0ujvtdvIW4libjW+1QSFFYZyN33k6ZLAiH3AdgaxGGbwE48E0J77X+iY2I
yIBc3scDlaIVY8gKUPSVJbua7CHMx2/Z7idmqpxyojGIW1OpaqvjjTu3O8C08NRDCYCUXJOp+bgs
QRSe7W8WfJpIOkpkDpyCmrH7hI6ztfRhV3FBChygI6oYY7zpGh2vkiRU1JbWciGWrOo6YPpL56nm
0UdAIkBEXeWUhzKNzDAxuEUQPtUAHEv892LFs9NpgCo0QKKvQ00WbEZxbPpDpR1QvxXFjWB0Km5U
0XGa5M9uiKu+530BR6Ly7oCf8MFpSPGNHt6OjjOgZJybXiIaxjFsE+6di8LBEHuBp2mz4kbaE+Kt
hDCuBAEGgT1+qxNWACf7RS/ASBDlhGI3BBmF+Q85bJ909eKWCXYEKYM5AtPClUE6w7ScjKJJigNU
AuCRksweop4v1qDJ7Uh27jAI0neSuhzPm1dpGUtXmqfUlDVfEdMcJ85fL5pnnNSqjBG5qkkEfO0i
2TPwMt649T7HoAey5c6mBcv/VA5uJZYVI3suJXvJV5kN9d0RLM9T9l2ZHNfkpAt4FrQuhAhDkNPu
jJfK9vKZ6pZVD8isE7upUxDcBWJ+xhM2Iyf4k0urPTlzE86ICQd0YKb4PobMq+xH1U8gbXRvIqCO
AeQAJwOgjmNaDJXpsNaGAG6QD077Tnm2JfHj79gpUHgInlzHgb7TqNIhEvINQ8N9TRNUQ0mhtGAV
AztEWNA0JUFYVqML+7pPEBtgd7KeJtal2qfJKQmd2maYnBtEUBFGfagm4Dx9C1VXlnkTqCUBB9PZ
xOZJEyvZQ6fgs1pqtakzzUvCnSl2IvTwRtXHMFm0mv0ootAMudDkV6bMyqjHaOMjYX7MwmejCBo0
PfBGr0lCp+J+R+SG7MFIFIMnARw2iHqbF+PL+1nANKqFDII4MHSup9XOdfWmMVNQEC1KX2RRzqTn
FPQ5Jgt4dPHGPdlAC/nVjHSw8se09x08RjmeR7qRQdZuyZO5CyGJ/t72twq+cHKzBBpWVGcEONZY
7PsYUibaCK1IcwtbF2jRE+lT+lob3t9uw9KANfTvcdC1GWI7ct7DkBPusTTX89fV89jACGiJgXR9
b77NuyuXPcVfnTunkf/5JFgcLq8Un6amHcdaoo8UDw7yWTQzCc6QyQFH4Kn+7e+QiH7Q/eiI1CIU
qztWvUWQfrnWbAcPb9/LLlTlBQCgPPMkpxAwOGo3ea7/xaUQJVDfcTxqXKHYcphjKAGsFxODyIjY
Csvr2WqFak2kHcjdKaig+/O1ynuQ3+i99vxrGF4lNNMNwSySyvUo4NUzKZlYShtYYZz9k5o0eyda
ZZWJeE2zWoSr7NR/iN6vxjIR5kWJDPfx4YPZ9pSgYEydQ3YftBUX7toGvOjCe4Xe5otjv9W80Yf/
TpqN/LbHmA28bAnaqU9TM75dFMudHLXCvazAn25dfaH2ORktIGRhooQx7M2Wk34ZRUpqtrNaGRsM
jlcYgs6hV7V6K/VHpEGwp6+83cFt1x5RHmqbzZBYDUeFYIJ/wmIV//qJQEpADs9AqlyWBbJrgL6N
u3Mo0+fYIJ/084yw4/GPSu+fijqRGqRYte5pdPqH3syi/Fc9YbPJhwBIfX0MYQwuzqw5PTCMTCgj
UWR/Ulnsj23gZKsWYECd+MNz2lcXX/SIm3yQDEyQSxlErygEHlZv5QlkissE0IqpxKOE9GXNmQLG
2JNs91MTTPedIAmsCc2KFCc0tN+Qrhz62MtL98Sgai1BhHUxPnDWLWeaf2F7FXf/fruX7F3NNpEc
Vb9QlukCkPfbXabbBdETEQzCt5TIpcR4ob06q5b8nxwmQmPi5gYAKfT0m71aqLCtmW7198xeUcmC
4dnXLumAEsce+lLh4SY+Uzu7dGnRLk6SKmyXbUec17gURkLDUuhQYQuxU8MIvZ5IUs9VAs2cMHLx
nYuAQiRdcf5ewW5K4qG0JAMYPiVCbgCUX1UpokBXOMwxaNaC0w0RHeoF1hv+8RLFueH47Q7y5+CZ
u0QHadRjhGFJ8jirO43rloiN0uZL9v+ZLxjbFXhIkgkYp5xwH0OjHWPJfpHWqhonopuBpI6T2gBY
3wU/wRa3aR5ffxc2w4S5mUcpM45NIo0EjlHDj32rtgWFe1thkihXkUsqFB3FWrhuByUJ5aQsU6mr
KtHJDAeCib974SXlNw1MkUCKqZ9Jdj/am92kc+x+x6E2DgopyNIcblHKlH8qIBCa6bGhuxX3gd6l
9HsMHfUrYOhc0tc7kNGHa6fGCf8nKB+zVzaQKNcOkHk+hKB2YiUwrHJ8mW2Lc7ByLu9HB0W/xpQi
l3LvuneNfqzz37nrlLy5qaDCYtsOVdNlBJhYAKwfCSC0dTGNDYAOZBy8PnARuhTsRguSNDrlAf3Z
m+Dfnf3JJ1Ckz/XOLJBLYuBmthkt33v2F7VO5ZUflZQVtsgPuTbWkquWAkFQlD8ZHBUjytsif3Qk
jCL6IcxkFVh2WMMygV6CcdrIWFIgmNqUc227qL5zRU36z9EORG+koSNcZFjDgzLiDjzGkBkWzYXB
fLLLvNphCYT6TM7wfNZYF+Stc3/Yj0K+xabfyOT6zXUCk/XRfQgq67fJaTd2ZanzhQFuXYjF3mnz
AuVJlF1u5wPPUlWM6/XRG+gccoGSU6wVzR8Svo24sh7VmN/b7VqIw3WQ+VSb29bKAXjkcx1mAj12
LQHpA4Gw8G5ZZM175pvkhxtS1Arbm+xqWuuDsThWLJWlNcTh6asVFRcwKplVv21MBfsqZXTODg3u
n8pU4pDC66TUIEnCTwIOB7UsE7Y74OMkp1afNQQWIhV5aw3bNZqBKmzGKs6iA1hEIrrVvaiWEGw+
1uOdr4p3GRmsHXA3Y4ZbqtkqliosIRh6adQ4LN8i6vyqd1zdkAbln36Me/D+6mB9KyMqi7ib9i68
IWPv+ADvtLbf8n2gRA83hl44gkoTXhnXW4YBW5d7DwtpaVD2l7T3rfW/bKyB66qQCwPgkGjtyxg+
9lZk3h9TCRlqiIUmg8MshVeVzqUw4qt3kt66ysD36jihUOZuYolhuMs7fQiq2DBJZDZN1Nw1LNDt
hVyBv14uDNpSaRzLtyKVwB0pbST0OQdUlWQ54QTolPgWUmbWiHD9BVUBKi3wUrCmoEEYSA9Kjbvf
pD7eE1dC3cIUZuTv6var2RYq0vJYBGC+EpODWCV40UN5howsnSgJtmibsSKNmL6U0il35UOb1k3o
xOuyYRKgIlntQgd/y+J3StcjGEdclsihx2aAhjt+HtE2yCXqG29T79LDRcPTeg5vlIugHUuysr06
6mpFOm/97U+xZ6+vGV7eo3sIlk/ZD+L7qeIdOHHzQK25msHxBM2nQGUaf/0QkRmwR+5euLMx6Uz/
9GSh5Cn1dz0nZOZjUG7MQDlvoSrxhIqAfXfiDUoLMrAa2dutgVGvUfalWpiUXWCVUjFwBIOapK1A
IbQyUd7P1xlBflreXPPKQqWUGA2OU+y2gC+tWNFGGQaiBEF/JbkWtVKghKoe5+xfFIHa0pJRcguV
ZupnqsCoyhNNbNyNDLo+ofPOv/Tm1DF682CZrTeRsmwVi+R4HvwydAmUvRdxX/Ox2xQIN755CtHC
O1TCXqEvij+aKKTPJUF0VQ1cj08Dg8oa+yq4b4QekXfJPzdogG5IrWz+kYzlztW8rLHqq/I+fu8h
dCiUjGz/g9qjkCzcrsm7M3LRapJbtBQckO34rykq35hKBvllIeidlSy6pNCdH7xGw3UnaiOQaWiT
Kgt+sXvCTiEADatvsaxKYxbyobvxt/HzLFrnnQHrLQ9Zf1ESH02p1Bip6nEga9KR2JF/xoW/RcMU
FHZSL2v1iNq30I//VTY5CkUJAOcs4l5CpGLj7iYOnExkhzRfGQ0EUYd2AJN9yCzSWO3/3FxSmdU3
bgX0C985zFwFlFX/42SyfJ7SuWqT9ldz7TWdicaNHGZ2vrymAUKYr+MCa3fZdLmQTeSQjRGlIGKv
6+HeifmABlih5r1XjqT+/IlrN/70FgQvIWC48xcvNrgnOBTFMW+3SXQrnKrq5ZdlyihNXXjsATpz
vd22mxhKXijPe/bEpZfqgCUY2kPi/NDw1MKkJA5P0yTxZH9Apk4lX4rUlDY5leH6oYV6TLH4+gFc
kFicUs+XWeKqIkwRog7KwsX9n2AlaXBzXwfwwZ05CDbTdpvzZ8LcH1SXV8W1+9uhrpQ6VMh1NHi8
g/klfq9WX4X7O9Vky9iFsNrq0VDVV2mrUqnofMcAy0Y7Dv9u2o6DMfKrEKK1k8XhrzmQLdachDUW
H8bJXzdDIKLOaku8wXugyoQinnA3Y5A52BEFSHEywmakQFLhnJ9WvHF8tw0/Jn/jwJPoq7DyqPoJ
BcdI5oFrDWApYH1hFSHx7ABgo34sR2083TEgoD9iplAfbHcHP2ueotIeKan+Xh2JLsXLs/aivEUZ
G/OX8nB83oEnx0kCr5fAL2nwCcXIEIOU2JTWggizeVLLS16l2WhAaTnC0IquItCpmHzVklN2NXNS
onoBBFyDZbsoH+HdmhXPnSN3hHeyDUx44lhOr7wzYE9DS8nWFyaZrn8uk5BqcRFdAxSap16rxF3h
uCg7ifF/sXHJj7stKfrn0/o1Qia8qVl4AFeHLoYYYho2hIRr4YcJOU7oDZGbkoLh6XDX/YWUqtu0
C0kfDF71ySc7453sJfe4QvwnWnxMYXlpnSMkc09aLtMByffLjjmZPGY74AGasNXyUdY78gGDfmL/
srTOiApl3IaQT5d9QJa6/wXolGoxVcDMQ80N3DjpKz/esCqyey2oNOyG5SwwpcPhgwsIbgOrsQa7
K9gEQVvoUPQiYla5XNTf27Yuba8X3HHEAOD6Et5MXHHfPAP+qWsvU74005r+rVFkiGnwk6fPm6tW
2iJmhEVT8596AzGvKe66JoG6WMBxFRgS0rao3Syy71105lFJscWcSiHZhyx/l52E+ej6f6pCKcCJ
V8lwD0fAnrUTpe0+cZkk0WMmS9pEpX/Y7WmLx7GEqIyIxPgGKy2Sln20GZ1ODqd/+XS0mNaOufEf
LraDrJ+/+3VMolwXtUdBaEFgONc4YAKIKp4Fckv4HOIfMFWNE7C86HXcHVDB1NBA8cRWRP9vli6D
46Da1Xz9ftrIO6UXjDN7HBX4UTtm04b65swAEQgfg7MSVbxAKUUcozE5dPz1Q9CsoyoxEb6Xj4Ch
3AXNDP4x+HKF7s/A79vWfKxE9FGvTr0dNXNJ4yHYUpy/GjPuoajF95/ubWH0+ASec7ocpLUvqj0J
4tiXuiImtR0S6goyxVbrBoys7xTq7Ty2ZWhU23Y8SEpA4ewTBLwq11ybEJKiNiEbXmqlcVePldhS
BmBlBu32QvUUzOhjDbmHXh/RQvjMxVQCn/cHJ5snSOjHUWyt6eM7TDLk+zI0ZNRRKCk270xyd2RN
Z5ixvbwNsHq5QdzlVriibB4ON7Imb0BrzaW8MmG+GQwz3DQNeK533UHQvJUCgh0SVV6Fp1UsvqZL
tKArwCc2h/WNozvZXF0vRrBIWr9tmHZna7Cn3GgPE5/z2+QrX9DOfs7ZWpiaKoUoxkCQDDQXnNHh
uhEwQc8yakYK5pMtfnyamqdorxZcEeU4rFlU21EHr+/guabUJ6S0Dk87uqfZWSN/5tsgwggxGwDd
Du74wCBF5nT0YnO0k3Y9feYiaUmdjNPHeR9L/M0rT0C9Cd4wQssTQCzcRFmPmUEa22OcmbRoZSUA
ArcU8RepxuXVzv+woBXFKkvMbZbAC+gjYBChLJtmdFDHAI+LUejpYZyjVQSd1SFUXEguub8RNnOr
q/RGUS6JnYnOnc/41Rfb8V+ifxZ1bjjUCfIz/2NEsFU7OApg57FrjieO+9Zve347maEMX8BQA0G2
oOc91TWrN7tFqLr6oh7ZT2bPVagZsQqgU6Bn0ak4dOVgUS0j4NslJMre9OD4rnmbVOJNDgpCXupg
AUpxDpIvcr+I56U4zJWHZIwkTTRst6I0X0K6U6aICGATCtfzTuUhABtONk0mLhId48YV9ceECw6g
5yVC8W/NIZ5JhwYvon8dJoG5/ZMjDLb5rFgeokw2StBHpJ/vMh7MsDr4A4dDECD/sI6NaCUObkhT
T+l+O1MxOh/MUMnwVOaDwaebK1e1ExDIPRKWoW+wLgs+aHQ9xC/dgkqcYTSeYO/KgUkavyvVlriH
/tgY1hjtjuNzNzN/UEFfVtovQ8ZUQEWvw14sXYPAAEfCOGynrgGNrMwCCv2KE8O0pGvc/lWGKKrQ
DRIwLJCyrzQBWkCQn1bI15XuX0yZ/vw6wjgiJCrLSpHh71CGKRzIOAj2cV92tBUa6eEgpW2onpIz
9hgLtX366HiLimSXJBtsxxVKiGbHAVyTkDGpNKgimykdnvdIIhM0YtGcQpD2GNXeUj7xGkMw7lxA
3kBTcR3lqDdKHqmhG+NnzJmBrQzN2SWV2UwaEy9xxkrWO3LneAUl7C22sa73qggp5QDpyvEgQHK2
0Tkg4Gx6aEXbgfrwfcoqaLtiP7pZ+Las0ns0LFBt5kFk7s97WmfRGh/MlFsBJkZ6lN2x5nZsLmOH
BVwwbelwegxw6iNr9gdMcGL3TloReEyrC9NBXh21cy1EiY7Eu9QoM5YfMCsw55/FIulnJN38gJzB
vCYEaKSADkOIpPtHEyGly/ywsvpWB6PYP0hK20C165KsJawU6J0D65jdAPPibBcEschgr4Z0drrO
VB+rPC/nT7eJpkSSPXTiAb8YdlkxhZsBAyCK7IOAQJ2OLuI+/aZhAtMntdDWJrSS/gNxJENavKBL
ODiq3hmUmYmaDXvrbTg3POzmB5m1lni+PTkrf0NEHvv583D+5qe6BcAIUt13gPrQdO8XwdIm3WcQ
eevFnsnG44s747uskK1WqDIA0O7sAeQGC/XCS4I2ykdw7VTFlw1h0yW87hCDrnyoG5Q5Dz9L+0AJ
qcqlWZjSS57n9liYA1idw5BVAsM+I/jD3huf8SvaoEZyvAA6QyBUH6FGOL8FOLLpFQfscS+VCm8t
OiK/o1DZzptdXgdj5ItiRmtk0XxqmAodBFg8wUmCdq8Qhg9R9SudQvpSyBP7OetFy6I48NpAtcVk
5fZnkIBOGxssvo1oVKjvgb/hp42d4ggm723+huOagHO8cWbE3WDcFF1825xv7v+pobUJuezMZIfN
IURLJpWmikXTJZll6+/H5Dt9lUV+XcWKmknrrMRmhe3SeJ2FPixqST44XMupZ4H16L2xVjgQi+V5
KQ6buxOWQP7fO6+1ubav17ahWs3JURR3g8rloNjOh5G42TBNFp9wRCRSsrnbsvMJ91JZ2oVCtG/j
xQ7ZPbtv4jCsyaGuvouBzi8Io05ruVJOLj7KJEY5zpGV9ALosiXDajH4Hq4G+KZed4cjd0lnXfGS
IuxRNYqyuGwifKVSzrKjaJm+RhI85Qn368XUUNxNfMMnBItXTddwmgSqY2sJigZt/vCDc/flfEVU
61MlCftgzN7hZrCww/4wiVWRBHlHdMUWjCvU343R1BwSwOs3npupTOICh2fgpzcPtQWGTXiLEFwT
gV8Nyyvk79ialgBMezVJuNSUcPiFi1IT9VqOd6p36s37PdwEgOAhmdMovZCHvO6ieg0CVNC+C745
n65q2GI49vDQ/QPsmxlT5ip4g5NIZjsYHlaGcR91B7r6uHKPBdIDCx7oBbZPmPIi+RIkOOF286wK
sWy9AHNx1WqUBDscf1CpjUfaxl+Uy2HLQ+aUqVbtsLzTPH/q69B6mRL/ykscUeP3GnVk7+srppTc
mgulvbQM/zKMdAeFWmBtUoDm4cOccNiAkPNSomyKHtIpxTrpxCss+7iG7nls49GvtgBolsEWqgTf
KUH5NMN42VE/RPuE5jQij3EHEFwj6ZZUr9O0j2/xylG6CEF7sETPQ9O0gE0QrmMeIX7gIXcukQs6
TcxPGmAydTP2AE9P/q/HXXe2M3O9ISGLYpiQ+osS8KX+2JvJtWFbIY1hA2JyG2YhczjrJ0rycE+B
40usd/RFwfSuo8VfEzf0WIw4g4H59dj0QY4uKUriuq4DDWYblHtrHTpK1rCqnPAz+TY3TnUIF7CR
sH9VROCaf5uyhkHJMUikRdwNyE51Inas8UkILl+Plnt3ZPQ1j2xbrOvStusd5b6pU5UjOYub403S
AjQrH9MSO8XQv119mm4vukuzwAvcnljyQMOsk1oLlyMLBng+k9Clb+ToR6T0YWddCG4BKshWyyn1
hwzXRIecORY0AuaG6+4VzaUQRlH3tl25ELOan+FGvy0yezNdVmlEWdFwwdfcie/1mvFenflCOgZA
rT/V/MIbWKD8wqY4s0eNtWQS7gVSMWI2tvQdeDhjcv7mLgjyxz7fjN7mKE7KowkFoNUrCmN0tiN9
kGAZ1nPrSapQSrw/zc0LkYklVc2vpKCqyxQqpp/CcX6zXhaqXhQNXCSMEWykW8nZ3+BuY6vVV8SZ
I1t2CD+dQwMylFRSEgsbycOZF5JGeUJ5gEqXCjqLQHkwB8z0S22vB3HjqOnTayh+lweX2pKul/s1
eYATnX0or1Eu7bRH5Rw4VM+EusFYix5lEboupNHXVbIy4j0B4f74Y4aEdA3BHT/PaVZ6rENnnc1d
yiQE9OmGSsOt/5FPIGsGqx7K7IaHI9ConlF8K4Q5IApW4guMxxTkERwDDqMctTp9alfB+nKC0S/N
5BAp5XWMm1ESnH7y3nGPd4SWmZ+WN9PjoStnuqIdhIj/7yIUs/6FIuZ3VeElG8MeoksuQYPLgXe/
4KZotAmrW0h0Cn67/pon1V3EMzOTYv+LitroZOvkibTsogiAdQ5JAvOQKyrGWtC8vCBsAr1KVpvQ
r2ePemAiiklAI+1kcLPk7IP1AIjrbVs1E8u7RbfxYYRfwnyb8Yq+YbBz/odC3Xq3DxtqDr0O3G3N
yhEDmkzXp+KzOlwrinhn6xlgzEkYPHNmIY54onJQ+zWnQqzV1KU7v+addV4sVYuqIhos46RJspoO
FCs7Z5WLfTNwgCQKoL7o35taQeuqv+n1sckAWzPXhxd35nurKb6CZfgJ1W4EycffJ18yspHjmZ3U
qDXl1owo9/c+NwsjIZ5FP7qpL4GRChFY2jjy8Et/yGgcHJ30f0XlNwmwi87UfiAk/7s8tjF82PMZ
Xp98gi9WoDk+tF5ieFlZTT7/9L6hVE+7TjBOIMwSavmAqzBRa2LAWKSXfsl3UQYxH/lxIqHSCNlq
Ej4t/8Aje2GVdR4jZ1u3WjBLS1MAhOUMC7D/L7UZddfY3E3Epq58nIKrplyJd6mUFnZRp7nacaY2
u1yi2KjMsjJm7V4OKdj15c5Mgzf9GxgWRto+I1D0PYlEGk6/UhRK5kRAw6PRdMzE0GqaSUD2KPrO
pz3wX8JOLN0cep+BL+/DgZpoEJVcBIXu7meu1Lok9zCvA993Eg2SYv6vWJ+OXZaj44MqUJiYbO6K
r59pQAqoeLRks+nKnqJD+iOsu5cREC2HHhzYXKxVbsG+LUBqlcvq68CyIvWTEySyyGQh7oAST/4e
VRc4XguLZPIfGauVThpjtNYzx4VSwO5Xo5foYFG2/dequS8/3hzOnctbDQOT+y6REoTyRAL06HOu
uHBnJjvNL7h+i5JHZat1PlHN0KX+UXTv02CiEn4OoGdAQEOvGn1IoCl8B0RZSFxidkq0OLXOuA9M
hKmoVqaZmT+mCVq+/bLMEwy0nw9ZommNISg7GpoS/b9vbVC+mufnMv3MABUfw0jJB2OtzV2JNQ+T
ePsbWT7kaZf1DBCh16FGObozbOhlUvkoJ/iJFVTPpjc11A3HQfz3tQ+UjBS9YPhGfG+vS5iXrbBs
9hHWcoJmNXsbNej7dytfV3wEskuZECYCqOGadm5KlqrZvKCLgPwy9dnaJk1QJfcOBjC2oPUtCg+s
FEW9bkll9WSb3bDG3XFr2cWjh4hwimQHkRybBmjZo8Nm/ggesk6p5HnNNDWEUXg67I8x5LBu7q14
Xu5XvcWRsYaw5X5xBvosuQ9989Y/sWyOSSSqv0NIznbAdJkv8hF8mxgFeBQaGtizN35yRNjLEo8/
KshpqELfZZmtJBFpL22pWdLzJ2M+oJjyr3P7MLyAkq4gPTRM0bh11wjYsDRk9s21eABODkQ1EMlh
LggeHORg9LXjkgaQ0ENQ0uRGzZ40Bd+YSNn8KG3WSuDIEw/jqV0QD/ePp+LF+tA4mvYg/x2HV+8A
dZ5TrLkt+qugU/4IbEWT0n3I/lHhu7j6XuSEG4GVZKlE8hh36wyFiBPIE9shdUfrBddMWiF1HTFs
VgbkX4XrySIluf4zzF3L1674stvCTDvt2mw11Sc6SFzj+eBvai9QSOwcW+trbjyhvk11jXKK6RRX
Em+AI9CJYzoQclTEf99Cwr7kBL5E4IaLT88CSaSM5cKJhweiwN/B8h8yQcO4FkokAIwbXxc3ua3k
k/5W6BeJRUKKQHwWb72oMFAsVCf68C2JJ8TtMVfbfzYBKQUtMMYm5TM8huhxPFjBnkWMFftrIlt7
kpv4pnU57YNjQwJub7EgnzVDRYcWDT/7lZR2QkWQbRW+TRTPwLWQxcfV5+RpD75evhSQzVCpyFHl
uWE3kPorPwF+b2+B/oWzAhg1QowJheUrKbtMppsaPVpej7vSOZbd3Ijpq4mLF0HPOdPZqpozjjQz
oHfh707szBXIjElThXXcpG+9HHDJffM5BXNNfUFVu1CeEq9KcqWwc9s9GgOrVDdpR1khFCsAs98C
sc/Z7Jp37LUze2nC3Ak0OvxlXTCawhE6z2fSxqTdRwEVYZNjGJYrGNsqX51r8js5lcDQoGODUWIU
0yaHD5SEp8R9PRYsNCnD0VMjITjYiCO0h3uD+uNIk2QbmjRy4826IgTK1fOWAfbZZJjQ1dkc1V+4
MdRyZ8mxl50mTstb5Fnhfh6a//fqGXTt/ZrmS5GN+ovb64PRe1g9qMQwhiGmqnQIXNEeCiOJrGk2
99TABZbLDNH5/tkWG1U3S+NN9KQRAN9vdZxVzzl3dU5UlFvcZZ3PdlcqBchFlcw9Ba/KQ26trvUK
YWbZx05gLDrFztmZHVP+LoUWvFGxsR5C4n+BXesn5l2cA+HAhbakEobRBJ0RNCCKVTZIFGrkKSjT
36BXBKE3TQI59yetpUbq8/4spgnIjHm40kAKWXx/U4Ygxxr5/W2GGXThLfSXjaqYq1ykvaa73CnG
GZnEgfUlMYBhB1mjRCtbn/L4AdzxCFIwV/y/Ec910V6qAnZcjM1krfinVASNRioavIUDbHpxUsQ+
xUd86kVjqI2ssdErkCJN58gOvKSGREKUUQ6je6lVxMqUwua/cO5sAaJ0wevv6fpp1c4RtE8zgPRL
H2rf9mVsRCUkOV0Pg/vOBJ4MiTF5nRsyRwi00/LZaB71bX7NgL0y9MR0tv+uP1YNNyLxIks/R4Ov
go+SUNf6BCzcVHItZmyYWA+eo4rRy7JJqn3gqeSRHSMM9+jxV+U9Lbv8ivCVZtti+IHpcPkazuZr
ElzAb97I/rf7oJddLf8eN0/N0Qg1ytzTUkTrqWdPNjErVj/x/Rj40BkeV7aySRlVnmUMwnv+IwMo
Ibey/XxDQUnrXar5cIE7xBDwK2VNniusV/iL5W/5E9Psv5kEwTHxpX+sP1YOptAtRsjp/58EEdb+
3sUVgZCqZVS3hhagAdxYyEf4djdDoQToaLICscrP3LuiiCpOPSPa6F7/HpRZex8s5giUhSgb+C5N
BVic4TAmmXMFqnbJ4I4a1SpZHvlkz13onJmE/Ld+PxDhHN/uZEVQ/ZixScevaEiAz8XiJ6pe9Q93
MRCWxmNDepLrkoGbq3/LRZByHNSRxeKfG1T3f6j/Ys2lFq2cIGrbjK2pHjcUt/aVh8t/ea2WhccU
IvbMT1xTR+aVum70XfggHoTomKhlFzzCxn2qBzYSRAsX4gfnREaAjworWwK2uTUijmHatokdsDTO
YbG1BjXnAtQbaJTkKkJAR/FTj+niXkNm/9dMGe9RcEfuvTG8N55x8S30kGs9VMRFXzUM7EN9gWzm
DXhkWLFLhzg060TSG4rIJ5gAAbIkcf1WTQBxqxXORQEhzjdC/642KDdBUWZh63sd4aYfrcY3KA5U
j2AY3FQ2ArRUml0xzEpRlnbHXmb5tUmtMWPhuzuXEAPDla4O3VF22KfqGr+UW1aIvTGcz32gN9Ae
uEgHlKU6dnRiUNYThkFqRatMRPcJiKUCp72moScx1i7AnODkNAcpYWD8kONV4tyiqcGpgnyC8Pk2
pfsqiXREoG+8cEIvsB/Yzy6ZBhnQvwIqOpbspvp90hQ/SVFIow1vXCBFviBE55QxA49GdQzouT3c
zk2kbq4a1puhlpJ/dJYwKSWJ7329Q3dJTlUhbrDm+07/vOJJTDGFaHmFnFRFc3hRQQ26y2u/85RD
/n0dizeWjkQlXID1ZdzmDtucE+3dba3Djt7MThZKF1desQFex9XxHbrx2syXrZzFecULXcBLdaZN
w28kidQmtQMP8cSECKFreuVibCvWisVOm0idL5LX+gmbpC7ByntSGMPYNyUDK377ZxbiWtF42fbC
dP4JKmU1LGcWuwHVi4P7x8thSQw8VXgSd0JnPXmCj6QJz7EFdKjpmPqKc+N3dk9nhZHykrtOAVEM
S7m4ykDrfP0T1cwwdwtAjB7C7oU3GM/yIKu1PRNpINCtIm90oUWQsUKZk63ZTdqmtQdZ7tSK5jmR
isKIuaGqNEKMzjY4LAOGUHRX1i1F0bs/JKY5r/4qzzFWnM/mBb/LfzZe5PQ+N18bgehdWHW/041q
rYCJcKn6U0m1d/tOULXn4Rp/D0GMxDSoFg3LwVzxHllXyY80e+ncvaYIXUTVUW21aJoyQKd7fdA+
sJxQ8nmCT0p2/dLyTb1eaFNnS+M4yBB1rSb+zpi7UZt5gKxRMam6zoitQhDfaCBwtRHFSJwAcCgk
w5ZX16ecAqsUBrKmtH6F7eQIpAEAuXuomz1aeR1q6sCX2dqU24f5kUrHWPXv4ysINbs1h2+Rnaqo
4XW7M/+QHOtSHxuH4c3vY8XjqrTYC1swQam2AafqvxLxhQemGpmTEAjnyGzH8UFkmOj2id+x/h4h
7njy4vuASd9Held1XHBb4U6I+5GjAumtTYkW6WglmupxskpHv+C912MNF2lqOsSb/gb5UsddN/Eg
eS/466Ld5YIBHy2cDCEokP4JqNl3VuaETuXU7D0msigL5SkRHOCDyeyQ7jkYPVkFFv9pJ+xbtcwt
CdoDcakyvGvVXH8JydlDzaQP9Q0QM0/aIIVAjGBd0uh1/mce1q0erKqrAQuiXkMhyDte8PJrjvOo
gqxe0lRcMUpMnEjGbIhbqy5yFoFbPd1sgkAvu695zTzZcTsps0l2WDs/JUELuW1N7FUuTRVjztB8
IiU71LnIMD3+shdBgzz/1vXwD/R2Zk1x4q49lzHjTjlVYpPNa6CBeQP/IxuRBRv3MfwrMFNiCVMx
M5zRWC91aFAhj85B+DVQYJuCEtMr7KMaM/YSCGKIZSe2ow58+3aHk884K/3qN6+AWaGXsGuUxqHa
keZ3apPMEUVbgdpNiqbAm8n6SfRpNZj/AE+PHej13SaANLkhysHX/RNgH1oCa6TA9kOyOmITA2LS
hAf++qCqHMTc0m/SAKw61pUoxqkqwChbbLX4EB1ThXs1XgwBPp0uXAYgZIMMwmwzWCDNSSac/Q3W
lkkweu6MQRTWlAu2OmaR74L4AaSGpJJAGn9bqnoHoJ2rH9ng9N969MQAiAOAzQs+RTMAAAGvmHfv
wL8KF38RUSoXF/oyL+2HkmnZ/FFEW8xfiAzMbUresqxVa8KvtAMioeUnZ5CBm6+WQ68sbFuSphjI
ePEFeLZBMZ8D56/bZ61wzlCLzR+wW12sK59vag1Ys34vXkY/Dho58itSAlPCrw+7fjw7SQSEr6DE
kboSNXrpoyRxxWpwiUCG3wG6L8YGYWi/BL8NMn1AN/ZlJAgzRa8X1Sd+niPBZppRd8Nf0I/nmZig
aTX1NqaRl6Woxtp2es3yrxhebzT1iWOca7BZr+ene6jOUFpcSrbbbyUxDWqq7tU8o5D0pLhsCWME
ENGUPaVRXvwVWxOPgj39exUYuzdmsby9yro02eqPsBGxbp0li7w4YpT1lX70oeVhHPWSaRDhaPjE
sTFPDlIknmbxs5W3w1Ix+OjPviyq+ZDY8llDr51qaUlq0EL8ZJ9vOgdb+JxZ3wiL6hzHxzckAAR/
CUhT/cZ4aTB8wx93Mp418cdY4uWFulilMWgjeH5Cg/0bNfJeMc/IAd/Z63O7ieyj4jxaw71js3Zo
MjD9WivfpZis5KGkH/Sn0nExLLnP0uFTctiZIFXf1nh83z9+CShXKrfPNV7Pk6CiEyolPwBiqKtX
ytJLxNg2a1dijnQJBLJPYruVnA8/+UOszcLwK4zUa7FmXQuHf+OOxTVuk1xJdpqvM03fpwYc7f1Y
m/xcQdVJ7H3gFG/p6aU/R5sm1O+RwetFQ3dOVLk1gKZQLvYGxMTQZv7oMu0yuIlrfo5aFC0bP3pR
HAK5Pm5bfyyQ1tdupYR5NdlA2RFp8t5IUWaDipFQPY5q8BpwR1NE/ElhkUQEI1lk++n7gSqQqUNu
TedMFJFkYnLAVcLrKtY/gDW280F6RJ+7lX5zqD+NynxRnojq+xw8nUfv9DqpD5QaFn9LMTb+jnLr
y706pqSy1Tzqfcs63Cl13jROuACYAVT7ax40PT4YeElUNjTkCcom2s90TWzG7loFLNreFvFNVygA
XZ6MuXM1isg8140UovL3ANT5wdtwQDZTg4X9I+dOLfIRxwNTnKe6kLuAQXmHRgD3QKwMJbxXcqL4
bwgVYKbpJ6MkorvTfTceBDL+igKXYd2z0VwHCB4wpt1YBe71aCQcuoxvr4gZsU137tzB+6H0cv2C
qhrNf4CFVDQGUTPQnqKuufJ1bQu3ix86Uzlem/Qp9BE3tiIA1IUJEBmmS5gvWo/G2qBkdOoiJCfW
C4T4c87Ul8ggvAx2o//khxRBeR/gSJKmgzfS6mDVHCwxZCBMElPSrRnvqvhIGL+UuynAe571aFcp
OOEu5zEi+lgZ/sidYILVXVSql4EVsVs9nD7IeQuk/kXrH/1kEyMok1XzAv36P29nmetY4V5LO5Pr
dePK/h9lIOh7Gk1UH/2RklaJz3uLnvLcKmr8GlY+YqATLQw6FHtfeuFkjXFejegQC0ce65RD8zh4
FMu6lfZqoXtLMt/7YcvwxBj8ruVotSkztogXMG2AMxeFPtaphfm8atBYb/YHSMzIq8R4KbEOwFJn
flr0wnhE4gktR+6p9GNZjGLJhv7+q210QGthLTa3FTrzOr+1Y6jKRmt1Cm0sUGsAAYYeTLzEg+UA
0d9rEfdzP+95zxCfJZdmnzSokH1Udf9wyBXavFbFkSFOxHiWY86ot7vKpIiC+APyaOzd52msIWeZ
JyXpGb9aB3cYNuGfGn967Jf9cyYTDrfrs5N+70WYbeBOJguxgfC6rgo8XFSr0E28SBT3nohOEtkq
WdNYrSmM72kTM8QVuwJXOS5711TOiDD6liZAH3V8UI9OTYaRdypaRnS9wWiShmWNZU8jp1Uyls0I
gw1pl3++60krp10fIp92JDuiY7StoVcxe7T4EflTMqOkt9IZo8QJZQf1xZA/f34W9WVXkDpYy7hA
borwzg1EoiI86ER/hnJF07SLAb9woPRgPr/axtALkKrQdzXiUNS2X5WseM0IM2RsZQ08GEJg3sGF
pe7pn2mkxs8oKCWosBPRmeNJcwewwlPEgLZUNlqy964NpB11iq1Lrjx2RiFuiIEw+K9qD5fzdYA6
dn548S3BFErW52ayJJfX0XqWjBvLtS+vhvts0NBBMJvpNz12usmIbL2eLecjSFCuK0bzaQlILGA8
MhUcsjXA9LJrg10a8CNdsFN+vQ62S2QWTqtOSIb6eXWvXxU48NWiD3wVcXdpV7JV4Ji7fGCW0dZR
7sJ+s22U4aNCQrBVYMQmU0unZutkIcedLmFGuGMx5rHczpFOk+iVnZCIlwU4GIQOw7dF3Stfljeq
N6mTjibFdS0XKElIVJmqpDLJXWIqVC8M+/lEUXHw/LwaqQRfoAVboRP5feJPmryZ9E6JlfT8B5KH
L3iQOWiu492NdkyhVR51PdqE78u/XAhA81kMIncKWpiSH0U3O8V4qsFJAGt45d05ZH6p9qANTZ3q
THXQ5aotaB6pmk8Kr4iqC7QBInrDI3bwGZWOhOXPYHIuJ8I5nmqrboGk9bkXtk/EFhjSMmm6FvmY
ytInDGK81k4s11K5gpxPNe869cei+SEBER9X9iPW2bCpVETS37LHJqGL+a54aYNmBzp7KByPRaHm
jKSmlg7sGTzIj/BnkVMs6zhDhyUgxg6M4xM8YDZ9s7siOFrXPZ1/r66DPEIbeoV5JMgGg04o4Kj/
3pOMUMniDewcV1YWHSq42FslBijZDMNmUEn+XNx3/P/+EVTwDaniLaAQjZl24BCL0bUO382YMQTg
61nWhS8T9eZrcfOj+TI5iUWfF1GKRcDRQs6wEzOWd9JFqaPtQs64QNwbkdSzkhesT9J3uWSDRmpD
eNj2EOGNsOs3O03qQe+tsFg+Yd6BOXh4le5oewuqHCZPxIx0sfcnvoJs3RPdCLA8vJesAQxfO+f8
0KC5wiovL+T8IBzyIF5tu2EnmZsRIEqqlR8yDbMPDDivw6aZgfAdt4vCWPzdiMOwScoqdmR90JLJ
qU6XCQ6QMBiucG5sg+dv5N0eOTJh5py5De5QS9bP2JCRp+AGniUwbP8pRGYKpmyvY0XZCoZibvD8
Hdr9/J9Glj53FDimGbjBlBVvtdPFEwSMQN1tpZ6W2TGM1sVNMDRRWtWXkQK6Xie0fik/B7t2zk76
qoP5fponINT9PqQ57yU5yLh7EUAp21AO2wFFb6VX/3vR82xZggwGHLe9MvvojyFBJK1/AqLrSk7u
ASpOj/d3YpoXG+9tqF+n0+cH76u9KMNq1bHICx3k/8hf7zzBQuCvWkxLJ2AA04HgOTdRdD9kGc0n
GUI3PWIIbuKeIPQgmIVVWS1OU1oXbYbMWdFdt1yGm76WduatyP1QK89feD3M/3ynE0bi6VWlBtTR
Iqg/UWPXWIyYDmJHYa1vQOI2ikMLaHezkM1vIo9Q5B85G95oOBu0TC2AzuLG4JRoTiZe4nHku9F1
Of27QBHNYMsj2zCImOBDz95dlUEgevOJgob7ZuSStsnbVxsh/LlpWiwouuMYJUy4VvqiiDW4MHTx
gBDLZHysQyDhuLVKzJgggcvxemXtOzNEbzCwkV1HhIWwU4PjbmE6YcYzZzJxKYmChbE1rvbwjhzP
WGPa+KayPhn/rE5aN7B4SPjccNgyXhlW42GkRCymdpdlUsoT5zLIAh2f/dYYIrZ0y6f9VWx3l05G
QaPQjX9W/kGU2FQ2yeDoDpcAUhSKzzadWInpAFd4LsAG2279JczECoyotkntVU2v5J5Hw19A5B97
GZmj0xC07FTTICtw5dyqkFW5B1ZFqYxYbb+1IuL52z369P+d/QJRi4cXzRP4hyI9c0mzfW80tOgz
NjSYViHCQGa0RQWve403GHpGAORNDx+JlXVQ5kQHneqQjiHfVViS5lYWfYvPqv2WR0ytw593Ro9k
Hc6r8+6QX/WgcPbEOk6xn0VsNeGIu+y+V02LG8xgD4vgHWtuedyW493pzaKAeUQgK9DmYZw+nxKz
IgoQEYuko8nDA2LgvB+PdtHAcJ7nB5wz5hD/pC8wKJwHOt8Fs6RogC/2TNWn4KxxKj/Ieq1LRlgQ
WW0gRis5SdRa8oaRLY8kzsgKZBryqE309FV0oRmOE7NiG/oEXcRHyilA3G52qT3u21e9lkIleCyJ
HKjbKLNfDwtgyKEK3czr9VoZOICKT3Hi4DO/3rcUJauMXHE9+uJkW2Eebn5VG++TlKxLCbG1qBbB
G5qtpRD4fJ/2Ex3FAL8j1VeGM9tSPNjeR/5zq1Q4jSOmtmYoZF2F01MvhUOYrW/6yjqLzkLQ2owd
WQmhk+EmqOTNProwIFRselymM8gZXaGDigUe2LE+P4b28Vy9NrUKMnqVa7GWp4uYYRGmIEurlZGm
ShSbAG8aX9e/oLMPXdTUKGx+2t69VaXtRUM+MBJTQoOuSYDdTqz2F625XYIpzdYjxAPxKzIVBXjU
FAjsChdi7jy4YjoAKVfL/0Vay26vzywtcCpLgsJ6dst+vWIo0c6VtoYInASpxDmBvPme7/4yOfze
QaDenv4E9Q/7Gb36d8FX4aFG8AeR14Vs/ZuZsswUv9pjGIOb0CeUzIszKmuvEyUnck7bTSNegAdG
2vyczWR52kOV0YljNH6TPa69zGJGr6Xb02fPBHgdRfJ5TADf2fsFoxemStv2Wx7mEIwR8cO23euJ
2mL8hiLWa+DFhFx2a83o7eAJN/Y01WKri+S6s0n/wqAOGderN2OdOlyHZjCLp7Rk882c45hmjier
A9bgAoxqq9LdUjNbslHzIapnTo24diCkqpqd5xQW2ZzA/eCIFPpYRfklZwf7EnDinvsiIrtlr5NG
NGtj+DHbhpgNXucRI42cFCJ5smjRWwHm7kjCTLWlz9Fd15lzo/fRjOIvWw64Hsw0HYBLa99B2DhT
sRZ5d8P+n07pYUduReOUKitrQ+Tv8BxfYeOKTGMZF0MhsfKvmTEhZQ6hkF8EOIHd5ZpHttU/435K
igNAKygJnh78Psd8Zd4tFdxZ0fv6g8zsFJI0xkSBffsTm2LfKfoOB5AoB2Jt0/TK3rCC46VrrSAQ
uhl5G7KcbYcMKStwiuWHYmS/s2ct61sWzznlgbmblX9sGEvEbuesUcTfIGEsv7EQNjxumPk18Tkq
HRGCwNPfMv9CrZeFp1UBmw2Br4bP4b4IlVGuaBObxsLYlxuEx2gIKOu9mQqmznkOL5dtA6CnsrI1
9hZB+55+8xLKIlPH21QGhUZKYV37ZaX4swq5Xl7V2apRZKltcW4fya3pd89MD2giCc5bG2dZupQW
EQfqm8BUYGK+Wvcc1gZsy8NMMqaVS+/tUI3TUUcPI0BTHpIRt/RQ5R+3HHs9BT7wdbQ/9dPqigvF
TiFJ+XiD6XaWlmCDZSLP8H3NFqBOJdrcmANoScyNU3dehPXcMfn19eljQIrqT7/pd2jof56WJt9k
Fgl/byFFVPhyAgXBluAtbjhsYDV9fmeZP/+Ib6h4wYiSZJWtNsRLe6m3YfJ3Wj+8um6SwHY73EuX
pbIlg/04xaWnc17g2XscMyu1D0HC+ehR+JO7D4BjCLt9DW33LV7LckVvjreoB1Wzh3QBZJF2RIcw
exkSCciuiZBl2WoVJB5CaqAgOIQIRsFhPCtge6/afwiv2/jO99ySOIv6rUTb4sJVqAaj5gAa9o/0
b2x9sIwSPZrk/S/DBN55886QIKdWQ7uPNrY2m0OUC31IkMjlhk3VFghNGk5YLIHxLZ/0GtyjvXMM
i5qVDW9MY4aqDnSdhOKDgk+nZ7KbM13Rb/pNccCdxO/c7HZejPcfLRWYV9uvuy6FB8LipZyvDk3c
f9uIaQtMEdciHhVwL3dMyWHWbJRtM+CWdRSiP6oyWZ873D02sXhbFThfINKiJPFAMiKRk8JqYOWZ
RRKJcszgBQRh/8GW7cQBTlU/7yDBdox6PntbxdAxvLRqd47F67VYFyDX7pPZQDESsaydGSvVzlXm
ZRRCYY2M/+/bBlDwhzWrT1W0e0N3ztiVXs+Vh4SLZzpKbR6Tr8aS8A58yAvvUHX53DviGkCkNy5C
Kg2MG7hJf/RBaROsigR5D09c/7qarrO2R7iX+GxjAd1ZevZ4VV1trptZNFcOGeYgpoHjMk3eZwh6
qZagY9ggOuhnW5ct8TpgZkA8d76A/qL2dOG5j+l61+kaszOfo1pPMv3ziJJ2fzoWE7zG0hffHDvl
ZIjtYhgkD4uCqrbnAOTsMuQx7k3BP2Vh7nUI/2aclAWr6yxK23SUohorLp3xLUdVXMztNwdRv/yx
EeclEBzSAr1okGuL4vsL1FmyXTC55JD1FzHJQ4uIY3mr+5kAwOG0vZp165p4zqMC4AmjkI1zjPTu
0vzPJu15XbmeLIDRooBJwQyw/twx/+RtfzJn7/b85V53jKTFgy5tGsit8PDouqR+bzXZxdNYY8tg
13Wwf7s0xptpt9OdcX5KDSJmGTRYyAZVGpgilW2Do0XJru21JSJtA/RRl/ZdOvQ7/7ogv/R1HMIY
UO8nhySvfHD7KulN8Pwctk+MBw/TrnKgQ2t6Bm9c2l8QoZoR62RgeheMRIuwgIBNZuOaFuk5m9Mi
DrSORcNmdi6R5D+SeFfR5LtWSuyQs7t3/4YxNYVFZLmT+BOaykg6QjCDfiQOvx42NHr+AC/K6rXJ
uOanwKZibNsismEKzdSVyiIcsQ/m8ueIE4O7XEL1v2LkQ+mWLRwvvGIFIl27wvuTf9eO4D9Es9mU
uZd4nA2YRKQmgXs6MD+L1oLlz64HJ6ntRV4maHPvpq8c7kX+i88wj6EOtF/QM+NhWZbX7n+/tl/9
GcMfTszYrBFGWvunCJjsNczcgGi7lrM8S40iy3CcYHprVSC1I3yweFDly2fWpwyGKluF97B7XMI+
6wcAhbhuh/zy0MfQl5CI6E0RG5bL1X76mdKNXD9fBjmj845Yntejcoi0swU/mPxeLPZos5O/aPQc
1yeX1qWnsmY0Cpu1YQnPOEbyP9t4Kz4gWpgBC2bemltNUsa400g/OYXhSHSZjOgDbI4CJtS91N5l
GimCsO/OlvGT4g43Sg0j1u/kJDGPv7F47hVP9+WlakBFynCFHQOzxvPOWzW895b0bs47gJUNXE6e
ufdbKgnmel1O+86WGKl+h6ikVhejqGU76/o9JFROv5z8kFpa+gWp5e0rOwaTJrL6Nt/EM8XPr0GD
eWnMB0ea9t1OzbL5NCkTi6VnMdqahvSEIlyZFjydeKsYEtnzXtFgD9dmfPxMUuIt6ekmQanyYYRG
yMouhCMBg9JUv5/3rjge8ehXhGF2UZkwOGmn2noDA4pCPltlFuNUOR2zMFQ0xfR/ePQykxNBsx86
1DTlK03dOz369rUzhU3ZuHSslD1KFnDT0QQ/gZUgGzJAIJsEgGeqTWMSvD0HbQFtMIovmF3Iixvr
/q7B/82k5JtVtziwc0TgzwBYcfDykn4exf/kTN2HKF4LfKSVtBhRAqu8sP19x15kpxH7MYvQYiZv
V8FMOcltIaHUnRI4Z4uneFMoNk9h3Q6LWP9768Dte0CylNFymwRxAXcQ9SJiS9YKp1Q/4mjthmEW
ohYp75MUtaQt7VM/LUXYqh3ACrvgoWqiDaWSQLKzwYuqv7z7vaRbhnqFoG5IMkSq/scBqpzW+5io
nyxtrHoUWKZYyDVH5j9nXl7c61gvnKebGZTtLIv3d6vDDxez4O0/h3CbsPu0Cfx5rnU+3FH0a229
6dGG9P5rEkjciqOb0SAetpAolBDtYO/di+9w2zvQEAJ/lG6RLSWYn1gOqD0dleOS6fRayvBes6Pr
X38tyIG3hAH6g/wBsAqglJklY7Zx55ZdmwdU9NsFJbt29onGwccq/W84X96xEA5xFXnki5moAAE5
iylq9tqOJDo9/bspTp5sW2M+kBtKzUt2tTlvXhL9yQW8vkoLSUG2d9FBRho1m+72yRtWTFsObJXD
6Dm8qhmRatWVjpX31iuH/5zFsHhGT3AIDmkvAMyFABJdag2Z5m7q9xzMt2atVDsEd6COwCm5IRJu
do4nfbe07SoUJbJFIIPQCbvYAJqPCEiijoSaVyTRYOUBEVHDM/qbrGv7EU0PKcXgF6OUe+5Gthjv
gxYjWHmUxiFiLQgFZtG+qLP34vcxtfWhYmE4c1AbIndRQQCbdGUrrPZI6YK7yJB4Dp+Ytvvfzd1m
udnN8dlqCeCTM9SubyCVoiEPRKRc3w2/OwEh9IRulwGvExkZyfa6Yy5h8wxNIuWH3mXo0ho27WSx
AUas3BI2hoHCS/dMzPZs5iDXQ4TpLyEmUUj2e2VZ0PU06xsoMKH02HErYLJaIWT6s1FZdMaDhSO8
4b9Faw/tUQ9osG0Yo/EeNgt7Q1MszOsjamqO3+FO1HoD7BK58GlDjhVqgZQZL6geFaSVS6QsUk5l
On59wVmwlCe1kBSZ/yQOyMdEmA5x8VewMPDmcyZmWw1S+oYQeEE/LCrEz5und8eZCfrSTxzEDmoL
V3JIjkpqGtJfWmiONFA7ApO/J1HwPcyzjMOUd97g23uVTazDYlbSJV+VFxJtYKazab2W8V8nOMjr
Bjw36tHJGdNh8Jm2BqX+ATeQdkpl3S+ngrnsHXX/HAJvaoezsw+hA6Sn/xIh6T9FxzLy/bGvSoyY
OrrdxT8Qwkay7TGsN3JxracqANXrp3y9EU61nCHULx8in85KxSRH5kBLC2YzhmgQP/ITQQx6EVFn
2HSUnrIWoLznYBHZdMAvZPc8vfV+6ScNHuvqpstSA1aus+8JCqZgcty0E/1mSd4oaJMfiYLzUvu4
JxHZ+IydMhXguBqPzW4YK+uGaxocWAz+DQK0U+Q4+ZzYaCpvXy0XXFPwkmpsQ224AryiMs41bmf7
mhRzWNUdGVJ3DlbB29omy7R4e80ZdW1dPHx2V25Cgwg46dBLHXaBLRuHH5rkplE4rENy0pJBh3HF
/ADRPwXjQjrQdSThAp5xzWLoHki7w5IN8/mxT3wWAjOGltKR7edZi0sDsAEaVPR46yNMsSdsS46h
ukJ3Qv1uDWLRpM1dMPTPnXTGP+G6Tj7j51eaAIPILH84836cIL63RhwnWG6MPN4PZ8AcXp/cyS16
uQvkizqZCAvQt5TAFmWFx04QPr+EnmqmmL9ujVSSI1VNisrzuBROIne4QQKaKsTilIWmol/Zu9l/
WEE+KO3rDvFfy9y2vWB4JMI/oLsAPunJyHRld2ZFxqEnOTFhDbHl0YPhevjBvA1g8J84M3ZF4AGl
my+2N3OZCkUryRti6PEbmbt694YW65q5vnX9z8R+p9FO5jJiCH1nNCNmglP6TUvrP+CNK7oLNUxj
kERobP/7i//RpWyq2mw3e+bxipzKlXprHxprimsOfNMWy1G6mMVueE8z1ZGogZrVszsbCUYofP83
ToRyp7e49PWbjKzm6cVS4AZCAegMkbWzeWNvqwYhDpcVvU7Xo06NoppOMfO5kNasib/fPH0EKfyO
0tIODDHY/rc+mYjAn/NbmdGP5mBemheqpBJ++JTtXw73EPSFKT0UcS/NNOF+PabCB48bcY3xVkWb
eQbum5hF8XRchDYRhrW7HO5zVP1MszmkPZGg33FZ21zJuSG9kACcDilmZlMzW/S8q1OYsykHhkgD
UNXhNdwnJc57sQHIYnCPyr+f5Dp+xlPtVxUckjPD4HleJtoHVC4gnksJBD/8u7P4F2CGFE0ICk3y
sbhouC9ZtKQ7eazmRRi1P+38dZmKeNdwMxOYaUsjUWTbOKdAak8Eaz5rt9HDYXo3I2rZlmC43lWn
xJzDxm62VUdmwoVc2mu9AJScSwGw6Gd1c4FxVKr1X48BZZXrrWItqoS5SZEsGprk/VpAQCpA8j83
K3RI8iS+sDxXx49/CaVlLnRhfy+YLZmyCfl2DTXJRTfMPSHcUOTWp9wVvS35Gv3sxIhtQ1covd/u
4/Ud9yFlBddCW6qKYJgXVHUhsQK1nQFg6xZYGMlyyKcrOKL5ZEYfJskiqRBGu2arPXLXUycvfQhA
pDEeYiKilQzqIhp7aXozCABwYmI9gnAPkwPBZb+tSR2eWYWYquVUZbeY6SIXYAunw/B+hciCz0G2
pDNVlDbp6Al+nI+hoOzr8Sp2USNrk/pfcvVWc09Rqm1SyLtSDaowRtNhrZUQc5xHdwSX56UYVFkE
ng5IfMMQQFobM8P7dx0W1MEe6CETEX0ryZU2wXRMJ7nvO8mr1PPJJ2iCl93W6RHnzhK9ciLC098D
YOP2h58TDFE48gkierIx/qP83Wu4oy4DkJaZnoJRFC+sBy7x8aW4J4yF+2HgYS4tJZ0uPiwaF+e3
uK3vNS9ZFBnUSfk8fUwklJ0/kls0uOeICDzd6v5QFNzqrwr4T8QThyiVG7TRO7l386WU+VwjZ73o
Hfzg7p+NCxksljVaZloMiOIKTZdFu+gzvm0623IwuuQTGDPzH+jGMtSN/qDYyuffcjoANK8lvLBp
pDtcLlVEBBc8SQR5wN3xqp/9bVtS+Dq+wt4uXBEgBLiTMXHLdLXz8168w9OVL1ch9NWZQaV6o1pO
UC5vs3Mn2yCRPTXQClhotYH51EajSqeJe1ariiTO8yD1pRIXsZ1cFftOgyhU5NIB0kBOrVnb5h4A
9Mzp/SkV7rXRjKmySgJJi3EiorBwHMKfC3z+ZP8aOoFE2MTyQ1E3kiJ4jtVk2U7r/DH69ucxj1lk
jWRhgjRXr932RiHdyZsgp1pg+/nJH4awdKN1khtMVcrgppvg+3DweFVhK77yZ3xE3j734lUqDDL/
hrVhaG1tkJn+dxM7HypuqNIE2qCqKk36Hv3i/e2VBUAqmz9y3wywVgSn0R21hjesHMZZpPxqQARZ
21EDvmxVo5uu4wMGDt05kQRlLl/2WT8l1YJZJOZ2uWot5pyFSGvOsB8EfGbUnR7OApO85WSi5F3v
gnS2JiEp7KBtkUZOecD1kpcgxasaiq1zl5HuS8hOhOFBSstzR8bJO6+sueEOCvVTrB8olZEFubAu
vMhJMbyRw53Bwc0/XEG1EDDm7fBYh9GazJwMCDGmbTFozFfnKRLiKLjMxfU+zQYd2Y39Ci2egvEF
7OqeXV39UDDuI/BZ9ft+9eDbxfubvT57mCwLco0siCp0M5AS1UgRSTqZ384P5QlQRZdiKBttPeEM
wYW/4klwD3R610dGPMbjjD0eFZKM/4Sy+LjlCw6qLhVjX54dmOjdsYIdRd1PxMSo4POnI1L+nnD8
l4Txqie9Xz/TMoQwCOBegB3hxSwPCZQMTiZ4Fv7Pfh6lz3nC5G8qbnd0ZM9PYLcVv9rcBvOYRgAj
R6cHUMG3TWhD4fa76JV7Lo0z5dI49B4v8HNBxmyjRfwpS+TU/WTOhwyvH2DpxlGlZS6zNi21LS9j
el23Ni1EvbPlI4T9N/NfxC9Sh66VftHV5C+Pep00VPNinDDnf82o7eDi1JndfAhoNN+q5WH6A2jI
nJ12Iyl9Hli1p01WkStq6rlopi/re35ZvON0t3mTy7RcacgUyT9N3U2WRtzp51q/smh/HM6t1ywd
dDphlT69k/gZcDLGy3pV5AQvsDjD/cuMDiy2CFmVfXHPScPvQp31CCaxo0FljhpIZwdsZlFGxqLt
M7isZIL6pNIUWWJpkAYXuEQvVnUs0Aicw8S2d8ZFNdVf2B0bGiciSTyMqfRFi7XKsR2viCAd+2RU
8BfHbpd2DsuLmJM4Lv15jkWQGQNTMBXm90n1yu+cxhrOaEiNdTeP53CFcjCdAssVtJCW7mAfB8gW
RlQ1PoxT9Th5E7zrM/k2LzVX7Xswjskki3I4QGXjpCbN2AKGvX9umzEN4a4jfc81mUKISZKc5Nse
M/kOyCZ2qAzqBBGXz7ICIkFZlpBc9hVbbKqhLaflNGM4NuzGlZGpl4EHuR/9+sbFKyZoPdBRFpPp
/W1BrgiYukKcGteWoG8bvUvbYveb4Jb7t5qRrbkjgwklsdMEPQJBapCnBl50azDipalfDEWCg0+d
zq8gG9B4I2FWY2qAEPzKi7G7wAcj2SC8JDobRKy90wFLG/wcFgDu+nJ9n/AVGVYnFjFLquEDGBoA
/AGi+7TEh6dxzNIP1zAmpfmffQBDKsbzhV6WjFJju98bHWZbUaEfEup2dqell3h0G4uXPe3B1i+0
AawnE75b00j6JcvEGG17Fry3gpCV9CKpMeSnqChjtu7JtB/wHJVRi5Y3BNbP/RekiXyqdxQzioOz
fvp//NyOW84Feuv+GO5v9KHHdWPgdmH69qu+E1oU7BBgw/JSJNrv9qJHn/emIKoBeA/tu2vl6OBx
Qk2N4Px/s0HEaV/T8eZzChS1RnxIAdrH70C8+bE+C6dFaK7QlFNJuCLXpGkh4IXMj9g+Z8Q40y/V
+O+ihdhe1h36lvaky6kcvqJbBiirdyx0gXMRM8+EzjnGFKNjBiy8rHlAkEMMNeDUqFmxWiJBf3yw
65ow4QDV7hi1+lehKMabAPNTg0KmQsSw4p6VzKGJetefxrvUiX6dXEo6GcNy+bney3hhhl0JfyHn
AQwWakz6j/LnV/MEob43LG4ti5kbowIneCUgamjP+nK36deIkNOXwLiHTCrWecg1nK6aW30v3w3x
QNPj8GozvyVFnW30dXcUm83WrxK3GBGsag/b2mHhEow9HP5ku1nyssaflUQeKQS5B2gwUAvtODpl
sfw0P9rZs7mIj6rxTcPDpoXvHr42G/7V6gwN1zy7l9YMFWb5asNL2G08WW09X7DLdhNf129tJAuf
S5qZkbzrfu4rXgw+4v7JaiZURBEnx8IDV495txe6/90m0kxe4Z10d357LSPix2cmgF1rMiuyig4q
8jAa6OL/C8ZAWPSFuiizDMEoOzTZe+FEHXhvVoBA/DuR4ol6WtCIt3dC+SHOg1Z6qGhW1AiVj070
JdM4G8SzpCOrM+ZPoE5TW81yLSyqmVEHaeeB0+ny1KctQUvsmolVahzpj/k55nk3TZ61ompaEPxi
m3I3xk780WxiQjy6VaPgt/3q4UpED14n6d/5VcAPTR9UtESKaSlSdz03yLwJWqb2re2lPVDgbAo0
f2pNSBTliVVku8uQ69BKfxGY4kq3twXsBJxBo7hFhdJAmPQWJ9gVWHmTYDcCImhkPCK+4iQcShVW
2UbW+zC3g6sEqYNjJ3lLVisyGyFGNJw6gdGgPwJC889BpugjtvulhqrV8jFsDLfZ83qWPvCdgcg/
HFKBHg0+I4JC65+RIVyes+oVn7NxSgv3HGfO1naZOPQRT2YEXUARb+cCIvDveupCxzyZD+zA4YmW
7IbRswM5cl+kamXbPE/0Am+bedhOoBD4Zkh33DW5vPmMXBRue9f//e729BYpYjzT+6gasYDzlcjm
BH8ggLILk7tYlsn6ZWhrX7RlZ8cw2iMp4HD2Rs+0++yJIRayNy/krUZyDGm1EkE6r0t4UuMfKS1u
ssYkv/l6rlh3unSI2FVtlAL6aGNptM6SO7p/smy3Vff6Zp4dMiXpJSwuJalef45BLDsoPUICL0G6
GetqoCoWuzH4gEln3cwSXA/NNQRd69qwaXfGW2sJZwt61gbTe4cg1mdbgb1D4TyC2B0NgqMfJCT3
DnnO+Mv4RsehqGyCryhqBaOcTU6E7q+1TyMHUQXhatHc7KCrI7PBrgQg5shu9k1EOcPs0I5LCngf
AzeqxRdp/Dv5vf9Z6/djaaVaW+SvnvChZ/t5Yw47e69BA8ulbQjdJ+sk9YC3hq1kL/sTjLYeMPgF
KL2YBjQrh+0kmJ1N0nHNotczFaMzJ4eE1B3j8txZ83zch8mZgYbPt/qDUE1pAOGhgobX0uUNLRh/
L614u0nbec63a9IhrbepnIboHNPEf0637+anMq2rrBD5kO9OwyuDDmwrjdtjnp+bpn0hPM75thbU
uGe0ZY32pv0uhCiXZYO8Unrb6e718j/yPe9CHGrA92pb7NUuy5uGAYGP6NhA+xNKngLwP9TtLxyC
8d4X8Mbgq36Qke5fMVPm+Mj75CXY2iIIL0l/6YmvGwWQEpwiS947JVfFyQmW/Ffyq4ll5E0HQu85
gNUoQkOiPAaU4t5GtP1HoDxyOXm2lk1SldI5Na17lRBULzrAm0L55KjexV+B2quzs2VoZpVOCA9C
FARd0DGMvoiKqOFv/0HMEIiY4Q3a0qBgkDHoo55/P7dTu8ZIFshzpO9DisPh0tGFtkinlUxMYUg8
cKyqTmp5mxWXE0V7TPw00rrZ0Xws8D1946XUoSmr72bsVnKMOioqRv3NV+a22n48mqJx+DQqju7n
D2zzrQOuKyBwzR3Uwn11gxHeHL+JBbqGq7PihezgYQnoqpKrGZ2CrH0RNQG0IaOqJ74RyfJtpkf1
SBLE/iNgFHHHBjn0rekEQXQgvCZz8lIN6pP/wgiWcp7Ymy5lcrQUCE4c+LB58ZA+G2rME5iNIv95
r/OBDZG2rYUPNiA14uepVludyUUkPmt6zc8uGi8v46lsHgkDioscz2JqSOqu6Q/w4eU91YwlZnQV
JAjh2VklW4eTkpoRYULB2SAcpzDFxDRGXlGJSPDQsccGJzjGqweq60HrnUPY2usqkp6cmUIDYiec
pm3tM38KDDNNa0SkQB+0pNn1fAh2iyZEuTbalVfreJelevnAbEmcRRYgbPFZ91ZhhGUpdTJKgyLB
Wy1mxd16uHehk3urZdIMSrmIE9u3V0TMaf1RhnEvYlmA+1Um1Lq/e4xJpPeb9xfXBAaXWh/MycQR
YW1iMSV1fCAjYxD525chtds20xTsUV/nyN7gQ9RWBjErhviTdR11zmgxcZ/CQybl2xjwaA/eIvXm
yJtQDQ0prfq6/siwmEt6lU3gb9vMxJmV4S3hdNXRvQopzqBkePAvxaaQlPkCimecMB5nZFYxtvqU
dZ2hg53amle9msEWwFfhF67NihpzYxed4gdmMWGyOR93MJjlnbzihsWoyAd2s5tzGIdmOgjQFfj0
fg5htq0ZgEsakTVmktNdDqeTRm4A2qAZX9VwA0ny0EG53LlYmmQZUPS0/QL9jeyvzRFY8OYLDjbe
USJ95uYsjzhYsuREnjNjxQ4s5rCO/OOCgtT8VMf9qbDjh1RJEgdZ2n/l2tXPdSFSlesB+1U38RV8
EW85/zmDJDs4Gp1zummN5pqEyWIA2sgp24x6GMEHVivd0/EZ2exieai0ORUUflfzwp4ha3ooa71G
FJKRXtCot5CpWoDDJD8hYH7fKcgj+bMHMtuEqftspIbkn5iHduDut7aIQr/yXnq0r1WwQ9djRjny
Df0/Ccun3WxrPgtsgFJU9I1v5zRDJJAHzVj7Kh+aKu2yG8pbaqyMbOP0l4i87yYMsVC8S4EHbW7v
nVTU0zN43N1otJBJIFhWYttdWCy5qE9mYR94FU3KeZifIGmErfJypr10yVe5jvsQce7o8+cSzSX0
qACs/kuN6xxklYzD+9KUQcNdBEGtBVm44v0knSHaK8F+9MMLlv9Ya5rYm9qDbZ7fjtA5UTIfKrRq
55ecX8xlkSmI1sOeOzv9TtVeHpuMAX+pExHKPFsXH+apJIy6ta/lxi/fhGYRtJyl2bv1JNZLUyjf
8bi4MRoAqy4fHSKDlf+Y6MBiTyzxcX+Ft+nPCrgMJjcD5OyAcpiF1I/G+WS0Rv73yFFEhWFx0gC1
z59qxf4u5971fr3yXURMZ8qdln6dDN7Ro8QbSS8K2/TbOuY5rcLXFddec0Kfigz7sFTRzViUSwRC
z/nX1A/bpCfabVb1Is27C1Kn70gJITeR4KpfzqXC1wQS2VD2qEjQz67VwrF3rtNBgoP1ehlnkPiC
xp84GsyaEO4VuV9Wc/cU3b/d4ezicyXVf19xbLnjwJreadnNX9FA1QJ1KpOvFM/1/2ZLyEQEgQ1p
MgedB7vX/Y8+kWfGsCdvSCgAf9hg/MhYN3jBEw2NNd57JCIDLNjderNBDMijn7u3nYotkUrWaoBw
XVddL/XR8w/eBZbg+MrvTUXDXHksF6Mik1UE4KIlhtlKbOoBxSU5aXiGgP+amNugTsZRc96OzVjV
aVlCjs4WVzW4D29QAHx92MT6ha5YD1Hzn3wWJbrgd+zCHB0f5tOSOP6OBMZ5BO1wz8wTZarnwAbn
ayRHj5BHCMkW+Pfjd36iMbFmVsJ5Fc1O3kOu9MVSLbXp9s9UKY+RHNiLAwNT3fZNMxBwR21PgFOY
5G/PIYtRDyJhq+m7MzLlKZt4CmbKy6fGyAURwNnErDTiYX6GRWMaxIUotazstP2wdBdbAaQjddW8
gT8k0NZ03QNczGBd6WXHbHX/xCqkI1MgQJATEn8HAG7cU6RUq2lTO8b+YVXC8JcTUBIRuV4GL8aI
O5vW2NaPDdMO4+eqigI6MrhdD7hn/qp4ltbDhZXCP4Q5KybvHyZZGzkAkQHaFQLA6Nbv7rigMheh
KdT8EpaFGWdjSQesqxNbFFpY72Gd0FO82LSz4CtphWvSiO6lvlXBYM8UQ3SpR6qW9vwSAVArjkZv
2bwBVJ9anIGv4fzES/tw2vY3w4Ba9cUU+I4dcsxT/9N/odG8aAPno2zTo6N52xuO6Toz4C5u/81G
7D+HCD/1hT449fjVaVTmYxh+PscfwC/pff54CrYwETqzU1px+kmbUpyKZKuZ0ajl57teNfgGuZ1U
qbFjuz4pdVgLwdsnZE9WpCrAV7SlSu7u7rZpABt/DDy9n38CtR0jDrT3L24oSjoSCNe2zMWZ/gp7
Uw1fkTV9NwxzUX+lBHTiW5lpTdlCogirlMqpP8Ij7z0WjSzxOqBP5xim6nrAytRWnHVDSWoXigQa
cx/OehVa/lyDqGlUt7/3UGhxEqw2hW1KRgzbl5fqFy8PoZ5RsxKaro9N7OQ4/g/tsWKNG5lxuYbJ
uzT3AF2jwiPdWFsOzeVIu38bS+mRuMRDyqfvBjBEr/k+Ic++DepPYC8oLUksbQ33vIg+57750idU
qddkAc8Gbt5a200zlgvaxB58ibllfv1adFAFWmZUF6nrMFUaZDg/cpPOo3HBhDOViYmUWc9pU5Oy
edDdctOhJ8LDa+x/TcngkkrRJQZLWpE7nC/gH8drG7hdYQ6rnyjhWR7xRfyt/ykcePuEoCX1/xts
SW6lGUN8cZjDiJR9Pa41IlK0vpHrgiKH8Q9MZlpkUlX+crYCtZEpStKGaYZfHM4iRbBHtn2ZzfEd
K/PFhUTjF1w5pnuQT1xpOSEnkvDqwEnEfO6jdpMIGpO2myo2rNtHX8PzOR5jHQ6V5v/moaHMp/mT
nCvNO8b3/T/fvOYglARvxgawitqUo52BlASWbFSL8lPAOdwyTkcL9DHZYeWXiJQQ4HzZBfEdumvq
IF66+43tSnKftSyuilT4GQGT7sfagJJ80twc7K5w8D7czigNWumae8Kxa7S9DUX5I0qiAi60Ny19
62uD8GnB5X6RsEM6b8pXTQOAgh+fwJvhqVR4TZuRQEvhO8zC75gx7LXh630auyAqOUeI6UXgzlev
CNtdZ7+j48fP1vl4ULytSaOD6EpFySOTJVEGcTPo+8xVxVGbLBCTzL7y3DQSzc/aTvu8NhwjFfMt
eKK2nFZO0Bbz3UGlW/AFIMbADXQSMUHVJrpdOoRu5v1N2ck1z+HgE/oWECU20k4xtXZyZ9Y2vNE9
Hqu/H+Dwc/DILxKMemVzumiwW3DCD2jaRJy83V8MKwc/AKD2KPgUyiXrvb12VhEQEz7/n/VCMz9Y
IUdZecnyHS0GDhd1hkVAAdgXoPCrDRExUfaTd2VlSM3rXqv926SwaySe418s+nFRCqW5qwLr+X7N
085tKyYqRB2wJow0fKyWy1Y/02HN+KAR7d8tksI5H46mopUTxmfXvCVFWt49PEqtUtJraHThBVQo
FskYEmwl67hbIM9lc/0G24H4kDfAycDQfMNbkW1BlkMsSPaVBW9JqrYLW1xN9WxOX/dqFJcnF73+
vz0+iABWSEkQZfgGiv70VI14H/48q838BOT2yUPuisfeMR+POiUlzZNXl+daBuYIyxogdXKN3f0K
LKSX3tJDdimgivjLhIjqahdnFUPDtN2Xou+lHa8B85lEMhQwo1L6McdEBRpkvsJV8rATqWao1FCf
ArDXLn4zLC9nZ1YcPxEwlsa9ud2BBcmoGg8Abqw/itW2b5kQGrawnUr8TbxNRsmIZI4kozvD1D1s
N6IOnusFZVQf3tBQeiEOtNYUxoLmSI7m1IbfmqKL1I+xkyFK9fIJZKl926T6HHp2rcg1Rrk3h+Uq
3QJW60tvUoh+n6aZ2XiXRsKD9Fltr8Jpwy2E/8VG9wYaG9l9i1gj4JUja3Z2nV9lqSPLZ65m9aPs
l629MHJCTefhh3ZvxSIG2V4h93XnKiPnutxCa7q3BsnrSBN4d1R4yCVHNKtl6g8uHkDIBtEt3y/g
wdrVW+80pgtqEOIGEobvMhEP1HVAAXP6OiwKAEXBS+K374TbRxtOh929nq2Qg1oTeaJgTPowfPeS
T/AoUwSW4rphVjRzmZIqMZneJkOo1oxthH8G1hD2ZalDaDkRW8UO2nietq0w286qEkcGLqkDrruy
S11atzvgvjDSHU5jdIjw9rHqlfZeKupmCOqOXqZUa9mTi8QHHi6lz/HatxVWlJ/JHnxzUyCZbIyi
dpJrPHTlUPPGR8bvqEF6yVHqec2Hc/aMaGrABAMmmiTvdwfhttgsp0jpDB3TYxiSGH14MwP0em1B
6PfNXhelTFlSXI/kp97XI8sInpIf1CAgDYvsITXYLGHiPWbsp+GDXFC/104RGlt6AuU6KubSBdw4
Q4OrRB97n6KVxxp1JZ/YnUrBHar3KBMn5hwJLt2PdtJasF+kRNhcg+OcB4Ae44r56PAtb26Ftjku
BpksVtJ77PuAKGdrgpidU96v69UhFbY+noAbylirhdaBpGra5Hy6/46096KjgXOlpX/gfQAsB4U9
rl5jT96+1F+ORXWkG+rQUc0/AaYgTRWWQRzxPRiKdCr9azXEBWAWEkcvRps4MXdlfT6ofZ7GbqiI
zSQF5Wz1KbrekFphPH8a+/0Tn1z30wzlegDfn0LPtTzOuzfekoi1xDspd74de8cwzD/W2E9A9ZAV
405hmyCP5VFDGUsavMiBkhXpfIX57zv/5wZRKA4PEkGYo8zW3q7PaRpVjTtMa1xuVO0acNhQLT8I
tIzgr8gEBkpBwdHL+GMBTTuax5ZN3pQe7SYQ2nwMUyTKG2ZyS9jnDZbxGyYmCYf0wGr/zNhZ3hMS
93SEIcWNt0oyWndzgA8CozMVt/zty3zq71YB5g1CLvWdWK8/OUQ2Y+Vp3wmxg8/M9Pp3cSLp5bcO
XU7y/Nzxk6FSRmNoyNOxvb3ffWqnhXMaMB974O9J9Tu9pYMwmQyyoPhfID7jYjS59leld0XJMgul
I84f6QrItf4o2xa+txcbMZwlWCJQDFU70wzMjVrdsKpoM0xzYB1XgMwZP85wPbOFsKqeICE8NuZi
DF8UNfl4t1n5iioIJz53qP8wrBsb9rSFzd4yMz0dDDcmIK3tdTxMxq9HHJ4i1j6fvEk9C7K4NzD0
0rjCVr7oZwBKgI391ZO56Z+cSsTc+leMZv5teiNmpMyJdIsNnBhks/CzYcK746xzffgUap9rqK/b
8Y+v44/STdE5GkduyjEQaFbTBVgWq763a3B4LLu+KdW1HHQN/xTkacwGUfync4nelJWmPj655EeD
hmzdeFIiZlbOph4+MxgvIh+xJ8n5QZvyfgCBZhCaKVqXZwSxU/gHyQre3nvCqcdRkiykyLz7nktF
8Xpho8EjBnLgDywE/Rjn+VrfZBFtwm6Q+6i2vxksQa+3URuk/gsuarx/ax3toQIv6xxWXWjod6IY
FJ82R/kG9VtUnpS9TpKasE3eW3AFz8OV5e9EVC2UFBQuZR6WXQTl+n2bhDHfpSHd3jm9LbZHRlPg
fVo83t5EHuTe9xfP/TiTwHZ+YoUiSpmWk8oRabqxFIhy/J3qGFn6J58jiiKX16xOtKVRXls4PiUJ
Oqg3jlRdM/0I2oADYJtVa63QqC5MmxseD5TDYPPOowMYVAoydxcMmKiThPJvf5FLU2H4Tv5qbgkw
nk/rqJO/w402ZMRbQv6XMIlrdEeDUYKaa2uCnV44tCIU1B457CJTrWzTPaN16oW//zN4xw2JEIlB
DR9a8zCkGAlGelnMK2jnHivtsWp7UqDFTlU5y/3gq9dMh2gOEmoveat2VQnYKZnKHfS1luyiy6oC
Nme8uUgJQdT34E71+R9VQ4iDthHpOE2KBfGpbSNJPP2c5j4Lvm1MzRHDBXaApMkVc4I3DOox6rqJ
LNkY+7j1CsV4OrXXJaBVBf4VkSTPFm/99J5zM9N5xNnNkdQbKaRzjRp+Vg9ZpiCM53HjInARyIbf
hyc6/Kc4vidBtLOR7XcVQSme6xjPCghgA2MD9lfIYad3c2+WaRVuYKDWF9f0R0mfgMuxP2za4qRi
Doo+mpwoH3q0/AoGbzU2nNRYBQZ10yt0kspO6utR0yK9HKxplbxmmQIqcpLJrrcgZXBQw7zotJVo
1344IJrA5Ix+PXg2kvEryOz1J0YZUovpxJU5BVhQaC/9xFzCoa1O8DvzDDHoBpljNMXWwlAm5PyA
gPL4CYALdDvBKhSjZ6Lw7TJglneb8eVNPUjNP4LIHNzsr+xaME1fp1/oUA2EjApox2yN6Hf9tkjS
xhyweqZCofrERikOTnOa6Nwg9rmdLYMVymsWTh36ikxor+OdWPeyaP2txA/mbTb46hBW/kIqF8Dk
NZ4LUL5k9tkNzIjDsyIJt0xPE9jVP9r6Rs9ZA2eI9ndDW4FgjgyeHsMfIkFrMgNYRqPCXeF5OAw1
w1xdtjRozerQfySS9qZS6ER+le4ES8L5WZYw8VRVwBQSX9mXUYjYSdX4tID6sj9aulSpFhzDj/wA
0YeT62BMvljdkaFxbgcs3CPrUv0ZbdQ7gbNyVVSJOgbS9XW7dt2V8anyVfwfEAJjogPBlHxFN7tv
tmQ7khf1I01fXcZY7+CNlj4HvCGpRXEMSdU5mhfi+FUHvh1DTbU7h0FXEHRecKGG8rHIcbrYA32c
3i5tNuWAp+oN9WCPNYDWFHBKuJ+OdKraz/xwSBgqdquAys9Di5+dtpLv22TVEyxDXI5/KfRmy2nn
7SEFR1mmvpSEpuigB17Mr6voBMLPWCJyqedgolsqkSATXWEaIL6+2CT0bK1O10cGvoN2VStavKwS
Ridec+HnTPjPBQ/BdYIxy6WK66qiQwE+J13S8qAZmQTKC4WGMyNZOqInTeJLl6guiSRLCiWSnTkg
JrXypGCiK7Fvw8PLmnJl2Zr1xF8SYGLm5Ly+abxi1Ekh21QAu/34Pwy7NCXTEJf7d4G7hX7zK7hB
U132erOUvg17+iDIr+XzNwJnjAxySBIxDFSlqoclGpdr81VwHrYbd/CEcXjcsqoSXuIBXzHwYZz7
ho4cHqhF/nzRoc83oLGJmrbyP0R9B57WhE0unsyuHGIpTDmBJwCYb8Z0keeZD9cOnkCUvETw3khX
razRUZKHigMF34owC5BQjLplujl0xi23Pci8LzduZoF7bV9aX1vYnj1dT1DQhzvBzpnITKKAhIvA
8McPxXhCLO6QQ/7KhcveCC/2OjuRsmujhe+N8PmqAU6KEU7hTb/6qrD5o5GgYm6b+bew7X/Os4F9
ehM57scFRjOHhEG3jy0fvuRM2ctuw5d8q/Y//bnKLIZ+eudZph2/V/NNRwE3yGmZ89hmfpRvpK/W
a5bmaHrEUm7Hr4zf7vZDl7UWNxwiAYFQ6//MswprpEOWXxvsNjdRhcfqjmRzvd4aCE3i4aygpBxA
pvjYUjnQa3Hzw0x539wXJviTB1vpECVPwH1rtEuGlVi/ByOo4HLR96WT077UtBJYqKBF3nTNYTww
r73N3E57uFTzbwWD4QJ9obPvTWqHXWTS7kSkcCzNpbDYMbtVBoDfwFDA8k3X3f1Evy/jB4ruEjYO
Ty9w5jBfVLMgN0CQK9B7PkYg/ZNeJgTgmkMktBzimZioUrX0qqLRrdBxb2X80fsE2+HCrWVJxEcG
bOngVLKaPpCKRBVsuxQNKqbVOKXLqSbUhagCBduRlFKME8jbrK74kyfnTIAwlF8Sen7uWLNGCNNo
9qQq8FuF7NjnXWnN6LXZHY50e41xjcvurE8sOHkXUk1rLQi1LqE43BhHL/wYyj9J8N4tSp/ohNTf
h7fHvXPlJYYWzzgEk1cvX1INj5Pd9732h6h28RBTBzJcNJwrwzYhXkWPd6Lny+yX8TUPk65UzxA8
5MR8BOesW/bAaK4OuyDnuZKHOhbBzGTdJd+TKNyXVqAZ8iTZ0FA7HChceAxI7R3UJIHtodkzaeYq
CLvvC/21X/sZg+6WYdeLugZyJqDS7EsGxX2+RYcp1pN4Rn2AmHjTggJ6FrCSH7ra1hEW8/AI8SM+
gKzH9U2RfMzNri/MFG1gzh55CxHede5/Xj0gclWNcINo22jg5Kur/QXSPi4qJGt/npcJ1MUE5B00
psAHSfowsq3Nm82tnOhas1fAaG+IX+RZ5YO8WsrWRTmjuVHEXFSauunChrD7gS4Ij7ukyWC77TFw
sx969r0IbgKQ3zITkSWusg1ufFVFK6s7Xkh6Edq/mc/N/Si7Jxu32JdhcwfV5c6XPo5gdxfnuuwf
q38cHNJHWhg+E6c4S24DB36xZiDz7OjZHqv5qXAtTXAzjGMcZEiLrHwNvIp6LfQEeNm4qroKiWmo
cCsVmyCY78dC2QMkbjfCm7XioOZnqXCh6NmBFRe1acLoXfCy3VvC902W6VmZwXf+dATtVUVAPLl9
lFv2dIlS6sVMRnYTDuOKD396q+9dZQawr6vcnq8fJfSaYp4eTqSLUP7x99iLqCOTEOyDz3FCoLwq
2+biq3Z3NIK6geFGrebeDHhoLV4Mw71JIoki29PrNsO2BKBbPdJSaw6VtEcH7xNjRrFmkN6vm052
qLI8epUNHkzIhy9lEM0wsxJXmkA7CEXRyfhQTlmJHrDNMUIi/oajXjW9h4+8H0EjsP1llqoMukXr
brVBeFOY+XI7jIyNGy7d0nzhtmriJP8H2lbnm5o3toul72fzRpoYMlC4Y89hTolC9MV9/VRJ5XRL
dmxcq255wef0rycZEQh5Z3CEqtrZ5z7tx5ch3bYvaGFRcsVE5s464r4WLSc5oG+HWat0NPCD7LoK
dLN/lqtCt8u0SLnbv1Nox2eIX/hQDL4dGQYjofxvpQ8EeeFXqVareE6T3ASmGiCIXngxsSFuIYtH
2qLKbRo5uDhVXiwGaql33dDfEf7OPeAanQRqUf02+rAsTVQYiYsWqj2WvMzQSZCPi1pPmqsZUVCc
uqDKuRu5e9GFCzNNQReQKR8llj0v+311SPHaNymEsqF0OtD4l6pXUgofwEOwdTchg8cgUKRoNYlj
SUkSpvz0VwMwkEef539KY52V5GzyQ9A9WCVU0+aEo74D+FBoevfhoJ3FxmwVZ1nbS8bvR7pcOKe1
YneAhOOMGBpNTzDcnnynAroGuh3xs4/7+w6V79gGabMzAE+bfvrzp/ttnj/7vmo4EqdFZG/ZBxA1
aduy2VxwIag11MplRR32HWrpM1pXiV2cwDCb+3t3gLuEX2fNF3KrOikbAY1zakxosqCPRmR33ARu
vJWV/IFhXiqmdvqLow2E+WuketdYav9QjU02++Gag7/4EPjIm1wKyAnFy9nQ9lNsnjo5GobYlCXH
6Yv1fomM5BnlcoPxfgRZyYhWjiPdp9+1zMeOkJJYuchrYL3ajoLsdCO6bP+ur7f4lJx5lfz0/VOy
HQoCugYUf4dYP+vE4P1iGXa4IS0UTelwHOd6tqtm6vMfz36pI5LrgmB67pj8Q/dytzlYszGK+5bG
68L2KSHHOBzOaxO1Ll1XcUoWxEyn/b8sYrTx7kg03GyVye/IXmGvCYE5f9H6WLEt62/EqF81Dlff
ghdPQhkCQwYOkLrgmjVY9/Kg+6IOXOH2+QWIwUcwzLiAhNKcu6MTlmYHGjgn3FSzlzhYTaT/Y8cW
JHYgYuA1pEjzCooiijd+wEKmYToWCeTLckLazAXXUUijDl1+HE0G+zXt+2u6dlCGlZu8hbfVpgkY
fonnG1mvZGkUZ+YjKOiAUmpunaEb+XAdWlsHKICR27IB//bQEiItjNWnWzNzlTgKmUdjwla1/tGa
fh5pN3qur/92Yeo9WVyaOuRmLDi6+Lrase9f13HztGkRrXogCxW68kVrR5Y0CxBYsG7+PaluSius
TEx7yMz8Q+JQAh5z5v5Cj5xSAhrA6wM9EhswD66Aff3LE4NpAq6EsglHjYEOXIXn2Pt0f/cMINHm
7yEf0CobnrxekCPmsahBTuuSbKB8Uafw6TtzQMKWOaiXvJs+6F3ADrtzqaGdWefKzGZMeFyCwIFx
pTxA6fmcFQ3YvPRqW+9FyfT98kygNtqoLBgnfbKjdlzHVHxpHf0Wy4Iwip5j/UuAPH2POCI5edkk
GYDeCPFqZrIvISoQNTo6/SaUPYSopAIc0dUKu8OZibHFix+n+kph4BWq4qivyWprwI34N81u7XbY
9dqqIkbYraI9q9YV5N+GIB/pm1IW34nFuIkD8BVy3N8vtKe02gFy3aSTi6JBlZUIZKz47Nc6VHbq
KgueJBhASikEknUQjm9xg2P+/3a31FMk3Sm4gJEl74NrSmrdB/lMvHR4vJ6grm7L8XxM0Ka3w1tX
bbraZ87y38HVsnfN/ruV2vNzCpsQ0jONov/YC3x4PWZX8N+wAldy+7Pu1tsYvinXsblTRB2z9g31
/A3DOJTvBDA9xb0XV6PMHNwq2x8i5eaXZjgisHlujDfUE03S3T7Ph08R2hW9KubbbKyw1l1wPM6h
6EE6a/GaafjPKn4281h7YXTL2czw48MVjt/+vcH5K1kSVI8Ei0tK7877lqkxmOBwBYiFVYhvvQyc
bdHVToJscdHRQuNGKhAWPU2dJVqg1B2daArotZxCb3kyHrBe58ei9UL0MW5oof7qv2i6wECwTTcP
wP2C2PtGQwBcTolglJase6M2/7nINVUhC7Q3eencrgdpGhMkXxBUkYiBK23wKbRl2IwrsA2JXOhB
NpcsdTtJ2HOrhmDqMaMkBgfn0yaPy7rBqlDS1U8QDaQsCP+LhdP56JLkL+WFPeKYi20bQgZe5I+e
mx8K+Bn1hEUyEQGwBTpPkCzhgFrmyDyY4iDneO7YU4xnyc3ugOOT2ycK7g0RZaXtRTM7ZN8373/Z
6LyHzgPFALNid3H4IwIYoGdMO2cq5jl7C9lZ16lgQdoXc3H+BB+iVoEPxf1UaUkHScbHdo2CBJdC
kmV2aUdmTd9KWgXoVxAMj23QgNQMrQjdlc6CaOMO9C0Q8Y1ESqs6uho38paMIWhy2vQ9THIcUXDW
gTcdBzJP3HRkGUZWhenZJ37blxsPRh5xEOlrkN9GXNxIw4+RITIX/wrBxlLJdTepcCb3qHehQsFl
UIS2mfTVD2pFGb4EJw4BuNg9HnrSptsGawHctmu8ngcna5B8DCyRJwYTbUMWbgG38FPrNKLfmi29
MxE3njS5Js+wJHalrJy0z8hjShBtje3r0jYsYRSRAd+MO19YkNI7O4yFWzJwl7M/n/g6gC+wwZYe
WwnoSXm5Ufybw9cBiLJ2wcV0WccMrWgsNMUAWPC5EfMq8c0I/WFiEHm3S//0MnR2+cVjq7y0R8Xl
lt22RudKY5In5Ix0o+ePejkzii+8SfdSj8T59jwlaW6optHDLoc5v7LXrp9SFvyEnP6l/ztdnYvw
HTw9ycPWHj5NTJAgWYshO2tFIO9E79bnZLuMytzQ47/SyT91OefoGdfxuASXX7fKBEUaelxek1n0
xonqYO/aEiR4ogCH6Bko7Fgu3MDlHrVxT4F4CUrf/I3o3q+27RvTYA6iaVqYzZw9XwNg73ghDZcz
dJ+zPuQifMHy42R1OowqRYj2mgp15zfYqolhC3BsXio4YGnrl5YKZ75Y9NzqABV6wWqUzFdx6872
kYHJbKeZcBo1TnpqIG5NgDeb1qJ5UdzmWksKDyXwlsJyZyeFzypkupmzRi1/6XEK/7mKSjjNtaAK
SspoxrrXwtS/DXCmUJQ5WY9rd+fmQgC0+FcDMaAyQNSdGTHr7q63BjSWjoY56Tcyp+JU001oXFjo
NbJPdHE3JkSqZWjCUaMYaJSQTAPmLbqkrYVsCLRO4WvysM/Y1f4YpeBMl84Nea4klHZitFSiPbrZ
W9IkKfLIwnnmMHGp2XJSJAvFKMJ7nFB5spHDspRWbYidiiyeFbMa94R+2ArRG28gnEi6uTLB9rfu
rLAce7V8afRpNOxhRW9+VpGMisXY09cFuxOd1u5guoo3zLoaeuzAP133zL9b8uj0rtNGIUvuJQso
Gj2L+zX21QgchiWfIQshSYBCgnCzxcLCADEg3NIFcqlWW9Bxrd6e7PQeSPJTGACFJeGihPlyq8ob
qzlXURppFetYIzvfn0Vsw71Gg1BpRYQRWFHUzVRw6D8jpCxlZ/X8QyG2BH081Go6SmT1SAwhO2kY
kL4X4dSbA6xQY7UWRK0+AYjBiQJO9cfX03w8DaKpq02pYXXBnJiwH6sYrWW1TCEf9jiQ3rh8tJ4i
is78lxOe0Aw3Sbt+SSam/BSVPWQY88RhHxgrtoafZIjH74wMy1IXopLYAnb9n/hTKj92v8Lg0K9H
F8mxX/rxTqKeB9QPjORnsDDkB+5v+Yay3v2wXDUgMWcJrNrPoJMH8JgGpWFB2XBdUQmYgSpAic8Q
tD/d3mwMWBR2JkelLgX8F/m18ogmslhMvUJI0tJImug12gqPG0WVDUhP5UNBGdMjUfsoo7/odOEq
DsXA+q2EuO5969+MTcZxpq1QQSk82mEDcBnMcte5ohcra0ivcbkcyekYYJrohRrEkLHZmyjijSqM
yAyMbBmGoV25XE/MJrshKLseYPfSMbv3jlG7nw2XXHtRDb9FbK0PJFBU6mnQJidGk64cBDQ6h5We
gi7Lz/ApVwnA/dg5unPGMhokZUt4PKbV4u4JcxgvO9KbRT7/NNAjXlgknCMvV7NoDs5cu5C53M5W
Npk9Ct1ugX4hwd5hNrIxaKnmnPk7uD4SSXi2fA5nsImgXprOlqsssmcJkz38q4BhpwZnIvY0prWo
2Io7YA/Ze9YYRDclY73mypdEs6SSuaMY38Xs/IlFDGVOG97ZkCDjDbO6yEidg5NuklU/SB5tCFNI
j+zEW4SJBziDObEPWMt5tFaO4Xish+VPZWsGSyi5aem80xEjdjsnrL9MwJsEDjfQGAVGgqBT8qKK
fnOt6zg0FL/aZqjNI8WNz4EFKjwSn+N3pl7yAf0xwPajk0aa5/58ukbyjSt0zSW8nA3Sq0WZm/RG
PSdmOrEqyINNpNE48eI/HUe3Q+bmnM8mPOHJcfyrxjIsdOO/uMkWtHBLl5zKm9AbaEyM2EwXzjgO
R5G5Ksri9eUf2PcQnvcHu5yyo6Yp7Cp/D1Tb8+fzRpMVrqb5ShF4QALzaaHBWFSrt4JUgXFeNDI4
yXUhw1mh83jsxQxQzDUdh/eMw96TOvX02xsthL2H00NoithL0uLXhZla0yLRj0yV5Og2cINFtvYg
Umt05SQAAoa+XCchRrHnPsmIDwjR3m5UslsyTPBvfMTa3PMnebLEEzj+TtldJ/wdocubeY14aUI0
7TNEjwwqHgmVpZZydJMIVW/frflAwMcCEbq3C4WBv6B7Bpceh2CZ5zJJpxhDzfKIOTyrhRg4xd7w
76L1QhKkSzc4hy+KWXBfDh0SeC7B7JozGzSsRjO/MsHr+3lZwGRiZl4HeZSneBUfwFMujvrSgtjf
x0FtfKFb0z8GLVNRw0V5UFC0AD0h07f6figULcDvQRBloV/NNGu3JVlt59PVuhySX706Mv+OdkAh
p0mzc56r1//PurSFzQwiTAJ0ySN0jnJMQafPDuzEtQRkKqvMcUL54aU1jdOdQYn4NEXFmtbcc52n
kXKV7F1Ye4jdQaUgpbSeISHRCW4wELIQ/J6eVbvagAO906BlZ6XkqzKOjZCraorUTR4Ir6lEW35j
LlRP/b0Ual+zSRpTY7zCQhZJP43p/ajkWXzDHOuw/mxIqeBNbGMCVBW2EnviT3B4Xe+GP90VG4LM
gNqnx8g+G9jT0P164HWeHVs7F/zVHQ999sq0uMBPPU5zu8uWJExzHV4xgAEg98ODPCGXQwGE3EB4
FsUyPAL1upm5iLSwPnqIs/sStydN8/7bDLsWdlIKeDJrSCbgHgWIPTlZJeZoQDC5eG1QPeegTo3n
zNwNBwffRhZBH1mf6NDoq6MjKFAyG8ViaS8AoBqzqip4lxwPw1TPOP7yEui5GUSZgeUzMZuU0mnU
pdO0QUldPFW7/e3l5muPPAJOade73LVMsKyFbUDF+0GFUS/Wt9JP3qgYTIzWAchtrTlogFiO4g91
HGakne9PTu0Ik1nNUMTTeFg50YEPbK07fGFg6hgheGPcWSUGKcwqXmOSq642qwDCJXgnNw0/m9FM
gcQDSrlDAMYn2T8EsnuKsQaoNt4DgNmIRWva1I5Rhe6p51dz0Z/Dwcqna0yAGu7r+xj+F0NdQxI3
Vjr8pse9zYPJvdpzBieF7cuGZSvtnQiHNgC5vvzdNJ738OsRYv2yi4FrjJ9Gq6+orBoCHnFadGcV
qq2HlmSMgla7i/k5CNuqmdr8He4NmPfEmkZHNywDMbqjHb6/34pmGWc8Lq2GQLomfoBkvbr6DfVt
PX2l5jK+JFuL6moltMHM72O+g/BXSnCltycGWlEyVKdtM5smhWIgjf+ApxIpSuHYLkFy/MatI9RZ
8fKlgV883IGjHDU0eWVh5Jt9K+GknrarEEYJfPnpuEb6hh/xOhOpSRV+zcgLDQyd5mTxEvfY60p+
/+GOul7dMXgY9+STnb2R5lOC5RwaMCrmCwVsVCzQRxdqg5/pZe/JhBgF1WJEoTwpsenbH+n4MnTi
WDFdAjHN+DJmyMpxTAsywWh21XaZ6VBguht17PN2gKEL5872bB9rXnj2oRPD+5TJnoYCnpsA/TsP
FdtPeJVs8smwStaUueRrUpIIGk7gqYDn4yhJHgvg4uP5NloaTwmjI7nD3IzwbFPkrSyHo/TRYj9j
+rtTm6DP3LF0PSHrtFZfSOe43UVv7raVpGV/8BroDSJfMwpiRu4+8qOPu9I02V6seNxhDqRWiRQB
fvAMtp6jXcPvAphwD7Et1ELLzyeez7I4HXzVOewoFgm7rpMcAZj7cxcMj1QDKj0gghPhqUEgrpch
TRgSzQQcR8rR3Z2QPl/qL10M3/CPWxP6ZMMYxjaaJGvHnJrzllLmtMIi1BjmiHYTRMHurpYktpAO
6CoPu0ywh845wE0piw1q+fXgWc4z7aERU6BE444QDb05OnoqMFtPkVrSi9yAqwk6VjQgSa0cSiZ/
sMyoXwirmXCqi1urE9/Si2bzXFr2lkIEPWXK4AANNbugOP6/5kZ61v5etOS+/IUbBRAKVBzFBtWi
P5z63Cy04XuFPXnTL9Obt7Ihra+q/eooGZyw2LnJHnJ6JlCiecgm9+SftGM+jQRK1FjbaxEm/F83
AWWKWGJZ9BFkeaN0H+DHAlOcDcCvg0VakWuo224c6rIPEOyVe4ERJLodpjw1Xq/th2DqogGbkNmH
JOdXFCalDAfG4J27VteMZuU1KNM2H3xeL6DmneHBnnA5zqhCKIiFHQ1lufizxbqfZTekwUNgy22V
f74COZ3mNCQGEccSlHGU+wuZQSjN/XmZ/qelev+nKoCSpmrp+Hmc2G2rj39hiN0Fewl9A9sMPQ7K
oHFlqA5RodM0/DPZixwsFyGT7awxF0qouNJNUgMYXM5yvyc2bp7MZQJ8tc4igRoIGlfzXf1GfYiU
oAOaAKLbbf1fgt3hEZTFkKeGO37QzRtly8ss9sMBbtiLfImTdInzcThwKqOj88xmnJp+vpMQcxVS
griB/etuDySfK3nobYP0XQ3nZARO4PW/iFCZR66wYN0d+22Tl7v1or+1e5NtDfn2cMOMBrkf+9Na
oW2uYMa0Xos7g2vS6cog6KnhGSKzoI7Zh4fLqcbieEjV1ihod7eWtvMXvnvOqQyhrLZexR6ZPxOL
I346rIKohunaDbcYy6t25wz6M4eyY7MLqKK79L1nlZsHvs89Z7pL43qzb7+/wBe5IvBcCfDH2B/W
B/XbCxjKXD8I8cEOux9cHoxMxE8RNLvalC/NckNg6PocvOX2gbM7YNpInPbstnqpbTsXIZXRLKHc
oFe6S8FytA1ILeBz0KhIamKIoqFxGH9LxwECb2tMjlQbidAzz0/IeO9cCxS/6Hs3OgdkoIYpah1F
86jRwTJN8TzLX0nTFvR7aRBWtsf3RBM8bWnhcwXz/MMqEPeqi/HhYXUPYMHynop2Cmum5AfY+8HO
KapRjdwf7iK8jVr51aKa7cV5+n/ngHTs44j/zGxTSUFnxI1IgPsrP49djv5GPX0zLXkbwlgSB7/Y
PcCseRGczjRdLNaUPcMBJa8blyuRC5ROA2vCXourrFi1HcKzX98XfgmQeJRheN5Q/hPlU7Nnlx+8
FefUYbutMC3h6cNU6r4o0tpgEKJ2MVFG2Y+vj8hQjrHgfz+nllrcCW37C1VmmJovjpGoFd5sdaJT
Fv3XfFDCVB2bggrM46EIPZgtB/Hmebf/WL78vzQePHzWGwQXJbwuPszdSi+IjcJlhrOJLsx7G6bg
6Gd0Uo23uqbhd7/oKr/j8cHQCkleBoqrY9tnQIB3yuZGiDnABgx0ILFPfLaudbyzffRLgf9/bghE
nVbFDAOSAyj2UcNIo9unLsSD0r5TkqDTx86MbLYHQfo5zbHgMmyWB/yHp3bj9NDUKDjMZkOa8RFi
sb88fM6pjrRYkCzz7WE4jC3JuV7zHT2NRMBu1o3FgtNqZRa9JPKRnAPls5Oao8GnY22MFoox4geT
nd29moROjJpgYV3ceMdjRjxKZfVy8i1+pOzWER3f344pfiT1AY1b+Gf1TOVsRYp1ULQMijibPWhh
PoDvMWPm2+otl1E29EaNOBEZEyv9zM45NHZYS9VuFB8BziH5FrSfgdRszWWv1B+yn0UBmiS8xv4W
O2wHHJ0Oj1lfL6eZQCE/QVkLcKYmPrcrJLqtyp2TRdk5nrdQ9qHntdENHl3xaFLAqBsJ1Eyni2fU
txvSL7sMMSXIbJQ4vqJLijZRYHuBuAjLQ7NS89jf4G2iPhAl7wloGSPOIbF8dFjRBw9MMH3JiFDk
RhjZ/OTyqMywpnzUQLJ1Nwx98SjjCM4yNwLKKqvfroAsbka0vyBl23Dd7FsS+y0lqCYdBZ9RzWWu
tKDUw9qLZr4JIdGtjlzEqwPzMWWOzjf0YVbXHzs0EXW+doSLpdYsTagHRxG8ZHvMahnzs0Y5isnh
wwFmSDH3cv88Ieirfi+GHWuyGQTu/AEAKVIFIkAUaspIiJXQhcJvQt6yMR0pF32ZOBEJc9nKynoY
EbGRe9WapqlqmN9pxwVWw13wJff9d6byIJgHUIqpHHmd9Lzvxx3cQJxyG2xdCCPcmYvZYzDxsqAf
KDcaih2MnWtRp4jB+Xr3ieDphchUmM6/AvVmblBIP0cef33R90mAAIQkPd9umZSJ+59SrAcriiWf
8gYNLLo7/OXfc9mAq7rWN/9xpCKCgs0+6VGSySDA1HkvU5FTfTpAKtzo9aiLUQbjOzB56+JqHjzi
MoSuEObbzyTBtostqiTCM4MSbqh22WwrPmQIJwNB3q41sMlzpW7HehlxAPbmVnx9XrX1u4OlyIVL
MKGO5ERhCHK9McSEo+TEb/6odkLzPJwRfQb6GvRgVDEr1EEHPyelkzyHtNrAEXKPY1Cz4N2LYeVV
RM9IeMJJzoN/ulumawOWOISDumc9eBjruGYOYfFjp3tD2SRShDHS4Ko2zgLFjqhkpAyRjh1VnzJh
tBWNRAPNS4MIpUgWdT5yVhxv1G2LUCf3jVvikmqB69UzLni/XrSAXoFrecS501tTLEM+KjLHpaC4
u+l+YThx0NpMY4L1h8HQbL8qb0TJHLkzJd0RBwKkcK4K2HrS5fXt0xDIFs82RGoHsBSkPTD8/BWl
Qc6q+nu9tPZzG+UP8zqo217vX91vu1PiBijdSnJWEcIFjdmewPgC1ZHnH9/5sai/wei3yKr6BuZe
jTaYAVy9JHStFTqRKCURySv6NE0CQC2W1VV8EvSBmxWft6S89OewlPkDGdJCEaqxlKm8HKL1uR43
8inQ6lEUMADkelxuf5bo0+CH2YnhQWWtEoIpYHAmJ1RzXJdteOOo9MCTBw7zQjnFvl/cTlLK7oK2
RVpv/jLBz/RY9CHNSFzfRKhJezd3FbzDxfFyTbew+/IncP8/oHkQ2M/dOTZVhxpp1vzzsZQxJKyZ
mGiDuhQKKeAiPwu3bXCoKNlEJX5U6LPNARIuuWYhukn61hAFA6uqe9k9PhpYRj+obh1mNBtN34g8
tfDI8t6OiWFlT30NqO4hbS6BTjKdhxw4gWYHe0jYZygbUwIdAn4y+AhLVywHQg7bMH1YSCxdD+fc
WKKOFoBKMN5aqj5pUrSYuwLhDmrYlTKfVuQSxMPVhseabwBEOyq+8pl2m6cxGQkWibSJoN6I5hjj
FTJr7Xfgcq0yuLuhF/0xENCmAx+bcRpochz31KV6njxnySI5BbhD0Yh7y3HAfIsrvZTqlirrqAQw
vWYHxhVSyn/UiaN8d4YG7pbRL2pI1l5KiQmVcHc2cym1dLZO7rx4zHcz00HtxJVOERAfohaJH9yN
hGxIVH9kUd61D6W6twbbErnMeGJP1l038FIXj0Z126HvAFLq9j4ExonlQDSjjkKI2D1erc6LWEM0
RURl7vfKZ69suRNgMZS1LcxTFEzfqEnThz8YcUxORJJhvu3FItZPo2DvYcDBY9nX1+PM1Ur2URKi
wEkbmk+WZvEyDFObDShtHiW7BsKf6Amumy1Tbi5K53YtolfS9uFlW0aZLqXsmHaU/ODW/W20cPvQ
PHv0rKgLctl6Uue55HzlHN+ooEF16WdHHykQfwr06K/FUL6K6myLZR60XmuX5McYXhC1v39NWjw8
TPB15mxrPaxeAUUGCyY3e6ND1sVvlmWUgGswsl/tpnp0f9+8kIUSsOrNf7tx2eB1Q3Q2c0eGE5FY
kXjyGRwMHdDOsQ5L50zJ19pzuzlmxxQ97+NymeCl1Y4mSRJvzyNMKKYw1nU6s5ZJgWaZairqqoJF
O/WdWG3726WLSPjaChxxtW2DHiF9ly9ppm3vEY6NQSMPSAUwBlg26oNMpriv7bNHfeq0ezBL8oOd
hhOnLRqFh4OCzWWB0Bo0uN+ZJYPtPK/aF/t90Oo1R7QzAHnp10DUvIaIvnvkL2WoLXlW21kg9LNO
MPDXt0WY0J/jjXAbE7C8M6HUSoQGyub2l39kuAjDH41IrutKVmDKxNXttMI2jHvPHe4DZ6AH7kli
rQzdJ6h/g8Rf8fYdG6Yno/mAYYDsPWwHHCn5oH7FuVLLX4Vy7dNY8hItmqdw0qeQp51QaSzeqHtV
/Svid6sUyatx0o9e+qv+be3MGbK7nJ19YR3gNRwR69buPY5xgxxhwKPPU5Gc/idNojX7JcEU6PcQ
clEvnsxdHzbyUzGgcO7J+Lf/gqhZXtDc2SEqBjdVW29UYywiHgeX1pH4L6qfI6Q/DPC+4JaATST7
CUtOiPo8kc/xt8JTEHNVTBGcbWG8M0XjiKA3EmWtTy1rttB0cu7Gv4DXS11fQLLy+kL+vmchb1Wz
Z/8r0xj90eNjNmUmMdIvDWa3pgnxqsorf+A3c56ONL7WcY//K1jGPHmjQ84lur4aXlAmNPP4XyHx
ccD7ljmVdZ4QhjxI+3KXioIRdJF6mbN/lZhDATJ/8xoHAIUtFfOkqN/pgUjCz4khszgoX4P4KXlY
V5uP2yV0Dvtfeu5D2c1/K0TNYOOOfpEF/Wd3KafBlO0TQaVoBm/Y04YHqs5JcgJLXLlMH9dwCjPR
n/DNUF47g46xnMgLul3kPTFrZu6+d65Hsao3JMWg6Xnwx0eRJ2DL09QqE9Cz8VlzTS7+ZFIWRWCW
VJDuSxCJbbqAnzitQj7JDr4T+2IH33ZQs2FUDjAbCASwpa/FTtn5B5vH19ZSDe0FqlQtF8OSyTqC
90j2ilerivA5N9j/Mo03m+wsc9i1B02F/FeoAGZKh81DshAH/UYoUHpiCjLTlX/4r3EkQuVWvv6C
/oK+v8cagBnQizjQibZLHg2hE//xLCzsTPzlqw9llz/jjIHZD77gh8AJCZs7q4rsBNpLVHbpv4uV
4l8v0bh8gq7630IanVeMo36Xgn0DsADSDZ3mOv5wFwrFjiLqBzBUHfjyuvifzr14ryvWlE8qR3ff
T8gRaSiJX4+K3qp3kyN5K7M8EK55ay+IBIj5uNx2LmKgm6gwq1FOUyRC5YuaLJ+0nQ2xNlQGGpZ8
+ehOHRF/fYBsBpSA8eCwn8CMcBu/2SsMjZmbnSQQogea0+8yLj7Pp/gibYxM+N1lGLrfCPTN1XbC
rnJ7s7pySNBhm3TJ9CWN1cNAX42j+e5CHtdF2wWUJ72ICfgvc20xFY3DAib9HZWl0ZoWNUCC/u++
e6Z1U1xJ7ao4ArC3/YKBq/czcujiC+AxrsCs2+HHGwkh2pcRengudbkQL3o/MmLjYRdFT2NKig2U
E6JvMsWZL6zIUN9n4rJ1tyGZrgjAN0yCTsYV7HJwAfN64fA/SSbk6u7pBzhzduOrPQrLS2mfNXQJ
EvTLUuMwPkbIN9aHLa54oh02T8mJsIs/eqpKwxqKJg9Ilqmfw3561jtFo6hHBi8TOx8xR5g3i+55
m+El5xJSAstSN97bMNiGXoCSVLd524hWFLAqdjtECnowAy1t9e07spZzAmLE51wmgY+n18i1txJz
VSQwerknUsmG82LoCc1GlrrTJUcr5BlSk4JmnZ65WJ2OX6yUvkQ0NKxLbp8t1aZ3MWeT0Zh3McWR
Z++CGCPHlwf1t3zFucTKfrGcWBEsiO4cC7juB8ckrFWxUcywcwR5CpS5brTl4FYaCzt0I0c9Hf5j
eOewCSs47Yp29Gr9HlcjqStv64OydfhUmTUFRk6ZTOd8cTKSR7og2QPsu5lfOW7f8StbcCk0epQs
Y7NX1i2JhgXx5ACgHfJ4mWAfvlbq6/WpMJT6Vv1Zk2VhUw5+v5OJ3+IGEZ3QBsh//vB9JOwmV9lb
6g+sD2GN7V/Va7Gki7l27Ed0omJJ5JrzMSppVMxZPmdciEW4hJOjBrm1+xeZphwyo4kdMM8kmzlo
vEvnWEAW7LpD+w+2N7G9iFe1wNnJGwpE+pT1gHG6QI0J/+rKs87NXEwyZO4hkAumdAbe4GdslbWf
78FChm/6cibwsei4CyjPf2o7ROU6B3gom6lqu/TiL2/J+0M3j/vZf1GSDxpXHuaH+VMhYhRc98wt
QLyJelEjgOYefno8Rgs1xvzX73ggO7gi70EKpcKatF6sNTvWjTq0HOpZ+h5y70joiJv7g0FVcF2F
t/27YHfBY+LHU+ltUgz82yHFFkNFsaAW0TYQnbtsWaazir4oAoENjT800d6Aa6JljJkxnGQzQnhR
b9YHMQ3MOyeisb7Nvl90Vnhtk9ZOEb17rQmxVWXg/oCpTsJAirDuhVfhsepbOgNeK9gIt5D1uqcG
NoCPJnbyy96MceThT6ghpvK0BBqivoMpwcJOqGsByM0+k7NOKGpk89B6QvFWaGWkkYTo6Uxxxm/q
WcBvdWlt79w9Uxbis5N56rAdmCBV1m3OohrrNM+KeENNSvHQVxcDJT2sB1rTKznUjHrUpk8bcpR7
QEA9d6Jfe55qMtAxgPBrQ54NFFNbaDcTnv7Wra9cm4vkso+wg6jFasvy5An0J5XkqaUrGJP41YJC
QqDOy/2kamyq49jPttxP1liOwG0W5fx/hDMisTBdN9T450pffMaRVcVo+uoYLrKKOu2yqNMQ/sPi
1cN65IS9QloxZfn8MdO8mDvQ1v77hitFZERLgXJyTJOVXxqwnTBiPfQeglXCNyUdiYBmTdco6OZB
ibtQ0CR+yTj1NKUfibumGN28CRMmQmR3RSyjb0d3yg0FOJigB/2+k/I2mmirY35IdzWPEoaVKd7o
CIuFAZ3YY+SjzxGdQj9wumpCF5juQqRwffcgawGs09tT6mznxdf2ZJE13YB+Wv3WZHdfwErxqy6+
1dope2pJ2S6e2rAet+yymWB/I52d/tNnrKGaGpK8sfQebgbvQ5oQZaNdfJQ4zA521/ZoWd3c8H0g
Q4FQhRb/5Zj9Xnde4TdkG7tVNIErni9QZDDGPl1PzUk8jFuuGtB3Lb9zgvpmHEFSZYoQpsSAldHd
s/zRrsG8zwRD2E49Rup8TBlwJovj/XOc110voKfUaX1I6QgidaJuVVOTpr1PqUBbMaZhVYgRTKS6
XvrQYSFd7DFtDcixU5eLqzm1sHQXwVDSWirpmWV965ndAksk86EIU5n+FF7LQKBG6yxNo76gS2Wd
sppIpEQ8GsnxPFBdDrW3KdzFSa94uhM77WajphGSNn2bwwlK6Yp4S/iaPIqc1H/o5xJL2+xOoi20
t4mW2aaXUm9C161rMwrTXlHIcfBEbJdcBC8yp/Ku84cr8HD20ZPqAsmAAPcTWplKKcs/D//DLd4c
WfHDi7aHZx8BebXs47DV5Nro5MJ6Bjd24JhtpOF02ZXHu2mAubh3NsJfpTqecfgwuOXdJYUr/b7h
tmx3e3w9Ao7eUKxtJ3kDgI+3KOoVzgahYAMBvIFG3+BFpiwpQqDRmHovnYosYAGuVJHWfLxVeOfX
SO3vUYNm9JRUb3A+mjZiUF0QJ+fpt8iTT4jPsQ365grfcjg8QtPBUj3z/witNfCaHsrPa8kFaUBP
f8YP7oOfAPGWOgoSz3B+lBsHhhgkfE5c5DrvvxAwdWxIF+hFle/9fJl0Httm6Cao7YKVE9KUzoUY
fOB6RkdcPkn1YXvRelFyWh/EwGVkf6xPew/3T+eQo1S4yzMJjCTOyB69ZrP1FEvgfCtXzBj+rnM3
JmwjV4rOnPw5Y8e5pQOvYA6Y+n8h5lXwNcPCqnIn52/hog+cnc5nQYexK6J737Yc+17u/rNjyXzx
CpT7Gg8uQHo33AbOFZRyA8E07D4dM9M7w9niGwMiv9UgfYfblGWAF3rBMK+b2pIFArkyIeEU1T3M
pF2fF6DtQruZCBSlkp4XLX+8gh2q7Hv/MPwaRExLufh/h9QBjAjHPCu05HdDtD/MhwkknjpQf6HH
t9vpqLS1KdLWPODkCkYzM+1oP9VcCsWy04KEpIec+R+XTL2iygyrF6dr5q/NE0U1zNaZV8b2NOET
/ympJNJGRyVhPwQTN+eaVlotWEIlcPQgTe03FNkFQCBxPeXD6OhL7tg6a7XxuRFZVOaVHhTsipAH
dqC8IRElTCCShdDwLeK53ffuCv+luybal/XkoTr3jCpsktpH/qiHFbLDG9+mahkaaTi+awM66Sib
+fOYjcIUMEwK8tNtGwOTgaNRJwLOKwAVSyKFqWpeC+nAqL3N0AxXzoMb36hdv3fFN7iz2HmdkX7y
6M/Dk6veHltaoJL4dOuZW9Rj74shtLnYtvLWPBL6o6yyQD4GMOpZX3DGxBXBDfd4w+kvXj7iKQ5Q
w+pn1OLyr2bjvl5H6YA8nEObA6QKA5v6RBhYzKWlyOGFdi8QAl5IS5ADAYc2tQnyPa2z70Tbj5IN
TSAnkox1UolL0pW61fgAB8KL59OhkLQxHCJ39YwFblkW+tFOajhVinPRh9Bd3FAjDXwlzv2xALLr
m6ao+HoQj99PmN31UhfBqcEZxAa3d3wMwN3CvlbcRwn+0hNylub5CT4vSQVnFMMQ9PDq/iSWKdmq
9hLTRytIcNCuyoC3z5jQAoMw7POXmDnBWJETUQoZXM2Z7+HfJpUDT5iC/kIs9FMsZtnSCz0l3BpL
+exF4p4hiVsHBHNcRBgU45bRPiufPPisYIDq4cSy/JrTtgfzrLxGBBEfbWrpj1wc2N6bV8YpXyVy
Sglr/hdNlOaWxT9TA4i8KI1kY1mGIAHodJaSLAzjVtLYHtpbnWSBTzw0YOpjPdQHXbENdBX6fwU0
DrcvP/5B2nYK03Q5epqFXYQ8K7E6IHWazmJ2ixN+SRo5vcBYNPBwFTWijt1Otxr7tWd/PkysHKAw
bjLqWWYt60CfiRPSLATJGTIvkVNmr90OAURvonyC/Z5/30CcGoVNGJlNwlGFjmwsTqQJC30J232n
256gSjkHmUOgrGHqc26wjBPCv6UV3xdcKLVy4qU0iZvHfUCVcsJ7HobyMz2CImeXOliidJ3CN71c
Mxnp50EjfpD1eM4FA4N8XJnYpCVXmRpC2Yeb/GtnLaY7B24JBA++LiyJR2Wdow7PQX551O0OlGj1
c4vabZHjOaL2eN59fxM7tIezUHZwJOEN5AX3Aw8CoZGWCkkd4+0M/CSX39AL0ixal8O15C8vcocw
JA280Nj79PJxAJgHV/bJCEjkm/hB6PRwqApfN11ogDS0wAFmReBS+Mzx5dZlsHHzOLmA5b7JugAi
QzDvJRbN3XiJWkqFj4S1YLQaKmrRFhTgcFBCPWfenJUbdA2oUxydBqsvfXr9CSK0JXsIR5OdvVah
oghAhl3Ex4MFhr+cX9rrmrwumMFt/MIB19pt24x72Kw4ImHPI7qK0cEhgtCK5SPZBi/S6D4WDKg1
zV6ouQtywGGfbO18UB3gjKliro2qRzXDU1NUWS8d5j/3jotMUZlDotH7sIStaPIGDmd9t4vBcU9v
7B6x1l3tZ90+KEVfE1XIUf9/e+jg8m7LfO53WSOZNwjoYkkHvp1KLz3EZ7Moi4fdwwy2qz4XGpU4
8+7CDUT8UVWKv6F9nhti+gp6pBlwiW4q8EjWWjoqXe+dJM5xOTbpNTUQ21JPCfv2GC1UtWjQBdIs
LgbYARvdGzxO5OVGZAsdXtktoGqBDpQ+inqTB0FjLzZI6HazVOm4aVrY1HcrhS1YAYG9OeLV4tCb
gMab0bFWOXarmaR9sGHR4p9BJpbwH9pTjLVapdM1B/+2RuKgreccLJwhaQ5NSueeHfjVn+MsKK/2
ImwOIq+L1Wmo3+15p+qiqKoXOpxTAPmW0bBFUg1DX+dU65ZzUIcgQefJxdTJE8OX26AGS+D05omu
/911nceS46A5ungKW45zC6xSte7MCVYjCfk7jl45vd+EIYO9s8EooGdQtrM6a0bRrUuO0td5eg3A
+UaIsrIhYhf9pIlvuIzFoDnFHt9bzvsn2fclsAQkKROAvH/jXzut1B98I3x0XsRBy1v1By8t2D6e
ZqbZBdqAsgfuydED4YXSpratcXq1pIcJbht9EXlmZ4Qt84lMlZb1ExizAr4mSKFHpHRCxdiMbEQl
86VuO0soNMj9zPBZpQ+mxCgkoOKK4pEoJmEsB22by3a6zwftBpRJ3H5PRRI0t0Ek9svDvjIpyuMK
EnqkKBYx4LbvCGlom4OANEUa6iR7GASFjdkmpcZQCUTckCGB92PlogyikI4U7ykCkw1xVXamTxPA
oof13pZG1hC5uA6jqv41poIzYWt8zcVdI4vaJ74AsBG9JFocYVW1uktKgINgF7FPSnKkT4kXlTsC
L5OUlmDD+ebp7vDwO8MGEQdiy1TgivKKRid79hzBelkcVd+SrR3lfy6VXnZAmi0E/Md22FN3O2Bd
GCaxWaBrct0rQeqGPeEf76LuHn8ezOUEn9mC411Y5HbWdQzjRU3PyBBdgSUU9X+QG8dp2f38Sp8i
vS1uo7szKWUAniilhoUcW6hHYkBgeqgga4LCUsK1upRboBPfPwopBqf946htyoGZoTtxqv6QPoHn
W80w0l9MSYdY75gnbSXMMLSmMPF5tP+ynfp0/6O1m3tl/r1z1NzaSFA2cL+2rEfHKCXKleWsu/Lq
V5eK0VqDDqZih2shLv+Nqkk/MH8aJtt/T0BlvFyBVr/DUj/nRJQ0zF8IeHChlJjZYhF3wc8SmjPL
JX12njDiugS1wTZ+MvflSBDfTNkUT2BCM0hDd1F6BJk5EGS6baB8HoWZXLeVyScxP4436HJvUJjo
vHfTW5D1hOKjM9NZU8NoiVeT66SyC1sB8f4r5O0f2fy2mDpxf4WSCRNYI8ELvg+m2nPeZobPZQX6
g82IulMGwALUVBTOKjRO6Hshk4yEmtw19WQgUIlHMweTixvmTL6hzpTAB+qW6vP5x+4KIC8ctcic
kH95aFYHLDMuMhJjXdsWc+XzpxR6pOiPPYW4odT9lK2IalO8VQz28KZxUPtOv6Lag4LQ9fa69xGx
NpoPOjOov9U4Fzrv41fy7nFn9nOkzcPXjdSRhK6gRgFE6LWpxaX+7lKH9xX8Rep7zdUtj2WZTU80
EvemxKe9sWwNE2C6563Z0G3o49JdNe/5ZMcFTrGR3yGs1Gg1Xsu1vtsJYRE4aFbdY3ie57R7rWod
p4zTpFtFNvXN/incH/TBvkFD7z87oALII1UJ+RlwFCd7JbmZHrZUYlCGcP+ImjmCK+uoHl4q7xLa
lWbjfgI6IunFIy/bZrT2dQY4FQ01KRhSZcWnpGVCz/sCU/z60djX5A/+CBvSvfrHBpRPJRhR6Er/
z3KjgM3kUxt69gwPi0YfQibjD0p7tj5F/F+Mj+eGT9gHFCD61tMplFO0GSBS+PG2myvX4Is3aXOk
vIFxlrOsdFmd3gVFxlRJ/dNbnMSHMpJ2KPaOXKsTZJPwMkLFp1Y3e+JPjcEGe5iOk8MNMnP2+Fmk
6tOVBtNup/7Kql5UIljNgu8KPTEC8zQJL6clJo0OmJ+v0Gx8VUCHXEC/rPrI0hAAZ0cJRElTUw78
Dy383i2GZ7l+mfTl6OsD3Apme9Jzu5PxhB0vYBmcmpx3v6ySZSJhGnwmI7DQ84qWh6uen0NKnDUs
4lBGmEYOKA6gPxDaQXQmtHZMBeFUGwx3/yu6Mst0ov18kuTsrkHC+FfS6j8j7rqHjTf8DkcLjZLE
nALUoSZKSrONgvJjMXTGsdrmdmfrBOWWbO+AHbIm2Pu61xQ0S0ZZQQ0Bhi6x3Dlwb6/0kxfHTOAj
FJDAyiqw7Kp8HoUCuKYvQ2RVGrUeXUp0D3fZOaGIWI6sT3FTevSF/0trLLvW3gS50BNppGTeU6eK
964RW+nfSj9fiqNdrKZKVJ2Lj47ji6US7GSRoUJpii8QTHU3zVklMw4JJFsgjWT8pJq8pFPj4XWO
AQOLNUWj1RfAH6vxYxhj+yD7UnXGta3Y/Z4qKjqeZpEN3p0DMYnXv1L9v/2WvCJkWWg2QxYkWzid
sFXZZv6esL0jwjJTKg2+rcmhR83ZN/Z19XRyPx/Q5y8Pw7ORvhSxAMGuhZm0o/4jGp6PBeExHXh6
YomfQX30CaL9U4Bei8eAEzPLkQQur61Zgqi08VOYk7k+EAwqe4UqwSdDqc4qiRaFFJAyIHB23iws
NW5o9esLlEQFGgIvtkIUwBHLb2hkDseECgKzNV1nZHvqmXFpLHGXN7681IZ0s/KJ62MOz9IL7G78
0qkxfGG1A5d21KZd7u0orO8qnljmi13y0luF/UY4BA35K2OpBkv7Oat6hQkvYokZsrzhsr0aG6HQ
QU4EHwR6l5RDU1h/dKhTRUNEcs+dZ1uigUi4OpSu9hZXqFPRmgBTr0t4LuNJWs/BXFhOpn0sM7Qf
tXmHivBWdX/9p2fL6jGfEXG0zET3k6vxX7YSxbjURXbm3gk+CDkW6q0I1UCQHBlS/VzEcQwU4kDw
o5pxrehL8mN/uMgs05nPP0WWwKtbCVe4I20Re3LF8fUAsmLhbewDH03Kb44d+pKRPKWOq3ooC1s8
pdsg7FFiTkIsf0cg7K/Yss+TNidd8M66SQ+vsFIH4TA4sdk/CB0JLOLKm4NntPmhX6OtfdvFRpVy
t2TL3fiddKS6/OLED60sLnXOpVvGGWBd9WsB+rYpUVmFngqvpAcIlVuX+C/g1TnWZcgurSvn4fem
Oe4x1Z4He2JoVwtwoG5mpLIaA9ZewcBsf9VQ9BwdIBYZM+B9PdyMdmTnmTlUKxFKlH/YabYFCi44
bB0lhmxgBUMzlHhjlItrjj89JL96ud1FsS+KwQ96qu5nQ5+EwYXri8au2onEfxCjCGUoXP1sBsIj
2CYogRTvsuH0hPUA3K4/ICGaY+NjHFUtT0T16QsxgYslOUoWBL23NdmWXjRUTR3XERjuFnRKXK9e
YOgxlnUGsU/prsiP7laGVUQERro/LmScMGaHxD6kciF7idwqQeIuP7gYXJyNzOGWXqCC1bUX8Gqw
B+04R2bspKewtTxP8SiL4fD56n+zTA6ceND+NyYdRoxWxnnSM2Eb5HzExMydkt8MoD9ZGDidffI8
oe9Eh+OBHxv4/aiio/3IJRnMud5eHj2QRJDuF6VJ/X5QQbTRxIXnfrHjuJfyK9fWHBsfUnkO1V6j
eLhV9W0MppgpV63qfErl6Av5VbZ6aiakxtCziSPV91bqxyHpPDcjmAqz5gc33F1iN1Qxtcuj9FMW
jDxQSSCcJp2gITDWQnJbAJ5r7z9Y8UyICXm7mOds5GYssdXU6DCrrO9XmRR0Ua32D2VKXUQ5Hh11
KXbXwI3wus0fh/CsDk1EWKBJHb5Ep3NofR6leyRtXT3tTjL9yWNU7Gp6NkFoMhWRiyd+OtwSZP7G
1/UcsxQ5H8Mof3pV3Y9W7HdFrMb0v7N3vZ3vvbP41iZ6YFUFvYO7Pw3gGnpPotqlYEJVjgORW77P
cxScIZRQ6rzMAVEYS0ik7/90jtbIgl7RByR2bMN4QZwOo2ib5pDyLSzh7/9A60kjRNjkroz9W1JM
qMaSLnv9FR8lwhxGFIyiuUwB7UumesLm8Ynti4SGyIQ2tJTNl5GYnb0uBTwjZl+z00YjK2gPFac+
CQqIrqZ7tTz14e4hWeqZm50v/p2xi89dZcRlU/tlxL89tipwhDNhID38iVvmczoC7JopM0udm8N0
IkvRqFIk1DJXQpHWMDJ/NBrPsBXD1Q9xLobKhbSpy0bPKTaXMe4fXhoGWeL8JhXVd8qAYq1CDiXo
9KMPXwbQH9IfmB8s7hCUCf7uLkJawKHUZ7hnNxAB7KQG7od3SY8I5zCwNjWE1tqBeRTtlUNnIjuU
fvTQGJtXcWiLGn8eHbNf+AYA1GwHnViKQgOj5D/NosBoH9RG4KLjrM4Qdp1TNBpyO0T1QzI9lWmG
s9WbbZI0LFZTDjd4i0uvanfMuwfwjFwRD310WCWY/u4uKQX1Ykxvcg+6YTJVRtDOGpmMjPirzLMK
uF6dB7sF/7+RdM/8PuozQqQ6tEuKqhB4+5KUzBQ+CZOdb/m4weXuwNnlNlgKPIsugK1sfjE0HGF8
oW3f1JqKga5oUogD68HuY37I7QeH7k5M9qj6+XNWcxHI+sdc+3frHLrEUBCBPM+2nRvYZpdq1R7s
F4Fu1SoCy7BtYojuWLCJQCcAaFak8YTs4WjGPTWQT6oqzwWGsKF0C+ZgjLl9hqJ16GDwUh9zjDzG
voPcLpMWg4lXsJIn/x5ziwBbbluh79tPCbXXWnVu4sUbPiMt5Ew+rnZ4B2TimbaMI0/I6XlDpzvE
ElMboCfIitrxFjCU6i5MZoRFaD/oMR9jqD9wrZZ6FrtJv7hLVo+lB2gqceXoJc41Wow/gB0p5Hiq
gkuFI5XG8fmmGCLI7C6pOeXhtB4N7c7hjHzcbrSLdYjBNL/gbuSzDAHlwY0DYVT20/PelSjDIKph
WW/E+gSaNXpuL4UkIYLQDhRMGcf3LfAW8pBJTvC2Oc/KviozHf8eOFm2JQo6Agru8Rme/7bCUn8u
kt5wltkyqQ9f3c8R/I1CVDvm+kBbeh08PVhGUcs70sI0CtO/OcxYoHEnQd0Jy4y04mtO0laA8cgN
JjrLyjtvN2xGqX/zPK1QXn95z7F/SFJvv9j2OschFBqyyzqjkD62ROvdQginOusHvNWLMqJDdjz4
CuTPyTul5BPOoANOrB5R/R3loXo1pz9WO4TF+qHRHoVYW80YJuwQCWFJD6v4VLDqFkx00Bg7XWWC
ngE9jIDGDZmrkoe3lUd5ID8b0DSWYfpUcCEDKf9GAxtEO8dzsw7QQTMYL81FN4/MMG2k8sAEzP0e
0yAOw73Kb9QKIQxbKjcGx34ysH2Q/YSrRGPoxX633v1xaAckcHfCrUQLVa22qhlQ10vGEGCROxO+
sv9Fpmib9nwtYgL73JsDuN7Oo6VFaHRmbanssdm7WdI69vvvyPDPKNSzcdB9+uZpVIkb7Lh8rUX6
t+Fywvttdqy2Ro9NtBBS6aoRUWRGKYeukJ1FtqYVzp1dqj9llu70QhUA1QKox8zuqI26Z12ZyjDu
D7boWo83cD8AqUgA/CGM0VhqvcG3Sw3mOc4XyTPZLwBIJnyHfHXrjrvS7oFLhCaRuV7ML0K6mLSb
HudFUf254aIan4x/dCIyVKpa4nj2T4A/knngqajg2asQSF3fPNFaqjZAb2Do42zBIuWvslRMsEdt
kqof8rHzZiHaNsKfarWkemKugD+gudVi+JhdbQHOD+RZ4WT1vIYemPFmEBO/tO0l0ez56VZBMag8
Y3//pBadhQGZmmXyh3Eo4RmMyXkxVHkRwYYUX6pgnpkxd+3n7Sp7bYdeFYphVRa/+VTvCLKkhtTp
u60jSqEuZeve0C/gakaEzFFTvyd8pLbqR7rAo1VTEnxQ0cpxw5pGywaOw715eRc0zvXs1UcDmLnK
/B8dMH80de645cOGEjMHa6XuioXtPJxiPzRN0GSLBkfaqPSU8yIX6Tj2JBLKO30J6W+1ahuL6U7Y
XNRiXQ/7mZ1VcVkAbuLAGdnZRj7dM+lNO419yWE3OkXfLqGmGjRYTBnWgDqE4cVjLS4rIkKZFdIP
TYTB1ScJElGNgVa+/FS82mNO9h8aqefpOpNKy6KOlDmp7Un2fWGT2ThkL7rrkJLdUkWDxz6Ux6t9
BsDn4D0AFOXDkitvWcibia2m4oMRVu3LSeu8+f3GfmB+/5iPbyiXHQ68CFs5+K8O5zAcsjNfHXfP
RAUleM6zwTjiHlAFC+5+VgpCbGCwGrOi4VFRVxKm4iSQK5NgZUfhp8WnKJ5c1h5TmrnSJYuUa8zp
aLlR58hXYfkV1rT7+AZLDGlsWU4+eOa2bflZ48LuM9BO/yc9Cu1kVHeg9znKK6q1evVleKNItTka
HoZM2m6Gus2EFWnUS96YxHLTRqqtMesoFkptvMcRtYoXe7YbpPr1DB55NNEu0sMLPTA9/R811JeM
dUj4E+u+boYFhqmfTmG4M9UKlFxbQPHzExERPaX5LVUjIhtzfdpfR08i8SLVkg6mqW/ZS/xOA2Hh
ZLYVefB1FgajT0O//uuXRAUMQP+9URNzsca1j5yJN62AxbX5XgYHdfnMcqad/4wnZ8HsDs9jky/I
McbHrh3uPqb5Pjrn8eszmMA2GUpBa1oqe3okbvslGObBhx65sV3D1iwiWhg+bQcw1ToJZunjs5P1
Sl5CANxPbuvAAqe39zYYqlyQofJMKflGMiaHAi0Gh446M8Y5YeiFuw/rnF70zD2zOly+watBuZbB
Q/4gPxZHmKC1+qE0U8SOq5EOeWeS2IkVln3fCoSNuUqNKOlyAFxeRubNam+oaNhH0mO6tl35g7FK
lpzNpFwWs9LDE5MjLsrXAfCuEZxZnd8ECz1JHTbV9qF35/apjG1YlsxInXun0tsFQX2m0wXrmnIA
eesVE4SY3NISivWNJV06CtNXTM4kayHGqI3Re97G+eEzT/uytf+rW6aFJCjSJgs3DWP+uJDZi/BM
0nUzNjHo5r5z2s+gDp7YjRkR6kf7J2XIiLxAuhicLghO1VhsZmizisBvPOzEQjA0mZNrnFIV3yjy
wEXbcD7wUPKZ6s/iuINnFyxKrhKQRWbTfVNMIqfVtr9+LhtE0/Ju/6Uhy585z41P+GHlC9ELS5AE
8t/YIqFzxOyzdKAej/3+zGRy3RY6NOY+HYUSaUKDJOssMEXGB12bfAmaNE4kcc/kiPCRqfISNO+j
0dLwZ1xxxiVYgam7jQn+qVR890ml0RYXUXHscRbGrs/+OSjMaUaYqGA/JHDN2M9Lm20tiJn4lZL5
dcWIWybbW2ot3HrEGcGBv9u+Rv136JmU8JH8/Z1OETpeqs4lK7cRsEFbQXagWFVFMr0IOA56t5uT
PN65kgAlhIZizYgEthE681+T6E6gvMZINRQkIGAE6inFD7lUWoTnbuQ910uL8zygbjt6SBg/thoW
0hvzbdCHm1Rzm371I4YW9ZiKDcMS3XYAvcSPldHOBCXcZ+PxKkxoDbyBD5yDHzwj8X7lQar5HjrP
F/yIR37HPzRnLK+fLt0casujfxtL7F8dfZZCPhx4GzrmNLgse341a1Ym5aoHQdW06+351J2d/CGS
7WN3QdWBygH2b9f+Bhg5/hxz286ovdLQwmppBl2vjqzdBi6MNH9YOIm2bQzqK7BuANAPEAN8h0no
Fi6+64TA6UbTfUxY9Z58qubU1x+1edKwrbB5kyW3lPyjtm4ETdnEnrRAsccBxJvm7PELbTHBWoPo
Ms3TWRMc7Eex0K8+8aNcDWwQ1U4gclhShe+r+m4cYPlEZHd/7qqfAdjTVw1wfrLqiqDND7G2m2WE
A227AMDhrEQEpb6R5l4BnKClnxy22mIeuEuc5Y8m9OlWJv4cBYw57IZJPjKdLFH8F17l25CITELe
wYXFH2c+DyUhO6JTzpUn4S2uQI4nq1doq4csBsHU9YxWMEB9ctn3YKk136DLGni/qTQpR4pr5+iE
oHD/RLro2eGEm06cyzMtQVP8UYPxn0Y+llGkD4gmyFVAezyekdbqE/xQveU0sLYeiv83M3uKNEJG
dJn95pStyxTpXvdZ0Uaj2owndRzLEJGdbSLet74mp3seNOnZTShcSuzKgElZt0BOlJgWl6KeK2FL
9bAbKIWLdIzRv9L1LN1WNT9FYk7s75Sf8xhKKE9yRemH3PlE6pRW+2ZnOCCYwPnD9yoCuXHe5JEY
hnQGR7CJ232IZC64HU4kq+VDApU7ejBrYRrRXn5pO2khg+RhO2DoUL0U+P3Z2tn9flFnsYVsKPS7
pzcnMWNUIhSKJSKv7zLjeqrqeWra0LGF9bTVXd3ZL1mEsMnCkSpaKI8lIa9LrpHQvd9kiy3CzIUz
q3pJZFkEUA/5HOVLGj5YhOu9mbjGhx6ywIs0/4+o+HDiTrDroL5k8vGvsvFaAH1OeBXLEZB9wjeT
6d/NxKdDwDouOJC2S3cf6+FWarsf1D00hQxaRGw/VMElKXw2ZasTlhHjQ+4/DGNF8YW9jTj7rVsw
x0VOXn0Bztr8cLNC6MxSsav1r/t2DYP3J32XHu7k51SDJwz2GDwiOxdg9sx/JyEG7xxkwuPYcMdA
59oPGnVuUs5Ad9wdzrrsP+IbulUEsAP6fhXC7G3oUerSJI2tUlj/e8dev0snhmitJe1HdI9Xqzrf
oh7rBBDZugdWpHnXzGhfYnf1jEuJ7TGDHXyij2BA+62VyjhCoEPRrnWrV+gXFYpq/8LGk11KttOR
d3/XLe7NSjqxFwpj7mDPzFwP0Ht1GQ+VGCmIQ8IDpvDRBNiYgdcw8wqABf9Rnh08YEGNrYJ+qUN0
uuJWjxHKsY3a4pOdGyhAsIaI9BIKwKi/XBaIvp9eDPJU4qiHf2rYLxKYt1lmZiJ6UgmwRZP/e0Lm
NxcaC9CxXqbo5yhs+6pFAPzFT90DLU0L9ZQbEuyLzrEtKxQxrYM/Acl7/EESX2h0pjJ1LRZnoAFW
hybbUAaxu5A3NThHuqe38/N0jCMdGGY4EyJeUXyjOecmvSTFrXvLispb09haX6eRNb53KAiDYY9/
2VXAHB3ajDPhsG7KPVE8qr0UccPQ4iJeT/zTWBRQYNal1maJT4eF76jv/rKZnJtoAIPfLmw03xuA
2kOmcigcwLP2oXkiPabrciPIsimmtXqIaoc3+yWvVC9d9WN1GZkaV/qnHzAaUFoaSDodaH36GJcD
nKF7uKuLtDUVE0JL0EKA7satmjBMRceTqEQUx6dpc7XFYK4+Wp7KebIPvr5BXTEkjX6dKbnTDigC
Fd3hkTUF9erXUdz+Tt7kDEjS8PSxoC683CjErG21WpgfJ4KMUUQXQoirCxLs/zHuaWtRdklmYbBB
GQm5E+w53J1OmmYReGEIEBmDYv2GjwKGUdZof3aHOyzXd/XycsLOKc7bTdfkBOUnuBLiYZDkjaxk
H5iWwScIXYoYHjk3qcQZIiuLws8zTiRZtTFaA0jeisBDddMlKhjkYimzk/icpdKDTBnMEzWqwMgX
XoJKMXmyDAU1jNv51fLdDNgJ44JcXSyXQmszpHLaUpL6hze6r2I/Lm0T3CD86E+uptlr3l8zh32G
ON150F4qjRhfJT39zx3BSXmljPfWN9kU/tOKm/QENO2QJVk5jYCnGXo80PL2zFRWlcGDlYrSxI4s
AnS1U4zns2NtLmP6B0DIpRGdhrtBLPm3SR7a5iXa1hBJ2DRULWu+PRC9pGzFoYgW8jTB7a+zA6N8
jH3f+eTBqENV1J8ZWA49ohfg+6PHg6VHxcYMfzVFlCUxdOZWhOmJHB3wxjjA7aM9TC3W+iB9gXXw
Hq9yNDKX+xZX/VfyiHnbKsCKJ8mNrOIn/04T9ZQ/Ly2ru3D1fRkU1BzBPWA/0zDlQW52OGSuLT6T
BQ7DOVw/eQlypM0Hx8ne1KffSxXZfWvHFqMdL4N+Q2xnuvx6C/GXurNupcv2QdWXl6a3cN2n446F
kHAHRSNWemVA6CninNmxH7WFW6/0m3qPoQyM0kfOkpuRorwn4xxCeIhSyHL9jmqSIp1h2Ped7pGb
1B5IW6fDL8oRpOMdf3+JaDUPeqhELtsD6pXVvgCHWiNCGNMJFv+zq1wQYho1gNA4h8hjyE+xP54H
tt3yIRkJDFZyNaXJEeWDj935oEMrdxa9qmz7nOopk8KB2ixH1znlFl9Ure0Eo2RrdBl6SEQWc+Bf
2ZoV/cTjx6Rfcuv83qPcabsm74YCo9lNBac3ASarbBfrHXy0Gd9OyaIxelzvHqazw7YRvC/aKroX
iePg7z4DBKviXzxYNuxL348Cq3JkOpdrTb8XMhGDiAAcmuplFG8J4ty3LcaUwbZaGivUOKOovkK/
o7g7PuvWvhQomNMuo1OmrBpRn475QRwXzXB9+rxy6YJJZ8uuOJ8qW8BvDvkOP1tATPPq/Kq+ZJXr
QbjrtGG6QD9YsTnEH97/iMk8i9XLV0BWy2oRnTWhROX0BfcmbyWfiHtV6mPV2oG6ZtCqpY55iBhw
4lprZ1NHyrFVsq//1+taS3qMjfHVcjrJ2EogMBd+Jk3FcwBetmim27Y9Pzku6F8mvZc43IN946fV
CWjti5tJgNQ4poJkH/+VvHeNvuXyqutaxVOKqrHqKTpzqF30kAnWMSrPuBvC0qsCrijSlHUa8kce
LicDOxKXkje/Qm12KIeSk3720HNgktunVK9Aukv7/tec0K0DqscDz7kkW3Htlq+2RRh5JVInt9N/
EFLvRlhw6SnKE4EScejjmmeu4VlsLTcrbhRQQEFr15IyWWIneLujSBQcxcvJqQ01KW/9esHCsdq7
6ott3Cu1EkstZ2AGMmxLAiYd8XADWr0EhC64D5DGbjgISdR4PVx/avwpQVEwxWCFbtJaWGcoCPpR
UgG9v32CKjoOjEeSzNmEFHQef5/CHCCVtqLoIfliGdvFeeCY+vctoSld7fznFfseeugjpI/KcPJY
vOb8lulQEDlb11YFt5B2V+fDt5tK3XYFRopmehbuxtJP0yjB8iureEToaPx4M3fmr8MYW/d6lT3s
pVdjO8RYSp9mQwXFsGWsGWNzI7fbpcUlE4e4pA9OFmzXmDnJsvNiBCod87VE2nkwgAYqZ8g+hSCO
HcfBZCN/CnXKLyAYhg02xqIHV0oUh+sCWIPI01YbXyGi+lg7JKuyyizc7H4u1dYCJace7i7fBkYQ
HqDr8cgSCSmL+QVdA5T2M87HCE+YKKNx9EY1Koq1Vnkvc/pzJf2Kr0k2dJrZkzRcVPZ+7hxT2O+q
2yGnA4ekxsDhgyD1fzF5xTmaF71Hwq7rXfZCnI3RRk/QmeMLmWW1JKFdzRhl3P3kcE11/S/BkZjU
SUp1VL3XsFWOjbH9dr4cJP/HP++ePuqxjI5OjSnShg2WBb4d9Q/IsDF7iAPGQkMaVtB9uj3YJ9hE
YVw1mg1En8hkOdsFRUSEtdI6FGgiAYNtnX93+p3uHWMLXpbVGQ7W3KY3X8bFSlNlLbvlGqU92Fqc
x7f/9nxdQfpgYFel5wqe4oK8X1UG2ccex4ytusxfFZO2mHVIeCcohNaGk29a1nm+nhAlFGzUn236
ctkUgRjCLIdKhZqmP83eIQh/PZyqTYmk4syt3ndXYef+AQ9+dPIboCGfiMKW1/KWPRCnWwxAwK2V
crgqylpR5NvJGkvGbYO1QTx26SwclZlAeOM2eCgAW697ZCXdZIr+7kSWYQAOMU36t0s1SZchgaMD
3//bPixLTDzZp2FRma5ZfAgnrJy46n5a6yUMOjVhnnZ2GB6PjX2dGfNNjTJMjXf3sCRust50MoDB
ktIZIhBiK42yyelfD2SZUgF/PSeBhyURwufD8dfia07a0w13p3MPhuhHEPUScVCvnhme780sazhW
Cr6naXVxhA0Q6fq1Y7Ycvj8guGJu9nbzrfQs+9f6qrqErW4AApfAiplDgDc+qkEJMhaF2mWDo7ha
4YggUeWov35LhEMfHJ65C1NUDnPdKzrGTfKgvAxVFKGkwcoWkTfa+Fpy9onvVRp9ErrKTA5oElnC
dzLXDuwZkOknJrb+Ve0pO+aQ7hPvbxSmWZJm4DLlqCCoRgXdMdfQdVTdJi2HMEF/5AtAtkR09Xl3
/B9bj8bVmrrLWf7TowY8wD1HiJZd4d26FIpRQwKOdAU6xPFHQwNeUzx3AQUmy2gkYN8ZKpRWn51+
0qMYx0pc9JWFCEopsxhcvoQtmY9mqIlBm0jcuQTNfMwL++JdDCPJIe+xZpYXYiMKL1G6iNela/3s
mpAqO3/V0wQCVVYxbpjgLJw8l1BvgAQuikVvkeVmpKORvYeF0UvUqTRq82J9Ws5xWCoC/R/gIS71
O5BNF9PEh6Swy/CDQ9tz6RiezAJjVxNvcUQfk0UJ8Wk8tMgul3PZuqtessQEshsnUFUKf5VUVmrK
bdSpG7l92mdUqxeP1o+Ec+0q111NvO+qD3q+EyyhkZ+BB3EVuWcjR/EKUVH4ZYE2xy49n+ZDyhTG
9ybgaMeThDKyICuDc6cPbEmQYdilMXXcwwEc5rpakcnaa0f4f6yXKc2+b12zO8PN/N8RgAZTHUOn
QrPJrfGbqmcXa2cdYake57uEdAjsSHOd55iNjSvMH91P1PsEdnkUF7aZcslf3V76HWLZsLazViHm
E9iJxxFqP2rN9ajK9D7huGwtWsbV8WG0tBLWJuAi9YQvKgzj2nvJX5aD7pVHgby9VJzoJRJXo8iC
QTv/XUdtu/AS/rMeTtm5yt5BKYI/B8R9SHORdc4XXNmq5AWmyzY3u6pLdLTO/uJr+QKcYJw1i+8S
ZW9mBgBVv8r0b+52sSCNgfQUdKYcbatX4d9Ics6avgWhhJ/fbkLLxUAscoU0PH5nOaYcuzhYHV0N
FxSWhbRMKUmH2eqpv1K9556pa9dNSsOR/+cS/GpnigFo4wyd1Rg3BIm+q1alMDsadDYVr5kD4CIo
07N4TL4aTUN24u14hQOIFKPiX5nXkBuIVUFLOe8rd+RX7ME6+O04YpvT2WUUoIWgf+EEY01e54gR
W3dbNoRi3Hh2XOf0+V1kaSrqbcxKZ3Oi2808VL5cyn6OTztQuMNZJs/E+GSumHEpndEqnaVP37Et
2rD0JPyN2Tq6Ev9iXLyZycraJkNflHACC5yhl+MlaKVPjVbYY2pYmNtYFHS/z0vXlF1aBo4aOAN8
QHFRa90WPMCGCEMB3wFWL+7lzJAr1fEa7dyu2BejxO0T355XTku1jX91kUtGNjk0j39M/NJFifaU
tjulRffPNdRhviOIIEYBWH4vR678+9w55XOsyhuRzzbafy/i7Lr16K0hIQe3thdGjq13/uyblVwC
ki/ncLdB230riXrnNPa1+hoFTJdRKBeZ3wuE40xcKT45TAcgJTVgURWhfHvIcf1Ur79EcbICNj+W
R2b3qDKO0Oe4Q1UDLyrmOAZMitmiJrjkl/pXjmSAxv0PrxdpjprHBmWw2hjw9sCZWv3ChLt16/Ew
uHSBeEyAYtHotDhTyKh+ng1wyYaAXPHT278Qp4JxMqA+U/d6Lo/W2hxzB+0ZRJJ1ayh0MbRrUyON
KD1Pv5WfaKOxJGOraAHlhg8AO5IRSdp1QNgAkoUNjaeSz7JlYQO0pu4I8rQv8F6EJid+cTaJY4J3
G87yr3iTiF/69tmFxwOo9rE3oAzW1TPmezWozyvHYB/iTSA3gvgueSoMKYjhlC/Jn7lNmB4GDwLd
/LxyB3GaQZ7TXTJM8w+7vUQNFnbFKkqtzKHe8GmVi0ckoD17AgdOuCYeIuJ9yj7a0oX21Fj3Gwai
+0itpcjmk5tTh3b2e5yyTNsINn/h0oj8FSEWKFijRjJh2KMKfyWk3nSxT6wXrGqHH/J2iOZmWxDi
YurKWQPwe3SGaCjKyh6kweaejO4WM3ajOX+/rXHU8D0nWucMFIfZoHI95V2Qm7dbCQIWS68UHA09
5Rw4wvTohBuIAvR6DVZ75vVFtUDUSZXU4IsyVoJxAngDX9hPefu58lHinxNqEK1/emBEkkRTmUKA
ftuPSGmCfOhbYtH6NApc4lNxZlvxOCfXwMbCVpF5tYpeSbBV+EeO84aXgUc11uwBgQbSmM5bXXIt
Ei/p8L86ICaNo20xIsMjIwEHIYQ8HoO4T6zUxd5WfXPkvEg8WCXSVGP6sO/DNk2SqSZ45nLvzcFU
IyjIHQZ3pAc5+68wHMEuDZO1IGjwJ1H3rII8GoMOESJd7u/kNpbCM4Ww/ipVZHBd17mTLjx6+Wz0
FCFdhzmDzzASja9DKdoIf1Y4Mpt1cJGTAM2UlaxOWJ9XoyfiHwRJuA6UkRhw4EFelvKj8bWY+jlC
3xE6PJNTG+uH3/iOseG8TX8nnd0mTonoq1mRbiZBDkmdjrYy5SCphaitKe7A8tlRM+vGL7445KzA
GKthVqPaKd2G/pdQViU+XBWIjGilQ58zIwu7bqdPgey4Zr7PkvP93pX7yedgofi+OdgMySs0/1zO
QN2YOxXllTWHCTC+7CAldbw4ws1jSIZvBJ7VBun5C3YUjppdwKh1XyrhV6zzXPe3luwyQaCF20BL
+k0COAV3TXxWfXNNy9gGO6UrV6X0I7HPZLjVvWDb1p0m+Ur/8UQ3sEbyFrs3+j5ruZBx9L+3ZgS0
TM40ZztLZytc4h9Tod9d7esFozwCbJqVaAWQ+T2hFE6kcf0mFcOijxrLySD3fEntTKoMs+I/khE1
qJJWZjVtRnphT5dp7gpuR1qsyIfpgegqN5SdEQYrEgryJJKVdDzD65nxHbp3H70+qk4/nYBhZQeT
NUceX5By6zgEyUcimdZqwLnhF1S0Q284GyBJ5b1ojnNz7JTnG4lOMi7nQpPROsyjD5kwD4tOgwS7
j8JGuSK7YQIuOjB//gfOY5mjf5pMw9kbcc5debgG85b4aCjq3hd33w7fU/2dxzC6BFN3P6CXudey
Ac/w2ij5/ez1qmnIhcynbpYE2ECfnliTlWRqxoBnCIJZfKmq+4VO+wb+C3FaXjoAbAGXAHQWR9U4
86jboxMfAaZdiKLQQGxhnMhpgptd9CYMB0SaMCJQi0eaz5CNxLLn+OYQ+3uKsOrhbw29d4ZD+WJd
WGGPg2XmgWZO42CKfJRMXtFInKq0yezueJkHkGM3SR07PWicWJd3UVV5Uj3tqhYLkyraaUmGEovx
lCAgPRGgyNv8HS24CGcSXmtiwomxCj8Jcn3wxrnMM3ASb0lbxMHyJCJbddDJyuIYL+mh1gAm7dxk
XH/LtTh5sOI2dir3VEbDuS8Tv5QkJVpDfsLFeIWDIdWS+mO8ui4NV04l04OmoHIZrOK7S2ooJnPJ
D+bEXNMox2Y3ItDJd1peYH9qxT0/4AjzKPc2pGyE7XKcmpCP1SaRcDODKnl08PlE7Io3mY3Ibipt
DJdcm4TvjJvoKCjQvLwYw8u10qfVsFIbVjJEBHFNvU+umconmIEGYM6EbJfqwfy/8r72UOYEf1ny
8CKRSPp5KX8ypesntOuD2SXaf6obUtCezgYgDpSbPmLXqvwn/yITVjSoJ1/YVl+D9WzrisM79eN+
7tXDRGa4pRG1CSej+/gLxjLoSJj+qeL+CGZYnGG3klLo4DkL54KYqUty0ZSzkx4EJXhAWGy6MNwU
55Q+MIS1TyRSvTc0HlLt80+wK/2ul3Jbu9LTgtcFcklV/L9LCNxbFh4LshedeEFhJi74mldnoCID
C4DS4qdtSDWzWGwMmvRTPydldqvqLM53nImqeD0/SQr/Zi+vqE1ZWPPftMVhUMOhd/aPzVyuQ176
A0sdMEbap7PvGA/X7PPl/ToTyf1zGeDrT5bLY5BIW0uogcr4JMvwdLOAi3Z8O6th4Ak1Y69FwoOJ
ltcdn4x5zARH3awuVePHHHK2QaCuWhSMWO8VVnXYfHHrtE+z8a++ItyyU8VZUcNaWo9Zzj4c8710
tuKrOMh/Aom3Yu1ht1qUVHvlBipNuhCrN6At9pgnLmWBErRmRZ2D6+nmqxyUO3P1VtwRaX+/31yS
i+dgohAoOMZ7l9WdEqrLAyc4sUd1/5scwn314nv7Cpa1tUZeErG19JK5YCOgrSfOHsgUD569ke+g
eNqTCwL9e7lUjsRSmrIeQpodfZYTgQKBMah1LBYW6kf8LBk/537j1dORcuRZoUteLzWEB4/qrfTX
lv9b24H+WVOmMmkcajoP0fRx3zRIW0WDRHvNhPneiI0MgMpCYA82g9aLJ1Q7KE7UJlJyi5dv5Vnu
14CRzJvTEzwVYko6VopOXn3i77VI7a7lurE7veiHH5Lu7H36vYE55KZmoqMLmIL+itXNC4Z9k3rP
Q6FWxkHPDnNoqteedk8afAO6RVTLUjnsp5qHx5YDrxQGCTsaWYSvyvwl8VYZpECmj10iRozAxaS2
w61+yhLHs5aPyT9MrLGq9L3pmDNbvwghy16Rnl59+FQud+DP9+qd2oqDNpsRzPIP44YaK/JpvbSZ
I/l0hGYIgt5hmD7BukQ/2HKTn3FyUVYqOCK7t1iFdzs3iUGdYgDXy0ElW236bq10H5SdgQeTNJ1v
cRopZSUkEcBg1+0Mr+Wysu7/PDW1U/M29H9eayaG0LQMjlgiKwkh8W2SGMp3H0quMl/mYCjdT5tH
WEN+7O0IcJAiBjIlERCn/ZOasPGWEgSp2fz7IqyiDnRpCCxFxW220x6g1rGKY53wrsjtt5NoLIKw
1ZdrUBy+NVYG08wqJPTiyXh03+KuFKSts8INdSJR69z2RyNXsa2QFKKMdcjXkr9r0ypluPSlDdf0
HOuSP8ZCYmU7nfccmOsYLko3Jpnx38n+M9AJ58QWTBviES/rPlnOR86g8t757cN9Ea31D6zVbMCI
dLSnSV+mb8OBmTzrxWsthmEwTIMqcT/C2GxxQs7GximW9pShy7uQMYlIocMSqug3Ptw/p7cJzvKE
l3wZ+XYk40dmwOHu7wFeNkswZaH1nQu1jmo6tyXPxrnO51DfBOCVpbmj9ySVfOpdXOWbtpwqmv+l
Iuw6Rra+PQgoRi5gbdmiJtg1VP5LNh4xnLHWoOZI3HDuxfsNtisbeIEozok7KqU2xj0oru3CiYBi
FdSL5ZvA4HPnuXOT9cvcvUGOVu7pCKXveCFcDy6DH7dfTC62wgOpn7CJr0zW/IoLgJs5dFb8SRt7
vTFhKYPi/Kf1huj7OjX64eevTeEtee64QamhWmaO+IpLT6fYJDqzlyS+WSpICopafnogeA0A9v0z
Qf6uVmrNu2cgO6rmwh2VVKrfcKaAhOr9caSVvOP6kxsqCC8iRDP5i/eSq+Ouua56/CDy3fOgdgxZ
WZHAa5iuXaf+7Vh5fZFKaFacSIG95IMuU/L+Z4ABtlOHz3yDUnrSyDtWkEFVIusEMDwD+2ebrj9t
LdqWLZRGtYAKqPsqqGWOLova5BZ5kHWOOa1g7b17vG6Dm0agqfN+N/ZvvR68+wmIDImDwLSlrbGg
yG/WnNToNafT/UU2HaZhWMdwEh9FEkKcuPvxmRGfA/9HAeq94uZZZzMDu7E1gzh4+0+Pw8FMsZ8l
QV4c79m2R8LyanP2015WDl27RxDCEBEsJeaZ14TH6flNrtR1DTyJS7ZxbK4KjhnDYg3g4Cl+4PaD
X1dZ5om2v/W3eqqdz5K5rLaOCItyBiKgYo5pNkVO4q3cRRqZNaoQJfIV8Jr9wcE362bts2+ktFYh
vOJJvpaP+dFevUqf9hfW3EU7+xv1gQJ8UkSz+dlIZ0HEXVAH6TCLQ6O18uWYIdJqN14ieSf9yCs2
lhZu2Gwo9FHMUETYByos0CHwL9Olu4s0TPJY0GxazKinngtro0Cpss6oe3spsl7aU3rZm9khGTR1
Pp0E5pDG3GK31Z0pCm/xqaMQRhUdlpiK1r4iOYyTcHMehB7FBHy3ZVkSMRYAsWdqIJVJ22GROEO8
jzu/sGj6l7T/bx4Z8EChtAd/+EEJAZKAzryADCI3ntepAJvTvtLrnnniFNp6e58UlbE3PLf/nQVT
0DRmmWHpzgE1yzeJpfDfGenr1XYVpZjgjQKjM4lBAfTOu5lKhUpASO2olDjLrC6MxOF4iW0S+3QB
XuLN+QaNrs61vamMB0uqGQ6F4PK4J5tjwEUQ4UqUr6ttGDV/OInZLGvC6NhCqHoFN2LldjZCNSNI
aQ+WYGQbWH+AzGgnrqluJ0VLYVp0SMLXqGRGNqeJPBlNLQfZPDFbUt3t8rSOVVxT5K/wXkNNV4HA
l4y8LHOnrqkWGqfI+PQnnWnbjiUrSZdEj+xXVPraIPM8xea6CKPXByV/fKMA+hwYF3BK2Lt3mSn2
0gVu7fCRuMLPTsi7TlzSaqAX6LzRnxTk0V7fnqTE8pRyFwMDXof/SUD9cWM4JNr4SyaycCpBcERe
d2S3iq5v/8U/dkn6kpFKaWekHCXlAHBdcv8BSlAKJ4OdZdqc9A7xVMWSGr3lneBtEjfhZB5wW69s
dr9p9in3+1gjOPmh0RWTW+tnJd+Yjs5AThfuBOxMuR6JuHu26vZskm09nSdqYpfoNhXXF4QqiWDD
1DIWlyBR891QmpVXh9GQS/93lRYZ1oVJe1T8+HcZvlL02HriEHBwL80QwpMj5Gmfxq1EIY1M4HyS
2+GsEZLJ017Ibwwltq+pb45JccJMOVW/NMSe0o0yiCmvEljIly7NR0YiOQK1ccdmSg38IVLH3/38
2QnE7stUZsOhYhpXXyGP8HWWjBsoX1MWcMH+1boJ8cTC9OBvusRYovRay8yT5TcwKDCnTRPiA1iv
aM8ErDs2kcaQ8tZK1PN5bscjjbAEhjb+Q3/8aA6oX5khxcqnAOhPRLQWWJzB0SlffFCfUO3g8oMH
wp1EXqxvx8QH/YSi0RFCp+zNpio6NXyfuchPZBhSTJsFX7+kpbWmabcSKHmS9hf/ifrigAlgm0aB
2zPY4yzh2WKHrFhKmdyI3GFiPs9bkmmDy3QA6B/q4kAKiW3WaRCihX0MRA/gPuTijq8mM8TV9pIJ
udWmmcro757Yd8z8Y3vhxnw5GFl7hV4zWBxLLLgnLuoSV0vMCGne3ul846y1VYBITUpZ+TKY7Yu2
EEmHl04n8f4c/wqGSJsK4cSeOqObidZk5eNZhiJroX8EaWcTeadBVNi1UQxOyDsIVhC+8ttZtNru
wyMKGFFfevEm8FHKvuErN2xOygcqGkmyhDko028ZfglxdePfh213L05FDjh3fR95XvLPALXdsZAq
+NK4m9YSOffjTOv9TorWkW0T5fID2+34zQnK0d38hFj6pS/Ye0HdbExpUFAONtf1q9d6UJM1h0+W
cLmiwERm+IdDqX4kuYku2hJdYHsDQECQdygNNj7jCVRINwyONuTorQZ3gsKZlzgf4BrL0uUbCR7y
KnyJiT8/Y1nBYscy0NycTs4AYbnZTZ/1kWhW1eb+LW7SkHv5nHrjxWe/uZOUM63nSP3bP0xVGYeO
9qxo6gGQ8D1+4/i2CZHgsxuu+5ZiQZWjgfNvxNAB1gxy/W0SfjZrqbAVr12TL8uJEJG+vqQq7LYo
TQ/EdUi9NlfszcyJ7qgdfLdqOapVsm5LIirSQWARtdkW92h2oaGuhhGvrzkcAHKR8zGVfTcaXsqQ
tlOydtq2nwK58BRDC7nvqs/9x21n7TLo4NzRxGsy6EtVNlI5hUpBt9v622ER1wJ6F4I2u6nF5PFm
bAxvnTCOGhjkL6afZSUJ1jOkj6jm9+H0EpCW86QvR85MFAqT7zsm5NN68wzOl3CkOc3hozIZ7wJd
4D5owYJGP6M2MX0aTNlsLBhmI1aOaxZ5y7k5vzy0RE8hWkKGI4sGKK8OoEDr65lyt3/dw8T8HmeD
GrGE9E5r3xPzFJ9cVa6a9k3UUCU/sv1+4aPJE3irYYArJbODfYGu/O0IlTaCGVDCfi10hvmCbW11
yYDunTMoqu37iqpAU9zglRq5HAWODIVaDR1x4u9MdbJTAqsfGHmbrDKmiMAqyktCd46AWmQa+/kk
pCwNTTPZwCUtvOrd4a6Jhw6DGQkw1QfS9AVdUHRyZIVKVoQ8zbm4MvmNvYjP+b2lPZNC5IaukFge
1F4ETA9whZc2HqoE5GKKeUeuANaaUu6tkMXgC5s13ub50jcOOVXXUt5HiRLQzkPVAnmqd+BYdh3O
1AfXwyHQjQSFLtYTI+5iueSKaxUNgMvqUEa0S+X63hXLfV7sBttwXR7E52sN8AOnC080Y+NU14/B
kJXMb+lbQTUg5yv5PCIi86+OVal2OX/7WdB99EWpdfhwa28bCxl0H+IH79k/Hd0mzLHVM0uUzF6O
TVF7c3EkPcYiYHw1ohvEAm/s1ezbh2XyrMQmMFIpsq8KYcQ7FCRdyktrgsLJaJfJ7IfndYkeMfo5
XMQgA9IeiUXH24+pTiv1O/OAVfPRf+BbU86riSZvjnBkaGS04HODYfJ/SLHjci6FjtG5KSJRIeu/
V0UgpMjIq/gEbEv3E3FBeMHJOkVFRb1esLKcP1XuEN5Iv+XZdBsBzulQ/liZat3xqAuoq0bTUHgl
smR/0dMlsgFr+GTLL932A98x0pnkSedXfXq93Yxe3zZuOtOZrj8wxVRGcCrgK3gdNJcfb+zqtLRU
tYlBwrKhR8fLjzAMETcqeczKMpqqXRzPc974Mpi6vHCe+RtxPYgH5CWtEuubpxL+fZwk6vEBC0gf
6hqqFyuNV+/c9/ekQn6qEWxd7VS0qDybE4qB1nOs2FbsEi8NiMc92cfik2GjfMbumSDtFxGvEydO
K/lcrfQD8OYNREVCf4wbrUraJzqJ4U+8lDXkQqkMOKCNC6gZh9KbEPrJh+SWt9RY9eG8yoO4LEfx
fS3YpYuC/hwJkDU/QUIkWZTKaaDK3228Y0plLwkRajPRQFq3WC1/uNayp1Bu2gBWe/x8gABhdRxh
a2SrcWbn6uxhVUI62GEPni5LLOrxeuTMYeMgo+JyINjBUAvHtfpiOWO0tbA4kUa0RgifjHylAryI
BT92+e6FTWem2gzgg4T5vopBTVetQMCVHp2T+4wzOJAdkz97QJJvBKY6bUtrGyiTqZlgmy3cAVW7
S49nu8Pv61Ef7Ef4yzvGUOkf9+eRoJ4XTAzNuTJ5ts1Jy/1nMlrgSd6MIRgBwVGf7Oi3wAyJmjkN
KYcDFr2HzS7AStA6k2Krlay6qPtCIxO/kp5LIYs3//BON5fKBOaho7RvGNMXWiLGSFPLdht8kjhy
CtCTUPiFBObOEeOgsbqz2SMdHUE/Udhuzz9OKYn6dkCInsMd0/6Ecq0Cgt+7ve3V3q1AK6mvKuB8
nkex4qGLHoByoQ5HGYZCTbwUBKbpNSXkZyFLj1mifRPvEHVTuYd/rLbcW6V+w3utejCE7Zt2FIKo
U9HajUc0Ib6hgNn2qQEA8YFSCNpGPHDhPx+MRrZsQ2DA3qdIqxes0HHglBA4hlNBOkIHezkYl7om
lw5o4+Ix5q6PaLwICLupo/L6+eAtXSNny+pQlo4RhoBbIyZXMuRjahu1Y37KT1Cvd+2z7mgU1D4R
mOr5FYTZth45Dk6pVjKRdkGaE51YdII2qNyIpfJ4i2SRTYDG9H0E/QUfbnMecbBXVELG250c0fe+
ZqLsqTyUIS4AJ5GwhPglbqeZRkGbJPbdUOJ41keU/k49BAevyTXWzfrlGik0J112kCqOXu8CjP00
prSoPJJc/3NdFCsDjjm+x3SPRI/H/ZBb5vQYPXguHcJoZHMJjqHy0CWUm4x4DGN9gFRyxY3Fh1ZQ
YIOkeoLMSN5LJLu/KmWB7nUNamcT7MLm+cEfoUWF9uP8oySAxVd/Fj7bqM91uXrYUpmy2yANScJG
+oEowvNzM2garyeK7clRR/clpcxJJT85b0k+5lejmuke9ZsQ18eNr/SkyNDTxAlzNs19sl6hPHAY
+3dlHGWBbhuKFZ1mCS/iXGFpEHnujn7xILGtM2uzPG+Tb+j0bVyzl+3pwcOuiFeViPQVycQF2wOI
vBs2hwget6GUWgTPfjkGaF0+qMr+Dz3ZdzR0Jk1PTz1qIqEJRxeYbKzy+JJk0cMO3YGhp1xTCFiV
exvU32Ouh/99AnPpI7ngvXiIRyT70gYrDUn1kjuERCfFANZBbJiPF9zC2JvE625O0/ML3/2dFcQY
0fIYNkhPXwXMoO7qZsdbQwCZ2z4ujYyGy/kDFwEj6w5NfkJrbEU+AHOI6upwtvLTw5InjauJlkcE
G0eeyJOrX6xIsz7lPu5zm29eNQ3xVkcM8Tz8SVKf6HAKsqbC5rqoPk7njZ+YStVY7rhYDOn4zgbz
hHB6ajv23Cd5f7iGksTbdIvscLtFPPjyQ5gLqMu0dj1cMAmc4ju0hdZ+0RyUZ0iAfLb0AKLUrapg
5KxvANOqWlrjB3lt/dGxzgIcOeBDjZZK+UrSIFB2vPduyjufBmSSYzNTOHoLsVGKYvtxc4gto9+q
5E81G2rQR3c8KcJbehra5Pb0TiN725Oi7zLGnPUNMp35DoojuWdK2kMpcCBTp584Ty9tHtwT+MGH
WH67MgIjNYExDWZeqre72LPk8CeWx20N0pWz/6oYm/ZJfHHygysDAzVfMdafrNVRd2AGPXbPxNck
REKQpnUmylJohFWVmECo7WIKqPzShPu3gUlX2D2rTjp8ymCtUhAw54Tcdjk/B+Rx2z9rcxj0VTWE
36ZqbeFFoLB182XLPNPe5wXPrHmfdGhXHYUbrWEBUR0EnAAHM2oDCER9N2MTFt9h1SN30UMww8z+
Tz/kcsaoTm1kKZo/dv3fLnMZN/19XvbZJSs6Xsmm1GVMXk+6AjS3/X5c2XLZBItwYPy3gnSoku2g
BX/9JE3w+ya2k6C0GTsd7sFcZaefpYswxx49uGn883mlw6jPdr9wObVR2y8XDRXvYg5Kp+eCBmLG
Lj4WMbCO14U5KLqotZAZiF76SLKwG0SFyZeE7/aVBXbnzZBzOunqkbb2+qhO4+jghpcIurAbNmb1
4/uAYlzYzmJaXOwE2KFp4lvXhkWBKPiZg6BRE1rld+bN7JhRiu+pXoYGhz1MvidBGk19WdlwITTf
xypjCSC9Z5ZP70YF3fiY2PS4E9s6FYnVbCNEahNPEbQFxtd2W45XOZfLtzfmcPEnmhg+pchQwExG
y8PvAKlySDKwIjEFXnd9rQkrhSMZ/0+LodrhinnUIJ0EV6bo4NACLDfRaVrJ1CpGZvmQjEU3y3Yd
3X6NNidg3HPzvHLJJYnZsKjiew038B1Jv5yxsrj+XWZKpVJmnyH/1plydSQsmbnwn6XC7Agw3a2g
M2hFMYaR8OMJqnUGcpmT6yAEhuGd8nc934dNbiENJFBsrvZyCUMN1MAuC+I5pHebU63O2uXIWdXC
sItIKfp2LyTc01my9yu2hpsq1ZBSGxHbBPHdX47Lp20OUTWDK807Ow5VaGszLIsWjhK/FlOdsRG+
WP9vfWFLiXbZeDIKN1Ve+JvpH7T7a1e/sFWTYdFaiUjpSxA81q5G7BvXBRqqEWnbEgH7kXIBvdp+
uhwV9nBCvDhBRIhtaMv35gtdU91R5a/G3K/bYXCNeDLgLWSDlE5537Dn9zTOfup1ywbuKGyeOrhb
g1lc+fZMANmdsbFrmcWHpK63o8oCN0iIPwQFe3m9+cJjEawSOVjcIl8Qd8OI4at9+uCYClsJbxr+
+NxRa3k48XN2EFzxysse+i218tLls/ElrMa4CCeIjxkHwewkvXKGKmZLMSCoEI+AzUKzOwYRnBsh
sz1RIA6KyRKauCgUSzwIPvkIWkwkrDZ7+jy8xGZsJ35eFpYmRWHvDEaJC3LbEXsAQ08rPdSu+cl5
JXBlmO5GzAijijAuvGpmLfilVFe90zrUh85BBo861nvfKzb7s9xTtEwHgG3GkSrfxhbLgPT5ujYh
eNJQuPBkvUyRR/h7SIgnulRrKAE5ftPYHDXtflgJTxejEQYc0R0wzHHKdS4LQfkJLFGbT6TCGuvE
7nmfYFncO2fCjY2b76TurLxBrGd/Od9zOBC2y7iiCMOr3KGGUcVbrzQxWGRlz9Rlop8yoQgC8Vjn
0HT0V31XMn296SEm71MlkAB9NV9CtvwoXo88LFJSZhMYNVxQNdh+w2w/nLTswVyYGrkvjuxSSkp3
F9ekKCUmiMS8dQE84Y9wbYIN1/RqgkD5btDX2koCxS/u/UfSTWa4LHBQvEQKYymskF6OfbdS1gi+
mn8tiKI9rEud4usLvgbYT2O/JGJWvdywBwrZh/WBUQGywdZmxhzkPsfl3KZgH1Y9a6g5OAAc4Grw
3dTInWbgf1MUUTiC4PYqftyswbVSPWciWJm9vmFh+QcvS49yfOPSq6Vz43RNS/1skk0fZn8vPHPk
WTihbLN7HEPK5JiSGrbSHnCPeQ0kztFVeRmR1QCVjuHeRUVSrRO2NSxeKJ8HJaNIR5RPfJ9JfKlM
tCNVbQw6cwUzS0ti59qf3oz1nzP9mpPFphhTiYdgCYDCVVl/Liw0hKsdeZz8BhMumE+4hlAnvLX4
gz2vypYz2swIQGlb4RyFUMrDPnMyIUOrQ9LGd5FemDVFDSXWXgMUF1WyYbpRfYQyz3KJGtYf0gXm
y8LI+UVx5cyPPd5tOlaLqvdgis3BDniCibEudojFdtxIABhRiMQj9IUFitBdoMkFmMazwWdFqise
+/f3u3BAvxCTeImFeEuLmGpq+vt3wm0odF+Hkc0C3D29107FVim+cfXhd2jjbZSInN2qSP1YzJxv
3FatbxvSReEN+iWuqbcEw33o53jZqTCHNLGd2r/k8b0BiUFWtJNwLiZz2/eQl6IDwbXEHXtJ7M42
ZJutXaROePNgrxNu61Fm/YdNCv7ydp6D3nfU/TIsMMEmdACTZaCD53LVwnuCeIA6pEELv7qhLbJl
/atSV+tLLWN6DmJjMrgR4orrgm1gzcTQfMzlCWb983oLV8Ru6ogPsyWSMqDMGbGbLcnp/rcQ4qR7
jfHy7jNoH6PgnpM0Au6CjwoSyk6AV+WJAXAYIav0CTZERLC4drdiiSCsVgssDXeW/ZxsLCBfFiHV
zI/2PXHcVAnz5uDAiYZ9RcTL2pkia5ANGe6oF+rBbgtNKmhJcCdDXms4SEBpQ59OLmfCYRZji0qW
LsGFgs0gkWJlt6WkcW2XCoU3B0Nd0Ox48RcJsRewk4gu0Xn6+/uVgWO1BftaIeHD5yivalgvKw4W
Oc+dliPyDV6O3QPsq/gHQ8o5hyY0EUpbdc/vWTcAB12uol/1mmnSNCsSNemUBOdj2+YWtl4wCmlk
Hg4f7VP2Bhiv/4PRnWI213SOxOpgc0SWIdFZ3Uwuy49vgFMKYY7q4pwhh0PWcDKUDThYwIJOKPer
GWCqRPguOkJyvAODyiA1s0oTyT3LB0rfom6klZ/9YlNk1hZhnsyzWEWo17EyGMABNidOfkfcvFwF
nhCCwoGj39v14CD5x9ozto30JiXosAvZ/3CQSg3qQB77HqsBxGE29NWdUXI01PwOBegcjYMjb2wW
Gokn05RaVrShyZRrYl/02peHdsPDSXruJjkJdGrOxJGjRQg8q+/Nz+VOLH4wYRsXE54SOVLMF/lr
+xbMIEzB3DcDSqRFJRBe93vDV5I2WtsauFQB3TCqCntSvcBFizHYMmQbqE3UAtjCZY+cXi8X506u
2/DbtSPv7BRkjOu8c0rspVM38bfdI+9/EmHEDQBuHU9sl//eKiPp2Sf8KDV/44hEUFIyZDrS4zq5
tkjbZo0rGPP4ieN977mgSS68P4F5324kcTvxuXZ2Rw/w/G+GGnyYgEaFWzl7IJUiOmqRf2ELSTLG
DvTk7OD76G/IP+kmfZH+yehfEQnp2X0kKrXQ72sXKN0DeoTtFn5wcS9Ow9L6LIGs3ypX+kX5Bh+g
GFzexfMChxg+yj0semJK9cYeqhLWjLKJ1zaCHp4VNg1NRWhYx10qiZtyV7FbqV6ec3GlZP1iIuwV
CLBpXgVVN7zJZG55/iN8w5Fi/oW3DJ2jRAVaGaRIz5/e1N2fy0aKycU1cjURusuEKX0t3l6mZ+Pi
NmF4SSMkWPjvwzBu69gG1Rm8zCNP35iOuRxlpWy5TAVcjYuRrN02plB6SI7DQKnXFpFl0GmXpepL
VmhVX9mNptjcr0kWM8bRnY7pYju5u0ybTY8G7roLvbUHQMUY23oGLkNjpbKj4T4VPfArmeDxAf2O
FFCvNC4aRNihb0MrcFpvPFEFRugXcIR43Igmx4GB7MErYi2MEXSA9KGt0OXQrLW2GWV4qgFUx9Yo
J0TwjGyUCgTz6VdcQfIB6N7+nT0EhxphRxBi7jJRpUA5MjByg1cyylIMfWmmEY3Qs0GMc9VsT7B6
ayUzmW6P3POenPziBlszGW7AnqnjTU2r+3JIPYIRjarjJpiTNoROJiTSer4jhYlTd3ZoP9ZnQT4l
5Yhqgnyu2RwY0Kd82PSpRZpHu9kKnc8LIHsUk3Ns/u2aWf5pTWpEhGvBhVnYz4R4pPmyo7kBxSI1
W60+ywmFTnAFnzGzuXzwheeu3+Y4hGb2fAQMXSFcNzZ0jQQVko1oKEXyvA6lt4QhWYRiLe/j/pwz
4KizY7TTgChEpHaVzKGhYTQ09JuEYIbD8wMyRRdbG5NVCzUS85wwpoheTj5EU4rNc6h42QdF7rO6
kA/AEo+ObiM7CbFagkTS0Eo4JUP5cIxGH5H4vrkE2oxlOtJkKyPuOjIp65iKP0l9d/g0IcybkKjS
5xP5jupRHc+W4UzaiWCD/Z4lgoHTCoZqqV3/jXMmEGTqpG1e9/dC3lKP1IC9o3KV/Qi7h1ClnZQ7
pGvikH4nfMoeiE6FPpZkaHNM0K2BxCQruVLkPlnQ4weCYW3js4Q38IXkBFwdBgkSVjLd/puRMrmb
WYj5XlX5euvHO+NWTpm1qb/JkXsOJ1FlNl0sg0Ii/mn246AQ13prpl9b5SKZL9AOE0VDAYojRs6I
zr9Lpe7QJgZyWagwsVCVptRBye2u4dLyTljiXy7sPxYnG3P5G0nu7XkOqr3ywqSRaCTJsDzUeQbC
mOZA2mdEvdeOSCF6q6HTOJXUf/QKgQCvYyZKczti7Nxp/hFVEOCYgdBk6Wfk+N8Iaq4KCAaeoS3w
gT2UptP+N1Fud0PNyyIb0PeI75KVcFh5SY7M1xsOXVkvNbTlo9tYNxPsvqEKHDENUWXPyXj1P+q2
5B+eoyyXX16IaFZyc+qrbaUCkD99z4yeTny1370/V/FrzqYsGuW9mgGtf7dlrEbas5xW9jl7uz98
6X+TjjPxW54lfkzDSx3GsLc+IikRN+J9jp1q+Qg7GA+PFBW2WJ9ShH+kZ7IN+76VakEK+Wv1c0ah
6ljyyQYqGnZfVPeV1tWBOdxWVMbhYmgpGPxTPqSIWKbqx7H6RWpQx8bPteFU57d4MjpFeTZ4t4oh
sOKrPxS5Qeb/ltzdQanEPRNmmPmKzF0H+JUUYT/gD4Xc9VcvEdklxx8GSax7aZ/o3HJ5wCcIFNTN
c5pAt9aLSJoaYwJmlkGK0HEjWf2r9swY4kIXmcozosyfsFTOyK8/BA0Tm9yhEmNy+QSY9zdahWs8
s8vCDz36a0pvxFCPRTeY4VV8Q5Hjf3wUQas8dkMNcwZ7tuawYuKyQSn71szoqHyWDnIIsl6yrMfH
hX8N4qwVKov8JqNy9MqtpzCgg7vcOnNZG+1mvjopctaFRGxhZjWbd4/jRpQEc7EcPE0boav5kz1n
8Wwch/rWl7qAHdoVR3T8u8480TE2niUNsFwdYvIdl+DMQo5Sfzl34LrRfeuyxARdEFAMDV4Ow41w
9aAHLtEP4FooTygaAzcDayGOSUxyf8gY+HTjtvh+SGr5uO7xXc5fWDsVrtsYJF4tU/t8QJX1tR9x
YougUEJnrxaSKourTNn5sfhj/sIrxuqARnaF5Kczs1frpAoUFpPKQhrVt0LtzwmKGwMdzJXqCLtd
pRzcO9oJ3OzK3KmvYUuA8wCaTVKo/hysvysMtLKAz9fQDAAWnk3b0dO7wgZMouPthCYhZAf0JEwI
A3H+gjVX2QIDqNELuH1iBpB+EPDABfxm9wgYWgbHtD3VJu5o+UKUdBQw9KZCoeo3UvxavZwHMf0H
dush7x7vZ+kFr1++YWUS0As+ehSk2gVpQZoGi3Je/K7Q+L7/d39M9f97G6YFMfQE5ADbryE4Rd2T
vqOvHqYzrzgmIzwjScUG5+ZhTeNnfuwuRV5jqfpc1FqJwn8yrSSAe6w8kIwk2PMiqeQaCnBW4Xkj
VMQ6p9w0eLFJ0NObFO78F2WzEXeVsfvRh0tYzOldNSb/EwKQJS8S6+F9a/WIHXW7t7Ltf1oqIDzW
hhZITSuQy4I+tkUbpd7jDjwRMsbaetr9YcNrgEpxvO4esBdbji7gc60nu30soyXGIlmb8ibUM7Tq
sp2DaI8SYR6FZ0QyMS6WaFJaaNI8rwHdaQUdUvQVsfdOMU7t1F0hRxmF3rum+IIxg0D4y4zeI9ga
83U0zutAXeHE/GL+TPuLIlG1CIZSj+vRd5iuupohldNYz4At8DW+hECEwRaQKIC2gErAzTj6zmQt
P1p/iyu0YrH/nneRoMQxHuQXe0ioLWewpIi+8G/RNhPxZ0wmuBDIwJt+8/CWF1VEvxBLO2cBBWlz
NIbZhBvo2JKfh1s7u57KpGoPWhx8eiigUudv3f56Td55eKhhIHxehfgq/gyUF97I3haPoeP3eL8d
pA8UD03XLBwkwidPcynTTLCG+N0sVQetw1fJPaFp0/QmNjc3k5G+7SjzAePCAvkX2e+3ytK3jM+j
6PrEvBbEL+shnKJdgk5U/bwZu/wKIWtxJKMWmMFuKIslqwKxPz8Y0I7fzH+dft2KG+etrrFnDC7+
Gxeq6b+32PY2DrgBKOZ4jncTZ3DEImtpkjCckXzZ6ikROaoJekw8bu/POSZJ+BSuueHbOwYcNqwC
9tc8lVJf/54qG/rKDRQPMvPubzqwiJslp59zaepU4W690U+ar9McpF+0FH/pcGiUt2chBqj7jMaF
wMC/XkPw7Isfp6tOD68RkZHM63cYD61BkAvCx/vDrl+xeQXXijVD5wsF9DacHy5zuHgo70dNmziu
PYv0UOyZVZgkV/3sie/J+QXFNrKdpLbGSK/DCnRW24UWjsGoER54CCdbmJvZy1fTNjjKgqfOh+Wv
nGxxdD9B4fgEDKMaL22qPh3eXCGahYTBbe3wVdCT76Rz0gk8h3si9N1SrDW4FPS28UdJYTEkECLA
jwOcldmL01zbuptYK55Oam9fA9c8Xn8h33c2lzhyu5sWbbSq+AMp/j2H9gZebfNDxLSRDWTUt2uV
U0y5CfYvjA85E3P3SI39ooqK2dM7FJZWnd0v0EhoHCisqU2OmioRFp+uei+PNeVTM2X+zvXKAc/b
OBOuOkLMo/LM+wcpMZEP1OLuheAnhyshGr+A+vwb5ZUnmKlZLsqANr5LqiorAKr8DCa2Ko7GwKlj
viqCvcrtf0f9SgmU4JgxXsOdkezuJusIgZnsbXBSTRklpTQhWf19hSigoeBu7Lr2HcVuv/Q+ZYMU
kO51YqpEAq3OafXrJEaF5iia/L/gVGti31xmA9Dqu8f2hyGzdNRjJFoXW3mysZSs/1irW6mvxCmb
3So6zKniUVHGbnBfENCiiJg2WTVhdTxFGYkBBTL4Zk2oEgR65Xs7IsRu2mL678EPE3I/N7zSXyeb
3MWGslvdrLRnziQ4UkQ6xoHizW7gn0OMprCujQjbrbKqR45+kLcDF074vNi3a/92sTwMEb/6XStg
vn7xCVE974CTjSMttBhPUAiwC0tiQpvPbzR9YuJvXrFGnwG8/t1pZNCpYoVhADnPjw/VTluzrzXF
eNC1k9sa2sYVm/jvAxGkJh+up65mkLUBWXU0xBnY/9Ylo74ShAjXN/c29+sqescs9w7Kp8O2czjO
7v7z/fCI5V/09/o3aBdqJmJBnIEtWaVqrYEW/qwNa/oFtMNuWDky4qr12uE+wrZm2pi1gvj51g55
cAGpRzUq3sZ+dqT+c1C/XC+N51sJJhRCyTwe/UBHCefps1Fg93uHA1ifEHtigf6aW8C1Uv56WQeE
es3mL2M54tSFGipqXPsKkdqQiDncVezf6mKDXhFA4Ze2n/HPwowiXGktwPSHXiyNOq1A40/6EIIM
5CAwOaDQMpfhhHlqiRDQwviSJXEzwYkhpgL2l3OPxWsqb5+361SLS0i4+6WT+3PRzY9XHEKAPrzL
Jq9YijN1OocN8zre3V62aE6ZYsneWXMu3MkdPcrBX7EeIa/aXBhprhMIfMeNzEjCuYiUhP7/Ek+9
Z6PJzRH5sXOOW4OlPqrLM4tfIxUqXubvuFfTP4qWOuvUIvlvEz/spzNDF6d7zri8ZJpt5lBduCAR
A2KrGxIOf4AePRC29/nBNVULvhevgL7DXJPL06ncu5iwmfuQDKoCCinfxWtwo72WuVovpS1CBA1D
Ar1AS3XdlPg++89286S7SCgUbWsXSNnRKK2HJa0OxaxtYLPqA/SxnfQkis8n30Eji/cHRD0Td8hJ
Z6uEQxN7y4r7IuMwrmIvTNqpCRMnkIpHxAmlGmvlCuOI24tubOAo1gPPGaYSl7EO2Bj/knuB/lWu
fkd2kaY8EL+8mlFg45a/zL7ah+upAb+1zTK0H5dkstd3HV445Sb5Y1o9b4smLYeVipJFPnK8+Ycf
Bmz+FIyIFTcMizSyaBX7TfN8tzmq9bJRKgb1+MHtH0XgeBqUzVNhAtZRuvzwnkVAGdjtsler9fML
3b0vSemWyW1mAxqk15UBvIV0ej0eMJe6eXD3x7dSHqxwGv9cdYs8i5b21ls0Zsmw/0/tAe48b6Gl
yDlGnXHzzEPASDZU5Q+lI6hrrEXewpGfNYnUKDqJ8IsRcE11U610eaUtdyYfRuyh18a1qowTn5Zf
ionof/INLbVJrGb6kN3h2SXNKQ02fJl8tmLu580+xu28ikWwmv/C/bJqeQYuuSgEoo0Tq93rvKxZ
CSGcMwIFnwS1DnwVHegHiMQR+KhykXmniNzbVGl9XX+DEwLjJY1QuiCdERnq8AIYHty6Kmjl+S6Z
0PWgT0SE3GrzAbSX1zaoeak93HDsPV2ktcEgamoRcmljtGaN4dBUa/1ygr6Ug3Al45/x461obSU/
k2TkeK8N5NwHaQBoNijrVKuVrYSTJrl5SutHJZyKvMpikdzX0evPNyR+COcQMNfQ4xLFU1RM7Vbk
UBR8MXyW1837eRiTAqC3tVgZshOhxGxxwsxFDI6CbThUnbRHUsoqbiSOKkok2h/iR7ySYYbqL3lC
TVr7UpzTmFnqqZubNYkRV6XmmiVsTu7jMhESE1nZzqezZcx0mOLnfFfdceBpbfAVN0eavBxYNPnf
Cx31DX+wxTc5N7XyxtN0Jr80asOQ0/m97u88/ryZryFHzWOCSoNnSOocHT6O+M8O31Cge/nnJsdt
ttAHhUyH03GF03CiGkpkOD5Y/KluDHOgkWI2BkoKhr279+Pytww33C2jURluluTAmWqJr/kZQZaz
RFhdMslEZzEhdLOfOix8V7+C7r9Jc7GXvTvoNSTjSdQIsXyBWRA2dw0tU8IEBRqKTqXI6oBbIFaA
7S/TfztUeud/9MmoQFFY5avMLO1tSRmkAWBFa69DCtj6QFaMIhGyLhLkzl0vFL3W4304P9ktE4FJ
Pak0I5fkgZViedQi96k5jpS+H6Z7G0ftq439R0tb8h4tRvvuDYb+lg/pafb8SFh8oD27h2mfufau
jJvqGDWbG2ekq8DRjCNb2F9ajJJEOe89eUAaJXtgtPeexbDjCr+7clYPrVKt0egrl+3Qy/Wr4Hw5
A5RSzD2KnaGj/6XJcs30LV/7am/W7HUHSUWW+2U+wDv/0ngcBAxYyY+z/+p6rSj5EoMTXO7TulyD
lDboSayUfbhN5XbSjZ7HtSJRNTdXf+6x4qj/OPQV2QFwCJVc6uZQr8CQNM5fWeD3Mg+K4YE8eVC1
IISXYh0OrEHS8wyJysWPFdHaUz0QAm8BMrWqc61EWTE7yNoua+se5ja6tcvOdC/PfONxKtvRppHx
p9vmJdGGmMR7u4UsfN9sFrz1MuUGejmjHikw5wZFpVCyFSABrzyiUIL/4r/gDOiOFAjIBiegidOF
Xn42KO2yU7OhfjVIdQ4GQNsgB+LATNT9MQHU6NV8FbyEsCBrLRgkZKoz6OGnhBWDqSE2R7IZrG4o
KracZ3uHmDcIteMUdubmmk19nN3njXqSBQH0luVjW5wmlQscD2MIqSp2UbGRau6AaOcpWPrPep9V
CSuoA7+SknQS4GimFm6BhgBI2mVQGKNl9riqhRDhWOaSEikLc4j1AZeZwSmM6ECIzvUKlbvwhmpZ
W1IEAVurB9+kwtU4tLL0jFby5fI6KQ7SuBHcLo886DnsmwG4XsDQmyu0JSxAVEXcx9ZISoXyCp/1
zDPn2Gnfi5Wv6IAwCUFGhz7uVfTexolDx09GXiuc0d3fFIlVwCatDCwH6dXu2YuIe7HZszQvXgay
RFsPPPg98l4TEsplnrlJTnHRfapDUFF46LJ9m8gHvU1iM8ZdTCGFUoLzY2kYB3V84EM73Oq5bbvl
BU4xbtahYmc0LV3PJWfMEqNraGr+rnAf1/x8BTX+mY3BQ1wJ5ygsm7eBHPFbXNp7rfCLMD709Kfv
E4YW0zZmZo9+LedBk2czBlgkJz7I8To7aYLluoCYiL0zskKxQESXTewRWc9vg+1BxRMbZ8O0Eb1I
6YGkw7s+dWWA8Kdf9RWlaAaDinqZbcMZYQhqT5Zadnj/wivU5mM3TDX1abtezpnieuPzZhHhk+Vq
Oe1yLQCibOyj0CvQ0xYJaF7Olh/NLFnUEuTtMz0mSNctx8rr15mVFi3F8U6srV/NrQfoe5vjVlnQ
M4oEftC7/8MSm83F0YwvitGexXRlk97qM+IA7cHHC6XyACZufoWoQLGlG7VHiWhzEK9UAUojtPKy
tZRT4Em7vntr1zFb/aILBIWb8a4LG4PQSZ39F53Gz4nxC2EVzXo51PV5WC9x8waHC6jlgL4zn0PP
INs5Nz5pqwOtVstKSZbFTUhUvKKF9b3uz9AXQY2GvVyXdT1X11GfCtitFnIWAzyonDhog09Ah8Yz
UvN/mKwgKxuQvwbGZrDx04Xm5kifckN+gVJzdS1G2M775qXBhFEtEqhqk0GvcU0aWVZT++3i/vVr
DcvDfRd+Kwpw5vJoXQ9AcDWjTOhghZR83gmsDlFK/BfIcbAxeSVA8FGcw3txdiQmHXA3iZ/PBcCc
F/Bj/E0RTDxHbKUTrf/9uQFNVuoErnfOIZJGevkeH9ZWpp0Q9BQsj0TDmz/MSq/jYDl/aL7pqlPm
dHQp2P7DVPOJl8VZAHqcVH4fh/I38vLTuCtvXz+Abj1GmFscqpiS5bkbQRzi7gHXziB6IuXRkY3H
a5Q1vYsSiYiXHZEPpTKXjbC+3mt7imu6+gxRcHdULZ7DGbhBsZVLBJa1kV83tKpIWpynwenSRkPS
Ik3ZEsOH9npDsUO/LqQZoDHt0OO3opPNa6g04vQuIKM1QUjif8Md5Dz/YY/DtTcjnWmtboCGzGfD
cbCyfEXKM4Aaxj98t+E29ewJllSZ5Tmn89fZkpyOhwRDWb5mZUvgGsMszjFCKALT2sRTJD/TjMus
hk/LK8UKDLwAXq+kAGbjG0aheiuLGgnUJ6M5ZKTx4X8dqt7rZ9mNgPiimKWEaTQx7lhtNBMhaVCW
H7bIqokLF+HQNDgYjZGpxjwdTGKdd8QeeJheACdjNsXq4fjRpErDs9DRJxdKtPa27n3Vn0JrL37x
/AhdN3hS2C5VXhrzLTfAiDVTmFehKX1xp/ZuAg6+36X4SHKnv3UflFpW95/A/fDhpwqrWA8Wn+1V
U3pf2w9Wth+V0qW1lqKkMxL8p/YwXssYxAwejD8PEpuZGMQjwiG28MY00cO2eUy+sP/kPUpSqxbD
dmTKYbJCLpt7gpaCu0yaAl3z3VYAKb5SagdPPFOEY+DmEVy5X9mriIXbpQlCvp+bFN07JmuhbnZ+
bNX22AXwCPRt1eJ99XvwJ8Gi0ZGejG+uQfhqM1rftN1Zc+s6HX9WGqNULSzcHWaH548tsLiYKpbd
RTJXWVh4MhSn96q3vf08ypyvKj4RY0JWYTyGT0VCFXYDvMK9dnIBQWai2ZxrsRVRZq/TbWa+qVvd
iLOzcA69qVnLW4PCOEbdUiwtNtE6IM3hj/URuok1USH2TtPzYJhdj9OdlGQNByalgRrkptNNBKbh
Czqn4rrE50LfQlvg1t7PQt0AT8MCOtGY9/imbVv8gXT8y49/LHvqPsuOu2Eymww3aC0JEJwoEex9
KYzW41ZrntX4a+JOLtnPXTkNA5P4LymiT+KVQblf5n/iaP1XrvZmB4WpO7yg3i9HjFLF5BnIT+m9
9ZIob+2DOzgDBJe1tPbID+RrSuPWfF+jXKRkrfmF4I/Z3v9edIVuRLIEg+dhX2rVD/S/uD2SZsTT
QgRyxWFdq+cRLsmOr5QnTOvl4ZosDT3U/3nx2A3yUIAMpLszkbo3CxoVIkThnqs2zZ2n+lW2uzSN
MthegWlnKcnML3KN2yrVo+F7UxrB1KMagDnPv3t5DG9ug69iDHBLER0vlRho2XkcD3CMy1aafMqR
Zmn48T7MfJhmP3Kx04qlkrHLVXta8q3HvbPBDWJkDC+Q7xxF6kk7YEA3zVEfvQHyAzYB1EHwXmgy
jpFxYxvGM0UKtmhTwnI3RBAulnQAsM8XmbcBMYh6qhGsXGasIQgG+OevY9gEfuvFqOqB1j3S2krG
TzF9HnUSBuFli60uhl9PRfjVaXFB+FGcqEl18kXCGO4nueghZ1UUEOQpsYLpAb2BtW+InZ7p3X8Y
Y+oz3lXIig3lP6lMzgTgbxExn+ZSlGv2+k365ZGesxTVjko8PxRQJQFyi82Vq8HvVP4h8A0bl4ag
zuVYt115FWjoG8JlNKaguA1a6Diii886iIIbbe0RThojVg86MsMLOKthC4RLnrVk8jHdIrPF0D2D
27M6bTmB5wH3svxUpBCeUzANz0quUKbNJ+osQMgGaqQSRXTZWNQcLyw9iPPqv9p1HeDWQJ3cOBLA
F/Tu996x4sH3JKXIR8JFEBfvlXBbqT5YUpfeZvYSWy7Q6LFwfF8DvjCV2daUi0ntJPy69pBd53EE
X52PK7hi4UpXueEAY3gB9agiewOoeNqPUGEdclmkdK1cW7vFuU8+iAnctqOFWsP1fShr4NdJiuPB
vdt3+z7lMzNB9pIWdbz0e8ckG2BdbsttNr+WRUJpXRcpEXrl/2rgmsAwf0o+RePg5AERC4iNgNae
vCbCXKjo+3sszVVq/yYoIRG0B07KXyGT5QOpuNs2GTzpwZMCUwb7sP3x1qfxl6r3oVJiBgy/bgE2
6N//nBLDHyH4mOst7PMFFJYXC0Q/+qjDCfXfcanamQe4KYHjPHof/K3lX2X0zwfxiYSDbJhnWzvg
EOV7VrKVGF5xDJ5Aq65fjcIpuThZw9H0hiF2pDrLT4AKZRgQKm/QCZxz2EqBaBGeOYIjaCxBvEP3
u0aj/5upev1urMV4TYprQRa+d4rK/IyDvr3o/9uXekr2Ul5TVLtNwHzKX3NDUovqRUsnlGnlIt7p
AoSmWAfFvR/C6sRpLCK3gE0sXP4YpTNij24wdvi1gcp3x+XUn8bgUrR5E9c48BYyYVXxNehJo6Uw
KVsTFkdQ40CIe4R5w0xtWCQLYpms1uT4+r0qa5b8VjiPio8YhcfmSwEaaQtWoGBASdwl4aZZFq+g
J/P05ZrhxMVQShQjLRd9+4vyHyKqFEpTwPr16BUSWRxFVlgF69Zy37JKm2GLxRl8is99GFdShonv
/r7zKE92PsIBGFyxwAWBOzM6S2rIe9qeREZng40dgrALVyRzkNcCPeaJqhoDZjn+KIs5KHaEb2Fs
K4iu4AktmU34hO0EM+SoAeuEpXggz1WqtfOmxD+vvdNeGhjoURqUUTD8fgBM2pGXZq5A/z2CiMdO
Z59Svp7OYrB1PBokkIbAOYUZq4bBjevA4WxuVz4h2G+1bA+huuJP70w4Rr8QJcEP/GSK5ZEH4oHR
5+354KKaTkwUoEbcpNAafWbzED2BXrLBnBiP5YVAEM5dpV3E1F3aArR3tl7xT/EF7SdNcQgLKAI8
XhZMIa2bWXND29BDY6k4ZEHoyiHUA/u94elAuFPjuvzE423xunV+H+YxRz9BMbj4DWZrlgSObkpM
1MpnCMVrimROcea4oFv5jRWprrEtW8MeX91zxrMcZoR9KPKPuUN8gBqRvrIy6sLjVbbNnvGZV5Gu
ZvVGptbivDmX7/s/PF7aUtk6b5M5DB545yh0KM2hWCuefcUTcnt9Y+Etu+6ngM8h232QEekmH+qj
d98hOR3kDKPdPp3OTYUgrkAGg88vaX6pUpN74GE1gCF0gIWdxUng/5a9ba75dUPVrE9D9g1VQksq
cqgAxX2u3PzGgkum1ZsR4SKzKd4MAlLI5yJvP8+OrymySAEG1NUZ2MloBmeEIDuM0nrCPSegjsac
zBfbSrPJ+hS9Il1DK2R0rk+zW6AB9hxJ6SyTYomMtIRNQ4bAOlfaLZQ6fWoHNqGxw3im1fV3QcfF
8zuiq0TFxHlcVDAS/UXDZ2Dmahj23aktPBRXlhWn5iYTnqa46UdQtX5KUZDRXzXDL4EEip2ofTrS
B/3EtB9jXGcMo8bMBtnvmBQv8goypy01M69KXwo18t+NaO2KmheNmn+fOcLiEqvL5OQomqZWFTUc
PVpcfFBjf1YY5h7pfMjyn77IpVDfuf19lcLPoiprXlcYpTpkZ7HA/iK5ltOXaQhonphMeHOmSpYQ
RcHmWVDrRcxPZraYFqBlJ8qenBbaxNaJzK/+SzRYCuC2aSjsae57/7+Ee7tj1lrtVgK+8y3bMYsD
A/2GLQCASVNrKoJT2sB0s3N8+Re/eoMxXBn7Mh7StEH00Pt85+qVLRGA05CXjGVrHFPj54WdpFde
l1ZqbOnryQG3gbXS0/qYor5ejokLW+YeMTJNufcMrx/PW67VE3YmtA5KFC//UkrkbUAHfr8fLnZX
goSPx1zew2Qs0XRjZBNWuWSFpkgvpAOP40Co7XeAvOOEPWU1nbh1d92fG1jOAwk3N0qk73v4M+1b
nBpWvBQKCH0RN0K/rM0nZcha+v3bfARqYR8u+ulWZ5w9Rc5N2qkmXvo00x01stNrWKgOBNpPRjEq
hsrcJw4wZbH2+Mc1q9iR3GdLFCQJBFtbMI7brRnJf2/E/lCec9hZlHPgIRVW6AaZqP3P5rPaIPSz
+k4Nbht0rpGBfe30LAR4GSwjFsklxkwRCOEYgBOtD6JrIdRgUAoq9oDbEdxsUBe4cnWP/NyqE54x
2LGyu11qah80fIQaxVmOJvlz93th5cyGpY4FZ9J5rRpSC0U8Zal88zduG1rLe5E1WBJ630MzhPYG
af0stkZG+EHiQQLeXm1vFUUjfhMEI/l8Y412p/uzuCOtK6mHj0WdTaCcBKF9WviwQOOZF7FZKwFr
fZ+rjiqTth6i2+bW53B886sqzeFz1dSVofESCnTL9P6llwzN7a0X+MhMCrGWGCFi4+H691PnK61A
LsnCzKyf9mc0q2Qusewei0ZKmErvkxnO9sGgojWat1Bg2o85Ba7XN/zMjtb9A+nKqoZqrYAZisoK
z9Db1gKIKaMIwrcD3Ak+2e7wi4Xgjzm5g20LoAUvFBLXIiPt9xCwWEAhnJ5uc3naTja5iCMxAEmf
vJ+5IIDuR0HSQxJxzrnqx0UpN6MTxOitBE4oEsa128dK2eRyASIQz7nY6kNfmFk+89lMTYlEWjWm
L2J8ppQuqG7lo5ipbMeap8rUgAmQBuUeXRYLGTPFKxN5FFvJMMCiaINNrj4G5UTw1jXH+Umcgr6w
0nXB3XhuYMiseoni6DThoCgKhG6LU+DQZ8oZPtJ12cTjikvqMN81KVkYG6ZdcffuiJsBpERy8wZA
0ZQujNbu/4etqWpHaARVIodSKYZFn3/rToyHqkhUB6vb6F89opaz0LCJIeYKwYCVbH08skoF6VeL
Gz0c/7q2gq1Z+TYqw9SqRD2Cs0SCy01oqM5g550kQ0khXnchVKOvG9C743syvNpe8J94qACmQNDF
q1yof8LEByWJ+yl1jcUGKdBebOZx84rnH/+z7jQlK/uNmMVPYLP68r1MPv5DTV7ur36c4RNUVTVI
T62k1B1QNRuFWu9tWJ0LIGnOZT3BB+eNNRnMeUWkGYFth6H1m75RsFW1LxcOuqb2nOL3Qh3VppwJ
+RpUSHs2DFDEm8Pm6KCGIufxwxe7pTik1toJ4tquir/gHd0IM5cJSzuwMI2Vq9/QITUEnCgrj4O1
Tzqsum0HtA6iacZCJHe8wuoCvuE5DUHgWwT6ZHD6GavFzT0SSwypWBVuiMpl8tYz9Tia8QFdu+lW
E7J3YwuTwW9HWOAjcpP1bOWJX9I/oHcdMoIpW4xkiq8OELR84kZlIyw8E+FeAz02CEOWPCJaoM4q
+KwqLeNIpmXRQABV9nzogMX4FnSUrs805Uh6HhPtZRmrhrzry/gnXIkSSIkwZTYx6MXS7wO8E+Wi
Sfrc8Aq3h6ouQm8ARD6xdqssf1Dc5ShQGp6TizahymgsHnvvK8cldGEHPxAG/Hj7uPKTAowrpWQn
AvOjeGDHicPBWY+GW/AP7bwtErKIyNfqgorWtSafS4yue3/xsXcudL1HZpU+X2UyYd+vLPmXQKT0
7Kgx3z2bbqPtm3RWFVHMJTAENP2qZpU4SNA5/6opZ4u2rQ6ntMDP4iJStS4raRsWJ76OV1vw0YyE
QdCqinSdjMNBBKqVlZO4OJRMYwZ+algRLeOWjUJV6fq0c7ejHBTU4IPpcBhHp9pzeS3OskpggtLH
a/PRtaFcXQJ7rvdEIhRCIUf6BuKV9z2IGI8NIPo6RycubfFf8OYdLOu3oL1OMaZYWAdhn8vOKtgh
WnqW4N0ZMFiFdYGaMo14kMWd42rGx/OD5Mtd5FUrDgO8lchOBb3cQ30nPmwBYIxxTykYa/5sEx+l
TxaE1mo60XaGDXfzi0Vji7Pix//mFDzVRioMD2703zWgl30/ztN1J3HMrO52x0viTZjRJErG1tRo
/x/usKq4wcCutBJD9Ko3i7+o60yc2lCdtnzGnzJE5D3WQqpN4j74dggy4cdtIw+SB4bkTlTXNlbf
+Fqw2uzu9OPE0+8uG7ki2uF/8gKeC9A1xh22OP4bdGuqaei214n/7lne37ng8i2pPo0lL2aGa3fS
Z/m0ejzsOw6DC2AOIpmaEAJJLNcF9muXcyKVB/iczWWpAmiz7JsnK4OfMvTwqweG0mZoujWd96ZV
iqWQj/HBTLa966Nj9okthAQ1fDFpF10OFEzCb/a6MaJwo5QPYrDGqlQjVUg1o/XefnGhykeAXrGy
vXpTrIBg6z0rtVVbOlxnRKCnmPDLM4MUkZqgIzwFr/0iVxztLA0AXxlBNtU13TkhWmA2qG3VFE74
qes418mp5olTULetxWDnOHCKDurPdRNDIAaDR5oIFbPCy480TNnvbj/pKQwllggpiJav8x/hCJeW
4JdY1SydY0KDQbNbySKTeYw527I4gm4aQSdcL09j+jNZCjssGPRu4or6fpZUZq+TrWYwZ/eSGE7s
eAioU7TZlTZqNnGVDPs4bFWgWosDjEf/y3j4Fm+GwxqaGkwpfc1DRSUfruSaCyujsPbqDLjxJyB2
1p42rLWy1Os4nW2KeD6ysUCu0g8Y057CrLpSEEIRr7eb4hj/WI4UVwGGwJQ/1CA/q2dRqeEaumdl
WH5mgLFA8HcPLH8KUd4F3A2SraQqTQbKDAT0ktDzOz4hwGitWL/9Yu9UDp2sExI56ST0b0/5D6FX
XaOobKAp+k8vbgN5ijuOOYCiylhkzEvFDKi9I2T26XJYRt6dU/zzYGPMEbmdWwjJyOQnELLYqHj8
i86rNSJfr9DEh2G6jQBelLk2CoC6tRffc02mqVWT7pYPlhSG7SbTd0BYoME1MJQaNJapZaXJ/I4n
2EfCeXoAgOKn/1cFbQ0zWMtcDUx0lsDWv4fjUMaIQuG9v1QVjYapcoRPt90NiVkiGNlaawiOqUpI
YXEJsg6g033rXMIeZH7e9EZ0SIezuZv/6w2qLXILGMhA0K0ykVT/6QaBowZC2jYh9i4MEPa/JxFV
YCLl09e2MAarGDTw+C0ekjkePg1JVVFDKqLZFfhDpzz3Hr4GKXkFRFqLuEcqdizAHzKXFF2g7HdD
W7+MkRvKCbr8e10JvDWkYXosUIYATRjZ91vi+AxgRPrwvT8zIXjQUjTZy+xVTWALYSS0/sL2xgv2
h78mxnOBcYvy/yFdQ0KybyNlaLOM8CfZkDZ6jTYTgj08N0EigzQfXa/JZj63IyeafdtZNbOKMSUV
KBhIp6Am+K+7MWKNlYzIQOGKd2fNsU/bkrUtwu4dixDA6Pg3jI6yu+tr7SkHhiScAWjGgfM4uo5p
G6haiIP65wW1P8xZjhuAUC5/w2GfVx7nYZhXH+R9SGoXrELuzBsFQAe/5uSmiV+Mfs+5UW8ZlUKv
f6k9jfBARFAjnnBwxAC/+XNp8rKo6y3AasKTgWyVGr76r+Sr8FJHUTe8Gyu7k0boF7saMUNc7uWr
icuZTYyxpI+q7bcsrMpVUXWUjDPZRVvsMCNq12Aq7/IsaUAdzNob5FMDJFRRQ+FHR4NYItmY95mr
nfWMoVvztkBuAfic8Oyy/edNBp3o1tnHqObw6w+753lOwEbNbLWbjkcV145oBBgonsvh1sJ4pGIJ
DBocmKEjlH8+8xKhvve6NKXjRWAC9LM1stfK6nPIaX09+2AR5/Y+DQguHGb+d+vx8jNuCZaDgyKJ
DwnaL8P9cr+Nq98vVrxss08cAE8U9iZFAa5wp8p+Zkzwx5PLcBXxekpTXbw4BumGEyeNderzF5Ik
hYbCco3brQi/tmCJsYBDhYvsLOr8eS5saHrR0FJTZ+nCBQZLzEPmACUhXA6V9C0Jc2P8hlB6uka6
moq2rR64uOdd06jZWB22Xs2iSQBg0wDX9sQajNNGKrLjLlxHOHB6ef4HgreS09zKL6XrBK2ilZ2j
/gznllAE09IL9M4AS+cF/c7nOG70Bwdk4Xbs0jjJbzuJFvT6fJLu5mDTXblQy1ekgH5392/qUvuJ
P8qghIYXab5rJcz/MZw1scGFHkYOXoneXkc5iJUFqGifB0gRfQ4bRf8rPcH3LtUWFy24jUzsdjr8
dTNKlKbyKEa5J90PrN+Zt46qdlAZqQTBcDiHp/AqQaaicjwVA/W/LmNGdIHhg+jxFq+RdhzrGaVW
O93aHZud5sOOnVo1vjWT2nGr10b+krKoMefrtV2qf+pZUwr/SVvDN3WRCXsD4ItIjiE7R6+HpBbf
jM/Eu0Hac+H2Zh/myX0Qpjj/OqPi3l/dT+SQE0qo4Vx7/G32c96feCO16Y2/CsTIC+v6bHX4r7qg
swofh3fMG9eDhQIXd3ypHiHdZBk6xgd2dr5N9RjX/H7+I0JAQiezhvcI5IBgkwnMdgSA3R08E+pU
SNrKJu/uoMjuvN5S+3rmxnbjFg4NErCuGJc/Ng1aSbxB7MRtsNbumWaf2RyA5UBcUeaN2O/u2yIc
JSeiera4xZrY9JTD9B2k6II1AilK79x3+VotdsYh9MdgMTgjLrcHh7f6AfBdfEWChE5kmUanSep2
WXOis1VyUio7pB+MfP6Vae1fbQ/It0GbbTPHWeIq1tPM2qdDMuKI6em7QirKxjj6PwQm9P1tBSq2
E0E0ZB/oVrI8XvGCLOBFEVF7c1wdrgj/Oije4smN7qpqaPgsyXCEjOFtq+FKKaTgW/ITj+SXXUI0
lHncmy4uI33vXSYFeiVtKkUsn2kTW+njbzFs0k4jzucTh3gUpHrFeoXs8APuYic8feW5FTATEK7M
puKwKPa5NLWhL/NSahf78VIhgfH7tVfZ3h64NoDRh7r6/VdLP0Itkcb8k7NCLQSGsgsGRAWeQudb
10TAWVyieQASvUA8U1Vc/FqaHTy2hpVVa7HJGOIeRagPIfyB9RrTQw9Lmnqnv7PoaZOFFfJ3w329
rDgrxNZnC7gJI+8zs+13pgnRxGYHaD3lrcJo5/k45CS26UHpuDPSyvvxnfxLtkuOOL+Q7iSjqGrb
SNIntW9WofrITjcEJxPn8D4kGnhJTABd8BQKBDltlBlMGGW4bZWAw2ZyaS7IIMN2ttTwo6pMQ4br
mT97mD71rfNZrbdhxlk3fXX8iXSrdBbgyAw5QXtA9t1Y4O+gB5dXeLloXeDR5KG4XPkfhxawAaZk
i51uBTtVsgSMr3Z5ejdhVabZF5ky2ElTJXyct/rmberbZwKUN9bmtgcCzoPSKPOuX6WdcntSFw1k
8oaE/rHuASxZNE9ICMuPr5rWM3CXjdDOLdN3xm3fmZ0u08yv0MgwlIKDJ88WABVFBfFxQjLgGjUz
0yIFfs+RlUYYAwrQx6jkO3xmIZQ7fhvdsD48rHzpUBsJMAW2UijWun77Pfe7MoE6GEDpf5GuCE5B
Q259Bm7JBzeALXhkQVpameyXNoY5KYqT0ImjJ6paapDOxeI3YHdBbayy9Yc4+kfe5UEFQ/OcwtRe
+Prg8PslKEJtAgO88g3Lsf2KZUdJJTM+X3ZHtJ9ynFqKXt3wxMeYgXiutVT5DXHuExYs23QTmlnI
dkMqa4znpgmQ459/tv7xto/xQXQmatFxNaomfQKE0xcE7ZamsVWGn5pfP198/HxwvKUcipfpirMx
o/oqN6VyK7crPW5EtwK9p8vplkb2rpdDnEnuuKqp6b2r8/evKVGmNodzaHmBgTvfLkFmkiQjjRFj
Mp/i7vdR9hmR3cH1GDONhEMQMHs30ZT5z1HrDgOf9D0x6USHH0vL1KCKzIzGX4CJGLo2H38A1CGa
v20nWqyu+QBlaQ3vjGaIMD6Cabu5K25UNsHpztCKZ75n2kSxqb5rU1mWEmPcTN24n7s0nBlM1uFt
ddfHfj/omDrykBsp8oYnVCJmQfMe8BjIbZoI2FpmqPXOLm2wTKnDwr3OvPM4lAmKZOS2ApirTz7A
59Sv6Inx9AyiGLK/dh6BCo6myyjJEnS8ibwozRQRaOz0sIXI/B7qBqz1btQ7rgCOa0ofmNU/lh73
Q4hJVQ5cqjlgerraP9o68b0BR/IFhZ9niDYrcu8hv7PX6R4dpzYWRzYfLeO/2JJt0h7a1rsVKwNU
wcGPSwSCR7MemsE60YPOqXeuuxVtRKG/IArKiHZSdQ3d3TVasuuqut40vdJimfpO/tFPFjahOl3Z
SoPG+eOLpKR4Q7hE6AhB9fwywuD9pUfHLslXjrJ7dr+LM3jddfqsMsRnpbrsCgcHAfZtIyXVhBSQ
XLwN74XD/E3m42celHHH4QuSAENtrw7XhsbTCXUceEPRz7vybmHIZSY0AGMDzQalVA9UHQGcqzFY
VB8DvBsMUqBIlOTkRSiGiy62i4xP/JkVWLIl4FES0ICxAbKTsnMr8/DfVywHfjIgZZKiSMNuL6oB
GvOb3uNEOxFkydUDkBFWfav5n8GltRaaqKa/e6rG0tQ/mNuvfh8ObOCJ+nhQQP2GgRGzrxZHtBgw
uj4PGlRAMU65261AhU5KjVZIC6SG3VzcpoidIY+I+mphuOoCdE4G8ICRg9RHolxGixlQUOaiOyP+
10c2lyX7sxIoeV3qN44CjwuT4pq+WiK5aWSnEE7H5ly8Qa+TTBDmgEX3CFfchZDLDS9ljLHKVdTY
vL7wrvGZUO43AfW+y4cSUfBzglGVolcHpyF0p2VO+JBm4R75Qc+KaOBLcIHV6bR8yJdufu8FAR2i
AhPRuZPBtXPcQvvEGc99Gzsfvk3rBkLa67uixtjMZO1MIchcaFP0ZrazFV/xKE3OCxsfl06PsfN7
DkYpytYJzbatUViS0tQYc/jlyyURESK9flUFB76nKztvpdGWYC7pudmHl+xEx/xBWYAygb3URvZN
6b2HsafFQiY07408XTmUXLKc18GbpdFInzZ7yJVhs7+qNrUlrgsQGtbG7gA57jAadv5Rl+4rnmbt
LxqajkGJq9A8tnHoSmN8+EQYz0TXt1OkDFGODlUGfPROqtydpJHBaMhKjAaVKEh8PJkphMFsO7tA
2mSnVJNC9sMhMvxJqW7WLgez1VmmCFTiI2B94CkurlbI1to1kfAwNqwT9Rv9fLuxNiy5VmkwawG0
oL5m5MUG9rahaCl2bsvBy8GWDJkVf3qtme62E6P+mmYnJxBZ92OiDgUuQFTPWdN1Gbu5b2JR5xci
xK2pYNVjupyLfv180IXaFuLNHpayYeOqMYCrsfCzh3l4y934ECDUmFwhEAKfOmJ7/RrRXcfiW8/L
xkV0jIYCY55emINzqkICXHBuxtqA4nJQKn+kIFSII1yv2SqtyNcVC7m43As/+icCKViz/egH7NWj
CciGn09A/lLEHTaNqzJjFcWb7f5d7nwARYfU1LdD5c/FxWhFXDpQzf5coEEpmIr7gPcgj5lixbmC
2+QpJjvKDpTmdbmLAXVNj8houu4Uw2g+y1HFJlI8q1A2oMQdw6MEN6Q+CefVe5I7PpufbZ8M3CpO
C5V8Qo4WCKvNnYOFuX+OLS7Mzc+cZOge9FAy0AxZqlgQ/z+BwRLHTcIJqI40kdE69it2knnEdFoW
ZK+lrAX/aAbI4WZ4tAXn5R+xK9a5ogiJIfVlksjViE+QalaP8ruDuv2SdJf+eaFrKCj8Tlp41F8i
y9zAOV/LmpXwSb+iyd/nZzI6V8Q8t4raaTMDHpLTfMpGG+vA7CtLUDBL+xq1akrWo2t/hiYyIt+J
7hFnX/szVAXnIzGMtHgR8oHx0jV4dwEfLKYQFM1U+AiqkybJgWvi59lsHqlpuvmNY3Z4G8rkbe/8
n6WR1g0qd6fw6en+JoMaJKhIhgbwJ7UzSYQC0A0NcF0Z/qt1gWOye1r2wGqdMNuCg/kVEOJaJisv
55Q8uTuBWRGMVTKWBaERSvBuPEWkBkzNalLtmRuPAPrjeZVK+iW9O32h3b3ROkvsJlgRUW487JRw
yk67WUkMaVgYhv9qHdpjxsPpDyQHnWb9UTGFkDfI9Ztb8DZEjTegk/QM0zvDzxYLG6u9g63d9/R4
ormqD7eYLFHa+RO3zkaltWdoWI/P9Tv32k8YUJDLwW2XkSXPCklg+FiyIfF9dv5AMdCxNtzFQJd8
Lki6F5oVoTb7IIxYUZuToK4AEvsd3VW2YscLBhCDXkkHGRihyodVygqhM+IQn7jWNRp1RLxctgWf
GUtjJ5SnNpH0ntWBLz2jFp+LT7XHJQQXasLo1VYpXiSyg2Lp06/VOjqMNyRbKk7H7H46sUaN9/kp
zk9tfyANCcjE3tqen+Jc5pG0anpYLsrxJ7qRANvLyA2FyDEaVUwlifnp5X1pzo4Secd6YxDVl9ce
uHDFbAhiq+DC9P/WLoczzBLCcXSIAuHqNqiThAXau7mtd+B7blpDtfbdUfpHwBv4Kr8hVbWO6t2M
4O7w8kSqJzPO+xgl0w6BVrzXff1ATpOBLZUADsjE5/6KHu48LpRfAr5X27kb/78epn60jGs7qv59
KYMr+bh00Ora52qHrQNNTyw+LXr6NgZsCejUdz2XQRw8FylT0YqtjipgYQ5GvOO+2xU6XwDSawZf
5z1Zxd/UqEgWeIwmRv2us8m/u5IicZa8REHTrgo8C8zW8f4wWbTAE9gpU5Eyev7HhJqrg1PZUGUn
Nm2HX8IRSyfTYYWA+IA/wG65GdfSuRSFxhkFSE4fgES4xLqBL37RtblCBuFFZjoBV3jj5nQ/MabR
0JmJo6RlRcVLOmUrcKKvhQecpTR2qLxfe6+l233DYsd1dUDPg1nxmCfQL2ImkYN6O8ROFt6+eeUC
xtT3YkaqVrQAPJhO2fsOEq52RddbWZk0u7HjS6s7P+mkUgrjW7xF4RPUWzKEK5arXWIH+MaZiSZ/
kAIgdXRSRZGnR1V0UJPl1FiH75xenijLvfsUzTESn/L2XrrSN5iXbJXPxVDoFcbnOc2pU33QV0X1
KCixyC4hCS9IuGBBI0JXqHWUKZIoRv/RX6XcgOQNpb8Y4pEIcp/Oqto6leHc1wiqVT8TCcwDC00U
sv5zG3Yo+f7YlRn2VTL78QfCOYTe6/iNyGR7yu2tfPPNU5EbZaMxf/+J4tMFFmLA5gk0b05ZqRxS
lNZaHW1Q+XjD7VSxvZxoZO7CI8wkr+jv57/00FapgYqSm+Pfbth22Sdf/R+iJcZ2pmrKLSvblXid
PhckFBdb8Rw/LfSsetaLtO4kjNHVggR6ikQrnXc5i7CDh2Yud1a8VA1TUUDDiCVTdSDOOhACAfOU
kYZW76mBHady8KWWpFKEPpa4WkbhABZ+wPojjvpSsMQKJxVPrzvzxPUu07n5MBGiTl1b9jMw0cf6
fszCxU0w0bJ0jMJCZMnxED9fMHgfV811LWp2M9E+xJ7E0AUEskPrkHK2F+T4m3t5xNb2Z9KEWLJO
Y9Y8tq+DzXuRW8rmtTYR5d1eWdR71R2knKi6dVV1l5ndMnowx1m1N6Olm+tMyQqQKSW/wgLLq1QE
avsrvRMyu/pJrvlxXNJ4uc8xOnQ/YfSVFSKNgXzUsFqHBcpG9pyW+wlSbsf8SlNmcAGAAD2nhZ+m
qeqw6ORoaDK2+kaIzbCUH0U7iB50c7pPAS1KOdW3YOsH7wwOWRWJ7RvsCWC/bU/AJRULWt6+PdiU
f10mAD7sXLLYM6Z1YHm+KG9pnIv5jKixb2BHCSZ4eCyzireWgoNJYzZS88DE3Ni4C639aRlT7MSH
BWniMImwXEy5WuQkYFykgP3Gh/8tH5pfujMIhChEWk1Gw47FLP+L0XDqJK82Q5ujMHCyxSBa9POu
MgUutZEBFwWvxNndiw+dYzSd6nL/NfI6Hdv9fSwRz0czOKYniuLRwXYYP1J1XbOl4F2BnnCDaKYK
MQTCtwF9HOF2pTsck48K/IydqVOUWwXmrfKrKdwHzJGN7r2ScJtwtF/iX7BPtd0OeMSeqAKi7GRz
nN2xkoEClnDnOpvCrJ7Yv6sRMTaoKEzhYQfVD+i/U6z+QQRYF6gOCxm+sikFXjyW7vyB+yxFJ9W1
NpLMdNdhowPFV6ds5tq/1gWrhN5IeqHO1uzW+DUc7uj+pm/T0NOsTmd+SX0huRSxPy79T5/EdN80
/qzmwuNThtRPndnWNHYw0Jp3pqyrMna3/TXCWGBrU5b3M6APmR+rioErx/aUI9etqv+jdhZf8qUc
cVtfNmkWt4f+ONDb2M4GCIxgnNMxUakZMM4s9X0/70GEoP3YvjkUXIAATvfX6PpRwKeSduD0eTsr
11fZ9cqJ2FI1hAvX3QUFPg/ptUi5duvS/lzVSDi4BuYDD4+V1JTLvLnEUvECdQBj0bw+6wI84jZG
qosB0WbJw0eBNrUaUlgSuqYh6Jn6Wv8Qo5KICaS7Iu4W9AXL5Df5Nz2qfmfnkGJ93vHEwzLTscnB
bjUUB89ypdkDTuwV7JeyKPfmsfwyAkaGzVBHFBSqcvM5WsITmACeuHUhhKse+UkgUWksEuyd2POX
t43l8tz2pLyDodEhKuk9TMU/3ZxbVPSOVE/fs2MeF8ALs5HHy4v85fpT7OTLl14T1v7wuzom2/MB
i2HFPQky2wQY5/anyxyra3YtT6WruTF19FT45n4PMlcxvaVtHUTSXnwMx0DJm400pBEiX6kYuI7B
55jhuNMFLvAufME4LYIZcLSxwWIfT6gYrv4bOr2i/4tXyqkSGtZx+s7J9p6kqpLYFkNKmz45Qhys
vdO2zbf4jlIx8l7IhdQaZKeBJvV8Sfwt7/m+dsm3DPx5riB72Resbgu2BC60AVZQtpJGl8Jp91ph
aDE0+sKjx0ov4P6QouSHI5EJFpqPs5Z9BuH8IIfba01agtetWvlR1g4U64beEka3iOx80Tl0pA9I
8/YeJAmEQ+rWIXWTptu2K1pyktV0VkX2BIAwSA1xJA+ODBpAVjHfCcmwyQLXqwjFp+A5PCmervMZ
fHFAXNB/e661lAuA83qBq0r7VSKB+f74ZGWEkatnGFe+Fnc5SnwRhqYjdX3tM6JLc1oDAAm5XHeI
uCqbqw0OhRtDiS2flxzudAnbsxDqc44GLeC77+bhz0bLfc7rF3K5uzfVik45tRvU7t5IZ5jc14YD
T3hd75Pb4WEZ5whOmf6yMkKqSqmCTJadRJ7pWkAHeG7qfarDQrKaQ1IGBdleS9wluO8Psi+02lrm
F3lr/9AIZKFz8O2JX6eaeLcYx1XUPBHx/lZIx8+jotzZKwOEh5nU5unloV/Es4n+RM+OGteKIU1p
06tJ/OcC/D197R1UlSkGQb43cK6vsGqYmzIyyiHxrnFszZyPr7YKhu+YvayIoAjwdL6O1mhQm1En
uKES783t/ey32Z7gXoXBUSUiDPhz2wHRyWllObaqe7c4jUdus/nP+BskA4BXFFRcYEXEm0/LxEKj
QKwAfZqCK2yJuqW0Askct+lFCFckoJvrDoX/aK2RBB+3iyMdkXzc5HnVt82SxeQoWcgsZyCb1FDm
IrH330O/AnTs4J/1GCnA3/d3voB6iunpZVKVWecxE+cY+RdK/ft0RUeocMbLwIKg2bwn9ULv31Lm
lEjGO4UfTB2Inxs41WWx/Wsa3nX9gp4jNDbGgCneQcmzJWFgtBNMj9j1mVhy7d7WuhuTXLAJpAFV
ur0p9XbEZqokfdIX1i3viXLwK7ombaNvf0EX+cp3B3W11ZobjvU26XKCTvN49s9lH6N2neLjD2D5
3F97buw28hOEHjEpzx104B0p5zRGDjs0liKPqFfvDLwJ0gWGspjb+aHs3vh2/+iNmrN0/Z0Qo172
tCbYwg8+5QUbd/R9vLPRWwPsEgXH6KB+2vxPqkQN0mKok5P462a8ztS6mLfP0Fs6ttSWFLOwKKbz
H+kUPFUOSaDkPTmzi6CeXhMCmF/pykVyuwL8QFS6le0gMqb+VSk7aH1Ne62+SbEth3PkrZc1I10r
JILCZ639p61bEctUtkDY1jExwvXdtnxtPwnQlGPUmsY/+2eSvgU0MvzAG8i4dqam0CuivHlleIzi
WVP4PcrqKu1O2HTjeefmVA9ioy9MQt9kMF7+p8lzWt/ptK33DR26SPEopzcjxkffIsc09eadu5ID
Aggs7LFlEg+mBIwavvAoFBWZEtiVSICCVg4JXYVgec241SpLXS6CnPYy9aKvfvX0e670rZQXJ8vy
OfbGjBX68iPTc7XfcH1lYJdKjIiBIUP7fu3Ih+VqszlLh3UmjwZUuJ5e89xUWAvYv1u0JVwVw/2b
SE6DNnuYjRgbktF5D26JZ6GKQB0MRDW0ia8jR407Bxus8mxaNPsnnjHQD4NIgWa7Wv/CSXyZ4kDP
doXqSmgV8+43RjYfcdJ5KOxDr3zcLw1ikw6YummTNMhBZkZCaFhPVjkzrVKRIP6ct+jmcTV7SOXX
xDWMzI4cfoPM/p3bi88XiH/nJiZr7U4YMOqbRXO2JHLJ0oGfVd7BFw1p0bMUYLMcwyn88hacajGj
NyV9Xgj//RBWU7q+XFFrVJnphg/lr5BnsxaPJ06wvhBogotjyxOWasBujiEng+kLG735RBG1thep
m+WFeICy75lyuWuS63y7evHzNJUxS7eZV48g4AB7ZguGEPMF8gwKLHqxDNQHDmfv5xzl6+GF94r2
p4uKHm/ZLm8+3SIORa7OFOVb2cbj1950qoOEQQ5ZLvmOWyVgmzEF6NrfKJbbtPpUKwg/yjxaWF6m
Wk/W816hhB4hcDHGdMBN4QPxnps8T/dIuA4FEKthvPAR3EeUILgg8g9GGXSfurZldniWky1wWL1U
M+MIym5mnAx0QnNo0dwSNqv/VmwHKadUCt13YFv2aIcrm6cdhSQLWe3Y9drFRmf7gJzyTbnyv2zi
T6PPcHc3qxNox/or6fbOEug7WFBOn5YWY/IMa7uB4BW658YCmlFvyq6RWhMc8rfU3w/aOeycZRo9
CN1Q/XSomOye7ieluNaw2do6jq72Ww7qRw0yZVj8J5j4nlQIrn2QU3eAtMADykD0sxaSkz7/rtxh
bg+OHczR4R2sLE7eQBBpDzUleUzhvKweXM+x6cAjZphfELS+dBT07mISkuGp3MlR4PepqWZUwZW0
217fXVWvyg8kLefzxH+tjXmxzDsepTdVOQE7TMdhAuWUiTHsCVBrSlO9WE2sVd+JRqnsEtnMldul
VsZ1jfM2hMhXdXfqGQZwsEpsxbVpKpWNCGxOUJcHldGpNi7XBh3TOt7IMroadWOuQD0N5XMd6FUQ
UGFpK/hxbs3jGVmwwd2VODhoc03euzjQuDO5sTg37DFsZeE7GtPySA4WbTYfdutpqTkbcT66W1GI
uJENajxwsEcpDu7I6yJu3ZJsyT3pRS2Z2brEvLYQ57aoGQxvxig2gXBvUU8kOhiTUurSTeyN5UtE
m0bu1EBKpRoiRLzJpnjiJXZTd3M0iZfCIx/JbRNWwd/E3PR2MLDV3lOuO/76VAU50ULZEt0ZM5td
z+KgXX2GH6Tr3Sk0SIPCOaeEMvcwkl96jEUQYbc1tCGgqjUR3sAg+Nxt2rHUyF8f1KNKGjNaJJoI
PhsGvbEQ4bPh6LqV5oZUdOXZd4Q3lpjkfKSoJCGxdmhEo2DF3Oev6Ypua9o3bVnNDXsd8IkbnYPZ
Qof+a2KeT7c9/IPv9VA96IUnfGjU8kKKwyTGCNs3YDwu0fXlu54MfO+C4VTuuAbvCMRei42vuQ+P
sJFMHZXwt6ffOzrZE9ltHZl1plxmsz84WaUC33msKZIpBvjQUR7OhYBJ4pUURKJzPLC3k0A8p2wV
I+t16sDLjZ26mTsw1xmXBt9+246zQVTCxuUJg0NY9XylGsKzdbM1MTBXKurUHogHmvc/pLP9jXyU
MDJl862QkqHz3ngLIzfADWBYk7eV2tSfchGYWkdiyJx/oqZ+yGcnqqRobjXKX4knK2T57G5q6sh1
pRVHU/fhJ2uENoqd7RQANXOcolpbZljDaygceZ/y8l2f0euG5u7vCtFtVktJtUw2B8ggKFTwhCc/
dR/U4BA0Tk57YmZiSyexbssFLVLiIirVJqmOvnVi3uqETPrJPUxG+G4QmqNM4QkVwlBD4RX2FwBn
JgFDh2z2CiLh45mzig3BH8u+M+/tJWSC+DBliaK63r6jTuvksxlnIKrUvpaZs11AmIcn8diwwPbT
RXKxfa3TW281xafZskRQKch5Q486x5eg6pJW/nSIi+uepEVe7p+96JbsJQsm2bGrniOw5stAiRcn
1Thki2tiJawM1tvzIyNBewPOmRB6nRJCtQDPRwrlWHteqgx72BTDV+vE2V1stvfYlHxl7MRA2s6p
MtOkByd8gwvKod+17yHb3JqBvVvaq22zLlqS1tuyTRuMnh+3Qk6Qz5Xmc6tEEPLXv9mFmxdenod7
BWWXE3hJsCmfrvAMS+0/e/HSj9SnZ9sF3JX4ru0KSkjWKICyERqYk8N9i1iBbf6xqqcyqbz3/6dN
O0BCQ5uOMh6Qr9O5cAEhvyHVi3BKHZnnSWO8I1+RXETEWTg3aJHgQGwxaopAz17bSSb0cJ12oV0w
NbAWsBypxEOoOHBFbOVo+eJi+PhfOmk6LxUnVoEpds3x7+ElnQpeCNUeRpfSxBBEWJ6f6mgqpmJM
ZtKV7YaCEHd5xSEGtTN9/Fr+VRG74B7bLCR6/pe1hPEgEdP9D/7JPpliqbg8ZdhB3XQyY9e0aWnE
xhlZwYtzjwUI7tZ6eCGafc1YSqN7FCwDC5sRI5zLvIf06bfcbUS/2UzCABIeAF/+bPaqcSjAC/fx
QTbkwtY+cuKSQhQZ1bE2PHD6x/NLUxgLsSE+4YuSp/FW/53zlaMvEJQzIZga0Kz9ZLxEQgbGr0V9
zZtjkoeJIu8c8ap8Rx8bb2GIQrdK2TiXWzdPMvhO6wLjsnapOSHxkzgL9yyOF9+AYDX+L61OoocT
qEeyW7FF2iiiL73LuNQ7vH47/MI9EhMDajpomzqq9TY6myXToc0XmxYJm4MNtf7xC9i0zhflXPhU
CxjDS+PbIe41USex6gvu+dvhiG2yqA6zI4VCyr3EBVWQUbUImUCCMaEf9RAHzoGpURg2ljqUxikC
5gHe+KnoCYDS8XygstGDdC1GkcNZ+nFyr/D5zcQLFml0QIdFurScXB0v5NmEeIt/mH/OdgqQIV/3
dDIppGL1sziQS6XEe8A7M95q7QRff8cd8QsG3FASvcAGhQWQ9NpiZnM62cC0pk+ys1O6WriqLksj
YXQM+VGJdIRhGM5TtAEfJUWL1xEGrtN/N7OPS4L6IqDbIkiogPIeUYf0dS1VbWp5odgvc5G/P715
MI9V4PxgEaWJUwtApPyI/3UlVti12Bz2TjiD6VP578zyZ+BfFQIa1GGh5ibARtRUsCPMRP/sNy/M
bTkC5Q6yANIb6mxdazJKP8cirNXiJUSEUOfDmcby8WvwWekA5SGSBXrpXQCbJKGS2NqfNnhniaKz
9uP52I9PBADl8occx4hwPVatp7LMDldLxxlYu459utnzaq5x5dhhypEl7RNT5bi1lRmsfmdRgl0M
tQCpRLY/VeeX706CehnloL0pcy/pAFO4KJjBCzkMgvhGZOsxoV1jXqbtkmsN+LL4uHZVzX96+WNL
QMzSie9dKeXCJN3utUdJFipRIW/u4it3qlAUJfdH58Lb2z1JvIS7OUDv3JlBdCS/MolB4oa+dss8
bLsjprp+7PgtIdhxYFq7N/rT4spceAdKZszyYQTPSgrtOiIckXrWAUwAKaw0edjbsyTAqPGzefbe
Li0OtHKsOgHyItFDpMvbLXDplLVe/0nXxdqQbo6UuyQ6nF5z1KjwDJBGcoqIg9+dchK3+vLmOt/n
kOBsXuBJWSIYL9bpjNa+vRFPvnJRqJ7enGanwHjbo6LnJTbgHWtA4JgEykUKS/h2T71dEel6AwmM
8HDHeZLGZfCSDLM4szXOcVnHAFqpNfX/Mpd/8wNNUtcsJFOUYglNQ15ipkGXWGRAz1FdGCWB1Gtx
dZ3xutu9o7jnlzM+FbBVo8WknrC0Uwpe6ks0RKvDPire8Bat9mer5FMiCrqNhJ2HktuvN3xdTHbm
Ea7A13bsgcaxYQVcL/GzYsSgLRV1c3QRFKRJYECwZ9zd6Ou7JlvgpYtP1W8HgK2B1InWnYt9EJUP
cAwIW61vipN3v85CC215TnO0VPqVbxmpPbFP+pmjGTnYe2x8GV9MVwFmmcLrXbDXKupF6Oor2V7l
mnmuhoet75BlxUTN2SaF+jptuC5ohwG3jXfQwCksFQJ1iRTmpDwyrmFV21YmQwYdFXVWEK2LyiK2
u0iuHLoSbTnfFL7e7E7cemsWTcx8cdErjjxqbQGK25u8cfKqHYit4gHo0MGaugWgzPw0YAi5MgH9
MNPvinMo5h0/qsUzzomvNGJHju0BWmgkvS6cNTFpFH6zMVSlnoOaoLs08YJ9ntcew0wRbPq0MHvz
cTzSFSm+8AcRF+b9EP14l9sS0q5X+VcLS1p3eo/d9pVbmX21ekgcmGuz16CGP91wifFDgYl73zI5
FRQcbxkb7RV635mg9TnWBVK+82vKvMzcw5Q78phobfkhkMPznw9VLXKlQM75QadoDojy8uG2kn4r
JqH8LqFtfnVNt669kZNWUJJCn/gYLNwlSNOqOlDqwVC5orryKAqC2t0S5jrEGFtdTzj89jII/l4U
6iGacDpYAkrzpLV6Md5klKeLqZxMOL2F07n9dRDc/ShCdsWC54CjXvTI+Gje9J7n40j6Uu7rtwxM
3rC4pJZE5Yzt1aywGovDy05+ftQOMyZbbxBwEBM4caDyKe567TlWt7sxAcnkYEJRiNqRwKsHQto4
5m+r3X6TQWINgbZGbiNWiq0AgkwU7X/VTEluoEdh93wjLfCQq/8VOh0UMbldDGu9Zkn5zYu8MlDD
OR9eXt8ojmSzPd15mNDKyVZ4dKnEQzlzMgiJ0R+OwZLxokPj+frOZAiykBgvn3leR35dhsDDwxP5
8uRQ7iJPIx0MLugLIqjQ+mF1drZmopECHdcjciWcTIS52arC+Dpd+CUmthSxsD4Ao1bG0ZjrjrZ+
EvEodyVaBC3t/glFsDCedDmEqGenSh92obmxKdDgDB6HYuTUJ7JRGgKofRE5ECtQ+D2DDJSb8uLD
DgohYEfYEh9luykQL4e3JL0XU98eZve+1G/HvsHoeG2jB0DJnGrYzE9wvhidiMhrSaiOUooq9CND
w7CU1w/sY81eRxiulkBDqrESgtjTeUKCp2EaLYnsrn4N0ddymZoWJZliIUdLsMJw4VzXxvPr8WF7
gpgFzXM2xBW0MgVV00FDi6zJzamxX2C+3ldufKbh91Wa7EK0wJa0YcQ/QIUt0lqtEjeNhkgvNbT2
Eb12HA4u2SEX1oJ/sAzDzxXl+SmSJS4hGsuQMOh3ANgE3OGui3I7x8Q+AXsqoPOqvpEKHyjfutdQ
2Dhs3qVoOOYWrQlQoDPd+cxB/T9oDYPrTTxWmtjHYSxiz1690RXxaLvXP1r1piN4o7zDzXr8hSFb
ZxJA/JEsnmewDp8hZz1miJi7JlRYHjuoodq6YfVYa17awImrxfORnJ6FZn6GIAMmpQMBiZA8tJ1p
5rMGutXxttTWbnsW5ZxSz160oTnf2oi08jOMt/fhCmWvUgs6eRaOCMQzt+gcnU+zrgl0+dZJBrhy
xQmnLyCZEh0ILXv1+oN+2WOU/wUVFrYHSkJdmb9yhunetQl44lizMKyBP9vyhDKW/bAyzTDhH1ct
f3IuVU5gcxwuL07UARyTIFWzD9UtDsqYNJZDYrU9WWcm4GpKpc+8KxKT8CVDYf99DzP6vWGeDNEb
uuteRE0Jw4NepTJgg8ggmEL9zjEcBM7BBHfPZg7ozXrbVhYOrgQX+QMb6kQ1XJ1AU9sW/KNm+ogK
9V5D7b7VYS2o2Mr6SIIuoMvDatHGJMMa8S7y8B/zt5e5sUJOEXhVx5yVeG/okO+vBCxzDCIx0xj7
ZnpNN4USZv0nAvU5uKh7zt9mEyKAH0iQ1fXzMGDk/ektnZ/bfuD+3p7s4wepZhQCh+Kl8u6NnZax
nKjJCWlu2r7t9W8Yi5RAiKMf5alNHe6Px8N3cfK9LL9SW5HxKWRjcJTRLaNqU81zYExF/A6zdEX2
lZPk5rlGwSdwGsXSnDRThJzWxHJmRftwfqD5/c9XMkeGA+OdJBMfJHA9F4FvVllE9xCGo7PZIY2j
gW5FrB8558r/53JL7cChLwIzY5Vewm8SCwEByPDBsAsf9lzTwuttrLhZ432eVImTG7kqZAOtfMqa
MFAGsS7VQBiVwcdbwyIo2jqDJMbJM6hcWhyOQmveXCjanLazM2P4/jaqAJ539+Zh19UevSkwZiXQ
HP8LMKWS0lZDWv5vOE48MB3yW9Pu1TTdi+WizIMG4sk2pSQIYpScjF8Ea9/3yG3NwmULWmtaokVk
wy9hzPYiSSLRPVj/0WaQX98qcc4W+GF+/EdSHLlSiK5skBsyVt4OTbenHbBCOssBAPkeOKucf2+/
YUU2URwEEYC9nQYMtOGOMTcyH+5EbdJQb+TALycUMC+lCOhxh12FK7AwU5GkqRzdpJG7LPU1E48N
Rvv5Hh0fA5s9cKBPyBwpdc5s2rz26ObjLR5Wot9dNlPXNZ5gT46xTOBND8ukjzTW8W+HBdpA4z/t
OEueKItG7ZOttqtcacQdZMgvXErGmOCoYIHhkOWi5Ja56Xao+6TeBjPeqssuVhY7dnDhXxP3fy5U
iv8BCcLqYobG+7P91Auv90pH91AYqyTNYx1bz2E2MjWNh0MYB89gxscxFnQ/XaRF7NejIqidOt2a
JNK2mDZKuwIPMAlja6cmyvkYZPWzYoOWML6Kj50IuYk+rFmwuTGJAeZCr/jXB4sA2LhSWZp4ekOj
G7i4JGtKQ2fcMD8fePL9AZgYW5CjfboOqRLiEL5TnccuURlTw9ODTWYFOvVU8kgBAO5CrbkL0To+
P/pbasCB/84FHoNg8ZDlM2Lbpq4xYpzNVG0EVPe1pAyFRGOWu2JEJIEjamMYvEi531cGCAuD/YnZ
jwFgpElazASLdQbTZd71gL12Cf2wx+uayWrzDSWg5skhtiXHJf3ze2PuKWmfKSWDvdfkh7LOYf5R
lA9k0IPwqupc/p5MxNJnMJaOFModTWARplMOYySdDkiOHnXmz+3Q6aa6Ir4aYOZxuR6ntdtuk9ws
qhgCpVr76jpKH2k53Z9CoM9YPL6qJLZIgUM0vx04K/bJxzNHSDN2LWrB5XCXRFb23rUQZiS83Icj
8O+zzboOowvEl+QcxPN5TdOLo1WQdirsSh7tygbauYZX04DDj3NqWPwPJiVNgnxtLojJFQDD/6Vt
zdOq/AZf5RN/ThohcyynXY/s0PIFNgln+77JbgM1e2tgoakA3F//Tg8oxpTDXSyiBqBT0RqM0pbY
Oes5k+HQ95OWROQdJ6rD3ww/NQ1VkC1VFgBe3mgFJAq0BAUZEnhGY+C88nH0+hM4uzEb/pdodvnD
h8bx5NIQFso6TrEeptf+F0j4ybbesDJL03j8noHYFbdFswpALFvJKm9UkwogLrBlT+0gLOj1RpB5
ixO0zwcqQTVJOmwqLX76Ag1w0R0z8hqSRdOyUa/ZntcG3Fkyu3UcOmV1+yx+4prjJAsxFNbpKyRb
T+7MOLeXt1gxLiOZkmZR8RKXMdFUlHnTL00W/+02m5QLiDA6MwjOcF3X+riOVs1nBa7WjpXsIAic
2Myt36Vf1hmbV5B5NxZY7Ed7b3pvqFFsHI7swoVHq8g/F+8DkhCyOtf/F3hKQc2xG65do+/nwHnx
exSIpdlrQBGQB+IT4KpC4b1yHajldaTEb1DcqxfKaTohGDVk9xRAWoOvkv2+Yg6t1t3P8bdy3dev
A6MeM4V/zli1aNE+5a3d//BxpFUn76qp3Q8T0YCyS6Nj+1C6faTe2GbcHSg9zhQgtaYcJQcM0tGL
V84AIXZjbrRnIhSJaWDYjNjQUY9NIhvUn/h8idM8oqgqaLWCs1nyJv9PSsMX1fcSC2IF6lAvuXtZ
d0hDxH7tLHlYkVR/CcQtpEOa25sp9DmxsqJtEq/Er+jrggem043wCPaAr6YDMMxeKrJNTQnrQKk9
P9v1W/GSzzqpQ8KGIvM1eVm8+ZTT/nU9kD9gR/NzP/A4KhuKHff3TpUdoXbpwbbJeaQ1EE39/Z4y
sxaG1SaPu5+CUp/Rwsm5vA9JYheAH/TG1wgORQHENHtWDZaWjPbEbHTrYFUH26lBHYtnvRbAxsYA
ueZ2UQVtns1o4RzDu7z7fN/8/atR2b1sR/laIa/LbW4/KW2E3cO8GroWECmleWDpxVnv6IMEZXHR
sNDyd7hPX5aOvUpqYCZueEaaNnVnZavzU23/EMCcBxAs5Pf4CEbN+ZO4cIsX+1SyoZrLMNdNDR/I
hunt9NJcZjkO1mENLYpB4kbNPkvwdqcNDek7YXeHk6nAjd+VZzqpawcAM0Z+XbiTeTVcJf4Ac7n5
FCIjbqYz5Pva4A1TpOFXoz+6dOdRWlKkPKP1fhc10wPDfQ6uTbKEOYdlcdhQGTn/VmKh9AjGvAfD
uJTSRkeWBHYleExPsxgqQ3L0RN2kRgnyw0YfbvsRPDWgwLspYMr7ygDyYJXy9qE3k0WbG94CTddp
kAAj1BAatTHPxSDzoDDQnMwrDQhHHEM83BfdobNs9mjNTLyjCGC6LnuILGct4ygNwb0lfYbC3wOd
aSr+/54vLwY9HxVR9nApBiR42A9MJUCtTORMXWidLHWJFpzlWBGt4Kmg4H9Za6bTmy2q1uoLsO+b
DKGiW35Seu/l3adndzsmtmgO3YNsm1q6eXo63sPKkIt58/YlyB/nUBvPmEGD0SRSzsBiXDkyyuDW
ruKJ72BvnkBHr5X5CLC4PLDD7fqt3BIX23h/5u7Aj3blrWKEuSKo4TdTrRzUbdkjIeCmHxrpH1ri
mpukiNOPbkg9BfPbwEc+P8rNN8pil91bsxW6OgoFeZznFB17lG1M8D0QGHjBdb/BQc69/v/BtX4U
vv2pTcAFhM3fe4X9E0TsOuyEq4e1y5i0uScdXtMQJdY5197KNej/axASlbsjLjKTUmYgYZThYjTQ
7a+Ec8Hf2WooY99YUKERvf2GpiRu4Gk8FTzGBBzz755cuNL4DJzwQGVY0diqnTqu718OeH5fEOUC
7HmRw7TF6LUhkzUxSMSHhDN2DIYrno6Zi6H75tPyfvmF/+X11+ewi6/nWhd+ZWCL4pdItXNMbW9f
cQmcMaiPu3CdoeiRYkkgCsSi2oX7CHCoa+ggrpRdUUDMwfrsBCBLrfhFYwP2oWBA4SsiUkq4RbE4
9mOkQ5O9BwnLxcizOB+Oox8xE5Gy7lw+n6n5mLxmWmLvpp7knYjKEBWucWVcnYlDBW1tCis2CCKT
1cgXfMOuhAc21NOgIV4CNigFw7gFJ2nEiQXMhuWM+HTDD2bBwj3ZTXcNHk8WthPW90VrWXJrs5A1
U5vJkERDXAwdn6YijylAGXsDkoWjYsuKn66OVnKuuNl0hXMmUDvN0nhBoj0BCUhBQuZ9J9NKsZgT
n6gkxMUeB/c2vnNE2K2Ud4Ol6UpWfLdZAevXqOXCXLaH0ieEDcqzogJJ3U86QV1U1KRr/O15dnLA
GkkhLCcXZFq0AYt7YyxTEOnArFMp5lFzqYIYGwYhZWjYphRN/4dBNhOmP/9nB+FpNPXP8JCnZsqt
zAZYiA7qhYVCGvu4ydwE/kmUxp3aAvfhZWTOsoGAT7mLMY6H2ZlRlJb35LeNarAv8SWzkNZMX3QV
7qVcNpKi1R1W5RbrU/vAseb3oGt2QohDR48mNnlsr/1NdSAw/sYKknke8DB6V2BJb8u8kD3fttM+
qu3e8nWxkJ3d0dt5/qhJkhxSHB2RLWWQuz6lyY708BC7EjDLKOT/PMJHHq7EAEbd1urTFC7t7sXy
/Lh23L4rOqZCwDh4v7mIRRHvgmCT4fja2FUWB5e53FeaRtWzMOP9ibRYiVNcPlPx6SLa5r0qxRU4
FU0pFBQ3kU7kSq0mIjyHs+roEzRK0VEaAy6SeWDlviFntf5feciGq86MJjVUAz2iHFTPART4n9sN
4RyWYMz8JsIuZnsSAKAUW+AbcMzeTwzkeaGfWN2WivKkCMNSWw8/PBETqo0oIUpiZ0wp9+7IdBj+
Cl0jF63vaWSWEh7Bs/y4Ku5QdJ702dX6pdYfeX5Zi67fIPRRiH1YS2OTsCsdHFPGeE3Oo8zoFnQI
sh9ifTxVq5V+/TunImdjliiy4AZxPtC8Sv3m6H6DWvk5hswilw8heQayCKikFl9KpsIC+UqMwGWj
ZdrJCGm8aOIWuwGnMZjMdhTg5qy9ymvk0P5PQNEnnY0hQjD84hnWc5Gc6bU9vzrERmXfJgL6fxiW
m+MppPuE97wstJIiOzjya8NG1t4OHvQv3nNVhbO6y7yj+vuZG17aIuTfvm0YwyDgmvecvgiHjCGe
LFKXHuTWU0IEtK1D3SVZ3je69Xu6K35sRrwi97+nyBoldfP6zUX2MF0oZYTHA4CDMNz79SyYQ/Gc
QDjSrPKdTkLLJ3/HiZulEc0Ix8Mra8Jcs/ka0IOxSA0JLplj1jviq8H40p3rAAqT50kFeRwP2/sp
qGDQ9go/4dYJAejc0ek3Xe/PuHZzcBSJOujQn8Y2JTh31eyB8cOk43xmtq+6/Pz5G09NpDTNb0mU
psDPgdPLP2uMpph2NM4mcOdZ2x9KBWtvkX0XfGa3UDXWTZW4pBWtkJ25LOCUDD6qtmizT04u/7WE
6JxjNPJMGTPfQytewGckttVIG7VQYByFJb/XcukKa7NO7L5w/wv/OsNpoKr24mVkidsiwD77beu3
G7l7AMatISHoAVffbuYEHsm/MP5jkAfPeZvG96Bhj3sb95yxEDPToB776eI+JM4pqt8L8fZDHAwz
iv0iUtVWwdx9JMNcpDW8jez288gFrcdgjOpKZO2NMVI/ojNmyqgnoTg9jrp0+bY7O6aSu4iv1ZdQ
Oy2FTpr96wtx/2cfv6h+NvVdlvvqoDVHR1viSLfHxOT/6thaJrWWrqHre9/G2L8+L8ejdKprwWMJ
M/sQjhgBha6MQv8l/ZBFSsiJ/fSCUgNHHPghmElTCchYwZ+4C7xM3qwIq34H+G+lBSCcbYizHsHo
6JY2zzvPMBceS6b8Uv21fkYjfu2p2F2+NRP8tGBuR9/JLp/SFNFtHC+epuzgxrj5RZMKpHY7dGOG
IuRLh44DxpsvxjdgcixCDKNUcQqhTqkET3OlUBfZmlmwq5OVcoq4Z3lPf9PgZDQfyrgh2yi94ZJW
h+yfOPtt7wUS02sBztSUO1SNYNu/O6RgFGrdBr6W7OznKS/OovbftntiebrpO1HiVDYbmWvqzUcL
ujJq/ELNJTKzdRCzfKo3XwiZ9j8jF9eS+SBS28rZpKtKRaNcLGyY5slayfq5XuELLABC5lWHbQ4F
MgpO3+HBcpt3ahl2auzT31ZAyaMKUSCpuq6HqM690nruyANC54VE0XpySXA0AnpEHLAu8f/An2LJ
ca/xNXVWI0iVNixIaD9D+jh6qR+EPmQP3pSXPhoeVaEjU+VBk/2kHw4bW7APsId2bSlnRHMl8wgd
8y9bsEN3NoX9qbDmw+8ilqKZ4ylwAg0xIk8rf/JR3DyEQDDuPKmD+Dq2o0CRM/12Bk1tp3rOlkL6
sxX1WpJfkn4ouEm75vYUYuUr5/GHtsVjC5XI/X/hrJ2JQiQPBa9+C/DyC5qVdPzB6A4434olou4g
AuNdsSq/X0NaVM9lr6aEphSdXXfY3Ngap42qf8/cWchsQ/n3MTDInOpheefCB2Uu/wYMUBiRu592
AU5ebZ/HiKysQM8W+OYFqK/MkzaQy+3nhh15n62b9sy1MbOXJp8qmSV1CFZRzEEjvnwi25Gmg3Ka
j1PuiPjqfbgqB7DD5eM5bKmXwNckAep24Wxs4YxrZbNyiOKBhB3f1mHIcmeJHxXKbiwKsQ1+cQ/+
k1YA/51KlWxpQCHynq/pVCS/yhfIgzB1+PFvFpibUm3t71/X4JvSBvRiQlPhYZ4ZnQ8HCpO3rspl
GJbro8WruQRn/DZt/GYnDYkKv5mE6eMJGhmlkhBRRytpZdzLsW33LLznCexlN7o7aKZC9KMRm7Dx
HGrwgVE6YulznWn3GsiqkE3+cz1Wb27vZsfoxVTm59Sdg5vkhHxkUjd6d5KtrqYoYQwnkHWfXUPW
hpRohpCJ4yW7vQFh1x6/WX3U2R2wiF0RKkKyAwitVrDy/uXYFiXs9trGdtoWczT/t9CST0us9Kcf
4Wrdy1L8K7rgVeg3nfkBIDA1rS8CtIIj2QOkYnfGuLTGh42aEjsaMnxFavHJC4WjwT3DJYWlcHVu
pLys3L5Mxx8qNLvMUkk5zrJdfuyTYgaSo1TElTPQkkqNwHBMR8AqLLhMW6q2OKJ5bqq7lb9jzINB
y6UOKY9gdzKkVq7UlSGnhL/2jCJ6u06tph4uiuE60LI0+tAsc0P8bir35oJpy6CaBrv0XOapIkb+
n2HRlSc52TJVU/JOBbaYkPtqzBwPjZn5r1rgMQdW8SBbAKou/7d37rFO/EubItCNiioPM5Be93Zq
6zwlnjnVeqfuv/6m7p+a0JdLeajMujgryLn0zUwp7dO4nhlm9CKo7U0MBAtuWDX0IM8moBqtIX3s
U0N+reyMziDXX1K1X/0WoMReAbp55trjZHz9k7Sz+ZLYlxLjijDoBWLY+Pcbc7xlSbiQaIPJW8i8
IjXXfMSrCFrwo05m62nn8yBInPtb7ihScr3C6omPl6XEw0sNFhm2ptmz4sPQclNEgTFJtZyTUQm2
9gRSXp7IZSOeLHFEnfXDEYDZfIv/zJl5CPqb8jvqm6XBwMxF6p0SF00NZqMo8SpXwOhwP6vSto4y
7SQ3JB6HFzqGG+H9fhr7VYvlBLlLdEFUX8fxj5Vv1CFMVTsXEWT8HND62BJps+3nv7js6uGFb1nr
WVld/S2GZ1aUkLVLSJYJImqLUA7SpYT9PnFHZqiO83Zezn1GTFVU971+KMvt8TL7Nk5KbGsFZnrW
/crv9kCfraFuCQVon6CQ/tsFmBOPumWQMXiDtF9uU25mkR0idHPJ+mmrA6gJ4JHGPQoeSXRVkJbM
1Dwnxyff2ucHWvTdWbH49Bwh209FRCDLFIUNdTgya/gbBDp3gkAEbdUv7NHNHSll5tAtfcU8Tg4e
2TUFOz1+S0QMH6TdfsCYYzsGl7mzo19VBTMU3JAOYB9EuYvk//WSOjZWJCEVlnLvLT2ofMIyl4q5
8p9Xecd+KrAxNvNETjKLtU01ma6lFnRlOl5HIE1bQVm/mKIDn2EgMxcNTFH6AhYvdr6r9zkC7jIW
doMxn4ZsN3rqUZ65cXbcIUjmW5abSfCFeeEAJPXvtlzo/eeFGIryUkTd09U2fcmkaEY9+qLYtVjL
Zzs3gZ5J6IMqThzAwo8RPi2wkNk6CKoNeDyEZM073M21agED4TA3rpoMTKnzr5kVg6ZR02xnJbBU
Efu9z4pvf3vvPpXHycGseeCCUjfXbP9NJpiap4sP++zhmh3hLQxbJZtyYEMZSlY1R4MN3NyJCZ/P
PGLLsCunOF/khbtOuT/v18KcrDjmPEcmW4w59T8XpKdEqWqHVKQYgcQSeCTdN6NOT4Ul7d6cY4LD
kqMObUolS7TPqtdQO43gJsoKnmwpDeJpg13s5xFZUlx7zbBeHwS4uHlGQqF8ZMR3ZcW6I5/CwUzv
zWlkv1qaXbx+QN7DAwoIDTDt9Kphe73jUv4xFEJnJB7eauO0huapSFiIqeYW6FY+EfTYqFUSkoT0
B1QjxxHqwHwBbX5Ooskc8abuZxsLheQ8gTA5E/oxpXp1KRQTvDRrE96J7h5AYYwpoDF89n4L/B7U
dYpbmUpBmH6h5hJPOuyYFmMBnBI4MhmyoM65e5Kmz9dUQxknUYhs9ja1Zss3CLkSVaM03WF7wcLw
9i7HoJ9pO56IBApDxZNenuLDQr8bb6yYqJyZ7iDV7znBg1GrAP61umtudy1d81MTQALA7+9EN+YH
4c6PoLKaaswVXJbfnEVLZVW35eeT5I8cUQf93nYnWsdJMpH7JKH6hMaxPHuQ7sXs/Ky3JJ4yA7GW
5WZzDKTCafMJK59izW/DweNvmTbvldrrbNcf6tjY5agyGmtOzrumE+Bq9lCUr6ejbTKwSKPC/0f1
Vn+ZHJxAvATcJmqTI8/3U2FXDyXN9mGuaex9BdLBnpW2ig4WMLq4ctoVju78zRP+m4opUUsRFRTa
MKSyxDTN8p7j2bB6zg21pakvG+BeC9uwhZs50ySJDsCLNyzXAKVpHpp8D1QNZl8wK836fQPxq9Km
y5e8mGNdRozYopWiUqWDn2cQk+6QAPnRX4B4jBn8CqjSZFwTUQnGgGqwCM+X9UrGQHbAtcM96ctd
Xl20830ArD5CgNBby/WM0D2fBJoaqEHhCI68mBXfROCpVDiTrs44tlpm7ZkXfdpGX6Mpn+d4KLps
e8/CzAON1TW5yanl+fKmalXFOJRPsNtNgsfiBTh48KqmuM4bbK0Q/KDMYSipib3D+bSKbPivJ8bN
DnhilN+SgNdh9mq82qye7QlvEq+SjQ5lSi9T8rP5os1/Aovt7BNSRkBntA6jFreS0VSRZnIabyH/
I7ZlNr1Tsd4sFpMjmkrVlLYcEAylwwPZKMs4sKrvoB47ARcaAahYRkEY/a6lLRw43sabtq/KkknS
uVTYPeut82Yyoj1cVvLzsbYBeAgJLFUR2L8SFNfrqmFN8yKDFvREpV+KUI2Y6NZTwyxi+CWnx2q/
5xlzAGj4OJppmcUWxGwQo89tGKA5Uzye7e67EFpyYZtN8fs+oir+NubErUScP0WqaEqwkOqIXFLS
wRdOZcLYWKsMgEIivqbMvAmt0ZPHZFB4vCY4C8NrcgEwJrHBas625wZ2yp3+sdjNN0+6QL18tNrS
Ez3MEHUacANWLw46TjQ+zBf/7I4SU3jNctVPwlv6UY2+CfwYF4zrjWAmjvOqb01YxZvTfKsq6dI9
XSOrmptgEiZbp5BJr1vxhxMA+iIhxTpEA/Sq0g+s7/8ouetQA0D4ntR5BIxYk9L6d+sASLoH+435
yF1QOV9u94bcoCVjfhFpkJBspKEDayPtnE7uMBlcGPN110DarAZoYprigam8K8NpV3CxSarPGseH
mQSuZhQnQJuQaM7J6ZlQCxNC1msZ3f2bTR5KdgdLNP6qeT2FfTtq0SHInEAqnJW4GJK6ukWRPQvS
t2BAcPfGrcvw3u2zEgft3yQv6G0XXQdEq/FeDjhr3MC71V8sLKJ4H9nJVfE/uswAvOl+2+j/mi4v
JS9o3t1px51nesZJybiA67XxVaRLpSxeV1vydfiUF8velQCcdh8UY/9RsykROF7pSbpZhkJzMd4a
6WdersqTqHq+Sgu1VGMcPTzlI3NmYTnqoynQzyEwv0ovdjLft03nPMdjbG7EjtjGPLMfnxBBpVYy
m8eZ7j7OSdRyAUvOrDfioq4LZ6Ek0wdoLjVHZ9NCZLpy9fcHKQxz2dsRpoay2b0pjezoYvnkC9mV
MNsZsgyHc+dAAgRnrLwKOrbTsXmlpSkGgFu//W03vA1t13nAzTJJvuXFDUjf+RpwjLL/mQeK1L7l
zti/KJNgs7Ajj/za4eun0hq8+cLlLvac9ME9gJVt1F6ID8/u8xZCo1DafagmUwy1FzUQnfi9OSv9
UNGjBJ1nZJcwybEIWCG5lw2AnyPiSp3v3+obf1sb3IvlmkctDQl3cyigL9y3qT0aMP2RseFbjGym
GYeBQPze6rXFriAUuOZVrOr10qIWc+0P87PkltmUGspHVv5DDOV7sutpmuGlpL0qeOPv0EwEdges
4ilRZwTlecNqqJzYCddqJnwc8EcpJ02trYPSiMj+KLM9HPDWu5E027P+RFsQUXWLo5bpYBYjqdAz
HVC/nu6RSeMjJF7wBHZVfp+ZN/6fJ1q78n0EQuAch+La5O4lXJLRoWNZWf6IZXUgJ5gHfE7sb7uW
7JHYUYJM+zVbiHchgYIfaQ+GFPQI7nGrlqj5GQL3jc4VrXyCNNGr+B7VTyrwIFhmn4bzHS/rgXe2
s0LuoNMGnN6hMD44X3JcFMlkiVmKA0kTNvj+289dKHZNoHQu1Y6lhAWITpUyNyZBOYUdqF3B7gBi
Y/cH7Z+qmkj5VaQBV5WDstG4DfLGhomUyP6dittsz42aKA0LbN8v1XJ7AfqjHKjRNBaa2iw0Nixw
wrBlZb8kLrMxMeHzlOfJR2K86da0QoHyyIIU2bTo/uxK28i1M/QMGEIthQWtoSgWn7yyTpLLpRPT
5ua45jNr7yuenx84W9o5PMpRdS1uffzfcgOYK1ayMflGL//NDXkOG6NWzz8KuOkokJMx230R9jXX
5WZ/nJU3Fm+vqruLh/3yJg5WMSG1fmlt0wTO6JHKbvTLNm7uU0q40IuhBvHffdlpER4FA2ErFbOL
XVpXU9rn1VW0ZfuTnhmzlxXGG/P8Z36f+IzcOOwFog+ksslydGGHSxXZHgPp+IvLsWACep8vyqQz
dkM9cZrF4mV81MPHJsoMfu5HeB8DfHmcldEb98hxcckt9O7oB3iBv6BHGk2Hfl5Xjd7gkkoVoWZX
EycjOmRcyO+a1lbzPqF1mhBuKYa9xAJEaY79XC4ERxSPEh5Oow1NVY5rqzVEzDAGiBuElqfMIQex
9K+BtznRf16c8pt//IdbwmF8ybdz4AYbtsaAiikcHmNEeDqjFfc+razo2KI9U3hC4h6llISKRNdl
K2xtvkRhtJC486B8r9a/ogfKaekJ/ERyPuVZHikgVhpu/PsoYf3O/+R85wXuHzu3/TkamHz5BC54
jMY2wy3BPJfy7an6UriozG5zKcmBCymKGxFZBJMBNGHd0Dj+hq4OVanTYANwz4YnW9+jBSROxk4a
nxPSr8JsMkVRsrK/J8HkjyICSK20x66GQKT3mqNVRv4PxpNZtUYCmJNdacO7M+7fJ7OLPjnH/2bx
JPTSJacd8/4YDHi/iYuCIIbKmq96jRoe/0Yd59N4coa1Ml39U0WFaJ2HL1DuRz7523I6CfKSToSI
KTQ8kF70wKeCQhNoI734dybMj0GuJO0Ds90z4Hn07WE+XaNOJ2ja/7H8A+DxQm7pl+YVKSnhpXeB
rBT0kCMaFdAoVdtEhCskB+ZQILxD1HvLZlBv2rlQ0dpiYh3SRb5+8fJzyMIL29QCmHxXFgWBOecs
lB/I9Xsg4d5ijRQIP1u3vWdWcli+mc90NayYnyTF9FwzQ+In6o46YTin7kN2MK3lxM5cnUUBQ461
W9p15FaIKxjAZepMQepTQrs2lGvA37Ng4EPXob+E/O16UTG3AvYRIqVGvjuSLWCUDN4YZiDS0ou0
cidp2ea/I/LXSL/3fPiX8fUx2FFmMF0/rj4gA3J/92PMm2T3vPokR9eRva+YXgtVgUsy0W/H6/tJ
UTsnSFiVgS3oJA5rMbSYJblZKbQIv/kCTad2uBGqfFpazdVU7/l7hZxBTJOVtYolYXUaQR9N+3Oq
dp7m0GzlHyT7HivoHp6kNQwaAYC40R2aCkxwlxnvRxZLNTi8opCwrMVQKQjQnM62cxS9uhJkIMRk
EWzFBxG6lJsK2qkGBOm9xDT/3tp43b5Vx1HG0+oIDbDR68PCiGYuS3CgzH1tS/wj4IX9rilC8Hn4
wmfXHcberb1gGngOxwk4Kuiwz4r+BqFVymhhpvb/Caz0T2HbmA/UCJ8foFCbZvdMzc2hqvJyLng5
GAsOG90aDlTjgCOuyv2Xl1Gl6Eptjk5ddYQpqwD8V8TbxPThpACrfzW5olGV5LaUj9YTzxCJ677a
uiUWBYQD1gPUfMvW6Pnh3CTpu7NyWUd9V6/RzXpQtAHQJEJK1LAzYK81R19Nyt0pXsSaXPqo7qVv
zBaMzOv3xiBGwPfjVMWbyRvSmsUadvg/fMtCGr1QqUQKhdkHEoVKBCyDNtgXDnh/VtnwXsfau6aV
ESPbMkqWpUMdM+yVVKmY/s4gvx9P5SSkZAuBSKboAi4BkfxRnE+NgRJCWeR4b1ZVUWahKVwFPfPT
r2XuncpMf33ZxXUZpe0nokVBLwncjs5pe8GCeFrp8dAMi9gkoUFv82/qbC+2Yr3LoBMmsDU3Oa5N
nVBFRwnjmi3cU9PxMe0QS9KOjM++JpMpquf4uMrIwviPLhUfiFHdDEozq0L1fI4hBetkQHzcvi1F
R336oXCRN9aq/eT0BihBhNgpCIP6vpcGVIQjwbNaMOJUVdQ3XS/XP7XnPjLOKbpjWYfdH+KJ83cw
sNqeN333WKfAUWGQTF/NMG9uOXQqY7AZbjmve2ElbVBYRACVoG4ZcYCQyKR30W8aZurPi5GL49pO
CNORNIStLrjikhuHUBXfekgrLYq1gLoRuvfKGHnAI35Aky0P4U8Pq+Xl9ICz/nIA1EBe2Tqjk/l0
A3ak4s7BdgxgRfDjrCU4WtdH2bsk3Fl3F2BFVk4C/OksLmRdP5vTH4p6ALlNwvfUPAppBaOUw90Q
z5zdwYeH+dlzz5xWMQsIM08KUlArE19CSnepKnUX37SuVvbuon6g8DBYSQt6NfLO9fuW1wY8Vipk
JVcbpn3QlvTuA+1zaLmIdk7tBNUa3T99zCOsv2rc3GEumq0NrgoXJ7kV2pD3aIoMsfFKzKOhiDA7
wn/3ZV2uMxjqaBNLoJdiMBEGygADef6WwIZ7yavPTQGSYV5eTzPMJsf6tIN6UtE9OETcUXXNWABG
B/YCzl4qF0mpE9pVTK8KqQPt2wKWExkZLpaxKTvF47uARAbzfDV4SEol5On6PMlzfJJFqIOi9gip
wCnT2awws/shxAx13prSObN8z78AJHRxB5uS7d63Dj1/klKisQT1g7vnNCHaUnqK14tQXF5EcIwQ
YS6PfguFCiAeZiPR+n/SOTil4NIiWgjhdul77vDfLO9FtxPasf8anGuIYSgjGcOLLeRE/h0eXHrM
0HocWXm6z0yUiSslyhl0W/vR+PqWu5eCQjNOGGKTZ95vp+CO3PMYnXiuiK6N3hQx0SSdve4LzG8B
brl7SNaIUZxSwtW9jB2M46pjzoJ3aQThVMp5jRYpMUPkbJpnZriKpVA3qLgLGWWFW0RJ74AITOPr
Xa8R/dSkNTCQKjMD+n4uTwAZ24qmO/eVDtoet3AxfxTs+odE8oZoApBoRVCuqDiuO8aB4g+3TrVP
mn73op8qNwX8MFFKqzmoP+zTl7OKcm5hE0NwUTtxgK8g2Ekre/AyQNSYNFzo58oQCzSHx0UK9QTb
EvXGkFJxwuc8kMXns07xufEZWyzIiwn49o4iTbBeIF46K3tMmyABOpCHLqtQPyEU9qQGjk0N4uCf
UthXX1wNUdmXGvz0WMeH2yEILtJa0dXMXpKBO4UMDxEDZ7C2HHrKNrkXrAnvrYyEllsrPwEC05Sj
wWiNZlme7T8bQTHLYZRjylryTp3QTMLh3nadny4IDthP7PxaVT+9ZWgDI4WLrb+eNmE77e1Ei29h
/8PuOiOnmtUQWkT7GQbsWauX9PZiZH3hQUP2d7qNI9Zdla9GjnRiHpsQobMLdaietFDHDBTS5Wxm
abwH+aMGPGkfdvekUwbn2HcIu3PpfucsoMxqxkagpXig6NzDfdGlb8AnlJzX/U4kJsrSQussSYnu
TnGRqGWMlDPFpfoqT+0mm7Hh3T1P9Hzsjg6sNTrwzNNGdWs0fqrDB1SOo8U4b4YOsAnfza9LRqKL
ruPJI8RD45o7CMQ3ZKufPt6k6RiNJxrr7Bjp/ikUKnejl9mpEmEmp0D2JTNYgh70Hiw8J66VMZJj
sszGc+aL4Jd9nUV1smXJ9I2ftlHkrSRyBumi4exmy7yRxISFrpmWgnsNWVfXOTGHo4pgxfJ/Yp/4
6NWxrB+SXOI/2m07qi2J8z26Ne2jWQREc2R9gRzQvNFjFUMl9KDzSWDIH/BYZON8cVjqTrS3Vcw4
c+vptfu21rUGo6lDi/mWAHjm/UGCT2n9q1VtkMIxbpCa+DpiPZ60xTaEbAmgrr4BSlv3B+LnDrIt
eZWJVYnnzMjSWOAlpWEE7m2jXJFsSr+Mb+RUo2HeiSAKQ4Gqj8jFE9KLBS63KzOfaTgcOv4CzqAE
NLFq5hQ3HTZzj/L0j8aW7+HUwVnbfThukglerrpDR/KM8qPQ7X5+FiWB3L38B+0mOhqvwMDdGlfE
qtYs7THOZQLyRw1S7zS4CS/YFI0KFl6ydRyJiiuSMFyKpt6cq3fkJA8HZAvnrFyKhh1tMrN5LKA6
z3Of/8WaV/7UjQU2VELgoriBAB4B1XcVAumlC9ECy0The3p2LNJFYnd0zD6oBppq9GmplqWRGKkL
xOla2mHFA1AGwd8TeMAH+Nl+g84Iux7v6wahTLflMCclre0ztiKPYiTI+mLv34vxoVJr6/9+GFKB
HosEnE8SFutPwKl6hdHeu5xYRjma56rblslrN/EvXSiKW/86+Bc8BXFMca1gQ6vbOK9QFKRMOaGO
IS+OE3gYdLJOUf0ESz6+N73cyIprLjI7PNSY22nIRE+kSwPd+4N4wdXb/5+FyfD1D1+IYLsuAak+
nkMYh3q4edxG0dLOfP5nxvi6d8FMUX88fN2sJxxo7+gGP/Ajhr7GHsrwG8oKz2QWGLOcHTYt8Gzx
zMYPkonFMmkJose/iL3Loffz5tlNRf+bBrD2kx3N3xwD8PT+hX2OcpG8vSFz3kmygsKPbDaTYdKO
1DZaLvikEdde6cwAOv7rcIZtxxx9vvuSi8C8HgMDQv1NA0V6i7IA8lnd7dcTfcFM8j+Vg5KAzHnD
FJ+56Qm3JMMFyrZng8KYiMSV4guzNuvZa7GyolA79ej2otnx7JnHETMsliNXwy+ej8tNS7czaUND
niQ7prk7zc8ENSZIJRRadsRWmS8ZmL9SDJ42IlF6fyogQdSQOn9OQ8zr1gavlsxR52PcDXYttb2s
oPPtGtPFPE4rW77H7kzTuMNKUyLSCTplPX0OkncHcJsDlGnINLuVA/x++GgIijSpuncM5x7fOxXV
TNr0U1FIOd4PNVBzaoFS5ICqvtUqVeXiU6SmGUCzMXKZgyXtaakGcUIs87fr7mseUDWz+n+tHBUP
E1PUOYQv86mBhAWtqU9s0zuviZuV+Je34c+Nd62JOHqMufqDTEokTBWKGShL2O+aV84o30Cs3GNS
BGKjXJBTAYbn0i+j6SWo9LmcQY6Q8JJgF0ZVssnZesCI5gabZ4IwGmQat1BuyFSpeFmR537ZQ9zH
avX/XEKjUAP2zkva2cDrcBPHYCAWecVhOIyLtV8sP45svJaq4K5v0AzFAi9Klmv6UmSFhlhbaulR
y+GbJ6Nzz0WSxaVyYVuOxnzukwHDur4iEGgTxYfBqmBOLLtnRo2vIcKBJvm5KgB0/iUg+oPYT8mz
E3o+z644rslE/tAMbJseRrn3SfA5bJ9AMwj/rp8A3F9n+BOXRQFKfReodBNFO7FNe+KdrQIfU47M
cPwxx/ouifWcIacEACTX6lFeE8Jr0RjZdwXdGzttGj6oZBzd9bLA2CIs3/xqTUlxEzPLleG+9gTj
b2HVz9XjxQqaNOQH/YFqdbuYXVub9nUvdu7f242oBstHPurbUNoieCbyi5kSwwkajyyXfHmbC9JB
LexRw84bAhkkV0l4VMb6ko54gK0+OCXAwFxlwK5c6wLriZimasD/4ngOdvhyrKj0fQiwqZbxhuwm
ruRPiJKOTCF9C/mnb+GrLq6eIDZtyKFSd+MuUkn7PpBdjIW4OZP/Yhf8oHb8lYx/XSx5XW91FDxq
dHtCUPwZR4UTgY0DCNTenk1MnBXxkLt15mz1wlLBRd8VkKZzKbQPJQS87lvtQ3Q9tbKaB90dkEu9
0BBdEwqbQGwxkh3ruwJ9vc3Mnw4O0JGJiu26lgFKBb9RrP/vIgdSLHe1zwYbIIFEjc9Gc9z2MJYd
dxynteYl+uT2TSoZJNnCWePuR34Oh3+SOQR0HUIxoqxgIk4DaDrZbKYSsST/Sbbw3Ai2T3VzD9kV
0SCyC0bCxD6hmjcK9XhnOyzcPR6TKtmcqVc88gXLn5rmw3MrX6+VFEUO6ACLeFdrz+PTxvIe6NB6
L5j9Ssl655WTHI3AOo508HpgN1tmzI9tNeNxjYADlpkDB6N9JuY27DPZhAjfDVXOoJlJxiMtSb6j
4J8bkW18TldDvmRNo2VOUiLQNBDhLA4ZbwkOdJuLiW5JB0ckNl3Rqo/7/lyNAarZD3h9S5UlSJOS
rohTgiQXnylj5K0D/WlGcPOVm/j/Flav5eLMAdeaH8eTBAjyWiib6nPs9Dfy7DPGQe5lGmxuRU25
5DojcGCqzvM5q825GCSQHmyJ7e92oOQD+UYfx8+E0dX1mI7Bw5LD6kAFGdEWP07iM73arPf5lw8Q
HLIWQc2AMgHHvEx0kdDG64kmrmOZFiUrRzJT10XnZJe0ZkQqFmM9btBK0mIqpx+14OHHT3zWyTnj
1+wyX8jM0SzBDofaWuIlxrSADGWORlkU+1WAQxxndh0YUfFH+MGPUiDovil2n7LYvf4VKefczrM7
vqiwuVWI6+EFacQ/KSBjEUCdByEpBgrhfYTFNQcrM8Lr6RJ88U3yDJGcI1DaLMNQevjfkYZ9lmqv
qmrj1aTw1QKubyjWlDimJPZ4USPZKNrblgzytN1OJaN0lJN8t6k9S6YZ+R78gVtFXhmkkHaeEbmO
LFCSA47iqHvIyCSATA6MqME6qV+LPMEbMfv0oEOzJfXCEPngqqXJipxAjBs3oESxl88NFnzZdfz2
FmVfokR0tUJTt5IUrS3Zq2AA6cYY3zmvVI0V42ibCNh8JFLvSRT85CEKxDnxs9ko7ylN2yEXpQpp
UXz34bBfk52YoGzOWi9iiv0KE01MVYxQaZcHrkXK/yH4EjgRWFrEA6V4RESQ+wQ2KyQdz9gWs6Kj
NzBlOalCy0GdZ1KGUrnfNj2iMUDg2+LnoNvSi61tCUqh5BOgLxE4LaA2qxQmbCD6GMaOJqbS+diw
xmrBAYl8sDX0Bnzbuk1MMo74fyxrh94+9yC7QjUyILZboVtQKJwcHlIA+lkgKt2H98ArdbxC4yUX
hiwRjjKKiwic4/jVlx05CcRxN+QGRLcg2OMF1TEWRKL0JY95W5m8xot3cLEBjK0+AUsMFpM22D4W
T2TLEX8/gxgMMVlHShAln46pv6XkaXiqf4T4Vr6OzwwSilQAhvpGSroeYvTDStCOdDnqu/sOxCbL
gu0EYr1GzV0y4ojtq5Y1nMgskP+cwm0B9oi5K60vwCJu2mpHBPKvKaaACT4daGr6wj2iWjJLCyv+
cejayI4GGkvVjdc6EH9NhNiIodLsuglOii2DyXR8+D7sbpVO7y6pCnH4GSbh+5qIs8DzoB2iGsoD
3e1MsD2Ru7e3bLW9Y5CVGd67LRgmBaF75P2l3qwMQRYgaH/nPjbqUp3eGyGY6H5EKJ+JZlq/t5dw
LLGq3FrAVUil/INL3CHZ6ReU6e8IXZc4JWBRux5AFXdLlg7QV5nQVQQXbMiQANLYulNOzdk0QWsl
0nPaZuAZ2gkgFPX+wbY8LTniAzeQmwXeKd2zrc0GX39L5MwsCBoYtATZDBuyJbNuciRk3M241pmL
8y2J2rF7w5ZWa1RNMjl+0QPhJV7qbmL6FQhxdNwU32GQVug/Jhc6asIFS3zMN7Kig506vllu6fOd
Iif9f8XYp6sU2+a+OlilAzXytvg1YpMg67wtTPIIPJ7T78VK6Ln4zKo0DFuOqDPjsNGPmoiqQFE1
0DyeaLbxWhVQhOCYlh5tJpDEAv47Y+8HeCy1PGAQQqex2bM6tsdSbefKmXh3MfX6CAQkcEzdlhqq
9/2j+IJ8VEqcilSEu2ztReSv/aJccq0T+HOk+LcW2ZsZEd/XCxmQo2RBVBANrbZ81KFlnm0jrv1U
PUBCDSXATU5OjVq55Cc4Ekbu4q/+IjtLHiA2oEvziun6fsLcdkJWt4jl+cEBcWu7JqJiqatUorYB
zvTLRfQQyDX5LnNpRUyOj0Dfo3SX1GzanSZwGd1PUO+01Ihgn5suSpTouFKHRQ0bmXu33eYzdfn2
NQOCPevZ/JwRKvcOqF/6Fviw5arYWCbK4knR/OHAdhxFP4a2wFk2gmFUhKapzDsvXOEp3cgR2uYH
/+XSe3G5pcldLcMKrhLGSWq9UUMIPE0oAjHujOW2UxyGwd2Yi8nx35QjrhZf52zmnqIGsXr1rr/7
x/RnoD5wp9pxq8AcG+eZeHTCEythU0wqqf6rqCzoDf7cig+ogv3delHvXrG1LzKoMGdlMb3bS0fB
DnnZBNRXIkLcryBgVPipuLwsZsdZVdtzUfaut4jGpjvqdF20xS9gBFednIcwWJBqfY8gWQt88dua
UFTuVqh4fH7mulU64LLSHByRBq5BWiSbO+F7YMUnt6qSSMOESqrLvWObKfKeux4LP099das1NNdE
pLZ7V9MMxa52/JHV4BjEot9AH00xJeqWRVH00lhRquKCr1vLXxEUXAV25HL4ySK8ijFccFmOzZ2y
sR5THWUD/QHF+r7VsUJqsCtbEPA+Yc71snfD5pswg8PGXIQH3iFGAD+xnF+qw8PeKc3l1xNIKDBu
S2L/Omt4AJsnSmHXKVg3mnQWigtMbkkGGMh8bV49a1HRk5Wng4tDH5VvYYBVoAYTm6PtpA9eIBPe
j8UUc4TsMOTph7kN38wGfX1HiYrGKQAz9BxZldhBWSyGDhhtlFx6ulHD9vsE11Dw6Mva7HS6zSYd
97dUhtyKqXejSLR0fRbgo7v4zGRTr9MIYJw/HTgqWruRRR6xwzngcA3H61AITMq6Nah+m5kxYM/Y
aEnFYkvjwEW46sVJ8TRTu9eMdXYJZ78ukFiVO0cBABwlgZQNfBvCbcdyQikXbls/HYWplpd6hJIP
2f8KeQrHTug7S6mdicO5rAMCCsFhA51tLB6KZ88XjWUyzGb1dU7OdsHzXnAbf4H8HBxTC+HnpujO
LvH2qH1kwkc4JpQrIoXVRnK725ETHeIR21Nl9OT32OOCUwrBSr0X9YXFV0fFoA2ebRbysxHGbEh9
lFfokXZrHMUMIf8FEZqeCG2RjFa/0ZbD5Z2jmGRBMCajHDj7ZhWrXuG6Ld0aJeaEdShBycFye2Gm
/f/6uP0Mhc40PICDGQMCpuMHJeGHwKJUCBFtU1NVTpKAWRkvoBOwHtsDhqodB+VoPGzAUvxn+gcF
3E5UcID3TXzHx3uFImXO2UqbKXEH0y6hjVbrZudvMQWKzHmQ9KVTGa1X9o48zGcwxu14P+46+ypg
HdWC8C+w+ePe8owvm1tS75I1oEwS/H0xARi67izkt/ikHEwunNw+tATU5FvzGhq5o4do1Hse4EXN
mEd65or0o7ZgiM+yeRZ/+bsLny1PNips+uN2b5wzi5X4vG/Fe1aHWWa7yK+enw7+ancEp/gOIIrh
uO8r/ztgt30ozSf2sQ5W4TmxOELQXDZbH5zNe8hcIGHVX96wdVqkXflEWsQttF4f3WHmzpJBDukA
d+XAMNXWEylIGweu5GxqqO5nf1wBnN/6luS6qPzd5BoMZq7GNSHDil0YJqPKTnNyq0gaPGipe4+e
e1eBkAebFRWnYgKiOcyEJICO8k7SW2WxyP1qVSpkGjr95dOkrjEXPVqbFW80IAUNd9jfsIw9Q1Uz
FNSE91XDhVOD9cylN8cloJKPGqjADqKUmmhvU5NWs1aV2y9fBUwI0Sgyc176Q2yswoUDerQnOyPI
oBOCVknKLqy9ssxa0zZM0wcVhhMCvqNx+5M6w3ywVDMI1O8LL6a5rTrumNs1C+zvBoCv0ZTBtdAe
TrDSjlGWhaYlc/oaeQKtlALOhRojQ+s58vBUqRCLAhXCKSD9UJBttBSumR4nCObeTKcVhNUipOKs
EdkKeKWDRNSpMcwTj0OXtXGATIQonEM4fZTaIqm1vThnJOfEbKAETsSzFqzpdL9d/3kWbJK3/EC8
JWLI+8amqxulE3+g9BzVLqgwcz82/zrktmJJmbrULLcJM+w73h3AOap5y8qD4zfaVZSI9dFJOQxg
YK58JJpZHKRAgDiLZ9gVae4puNrsDvoAOZq7bIlD2Ywqb26v9J/HtPm8lHKMaTgglfUWuRz040qV
jjGPE3FzGtB2+wsMnkfu66uXJKlOiAlbQeYGTqiTUPK9CT4vR9CLzXFs95HPEhF8u5SkQ4JyUMDa
6/VUB7RA+DrHjUMxwEXvKeoJ1fMInTSxydRAFmmIue1oIfik/Zdum5fweeLV/rSuBUX7NncRj6W7
UVdJRmFMol45wM6/KpjMK1RXAC4yNjevrdXL3hoXsXuhvgUqXy/3dGRx+QJVf3jC0kUkK8W70p1l
GKlfUrbtY8849TpyFIlrABCwLz1XfCXS+IjXm38bIZHTdzT+eoBx+beTwzQvbmVNsqCslYZ+AZ8w
1bP50zN/HgmO076JttxoL6+Wfn8HbHpWVWRfLZQbtRuUo+w+t9pcGjCbX0GabS14rkFZj/5NZJdO
SP2084ZYrRracuJzipsFFALY+bP3mBvzmZQcfvyYv0X/Ky/NxXl5Q6xrr7uLY2mQrP7bQ788xNgZ
uFommagpTg0jDV0gpKnTxDOFWfpxbf+iKptdYFivBo6cXVfTs4JRuddZvkHlRaoeEcp9sRHDvu3c
bfZ4eexyOrFDGYCEGXDNMKQ95TloFnz9E9BCKqBSInzBFKCQjTfl/7yGa6HVRuhyTi6Ocoe2PHAx
595b+N6AUEthZSL8jTqVk4feNx2OgYkNJ5h1DX/+tVvuLrVWr9/i2fZ4VIY5bAVB5/UWa3gf5vaP
84/dxcUi7ToM32KhipPBy62U2dNIPM8E07gv3IiR5lOCN0PUdeR06uT7tSz0GgG6RVsBULfe0S9k
Dpn+eZ7uDSu+xw6eKMpAkR9OCO5s6//u7y27Jit/op+kzeO6bKu/58qx4CNwZqa04ozRhP1zBAC4
8/MwOtog0fDIXKtJdyDoUjHHpBKol7gHK+gA6hiNBxuCqERL2LICt4n34tngQk8rlyrtH1LeX/sX
d3SfQnBvrukgRtvnJVjzL4B12dIm2wJDuGtapelvrlPbojcGMyadkeP7iErj7zWR7LAuSdcHnLif
Azu6Fd820/sG7n07UmiYZCYL5CLQJqjHeO4NK/um8VATl75LEqKrxlwveF9ND+tdnsI9tcjF0FgV
nlHxMnKBfZFcgF0SieeO7nRAEyVMRRE4sKSKh7OZlnWasL0scO8U4FtMPGMt/m/B/C2jVFZxP1yi
I46l3lpOdxNe2CrEOSdRKuEcJUarsQgxW64JOO1MArFzG9j97Tgbb/ul60kl+jMARsqPLu10dLK/
LVzAFDeMfaEwupA5JpbrKv0qhnAtBQ9hgl/OK66uIOgipGyto/vf++4cIJ2gcKoU5401t3euRxMO
3SDm/ApTU1s3rYuYxNm73U8RPxuaCy1yml2RA9tj78fzhQM2YGUolDUrSgtpqyaa2thRloOgfJod
j+M+f6A/6M/kI4T4ZgVCyX/BQfvy8mY+rxJMWc23kESW5hjVlVCiXmFg0m0hk8sMVo0uOuVrQ5B3
V1HPimGdFFSksnfH8uXC1j93USJeW2t8Y9OA5Wma/6Uw8BM8mrfCiUDlSiex5dz4wd4QBdai5Hz2
PUGvmaqikuTQpxVHfA8QN4bDHNDlqUHQBQWQX+DmTbGgfPQT9jWIGc5Tfw2OXEVB6BLKQIDgH/JA
FxZ0Y0/37kRLFoxd8hapi43/sglTwqKSsiNe3UbInfxb1wrqA4WAj5GieOGlCkP1/atYsAXVT+ds
q1ANPhzeG5e/Bmh32QNnPRnisYgOw7c/f6z+AH2thE+vsrqER8RguuWIgLZcDJsdHJF4opvD7uPx
4BFQL2dAiIxEe2X98Oj4PiL87dBpSKMozIrrvzVlJPkQhl1cMd76fBufjGka7OTuNk4ASz453Kic
Yex8EQoAbOzpZd+AAMiEaTx4BemWCUIHFJar0udwAMHjTiBgmIh6TMvIFkZvxIqLRq/UiPh0oG5w
4u5xxU7JS4ZpP9PVKbBF0ar9qf/aDYb1eYoJPukYuoe/FI7w3PPOvXwwS42cdHDNOUkJ5uCn15Eu
Y3q3MDEFy91wlWapqcKNnnDeCqaIBorbDr+2gnp92Wu79pMs3Ip2r/aqzByAYfEHXfzlHB3/v6lZ
mIanH3vEmjFeXh6skvtFddbuHQzjwT7waChBpZ0jp6MXEa6lrkXv4drWly5ub8yUhjqbRL02v6nS
Orai8WdUL/lUmynW6g49xfD9L97Ns/guTfddkjW1rVdWCzwC01jbI+5c071wbI7SuLe5BiAEEZ4n
HvcvGiEdIuen82UWijnRF7mHuDYJeDQuK17LcMVdFKVR9u0fv14IHJkSmeliCt49fNGFmjKSU4p0
z8aKm8zSD2Z96lHKMKd7CB8pJUCQLVNZ8ALfkC/4M3WYCEFRhtEpetzzL81OkSEfSmiJtO0m0k7P
YbPILJZU7kGzAwcnsJjDLttq0wESkJGHAzYbbdRXEcINRDRAF1ggbjP/qRd7S4MsLpxh8qsFdIYp
xdTRHPxVWQm56zd9yka6ib734ssv6of/UkCfE4tQWczMbHChVj3FKkJc2NNeBn30mfqyGdkpId/a
vLLizra1p5Pro8vphuxH1r78ZL57j3jQYY55RgcnII6LnBIfGoFg11FCTp/Ht/VISOGRIfzojjvB
GvC+mI3Hur2FXZDLhHS8LIK8mAWs6sagsJ8FpiRAMgy/PV1H9BQ9bY5f3c/N/JtgVr0DyLB8ABsJ
1hSSf+s0Erjie4H1tTQesYWDS159Gj848ZjuaMBWe5J8fP+fNbghv5f7hZHOGBakgeG50G2AMbSC
T8G90jwlkTT/FRZjAlPR4coXRA86og6ngBSbpxxDHq2y6hLp/t5umWVY17E+R2w4LEypqHX59djT
CqLu+3RXDzNEIJnnO6+ZOeZT3+bv8ck7TwLGZ+Yy8jKBMhiBfCRwdVLME65w5aGvtdu6kYh4h7XN
arYuTt/ncUFLkf3zVT3RKVxF3x7iMwxznc1VJAo+VVawb8Iwbb0h59vNIllxx9LBbsX0BNxu293I
c5bpBc6R7B6EPnxrr1Ie3dYPQ1pAPUBeUMvNAh5sm7f91ibVDETSayYr5AKkBYrf6dA6/pZ8oUEE
7aH4oKmRyjvVFwtta8yniAjDFBC0cell+QIeo1M9Hm+ivzxeRR84ulGGneGc9IePm15lSe0pzxjv
vhtFLtK3HpOqdK9m+JR32mHxX7kcO3uiAvc+cQo8FIOUXAH3uz+BgMFPWTAZimFaTskLytoroW4H
/kbBHTgj9Kv/ki/aPUqdOv47yZMVebCR7VRdSTcDGfLb/27BUkq/KSYaGdK7RlneZKx5C1lGzEsC
MIwBLuQzTVPkyM4xKSRoQzziT4mkBFHLwMhq6hQ+OwnIlK2Z5g3BUTwIEIy7yhzOKPoSovTpAR/x
BeYz7Y1HYQL9EKHv4CNmqt/JZnhTCLYjRgyufNC0QtcAuWga/w/mTRiHt0y9+6IlrUpc/gEmGzNQ
UmTn65AocNBMc5ddrPPF8R/dUWcNNEHuAuyP8us16UCM/qVUPNElGIEtXo6xw/DqpfFkNE4BhBb6
cScxB9fAXen0eVn2KhktO8LV0/WpeylevzQsMFyhHqQ9cdsbDb8dhWx2rHVOWj79t8mb0PyuzuaU
3cYzo47m0+h3cmZCYT4Svju4xVjPCd1R/XWs+4Bb1vt4mWseYjy7BY5dd7RxFKbR46pnkKhefe5g
nfgZ7RrCdNKKbJGCJby2s1BbeMenz1/JxIK5Md9Vw+BFEZn0jx582fykr6ojI+JyEs+ve1WtlGiS
ImtGew0bqHqJX50S9LwdbwJp0dWFXpsHB3NDZGlbyeQmKGKjE5LB5EFHPiIZu6B8W4iHdjSfWgTB
cLFQf1lgOun+8IZXS9VQfQQnph9DPDlS6QXiLaej06t7NMx7S4hq/U0awl/2OV4YCxMV/KQXSS28
qKhq0B5K3I2lYzkA+47znP4kHnaeMyz8BAcmK34lYyQzMMmWMwPBQFug5paQ35r4TQDFSfDVteZm
MkoXXzYYS2ES0TI3NUnbW0a+yoT7XmOPyTPF2tq7Ku/rtFpFETzcAvpT3NmJLU4AtSSmFT1rlmrN
P1AZulNq1c/TeadmvFJZ5hwG1Gl54pF529ngc8HrhYfWIFPhzviFEmx44twgvyNaCS1JK8nAU7wT
G0ZQh1EWgB1hXpuDFTqRwv9S6OGz+JVcwh+8qOttj3XlH/qrnsWPDuFbuHLIJLLglWSk16erFwqm
o58W2WZbxsoaUmkkWbv8pMvWYjxYwFOmn27CIWWFKIpTMcxN5jm0ts1eDcU9I/LVbamhzYF7M3eL
pIZvvN6zjPmwtDLYeDdl0o8Gt8YcBkdz+QnfMSHS67sixTJvQnKWwqvlMNZykYDJm4v/biNihCd+
5y6Iv7JmXZr7ad7E4N+GGbZuiPjlYHxSy+o/6wT9+NegY+4wLXoO/T+Uk6OtrvrtF81qKW5k7e4i
QJX8gS8bwksxXaT3QvH0W0q1ck48/7abe+pjYDKoH0RjEMCNxdbmg8HRr4zB02DoXsibs3E7zHYL
n5AbP7dyDhnPJOQl3wnUcTWCjTeqkZkZBcxEzh/JTCXTQcgZwSWDiPRV8VHLRPYwcnIzRJpvx1q7
MhI8AafRvXfAjCWO/0juQYd9uppmaVhfaqHTFsu3b03kmuYgUt6yujCJ0ye7iWvCnk11yZjIBQxG
4DMymhHHlk3BakiOuKZoPQRUv4UBVF2cgzRkqEDSJWRSj1qE+FcfUYH1SEq5cq8cTL3jvt0wsZEt
MIhodrIKJ+hom963VbULbaS2tCL14pJ/jBniBEBlyHjv3GUPGmGeNI04d0AUH/9uKxbz2liVkJcs
WG8pfULXtZscTKubuF1TnyQmFFVQw2BP3FS5qycUEGJoYBsovutMb3klBKlQyxs2GPuNBMZAtQQg
lSALuvdJT2d7fk2gXVsUgFh+I7tmvrN8yiQF1ePvtd6FkRqfyjyXRoxVz8wmuGStfdpkAoJiXKgU
k8BMpYdltxorN+z0OIzQlqOTqLjuDmqeJvTEAcnDW4s1OhwipuI7prOUzkb+jlmNVh56LF5O5+/C
B1uMnfsNnH/KmmREPAGtlFTfaX69vqcY/qtWG5TrNv7fv4RquhDuuPskPGwzF9MWZNTA6RdF1FOw
z3GfgsUbzbEgSyBMf16y16PrkzbzAXn9fSMwuuhc3h9M/R9rDPfae9U5xMb/L8pb0LNw/xmyLSQc
BdKHZZZYux8usPTYq8zX2xBVtiIyHisWRo4hF7ateZOsipyBkxMNfglxTP7Jmpt4An2s9NdCmA2Q
BVFD6unNAPyZsqjEeDVLc+qju9ZG+gKI8vswgbDKjGgnryiPLKcRCwu+mIQSKtchqQxIBYL+Fgko
Y8961LyMk8PLA7dLmq8ovN+0oZwkNvPNQ6nlswhQD9msNY7iNhTbLr9dzSO6suylC4yMEX0kaIG9
rS9BYWtVddvyGPAqj09FLe12fBOpXpEnNPeGFpLTgwpkMEVAa3tkk7KwPEuS7eEZjiz5Mk4cBexB
PH2tHfuSFVnXnDKPkaYqyRE9jxBiM1jixtSPUE1IZvO54p67PwYAacEpffVJ2EgZo+aiqfoU/NGL
+irg3jkKrTYqyvhdFJUqhLfHJu8lnl/KJk9YUbjXbrVrvCJJMAfE1dDwsBBCx7N5XpcbkN0MDh/n
41eFOThU4LtNLK8yQRby4LXEvCurp+oha0vqymPttC3SG0esqp4eUVsEUyULlQdwuPCy5Lc13SfI
GGPmT532G5FFuMESI5Gxnt4/AUKhAJI5qKt40eVD5fXGNHikUUxmaxcI7xWa8nNseKpCt23ZywOw
MxV5SnohDWniYhNJA+lck0U6TpjnIlCg5vJyvGdiKltr5S/H3XOXuZT1SChVXHU1mbX7ulZRafhj
JpcDbzZRy8BpVYWlZ/jkPLW8QiaZJeQhoqdOlWngu0ShduNF/YfzKxbLkBO4ax8ayHrJ+3Ai1+cS
5AGqVutsnj3A2aHHZGNFrUR8X9UIwtsipC0pIcXbpza/XHBwqg3K7KsqxcDV40j9Zkh6HppvGgwS
HKO/lL4O6/WtsHPNr37qj6ybjSOiaqYYO9AlYMaZEHSdU/J9SyEnbrNJTZbxJdpB9ba8LwO/j+mO
jTPfCVuP64RoQK5yERG5K1J8RF0zdaEE5cAMubPjm96sOYtlCHPOHV2eakhI9rRf/52c4S2ejMhz
CNhmWWh2zwqgaFlAfrUnC2ORpwB5ODmWOaOK+QbHTFEmXsfDX6My6um9A5O+A8c9karQyKLDsp90
c/589Oqagv363RaafrQPqMVP+QRukI/6Ugic8oJUj4mkwlY6oU24bvJKFE6Hcue87F+jrL/If03F
q0df4wBOW3cIvvxki+766i7Dq8BMQ79o25vrRu/+1oZ0Bmc3KYy4CtWGpHLgqKKpTppVvVjSqlC1
2Mrmt09/hM8dv9WaZZl5T6Q316SP9Dd9egQsQfgBTVLmS+e913e+hO0/NL/neYeBjaihcqFQ078g
OYM0upaUJlcHHfhDD9w3JcKUldtcs5z8IMG9oLfWN9SHj0du3BAmYt6dCvB17M/WU/TCRl5d5LdN
JU3HhaHw4wyGohwQfFz5JJAdXFSBrQeZE5ToQBfnypoyyf/v8cMMdSfTxH80SqCgvTIlP5c59SZy
gIuLHFkTblDHOQpOa9Sk83qpNGAdC4P7C7vapJgWfWIMIB++HjyiNPvWE/eHLrq7a1T463on/+dY
AV3GPj9NzBPVikbTf0iXtM9SKgW4Gh7HK1gI3GXc3/cDOOKI6ov7dOCetQLaFiPzwX+OhwRRaywR
PydO1xIZSvjyjvAybdj6w1nyh81JoLTuJY8vuivkL3URp2Oy5VdWtiqBbwsqmQwJt9E7vMCxpxjs
LpyY7jfxOtm1ne1yYsMpZu1iq77+5j9lYm9bw9BpjQ4PVOuwATNPX8KmFpvmMWuaQ0MqFoUqjH7Z
y1HSy6V3TTmf0MNgW6keRw0ZhKemBmNwwi5IH4DrrKGS6+MLv41dj34baRWhONE23UOuOWYV0evs
TT0c99YTXCWivpbJvmnb2C4aTzSmCgNFddKIihpiIyJUBejEdg0qf0oE+sKqRIoouIGDXKGWHDo2
bX6kEgARIrev5A7lv6oTAUIiU/CrmhCfNu9oAivXbbWpe+5OYbHSQK0wEpm4dobnE5GCVJbqGfKo
CkpEqYEA6O775HyvmOOxHdnThfkmAhotUwDl1bXMMmUya4XANKAIUd/smikutnOHsdhOCT09VjcF
/ASYx5Wv0e4GlzZzTfM0RlcGiwCYHw1pfnaVgYwvKrSOWtvC4sRU3siY5fX7vmuRaUc5tlJ2mJOi
f3zHtCb4yqD08RWvBss1HMXtpw8UahPHYjkZ5rc3XAZev98mrIgVvJI0ka+clypWZZsH8J27d5cv
5HlHjdqegloQa/bgsc0Tv7p0k3FCJTVWLRsnFJRewNKF5Q/WGA9Rc4e9fq8m6lqCZB4Vlv0Gt/pK
JrRm54hyvH6+EYar1I2apbxbsEvT8MV8zdIxY5fiMxaPxnrx4YtUTdmAmQwGA5wNx0I9BfIkN8Pw
QjnInQuPGbwf4Z8b6axTOiV0EFiBqMdQDVRj4EqdKAs1W1fTNZGU1ImlmbcA+GD8GCcLvFgJWJcZ
Ih3dl/UqJq4MD4V/raLhBAjBn3GN5BiUhN0KccMVOpbqcSbiJoqkdXUlEbmwbNJjIVgUqECXnae1
/wZZeokemg1yXZ920Y2TPlHiMCIDWdg9rO+WlmXBqJNZB0mL/OdewMlTNHG7xSX4bKBqWsfu2uay
f0ckitgo04g2N4j/3AuPTx9aOzdgt0ot4WHCInPml3Gbvpk/58e+AP9xNUv3aCP3XHFBiHDywivk
jDXki570Adhp23RDrIMvocr5JqEbIxYBgSzjj5up14TJRIxVi9bYqiFx1ahgDBJymOycCR6Y26Sq
vTFWcIY0kp5EpLo9JZnvhTf/koCggjp9LfYZ0eBHJVCTro46q/8nvzJav+nhGcsPVm3dUqiv5HZE
M+WwFpOnCMusFj1t+sYLMHe1lF8iSPl85f+T8WseRDqBPQMbEpfjNlCYUt9t0+QGrCTKtPCboG1R
lhvMfREkQzY326mzlIcD+ycOkFamwU3GtmYQTCLVpKU7YK6G9ll6gDvdvKZlfXkfNbvHmyng5NbU
UABuG2SFlK5YmKRixyIoVIL8HWPa1hvLTF1UOAauFSxgYvBwzxHWBF3Bi9UhzbCn4HqxG/DeUxXS
Khcz5R+c1dgDrWClVda+CzCpyl51iKTAiD0/YMug3+2lNcjmcYcsm0aoRv8sc201nLRfQcxu6/ol
UvnaheO/GPwQ1CEU6HR1jOuSfcEdcMTCc1XjgBOuSimGRYGFhr4eryLmAnegDRdSYSTIFnFBFUoG
b+wIN6ZBm7SWT7xLJQcoLLkZqW/T2s4ayA5mf/OUH1f+VaxlJepPIVERMtYsOqPOmzFczhn4339+
vRKPqHNGuu0wpu+Bnu5mwYTdgSFFny5yQ88w8cQKvYKZ6/KgUZPeJf9mIbiqfQjq7iy0pn7hGsl/
Qgv7piW3FJprW6JslljJ71Tya6AA5sXGXF/DVyPqbYLvEzBb7d172Uey9hxU5bNoVwVWCDSd/BLv
ZeKNp+XZvgbPyAVVOiru4QL72QWg+GtsDwpQM72aCEQoRMgBtUcG3x0BVo5BipfT5C9oplA4dGai
LD6cOXjUmzhncSrk4/KjyR8sT2zPOWHTkdXbrrbF/6FC6+ZdtPnMnbpSq6rCXiL66MDJvc8F8/33
/TpwP4nHlf68YVXa51ReaN0Hv+l0it811OgQhlMSEhLOMfel6++lQH8Id6dgFDBdfInkHyIh1rVL
DmBJufLKLlJcrqMLUCS6YKuAkGsjmQwgIKQP/b389FZ+4ebGy01zyuxiSm4Hmu5Q97QlpwHo5JJD
IGuSeTjLO/3LrchE/ry/zryg/9GygMf/qz1QCYxqjlnmCdiPJgFDZTrgMBeMofwyle+MfFU5tqPp
dAeKRfCjqOeWKyehabWEQA7s54fgCAgtkuyvRK2Ms2Ql4tGXCjikxtyXR5PbKnocqMLYM2hG4Hsj
NZ+GF26AvKu5I6uobQSCnPqDAPMWqJ/CMDsqSgfP08U9absQd4evzbOjNYXVkiZsJ/+Y1v7WfrZQ
VmtLmbNc16OxQh7zS9tFQOXbnoKr+yV5ojj/lXfNhOL3yVb8N2L79Px5KV2AdRStBp+Bzxbrl+oz
HfOWE6w29REmttgXQ7MfDkgqBHlrTbe5FMCDmTRqcTxu8NoShf+dXRuiQqIEcK96yycjG+mzV5Xg
uTQPPzUZ7A4VUM87FeCMJgxtDVtZrZt3aydvi4x+R7itU2Rt1Xm82l+4uvwsYs5ODff1YAx0HhUL
igDpUT4UOK4S1icQOf8/yxWFwMXMjsJeEOjZwWWwpAAr3rNuSDKMsYL56OVtrkCJNVy5ZRPa6klq
/8BrSYTCUZWQ+XtZ+cdmNER5NHXlq9u6e9Lxm3Kn1Kit3uCuB8Nt8Oi1BV1hcFRL/OTynmxKYJpg
eGji14ixY8zVHd8wNEm6Cr7kW+v8ZoWGLN3A0keL5EpBqHRBi2i2+m7WHRyCNfiGgkt+OxbGJX8k
ONmE/gNlWPO8DK97tsN7ln17WVlBrDx1g9+ywbwV8f4rDx+yQfGx+yHS7UaTmOVRmuO7oYryidjo
gW+7zaWOkKY+dKLB3ZfupveAq2fC/9EKU0fHfJhWrdbDana5ga25MmTDjBQaj+80EW0qEgx0swkI
un/Oa0Nx9XXp5RNgQgPtK5/VVKNdcA7M9tL0GS/MlWrq1JuG2MlnFXfeWX6OirFGGhyOLtU29c2/
gGMgU4R/xGJQupdp7AQYD7ss/s0A5M8GGdsYsfo8vWnuuRh6XowcZbko67k/qPXSYPDL/8q59FZF
69A3HvzZ2QKzf63+LeAxfCcjpNPCL33sYSBfRa6D1/rrSLht20QefynWJc3FGahuuKzST2rDf3c/
2QtfSyg/6kNG38bvJidvVpLuENgWMM7dJKY0SMlBBkHgiOERNDDo7FnuXZUgqBqJYMPUl8HGzMef
qW/psD4o1JSPDNP8z9N2tyqEvaXAiuK/41hVrGDkpE0fAfYPX1cte6GLW04Hg0Gn/Zekb2RsOp08
+1oSZYMfj0lLU4OkGp83NX8e17AZ3lPe9Smu3mRQVJvrdnZhz0qsWDf9CQjHV0hdM/yP+VeoKGwj
E5l3oyimnYDcG+XBuDL9Xqi7GqIqUCRlxw4pQEdo1iGYAqQVVyBgN3bmEomK0tJep4J5UmY3gqQE
U7uYglgoC4ow8TpMmKOzZ/wBkt9C7+sIN+ve7MMjDrw/luI7bNt7cVjZwEd/1h8Fmsl6ORTUYUBd
d8wbFEQExBkfw0Gjddf2wsHQ+AE4x2blxOona6VctbFrP/XNg7K/itWDZw+BgqqmQ3z6bcw42Iuo
LAs72cY6f6YjKr57+VKMQqjni7pQ4B/4IXe62WXZnNdHVjEMa4q1w6i4+/eZnFrM1HHhpi95kxDq
tGvf/5X7BlIJqiw8jTDLjRzUMB6GMWbtD45Ma+d6vyaoQOeUE28riZAIdh3h8MdVDZCTlYteCn1n
bQW+kglBP5wHzj8/nvwNU0b0ZMr+n1T4Xcb4ExASmSRjPdMILKNQ8MNVF17m0wjfCLoD6SJlyPxR
MBFK2KbTJpnPgbu9hsrPE26ymhQJrS40WrOq0aK50BUpL1v0O7rAqu4vPjOnJbd6GWEg4gKaYnuh
ig+dzwA30Ju8IwAteiFtTscoTXWUkfKn5BEslA2qeLbGC4EbVmrpNcZT2DaqLx651ipoxnH23X1K
M9Qrrr3rhKkmUCJA6bc1KKPmP9fWpvcWub0d1jwoKqf8QGb8hZ+sqvZPHFGjgIfmVEb4Z7MjJIZQ
778dR+8qX/BwjBgw98FFLs/aXBqGLB5YQnRSl/zaTkaa2mZ0MFmJ3Yjqp8DYHDeaTTjGrawg7OJN
g3dIdyrEfyu/XsELnZ9qB0CbI9TwRMuer8O+985eR7plTnngdopHQVv3ApeUMJB8alANjFmfGSR7
iXq/dux/6bZDH9VWE8Fv4sXzCrzf/rkrRd6dqWvY0nDm7kUBGZxFqkqU9iotsjq5Pww5gahRb37Q
fAGmPzGBvW1XXxHnZz+6k33ZV1ohijTco0gmMDfrMOfJ0xJZoxt6QuoxHq0CT9EdejpI/tdnnbln
xY9nhx/pHbbx0/31F777PfMmOg8MSIhXzEvsnWZIbo2THbXpywpuSrM4Nlp0IAsI2cGdpW+t9syD
KEXy4jHnXZDCzXV3PNTP2Q6h7mSXnt4Jnd4LWJvufhghpJan6sxHb1d8k92Mopw+u5LCA3has8Ea
xpwtKAucTKhxvHq6prmVwZXO5FIRmH6cn7IDXJtdZ+D2biB10DWKnu62x9Kn7ADXvyAEv9DoD4vS
aWon0HS1qZ+D/fIyCchdBfE4K6rmkDuIIZR1BYIYDPn36iZro8aFmwFSCVFQDfjKm3nYu90+rtin
I97Qds7KymjV+YbMRkjP3kkMdBVtprw0dMWvYYFyald5gvyTqJfkyGolQV0kKxf2zy9dgVBrwmM+
ZBtRftj6fMT7jOdOCcdECIJtClXdBbFIgFhbdwqAOsbFUCY2cI5qDg+JL2J3jAsgqlj276zYBu3F
NSlKJ/z5r3N3byTG6YKZ3IWdDhjohfO4+5Dol5jtLRGaFarekgCul8Q2o+h+1XAXh6tiGSBGq0dV
i1t5dFx/W9ppfKIBO6O8vedtypERKYIDOrGBiEXg1EhkgvhfxzaobbuoPuaA8u4AH7W4qytU/0VY
jKOMG9Wp/eJvvRPqFi2WtWlrUSJ5lcDqrqUGrZXtrrdRHWMxWIl+MKMEIT1dA1EGu7g7QEOBo07y
bFEUkXlrzb0cAUy+SP1XvGlEoxfyn1u0U24hSw4WtD4Pj3aG21Hrg2MRGusl+f5RZAguWXusfPA/
C6k5EKiGf9eE03uyZ9PQdLE7BC6IcKTw8EBYWHrv5cQd1aSjN2nseda1NCB8ZY5MNTIY7NNja8zZ
9tIQvhjvafVo6ccpcO7yZj+VN4lyo+RiecVg3+iMBx/UR7sS1k9ohiIr3oLuMbgI3efAIcZ77xZq
LQw4c9HXfcZSVerD/vvT8BaGyFEu1VgxSvIMFoir7uVkMppQRwhNd6n/Fd9JZMHWq1Aon1iVnSrL
ber4KSUCwryH5//5zt47n74srHPlrHgNMBIhN5uGRquwDwV6p64JnX7ihfFMJWlsBYhmiVeEw/+o
pYLrmV7Xz4w4SBe+RcsprChC4DOvtzrZ1L/i/EsM1flx32gSeHE1N109+KAr7uEuHo2xhUuJfeb+
PeHiZZgPd1NZSW+ZVQnWfYKo4Ul2lBTvkOxm0CEnmkvNA0kwR8+o5/1uZcY6EtLLV5FaBoQriPi+
hJTjS4U0Qiv5TO8ijUFbbwQ+SIEWU2cURG+cHbo7W/KOIMU8C+L8D/4frhC/rPagXggMmW1WnkFP
17GZuh6UiakESWtWMY9Bl60yVbtQ/+5cTW5XypKGIgkJooh/WshKrgg8p7redLQNaw12Mb29xwJm
QDg0KOclvMcGVajOPV75EwF0TVT+ReIy7TUBHCDXmH25AjdTjWfUsMNO3WBiIKEQi3bW8uXmsdIc
rguYdFwBq3gjH+tLoDp2eT/wD2PeViqfuvja5sAijbrbjRgdlXjapZQzgyITR3q6z2hlJ8OvdA3t
o7bo06DmKEdCTIZ0bSl4vnVNVNbMBwe8XGrpPwlxC38SwBR1JF3yKNtLVZqYjHFn4WKquvagEpMI
32c/j+t3mBhLQTVgMZxawPKC/n6d5Ksb/ddm9D9OwAlw5Bmg4xwu82oJnHxIdfplZeG0+ZfofgMa
gPCpDnwwNinUWDtyoqP9yQgryZDgh6N/+TVEqdlbmS6DYX1eCtC2CveG8JD8s0k3UtCsOoLkJRxG
qlFEeuYm/Kz6w9wDxyg+/T0TDMRb/fJqNLGrRq+vm2LWr62IsXV8amm/n7Ksq3bSm4ZzAdixBIz5
lkHLPy04Ydk4VtebLlbjz4oCYyWunsV4InQmXfiovDPurCfJzFmWIIabq5517bNKoAC71CdH7QoD
i8O17r/wZdfIBbmuqNNDmVzgrbW5gLBGZpFvW1Hp9vHKd65NUeOGmZEDrT7WUuzPSN09PXDebHVg
iaXPgGK/Npq653t1l8cnXFo43wBoE4WYeMQrJ2LWa7SgnZon7F7yyZRbDRe/aXrrWI4mj+Ky8+x/
Y9444FlGgoMW9FpFFq521HFvn/jfF5fHorqofTH1LsdVkWi4yDdGcIWY7Y+HYB1LD+Pzis45JVle
T0lEsWvEH1vE9AOLNW8+jR4nzlVsrv6j5HN+uxAQj82c25J/HhXDAQU9264E8sD2B56l6eGJwbh2
u0Zvdfigg2297dE13kcYW4kuCfFbdlzuWDMTUq97dGr5uxC66Y/RPfINbHK9HaoG22KjF6TH+EFm
IQceRdoU704hWdIBLeubmLcXGtv0J9v9/nhtEDQc5GciwRdQHbIKa/IyYi8fTDsSiy/L74kGR+YA
FFrlDYuhOG+bwdrVYrl49+6hXOgE+mB2mH7ND91zfPNOE181yaErKsEb1Zlhxj8IajXerhKxZAzT
B1DfLl06KrhRJZXQ9NLvjNUKtkERvlkxHupsrx1ykWU3aB0z/PnBBPVp5FlZvXBtRztf8vHBmU4s
mKBFhWzwBSGVArRcLmr7fIRu2CUuj5Vy8yyfpHSev/K1kZWuvwFn8fAMuwY9KMoIFPjVaArspGrk
IBDwVvl9ed27mRCxgKtKGbl78tP6pwSaeL1mXYuOndP63/slVpO+EHIRwchcohXho6NctCfWLm24
MB36k+pO4PfVI54NSs+2LPgPvbSmGSf4cIrCWibBrQnxlGFFwOzUFQ7sb2EHi/+lXe17Qb18ZmrE
oGBwaxOeggNC+bZXYxupWrTCVIZPxatuUDHl0E3oOjnH6X0RdoBez0aY1wYRp1gSnTMjd/fqeele
npnwZO5/STHCxF0nHYcySGJHE8Xgc8GY+xF3GnixoWxnvODrcnKmRWty27XdAjQstjugosUYwF/K
+ZNbCoXDLN2RQpLIhmi0KH24pfzgflBPpnl1DOkslCc1F5V8hIz/XanPukDP0n1LV1lzKw9XCMIl
E4FHFhG0y+ZNgNyhcWKY5PU7u6ETqID2wmH9yYhu/TQMaZ4LDFJm1DLpgQ8D+36K+ajZxS4todjq
JvXGM06lj1bDWaQr85MrDI2J2LPae0sLGk0esjSqc9Ozhf87pN7tFEDe5PuaBMDekDm5XsifmWnG
4ygv1796X9H7D13ZTKY/aUkLmsmGwHNhVWNkI0OEy3vJ6empxgvm1b24tZU1isvzlaOjg/eNp7pj
vtIklhWpRNEE6DO6dzUDYpgSrQK7t7VbfBwkFKnxf0qUQ0zd/VzRbPIt2UqAU6EM5iZGLxkN5MgO
t+su60q6clQjHUKElJSyOa6F81YS6qt955whNCsKHTLv+XIDjCHn7I+CYymt/ICJ6IJaCsibNWVK
xBdD5fLQk7CWxIG4CRkVWqnr+om0bMKMbFx9r8tWzrGKBcSKN2O+LD8PpKb/TlpfdVRCYWWLp2ws
5jdmL8gOWr/Wk+bzZcVqK3HMf1ld4LHHOvpXXv1HMMUkQvSVnUu/Np162n9ELyENtQMvUg1uT9Z6
mfxyfnpnTQSBY9XvMyk5VYK1Jx+h2rEPM9GJWeIkGxlOBOubbFKGFvwsuUDP2D3AJKzRC57MYHsY
sS8kl9A0ZsUlZNGzhqmMBT3SkFtjfD2YnWS+5k+Gr8icvCsKY5/N8lpXtU8u2CtAOYLXupFp1Rq/
urpkj0NEPifPIUAhUdi6qyF6mpdUZ/IMd/GDvugQ54onjpAZftBWqxshKTYFssJuBNfdzLWh+J3m
lj1CHi5HBou+RHllLHA8VZOiBOkzUVU6MY9NcXo5fCdGGNbaS7vb40Vo0exj467PX3xIcfeMocV4
mh/aHYgl7oaMilsiVLQb5JhzH8Al/808CytVXOizbeuMbw6Y5whFEQTpMzORtfMP/veYzY1HW//f
evX5ii2OXtfteoSz7BYmBGLM0sdbs082meKmpD4WJ1Gl1oTlckO5qxwDyqw7/jVFdMnLaf1/4YpZ
mrzpFlErItdD2889BMMCmue9UKyxoNkKm6MoP+8YKiAS462f8l9YJyBNi0HcEBP22E67h0SL8uXp
zZ8+jN+gKQsemQ+TuDrM09aguKAYzE4kVEd2Ii6UaJ03w3PUPTLOI5wzlcUWp4TmZWB2m1K4kDjL
flpUNRgpbKLHzP5wKpAmFeLNOKfrfpGtkU+EYVwtpiPZW1j4Kt3eImRxAsE2MNHFPDLwYSeSPYJ5
e7PoNhnOJvAkpY6Y+GJ4vuf02yPK8Jr9nKGavhTrbtEqV7hxf++P8fiUC+q/OCasEaXNW1YTQb4u
Bf5EsLljgXXs4PVSWnD+OPZYg0mlii3QvfTyeZ//NIIBY9TQ87Wl1BLw9ikkAVcjk8zoIC6L1sjN
eKrduf1hMpyeHS3augJy1iudx5An0yXfobvoN9F9CjC2OLw1A5gEzvQ3d9HPt/TnnFpxOb90Wttj
uUdSsvkLhhRMc59HNlBSyMgn4Z1fGMdvluyllhFiah783jUrY1pc3e8tVYBbNS++9pkmSX8IIqMH
3wpc8yfjZDeFBU+n6widT2wjzxg8ZCTml1Lcoa4hHneB0G96gPC289n/lxGv4ez6VpQHtHJW73uA
Ye+NT7/hQQPXT7wej75nX/UPnwuZj9Zjb57Bfh85UjTAn1iv9Is166nZchWh+QxcD9NuNBWPfouv
VI58djCnSxYA6wt9LTGqN3tnZMed++xHlUpTwxIBCT+IQaCsGgUUUzroCNZN2PPmOdgvyCgCVH81
IR7mBzzmBCxQeAiZwp1WIBq2YH2AVd4DSmE8xpgMVf0mfZsZmExv//oeJn3JUrrw43sJtdNsLPVc
J2HhfVEDJvC5nBlcCa/30UCczKDhHfm81hqr+XWVis88sJHJ+CVH1pTIyBWofzuLrzJ1IOsiejSy
lkpgqtLgsRchQWFhGupAHkmkzWd6rIm5XWo2w+20eJRM0GK6eOwq3SnWcclotY5/3G1oL/YZAn6u
cJhguDV1RddBjp0B5Jk4Xd1WCgn3M9YpmZs3kHhwdZqQJ45CW7ZMt4UExYiHO2SosvXPP3zkwzlR
wBgNHHj8D/cTr+wYwDFosTtkE7qYKrqd/ekuu/4h/4TQHnOyAqATWaAYLZQvuSTztm3hcogI0wdO
cnDWWEdcepQTJZxJbX9cfActxH1whJDuQ+aAGn/6ZIiQuy3+223d+YatjJaaADLbXzgm9aDb2ieZ
jiA66v1lAk8xt2e7NFPonMTmpA1QVTkgNsMRa55RFDdW0uEYRRiEbRotdCdsZDjBWhuUyR/KLtDX
KvaIZORFi52sLkWSkXBDnb4abApHuCRFdXxnqUdzUjYgQy9lr880ukbK5MbXQ+IwkwBikh211jnh
Cs+nvNyGTFrzZGzl9S8JljxyFkqkKI1CHcWvVv0OZMDVqS/DLkJ9tW22dLBtw6SbkKF9AZBk5xvI
O/uggaFIA8DN330jwQL4vmCL7YWvUGa+Y2iER5GuZ1dzEJAlt4YEheCvZpRNpcNaB5oy0C73n98u
kcYtLrq9cJxYqU0aDa7y/uyUcB4XUfMfunigflwNBs3HAo7vSdm9gXKIHX/KI+oTT61hh+MFMpI2
q7D+hAlmpy7tna7dlAATtporJtO76lUaKROYOcG0S2bLMX36WqEPeRULV5Ntk5Z6kQc36iM63w++
EzNPQB5d7ZDI3QpNbRoCbtCAUGbMGVKfEs12vi1rnVA36ERubN33er9C8tMohUjvmDZNIq6EXaKA
8k06akZ3Y4FXG5+T4LswFYaqTDeetkRBXXQ95dQkKByi81+RhEwL+NTI/uSz7tEqLfg85uKGd+yf
iPU7msJJB0DQNi/64c9vNHIXX1RN7l8gJI7npl3+2skFch4pzArAXnbEl2AOgmW78hJwgMTOAYLc
LAyAoZJH1mXtgJSzOvf1VB3lPYECcSHLTxluG6++Y4v6reQBSDjKMRbpXee94Wbw6rwXZgIwznv9
CmiWbhHzd9zxR44u5Lp61N3G3dBLO1T7QwINvPi1pC1PmYvnHHfiZam6SDIHzlJ375LfCS46otjj
8wI7FOegHLv3J0w3n5aVMZhLZrgXS5GbCUeEfzgoeCtu74XIM0dsLyrC5DY16bZZW/S4kcWn+Jk7
uwJOwxKgcXXqThhNVG5iRfzHxzmiM/X58uePU2M26laDDdgcPiwkFNbwyP8BjphQ5lpxH3a8TQrW
jIPy0LlDYPixzgqfOglGickHv/tHC/bqTvsxEVT8sP2HjvRLFYLAX8BviXcrPUshw3yHD/f3CDyB
s8P4dFU4mykqrwGSvgvhaArjc3WsMjbFtYgFgeMA/6UtxageSaOJFy/nkKl4hmFvp9rPZlEIT8S6
i1CLCfOVXU+37NESqd8LNkMEH2fc3R/GEN+RkKVELqc9M8adaCfc09D0fU+IO2e2IRTpN4nTVtXr
ranosPcrwXDXK+vm9lIiuPpAZotG2nMWgiw/7FNGpmiQXDrtG/ue0TB3OQ+lXREOrEED5tAu0NMp
FFhUZm/k3ntnmuTvXozzvlCT+QFTr6NFTuJR0rMBPzOLH9sCGWHPbqzewrbABo24IhnAtETR5XQF
9awTuC9kxmEeQsBREFxSH2BRJy8qmsMoRPerThpfIbyQbGN93Y4GoO/UrfNmX0fiExVmdGQkJzT8
xPXvtGqlAl47MjQBfz06sV2Rt8b2SLWZHC0rp7ice/6F7uzv7cb4Z4Ic3rM9P1+q2I2P8ncSWf8N
r4t7L0DXBNcwMearIwn9686yDgsfT6ynWfFRBjotCDzO/JAII8TJGaOpGTw6jqdN5lVqR5ZesVmA
040zw3tGq+7JgAZKhaZxQMSnmDsz+oZqsW+aGK97fdWTCDK8Z8E8SFOdHtR1RQ9+P5k+ukoNGlKH
EfHg0VN0G+SloMXYVY6bZUKfpKZZvb1jGd3unpy88CZK1TFhA6mc4cz2Gz4qAeQrgq1zBNWG0CBm
Sw+qr2KDM/Wvf6zS7+kamGsm7BCrfKc+a2vv9FyuRk+kmwb0oBqsICqVDaOoo6J4kk2wciI7hccP
QXZe0LyU92GBEp7gCVd0Wb3SR3zlN8nHTOUl0tzSGZhRX2/Rtqjm77m2JIM71o9J+I9xT7S09Yx1
lsp7lHKlJhOv9rwlE6h549bvGDv2l7JjiWNO6FpjEnNLJCKzZhtHP/mcgwyWIXILRbiB+1vDF8iC
nOnGEpF7Y/ZV/s6bPVSNB26u2/yrQymOFT6BagflqSsWWga2ml5hErnYGRhGByqf3oe4qxvwn6qh
8RL+InUTLREed43PvSnO7DsioT5S1WT9H6FtCN95zZ1bi6yvlUbmjMCfLYFXIufmCvCAccJysRBT
0YZ2qMNUDFqoBM6i/OUp7UyjlTSk18xejQIw5UQXRRLcwcBgBL7W6UzRSVDDdGzobvliCVSuT6Jv
GLJR/lw3Zbcp6SoTjPIO2/tRQ1B2DkgapamHxg4h3qE6uO0EzTH7j5oGqYmCqtTJzs4zvuEn14Xh
BhXWAYjVlOUji/N0O81sZvK9g+Yf1aT4pZ/szou4omJvSFVon2dT5FbBrpDWL19D+mt4BxwSHBXU
xWv9XdnmlVqgEDUQ/PNjST6RgsSaDD1sAvGBM1bvw1q4HLYy6RfvRL4I1SZi3w0b2Qb4sao0y7Bo
wWD+uLZZ03KMorpKlSBvkKMW+krIe9e3pCzGAiapxK05nZsnT2oRSEMc2VpillUo4CPQ3RCmuc28
0cXQJsTEfJaFpuF67kAgRxqVjn054BOq/eGJHg+Fm5lC7bM9SEYvFGxlDUJuCcYCdSE2ot5JfBMR
Yf+U6ObQE1HVE4ajQXNQogrQ7ePmKL7JUPobn/1k46+uNR/b4+KWAFDWHoKMeO9M76wct0XlXLNc
v7pC6EGO8aM3uVSrK9XqXhfsA8p/LfFukHBj2eMgMGuT1ghqXFoH6YLrJJNE66aErGn6QO2DZOsN
fgB/lf6Htof1xJTT25MiJ0y4kIXS9GsYrbfYzFMoydETbY10b3QQ3GolobX2ltE9Gig2CA0567SV
qUz5w0LqJ18zaXe4KWZ1148jt+19kvwagap+BSfFpUziRPk7x+RSo9bGxb7BlGyzNW/93b5eBX31
320BjnwAtqiWHt2OvnINWZqKypczcaFCRkhKOP/d3My9wuvTxMQ/vSslOotnbs/FCN/Xg8bWEC9o
9UsP48oBevXIhZ6hmpc0nAXJPyLz7K+hF54Tmnf/ButRIOvngvwtlh4kqlA2/YgZLGRo+IhN2CR3
XezikXeSAHeAjIXfRV5mbTDMRs6IdBwslxUM16dV2NrQgJfSP+StPQIqIVZKGdHqAJ+yuTIm/rLo
F3NKjVKTA+jDcF+qcVvx3ZQe36XUgD2H498n50F9EDbx/aeGesnUQsZTDZaKe2y1hWr333e7/iug
5KOwMMVle9PKDGgOBbnA1Fvs94MZO9B61hZ4KHtnHMrf65ozI3n5Ln3KDQ5VGiePMxCEOeP/Fzk1
lKR38y2Pbcy6Ofjr6g8TcB/94AgT59x716zcK6R2qBMlAtkLvFP5juzwIdOWCMEIxKPvmOCVnk2i
4ENoDr84kzTOlnF5HVg+66nqbXLxXKM+1RO2I3mlXtLu8BV9s7JnE7oOxsRe3J8uCD0mNEFEgdxX
hfWv7dQfvk2sUm2xu3JcrkoLszTHmjsQxAuy/zrL34IOFVsjkf9xKVIxe4C1qwS3HBGevSloEhmY
eKzOs0QlNXMLAZiiSFvk+8GKtg3I9YUFltePWlVNUql6itqx7iWGKotdzQSvQkD77iPl+E1c+6GX
AC2zIDNf3GNQT6Ahc1p1vYP2KYC7wYcLIt/BOkXqAe1IWBDJvuhNiD/XjQ6q8Ek0qQW2NR1f/0N8
bK5LR7BcjSK4uYoteie4Pz1hAPnw2kpO1FcMqI9Y+A52zodggZgxMOpq5f2hM57PqVdPhVQ9YI8n
h3L3x4cJAiktnIyIbXk0jIoymBTKE4Um/rcKGQ8QRIBuuoU+LBobffRXONQ15yPIR6mevgixHf9K
LqPkZPOUM4SbpUUcw5x2cGKF5rPMXzNMesDRb2Pqq0FiLRpDQ8RHFndQ/g0lAOXXbJ+mN1/cSxgu
lm5yG0oRPoO+gtBXKAqadjD+99II6zrVpfIT59a7DJDsntj3fRNGb9KuV6T3LObBiC50cp/67+mc
DpgrNYrv2/QNxqKKpVOnkVgspHYzGsPDT4ODlumhy2DPJa7BbTSTgS9JlUq94fZC6OQlhodnJAup
t+Cd0iw6TP/N0hA8VKbZGqViPiMLH3D2792uf52ardSj25HNNx0XINdqPYNeogeChkcwM/PQ8Zvc
8vmHzKmKE6DNOvw+rhTwnGxGqixflJ+sJ2SfFHijL6MDkWEtX3c1g9ZGwuixrwa/Q8UJ4Y9rbBa4
xunSAAUqEGBUlcm+6lgcgxWStxdAxigS0CX53jCDy6GiC4lrPFle5oFQ+Ek11p7c3txtA89jEfoA
L7GERcTdGGloCYzdwiYUNJS/6gDmP/ehYG6vtxigAiWXmlcvksJlNK5Ah/NjDMrSScR5jwL6Mh3c
MCfgv7WVdp5f+uMaGyzhxA1fuA5lW3oVus5FJ1Zintr7Yyyj/jsdoKDM5Z1ErtRH3hJC/UVEanvo
jppr0VMcil9qFPZqW/KL4Lwbrh4yafSWb8P4opYqBED6OsVhiCFlcvmQoTZ1JC2jk0NJ2jNS+t6K
Jg66uzB37SF6gzkDJbWaPi4G7woTB0IBr0lTfoX6pHJ9Sqm4xPRH/G/AlnsFZaSPDru9g7ZNaVlE
aXMuE/XBxnL+oWoWLYaBDeyofGLaSCvTDWFCkhnkwXORs1oGsOHLhpXk2mgTQFtjjhBODs+yNUYz
VhHoCEbvhXwNXnTsmMDuRJqiYORNISsC/eExBvBBQa0RhA9u141Wdn3WS4lGmgIKQDDlw+BMu7ZO
e+oEolPFI1HL8TlpQExRybvdlOPhhQevqeWndrhk0A0sIh9FlLylco4cIMxQT5DErSAwEMfLC57H
eh7AqCYA+u3aw4TsjPz9sa0Qy12VWc9cx8Wqwgr2dadnH+Ux0hvnt6TspIlZkngbz1VJ/Y4gkP2G
ZtJz2wRy61gQKT2WSuYvU6rfrJzCf0kJjfiPNxeYuqMN5xDl69NLdN96fjtdguaNykBwT3o6BmzN
dRuwZ7g0XtGmz4StXNr2lCSCivAbECChgAAZsn4a0PQE5iNJeph6XlHxEYQj29vPXiIj6Gja4D8h
fUuiw+WyPghXYlfmqbqJ0eg/HIm9QgpH88H5vn8E8UoPZ+8J3XhvUtfTpFPOnuIfzO4P+6JTtro5
UV4xiX1FQOMsYPppQhvXxeO172OAuw/XwBpoL0a+gOvA9YxcnRqoKhulkikNdKVv+KKByDWiuSRa
kxCiWfTku+XxZEqiqfHEfMYoNeJ4mZcjjuaTt7yIsEodZhP5iC88KLSBg213+/nSh8KFyecDUD4K
g8P5Bk/n3Zfcf7PcMWxeRKuO+y44+jK3eVl4ucMWJ2x2nWmLLbRJn8PFUX0ztthlkrVWV7Rfp9nL
zOzg5b4dUohzBnekyHXrXG66hfpRo+3RV1pOLudbouZmyGLULVtOc2SgRmfyqOX6jAnUt4sMrPX/
+GMdlMrrbcg1gZ90MrT4fkhOTgZ9+o8NJYkyIa/FkuTW9MZFP+Prmq5pZdHoff0MzuzVWbntoh3R
8GZzWy9VXM3mk0UjZOCVN0VKjwwc/GO/CdeV/vPx8xBxGR/eABJlG7L0YntjAyvthwwyaUlmwkW+
I2HtHx766ivcjwf/irweAnLKvKiD8oES33g1v3hIzpbOH6OyHW/KZvBszUTdSkyJTi44L2Z5d17w
6KUGHwsO5+++nulzqo9ie6PsSYcBnQwos0YgYiBvxSnVtRxsHTQYmyz62ZdMsSvh5DZfNlOGDhvE
tO2OqE825z9ZV+T2GLkgd6pilvk0ZovuJCR2GxunFdqkL0gios3u8DVvCl8BQ+LIuRYeEZ+lfNem
GQw+bFjmqX12/oSeMbOdrejbvK8Cw1isN2TtWU/H5mIst3T6kdTD2vIo3wEdq0QESmLFfG/AVZFV
T38eWl+f17kwti/rc+eozrw920F60KlHnUbIaPdonNrYpfNtWbhY9lMaXCzu2uB8U3/cJi3GdEEp
wmQQZnMOiUNtFxTyJkyryEsA6ld0F3ux9q6V/ltADOkpLzEXd2h2rSXCUcUonxwNNBoYy51+ycba
Zhw9dDcolsJQcGA6Ttw7y0mKb26o46bEPspZmuLdJiqCQD91/ZxK2TDtbcgy6OI/Em+inKvKoVhg
3rqVOfAAcVLZmK2yUhjglEdHefJND22KXMu+rnCKF6+sqn2BBWDCb5sjqVMMeITx4TenL9t4NNsr
30J2wzHL3yZpQ1AdMA3uy9oe49uUy0CedugdEcZVYUUvEuoaQ59OMQpabgBop4ImCwpg5z4LEhrQ
+nH18+tPlKCA8GhXfy+JpHouix8wVOPcoduqyHHx3vW4RbW0tctOi392MT9yWgfR/QWKXiEd25+4
QiSiP6KcC7mqtRVslmG8DrTrOLwJApyvS0sm7tYw5fk8aTo3glW8KI3ZQY/gZyBI9BeYTv72R0np
Xw/oushwUrTrdHBuCjy0+x/Ksku37d68+9sim4EsUVIC6jyDiuMjvQSwNJ1zfYUaAVNauwiDkwCC
QgyYuq/rivFUwOGmahlweJg2xtHrtmX06cW1cf73XHCaonhhorYw9DsQ09b5bma5B6JzGaj6/zUk
ao+rmwUtLX6LvTdnHiIbYNo2zxhkruAWdRoBEXEf3xGS9wRv1taSErJijXpNXLf/OUDFJsNdheYq
4BgCFea0MwmZXzsUPkc1YpWtvW3nlzzDnZG9QKX8z6+YTXJ8ROwC5P19cx3+7s03mM6Ma4bMaBoe
c8VwNehs3ETOgaXw7lP7Mdn0CFDuxNfDIHyDOijfiFyLkxOIeFS0f7GjjSjbwNsuEkjUXEKh5CJ6
2mDh3Ni4BfNmwtIPpdTt0lblVjvwz4gZ4e4CTucD6aFPVPZgApKHJ1mMo6rrBfNZWpSfGRUQBzzO
9oxVP/gtFEPOjzc++mjEgGZi9ioOVkLmSj5/lIP5X6VFzTkAPq5Xw9eGEiSEj2fDUxoKbEeFyZqD
uKMTAav/jey3m7U4gdqYogpCoyBma6Uzs4Fwp7VXEyIV+lVv0qPth6zKAgSUHGoRsVIF6V8iX3mb
QtgTJBC5WY7AUpWLm3UO1TABHw90QcmBgn/cYzCkgx2JSGeyyckuTmnvT544kPuPcOeb3Qib/r5u
zUx7Y70U0r8xvB9J/01iUeniQVdwggoP0i/0AXAe/rjTYHABM4vZovtVGH6UQvUXf7Z6g4RG3uD+
mkZkNBAnMBgcMYOtOA7Y6e+uE6iJ6ZKuRFExyldil8FRYGkhkcDmK6wUNb0PD0CMpXchAivUCVkf
c48JV3ds55GMmPq2GxHap7UzspHkGEufA69DL2ZrQ7EP/nRtGN8XQmhWVoBADwNJpbre4ZdBDsIM
vs3S/E0LJOkPe6pBemboNbVTG8XT1LW3Sn5qWKia/NJDBCg3bJpRrrBlQU0s2o+sly8XS+syIC2a
S+qhCtWOiUEHncEIj99H5eksxy3UbUbXIJdBv0vx3Wt5cFobZQ9dt0BtFZHpqYMj6Hs65Qk7XDb5
jMjyhnZ4C4OUwEpgyKiM245JZerAyLkgDgR9pSONlLfCEQcG+jrQcQn0JpTWU1cB70Me+LbbI5FO
kd+rQ1c41ALfFsq3oo3tr6ojT2xHGwmrADf9+znqzT4c18XwLDqKDqB+sH0FsfZPvBtQs1O62tGu
cKqd5BgBe3f1DmHwT4UArQBufrmYm4kQzrCse7m9PGrRXPTBhMXhzZHVIhJ/Jxp+AYlYU9y7ybZF
Pcu4kkulbwlCv4lyEoEh4+IcE3age859u0k5BSKIEJc5QufGl4hF7Sb7AhlVPVTI0g5yZ7KQ/SNU
8eqGPymQ53V2PHbpB1YbomLjA+WgEncF5DUvzdBn5xu3u7uhoctPxw2bOgF0qBxHcM4ob9juwlTC
+w2dFVzmVShhJmXLegGToZkg0a5RHOuaBceOw3fGoutjxr0k6lzHw6d0GMRZyXJFYc6+LbiAAioY
gI6fT2w3lGribEcOHq6HmWLMSGQ4DrjEv5jwgoZ44LxLZaShnBFKRYeP099dBYyyLLba3HE7h/LB
aOhbz67HIkMatZ1PuOA1/j9/cDO3vIfeqFdWt86ComKpGH6GhR53U56SuPU1UjlM8zbFDuy/EQee
o/xAWLaooiUWtIPllXS8D/xZz+Tp4lVGyWeU6TxqZ86kvDJL6Ver2Z0Mp+EJB+RjrQi194xwcRbu
hb+ROxlcQM4lf/CUAO+NODOhSGXPvkGRUlVtdKjRcyQ/rnd3pY+2L6xjQvmiDdyKStdAY1CyLwb1
8YFd1rqwB03d2kz+E6H9sDxxBhpBqCiaS8rRY7ibS0Dfn3A7bWyZo7xRBo79aWlyfatB+KtDeWTQ
QoKsiDX2auh9YpT00vcPJUQV0WrtuUdUzJt8FCKSnguHiRwATjBQGcdijQxDpm2g4xARlxE1+fUV
d+4O04fmRGq78fNyOmgvj8NESiDqltGDyRB2mKBNxiJypmg0/0K22sbIVGsFnU16Jz1XK8wI5Mgq
KkENXwPe7axTztHKOA9xZTvx+3y2DqLsjIgRnlVfLf0D3ScjHOvUWSb0158q6RxPyrmN38/6XtFE
rMmOBy+p7RVQJENwvIgL98q+yid7Gt8BNIoGxcIJ2RzHARPPSOKEkkKKn+VExcCP6KHXjvidYgoT
Gq/I9VTuM1A3SzDpPDuhiafubwKXf2ivtyhaeSAPk//RvqTAk4Zft+DLCejqJgKTwBBKeNmHaQz2
SJRIvs4hnFfemolYPRyAIL/GgH+4NpF6rQzOcn2AHTH+dZfOFj9CmNg4HqVA88QZhAvF/u2N8XCn
RyhJntVm9Z1WDyHGEquumlWRBgxEi2Bs2T/8tLcXJLX4HsGnJNf3KgujSH9FxDk64DYxKIcdlo5b
xKjaeBjP5j2Msb0jmqfLssCXExZyAB5Jf0KZADaBiS7VJVFaf9y8eOD2F8Zd8vFx1EimC55Cvlb+
ADL84UjHiKIZ7eojv6SpJIwH56XLJWf/cICFE3TtNmTfOKoOkCkweRnS/hggYPcnh1mvD4sPq6QI
48YXFe3fPvF/+MQSFajeZiYaHh+fZh8C31FXXtvXbTv+lT5Typ/wzM30HItFJp4l8d+cvWRgTtZl
cKbeHXUB7KD3BQ8DR0qGZY70eu+MeLJG0w6QhzB8DU6SmHSTYPaFRfFIkv8eABwCPAHe0HVN5tqp
8mgxgId+a/ZEaed//ebo+AvPnYH2xabnJlwV215GTaec26dYpX7DHTx5T6zAMacQCzTnjvlmE223
Em+p5SaNzytljufMTUugQeo4yk2lPy5qUJxxacC4RFJyiKmpWbTrt6pubTnIjuzvxrY5nOT28Uof
/pN9NkmRtncmO1SS4AK4AbVu6kDppUsIjvwXEW7LqmVNjFz3XQ9D5Evqw3xd/t6SX7JFchTXPAB4
l9BCtQpONgAHDAxgXiUG08tHaDd/ADEIrFUPPvfoVQXBYSmGBaHiuEDHA8GOlQM3NuwQbLEtFfAh
y9g09vJiATurYRKt1T0+V+9V7EhCHitL1KZFvZOsYFipDBejg9NtSV/kRYYFbBPtCueOjD+3huI6
byQqYJmnzuKz5h68OnIFBTKL2CSql78gVE2B8+/P06IPvEZMOoPpUIvuk8LsPB83GczKR0r7dlw1
YjQcMp1T03rk2rqLR9JJQw/C//tgR1V72CBZ35dAsNSHtRo8NHkbbHKE8qrCuyiTRKrma80npvZF
nBOxSCNxYp8GMH8xPXj5hSbj/TghZzonIBjKLu32Op306ohPOpoW276w+M9QqK6Qdm8BjaBch20t
S21/4O7L1JMiAcJo+30r+8m+Qyxx0ZsEvy6eO4UMZsZAAD6OdCqncTDtQfI8tmL5UAs2AGIqyxCO
wFcQM/zw0GWdD4jSfXOEhZ0VYJ3iL1KePkEidr+DEvcaJqoNw0DNTykxiJIW4U7VWO8ZODkAf7fO
lFrdsCu4ZOYaOCgSiujkgvu1xbGPRHOqUUjLSaKrMrMc5kfN62gnEy95wBoagf/K4doYyqceWXWH
Gp2XpfNBeaS8c+QCXx3iSVrn0nzzgKWjyxLdK74wJdecKyoAE+8MLTBCAbIN8T/btejxTegyhOiW
wVnjBCFe6ko0FEH+M4VKL3SF48LGTxjAU1CkQTt83kUIUG81XGGajuuTXsmMixdbFHl5HjQecll/
AO3O8vZPm9TBh7wJsqijOIgP1gqH/g785AEmIzEJGHSBFsLPnwVXREi8RfnkiKK/qBcha9Hz9eGI
gTo+ExceUC0zr1927ZF5O34ih3CxsmRpkk1Z+SnAtszEyeKjEpW22n8/HeDCC6zNAPE5LbQOvWMh
VQW2HcGYf05Ju/XdmBDifxx5XZLOWPO9eyQktpUajYdMPbUsjpWRDJ9gm8Hpsw1+v8UkynBj6xzy
BHqN6ApaTeEDWCk/w5zYWqnOoyhK/k2mbJmQCha4gRmRi6G9jqf7MJ7I6tcH5Zv6pqY15lV1Usyh
91G7YfUdG1DNiAjJ8Bd8k+tJY9yRcjrtEzDM8YlT9/WlaOSTEJFIyG1Xy/+bAOmD/4BChBzz64h+
YjDp50zWClQaBSBh/qEO7LTL2Er/ZpYRep3FlMuJWFGF9VtF3lHfX1NzoILc+G+3fJkRqC6kKO/Q
r59mIXG4hf/dHL2I+hO64WpGfMGE+QJvRGLEBh38UMK1gobew14sz8HfrzD+kkaiYr4igaNuW96r
AHbRqNd7cUYzyjPlkJV4Z/uwew2M1TCP2D2s+D6Q9mgk9vk96bKn2zgV5nWFYS/qWCVGK7CB1QGA
a5ffjU/wIargE6Cgn0i+BzdUY7JH85HEtPESuBytFskNv5UKEXQ/UyQCZ021zmiFTkm5Fvf1pMdM
StT8WyqSyzccVoj8M70Fr5ojA/081N5RkhgYkU6BL2U5GN01+1k1g6MuQkPb5VIVjga/GaOP1jz5
chAtZw4JwQbrCh6W2mcZWXPflRBhk3GtD7NSf8aom6pzZznZj9z4Eg9muAGfCuM4JKFX1wnpKjfE
NLQkAt21Fh/FCISbX6Dm6hLokgpmUByqqyf4/w7j2iiYST9bLYImD4XS6dPPTp/QPinufKOVqXtZ
mGdrBuOJ43jeQC6tzmtY/7mULySS190S03ZmEA0Yw7b7Pd7u+mOY+5egyQCpJKr/Odeu/kxnTqns
ojj3X9DBQGmxAygqHuYwSCO36wHyrunUydK1YK9sW6YiK5gxxsaunic/yIR2tvP4iD63XI/al0Bu
OVzwpymj9U/zJK07txgcOVwD/9ZlAZ8VchvV+YJNe1Vr4HvdojgKl+FMPjs+EFs4cguy1Q7oQ4xd
tZlXxTVKKh+bFCRFdKiWSZ6CUoHh4McT+QB2OdW5VznFAr5MKxpbENzqDs/UeGhhhwHZjEtC2Axs
Uz2YrErE4ZowPXBC1kKPheBBVVICF6DvQB66ISzb25by9dwEPiEwpMasvzQjsjdLJUZ1O2pOo238
vGTM+mfI/1awZl1blLb8mAwNTdqwhMHIB4SSwd6SZAY1jWrpBSp5P0hloeCS44cn8hI5EehhDzKw
YeXPh93CZPPwGKAeJ73hvZLnc1vdqfZd0BCm+zC+FQerBwv0dvd5CK8K+cpUMsfbfD1V5/ThYhPb
1mXcywtByTN1bPntJ0wWQcj41wVSOMmhHmxUEbjgLzI+bkHheGlxp4nZIxnwtANhAEMLnPlXdVCj
fVtCktLddigsJl3al0hHtKGmuWWM9dsgc3pexY7+zyp533tfQqbJB8yUUSH3/oyO0SKyRNTtPfrI
7e3NZkxVK3GPXPutzoalcDOGQX8e/UrGBqrSL+9sEVsfyWWnseVv0V0jqMpqnU1Z7Fo+wHII1362
A2KKxopBvYMLYDVUEUfgm0GBC8xRnEnYnD8CZsHiFWel1Pw+oHcVUP941SwPnyD+bMrewr+Amy97
H5RdK6RJj8lBBitV1lO9csvYdSPIClcPbzJDEVYK5nh+k00WrNO1cfV122iY76dkUtxZ2jokznQl
gvuJyiy4lqpMoeka1Roos/QtiteHWT2IJ04ukaw30nMBGytZodsvMr/LXnwnX82/qXJMs/E+wtVp
B60UY0ULjCCBlqjmxPXqjMiDKNK7xYKVjzdQzT05aUPfOCjvwuZfe7mGc4ckXMH9wouYI0OouDnU
PZnuV+na0LisGYv0ACUFZDx37GzVXb6VeJZNtLicsxnalA3Y46W+mtt1kYeCjswsIxu0YNrTOjDV
HqbLi19hwM2Mi64TmpnUEv1ftOPptCVKJeswKTGUPWYEjCI7c7lxTnE9a7QrmlDCVEn1lovMrZeR
50y7HRu50Tv5K7tPGisH8XiRABYor+9MHPgVV1hvDMdbtcD3glQLs3Hvh97ueVtA5gJgzIUjGvpi
1J/Bc+fQS6AIoTDuo5CzFfsd2quCEInFiMzoKD4oKY3KWgIjdZoPwfRrffI9mkWqOOCcivNRTB5l
3sCFjREfoyXVa8cMpMu8uMIbiyJZ6VGv0y2PlmQ3V+lAaTxoNcHipuWyWotQsBJFXeqF/GXJyV3+
Pwfb32g5ZN2Zpn0mGUCZ9q9uhtFqXpnNmQtZfjMOIdwmj7iAjjG9SBTq/U4pW3uqg97HCrqQEKYc
h7ZGKL4TlT1WsQXEmH5PIJJw9bnPIcmnXY61qK0r7s3Xx5TkmDqioluoDKptacHIiPrzlHvrMYYz
57YD9aGJbtraLfYZsHTZnE+o7Ivi/lGdscrf18Gx+rRmn2raioy9jVSI0hWqCh3Faam7ELVzRREk
z0rXfZ5V6XZwgTsgSh4xgrJz2cHSkcD/0MXKda6Q1uapGkE5fuUAuyByCePpCPqlFeu5Irtawx6z
Y0HijTKkxMzboesUNKhC+yVm+mZNBnS+FpC1Phc+u9LVniKYyQgA6CdnFkZlE63Xa+IgXaCOELbA
S5lA27KAw8H9W1xyrH+2F6WmL8w2cX3wsW0B4QLuqVUtm/lVWBpzNyz3Ym2h16l0vlFjtG5c/dO3
u2Y59xVhfGJexrDL96SJjDVZ7vKWFkY2Eny4mQwtGU6qyl1KyFSucDhzL9WoqB4CTn6bI80QcvtG
NWFlSoBtgE5421O0DK1eYHclITTx88i1dAI8cARfVLRBtxchlVVVbB7vUKdEX0fEl5NeWgHpJlOr
BiJAlbTGXV1YWokRYp1yVMtyawD+vqlXGpfowLl/0zzQLXiTbyrfyJWAZN7QmTMR8FMcCYBvNVBR
HvJkOKEOz4sJkx3vwq4HiVgvoo6jXJjxk1taJZOrPGIYz+a10v6MRA+bwb/3mIHKmE0SGQvXfKDH
rTrD8DBMa/MPSAOauZhnxFsWvoQgEoKyFpIv5xPGc3lBVgQcLmxTmlsMUqMiZXyVNDd9wo5+IH+o
rW/YDcQxdFmHXKla9jEqauYb5li7xhcKzf7Tb0Ofrnu0txPgXcRXajGElmFrjze8QYIuGHfC+iJR
n4IvxUuVT4R/z1Cqu/2z1Q0u+cUE9n7/RCo2csHFswcxA2Dtbuuu2c9rioRRNE8w7j29VIjItiEv
NXOjJ/JbITvTFFuLK5XOWGFqj70AGaqly4Iu3fkgEzBBWd0b07F5TN0eXuN7SYgMLQvLlFrYWVyU
MnLWRPKHR6X0QXwZgVeriUOR4XPSwOyK6N5T7Lv54pSZgXWL8Knndh4UgHILldbUpmM+4Z0N2P5E
2dbw7EX5Ze/VvrO47HThrJ7rx+FPerXIVBgorbQjCpegEGzrAzGTn6ZqC+9droJZSIy0CFFwWLXq
GHc1rWCQAuKtsm9asUFxS7MwB8RQSI522axTQGVrikyVX88VcELOgpDhRmLabjj3euGaXfjE0HCc
evUao/rZekRxFcetKb06kNTuBjojUNx2QrQJSRltxia+mehpg8peryOYNkQEdJg9BUkgeG9INiwY
fnODFdUQiI8jghAH9KBl8eQDPKVAwZ5gsOIgkgWffr2h0Fs3tVPS5Q+jyQY5jzKmptmhPMbo1xMm
YymIXm+SOx3NHmop9NIqHptIR9IFJBQq1ULzLQbRm5judz93t6pvQh4dq6vcTb/NGzFrmPFMkAoz
HNnyrn+BYmec5VaV9mxpoT/Iz3C5qX9ogeyBHImx6wXLrq55w8U9FAo9bHCRouBYxtlFw8dtg/lE
JuRJHplqdkHHRFk8l2P/YjkJjrQHzEfK9YvDXocUcd7qshpHIDRwYLUrojBGDFeJm5wwJPhB5kgO
AnnRb4xrQasgHy6No5XUbL0ECc6X6Q0HeLOj6Wtngp+m9b5nwZTe5/AaANXQVuVS1xbENd5mgCxq
WEFeRoVCODAnW5gUP59FEWv6E9/jBU4HDA5zNDR5FMVgbWAQlP/b60dQLHl225qbhusrEOIgMczd
5XsjTIh7wn2PSeAuShgEqDMIb4Bx7uQ/hS2RU0jd6W3TCPjfwlpGY9QPBx25FJdgMbrDa157Bl+6
79qyJYW9yGNzfnIPIXFBz6Z2/W7HtwdwiayT/DYY1KqXj/gcHTFLmBFC8fqEAJh23RSocLP6oAYX
J/A9eUkRcgu66wZHhm5U18fdM0hXwCma9yRAktle0jqXjtfnvLBgCagvCqezujPlJNfRT+xB6lNn
kSh6T2u9IKn8C4QSg2lUhWvHAfHMgRmVf+3kRsuLCu4K7GrOVNArWuYfkMuOQbU99cS5lr3BWv7o
ymPZWiNpjH7rgT4liBAhdwbRZHVnr6Cos5/cOQTu8u5bInAEkMdo692BrDwmJ5SMoD9Wu/KRjWqv
XHQrirE5Jl4QQf1ewS/yap8jOpRBeXV/ljzIWivvmaPLCeCLFL0rp0fcob3WbAEeoNtET0cmYF1m
Fo+BhTuPjSXX9Lh+PNZzVZ1qsf0DG0HawMDnewepy0AoDOt1NlwYiBgL4jeIOCwgDiVkxunth3Dq
AS0sAl6dQL1SjVJnO59EvNCIVPI7Yx3XuQbEErGVb9tI+sbVv5bcTI1WMlk5covwMhavDQyGPJfJ
0Xs8Cc7veO8NfdZ0HdrKjaP3tOrw+tnBqeFg4/BWdsoX6nqx2bpGRJvUN+hjLp9XbI4KdK4BEvpf
W5bRfsoN2RwG2ifjIiMznzsJf/6CrRvgmtqn4upXkxiKKzCbx/omXtDuAGZILt4sElQ7tjr63ggA
dfI0Gat3Pltj78yjlCzWatgAU2BrC/s0oq8ew+xDSBhjKT3HzYYmuaubngvvgLaaSRD386p7Dh4H
8pKGQ/GS9L/0lRnCp7fPlxDrEjnSiYspzw2Ohq/hEDw8kZiqej/Lqn1BW4ibgpbphURHVlNvqrac
4W6Jkury+HAZbEDVKo27zDTmE9RpQpMXDgAlB5orXHuLp5HIEG2MUvHR8zFI4UpEfDsEiieQEASB
blkYBop1HQH8PQ19NrIvdq2hJC9VpMOQ1Cp2AWz1coO3d0bAg2jn1TmcobeQTLfv8FDB7bJc/PzE
9+XdOez9xlItb2HgZEIf5O+55/OAMWcKxsbo3xqI5IvJDwUlPkegXAjYlH+4ftyhiSEluB0Pyl3f
um7nFc/HjuzWlzk5mACN7wl08zX2QovlDEn+oci23QToENkiBcFpxbnaGyCtiwr4G90GnYelDtT6
GdFcVpl2RRIEC6HuEBcisFvScbwD97y2auXrC9CZbktTYXHrh8wVcM8zNQ6Pgp0mI5tzWZBtT17r
W72YRZtw1BoT++a+3wV1lprz80+hOD0A1q97yDUouUn7kg3G9BC8jlFFolmm3bCoX08ROo2gdSMY
XwHsZDj7FVLHzReOja+LZq4kAIC1y4ZL41eFDOhPepYvRAWxK10Yq/DAq9qmrc8I4MitI/Q3z5YN
UyNq0sELmwaV9JvbFxfpbhMKYP/Vc5T+tMtQVnDnFHHD7gUJUVV+FJWi8EKh1udE3f/tpk65HmA7
IWUnSKLGhupaIE+ksPmFy9uw8YN1rKFPM/Z4xZC6O4N7EtsGRSxrxlw+os1iZ/9kzq6VZWBa5h0T
UIHJsaiXSzLb/D9GVdPEONtaskdYCtjC4g24YvgFMqp5Ad1vB9WqYFRj8+kYtlhKi8ypxNe6Il29
ouRWO24KH8Xj5of7vWX2BspHocCBZv8/a55/z/A6f+J92HEq9qbYYdOQb5ZZFDWMaELH8GOcJS9d
IsnPb89Gr51ujlyGL7PEDNuKmkufmz1ljRcfJknFs2tdlLV0EN17wFa7EHZ04yaIGPLWpXjBXGpX
D+cVoNfuXD8aC3I2h6erJKIQgTqAVEKvOiISrsRrkJBwQ1jiGFcQiop3h299mvYXkTQED9Ok6CuV
MQm2cO/Fh3y9kZrmZglOri78XI4o+x5XwHS6nJr7AfbBywL3OfBIcHvpMj/0vsXnZlqbY75OE17v
mAiWGM9wHEWqcDPbmn50LeUQkNs7S/VeXS9DDHNfqgH0Nf/GVEKttuN7LpCtmD8WkJwJo1kVZx18
/h2TwFLd8HEv1sABGS12r3DnCLNBDBEIje8R+uJdFnxabfEYvZwcCf8PQkiAfU7zTR2OV9+aKIF6
+zASaMQr+onJlI1M9oEkDpqBrnV8SZGKW5hBtwFOT/VfN0Jb+LLGQ9WLINLjxaALamGpNecGdOyE
cEFPO+XkXRkpGMOzyhwrLpqGpKl7As3hKZd4UAP4XqtDFpDeW0OvY43ejHHH6JCnWfshSCDqesi6
Ln3M5QLnUhjcIYBkjkVqAempOMI82qIn+O+PSyWYJvCAFrgfMaXr7LLmL6psSqTwNoeu8AxBL2fI
20Ixs9DqWuXPbONWl/BSPRpweLmrdPSDrv5kTBiEknHDJQkxxI0GsuE3n2PLnwywdQj4ny2fVaAu
maezEXJUA6MRD2EltfhP/bDuBI877IH/NrYNI+39/i80YV77QbzY22r5bqZN2Zhuiwcsqt/3P1M9
Ga5xxm9DJx2yCO/ya5x9y2I4LuQxoB2lV8Bdh+2kElvH8RPiwS6GpGZc6cbTjU+/+ddPPDnEMbGe
8V5irBfZ5NIRn5NIfRNvoJdKfS6vgbDwAIBNS2KVag0M5Or8OuErP1w+xXvmS51ZPdkFnu0GpoTu
8ymB0KOK6RMdSpeNAKeL9BmFbkEDXwjl2fBTd1ke2Vb9spDZ8s9aMAIwfGt7zeFTwDLbIyYafKLy
oZkO22/7wP1fpiVOwik0wPEVF9hFchWdNHgwMozA7FWA6O5cxkBfojvxvagC25G2VpqwZHOLDBeg
eVyr8UUoKzjUJ4ZhrQGh4s+XO0FdYJuJpbKDmXHs9V+BxKYvdky6QEbUGsufxeZhnkqJbrrNfbNh
6AtQj79cF8c+AyctGhZtLZfqaZVLNlkSAUSyfiGZr6QEi4y9bP0cwdzdb1tQc7z2lE8NJeucUH68
YmMvIOrc1Ep38edKPMiYKzmNFBDoclWVKJe0PVyZYHCYlcXKGSLxKPEsuYx8zsA9/FHNgeS3oLaD
n1t9T1g2laOU2YckK+SkbP45dU1ADbKsY0mCPm1jaXvidtoz0f5RTw0ZTks740CtHyh5ExCZgIDK
d1m4A15pCOvT8uUmxioAuwCcvSm0HA5obnICaj/meL4OvHIWFnA7uKcVdf5AkXJfB1KQzSPPiKMW
5+R4wcFLNeoziEZ8wm7m3hqXa70KuFHWrrYBIgNeoETQ2hvAQSJyK9RIILIJD0d0V8rfxIPd+BAa
o53tIYkRwdICcSImoTeEd2f69jBb2atmyCjaLUV4Xgvp3hkjoqI+pFmO/EJuSaSyUSCyounhMC3u
xxNJnOAPYOP1tmXM4ud5951xg6FGXo47oyKd2EDkBeAwOUuGdzTdPl2tLIxpIM/DVOg9eSQaRg/f
vB/IfzHvz8YOk3t16bn89Phj+p2BzV4InacySG/KyXHNiErPb4yO2jdWwNlciiO0Y6v3kwj06xtK
wGi1L3IYfeW5PfO3VHT1+PBd+pLHYS2+9UeLJnVGmDK0E8YQzgzT2vjLeU+59Qw/rvktXiiM27WH
dPbyZn4CDXPovKSZBu3usjRXDV6/XN4Gv77RjI9tShR2Lu6JW7BvJ4kOGq0Ni8y1hOT+KUZFgkii
AN7l9x1VKqjJQDDBcWDZGW6to460b8nI9fnq9w3iZGyyZ9KsmyR7KrFVm+wG+xLoFenGyz6GcXZt
OeY0AGQdZem6qUJxLM28j8KFOUL17LH4RLUIlNYqiYpIBVWQH2NymHgzj+2XzvZPFB0SKBqY4nYZ
DMZDNTqtMtCXc7kTc213to42QcUmeMLBIsvotzDp8bHOtHz7TV9qL1HtAi14vRD5cRkYr+5ZJ4yf
TBz+pLwkn/PnKWBoNlY0zuuD6dhmLvvIcysbIUV/cwWfHF9PykFJ1o0W/SPesn9rY3z2GHPVeM2Y
heRCubJ7S1DX4ySfzs3QkCGogV9gixKa+rDikERvJkptd48ClyWE8fagDgTLOcgLmdopgXUE1u0e
wL/9HdFmd9znqFdMWzaOm/kzAuMJDBZiWPkosmQNRzQmYzrRlDZeRF9uPdQGo3VR8N0WBj5Gvbg5
mPXWFzjnCdUrwCxHJIJFaBVvJtU/7UbD4ZIm+bEIP0CE760UcOWbZMtVJuyKCAXKQOEZAMl7gT8M
8RIKUMaflHSaJH9L3X10HMxDGyKlqciFZJsDQWY4kJdW+6+fNLAYwhXoG3OMBnxYWcVyp5mCAlXv
8ApFETOCaPPaEdEM+oxTjza7JCssW1fDpKDpVKXpo96BhHhRTxqX5PIeeZE+7FCXdaV9+72tkE+V
UN4ac6VjEeR9I9c0l+em/QGiilc/FxPYEB9OeOZsDFOqL5wqeRvsEQ0j+Z+NccSJvIaGKYFQyZO1
jfBuzvPtHnWcyPO1Adq/ZUbU3kEb1wCVnLueP4CHjZmfVFGYj1wl9kZldM9s3I5vMhODjizEuyRo
s9Bf6Cy7xWC8EmYGulMhiNmckz5QDiczRfq0tnH7nCqi2G/MQHgdbopVoVOXzPK88VhBZohu7Jmv
kcIVh9eRzt/2aoBeu4Gq7u/Bvm0VT1rokmnqiLP5eRnx8DbHH8OdRq1CEqHK202OzfreH8u0mXpw
83HAEVCtWhromNodRSWHt772dLYzXbLdVt3yDtjtNfI7E7A0HcYbfsclWicYKfLjvD7NUWLh6UA4
T2Bi/VxQ9R1DNLVGy8KmlJNDUqjCTXwyeZujbrDDp0/h2ze2cWt1bpkWurR26ApCunGKKiFc4SEp
DfirwlhzKQ+QLSDp+aAOyiEqIsIpxHgsMuPybQQKg3+/CI9gcuSK/avnXfA0X1KtInlBesEb9KAq
XCPJWZOmppjCpjfIm6WRs+yiw07DdXdDPcksN8WUyVO33e1dLfX+9M8mLrm0AV16CQatc0mzNGdh
56nbBGMje2G0ANig01rNFG5A6vdzW8PWtT8BNeIft6VuznIhQ8Wg0/f70R9KWgD7rin+1pMdM2Sx
i42rDudkMqBuocFiaPwJzUlH6qavqDp2yKZxW0tNcuxXGj7ESJ4xpb5F4kMVNI/tTB4mjKvtzaq1
/CO8LxYuCtReGwYO6YmRWZaIRG22Di8rF8MbL5gEmTMOXaRVl4vsmudTTydbfq574C9/raDtlSLG
+pv4bP2CVp81Q+Hl1nN5pARAP4Xsf7LuBAHA9mbFjftiitazf+idtkCjPnMZP7HaE0GaeWKaH7NR
JzzkN+cswFMqSk9HNqlyXS/8lSYqf3clCsO+pO6XQMbWqj8Cch1jHY8WbkaLQ2rWxvzJceWd+j8O
OJPpVNuLaSON9tRrDlHn8vWywFwVqygBncCcyApOCfvrF1aChNDYGgxKviJQG1nDr00lgQtzfoBr
E3lzqLPswKfFCQBtLcBlT8R6oiGbq8YVCHmvsTIbePAXsnpvTFSrX3t9M4bp++97PlAlxxQW/fji
69pd3eXPELFuMWIrsPSm5ZToZ2o+n5xxUWPOvM4RuAH+n7fsweCRWWBNW8etxkewUp+R5Z1kuNsy
yZF/RextOZDKBQaN5sDQ+/M48P2hVx2vJxHG7ypmRK9B75ziQs0IX5wMUfbTB7F/nazHAUkT2iJT
URErn8teLXUoW7unA+vxflt6BDVrX2WEDpXpDwcaaVmSl0861KIsV3FfSgrNZuBmgP5DC7f6HcKR
Xo0d9Hku/HCXBTDdNfSMYjZNcPJW3hy9QxWlyts5e39MpVGd8K5msjoWEOyboHjZArxhN4WvSNJE
bFs2tKpraQibHOoiyz5lccLZCbe3WiUWoONonFlcmP6PMAbA/d78Ea1geaD0VpwmQH4v3/YvIM1k
3l5T6lAXXvgKanejJmUMByGScvzzfWCpFUraGD7Cqu6jbpX2/n1W5KVAawFYHHnbJFD0+qrBX8qn
79wRaoX0PLcH1MYlQym6d6vIG2BLaEOlTMURW6A62/YV+BsW5dLQTIshcdTQGr0jdaFhXv5Ie5fB
/Wy7tVfBhKwCWz/U3eZk8Y7kPUgQ+l4pjjwIfBPdI87KdIYrsDOlkARIO9IyGnKtrvRnldYN/y6W
bZWzS/OOCcloeHqRQvE7t8x0N8SfI1Y2L+sqf/01MqJQkIoFwcSdraie/q/QAGrMeFafso84uxI4
lruiHeMliIbHA9lGjhlhIm8i38zI586FtoisayFe0a4lkb1WxoyKj1Az3HLWGv7YtPTWksZJX5tj
ZhlEacoejdUSrSoUGm8yY+iPMoXmuCktSeB3DJH5rxtN/ZvsusXFhBAaW1nH91li0TsYq5shaiag
RNhWiyAI5Xi0qzwDVA2cZGDdmWhrzQHd4q8u0KJgzQpjXvQad7qC3PdWEeL3MNxseUI+MpqtFuIl
Rm2SrleEldtOEv2e3HHb8sb3FB3j1mET8YQky2G2wbz9tRsT8yKmjsnOqWHtT3Iuv/6X6PcIRrXe
/p06cY/qRqpyJQapUZkz+vrGIQdG3L8Ksf8Y7DfonE5dtoiF+a5BPQye+O/2yjrSg/6HJH/kAHvG
yeTc5lJd1uuZ5iuOqB0sTNuR4KLoowkFHKzcGhEvObW3gBPBu2u+byryz8fyvgEswhOI1+YPs4wf
4x52hYqDWxzi9bsvXELyQBUELwxoB/Yfho7GsfPCMixRdihdLlOfQKb1s46ifV012cUJSRQFDjRB
3J39yjAAiHb07SFPYN+ZwRBBLBgydrSJeXPmJ7ic6gAmA2tiQq92CcsabUNkmqphQjzmZqN39vM7
9sS8V4WkCDxUDMy12S3gdVIk64vI0pzOMkCcd+4MMqghLlUj/S2L9kWNnMzMksg5T277IxhIUyAL
RU3F9fh4GrYVy7npjrig2H69MUsFCPCoKTHHJKPEzAv90vX7G2GXry3hYGqEeRnG3XvACO6gYKTt
Io/8wtIcDy8+qwEzsoUDRHEgKaTITGcrcSYCpOQCrTUJGjhI6OtkTmfSMaZGKgBb2jhxWqaIXqz3
yIoVrI83u2ClD4+oFHp/04BTKk0fqOZmFYc8bGPELz/raxpDglOGhIt5ouz5LVv7zmUSzzqsGsKC
tshk2XDiD0TikbRG+626o2C0iJcM5S5Fy7ww7EQfhyKbZPxtW3OwfCK4HWqe3jSnt2qx/E6Qy5ac
dY8jlgGQZbnWPzH3w+S15iyUKyMi9cfY/QookdXep0Nuq8oUbMsj4QGf30c0bpQ8YnjbgEy7bMKQ
ITakgqdlrwW68iQUdzOjXeB7mtz/kBT8R59XvxyWrZ2DxNr1Nt95orPWX03S93drHvUv88izIT1q
Q90F3hMxs8Y9YFeRjPT55PwakyXQ8PCje8gzEPE7skg6auAt/fiJ1n7zf9wq1+kGJlzxdnes38/L
0ly0XfFiuVF/ZystEEhdNXupV6xOWJUwROFHprhxx3LwCEt3tn7TFJW4RAv5CefArvMb7Wjax2Kk
JKKe0Vtty64idLy6eqXLodK83gV13Owo/2nc38h/ZS33JY2KjYa6F9at5A7+n3bSf+57Y+00shjW
LFMqUeDtIjrMRFLfTRA3YVs5GNx822Raw2n3UrwEO+r4nhYuEAzoUjFfN1rvdh/zj0HmAfh5Nhv0
4E4FfZ0Noi1UHrPHem/eiuup0XjBpeWgyODn2M/dj4Po4WXUJ/daenNUaG53xXNjR5jcMUdS03Sk
7JDE0PfWJBQTxBxgxj55bYQ8RQvTBJF2B3bcvqfz6GvOpaFDluzcZP7nvnMeQnAHAnCNeNk6z4q5
QgvUdS63frFyriRCseqqO4uK+CHaslIv140vXTk/OMPrhIUCmPZCqg+9NN1nNawNGmwCyPz5eVnk
Mh2jC7OtodG8rPpPUXmcwwy8jGbnp3jaqkn6TMQXxc4bd8M5/T+gBFF7fHJUfG3TD+Vv/QZOTwtQ
PC3miwg/IlByis8NVX54r1TFjUR4vK4qj4LFA0C9zP4FdDVeMjCFlcE9/Ect7hAzRQUg4+p4lJSM
bRG/qN7mUjFBVQtnGJh4U3I7RFW2FUhIUbgI5Mg2q4ODQuv2msLlFmFeNMnMtUEJqA2i3yfCRNJh
wOYTOFnj57TR0fbt8pcsdAW1FAvMqfjeVkCs3Og5xoj4/tzVkmgmd1xaYMQ8hyZx+rwCcs1sl90B
NPTp6KpFwJvmmwVodBPs5lKzGE9ef3fSmxbz87B+dUxs4EqiA6aFtVGIuxShVCY/gi9ZNwtra4m7
bZQC1aKGq2n2szwrUGiTVl6PHgCI3aVKnduAoyQCjUoXvY923S7w5B++rgVby/KvuwWbABrq9TUP
tgAUSCwjhJTQ0rBZpvYsnj0W3PDmLMRVzNKx/95Kt3Py0yMuqTakfew5wb9NaIag1ugDY08Ax5Tu
S9zXGqa+YGUwHXBR6GknpQ+YPak/nNzeHrj+zFV2dLDFcqPjBNWvA8uJMJ3EHqZFca4ATDVBMcB/
XOltmuSgZTy7KyLbdOMi+HJkX5Sp0L6bStlPKfcZQY8z6G8nbhpcSwcvydiv2lammxMX3QegGvrm
XdaRTLa0dIkE9MxPw+M9Jex8NhjDehes5iKUXY8bdcX4fyvt91Aynp0vl37y85zQZuIJSubG0jUe
B3Vgnhyk3mpV0tg8WTcgVPOSaAlaQUE8NybuRAPoBKSyH/955bbtWWP4qN4r3ziZu1CYxTNANZqq
Un3+S+hzSp5uVyV9Vn0NxqgmHu0m4OLe/WiwiFjkngR31V9UKYQXOFasfiwyNxf0lYPmHKVgq8Z1
mLv9fL6+zwrA6slwceBYCtOvOvQvEiI46hcHrtPdnXCft52FpDmEFTxDmWOfL96ctYYE+PZym/Na
jP1coxYrtHIiNuSK3dRoetnt2D9aokve19py1xFMXJ6P+cOG8nXJhSFBIVxtZrZBB+Wyr76KFFvl
EAMRR1ijhNUgRHwoLj4aME/5qIX1cIyCjPkpW6xt9kosafxxU8td4Fz3jfElg37H5RI37U946ked
mrEQqG4SgLzEpeb+HqMR/koT1s/X4VRX72Ak7HbjgswE8EDiSRz30HY8bppdYAIwYUhMHI0s/opk
/ZfinqEQSkECFhyd552N12ZH6M+OOxYJWP75ZenMf6mZo9/EmelG9Ulct1IBq1iXhSTr/h5u++57
jo5qNKIwB6vN515X7CeARe5/lg9kN4DRzJP9PK6Duzr0anJHL2Y++uXyo8ImBkFZrkw6GJzeAltR
24p4TQKCWWpgD0xnAAY4qEQtQGg3ojfTmnnk5H1G4iezpOUp0tWIKo6iFh1m1H6I9wmFuvvF36p1
p+XxH2hZsHqEEiwPzvvmYbo2A3zXDvlwTV0RvMQNHqRjlIjE6LnZT20ZMsiDwf9sz0Ta2Q5+XNmP
pfkZvmxgksXQgcP04aKckk/SPxdLFyuwYs8FVWEArSqKhStLIPnQewfJ20B1c19bOyei7n9XYpKi
6EltbQkDPqkcXWjlLREC+ppjiYU4OUsnV/OEhvsiFiKYcK898LdJENoZXRY30vOW8+UuAvOuOK8p
Rb7U0ek+fvnJjYD3jo6VPbxvfaIL7lTucxqhixoshM4axGNOIFoF9R3lIOiH3GNgMY24J+CRVfmD
x3zSITsB6dAKimIhWZQhFmBOQq/TaKIhJtRJFnyIbE0eouhuPmCwRmOU6iHH/mKkgMQiSf+YCjgA
s0omQqK6w2jyNXzZOtafP7p0Wx2zUrAwlmvAVkUMHU7yLY9oM+b7QwaT77eVC1HqDAAqSPrKw6eM
GFUBBhpYRtLinMe+Qd7BXYJEfKw+J2BymbHvOpH1sSoylVoN27SfRD3gHImzTj7CU8h65ZOSgFpu
6O7hk55dA63I6YoHZCX2d1neEq03JoClka0oCGKkqp2uNnqatbwLYLVtcWx39V9SyrkvyMet/buY
t1qwhOjfJXpk9qyFiuAy6eDpEogog8dKZM3/wCdt3y9YeZe+3SQfVtnFmWtp27uXbCRg83AjKb1x
5+fS6UYGv7NDPu7KZzNTfVdoUbVhe54tsXn/nujQIASgYCQBG480/SRdMjCDRqkq6hI1wWMrA9T7
yLjNAAIKCRFVWLs+83VlLsdI/mzjaRdqvKIwCg4eNX4346D5ydOLeZlb9vBi+emh6nOn4G2meRwl
7DfrpLW4aWPVKiwMkavu9VD9jOpox0aBgXk6cmn6tNXiWks0mvUuMVjzz0yaxKUAjyRG2nxQPUAQ
HA6f/n31t3lcEQRXC5foTFJnFxSVWuH+iFfHlWrhfhCrCxvyKqsJm+sygi8QZLkNlLSqhla345bI
quU1txu1jU7kTLiiCXKFinPKnDodVKv9a0941GRxGyy3q8+Vs4c7KSv/aLd/dsFHpynBSGgJbYAo
HvFCtKDXlHsuCt7HfYjKnVKe6CXgO/Cym/LJuYdu83QeE0WaxVgnRUoA24RlJFcVMkiad0YQax88
mEM8+8BP5oRumfMjIbV9SUyaY4wHB5KFsFIQEIowsB8Gc6BoCdrOa2m5F5ofW1Eoh6OyhkE8ldlF
TXaP0eLZRCfL9wJ0TUyHc9mvncsRoOPtqRirFh6e8ZGNK1c6J13H/KmY6EjSmHk/FWMIaNK+Y2Hp
0ZLFFeYyzNqTqlcoA8UqMfK3AoG8CWs35MCcldgDS25OITYJav/8Gg8+zVTk6YvCfTu0s9VKyCW6
e29xC/OCGNsJGsTWwu330mHJyZVWw1aQR9jSyyxy9piS6MPSDyd+CqO4VnhDrDh1qhhVGYWDafo+
soeEBJ896tEO3KspWmcgb5/eSDzZy0RrdCNL8C2kgIVPTn4VFMQOLRAqrrnL7V0ITyAKjgTTVxk6
VTA798+GYOgdu9jZ+3SYVeWN22RH5uFURQelTLlI8h0lzpKqA5y9yxeZpQxw94oDP7C7YEbMZSXj
hAz8v8YVlTH6v89e+J5XKyLypifJOns12BiNtKnFy6UEjLFKQE0KF+n7Sv6bHIarG86LqANEzBGt
rj+BzAWoDTaY6WQqRKck5tnRWeCj85Djqc7zgc0FsNMGRyMJ5g+cxS4hVFGdt0gub9wj+eCUPS7R
Iq9YHQbG5FV5YuPFdeD7SwgM2d182R748Bk4tppH2zgjIYobCBWTcGnPRcK5uwW/YDXIgE+JmFve
5AQLDtZ/Dps+RFqQeS/q8b+lJzkGqQLNBbmcKNfaM9JYB/t0K+y7drP8J8Ajm9Xf4WHMoNDc0jcK
86GWbVPOCbXo+2Y+asxT/37n4vjQEp0n5yZeIvCp864D18h4KMh1uP1ClA1ec5kndnBdFJGntW9J
2t+AzFlIlSA4PXcWaTEqbhU86dJpqXmqH8S3U34TJrd4YLK5qdVrH4v3zyIVXfZ7/BXnX/B5tVkv
Us+IH1oR8WMQdcs2YFgiI/e4Ix71Ho2BehZkUkfoFCmiheK1vF7zXuz3Yo4bewKzteQrxcn4E7qP
lLOs2OcdLTh2cepaddu8riDdniu5RL5SQKtaBFna0pRQraA6OwhPXXHJfK3B+xH98pUGMlxEUsBl
lP8UbSxcS1FKSPGrnSpQCrPcZzpr/vD/34jYmv8+07EHET3rQ15jk5Koq8/1mOGR3S/rDRK6fbBp
pcK13bhWe5gM/b3QD4y9SXLasCPQiNUdejN3ThZcCmKLZL3yTEnI8Qhrg/LvnxO+e44iEkiydj+G
W4Epu4D8z+iUB0RpZIVyHbz9TXZASvWkHOGp09UKjph2i3NxLjJLnXyevPRngSVxMQKX0bvtuoUv
HsS58tMmiw9XQzAB87OyGfMijFZaPa++2z3UlU9N8jiGIW37LNb369+QEO3K/6aI9n9bodCKSosN
8PgKg77lU+ssZWgEGund+56Ss1Yw6N3oUVOOhMv06YzrNq8bNWan6mDR5KAAFMQ67IcMu5f7fHr3
Xm0seQGrQmVmo5AzSwjwPYhCQDg1k3gUL37ExAc+RbaD8b3/of19XiuekN4PJtyHeI1zOKSqWJO+
jsBD9zoVhkgo8pfGGjq5a/zwe/dPTJHuQxCwLkUrYnyDvd1w1/M122wZZhavsUZuf3ArYuLX4mi1
7ny/xmFOw1bGi6AYP/wVPVxXychzGuywOa9+lrGBUA8pujMqbKzOOLknF0uljvH5Z6qQwKATn5T7
Hj0v5XTCK7IhiwFHRmpDGtGJany3ubEdr6X3j3HupqlIREyhvLDN9uYtIoyNWDv3+APY6yZ3gkbz
9e2FuXLoGKk2qZLI7sKnGadn30bbkpQYZ91inc42gLObTZNQSmj1RsX0xJC4Em1UcEWE8ShAMA7A
xMvfg7zVnSqwDP1eSXml+y4y0OK08Wqmm7wdFroDCL3fi2XU9DLuHd3GdHj57KPEIdh9HulBVA5R
LqTBtRvVIjl2jnZDlS/QUQasV43FtH4zXh8VOnPZbYWf+IVjEE5mJVPPplkyl0g3hW2mni/u6JsY
pvCYUXJGGV4ie2vCBVcCthdrDPAt+0IzNUmy5xExB/oKb25Z+op9YGMrrEC07KejHZpqrQzC9tJQ
VNeSu3um6LK+Qws1bkXWXUHANvs+mjdEu8JJwrNbzVe4wRe6EJyWuqn992jHGX4Wwi/TlJDcQG1H
YVCO7BqsCHjn4QKMMSDxj//9nlxknkCGT+WIA4bvu7fJ46UN6ul6zOttgjOWyKNTBxN2Naszbt3F
0w3xCYzbXEFqVLZ5qR4ttp/QgmhKz+EFrzcqHAHhmLV7V/VdsI15mCFG6VYEub3MCe37hnl4bVqx
GhDhAbGazaQkNgI1ZnM/jeEb0Hs8V6MT50JQefBfeA1o7rLiiUMLvE3WRuzokzKDjmb6Iu+m2lj7
giV7r6cqbOFCO8Yf1HqPGaA8c4RHLLm8OLsZsxkmNr9yh1ZpZuPr1TtT2jO61MK4ym5ZCyX/0ZHJ
98WJ7NwbsmMde7xjX5bOu05XMpqqspC1HdB9JCpNgn4IiGmznDJFdmM6PEbmJm7FvATC68AYra3l
WpJgOjtAhgu0qjvvaXmfWKaxUEQXMqeBGiEu1xp+olQUW9ZOawhASK3sXaa6y7y0VFm1hhCk6tjS
CGEmQxi2FGXOHzB2EDDJxbQk3ZRBucwvmU15k15E+gq7GTF46mya1pPnOETdFMvcNDmtAymtW5gz
bciSb34d22JHju98KnndYU8mK0qvaNkM0XexYT5xR24OdbfRkemHOwfeHbqKE9KqCsvFJ6DkgKKB
amat2LcwhBb/YsQe8yZrMa2tTJnntZvOvD3Iu1TKhyQpZvKmpv7C0aD3OFJCK2ahj5UVbQRrEl7G
zLvtTYBEvveqiij9qiUUEVuM14V8cMhR3HHZ5y8k9vtCCHh9UdtK619SFEKa/bjyw/LMAaoXA+fC
AVjpIP6bYvbyf5UA195nYA6PrqGtSKkAF1YbR9zSOG+2NjuKM1UQXqAO5SR6ygn34v99WXeJ+S7T
aikXxJ/siL6SsyWiibjsEQ2B4MkvPLw3lVDIGvm8SvGB2pIdmyjx/BDt2efY0/E2ZGDowzvoSCPp
YE2LW1sFfN0qYePB3IgzJZ+gjPjowJv7VFixrykid1P8Dh7GbGPXhqeFOvdGIpmHRTOvno6qZyHX
HBbMMB9H8Bh2EwImyXzKKCvShG6Rd9TRQlNFHJeLhszKg17wxsIouV7zbkzweOB9R6Ouchqqnc9k
6k+0BcRu99SLI7SUUAsFfTdgr9sXBQjN6vUq85ZbyrEXb91iujjyEeVPrJOMYxB48kUdJ0rjt+tD
0/gtIcNQFwJXfOmQKhch1lspW0kxZ8luDbZS4DM8xd3Lxfb2SZfspxQ6KbIqDbQMKlL6spXY/IuI
yiq2ERH2uKpFNcZWjlKEyxAEyB1+x2z6j+zITStU4bKjKEplEC6uIh5XkAtfed0wq05HF31IpRgJ
wyDticXNyGKlqhRmWgipDCwEYGDI/TzgMj21ps8gQB8t8EQIK/HhPo46fXSjli+FlOkNWpOt6VH3
Am+Td+mSQ7WQ6TX9pfizUEBOqtWH3cwbYSXRdMHalwRgIZV2mhyRVEJFjI1IVlR63x0ZDPsW8uaR
lycWz/atVDUHSocGDVqoB5lup5jinFAFUl76tvuBtZkiQ7+CLa66RynLyHxCYWzplEJzAA0A96/P
a+n20WXwHqCGrPjr9f4WYnTsVpObWOCAoJ3t2/+1hlKjq3PnuVaN5Y72HlV+I6t0aPeDjbmYOI9g
mI25mCG7ZktBJ2TqPDhlXi0hubGYeV30vh41b5aXc7dA95Wl145UemmmoxyS3XjtoRI/aWNaZNpa
ynKlGMuyd4wMnzU7vOCmjz8tFhqx+AzuyqM2VLQMldZNaG57aKe8MsPReZIPrDMOksP2RQcVEaBa
TUlilNe25imsM5O2xTrzB6cFpcNCPimh12UX65bsUJAEBqSxmxNVxIeMZDV46KtM0zJVMiQhBTP2
aP2y0liCxvMNLJ/0uyvO8mo1yssF/sK7yPxQkUsSYxwTclS+P7zTS/0Po7ir/boGY50xymUnRU/G
Ipd4yx5NN7/ES1KJG4Heh0dxjVykZNK04Lwo7lUgSZvpDQrGzOrmNk2yu6lpaeTBWSRwBgcWjtVC
ommf8lXg1B+ssSWA3migIjqM4jIPf8vvk8cFO45QFqI+RyFG/8HDkITG/doSNKbXe7h2EzkygBnW
EUUa4fUNWqgoNkK7jOF4y2hydxhh+DvS78DAPFQToYdn0Txl/3F8CCOwirAnQ8UEfweBvwxilGGR
MzTtojPGzMgr+++bkCXsQ+pSgcHz87Kdq/zOxKaswEzwoczgWyPlDK18Zj0oFgNn9FrYKuQ+Q6qn
TsgLAe1Gsiv+LT3PUeuX58gCoKR0yFsjtyVU4bcL6POUrcnhPkt/FrvPEZFFSQgS5Xct2RCYVc7H
CJvqN15Iq9bQFm1tuJs39AD6ed7WSw/ulAkt08NpMDqZTV/meG4O/5JK6l2ZU5oBOof5wRnRR+zg
s5tZbD/v1oKfqgmhX6HkOi7dcZ8GPXzRNxGBLT/KNjAMH1lAwY+yFD0jL+JAxx2RhT8ZkSoKbwgj
YkR6EaUMfpze6z/sUnWJ/sL0EIgkhOkMEryZurGKxFpOaJ1bxUBjOcx2wl4qE90JLlynq+MCjOdU
CAngXyVuaGWbr72XyImZK2tlkl9/b5xK02M/l/SjsoUkOzrnnOadFEISUWhSbp4GxgPL7o6kKrsa
xR4v7ddZv1mP7bQwU0vXLExL7gQ+r1jEk9ZL8T2hdAkfGLk2jB1iFuinEaTkBlTxcceVsLCtWLLf
IzCiVWNCpgwH98WJ1IW776Ewqvjnq+7YuV6txCrzFsxPQ52oQfwwwiUcB3G2oMjlXz7kjwyPUTLq
QQ2YpwVwvxRjR3IJiTKefAQEBhoXIwuR3g+oWGf/YGBnQvnazNqMDZo3losVTgz4eooH/KGDs+Hi
ZztJWcIK+/OIAHLYpA8wm4UY+GA409ZRy8jQ9HT8x43UzPmTqHPHwFsk0TCHPnRSPX/gDBaxXoQF
I8/MwrxXMBVPIETWY546ctLo0+YH3oBh5UKcBSZzi5ZpP9wnySDpQOLQC1Pr73AtlpBNJwfbdXM5
1JAbsJyIhW6p3g62ezjx/dzBKAZfBk1y3wJaMW0Lu3lSgO9gJpcLEZDL59Qo3nexQd+czzJjQhcs
ek8vMCp2PRJcL4r7XpVDphHgfl72OCq1FpB+IekGsErB8Nl3NuxJ2cuHSgDYnZvP7m1EnOF5raQt
qYZtiht2QwMRHPRgSJghtFSEhumEdatgRJV9SogXkZChYIupFg5w13jhJMeyo/VG8U0Wk8krf67M
n6EgdlBwLpFEqYHxJPGv+7W1651hCqEPwKmTSqvDKi/U7wEiaq2n1EMq90nnBK4WqCnjuluwvqK1
5E5O31ZMcObp2mwIdKJrhdrHKuMkxUjKB58d22KCh0X0MqRTYPTG5vht3hJEuoWTsrZbbmTE92uT
Q55A/5r5jLzDvzCndY6tkjTr0Td2VKZv6iw/QO2We8qSIBXAu/0fkpuAkRYG8kxuDvHvmp67e9zT
SAAtYWGUEgTWPHM3zmBMTByUL5+oZJvKXdCP+2PPjnQJtN1V5tTawU8ZbnkGueB7cyA61gvdkYS7
zx9VaSOFc9L6Fv5Sd7gHclpsVuU+JPc98JWJ5X/Ec8iGwBycx/ggCu/WHxSO6fPvBmbBUlXhPN5S
HVrmsTcK0tB6dVJNQ8g2HZNpU8nxQfb5DhC4ho3vUeSryWkUIGFanl7Pq3oV1pqb6ZgDiC4LRPpi
wpDWXcsDrd6VTqAfk9iDJa4LUr4cUJu73ZallsXBaysk6kP2GcC4USipB0veYNHhKata203hFIYH
fnsinvOJhS3Ru0EizioUZ1+DmAJNvoZsHCQO1VyhjnhfL7+r5SKLWIcFVHpKqXcMguGjDvif9k6Z
WS65S9jsQ9yspL+hQDsHRs0LPB2iQkAQ8oSzXNxN0f5MhyLUUXlxx62J1NsjRYKLlgsQ/vVERXpe
n3osJsyRN7JgLB/tqWu/HnVmrUThrVhFp0oFwS76LeI4eTP8iwQihFscReQp07eaZJ3Qhj1INKMh
svFjV/rC9lWROyLw1Ulnh/0OKWdLGGcQKuZIKXnoLQgNT08RYz7hv7S8nTiZNJbGSXZ27Xq3/gkq
L65g+iwRFwaPL83bN88viIY9AcTYPwx5E2LuuxyUqsBse+m/Dbh00PLPoC+iCBXF+LrT1BougWni
5CbpkiY2AZKRZSAI6OVUI/4T54wmcrK8tIOEsq7n21wwbc4ea9rKdMKOYCgBvhx3sHQ+clVBTPYN
n5ZeEfvz04XiPcXDAS7JkqQO8cFQOtvj3p0uN0Le03XCKkVdZhaKuVBQ7TBRy5oZ68KdLYRmF+u+
qPb7fgZfsaTM48ddUhM+1lBeEIEs4Jq8T+vVLd4yWtcnHfk4dVgIXtxtALFqZtn5mZ99lQ2Rzyua
8Ao4dfE+d1JqKvXRuqEUWOjoZgXMXdu9r7EzWs8GpSuwfC8G+Ajeb0Hu5eoD7K97evIrp5x3X4ex
NVpW2TAWcrb24HwHofNJMIVyPGL3M6qtLMKIcjqZAqUjSYysSLZtWdvipybzJLy1doaz7QWKfvra
iAiTUL20nzKPPDseu7J4ffsr5SdgZmlf+UnYNfBeg16/VCdLqTMnTzbtqfVlO2O4IPdgbWQp7jAj
Oy31fXKaMkfiICEY3tb7lpVIJZY1HhXrZ7abO//2AmPrF7AeBv8lZTieyaVNO13Ica8WSIw5NkHN
JBRxn0MKp/bWsBvJdRh4hKbnZB6sIY7I3m5zgjx28C/Eig0o03iCiN5pdc0eTitlBtYPDdLdu1HI
UkZ3rOhYRxBE2fTbhRLTW1t2JAj423txnnwt0p5cdV79G0u2kDGA7usvtzX08WjY2PMJulzfK42a
BRUxtiYs/cjs0ncxueO0XW0vGWl/zhT6bTaaJ9yRBHrfbZMcFUgcuNDqF5rSB/hBNZU3e3bmwX37
/TrZ+w6Vo6h3LPWeeXuPSAxnO+lCgGIjUjRzza7lBFqhF4i0m9xWbd8+tjZTgyRcDxMBzq3DOq4v
SZENvIibt2KV733xpzTAc+Rj2BCYHRyLwSLUkAghR2n6CHFvB2eMaej1mCyuuXmR6lD7DTm1TPW7
kkefbLoAnHqV8UG40KawMF7gytc34szeoV736y4KPsL2Ja7pn7t7kjjM0hA/qex9fVT056FltLCm
oe6HvcU8aSHVank8s06g5m97apVMeOmjp2RQTB6sPgqXF15Eq04XW9Ef/5cp86Nvrk9mMlzFZf0E
yN+U65GQmLaQmf4jP7KnIWqNd3nKtsvpI14ToMVUTsRNszpshQRnOWyBTstrFLoCQF98mfFBs98e
MeP+B7fmDx5ty3DCwghRFnyZ5ulO//ElJO/uo8nTvNlHifAfHre3r7BVP72KkHAEPf/3qt3dnNfu
3DPQTEvt+Ziaffs3fwBrOGVkzgkM0UBfsCJ+tUli7+sP73PfUvsl0UXaRX9jScT2mFr4Z0Z5QS5L
x8/LAroKdqDNe2R1r0kijItVG11YfJ2hLbCoTBfuFCV/a7ao0QYMG9zoKCuv+6wnEEq7t9kjhjVK
/UH27nzhERgvg/XMza+Q7Os8L6zPVeF8CUqJP5XU0GvRUlfDTyFZrlOFgCSkDN/uunGQejdaYLif
IwW23UJHAiRERQrPdCV5sbXcOJJ0mP/WhL28GqPKsN4h68g4RKOzFlDKgboOILFLUMBdwFZmEQvx
Pl8YN7fZpmAm3TtC86WyTeXsDGTnbG0GbFQWfbmmZm3wjNnvRcu2hBmHH4l6shz5ljz7txDCmsMs
eU8MIQ36Io/rC9wZjUpWD1omUExlbBLb8ehpZhXtt1zBtpf6rO5CJZ+SWT+hz7MjeF0fSURrMruY
Fz2RK2LTTB5g6xBYHuAOHb0fcm8pII+waQkAHAf5cztpa4wP90GhGC/JtSw8cQ++ddT6YhJsQF9b
edaNOAEhnDl8vLALt/Deh61uCAKfj0aL0VYO7/otX+PcCHKBp4fTWMwg1u/vB1/g8vIuuxgBbhvg
K1o7sF0Dv5LGGQYiigQAtpIndtYSHzO/w4VBpE8WocrtYi5jaBa17AM4KBGlUCFEAVk+NfB7WGsF
pXH1biquVGnUgKkYpDETpTYssUI87tDWLzh8IOkCtXhoBlppYmkMq26LewxHnAC1z9lNvWDhNKmG
ovxh/9d8+crCFpjZy84YZS2a9ybMHkILoJ2uiTk4YR6jNG28v6Cf6//VfQl3HlTGKvOaHH9JmVA2
qMOFrih3rflCydJ2knS+w8NQkcMXxBTRo0saaWurIpMXmjDQ9pu6QuzMOgr9BSdiQlZgm4cz1/w6
Bq514xUV9KcQq1fxNEBGC29g/i64NCIHB/EPsMrraJHIhaMYjdkFw/V0q1sQ0+i5jr7l0maSVbfy
5P/iIVGlsBJUoHRkUvx1T0OzDCfb+3erty+MHSPPWymcqmu9Lis5NcMHMEwPccSs5p+CFQNa+nA3
gm62pre5XJduXKdY432njiX+AYiFLNmY8SYXCN2O6flCWx9AQSShaNZPzV/Dtjyfh7ti+aYAhrBL
W74WiNeIyKi8kpI4+m6bMEXG4CQeVfx4WQPpjzEd+1jphpJjRwjppdAlA+hyPz1A4EE0aXSrQ55m
j7QbTmmPoKMhIt5QTj8SAZx+SKJP+sDsQrQFjvnTP4d2DFaFnX0IaL+L6lXYWH/BlsBvuRG2zkpk
6HukVLuTVqUAYtUyy2CUNAqiLUhQTXCD6U7TS85u6yTp8Dxjh29l9LPlSH7OSY3FfXgM7AcIvHrJ
w1GSZHq77EWQ7NJOmb3G6zDqSD3KNeCg13EyBDY419vBru6lsnBvVBEGcuRMWmN8xt0SDyMDCBIS
pG6TLFjmSErhgQW6T0rs59cACy48nUOjPnkSqf8CH4Pthi4NZUegyRTM12roumyT7uaV5Yg7Qpej
Qforv9Or5p0WLcLTP7FLyF/RkZANYUwNX7QVGX72cuXew4drz/D9KTFMRBgMGTFCtsozgu1gO9Ua
OpHHdEPsN1+LY4VUgDQFGi4IVcs+uBpwViMuwNaWvV4NlfU2tizEGFSaEuTmcxhwVdAr5YhPw1lP
3sSqBrYG9/63EhkMwnTTPm/rU0NgywoA0tSr+QEqnHOL+aVHnLLflgiQZD58qXGv522gw+8MvBv0
JbUhCk44c0j3oCObKTtUihrhfm9xjf/Wmtc+RYR1esDcXPgOE6QeaugFhszFifhetTJfv+L+v7LZ
LgEOleZHgKkp/DuPzhXviKvlhGlXP0PNv9dQ1xfGpH4THLLzTm5YppTX+OrS3NyxoThEd9mTjF2A
EvYfifLuru+4vgQASB45vTG44SSdjer849Lpx54Qn77fmJb02U4HrM7WBvjLSfIZRkGgkB9v5wxo
IQcaGEDv4Z+FU5QpWS4x6gGAuW2cMPc1Jmn9ARm5UvNrBuHaCE6UXhxPaLNxSAikJX+Wy88ES+sz
ISPyEA4OrjIlgLBgaR5cXkw7pGupVZs4ql23AXh5g+HvA7I8fJrx4hPFdfBGXhKJaOHdMgeKoieF
nC/37DpFaMq9f4nuPj3nhN+dr+VtBbfEq3QhCz2tC39LO9ebYUKmXWNB0LUVs4RmLqeyJxy6a+Ls
eq4nWSUD6aFnZdb6jptDF4opNJGErdSDCGO/j9K0P5lTcIFjIQ9seTNlM+g1CgMhVL1rBrDa4pEq
zW1j0R3zMGHINfJ0TqkV83fAxVLdUjhqwuyV0sJZCUMfCqy6peYrLVnRH3OM9SYdS5h5yh4rkhah
N5ATmPs9ehC6mOKriSQG1vovS0MgVdGsMmQvVH1sMcUnw0Hx+dlD9GPRUnVd/Np4HH2gLY5ejWGM
5JXtAtn+9+K5804WjBOEgIYa5rFBcIsn/G1Ys5xii3XFFHBXJrDIsZVFbzku/P8VHBPj0KZjdzCH
gea+iZrwtarmzRVirpSOmP0rCGaPkeGpy/M9ryVIklVsHH7njnZl+iJOSTWA+hQ3fbIp/6gyn+yK
TIxopBvAGY87HYp2giDPdYkkCBEW6OnhgyfXmOxyWf+VpRfTNj2QuQbaLGS1LZZRFIQyKlaeJqok
4WpsBHvdjA4wFQNQFp9Q98l6I78y58nYCpwaFDVzaqBXs0eXZDYrVU63dG90WifYRJ5m08TP1gk1
NyRI/KUnUxtWfdI/jGPc9Vnp3BGVpi/rWQlspOM5nCJovlGyUTvhk2SMtJ+WY0jKlPWH8nDdu1T5
E0EeKbvSKJOwrr6gTTD+iGLiExt8k177KVFSCD4jPTnkvrxNH1WH/ZQULv0etNjIPpIlhuoqjItE
sKat1JPQYUdg9/hXteSuikgx6ZuBFCY6TRstuBrnYdC9814j6mmsGkqZ7pr1YUnbiWv1cRbtpE+A
Qq9EWNeM9zu89fP908ZUzHe1Fx2c+oAFpIQ6t949asDyeeXgYG304+nbnmkCFiWAhV5gFpgyG/Ah
chL0TL5pvglxTlk3fDBBT8VwMUCqbajBl89tqbJnqCZ1auWTJrEHbevvAicq6URS3nzhPfpMlZGP
f65N5eZWrepRNk/m9K7AaHQRBsckVL0O5CLLHnAyYxvNXaFEDYZYR6Y/B/N6Vwy2xJ7PLD/eo2UO
2lUXfLJoEabEWE3BjyQfssLfni+SQCT1FxDJrJaZvljME5u6ea4tRIXkiNSqM9lPSyBBobnvNH+q
mNZx1uGSBpw6y82QEeynkROfK4PkAddGbLs/Z5TJkVwEfgQc76x+UcvbL8ymsK3uFp6xg28F9ynf
5HiI1nihLzR3CifkfnmnzKWWNbHZ+EiJX9xl4CzrHQWxjdrf8i0/R/69t5TJ3rfEpl7okl6EIF1V
1Wmw3G+CWtfQyZ5ItX5rQDCUmuxbMVj88+6xmiFcWLsQfFuMwQUZtL7zcU/o/bWtVzobxwxE/1dO
qYy6bicqZQhFD/jtTaQ/G2kmKpLiH2wyFmtX+1m47vvYNQxF1Vevd+CwQ1wPeT7IWZw5FqNCHQU3
l0GHSw8d9QG+SQNVQP9U73FJMX4vI9c5T96JHwKvce8m2g4+aQ3UfSJxKUPT6JfIk+DDT3ezkTVO
ae5+oPEbbMeTrVhdK3+DUqxxe5VsYFpwtqo/19SOE2+ttZeAsVN2wydBh/NBx79xQYLUHK/hQ5ii
wT8Vj6ddw878qltDuEMHL6Cc1aAc9Mff1HIOUcoqIvm+ZCnAXNO7NGeSzKDdg5lGx2n4bpjpo9KA
DPHxP6lRWUAXPP05Cvd1vE3Q2BrrfjcWBzWJHwips6SIM2+ZQQbXW9eRZANZ/eVWrisHWXx6vo1o
bUtCTimpHuAoLowf5i0q9mgcCljZjlJLNLvr6mq9llEwny74EZsSFB1jVqQ4suzXKxMDeaaS6Huw
chgsBsMYaBpT6e1ywX3njsU9PMwKGzMzaTgMj6YpMcpgiK3AZy5K1cdjOSz1mz2I7THEaE4xUmWY
ZswY3SQNCEy5O7fucroK70xhCokcue3/gVUQLeB47m1yvibeCsYzg4506GayQmqJU38Oo38/uVdm
LoGbTw02oJcGepFg8cH76t7kmCXtSHgXBvT9RIFyWkkYYY14Li14sCzgc8RfbuBqGO/72IKN5A4l
Mf7vp9sy3CZemE8AWcWCL8A3uhuyvT48UZdgodIchZmvsjHn45+z01/U48G8bTluO4Dt5rwWhEnu
2z6Bnlg8wMzOhIzh5MouwOZeVXmLpCs5o0il4XbXH6dIEN9s1mmrT1KzndRM7cHUlyRe1hLy5wuZ
/nbfN4mpGNcbzYKamPLtVpgeR++pyyQQhvsSjoOn8k9pqwdXsiwGuRVDN0Gvn3biqSXjWPZWkfd7
XtE+EPZErSWZZkDfWI+P7cB2dNUVwDDRmolWSQJSDTtX6aoVp3NfpWvFtsiwjL8O/xm+wWrhp+su
S9IQ3gJh0xHhOWv/TfusfPwWnARRBqckYNwessypfgPCa9XxWuI2a1Lom+xa84oWa1xmMJZJCzJI
kD5N8ses9eTqBBYThM6z0BkMv4KD6j7B+CDM1zhmTmAzvLxJN5y3qEQ0Eb6MJMjmmQkuaSHPD43Z
mwV20JE36TGvaL8tUYygA6b+C3I4Uw7Xi0vV/kjvG5r9UoP4XgNcwr3G9abGCB1UMxnYrYWiUzX+
GyWGp+88LKGlNHwf8KjsCBnuwhO97foxs2KqBhry27IUm1UsiLDTDs1wbMyjB+PRnNfE9oMQJeS/
ie2PoyIBHAMYk07SEehPSWgaCgwCKnRAgQUisraAYz2ch7wHTR/EAqQo5yUewMd9RRBtLpwa43UH
+ClQc0J2TTpDHNB2a0zZQIN6veEkWGooTyXC2FsOWwjeo1fyXbHSDjqOh0ZUy2RoXv1YaKQ/0xd2
kpN8O5Fa0WazgSKaVo0251pN+8vhHTEXWzJJOCxW7rNDdBNS/MCw0ApYqsGLJOGgdA+d2wBsQt1z
+i9F8S3If84J4vMDALxq2Lw7ijhPBXOQukd6p2hfs67tf/T7io7hOaK/anr91yDyBZc15kUYbTIy
7L4ZhnysmekB/TB7OkAFvFH1MbeDuHuYht+v5pD2eXb5AplmbkOi3z2YR70SeKAuaAc9RGBgAZRW
q6n4NLrPpVs4z7otHoQ4uxOiJWu67is5qSst8jcmsuqfQs37hupIpd2EfuGxueBx/cCYsLZayg8q
LeKQUgkJ7u72gZaxgt252nvovhGYCaMKQpnirzGPuBpJca0gN33MH1HEQfnzySpQLScEUybFTmAK
OFP1h2pqGprSFka2pzruNSWBaA6fFoCKMtHA6rXMEJGTCzNjtrRq3/LpoBogVVxwTZFcD0FNsh+z
W1W/BEDwKcwmdiJsgewoFkCM7+Oq+pvdhGpWABfNk7/4Pt90z8u3S266qlpDeYiKpoojYrsk1U5m
hJ/KUyLnGNT+fMaeFDoOIEE0JswngkLlcxSPpWwouawbe4kvf+8gOOjjNZahsGmUFRuMx2dJCx9E
jVTnrcugVuJyr9mpjkT/3PutR/IWyTEweuaojPwlViup4pWscWGs7Tw58bWzhrpXXQ6tAPaHU/XU
eJL2DuSP5ziPp34jwUEVPOzVStZFnloFi8/EFvX+UGDrTF09+8zUlOPDj1pRg7+DUTXV02D+zGF+
3UuhRbCKSWYP/Cwl5Z1GYPXszCof6ugEqsCwCZyAgkaVNJ7fKoF4UPIH5dfpDhfOGHhbfKTf+Hb8
+us23e8kxp/EVDuleJkJo77MX4+nJoWixdq5yWS9ffBZBEBVcTvqK2iYHRbN6BMaKkWSXjWm56VY
QTpbbF5UpKTHselgfTZKei178PZUhevQSJ3RhIvdxawXwYh+Gjv62y/TRWzvGCl1Ran2BwreBYqp
eRo0rXsm8YVh8996573JkLa2KXrKQK9/daPPTJLqS+jk6DThLtfhOUNH81zInwnvI9820pAGlL54
P6KOpijn8J8lMzFDndKK0lxImgRYRb3/zb98zLHsQ2NMYGpWHYNCbAgReyJYd1gt3ZNdeSUQKyIT
j4RFvt3oKYCbvopQllgzqqBAAuvhYvyOpLGYicouUSzS/mHOwbL/xm6zuX2NGZOVq7NTryaacTbV
NKyT+ozTQF2FkgejtzVuIviG7o5Hw0g/v1hcnHcQK2ZyMKQrMOq5q17odhuMlkHMsYCGBuapAqMQ
QbVJasz2AWsKlxQPiO3u5l0P655wW681xzoRWX9YUD7otX472icB4SfeBWtI8zItHdEqBHqWA59U
LocwdImHiTSK1INmbaxqzbVYWZYJyqDLUodYcgrelfiGqcMWeNPdKTofj1C5G7qAdWl9J3SGcuWl
Lm1ciLwhrf9Uw346eXQHwg1w25TZRVbQcyubhCTh/MKYLDAm8G6Lgs/tsNPcUTtMaLi84XTuYSnS
hLMOIe3FPVZXjDXk6dLR28BPt7l2zW/W7xhY6RVjYqwMZSWUMFqEbqCkV/gBjiwzUfiH1ERsgG7g
CpR9IviKhw+tj5nGvnTaDpmqIJMktynG/nVq7yZDJz8dL5d5HXJT66EC1EHYVg6kbcoamdxvyWYr
IdoAMZWvRm7v8ax1ApQNySG3fvHdfit41tx/Y88HzIcJ9ljawO+y6AUUTxPcX+bQITR5QsVT7BSv
2FxrLtY4PryDlJbd9/q7HQf9BHD7RqllM5W9gxwxtYy+rvKhJRYqZMx/GHw/9N4IkadzrBwxND1j
w+2mh6dujfL8G/sv7dNyA4Halyrb2AnzkeoZvSU5lPXzKvMC2e6ppp5SXfU7c7z+hjxUkhVd24lx
Bk5ChWnF1WL3Qie2J1t1OxO677cxeAOovbHP9d4+S93IO1sgVTNf+pWs5kJtkdUIzYA8C+rC9Pic
kcN+ID3oFuVD1Dl3gi20+RSelqj0R91GPBxSs1llPKD0fjhnWZmJwk/D1GF1h1qvwE0hiYSdMYC1
1KNHhiXnwcWH536vmJJVPUHGvw9SjhL2KX9/JsLGLSdCIM67OhowtL+QfiN+qm+X0NUeXfgh98Vb
in/HBYW678j/aU+7gQiQnqzJETydA7AQn6+GVKCzCDuR0l2MiIOMYCapGd1o5/V7JpLiiZnqzSGV
Z1dZIvWegs8Qn36S/MyWg5xLWUBlnuqJjJ5VA5scpA+q+uwt/nn7A7QDVowRsTUtd4gEhQ6eOAh6
gC9PSPsJmEMUX0nLech3sp+N5HGpxxvsnHImLsLGELiaMfz9lL6FNjozdTUcSJezxo4/uuHKKZ1y
M0Gk90fSYVParnnYhhDv0Y9nl9DVLOW6TVMPLMyd/MKyXlk1eeAUYvyHJ7rHL1AAoADqz2Svmjfk
9OO9B9JFAtgZO8IyKY6fjf7SCiKzUPf1/sS3MokkBkG2KXVi29DfPU/rv8m2R8tpxa6t4CQZvHMz
QfYJBLUCmB3BYGprD+YDv6qaHeq2SB6tP8nbnEOOFasOtEV7XbUFJZuYPBbZ+euSV3NYK0aNlKJ1
iDHG05PJNQ/cb1zHEJFISK7D496Vsq3WsnWg6+NitphWITaPQtUce4AXhhHxc1lkjnWb0duWkMJ1
+crJpvPEFEsIV9F1kozwjIOehJrHbwii5NSGSzsEWMGVCJEgP6VBK2M17b02bZ2fayhGj8C5vJXv
RLTmdtDv4pgZf7TYpa+jODe5ytxhK072GZs4A29OEm9DhZx9bxqLxndEQBob7BjNWfAhIpfOQwi1
5sd31u9HD62MKY8YIeQkjXARmUpOjKHXo1BhgfW2LnwcWBfyzf2t90hN9ZQ7+leCk5FVn1Vfum5f
RG6/GN+LN3XNgXepYej2yluDBmgOlrbKchvZsyO2i9bo5KgAAdExJ5zsauZRHW1pSBt+9wd8XfHM
7l9kilX90kD7o19MDAG3RKs8f8kgNedD58q7aPvw3xgvMyckPdOZwtVMLe48A67/IXeHdjRyCnFb
wkJWbuklnUazRkPNKKa+CL29dZcBbqPFgHiv1pnDmYHFMM7DT6eoPiFvyGlsg+YVhBDCaGwIjLmm
4P220yrQUIwqq0ELYK4mJzU1A+JVtaTRhet410kFMDVa7Hqh7tZrRAN3bVKtHQqz9P2+tohavdj/
iVcSmCh6I6KyaqheWxpGa6EOcuwm7MTiAKMnJRQctSK7zsX/Ew1yfwgRSMhUClYB6CaRpIqbXS4W
KD+zu9YsQy+Pgw28U4n+GG6wx3z489AQKC06VcpdXZ4Er4X2Axowq3Gcw0+9UEpX5plH/YveP1sX
0fQd2ncE560nJDiObH4uwmICKCohQqmW5FGEio/tf12EP28TiVWr1YZ8JhTHbMNUS2ayT/6h8jMF
TxN8vPFABiDNvTE+6pv6gWM3bESnaiY9L0Iu6O5TcNu4xhVepIorcARJQr5T+Wj4YHKh7j9bqqKN
6KDsWdmxUR+g+DIBcjK7+Pib8g2Vw/VMbgPBOEPd5I8Pzjuhz6BWTa/Nhd/97ZL0kb5bLnlUx8GB
BonVfC6FrFPRKJvvDd2G1a6DsW/I133hF4bPiG6SKSfzsxbCxwJCpJTavMLjLwfwJo6ircLW0oNk
AFv3Ku8ePUxlw9IsHMTl2OVjLH0p4ikXMkQUz5zBX5ge+ED2a8BxF8g2yMoZC0C2Npo43ddXQXnW
JGeWrrYsDf/UIl5ceHG9xVnMQECPWVgo4P77o4ur3S6POh8q6D2OGYO+vk+G50JguvOgq7hDrbo1
0febQnBnGFD5+ybp/jDjpcvuK3rdQBXuQHUa8GbMjb3Qy2A3r10fcXXQlHKOgpZkYW8eK69fwuqw
84chfLxQQOoBqde4OW+7jl9FEfD8jGGYRnRCfwZ5SVNEU/EXRqkVXYRkHuHWIeVQ5DWUf+yV5Iom
YXrVXSB0qwP0Yu11wRk+N5LOHgwrSLdICTzHsXk+q5Ri29rL1Rk55qUVRVZyYUyRPxzaNhVxKX2J
oNUGZQXcGeYa9QWxLXt5eBqgVh7L+nmXQEKKT7/VnldEVa0gDWC1HPgGO+rRLhO9otgdYCEwOqOo
mtiw4hsXEQyWrLasVUrkPMSFKoAuYrlF8Q0KbzQiiyngGm6ZkPOuDznb5xud6mMi0mG2BxN3i2kz
g2l4BShu4YGOwCE2uOZRP9xYkz3yEvKJP6MwblP7qrblaFlAEfWYow9Q3WEbmVVMfOkfD/ixIt8/
wB3H/hzxZXcKvnQFqrS8USsvePXNvsJFBw9xqH54bV2fJxvKK7xxdS5/xgcJ+TyF39lY22SWxDDp
yuGDUldTfBEKeqbLUYfjBtWoBZ13ksEU/i4FhsrtZmZoyQ6NJ+g1+ilgxgnmmRmF/5FsONeQgFMe
FvEJJSHNv/4MQMjzEy+erF+VmQwPavrn46Spb1Fnf9H1FdMfp2hf30r9c5gX3SQiDPJs1KWNvMUI
IuMz5Amb/N7kO96Wr0dcOMPTrCiSz/syQW4qfoPvojoiy1lya5ogkrllgfCju5GIEbMKJew7PCOj
7B2rTBrkVpom2zdFZ2NlOIBytFtwSQ50AOQrRZZUcIciW76MLuEQaMURoC8lhU9QsMz5NeyTKFAg
ZUH9EWIQGnxjuKhtJp3kEMpCduKFkD+fgmFnFAP37ma2ZudIgtslGtI7NSQxAbhM+ohF4buESVQf
6HAthB9n/QYMoegxeASMnHZ5Umph2WnIbD2bkNAFGCBS5E1zW4djb1j90RKP/o0OXLEzsf+Ezrhl
q0erYGMEbu16Q40V7s7Gu+ZYkBQii0v7h/Xv4ACzjOofBE672+GbPNznrAFz3uUOLhUJKR2n4e5O
+0yG4AKUUBs41Vfs2mSvKL0Z1LjCmcI3w9EP7FRE1wlerywQt7Tk3R6bSz/qSANUdtBaN+nhtG5m
g76I//GBylywLBbL0wX9VtuxEAT6eQfPb2E4wYds9YaBV+B26clibeQrN9+UyQqeC02HCjuCXbAX
TfPuYBPn/xM/E1Fy+5oxrhAWI+gMGSPp2MHEOm1kCHrvPS2omcG42H6ImsnNPhRXSj1wMseKIKyn
6/KQM7oJ8CB1vLyovTEG9HTSzg1URyAEYnAjGTr7V7tomibqx3p+VmVOUxxTDCnTQqsCRuGfck9C
B71f6cwMyHUlQXoGnOq4ZHesDf8fS6eUEAEGNYo9Q7YzULDjMNy20oEHciASFAV2RMRjTI4MYn78
ZVcwRVsUdHoRTp1qxriG7W86ANZig6q+8BOztSH4FYAuUBW9sX/dWJDzgFPqaJ4N6Y0Yb5lHPvwo
9oMovw/96d0mHCdPUwTV5Xm9lApVnJJk/Swgl3fVznd2gBcEHtj+O0uY1nTE7/mLUtLqDKQ1jaC9
tHqww1ud2PDoS3XuRcPD5jtlUXw1AkyI7U3YkrIMPLAvAXw6GVmGheBpd2Qlez7ZjF5sSqjz6ff5
aiM1Ag4nV1PBsSksE7ZAbkmTLLeKhhai24xmfLXIguqjBxyZzOGzBr7xwpWkrydunZ6WDz7vGA0h
oqQbKQPtiMGx2mtKLVw4oWOyNSNfUzdyWW0WYUfKf0jW4ZcybOwP9D4OOxz10X5lbAQa0aw+w8iV
M+1mif8I2Mc2hG2tPFJLKQ8rInOt0nbjzZTOTv1NLqeZRWTvttWI3DwWCBqTTaU3vtN/pdFX0TJm
oYUDx0asfB63ab/9ZXJgtrr2gluP3uRegXvFbDd5tOMNrRyTJZ4tq9FSBPMN/H2Qjgn/ipv6rGg1
BANkKSTRASwBJ5Zc2cv12eS1OlJ9rotZtWEI+waW4cY0xZVTdCsHloJpcIXDExHhnmNOIxcJ+lQ5
qN60u2UjmxwLKZo16VS9hjQR4yxk4C4MVh2glaFyEMH7op63GCLs71np3qNP/Qzpwim/6TmXs/ql
7Iu2tVANUalkbdYPouo0Z9y6yqFyI1tMO3+GdnYUktCCFtR3px61RS/MZmk4twaBdOMwD8A04Nwg
T2zoRnXsS+6EWzuXcqPNgdjxSTsrVJuoGGtQhiTnPGlLGP93MjCGg6qo9ktrmneFeHk2yOD7Vc26
PG+MarG/kWlmhtt6ZXLlusLPUwV9+FJzPbuvqKV39q75JmcB8KUcEaSt98cHafa+rKFdUQVmqvZ1
KhkWef6i8Sokj+dDB7RnIHTq62Ob94MQf57dn4vGhPdB4sIMZva4qXuqiio7mE6OBAmohCxERyIC
eJ+Vvd8PiqH0fOPmSNIW7M6RChLCN2meCgkShh1Ar5oeYoOPeYhtkzUml8h40oKSdHfAanTB2zSG
+dSdETEHxqfRZ+pVC84ULkjuRglkg2TKOHiNOrmRtmdWWc8D813iIN7N5pa+kIxbJyvxcXHbbTCe
MYmSRQtt7b52k1sugpjXClH3FheHtbh/NkzLRucFLbPkZyd5E56qUTm1SncvPs9X2y9BncyWBi4/
45niUWpzcIhENjz1XCtILITzyhPIzDZZAPlo7BJgIN71+v0OxyVLZ4/q2hT0/pDo+GfQ8HwHlOfK
xy5v1Vd+Or+iStrl6u9b9J+lcB3oKieyyHimOGpfMZh1ch7Ui0daVIh+UMYvP8JsaxOBWOtuxyb1
x4xx7PBA43CEhC2xbGckvyCVfQ8/m/ux7ynkHGWCmt8TJs5lmODp724B2VNxCXnhd1NOQYDzcvaw
Ix2L8FNlX/63xv3/1nr+/YD1j6SYjuKdp38TDkT42Eaz5QcboBb1wYxoTNYxk4ObYFAG49TJOo6Y
qU/+N6Y+s14geAJ+K8zOUNB/tPiaarLexz7KmWjPwianj6ILorutYQsmgP4iwJcCXlhbaAmYaFvJ
/ESy9W2sCD2UydDtk3fDBc6eH/3MVYtiPMe9UbSb4iqqZdl8uNFASoYlp9rPTP9X0xYELVZid4iz
1ZIAXSobekNFUFX/Se8mmJEq8MjU8wndvuqZdDWw9orYeFuxu/JlBxlSG3dt3wTp7M1c/IjJWo0c
mNg09YS9dkX3VOhHjhzRHaV71ocpnJ+9+lAd+c0xUS3Z0JM0YLnDxFA9dhHbf/U5aBC9YwTv5ZTD
mLcLpBAwxNc6unxeIvcMEBcA6QyigGG6YPuJNaL4HeodB2WQar+QbDc4QByzhNv4Y9YIZAT3aZO/
TyL1ElB9y109mF9sKKg7ian42PnlU+ACmwgyan5lM+Kz/WXAZSbngWr29dwv+yAbKMegBjkSGuZD
wsAR84JMJ8Vd+LeJ6EHs6R6QoV0a/rQgV7+sXJtxnnp6K0Ncz+Mh+rYWdbb/0XX3jqFk3EhlBvfN
3XnmncpWa27+XMVkTkxj7XhaUDFjlHAUkJ/ggWZba9kKGf5KdwRze6YlreeKdUlBklk/1FqAF6eV
Ip5cOb6fjKXBgSSo1YAF3fR0lwDO5IV44kXepxrLivbQCas0YjL5l5QpfexQTjVev6ofpJZVfPeA
z3N8RD4iEaTZH7ZvmB5geARXsJN28yiWuCGjCVStRn/UvAFPzKdWt4XAi6j7aNHv/uUZcUxDS/7h
qVszrGNTUQ2+yc3LTUTndWSUR1zJRH6MbVKNFCbSRBableoquApAwRcIaig9qckDlEepULF9mORM
yAuSw3cqkKvkBcnaqKHhg6XgG14okD6y0pZtkExiYjtXgrdWyy3lzxbyLWPWmh9RaydgA0vwIIT7
Z4g7w/1ydqANVxmZKcXCqPaVOSAL70VJhVUWbS1/IyHdrt6fWbZ/xQt01iZKx0jsl5GcCsvF3Kmr
SjB8kJi4YeIGhOTxQIUGFjlixnTIlMgSX449iDQSYGMiBLN8le0tBdjsTir1zc92yD9tiOZRLu31
0AFo/NvjaLSIZpgudRc7jpuPual6etx+mZ+NZjw4Jv5oYXCVM+bNyOw1gsGaSRoTTQDowGVIqkG9
3+RkkDOYt5E63epEGWopy7BINMd4ZRtBt/9juEOnU8fZRt0YXVkNhIgWVLC+CxrB2GHCnDD1YfqF
OWEsBnN7dmmEnRD/dW1iQXCB6BTwMvEr09sJ3BJlIecofEd04Fpu3wkWalIxqisnXjEuQnaPe4x3
e6kLMwgmadbFKXz42nZCq3DrViG0KgvMEOBAoPEWi+eleDruOqrVCnqNCK3qrAI6uAXkvkjBqWkl
q2gWrFyFyRk3uaTRHQJJO4f02p0Ue2+RJwiRCieTZwmGJlxxt3nAHi1z2BOu22uPAPWrSniOZFB1
UkE+HVjPPYAEpMMDByFFEL7actCkvOA1oz6qKqKqTS6yCBWpY1x6B/PV/fWDNi6v1I1o1HaRjNTU
jHSwZYdFxHwN++/vDOvuiEszRJYCADBzcmAOswWHRLaKUjmng/j2zOtaIuCHPOnXJEi4enWbuzHh
HwdeTB1McFyCaqTaUHl1YXkkpdQV0NJHuTgeiNAdt1qgw8oS2WYabJKhiTCdzaZB5fIR1jT4oUSN
gLbSOV2BpQhQDU4TCsFy5XuKYTzRJkqXVJo+U1qss1X9dJXcEKppnjpLzJXGfK09TaqHWh1mmgEv
71o106VxzWdr69abhHeL88g45G5ULXo/Fb1uVNZrB2UjHj+8cuu7q2xP5+72qbOEDGMcmXzpMPzr
REfBTYl4TOm/nufwdVHLf9qTDuzUgIz2ytuTMIY+HlZuoYYLw/JiVm3LPJ2ouTzrXTzk/0VUTHVr
sWFduZD+wIBZXyBe8SjaiucSbzQciHFqDmHO6HYV/M8EvWttKXLhE5u1hYmCaWAlmdEsd5reO68A
W1HpU0BBwN+WYmBn/MaDUxNpDU1xnniJyoOzEzF/X49BcqJMWI5H69ydqM/kVSpvVxtA4LkyIzCG
TYcGZgNyjmL/a3vMIMs21GJx/rMt1/TQxAbhP+T0fbmXq9JQiU2ChKK7TmCN8yg/6et1FKEir+iT
vg42dViM/TJWGjoTIzCCOjkZvyYmk/2eH7yoOVy7L5S1Vstu9wFAT61ksOIU5Be7SjKbNz6C9Oe1
biwarK5Ue+zycv0Ff+J7DYlSSJEwq9StvPyOpf9C/L6SyB1d6HDCIqI90jUYOZmhrGrEXJyUtDr2
PyrhbIBaXI2XlTjgG7A5z/WId47H3q3kTNOIx1uml3dgJSIf4fmmXt8sh9eNxM2zOqCDpgJfGQay
YUhT5iJA72oolwBQSg+z07kmx0BqJgXmROsFzdz5WkajVT6R8BlraajYQFMm5WpyRnIRvisBu4F3
gj6k7FN81M3w01CYFbcsGXCuTzwJPfDbTmnSwMRoZPPeqhv0BmrYnuY1LcfhmL9VP7dLZV2Xbj0f
s/+rgZ0PkYqXeoKsUq+I8o17uiOFvWCbuxJngGDddkNdkJH/S1fvhAlXc/GipEu0pRXnD5hMbpMV
6CJj9cV2P4peD4byEzWpvuS9HWwEf56hxBETlNLD5nxgGqyXchfrJeGZPR795t6/KoY3VijiCiKV
GCtsv3P3ShNVg7A5NhsKdrHexXXFMX5CpH3AOskCRjY4pQs7gZp2C6zrF8qyOXG2rNonK485uwgH
srt/QoVp4VXo7Utkq10YBr+RbCIwsdklMd/Q7qHeAhO/lZUzVsjb4Ob8jvL08AMfy7HQ0KN+JY7j
yrGMm+L6Y3it2xueNjhphAdO4ZNb9X0JL2JEyeD8KQNfMs+wgg/T8dw2/51X8r/0CqsPyrP4WmY3
iod2dUFZrJCQmdq9X02rXFGNrlHLAMrYrteIcK3PfcpWaY1o3b1kad8MXAESPA8Fia0Edumw4HML
hjqujWdfmjfxx6QCDeS6j47Cr95adukVuZeQvEpCEb8FHpa9gFqpwaf+nRkolWEpLV91fm+Yoaw9
rl6URnuTZZuONMVki5nRrILdWG2j+/zBQox+S4vG9nufcFCqUw7B5LD3ikayD0QYwYPsOeuyqxmk
cRl0bw8Km33Cx5GUvJ+Hew9jFuNaeXVTv/rI6IQWr53Fsslo1C0vWkDdoZonb0B3fXlYTH9UMcps
BokxfYj/pIX7QScsR8GpJrV2kWQFSbVSFnjovRGvpb2p4M+RUUAbPVpeL9lEmLQ1FvIqpZ86XpGX
ErzRRg7lfbcDHGShoNXyY7HiKWo2/IBe+DJrz3lAEua/eDXE9K80bHFqYrfxZsG2HSTi0ih8Lv6+
WBxtxDGOSu2Dt7uDY1WVYjPxO37MPzzDUFGnywBPK1oFuSFAloRzL2xTzYA2lceA1kRRcuz8h7Um
Yqw2xvIe7315h8XKuAh0fg8DxNV1viBAMtAARrvUMMymrRTnCW2v5GwTmrWfMP/H/8XGAYcy3Uin
4Nx4B5PrxXfDFm6loLbLWbZkvBcjY5zcaha3ikrMsiMDm7lKbtSPspoI4oYzK0SrA4ja73A/0rkN
UuWOBMxrHDArIXC1pAupaCsDtoSnU8A2NxdrqRWosJilFdyS0wwfpDKf9fa3E/0FYNc2ADl8vlAN
g5V/+VzrBQjSccrc8sf3jYmsHbxJm9ibDKJObFAINsNyU1Vu8xamvtgUOwgmkpKDbhDzWBOkkwvj
EVZAra2H1uIlvvyzuCCcUNHtw6Y7ym09fz+UJnHe/AO8BaObgahSGQxVNVb1CJ30Xr/PJXjVodWF
etnPFznIFTTdh/twZMShr5Ww34saFGKooKB7K7IFotPAAn8zb98GT1uRFeHgWoBxOW5kW9sWstBx
CM3Lur3uLPkz9sThWAPls9WuqTlhrycESG+clW1d7EZ20/a701k4FfYi2wd2KZX933U9vD7xFQRm
1GZBrfrrbebugJ/2YZ/HAXJaXxVyqeiOwSv2IKr8n/fi7WhCzYEH/MWpBBv4PTLbrWxkaLa74T9g
0W9TTdzdHI2WRXITSRdTHL3XeQhppB8rta16VGLHCgM19HGLQh0cUhfV3LXrr1fMr0SKvGe9KcPM
6auFCb4taXuEg0KIiF3r53r/REZ6t81vbyYt5s+SP7KeK4Ccbzt1pDkKa0zcvtR1n2MAPeWo8odP
amKre+tgC+sCDwPDX4EmjWwlsxsArTR9KfzGyNNgn+ZHsHzPNS23M7C0uES5j6Fp0UVtFeLwkk4s
NQT58sfDXpDB4xVkDwbe1UFqSVH6Adp3TXa81E5GpqjOn2gNp8ut/mNwj9iQTqG0P6s6PBgUe+A1
LBfRcAgQvby9NCyNdUHA18blowqIUqqzHn07Ze/8gJD7O6COIJ3/50z+/0oBRpMHAJ6toTf2mGHg
AiHx3NfhZTMsH4HGTCI3gTUWBqu/b3nIGpWfem5zQ2JNgZHiEO/UBv83dF3vzYCboVKjXO2ajXKm
8JelO2r5vEpd/JmDt/VJ2criKCZ7fxyLDzcNOYrfAOprZUxVI7PA3wPt61cpzmdX4hYU/ld8sBpw
NW0QXvGOP5md1UGSL2JtuN6d6EE6INAUMtp5Zaxzw+mzH5R7T8SbxV0uxK+JpfFPMv9cUQZe6zlB
fnk2QAdYr7Z0L+eKKE35kMi8ZOVXroABO4+YipFjc9nRCUBvLSylp4IsvSpO1PQGnCglekO73hDC
JayZJFQANgyMZjawncypJ7iNR9okMW5jGMHP7+FtzTgmnWlceu16ugBiji+a6rUYAKrOegr3nebZ
DibO5G79yrc4WHBYKsHzYzJ1c5N2q+UR02+7I27oa4+qeHgCX1CNOq9kGY1KLO0L5NQZquXqZeof
qWHcfsORmGWIxU4DNRCxo/+CjtuQq6FmzLU9wFgP0yYrYe5/3LBMe1Zktdcgj7pdy3t0JGWznDHs
idyttyO1MsWGnlozjeM28ayvv2Qy93thYTwdBpS3RODN7gaKnykAgAzeL1UCEhnpZ1fQFGqUIpw1
Za+udpASIpWWLfuuHJeAo3DFqb83JeBqRA5riGkDKeAy9T0mpmrIdMpa/Nu9WuyqakB7o1iD0aV6
50bDLd1so5WsGA5LQiNaFZDC0jJALJdfMc8g+M70P3HRgqqvFwBS/zjeWEzSBXZJfDHLBIQtgRHG
9r7melS6ddfSaKPcb5C9ihQtWTJXaRdMMEfNi23GEX0mKl9Qkk51fMHP0QQbU7rTJK4Lj0f/PNEM
d488Y62eOlPOgfPQ1MHRL4nsAm9Zi40nUi0FulyOVLvmuQvcfz3yzED+yv2r8qV/epHja1jrMavH
n83Y465LMHSfW4KFFQb318UBSkeQgmF0p7iqSZblRQE6xbcsK1uPNablL8bKo6y8SGpIgz1fOXXr
bs40vAQJlB97WhFmd4m/d+taxWU4DWZOIpuXyG4ArOOxaIR8e/yfqIE1n9LjbH6GjrlvdQVnxsql
XSUyvW4yaV10hlyGZwcYWu512Xaw6RqlIL5SxJZHOB3Duzd84h/M52dCyaUqf6ZIMoydHXYNZpk8
7g8Glg65MuhsbkdiqHUZNdzqT3OJgJ3KsYKVCQWHAGX+M9uC+ewSDN1gZ37c0bWYvjxC1vFYr6iO
8HPwMqYpJqTL3SxsV4196oW7kPKF/rmr0aNct/o/HGAk1tCcfvyDlGjCuB/PJJP0YgFsi+5efVbQ
nNDXNZqypB4qroevKO7riGf2MHo4HBKKhjicVrBi1qQmNp89qCSbCmrt9lN+5gMEszdSp9pZDqQd
ExmYParbwlhgeq/2UsfmfirYAKHSlHQ2YqiXf1rVOKUPue0OpaXP9/rOrShGZw+FV6PzukQpFl+0
y6Mxf8wRHogpdK+SvyhsksoCLuTBMXA+8a3pPidfIFHMfFWXMwvhADaOJM9y8E8a5mIQINSgDDx2
kfBC8zyC5pmkV2ZSYgl0phPwdhE+ufohLRYSIPnKzo2/eqvxe5vpcrrUaJJrURXv7LQNhqpPSLQZ
5IbS/RIe3vhlz49B+UR2KyCDAUMSyDmXZ1v+hyjRqyi/IBcOW8zMaA0oNyN3AuJfwofUE7uiOHkJ
gb5oj84fE6i7QKUThbTHm6VqOovUQb9buTnBjCuQAXst67+qwImrMpyZOBKVNwCqYbAzsmwLt/Jt
Uvo9fq1oBzp/D9bzB30t29B/S+g5T2J9KoFHOUWFaQvMe80mYIru+AmTghoNn3cQIJ8B5WLnsCOZ
URXjMM5ExJuXd/Vd2EAvoM+hWlHcRfxHJn9fhyiFcQTJQ1mastqtV2T5QsflXpjHoZie/yKnQAGT
wuiPOkgOf9qR82pYQwKhZ472WzZmW4WxBL/fGgNMTqg9sZm18Dm9hnzOiKGzvtNgFf9dfbBaLNDi
xvK797PtTEJt4XAH7VWZC1TaPK1p7zJTXxhg3I/0oLdDoaLoP4NoUfeCjvBQeFFIQOMPILdn9XNl
3Ezfw0VQkwOnQPOTE5L7JFYfP9JOiMH4oyNJo9JDXPtPdctbTvl6APouxkGywKyrRZXPOVer9Q47
YCtIoudNoopO+jPgoBo1N1xsf1VG8Wv8Dp3CFNc3/IyAKc80padyyOU3WvlqmTPOCYXrIKlZXds2
SJstV8Dzz8X2hMls5t6GLStj6k5SHsQS8HUeLHBO5YImwWFyS0BSwcjwldcJGDBvY2u3dpP6YrCv
Qivy9atSP7h9RyJAjvTyKVmErYXHVcNv1V2JidCN56gEBWLADLifcLtMkU2PUUkQ+OX7MxZ/ZU/R
N5ZdpNlpEdI6cyfTZTMg7aAW9Ikp3uoGyOWjuUC3FuTTvh/S8Tgvox2szrG/wYaWqDTMtct2KWeU
t+aq4cECYHp4VTG1a4X1muOS218j66pivmLv7Q89lSSwHMWMAGUFPYi8JEPglZ/BvDe0qP9KdR0T
cA+Zh5rbBoFinttjQS6FJGG3PFxFAUAgN/ssF0Ww6YpbnPhQjurGTgEwF2t3leCiSgCNDJRVsaQM
PbBBkc7Ln0wKGLQXrqw6j52CpBThE5x28V8mIeA1gc+rJ1EOkSKJoLH2E9AvW3WRCHZFRi/30vIw
lxi+NMUzsxomb2ldsnsJrL656Icf1kqZpCxkua0brGclvlNeNS8Y6pO3rL8uhFT66Kl2HtDrbCFG
ibM5p9KCDOby5C62EBoNleK+XkiSkyxn2tf8iErntEWk9LBsDOZdeEAFO+n66zu9IQj43Bgvvwck
OisonZTmvuG7dIi20CXPNC69ox5MtZk/U2CjB3wIqPa17xQcNp1kYngXsDKADp4d+noRcHtHw2I4
/XZgesLsw6VJiqIMPSlVZo3L/7Hf3FzWlox2IMTQ9Jhd4HUcvupjO6+PJqWMsy3qcAmWCsFjMAdx
tUYp9aSN6a3lAYJ8y7HgL+fjV8KzAYURAJB08Ncee5lacIaya0uOs+YQYQARkD4CnlPHTCR9Szre
DWnGuKpo2RDnx/BIq/PpnHOaTJIT0F0NhlKYlItt0qU9zx78B8rQ03y5gQRmyJ/eSJCrsTo397jn
9JPECViXFt32Pos4SKBj2QI5asnQAQurVhWM4r01J/5HU6VuPtfnfsfUg9nYfF04FhVoHHPqOr0H
FtAIzqXXXZruG1DD169cSoInUlTXpLitPLxiUjbUrBoagYKnhfz7XBnFGKBn+dpbDkScmDYi2MIA
vJbnyXY/mEErgswQpGv3+5Tm6PYhtuJz6kAclw+nYnytnwG5kt6jPsKh37UEOm49G+0dQFesCLRm
kVZpCU0qYquc0RrdEFpLfCzVytqqMPtArsV/xew7GDKu+BbXS4CkSePd+80IEyCE8LIxWgtJbfRn
xE8m/UE2WssyV7J/wsRmptixdPgu3zkHP3B8fuU0k1mKKutvH6vFf/V9S+4phw4s15BAhwKZa4S/
WF9Gn60UEUwcpslo293XX/wNpdaOlS0+RrmYsEDLOvrzXFGXjS4e5rn9HVqsAbYYmH3NC5TQQdle
IQS2ELfcrqiQeDT/586wzfJ5dRHrb017jCmjvIiMiz1yWo8OzzketPvHzTdgbN48Xfic3mZwrrjC
ZwKsDuobrrs4mhY6aBggiCwSnFCXTCXFZssFkFLq2CAZU91M4M1nNbtus4i0lu3dEHjNsotQFj1i
/LimEKebVihYZqFBAOHGj8rrjQBBdgEtayXRu/fQbJKkW9oeTcfpXnN0Iuwh8ZlkoVASodYcatp3
Y3zaxbGKSkKwcORiirdo8Qp4OaU/N3pcSTCR8gi1hgjchN6cztBoz4a5XrnCGHi6PtjHiwW23FCl
NuCGa0D/jo3q+dpQERfkSUQTnCsp95zm+/MCWRas1tJEJdtqc19ifniuimlQFdRiWXsD1YUqIbT9
mreQfx01RLVAkiZpHOetyQq3lbKyBWH+ORQekRR8FG2LfJ/2/vRPdk2K7kruyIEpW07JBFxAeG8v
pLUl0D1wey4zK8Lk96Cp2KuCGYA7Vqij/tvVdkKhVMY6f1ntRVdNPI+DHQk+ROLThU5TTsAi9F2A
ataIUHuzD3KAV3AhDoWu3ZtNPtHQb0jhPv/Ib0KSJv6HiS89v91ktQ4R1e+W3HQqSRpMxkg0kC5Q
fRSPXwSZxw0MysxuP9rHAsCHpKsZKIVhEWNor9lDddi7yghqdyB4JeTKWT6Lt2CQyxdJyxTmzm2q
mkmjK1vIjmb/hraejTM9Ie3w2q739oSKdvrvulKDBwHXqK90ci8rO1sggy0uI0Ftd8nlxy1WUGpn
EZJPvl0KAc6C+y3At+oy91kicplGnr3XTGRit2fUJ9gFt6GwuaRlzCUMbrAxUURMQcnhcP6xG3rm
r+3XZpYJM3cnq9BIKAQYxLWWshVg1owKjKScw5vUrmwFBiUUfi2QyOYdBoQ/xfB1YjBpCXT1eHMo
2dXZeTROw54tbEPmHd0GjR/SzE7P5KaWkTd0eBCocqbNWIFZkO8tJZ9yvCecRD0cMBzea/BNouC6
YaTHsPbZAqva8M0H53YPDZo2A3m+X358MO9bJvAlvqmJ5cZiILTm2+eUTkxoPMWb9oVP+V4bBwRz
4H16vhs6UFyrHqwrqOiaW9FiG4T2iHCfNVKFzeoXuu2XvNgPPLLbcg9pGkc0/FvwAI4v3/Pz/b+f
Q8bxIDgfILbspn5GjQGxFBheHMHVXzk9tWvJAhwVTJ7/RccvwyyvtBxoXZt0EETcQap9tAY5lNUd
dE2//O6YNDOpkD3419p1wIsmSZzND9DP+ccWOdWPpw2JXS74bN/yb9RqyGENodRHxNsf9JWvA7Ny
YtR5jME0XJ8MtSYU2r99UMRcPBYXh7DSn0u5Apj7LPy2OwnEvgUxwGNxj7Ufeheu0p3ACj+HB4GR
4AjQ0MeLGyVYHlk6y9X38hobAkktp5OZHqopCX5cJWkgab8zKybEQBwpBp0MmOv7axgvcLRrprzi
tU1iMXt/c8e5Z8yUfKeWLMrr+UdQ7ObnALgQpy8E4oWsCb1xrD/v3gJbGZyQX644GLmHfV0woQ34
hxim4U6fVS6L2CN8FRWdBAk/YlWQm01CUUpIgW9LyYQSuqfGAws0afvymyTE/uKxF17K9KNf77iB
pEYJWSFYVMYTMs+NcVQH56eKDD3OYpaRFDk6l91jwOXuSjddPv+ZgJEeooMi1p7WSCpE8c09jQxd
Z5AY2wpia/lqeouvcjeWRath38ABgFE7Nj+fXnyvwif1I6grZW/9CQzK1K4RjFMLn+XAGWKM40UZ
Ap3sOavm0/vXi69F1E43PjuUCuAwCfbkdOrAPgVrn1qqkhDgVNeylUi4NDhldXxZQjCLfqL91LoH
cmfkkwBxjbM4C7W735hP18SO3aZDlGwcjkrgMo+YjpoQ0auTz4xfEwX0p4eu9nmTzsuwOVV4hNPx
JmWWX+Ss8kq3GItj8QCSg/5/cZBQsR71mpAWX909w/ACilwDXfaJsSvDojrYqAiEqXDOILN6Y6a7
DwBm66kVHJolx8tExFCN6NWyIKup6o9TpctilFfJVER92m3eiyquJauiyC14bfDKGxdtxfCsVPnz
8a/lo3Otc5gHSFfxW+ayU6BsbwJy5BD+bJac9NKs0+34mQ3LYNFzv4zPngVVUQhIm76b4AyfvAFJ
NPffPOVmbTxMjnMaIYEq6MXsrzV8nCZgv2rqH/d/mUJ4Tv/cVM86Yh4KHR6W9YauOtTxTPcU7D2W
3laxCA4VBHrjzR+TZ6qUzDJSJr9LlcfYytoWIhmEEkQm0FE1XOL12I4EahuVrrMgMbQraGCkmlNB
nnsIihcyJDKbkFHbyOO/SRx6TOu9NiKPec6jRJNXIPjthaIrIW8A38G54Zz8UC0ggEaaFTqQYf/r
6UDw7sdMYC1s6WyQ1L9bIsBCo9cCTVPlXsho7x6nfXQXdt8/yWF5mLMu3leEx4yxOo6KaXZrSrte
3fF9Qa5jR+rr9LWHuNIrPMUnjKIziZEj3iG/r0cvHBfrXRXim225Ca4vgeJfcJyqG5A3snaTF5hL
wg9RMAAo9WY4S6GHbDJEv2P4z7u/kQlTQh7kWI7p8tuOs/lYPelRsP0Hg3ML5Zc3+bIeqUn+bKui
mf79JldbTDehhzm3acMwxyeXRvmx+mug6XxbK/HT1++hNAhzsd2O5EvP2UuWrRaN7CsTifqZMAR4
diw3HqgX/9N+AwVgKqXXEfzhVOOHmX2ZI7YQ1Q/ZiXHlztIN/9B2YXVcNhKpd7gQkNw9gq9tOPdM
uJjTUCiN1ABwozKleT44HDV5qzV7CTh17TAXJXhlpQMwTcDQ5a+ujJ7teZLKLY3iO4Mf85fZxLbV
RIOiXUIb9GAFRuIJ27CK3ITuqP1rIi24TFOLufG6dfhQJsJKjpYV9ZoTu7Zc5w5qoKVmfzwY3cYT
WpGfjBt41sgC0RK4FFQSRFK/N/RA8dtqOkROGNvrc6vLPF6n3vT5U518kMYMiW8cwrqi1B/HrmLT
eZhqn1R/iF/47Yy6AaOnuwghSnZGBazioEvAW/X3z/qbqPEogOG6bB/EKsg/91ARCCozBlTxTO96
uUKjov2kSn9bBn+wTtyHty/SaNWNg2/ped8SED6YArdkqlUVdNb0Eg0y0ulf/QqVknBGlOSkgM4k
Nd3e4JlAuyGY6/InAZaiRbsiAYYXOAWxFalX4YhrJPEAbDqnoYlOQx7nuiHdoOCdDuF+tmea0dxf
3gJB3Q7y9H3Nh7e1ENjtcVzXpSW0ybf+Htx1sDUtGzN8e+9jxUA8Dj9oRI0Lc7LfAJBl8bJd/SL1
iXNp4FIaFqyiypINkgveb/pS6P86No/wjC2EzPejXJaHunALc/4kFNFH3w0SqigAOOxzGcQwBPLF
ccBJj/mymSvPhZk9hjBljGgUG3gRJG9W1hyN5aD7Ni5ZEm7q1FHMzxoHOoQEZoZxXmYkRm0hdRYu
vimdJnwMHRe4N93HJIBqQBIDVQHoFq6Or5M8SsGLfd4LvT5Ll20qKG7nZZJ8pvIr3afFvhzQSLCu
ahL4/SAJU6GN+XOFgNYdyHZZUARhP0h7AT08/u7o+RGxfnhYyRMMFIBY5lGkT5fDM2okCcv5/XL0
x1c5glix16EbBKyZMw5nWHc0Si9N4tHtFeSInq0Rkcsr6meqVkd41z5/1xTFZGyY27+UGRCMOHZr
nze9XROkPXa0UpXCWbkp5zCXu7piR60/VJwZX9KBRudLQyG9L+yD8uJptEkv4CCzQdDO/Z2Q2FWQ
JL14ubEng4zVjGUEZyne5t2kJdzbt9k7E10tFiypJlutJZxq7SAFqukBedrBb7hX2xsYsdQqYYN2
pAwPjPqsxteVZMCBoQ4T2tONA0rcFSJdHuPkNftD7ahw5M5bYALm919Hkn2RidOs/nwG1m3IZ3Bh
OxM4pxMb1wZPUpBslMCOBFj5NcwPpao3wV6lNv1CHCYS398mewJq8uQkjVr1hPX0KGGDT+FISPQE
LcGDVmVyTygwT1U5pryyLBXqhW6o8IMFtEMa1ALeWVMaWX75D2ECDmFkV0Xhz0kJeNiLy8+TlUcA
in1ews+3+PQCOUaJLZAWtHJWW1203n7P9cnHQSMl/1aedU7R5o277su3O/UxaqxmReCP+ZLSpqoK
EZ0m/VFBIYlLfqN6V5aaOIGOYe67dSl1usbkLZHXEBp7YkeQgv+uWvU5w8jsE+XeklE2vgbVuhkQ
i6MueyKRWA9GpVxm0v2Dm3SmZ7PIcC9Nc0TIEOuBEPakx8gUjLRF5rytrFQ04zCHHq1pZlVd4nF9
ovem3ACFVqSfO30WBlRfUnh3HuCTWXcQnerGfKyixNiH8lqNTTj9y7P6zowpdH0vGu05IOJ++zxW
p2SgD7nhIQ7y+CradWwb+1SgDCdvakiWpycqbUxmo9TsxJz6mcPXICOtHC/JECxG19MJXBXvyDfF
M23DalU9GfG70XDSONbZjvayre5y33UIO+e1mwnfPMKHYekAHkytJYmI+KG39y7MyWHJ1YeSorJS
2GLTFggsBIZiOOZ4jnfjSTC6q+ONiFuRwT7FJjBGeja4ekLNNT2sTbT+gb8TcotInJLSYPGQHqTR
RCrekEJpaW/hPzORA3qYDzw6biTtdQFOhJx4JYZ7y7ChaDHnBER9FKgGkg6LMLO0VAMWKUBlhsdY
zzZiJKTwC6Rh9CJPCLUWDN7j5spobzqiDjv2BkEODHFrSQs6i5G84dpwWFG00eJNXYCgJOk66LFa
hR4+IZZ1zQ4XNvEPEXttcLWxnuB8j2amJxSb5YEMVjDSBxefpgT8/Lgb/YQh2xGKpYesWttRIQdS
rqFSkcf+NEhFqEAIRzNsSVHsVTQ8gVRtt8Znut/PtYKSm7+Si+iarefC9HCBC32XYWBRZVeEDj0D
zj+CXQgN2QL7+M6paHndGyKM3dY2D7mOiVp57kSdTzauM0HX1zDrWMBsXgwkz9vrYibrakn5ZAKY
ZvdbfabFFAEC5Sn29oD1z1VVo2ILfKRVPeNxD59QTevIJRbgs77p4B6370hSY6mXejavnRnJxnEA
uUNIMStcEriGqer0olEXzcA5V+1IExef1II4QMHNR0CLK/Fa49RyAwdyKEd6WmbwfaZ2S5ox5ftW
KSSRFVVrrxVGLn5UlXRSYi9dLzVAFiQqZdY+i8EBM5gL/cD/cU8UsA9ziZIsOwfta8NDJ9DhrJok
kreRfYqvyk7PjtD+WMlptQv3rPHUcd8ZWJHP9FvUIAyZw/vQJ/Q4zexn504JnpNmI12py+2Hq3yk
Ptcrd+ywIU2qZsGzwuJPaQCrSn9gx+S4HO1zZ9MAlboqXVul3eP2RVic8/d8hhVIr8jOEGzRo0zu
jLiWDJoPMHaeAMoRF+gF3YN7Q3lDr+YNgf9D3QjTDaZYUTS9UBjwDGnJVLUZCEsi3iQ6bwLuwMVh
1cpVqNgzbhoITb+o/nl1ZdLXmaTVwXdsXl4BnRNtWo/HgR54WSeGdBhyxGD43fCEYBiyWE+wzQeq
azdTO2U3v8tX4TFaY189CnM21LZ6RY0U3DAK7SKPX+1QAH4dyXZKx2Oq5J2QGbc9gGSXTO/3MxBn
yONRIWZ23sb0y/5+Yr7iU7AD+fFaTcfTgR8JWKuNBYG2HOaDT8Bfwgsi+uEC+5UmDCanTdZiuttg
04Cr1x8dRvqc7lwY5LTGUdy+Pu2Ecog64RFqeaPbLHFs3siGgxxUpOu+IfR4/kpew+L2u6yUEYH/
4XNNgmL7FIi+7RDzUHrOyfEZqUSh4Yx1XhFkXvTqd16bRLy0Z8IQUj856Rt83WJ4N82/n3Z2hGin
OjrkmqupRbWnkSsGbfTXGanTCCc/gpDhFayjBogUEaDDUSDElTLElVIdDiP19W3dLp1E/NqJGMYR
qaDWr4PCJW/AHTgvSmVAIAItU7+9PjwsW7YHTJwZerzwJ6X1GyhN53SARxGfllqEoIK94I/MpDBX
+nbM0Sg22j2rUmGld+4lW0QiFAB6Ha2xemreW54kDI54XWLAk4oJoKQg+C2peIF+/qqyp/uRnEKu
Rtc04WRlU4ZfQcKdYZlO62EVfoSWbmX0MTo+3LRIiPuSSPa9bF0SWZzQoFqlo+5S7oeRtHn7fYCY
eVbR1ytMqtR4C6q2zOlYSBstbaqv9+zau3Lfzo3+Yl754QDegVy4WfgmLggzV/BkpeAn2N1oBJ+6
tZXb5ApXSAWFbs5EY8dcLXugAx4rjQDgPyUOFT0OkDUI7uhXIMsEQ4UHQTNemYkvlnjuhygjPiVy
/7JHZ3Q7vS/2WT+XRGtPu6e+hZm4jRJVKxer6w33Oh1W8l8FV4TNtKewPXI0+vHg3779bHB3Bofd
JS8mtq1/7vGNP7slh6vqEH/tDKAdK+bKFdyRwPCQAiRwt1s+P/vfDNh88k7xBZOe7JWxuAytjJ29
Q9G75vuWxw8h2zxMeis+Hwy+Y+xtya0Q/+U7QuZ9CHSq0UFhXZgK8IaNkOMCK6jsXId1kyD48t53
SjowGciPPHmUc58IZgDjBnR+rqT2UKOGCw+yqJnOfUsTa7UP+Q2WBtD8nicdnqvr7d3kPq8auLRF
VRrXayDQyAV82vPIRgKCH8u4AGCW5kBGekb5EWIT2QRrJXIhh1kj3tJmBC/zY/qoePkRXF2NyWpJ
yDfkhnDmw8+87u/LuHz+mtio0DPNrIvtDm1B0elf077eU3ZV40ZQvo49AeZbVXRjips0v4GdynFs
0aq5f3eGInGb+bnqvchWKo7RvHI6AuiabOhZvuXG32GR3ZHCOFwXcVlG50fIl89r4x8PdkBarDfM
1/TB0U9C1wWT9DRSqw3dv08iE7aTzp3YHjWtSPwanw/AEj79JYjFuvfKPYKwWLPovX/W4syk0fj0
aqUXwhnfrLTpOGrqlsKls8ExcUovQCeCyWWH06drrQDLIG6cmcVMbaA9T2lSrvGGHQJeFsr2bbbF
fFVfgd2lvwGVo8ZIKhjj8KplUfXH/NmwnUCSDUklbGB6bp8YSdIxSqjbudVjMFLJpV/sCCli9CNZ
rJ8sbjetVO73k8+k7hB1ceT+gJ4pJAiFhD9zpHmNMgg5UcBJPIoA+Kmdx/YNbsfdSJMG0/dqUkxr
aiOW2PWSBwByanrYDxdilX1jBGTm25FHbjO1Op+4SuxIToJXUYF8T6UOfQSUeR+QOVbJHBfaaUdn
FFCBb7jB142LkwZi5JOOuLJgPt4Za9s/bdLKxpKatyMmIJKrLWf3VTvUTIA6/s8XRznixQuOL8Io
MiW7lRGqQlCeYpM1WH0iPDUCgWHAOGZjd3wSdG8oqtp89vrGsW23usAqwYi5HGzHs1VBlKWTg8Ov
PKmm4lteH7CrgzX2LpHM2EeyGjg0d9CnpCYaS/kwt3T3+gCshtLKC8/ztOxP5WsM4/1IK5RV4/Qi
TJQL7BDU67qFjMCrmQHJt5Gl9pQIX3q+DMeTENQE00XHH0l30skebi+cg44Q0Y72Do5gLsGKo/wh
THc0FrjBu8DU+GzpD1bH5oxSUpclvCvat4M4bl/JHGGTthb3LRiT0tUJwzFkD3gsI77fgJwQDT8f
dubq4t77GBOdqM+kabaCmcG/39WmSxxWKrXfWbLzcxDfmlpJaYFqyJ2b+V1K+M0dm9qk7wbk3ELa
8Xe2VNFEyZRAIByR3GyBx2jEBBtsYsKdv6Zb3O4626G59rJcl07qYNCRlVFo5aLwY+rPB4Ri0m0v
OE5Nns/PNcvUydPIG91ykQ/l84og1jRc8GSM3CPYWA9NdW4mW4tV8QZIm+JFvynLNQZfRNxTxV28
iiT93zBVrAke9Ewq1lDo9aTj/D/zy4NfxKXKuWe5W50zodM21XkCQlmY1kYE04zYWU1h/C/TW5ur
bBUudfrrUC0Bz7M5OmVqKH5N5xrEWvE+GIvZwNJSfb2GM0ViFFUmpZg1tO1O0vsmSKWRf7SQiwNL
DUa45xDY485MVP4PmCMfZKox/y71ELgyu2A/tZoaBFzLx+GxDxWNhv0EsiUDR2jbNGWz9XAlH6WJ
LgbixDjtgkclN0C17yhS3J38heiZCteZJk1ddIW0lsiC4FvNwfzjGABMbVZtF0UNDQgV/t9moVjL
fy4WdXIznCA2r4QOKFxCzyCnmQdHJPaQLen+ro0IQscQ4ORHoQvZqaq921mtnAvqPoy8SAb77hzS
bNUM1dWJA5l77NcdD/uRXhEi6h230qy2lyFqoMW+Yr+LZ567MYD1JYBD1Cskgt6bZYE7DWbKlTx+
sXxpdMyDbxUhvEr1mIKorc3xqG9lYRhbymOlZU0TWXQzcOgOhFs4gnJDc/1HuCpK9cyInVU1UIXV
pGjEItbEeFWq98nLu5HOd6ZRf//0YxH9hejlqqZ44/3lqqxTOwvgjokvQGXJc41TRqM5Lf6PR8eC
IBuHbkSqYmM5jQC0RKaeNF7A1H4CJv9CPIj9OzhIEow8lstfodKufz0MAhNbOttUSRwkRfwDBsSm
MxZpn/ashG0BWw66jsyH1YRVIZLEeahWVGXxElAbrRiYo3XPm16tpXHNBFz7JWTecObPkpfYoahq
2YXwPAERJ6dvI0FpAYCMydnbuPR1w4+qUZtjDCNcDbLs3Q4O+WKihgOns0N0qaSE4xv81OoMZOdQ
BdZeqG7vxgZLHVtwEmLwER9rh+zjlQ01KHA6K85kyhxHyg0MoDoOga3x52NTvJba8F/FkUIvOYgx
mboO8JuZr8dpPKUKSVXYcH3+yYMG7dMr8nqYv0FFkqAEMYxzo7jZ04QQFbjORLCqq8ixUypCoo5y
dLT4KP+xufUZtHTpXC/03kG7zZ8oqeSVzArFUAh9SOsjSnK5OSfpkK9piG4Y0REwWS/HEoxdRBEh
tEb2R2xHuQ0y2aHQfomtPa0aitqcfNe+ApiKU3ZBdAJ83yAwQ72GkX0EzMFdVIpgP6b5722/d6qx
kTtUWlflF5T9qTZNAsh2/xv6lUJ9hq5A3tHSUuK5wSvmRaAuSTuinPoz3Yltl735tTD+Nz42O5XE
cPyC3b2t+GG6JV/OUD9yTGO4wVVck8lRYyCkCX20sFuROdf/dvPnkE0gqDOZy1tkXkZx5Vnjswld
N6NmZ3HK5r19K2gbibLvLtkRrK1c2/nR0hj6C6lMih9uKfK4BexcEGMFQmy0K3OjcuTWtSm0CdRk
vlVGC2Xyu0sEumSKpp77fERb5Xay7oWmmh1eXT4pfX6XJyipvOEaHc1fdtE2lsXNrHdwzI0SU3fb
CX7dvY2tbfYkxuDxxqx2sHs0eSXscm/FVer75TablUw9Y/yNzGXdDFwHAdE/JgTOrFwqm2sYDDey
610+eUCxMTPf4xW5kZw2hhZ9HxdZYsbGnn6Z9E1xyzGBxaiwCqyrFayTLdRooP/7I2TjsZhWykDT
tz+oX5aIO++p3BWxhBoiKp90bv3Yy8FvGRhA0Kj6c0BJOQV1FIwriJWmv9TWxv2FLSvUQfYcukvp
hn0fphkUJaXyTMVJA9wzkFyTRo6w6n7wSA5dpG3nfVWdxEaLR+Kkg5dnmXTqEV30CxFRkVyrSbvC
j36lM/WBOqFc7Za2fy7LFNCfVzQz+uQWvGOk1r8/ntEzfG1zRpGasLOD0ER7ARXmYExwCz0sp9he
RLjMv5amP4lmbQ0mK0CXDIyuI/P3VAZEQQAojDWFIlXqVw6vV1iCqBkQCcLLqIdlgK9kLrTPH9Ua
CneS+WmkYPF7UPQqqYHrMHQ9P4kJPKvviY2WW+LMfrdhn0bOTyBvN8srpe2ZvNxBDSyTY6EJ7+vY
QxVd0OND6Lm03s95d+EoUxH6pmgx8FFciUTt/DKjIejTYALxxTv4DyUMXfBFEsZ4WLal3z13Vzlc
rKGDSZWuIeIg0Yhxg2IsQSWRzYSxQWqFblgksQFUg5XIBVoL3FrSysThH5bGQvFiFf1pGRRi/aAF
12DVwqrn1DfZyc1vM0clmXs7JYeVMrO6qMRLcIhs+7epjX0DNNbU5I6dNplicZzZUJK/2uR2l/GI
eZdXdEz5aRTeMBz2PuDyGYUJCKaD30z3zaeIca802hQbRVtUITYWufhcUjU+3+VdVZUoUa2auS3H
I+abZFA6HaQoLNVVYjMAORVDJbIRfa/rTjCMfBlmukrofnvniYZwWgJI9YfZOf9c1NvAEj4DbfIR
9+yNxCO66zNidhiXutyLqdAVGOmqreN4AMCAmqbDEnjhZxH0yrNl8HZUrpH54TP1khx5wmK2TICE
Q4Ujz+tLJA8JcP6WZqEN92Ouf7TFE86DOYtSUz8tyCCcd74hBXMQBGDiR2ixNfbrPcd8LdlmzRXK
DbtNrxgGvGDykPxEegR3u11S7iUI7rMLsOTJvi9T9w4gBn0KJSO2FezjwVgL7QG0LBtd3H7Wz0aJ
VMn9E+f0LUG5TlzC6/69UrtqR3BwZZCkfZiG5KX6XeaZYtwuA9ZNe9EzTvCZKUteq0734hzDf5Il
T0i+pEH+JgMfP1pCHSbtDal8u7bF7HX+ErG1265jAV1XjEXbvfbogzeces6re09ULgb3WeXGUCHN
jlYJXqoXrARdkuN3M9Ex5PaRKdnxkylov8lPZ9GR+Qh5WkRJhVJ4qvjDkY7IbDN6E/Ri23Oi9JGT
FdQwXQ0rPNx4HRQHabKc+IDR8XnP/4vZCwbAgWBllyvbgxftlfnZmI6sgRdRaidIxy0HBLFkyrBC
q/mjctg44iQsF8Zo3OWBSNKdTEfyQiK91A19tZWBFKItSaNe7X/3bdy+8mxwwwT+g+iYxJZh17sc
rJF9Ufam0XBItFZ/c6vXWOQt5iUwunCBR6qzKEpfXmoa/qsEww0RkI1cg2kSB5qeZoaFHD1dwE8j
XNaJju8UOWcppG5LDXqP3bkLxT+Q89BJfWDqq7+46mbAlWiWwzvfM+1sxM06MDoCMepBxAsQNygq
zxskZW+CIYpRPmHLiT0R6iVGVlGf+wz7gb6oTStuj4rc1Jzr8MIdlsdZyXxpSVI+Q45qPQYb8M3z
sN68nxijMi9CpSXs10Ktmabe/ffAcm1mjrQpNhv672kbTkwzOUwaMxl0ZbEQZxN5S9VI6GiIkGIX
S+Rgr99B5X3r3ZvKT0nrI3RoriUwpl3wh7BriS81z4V0IgWcb1IGVUU6zYaZIJ/FPDxVWxoH+xtW
e1sm6FHXf9J2YhNeiQxUEmTmmRqDYluGoD+TvlHzPgQDs8P0UuJ/IYrr2mia8s+397+Rgmsv46D7
Ok8f95H3S8iUJZIdR5StZ93a0T+J2esw2J3w6/FvUJrLz9jLc/nlnaDXRSC0ahbFh3J1xfSnyj4j
fqLO8YPPYMJi9C7ExwxX7aRUYnIFrlfVowsOtTMCumNQyaGD+nCXhaVwt+31KVbeNpyjSvL1CQ+4
FB3FAjN+OZ7Q1wvgzRLmboiOUAOWpOT8bS4ZS23oCyuzPnZ2DOpSXK3IWfo3epmjBn0G6nyKuM/B
tlBWkSINBMUZvxm6X7KDL9cKBO1CYX3W8NdaXKSNMFSnYR3lVtnir2LHa/6+pRqi6SEL8yU1MXtN
P2kgCXNs7eLMWQCq+E393jgNa7Knf1/Ms3vLRO7q8s7cuoJQJVZQ4fKYQrzb4R8Tu1NgU68zNhff
auISpuUiG4PUVHNd9AhWmYJxKv6mS1is+USZTiaIMhE3OVd2MeDTsPqJB5stw2RAAsOEa++gkWYS
pUZMQxdM8/4beOMDeEteA00K+TppI0giea3gpA31Y1CBezt5RKmpBwyv9Q9Ye3IurXaBhw2FrNA3
+hxfTDVJFjnwqdSS1CRj/DKVi6zNPO17MefWLMZFISMcqyiozhqSB4OrL2mqI1myj+4wVVeHBhTJ
tX7t2Cky7kh8bwUvumJfPAlW3qVgkJj+XDDQe/F53obgHU+qEr36MUPfPC4PwPEK8bi8hhKpjARW
IWHqifHTEudDeq2Je/b4/dZxvkz2hp/gY2LJOcim9r9JI+BRcKZOvuspb2GF1gafycG1kr+Vnywr
b0O/06KnCHffxqiYa6IExfKHfHeLhJdxlWeZuwmf65W43KljMaX9zFjs5517BabfrrBOEFBKjih1
xp0uZQrksiDMo4PNaSBkcbLVl1VlO4zFmRMcELz1MFWjEEzFCedOx1p00zHApskF6ia3uP3kr477
oz+iBL5XhlPomaO1r49hSmvF8uJbeIl8+QSMCsppQSFb5L1oV2VTh5Itk2pl9JnKesBxSjjyb25T
lmUhthfT8fv+GjtfpFiiQw9t5vL6JWar7Ag/OJXplr2LoQT8brAEh/w8ZHc06GXkhnJ/iH2bN2YE
LiEoddJUpBXgLiy6jw/Kv90CU3vfDw0Z90b6DinPKz+8meuN/LUULnUeBzIMTFkC6IpEQPUM8zDh
2sG17ixN8oSRgOI3joJjVaC6B+fT5JyIhsD8NxXUSUfbKZtBKKHLyGLl9MMCLWa0zNgVBScpXskH
bR6+iWEpPk99IaSsbHz2ZU0YqOZmVSs65mg9HupHzhxW67hmEJC7Tom9irr+xMJ9Q7FZZvmV8VN8
uUQVoVUGK6rS7b/vpPQp3kxrxWHUYrwDAJnE+waEZHq0+1Abiys1M/yySamXBDzETT7SGopZHEwA
KlCmwBVJnakzy0suvw5tFylcWNiQP/uB3PfVnBtM1G3IfsTDAJu0rBqaBf4Xt9+FP8KdGFVNKFIs
7Pz+2vx98ALv6cUJh6gJSdxnX+r6qSbNiHaP96ESaW8OcCDpJsMYLV5+LsPJ8ZgZSHJcuhrkdtM3
cxD4/MZy8pCeOQ32RJg0yYk3W5EgXu1ldzl9vTTUV5+lWOwba/TazLuI3aoHHky6lXylvf9RzTW0
Yfm6J4EwBhBqG1vlCFlS/4zgLGtuBu4Wp8e45ib7pRUg+RTcTksLSjq6k/1xoImYZIjuagXL8U9J
96IxPeVeCnLJgRlE2X2H6u3TbPUxAcxuNao3T/ePyRHg+mxUSRD5vyo0Yt1uoi1rRysf411gKHJk
ouhqz9Ixh434D98nAsPUVk26PQm4rUPzdNgnGKFdkXPXw7kaccGlr1PKst50e8bLiIg8AndRFP2+
4gTxaZr9isXFXrAwLheRr9pP+J3pV7f03CUV3YEZ2Y2b3wzhiN20hb2kCNPxMGRksOneTp+8cQc8
uIOGR5Z4/daULOQcJ0ojPd+OjsSEPjh8+4gEoFbYfpDcPaO0AqeC00ZaB8ZxSdo0iUuVG4vEsq11
Q9V0A6mYQdP88CjQXAZy61hq7lzNQin07zTdvIWL3OQFz4Dq56VghummfhufWvHsOChpRiVTVqpW
RQ6Fsmq8ZdHdTojlCac9io1Dcc5bXVeg3unzSBB2NoMoKvt5eiieH3fccnZc6jp2PTw/B3GSOd1X
5qFnPCamai0ljfHQGBiEc9Ex46Cpi2nsqwBTvt+3CH7d8q7QVFTumsAoTGl4ZT6/vZQbcaGJeUue
wJwpuPAmi9cK59V3FVezfZG2NRVuDUWAXAqKflHc8V6b2EatJjR+4nPGR05oOCYB5AR4lQ6h6GgZ
aszqvz90It5WikuL9p8Hdb3Z0GTqDS0vHBoI8G46KQjVya3EZKnL7zfQp/kOUmV/s5AJQA0VUmjQ
wAXhbccVtG64g8eicH+p5U0Ktm3+jmmRM+vIZRvRWpQx4Z4WsDOLWAAChwwDOEszz3sMRh/dHAEW
1MLUcn6mFsCBRzNDYITY6c8mUrp4DectNfwu4wh7VCWhU3JGmw/EOJ3A3EuQoQZk0AYV1dkwvl6o
P3XAOCfA26HUp5+HYbdsfDm1gAllcTBrVp/SNuJKgC0jB1PCtviuZCw7SqrPud8vvdje4ZmdQfHC
Ll+GKiSKfah/+EFkFP5x9wkUEIPknFJgDbjQP/5qQGj4Iwl5QE81uvqZV3L+gcmNdnBkvfnx8Oyx
nTlEQpcgR6AxLpb68b1wLq8jNSnGs5xH1RclmX3527PgIRJejzFdI9nkoZ5gDKTjCekFH21iSS2N
Vr4UNYecCaM7Ell6uVfPhadfkfh7oP869HdzKca3A1y4hWeVoEUshCmka57APhjMfEBU4iMZ7irl
xRFNQTcyoxftFhhq2QUrkVH0JzoSkq/XOl0K51M4vWngrHOSU0zN7CXYBEc3+Trz4/Wgo+0j34D7
ocQG/EefeT3c2hZOvjKGrEH97XzM524PyqZuALZ66TV3nE5U0OFNzdmXw0WH8Tn22j6EYqpbMS5d
97kZU1j+cvh9H+8QOl8SxUz3sqNen6fAeCu9u8C3MZh6R+Ab18yKIR01/SvF7aAgTB6zitthM3+x
aX5C9rVucdsThZ2yqKRDM/mS74NO67ms3+iDmQ7Jkmj6EaO6hj7RkSWU9PVmgvPxrbjWhcHjcHK2
ipSUWSZsog1EjOj8p1TljwiiDqFqqGlN5AqTLtlnmLcqEgLlbWXBjGwZ0GF1AUkT618JS7fcs8Xc
0la7TeixYDVNV2Ag7KyGHappJyJoaLylFp9an8nly80Fnt1YE1dOOIKpjY1E6k5HvbYHOT5QL2rT
bAH2m+JucZEtBq3I5WAvEQEMVLHUg+j6k0xAKkczl4jS03JYcOMJP4BQKyUcn+cpJRpJ4xSnEc2B
fBB86b7fjUW8wYq4cgKYO9ZAZ0bxk5gxthlSyRbQZHitPMR15ruRtwZ5nUSa8Ax/jPbuf97iyyvy
EVY86FDJ2XfyaytPUpdhtO5e7w4HufG9tCpwDE+v1zmdrWJQeevemZOXTFAa8KJO+C2ad8hChkZQ
lloLQul8jPEYiw4YwDCpsZd+JvVpVtOLlT0Sqqhqr3vKZMKK6N/eN9uPOSp9uIULZVPPgMVWwYtj
B0mUkgRV7IktkdVeiXwZXLbEgu57cuakRiGji1DxLwlfaPDegJffhaYwYbaQlvqjlVG52wCcvOqz
vrM/hFf9NRI8NZSzWXXUKCtW3sroCSRIVIyOhww/o7WxcaGn1FIr0pAxs3HY/ZVidM58DIn/5CTP
fMcDdIXDnEMLLdPNG5AEY9mgOkz7uno8GtD/6H+N68+qvP6P9NLtJzmzGJw6k4MQpjuDKWYGIIlD
4yNSyH8MIx1KQ06XrRlTPe43to7rDlG2MZEP0/+FriyuiWgt+jr7yjmeLZDCNbvm6IFYYsnDe7V1
hLUQ0vDF39/DxMFfHBuvuuQWVTFUXZPOLBtQ7Gb9waeaWfRMqzlwu5HpHwpPprRvP3BZBB/m9Kxe
Fo/k1VvtOrO/eCElEywtwA9nSRVk24iuCA69Zw9Oa+p/e2HMktd8rQIPYtg8yTBtcsTZjpckBkaM
IoY/06jaQnSZ05Io0GblFAVjV1ROCp3EzRicERMO5Ssdst9TXMS9v/oGB5WCYfxvdy44wUuxE2VR
H42OA84dEcxdojwDFNuzI8zfNU0TpH4Zq7ae9691/nJvqnZ13dXA53LKPf67uWO/xhe6t628N3XK
Cu3Qea9vb15Q61R6OWtsfLNk+1uTMo38VqcHMj0rjnPNydeCDAyWc3exTgnVokDfsGKf5zuT2dMn
9jHrvafKZpEtZU3bQImDbLodRAMCNvXwl6gguKYBpUY+DpZvyB0QSctp3Zf3FE/6twcScI+DWL1k
F/KoSvOxdkLNnabqLSfZlfC3W6tW1RnxJg1oGU0gOTiWnjAXhDMVCs3DBgk2rkuvhkBcrATuhil3
wCoFWXSVUdVINjZy6xL2kKee0a1BAa0YFZhggBlIhreVw2kByIlLLel1s5QG7UT4/Zl2rsW6iuBy
WoeTC9KrII8MyRN/krn0sTQn3fPXNEp62Q4A1I/PRrCDpn3z454jdD2V//bzvAD6xtbNHvt2gvpT
HgdrI0osik/FuwXfa2nf2hLtxQKHJnxMgBmgloQC4gjH3jgF0Ban8cv4/dHf88l2XX1EzFRMDiFY
OUe53xYsEgx7uLF4gdik9yXz7m+bHoKWT04pWtpnhKssaO39pZDxL6uNYZXaJUujcczO5k0pWalx
6EC6/NjE4ImLx3CksUyuDzVjAQWRGOLLHmE2cKRgt0naQYsGS13HT7HEmz9UJWej8HCW3JMmBHwV
Z96heKrUhW3mRpa8W/c4Qn++3hpq7ODDIywad77grlR5pYbuSlfpqD9BaH4z/r1S5JsLS/iDeKpg
i6jQ6aNCwb2GI2EYhSX7cwCtC64iLeiDQ6YBpc2vmG0HRExbIIzCimBYKaVBUZa75B4ropuLYN5Y
qqGlflLDZoqkOyQ2a/DWBGt61M8Jc3O3GN1fVKB+2YECS99zTvRLjwgHYOWN7UWd26oCjwob5/wU
qn8qpxkLMN7VgcvgD2ws/DSYD1VEZCxJYSPzX73e0xXpTmgukSrIIuLhx1Cw3fj7bbxTTWxPqQKw
fZDZw2sQlXdoQqGivx28CXSNxzzgDNWeAq7+Sf1X2b95QJ8y1XpOsbiepoWEVT+EApjDnSZMYCfS
z+jEmuolN4MZXwO3yEIWZtW0MpDzWlPCzVFO5CBk1Ko7g1phCtK44YDONKGCaOE1orE/Xjj1BXPQ
TCBE3T0CeBUosf2Uz5+37RiEeFYegEJFGQ8lqmr9csAJSp2Z1/d/knDsk4UeiwzPZkjY53WzVMdw
QXX1IzODGTi1GAlgrqsKKjgyIQdArHSVT4uULgwSWzqZve8OtJO4KmuoxCREJ3pQaL1UE9DM/LZ+
N3FaFTScmNDUghn5N4N4XZHz7KjjdTJ++fafRgVQDnZC9TRNoOFXC4yPy3531441fz3QOB+vZKAV
Fhlhkt9OYEIqUM3UMDPuKE/V5fsUnL1KCy7JWkwq0NwX1M0y+3pneI0C9BFiTl76j3OcXpKp0b1+
SjH6eKxqc092d0AKcr1S1alKL0X+/aimhZOC6qHhG8EIG+xSg4MnYIuAMUKkgIIjjJD9J+u0NLVw
Zaaf2eMb0RxocFtfRqU8SDKuqnpJkFZxfhTcte+/gtC+QDdhGLbLK2XScyqlgH7Gl+Nsy0FIh367
iGgVBCaJqYB64Vkry4C27AOcJw1uwAhBQ07RMUHTtLnn2AhTr9vcB69TZ/5VD7NZ460V9uEnZyc3
61Izkh0tZa9koJXZv/UiMzSCH4O01/Em2inFFi+ya+iO8pLQRzmgJ50VN5zHO178o5s/WbTeykv9
6lyUDNiGBru/Krd+rLihFF8sK/oDHDscI0aRWOH3NujBdzn0ssR6TKnjNsyA68qEeE4zxec4YoD8
7uhLbxy/NXHiZcdCg0A990xU0GZOu8UpbEcmQHuVh+/oECguy0kfO8fv/uSSlIps8AJIrJ5M1trY
HouOEdjgqfx4dWmlFKCzJd0jZFK7y/X7mwPi44iWzS+kRG8E7CW01q3/VZ90ntuKEntQrp84o1QC
A8B1KWIhdMGC2SBLSvmoqWGCu3e9Lz2vA8GGE0j2EErGQGQ9C281kQa8ZLPCWAu59KrjLSNy8BhJ
GAMddG1zVEABMe46B1l7kpysiu1PbON9QdneCJFOxCr1LDrRe7Nna1cdvBuAYcprxPlyo+nAjUn+
w1ZuW6cvQNadwZoexql8uiZzW1cYa9vM82UvDrYrvUhZTuF7mWGy5f3DY4uESn4aB2Dwx9ViLMML
CJdTtPjp+IOeNuaHg6i01ediERuy9Qry7Ocl+REfN2/XzWcQhqZauLNICEimT6EAEbOErxs0RhZi
j9w06iEMuN0TucSEgpFzT14w91tyfuPAs7BlXuKqLdEoLe3KALulg0fZuLGWei2U1rD6I/muJo9K
e78GCSpC9ac1BgEnc67EDDM9dOx4PCfo6YKHR2fZjP2MTw++EGxag/Lx4UO2P0PL7/8jtSCgdKh6
h+7WQyp7n2JY6eJERn37O6oSY8HrmtZ8dV13sFiSRH4qNqMJRxbA2SxjZBlG0cfhoIpnPVKibBt9
7OadHBAynmGB995B0TTjgXjJdtlueTwFmzurN6g7UHpY/GCHaKToKAK0ZqywGjCgeH/tcTSOUEh8
SECy5jdLwovn9bi+PvCzpPpLRWzIHC35W09iFlXj1TmYVGvB/6BUminXKVnzMUgb+A9lMrmeuJHN
3JXsqR9b/TdP0iAEtNjawFUX/pWHwCicd+zZaYnO8IkpTmc2ULh9IBiAsCLly8yIVCAliKRayNGv
BClpyaZYKW4QLzaDccXuy90f8IokWXtUUoLkoR0CX2y1Ucw6yXmbhglq7ij+cMoOelbXlNRtMEiI
Ri/y6yrMkABMFiimd2j+jPWOFZBh1f4kv7Hy9W4B5TLy5tlpMNJgkErlVVTXA86bR1+E4gqDcieC
+fyS/Gm6Udiw/JaYdA1/BcXF6CsxKAnL58QJQ7OFMsS5NG4STkNEFf4NP/pwE3JqkM8J9p4vgZy4
qOoSP/ZYjN4baHWSqh4qM03QkVvwzPZadyJGzYqh+1MVPl68S8UhC5MARas0p4EiPTxxJ701Io3d
nVFl4b3LNyqwqpEAouG6LfPQFfI11lV25e8R1K9L91hZm7wP9EuT1v/rz9YLgZx2jeg27xXMA83x
RpAmrdFKMBytaoakPOfZHxL3AsPnFJmL2ctrbrbgTtXHk3GSU/0mKQbF2fAJeIqpUv0yTDgHqm3B
ANlGIhOQjoic91r37NrMV079SKOUk7/QrzHMcQTZ3EHOqJp/svSP634zhKV3Kf9OFn22GJGyODxW
P23CYSBTfcv76aMYbYv9/VRFN3venMZ9UaQ3uJXzTJK0yZ8wNouCXTL/zm0BrfZNxiy4PZTm8Y8o
JZSR10DvEyPz3TNpXFCsbzok58MtWl3SfaR2g/uEY2/tlFHfXNpmGokZVxLbdu+Qq0e77JBTH+bO
XkKcOzxAdz+5/e0gUxWDnuKZYSHI+ytW3A31gcQz5ca65f97MN7J5QLQTdLdq3/aR/Yb0/Ekt4s2
n7Y5SSBMWOULhmNI3sWFG759PGFvVMJCkXMWCEbnha1898ivYd8RL81RYOn/SVtrEj/Ioef8tsYL
k5f3Ncw3x/4UzYdlkZigMbJDqsdRgEGqnf3b1WA+uPq7Umr+Bw5X+PFVZ8PP+Y6oQ1i/BUiKVGzT
YLhgVXTESdF3IBExFeMlWPRzs0sp7xvoLXgKQSYK7u5S4ojDpN68olX6FSHWwQTtBiQVxYT9alNC
hAyzi72tIiVeScAJ3BI49zavF/I0RNmj+ylTn0sLZQFQgQPnaTQK6vdOn1O1HULV3fDg5ge3PeeH
x8sPcO9+2ihHJqjjMsy0caRD6Vlm863R+DFBAyUJHJK1DQc3v5wgwDWCNNkfrxBz7JcrffSgyUWx
KKV1BGB04g48832pwYnebTf9mx22WmHzuvbayuKbJub37AdOCD/grqtvdZlzvA/U9SsHlQofGGtP
Q8g3ASOcKJYQFYftL2Y8UhzpEGB4Q2G3loY3PJKPYyHoTGRxrEgJFusGYhmFVOr4EXJZcU/G9LE5
OclxgnrcaMcutmbT2VdTLEdudexO3qZuCRLVJyG6FUxrdvfS2C5u8OxyCMNBDui+rgFLGBrsfx4y
tVHpHyHIpqCLlSw6FKTKbRof9utLLLXfMYwpcaXp+hHPyWMZyHyK1s1EoMmoyig2qWIZ9TCi90M7
i1KNQVGvSsG6b4yqlZ3ooHg7gPDI4UXXUgAvX77mo1hNl+ao8LA1aViprEtRph/UcaX9RC2NmKAo
d9jiNqUxxzJouux1Og+pGnXSOp4km2wGCBGlxhYelEjHtM2D8PcJrBhuLpPWbcJ3wDpZbKP+0MjK
54NIj8X0pPlBPgFevO6vPWjwFohu6d3OCu1tXmZDOe/yT2ZQJyAwgz6QS53D24ez/CKNjbapU1ML
nKkISS2UwqOWoHNQmV+moMVZeLn10WzHSlZW+yUcHId1kaxGLj1zdT9WgpfupLa1I7GEQe8wcotR
2/tMaZchR84fTnPyA8yET+TK0h595QVv3g0VHz5al/kmyIfHebC3Mzrz4r4YFKKo2695ASS5WE51
rM5HkvZ1VtlrSLbUhudmwMp40fxZZnEyfKBRm/GseB8EtR6UhioI3HAgisNL1H/qumqjxpoXRQ2b
aGCBhP2AkM70WLx57pwdaDt7XXb2dsYCOqcUQo+qSG3haYwJaGoGk8SIE/Jd6A7Q1gnBfPbAr0NW
hF40GGDXQ3Mf3hy0M13zazdUhyo1Oyba533llpam99Tt3Ddd8NS34CEJzQt2+zWvRwW6yRPWoaX5
Hf/uVaq760ZWlP2ES4Uj49ZMvUesViVxkcrKSkEze303KdhSKB5ot6aYgOjLi9j5nL79rjA8AkJu
9Kh+PzOyg+jfWydhNwVJ7oLOaSXn05PR/MdYe0g/wQbBAC8YnCLKotO3Y67QCh6fUyxu1rukw8dJ
2OcRspKUxcVP4dOnv4Z4nwYBi593zNHJDegF/fLKW4Ui3wKpTTpQN6u49MymElsU5u99NIOKi5Vr
mfgasWTfWKnNG1VDARJJVEVGSP6LgL5Mvsbb7kWd5PLOT2SrfiHUb594yLsFP9HP/uMorBnGan9h
dBVWCZbq2oSXrOLAA9c7R5untVaJX31SkBhSx1Rf+ik0UBNG/xdY1m6HcmhzwlfarwdN0mZHiJmI
3jH1Tzd6e28xZ51fEg7WdA8jwq0+NBPCCEkNijAB22BA+H+Je1y34n9OJza2Le3WrEvcMYlhFkNY
FvrYIJyvjPeyev62jrxQ8CtSMWM1Z08JhN8AV+9RdhUIUTH/SlZIzL2gfu9M/GlFw7ZwZfF7zzXo
w2ZfNzF2ir+UVD3A0VQ7x5KWcLmPDOkiXSfCLjNhWs4UW4J2Y7TaLv9wEpTNJsGOdRVf1ngSBqsr
fLOd4bsD3txQ4pNinsSuqZijQH1KqHqtdTN+Or3Zhlre5MxutwOutTfvy7GbYogakb2608ciqzHj
iypKQncblj4pSAiria2DEOTS04rIHK8mMNOQbr71/qUMZR2iCA8JjWBLkQU5RUXd/VqAz/gD2hlO
wD4flm/5RNi3+iQtgF6A+44XKlkc7Ko4sNToC/JBHAJMZymVwBSvUjGCAaoJV7XkWf9jwSa6z50l
bqA6TfDJL4oRDsU0w4am+eYJVRvWoJLmVC7KnmL5z+N17DCW0iGze61km+EEdwegc1WwIpMQMS26
3RrlniBr/eN0zcUwabo+nlRNQPobA0NpQL1lpgwOtkjiuwcYxOPHojDFi66eZV/H4FrHbEXXL+MS
Kf3S3xlO71bSPYHzElisfI9wvU78guIUEJI0HQIrD3iwD6MC2n9XNJ3Rykn6WYKhi17m1lLyH148
hnuF3NFMebhxsZt3mtjtKTo6zo2efb3Hj6bf3r/B7ikI6Eh3iGkqjJ+JmC4BdStuSzNt/GioUoyv
MtansLvhahlebYKNqq6jZ2fz063v+GhNUNJGwCtgBrOuXzDI4mXoJN3+fvqM3DUtbtwLqKkvlfai
bMdXSVvG/HbAvKFM+FRfns9W6jgYzyYTRVXasP9ZjTyDOHwaazoL1cYfCfyle8TUC3JY50ykGapc
IBljG2s08Lb4JIQtEVU8yT9s0EzmsF3qsTHjs/uAyIIqIZusAwvrk+fSfl2HiKGCtfGXHyQ+r+CB
A+vhZ+OVfXm87ctn30kGTOvY/6A7MEX2qEbqHSDHVh02pXUplbaWt+xYZ0i9AIHTekaOic4KdgKL
LfAsHzvvypxAP6mDHEJyFPIJXXC+mzNT0G+sQd9gKMpMq/IwFGqOEzP62U5vI6uhgeyrytyxCguW
bWaXGDmjgtD0Cn6qsGnXam8AWSb/eT0i1ZNPoXy+yYI+GTOp4gntnOilecTkordbMpn9za3BnESE
6lrsI6ksdiMvRdbRIiXAhnD8ggenINrVQgd2mBga8QVkMWFbleMP3FTvao98u1ShN+WWSyk7hbYM
VnWeelLhcbhA/262yCuPQUVmuqRZSWjyMHfz2a7zXqoYRQwWWKz8pXBXcVg+g9PbemTDJZgyr0Wj
Fy6JmWndfFUgJepNp0H2EEPafHBAu71sfvtqbYPOIK3SyOYj86pp7IzQWdc/w0icRAvQ360hQ9R8
HYqL7AEnBYq93UGgaQQX53LEGaNfHTYCybuN9zSftBiE8y6IURJt8WJoKHHA2tGwfos9XqA0Nitc
qVGLahRY+1AfRhcco8RkNcvCC8HhSFviOseQIWbbm5Sh1L2o7In7ytzCo1cUTJrKfZ1nPUBb4PJc
yRsfkr9CeG5Kelg+Fr+6JqEOtbprl8KUFubUbcf4hVptmEEl1TMt1SFD5Y8/YzYVUfIwEUAmFh1Y
Dz2LrSDULsWaSTrAKV37XRP33MWVCmvESWhnrx7Gp3/8AVvv4E5o7cnRpAcJ3CJwARmoLydVvriS
auf0ieEypXaQe3oFcbgHMV455R8FsDVT2W+aq+FTq1YtaVB142ivXqiEObVTM5eJpZtiyC3u6eeY
NCh75OV8U7fSuOAk6HRkHRFwsoBfHY1aaKq+W86c6/U0563Phhn+F+ahbcrFOTfpE1S9KB6VGlaM
b4k8Hhk+1pQOpJ/cFaqCdZ7XOaaRLESjCdwPqZXn0IbDcbmd6yhKuG9+I1rdEd3EKN2raBTL+tFE
hJ77ZNTuQ9MllbPeRc5Rqc8p9Y0RsxqijnRKDN5GVZr96rufuGvXMuoqmgEF25uo1MBapiRWWIVm
D7qYNdfrhX1nvO/o1vfRWK74y0SlfBN1WL6cus+GUH+2PkQ4IwcEOrWlAZoSTTIfTFFqIBgPDjoQ
TTeeRfO1d0ynKKzWD8kSbdSVIYEojHCSM24O2nEsrWbt4XW1DjMgDrjB2wn3iqr9nqarYisEHPZu
nyRtJkxCC+B40QTkWc0M8s3W+dR/pby0QTZHwZDKr0qzpn6KimVZ/b02GwbRQ1NngKOfW2RNIZYz
SDks6HuP0Yl13jdhWlvUN43w2/cPSkww0BSSsmS3LWWnZZLRtMFXwzbnrUQYHa2nBPeLpXPfQASS
FzP4mELWRrHYoAAgmtLXsD0yawuPATxVKjSzoEU3V8L1VRdDknu2MdBBRbL9ZME/fr6zLLKQuh9Q
39xIclSDPN1tiqDaTSwZ8paSbErmeYma2lCJX7XGcE6oO0afbwYCaWDX2NM8nTnlqjVobC6nGRLi
ScVtbiRuDoW6mFYfKKjVajnerDIGI9RkN0Np/bkMXBF4e0aYKtUaAQ3ME9fNk+KiZpcbDRBQk+8f
K54s1RVxHxNXZBuFMTVgFgrZ6l6e0LAZQgyvtTZKDBmlnQrrjObqabYql3KtAiLTmqIbiIFDtfpX
0sqmHjzyP6YxNa23m5H/LhKk0F4pUgyjWdFEXkzuOKHvO2FlAM7D4IhkI+UWjR/FOPprLJv9j/tS
V/GzRdHAp3IgnYEovmHmIUMsNcuvPVPJKdYlYGa1EZDaLjTFTKruMAK9L3vGuffFSLiMggnI2te+
v8wnJv3NVi2hSMMMd7XGtwBnLw1XrJKcvRmbk0muRSiBHvnwxMBH0yHFgl+qTXAOja5XITY/skmS
z/Ydwz2PSU+QhYina0KQgwKt5bVWC7DO0Ox+F0z/+cUsOlCCfHPODDAIEgNi4CtVk0Ue644YXhk7
jKq32lP9NqMoAb4gD6zTDT0EtNB2EEukBIITiWenbpr+MTX0FUgAwiQk2Oe4sSwwwRKQUhEkYa+6
PPaMT9Q4QE5PJzkaZNwchOh3fKjq34ilZQQfmrZPZtMfRGm+2EGANNlFypMzORqS+K4NQWqfcWKC
s1dQK2QdcrAbiJwQxeU+dkIYJQhN/jGE8A41z/QtkRNVTwUdHYCYZNAKXCYFgdvuXsT8HWy7i5s7
nqFaN5/IQH5uB6yVoFlFLw3r8WengAlpCM1KthS0HppB4kxv71x1paCOs1ddi3vflp4Gh7cSm0Rk
dRX/ManbV8t/AZOutbEPq8TYXtXjYJWP3KIXCF3PDaDGHObhSNICJut5nNi+lJ9rB1ZjFaZL277v
HHLcjKUSxNIR99H1iAI+keIJclb1jzMeIP5FCPLjX3g9XIgwjwhOrcBgSGc9bgOO9sKP2S/DGDtM
OUN3VR16Bz6y6CdphgkPJDpPAv5Whe5LLPkhe2bwiropvHef+dz+utY/tUw7Ij4VTnE1eaeM51Cu
mEMX3As2dWLx3D2XAAPL2yF5xw66ejBKswwbwoSZDsJM6Ks412YZINv3ZPf+2BbzPUYNNceS52DJ
QTYU4xCNTtiUshhjBQb4RL+DX0AMHi9oa4eSR0Hz38ANHgm0pTXrqlt4JVIvLroMZkJnkcPY0L5h
GRNehPH+cwmAXj3VlHgEzUF0lEEADmcDiUHyalsj1GCLkcXzOjzCAgfUbr6gxZbHOaRFH0WAM7A9
eUgSwfxqXMA85WR+gjxla4JhaXW7RSFmpy/CjKgT/DyRMD2572NCqO6dCNRRsiGDGY+fB1Eo++tH
V9Fa9MRmOVekDf46SJEHZmydeJ1ds5fxeDwSNfg+lzJvIJKTSnvCOPG2q0d1X1QljdVya3lz49Sc
+RPHjPq7urYGdrwFMcEtwWt1aq521oik/haUENXdj8881Txaqer3S5FKxpbFW0DzlBe21xJMozgN
sto5ti+QLJ73f4GYbzYmkdJCSYazHWNoCCmsLOGe51f2x8X3AbFP+OSnwCiDa4MxtGjzzoJBaIFF
b41/3E/SnXoEz0LWE0a+KXBSMogAG+rYiPHlNslSUGE777o4FtjDoiF7C+9igER+kNTQWorktCvQ
BoWi05hQJKGzGr3a/FnkGloPdK9RQqs+Qcavyao/9iR+sAvD6aFlk76b8InAuyenwaNYTaflcWbV
qqcucPjjZtzDZXn7woOoHX6/bM3C1cVoQT/TZUYROB7LfwOsCLaQG8gjOo++inmWp5VL3zMdH0yl
vidXVnLcuKl+mCIEqjxo1X96BnIENcv8W9/2d+engTspXLx4cTTaEzxrdkyp9eJFh8whtG4x381/
hN3EWcDL6dQri7fiAa2FMVQevKwlyXQWJ/dfOFtFejLNL6KevBhOunFFKVO58o2+Y+6BaWEidtc3
faA10V9tw42xFgLiFCOz1U1JkyskMhBd+cu1NDw8A8VjKzvIQ7C8KruaZADV6MoZBs9ngHLvMs22
wUFhvqtJHLOUdVyi76BF1lpB5O5Juw+A2XUfjT9KclCzDxJI0ICOyQSEm+1jcnF+TkSky1l3Nmdm
+NAmfuI6AVGL5d3JklWzGERMRRRLPaG0whWSRxPvUYr2MiO5JmL1XoGJoDUAc77JOu57N8zef02s
zVYf67/DpsO7luvo6OYWpe8uZD3rMPbqopRua190xDCvL/bygf5Xi3SMsgKTcZKAQdQuHeo3WJ5u
tE4xtpi45woUvMF4aiGthsJJ19h6oqjbpWz+ekqY7DF5XTMNYj64OswBwXw1JBKOdD9oelw9zJj6
wPq2HhUJc3P1Stu3kCJSlj0ZOtYYxksU7gm28ne3DjGRsRtExErCYyNyFQx3+qx6ZcIVG9YiF38E
j4vsJO5igRPvi3hyG/QwyGwefi1Cqf8pUE0UYou/hsS0+PVDVWzB9zyhw05Xs2B189Dk9A4zJ1yQ
jS1obpqpWvtgICqjUD/hM8hOqC7wIe1JbZEbaX3f6sadYlLE+3paZ4Ixy2ADPNZpkfuZLwctfeQu
/6dE9U3FG9h5M0tqoEq5bFdlggZ58BptflbPCqkZKPSiXT4nDOzySf/1zDWaZX9HtWPYvrg8MnNM
QXkXmuSynuQNMLM2iU0WNi09DPAcpiIXUpncBRw8mXLD4Bvd1epjiONvN2MLpZDA+U9Vgyhe2zRs
IEupJLQ1l9uOvVmSzwi0Ux1ZFFloNlCmYLOdSXmOQWAV1PuxUPJWmIBSh9qmT2RCS7QecsxS/izy
UEvFCCBy4XIAPQO2paE8l23VuLQBkMACliWEQnn4Dw/jQA9+H3U=
`pragma protect end_protected

// 
