`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59696)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeyblCbQ4sc2EXaQ8alTZCMIalsJOpBSZVsirfkSXJdD4P5d6UhHvUoQlAf
O34dBUJhL8/70VbWhnTR7LoE5gUffb2vJvWn9EkYGDb5Zg9yJt7Nxj0A8u0RILQnSCzKuA54va9N
4kXozhAIoCLq5cndhZz2Vlp8ViJNS8APwW9XckJsSrdFGgGRCyMGQO2ivQ3jJChjzSTGTRJ4An8o
TWHLPamfPOr+rPAO7s8fOE7DMw165NnF4LypmOhpB1U+tn6mBjGjgWF0uBLijRQfj9Ej1dx25TlL
8gPq9mQDBFYGs6FZoFR0MGyB+GMpEIskMIcN7OC9YKxbAuc2mQ0CNkdzbwWOT82/peHWWPNRNdx0
jn0fzkNzbnCtZAYvkzTY0FEW+M6+wVA8iv3y3sSZE5dRsdnggaRJ6JCXjTpYC+9k9PSy3O+4hIA+
ZgLw/ekdxqtC5YJuA4ryxXsYXN7iXEUCaUo+nUcrnjXPTRo7n/IjaCpz0N7Dc2OCoFTI9VYHj4t3
6n+AGbTFI1jAPSPlkz4esspR9emSGuTEOsyMRkKAhWj8TDOEu/bfyKq+hbu0dFhMbXc3rM1YPYeJ
rXK8oECcdrhhmJXJzHnKKQgTxt0pkt2PDjx0aQq2U5avEnGiMQGqlD37WwMRthhhde9N4rvhvW6p
+G0jYeNX/6xSF2oGpy9FbeEnDTsv8QkRnK/1rcZ4kQ2gC6P4sintZd9q6jp4b7Gg8cNGZO1oCKGW
R64Z4cLaJGq3Kuaf3j3cMsp7poaTncdY36kaSEmGcGiqZVJgwqUhOhFnk5QiSHvFKqqHMNiNUsEP
pzeyDPYzTafd4KDhA3y7lRFueAJXrlqueXq9CBhWDbo/GW638SbK77E2Vylzm+HOMUHG6xTQW/Po
TYllKCDhLjzfu2qvO920RiwV4EOhXaI3ZLPasZRhK4BJkx3uI3E1icWaOXa4N4jBBibldSb+DfV4
ZSq6rqdCPphLlpaxXjW+tPS9TSt2mXAwdhGF6XM17UNK/QZs9BAtZUmKdFPMHXnQZju6Of5fdnPi
f3KtJHf+Dw7dmp9XxjY7TmJ3dW8O3P/hsKw2/r9ZIy82MldzoQf9IJ4XVwJFRVga6vyG0wgxLHvk
BePPcbg29Or4txr3fS2Bm0QkSjSpfa3ud2glxilKg6Jvx7jzmt3W1Sy4/wWLbMLdkCOWAjoD+KaO
XxbvmkM8WJKlWYZdfKhfHRLBKGdZJzrQN2vFldVmKFdbkI2JzZDtTFtK0ggyIY2rIM0IEcTznK82
gnt1FZTQqdyrDQ7fLV3TUJ6SjMEVZWGqmwTh1Byd4yU+5A7EIoqqERaFDf71o7KbxBhh3u4b2THg
aiCxkXDGcR1MS+tEtloqh2pfNqa7qXCE7BM9jt5VB+1gFrdWHZN65g1JXbesoP9O/v+J6aoTQMEx
1W6ZGy0cLiE9ViEwkXcy6Zmv2Ieja0Uo7QvWCBkVtJ2z7iS7iCGjnCI7Il/sFEwbCty3BHo7G7Bo
lZb0uz3z3W+eAPCfUmPyvqADOOrWtQP4Mcl6whv9pBvNzDY3N0NUY1dQH5Wna/JsS0z7UnX25VK8
TZcHxDtGHez/wj0il51c9qbwXsywyZ9Kp+/3ZluY46rq7ULz4iE20l1n/he2OXZA3M6xZJiydphY
Qa+RF+75ZTuzWSsVIpaWNC9WxUOGje1gTH5/CcpdLyJkvUeyrGu0Y1Vi4jfGa4V3b3lA7D57rrt1
VNTZM4U2/diF+BNb9HAkYJMvS6nvAIsqohrdM5dnY7T7sFgYzFt9olyvUFn9JgaBcTOXGR0+h73d
3KbcDEHoWbRDrHRB0m21O9glUnH6d+YZtIS7TkvkyKtKJtakBRoFygwQlyymCW+8XndMegaHJ23I
blioRs4XN/QkALjsN3n4Ih5iOOi+wRfsSSDZ0jU8RS4k9ABPM3/T1utxbkuLtFuYYkTyxpcCyYBr
eMjGgTVFk42qFnacLQce57oS0EF6nYsZzvD5sFPCLel+wdFOLgwb75bDX0czL5/ARuFarSUAFPU+
g4H45Lw81kqxJrJgEVEIBwX8a+Gd1S7tcNv85rz3yeZVhm3W3uAoE377hX/Kik7p9J0wrexGF3YZ
nRxklcQj0JZQpEQOdBjdLH2NwmsC02jV/2/rEFdi3Xw4A0dgW2x2mThBSBy1+RKprR9nUcr5A7mM
weqv9Ljd0oxYbYonCOCXWaX5j2J1MvpmMhxlCL4Reh60GmqnivKZDxGpHWRsZqMcH2z87JSqTeJX
+0/YUvn7QiBz9dQdJngF5+4pOMjztPPu4PeS9yDVERqOXcqky3gZsAvPLRqNsxs0nu5OpnzQrITf
D5+sDPrQpEYQEARUbkHnOWvp42boUYcFGahnfEfl1PEQO0hFsW/SaYj7Aw3cJ352z4KK6w0bsPSK
2kfyDPO/E+tzTOUJgteLTx78xfkBOM15h4EcsHDwR8GQPGb9n8YFmRdOjdaD3TL5+RnTKKkkuDuF
rEuzuv1rTZ314793D5TtnWBQuuCGPKRKZopCEZ/zsMw0+CDo/7tLO9CmVU5r383cDHEnItOp8xaQ
sv9tKZeSu6PFHSYZR69d3dtjpCWw3QvrRhc9ZfYVxtNzejjPn4y/LjlqqVzvr/Lro6GN3wzGNigI
YV6pZCLVlJJLkjlUkeCbKX62JuW/X62A2XvbKSkpxx1gwM3NhpHR4y1SaAH403GQIsbM6hH1rCSP
zYNuyzh2cBKGLKY0ETSYebMk4248/KjcjTjhUAaUKVlbZszBB1i6CNtnLaz2EFZvLLe3HkQU6+RT
3+abI80GUI9pbNvAbvVkXgeQ81YisWeSIwAJ5MGNwysMLdrcALH+pVlVO+Yvk0ZIDtFaHle5If1s
HLPAHgUUI/7nbdRTGccfAq7bTVEGykdw+Y0ztaHpN4yT5WDf8lIcCp8ggT2VdaJ2iFvuDeiuVcqm
uB3W6TZFYYeO+IPtkguVh7o5py2YJ3ibELEjN/9reBJhtW9N7TeFC0VniFO2Ha9GNe/71Pi6Xbmg
JuqxJ7gklKVJjKoAp+botjk5TlEylC9rOO4Vs1nnwkCLtZdNJNDIQCa5Y9iywvrSpA6vaNblExmI
E/iNKPFVSDXO2NjAbZkSTuukfTEA0yvv1o9vbMCUWu8JFHQl9U14g9ysm6FhgG6EoQDgirY1GBOu
VR2p+LHrTlkSSAZG3Rr7nDdtc/t+1BmEmo3hkVNRLuFBUaZQij4jyMRHtjsS/8LErh8iZ5SfCqP+
2aZNu0vrc60CjhB2OgFGR5X/gGyDX4wSTAnW6jqH1E1Rx8N5zC+uqshI8vs3XQh3Jk6jy6ZeMFfX
yNgPU9pBVwALjPmBFjtyg9Fbt1hwWdj4z46jcQ/NyxfF3IeFbeCbvNEltZBeN3Cw1ZXqQt/mbvhh
cdfOUwLwLmAWQokwGTEwDsiA/4H6k6Xui8BdNb8DmQqqPtutwgPz2dcBNyrisrswhwrvrbmsR+yQ
GoFWLoInZ2TNMwji085E5oXYRxymzPa1XhdRlZbLuB2c/pQgBglhuCF++LkKX60f2RGZb7fcjwSl
auELZ1WOLg4xcYF0B3JFDHqj9jT/bBkkosYJe2eYL6IxRl7dXtgfXjEbev92NT+hP9hmIxHTMsiT
zJa4ZhjxyesjpH383L75GUdXjJ7VVOxOY0fni8BGiPlokHnWtq2LTO9aBe0TLNN2lcgT7ZCYT8kG
Pawre6j4gv7/RdG06YIW0mVh0NnStFDcx+PqTfc8FU89G6v+qkq7aaDfQALwv/eztHvqisP6yKYD
8ctMAl63nD39ziBvEfEHUkSCqofK7QNy/zkqoNdzxJZd2ARMBy1zJRiknG3/55x+L6hF7XWusMaL
RmH1h3uyjWtHEZqfk2ndEQf1mN21GFSTc2bMCtwhYBGOfZpf3Uw5YPZaCrpko3T0W/vkZEZN5FOt
R98w2O89+136/VbWXN5eOpMkh13XgV6ne6WRquTyvhJ0hBqQKsXOOYsaix4uk66VYTY7bPBSAgLs
bo78Wki7Gb8ppcI4Rs7Sx9SlcMsbJojoEJHJYG/yLBG1DNR4dwriYIqYzMDEqGi38m+sZzrNxgwn
KMFDneNxHtndrR6MgdJUjEZSw/TTSes/puaHVyBGNXyO443pm4byHfoyHfJVl9sz4Bqdsgg5kbTa
okNoirnDRyF0U9bzHA/irulO70RAD1w8CvvVA/NCcTQKDpomi/3kr5Up6DTN22v79Eq81sF1fJgo
im9GCKN4HDFQbhFIYfJJ1SDzfqe2SXdAmQgylTGRIYpvbCDE9Dzj+bgn6+ApP7t5RYI/oBxyncBY
1XLsHRRk45TSBJ49I8d1HBdiBxu1Oidu0+OhtmdHYS+/QA6M9eAKmckwCvyJVpbJ5U+DDyY0S15J
6vGpfTglnQdU8rnC+YY9JrKTU2w6fGIPC6h0lMkM+6iBnSTNT0p9GqQtITNaWMadc7H7uBRHIhLt
yZ9dixdcBaLCYDx9LysU6wmvhkTB7z40+6odNDQmLGiQENchZ8Y1JMmFaS8maE7uHlLocuEhRTg1
evEapVF5Fyz3oLL1pHbgRbQdmxG3E7chRO/4xsZ4QGVm7MvnkWu3Lt2Xh6JmpSrEfsnMqQIB5NfS
K8SA7ANx02/vSz4Iv3GpysafRPDpEdnI1Vmaj4v6ey3k7+7vZuNB9cztD/ktQ0mf2RIHZ86er7Vt
SdZqlksiEXCuJmiE7kwoU/nCkXxE8Z/sl085WGU179mXEeChFNp0aKZ7RRv5hXbNvqBXtcdCNvml
ef8lIgMrwlyvF+P2ceqdVv4Zrka0N1X5QR/Wi8KVVAZCzfhlZM7uNmnoUpTpytEqJIBtkVZ1a5zm
EQy0EaZ1a1zuV/2k0vYyAs6sNd8286ewt8+UFYIqHdvjj5+cfIKPS6jM5LJr/KnIaRN4YTQsiv4s
U3JQcp+j7J8phglDEiGfTIG7k43Ww75e2imqMXszql2cy/sL7K0sEtI4BFMvHGxAK6AvXYvCSsEa
p+xJdsttN904OaVKyO0G0nEkdjZGSRdgNaAPNXCaTknpNnpyWYj0jJwuIGPsLxg1oUdGfzgRDS4G
Sqvf9Kd2Tso9ncUpSlilA+nJHuPc/4AcpYpi46NAQdmPq4GkPYRuia1n9XUxJlReXM021yG04xQ4
UIQBVS3ckLtZHfD5I7aNEtNPVB0r3uqpXcoKIqxilxYe8ABV1grwyWvH8bZzjvaAZhx6lepi/5pM
eDlsEBFdPmMK6j/4n3M9qiqQ4zC+sPlELl66JfpsfHVc0TBrDK/dqrkYR0udvEqlTZoGkgSwH8IZ
YD3x1r1wezpQLbE8Qo5WDdCJZOvSjeqEQ/ZCcJhi2lRZAcsHu1KfxfwwtAFUyGLkwzbh28F/pFvp
O/xHtY6kbIZ4gWZrS7ktuP87dxxZs9o9dCYyn4AKEaclrJvJQ7J5HStkfY7vevcFeNzuq15W6RIr
oRNUB4h1yDmHGh9B4aDjLFW+kbUtbgDVlB7+9BHVClGmBGkfL7XmC9aFiN6r+oHTaDfEF6bjF7Re
a8NPFztXD+DElF0L5mwvqni5c2jxzs65Ztl5pXwfm5Cnxb4RPb0TVBmnoEFOm93XFAm9ME0Jkn3q
oz88u005cl6rQhCq+D0xWn/A2bTWqCYZTdu/Fli6aveTcqZqtVqmIIQRzGfvTxqV54Qppn6eFlkX
ZBsmNj++Rgr0U5SLg8XftGr1TwdBZ5KEkfDxJlXt8hvACooaKuXYjhD4LqTnq9oqbaO/sdekPC1P
cDqmAKHlxEfCciTqUQgUpcX0xy1N9/SkOJ8UkfafAdgmAzB5Els0smUxiszfG8zABHh7H1tFpTj6
aDxcSmhyUQ637TDDCyYbENJqelMik5xFa3BC0Tt2WF7C6w6XvIk9lSm7VBqIqNMi6OveCEI5fWmq
zxkXkOWqGXSeX7K1Oo8ETDFxZ5m37G6KNKCLkhB4s/7EN3dymiTAavt0YKKJKMFCHknVRimsKB6b
xmAGzp77rzq0Y7blAoihe7v3BZXYLgrQBSh8o492Tt5XG87hf2bl19f6++93UrcgehcTap11AE/7
8l3Ejc3hhXW1W6SPrc4nTw4h2cPToAbi2GHU0wYxuGQP3VNky2JdmynPX8t4JPKY97oq1w7GN4BF
Q+WfM8YogPepTt5hv73yQkcycjmJDZ3fAjfnWmFegPeHd3ItU3+z9hYg/dLRaHML/AmepQfo161g
/3DrEQaEO9UUwPZ1zKRtMvjWPu2VzayMuoYnXYEw4HVoEavLBpgPyFYYobIzEKlISExJe6PUPpA+
6DEzcJK2VdqfRy1ZdzjZliZkvnmVd6fSWcTAPwhjZRdFYuQzBK9mws3qP0kB4ytdw0upTxgwSNzo
skhx5y1pe8quKInt9BX2pmq65y7nyv/3S9uPscGW3FCuDUDukcGp8faGW3KpqhJwfgUrh3AbGRXO
0TEL1nQFXI/QSC2vZmoMevJwqKqh5iV7bmjZai+geB8qkVgicsVB1+VVJwkMKOSsbJsPHpWi5XCx
pytiQCCckCyhQyDCBFU5BU2jMPNIvnqeG8w1b0slnB61mStkRwOPzE1yWwJYhbNszVyhkWsjaqxc
2S97sQreiAyAzbXp/Gqr2knBg2aFg5G3Pm2pNMzhp1R6RxIcmrwFIrPk1y+kkERPorDlarDCDMsS
HIibnmkglEhflt6ksaXOjRtdPd1+htRnunDnuT7Xp5M77EOafIr6nHUE80PEmwMKGxP/juoFL2J4
XdZG1SzE6SbzxcQEb0omtGlIUQsyovJtTy1RA4se9706MTB+tBjFoQ4wBjOvTHab+I++zsTnPJZy
CxrcksCTZZ8b48j/RTpTkG2Yg5YMRVeGYsv53oMu4WIuu47HqTn+WdqW3USdzkl6zjqHNw42PJuk
opdG1+nbz0oMTdu/Ku3tpgUAAyi+Fl0jQfg0WnHmDl+n8v7vnsjVVkg4F2mvG1HHvUvuushVGCy6
Oo6gtwzakWQ0yo5v7pNKoIuvci4JuOc99wjel9eprrQSkvKiSC4wfFMHkLzLeLDgOKWWC7Jue+zK
x3u63u5U55N0LJj2CaPQYJG410PZOVKSGq51uvw7q3Bdi6SH3hlauYlQPy3PMQ5FCIt3sRVCdAfT
jTMTA0AZA8I3iPcWlTr0X1fVl3i4bI15Qu4aimFah1aKQT82X5G+Rag+ysmx3/Z59q90rdBuUva3
GftMc30oxh6gZ1Il8SItJEMdGNMxQ23B0gbxpwh6NowLrwVxYoPjT/psA0XIx9FilfFLzORfs/bB
Y3armCOTssbacRajfMCZmhGSmc+ipsNdW7JqknOlJ2+4aGb+GmLxTeMShEGhufOEsrtwGNr/tF3h
IJbY+l3MpfehXr62v1wcO9FYtp+esRSrYDXYXtpm6GnBTIYZvVauO85ByN2/JT+vxI/GYr7JpB6s
BUtJXdoyi9zY8XvWzSBwOugFFzwQ0FVLD13uKpf/bcd5TmcZLPzSWT/axXwjss2AL/m47UEQKc9/
t1VoY20VyfPTW+xkQyiHGp08MDLOi6N0o57uwJ/oUfmoEf+9jfiXbgxSSzeuPfCPNAGxMOqmpiza
vR1NOEdnhWpc06I0rXf1wxyVNgLHeVylOpAMSx3+2VtILIsD3yv34UyDjVi7yrOef+jvqxy7VEh3
HCne5CvhozzUvbcLcB1Pu7EFM6eGdbaW1FpvqI2o9mxMNaeMUgGQ/doIKJjGL+SNQuOAb/QI1MOf
neFl5cXL7wd7NWGXXRclDyJSluC952K0khBuDd0LeF0D6Nhtcom00SDaKllZ/E1bjZflewZUHqBo
QrJIIy+Ig+L/r/w+Eqh5TyaaEt0l/2vaxCPiyybrdnbdcizvhFUoEVrnZGRmb0F6h2H5W2zqVY3j
hd0BohEPOitrwPlpfU5i7SCYeIC7gGrUO7VU8qNLpihipaOC52YBK2+uLjxQ5RGphnfQL60d785X
vI4aHwjwnKib3BNHOXWAoNTnIRqofM8EnCy9lBz8D6Hqjeu0X/ruu2kgZj1h2HdVsZ/ELwQdJumE
/HxdeBqXE8/XB3chUV6vcAnfRQ/i81v/V8dMNP7SJl6s9n/azTd13+ZGPPHBxqt1ECSn/C9duuSV
4M++IZiy9I0L462HaUCG9YEqgDT8WXlnO7k/MB1Q7SNX/qQoZkcFzpekA66Ri6isYBM+4edddJ+k
fNnT9PHGiy5MIbV1gPdVFKYhYYiyxeyPJ0GriWo9K1+vWYBy/Oml5yeSH8yD0qgzPM5e03u4RLC/
RaKpk8LWa2xZN2e/jNQK8Qs3S4zK8/jpC3efKpHcoiKMPTurfM4hI3hsMXWNL8r2fA+ZOnO39puF
WSpcemUf9hgCVrtAogShsv1pPU+NTGcAjz9Gbp0DIT4EkTVP892Gd3seKJP3aqMcISFVpF/iNrMP
N9a11puVQjr2hQYoER5K7U22VQB5oDZohXrBwfHMQElIosIMkxtMU3Hj+wStgTcqadYCPYvqAia2
QWiO9OhAvCQCBZH/D28sxYxLh1zCDAbMqvBlx8lU3rmjlUDtv/Be4vd4TEWqTzKBF/Os/YnaWQIu
e0RxMBHtJ/Y7hpeEG1NMHZYYbCIKyTE72ZaqdI4hukGkomoxjmZMtBIwgZwqGMLFYJLkxAC4VG7R
ZpmmPXieesk9NcBz0NnnK1uI+r//KM/rYfl3Hl1tXHzvy83K1Yx02DbzG0bNeUi1vh2/F9Zq/cgQ
4a3v1a8awEmyH2VPfeK4kpbhgy83+C0aJStXk36hadfJ7Zwho5CxNb5cBw8nWcPDj70NTq41VMPF
MXR7BO7BvU4hhwEI9UEKIbexVrCGww55eYeAbAXUg7/t6d467ZaayvvTLo0ZWg3wwWomvfEhHtup
lfE7oJtEZVAk2puoKeyiRzbMtVUgiASoVCEOz2uiLZCEp5+K2vuA9CsPULVUwA8efFBgBOabS9px
np4LBAnJInRGV5LLFJj1uEO/ozPchly9yg+jt8xNOhuJV6yjH+WbXGb68XdYQvujFAje1Jq4WZOJ
NFw4reGFXTfE9R9zzj/82YyHtEWd3eVknIF6SEjHXNs+thhb039q4TYWKA5FOAewbsvpGj90BIj6
0Jh+6rRMUIvVJLxmCNGwh7e+0t5EFA94FehdFzT9rHk1UOsf9D6b86j0obrXd3hd7v9qdm04xA55
LGlTkDxLGytRlCMg6DLREZR+R2NOODzwA5+blLdQDfta4KyXh80lekDfOAs288aaSsv/d0+2X01K
YJWWqaY677k5rM4u8wzibmgUwUA0qeJVBYPctK1DVrQRq+U+y/WInNqx5Iu2HVMsrGP3+VoIuv2i
/95E42mPoYp7+23W1+6ZDpSHc0pqWckAUfnhsqtRnqlpkfuiGrOpWlfxLnYRmvG67dwBcAYig3KD
kD4y3YdYiCApvDbG1098V5D7vrdkr7ENin33NSr8P8PDwbiuqs0UVd1/OgYG97UIelOdEpL2kK/Z
FGTHspAK+c8uFoCXK57W+rhBzEiOk/PbokRxFSDskG92JFSwf3/oQ54GZHB1iWVcL+xZ3TjrH+Ll
aswVuGdqqmdLWHsRLI48zjpLdpMfcT3aaf6JowzsU9afRhaS7Se/39EY8qsZ37M1RVFI3XJrWTbP
9JF1248dmPRFkAXAFYu3GfAyLlVKO7cchkFTCzY5K1SfGo9vi5FsBqaGBrKjnc1O5SRGCurtjPVw
ooVbAgR0ERzZcpFwb58XPh+e1bz8d1PG7P0drjprA9K7Xs9FgAAWldgGGebFoe6az2dXxZ+eaUK1
vcsJW6O26BYyBxIFY42LZ160P19B3YVZlZatz5XIoV72vZ2JpLeLkyPXNnu542+dFJESLrfm1ZNc
LVhMf9z1KWZOPcBFVjaCPbTQv84cWHYZlCq0YxEKkU07BRAgWAsQDTz/akMq00OHo4XHGEr3OGBM
lXd4qD7zmVAXKSj9iUFi2vbqnsGL1x4fQnVHCEss56+B7PbO5TTSU/qZtF445wLUISu2J4tH86PR
yd/Qt2CvNrPTBon7T31MEt/k1lH6CX2QRlbQb7mZdY0ZXukpo1Ax7sq3ODXyTWWla59sVui0s8Ft
k3URjMeCJhlS9xGe5jgW06JWw4JimZ0LtHUND/tOJY+3R4OocpHAiyX6sKoWTkI5UtbmM28QElmy
413iol9kH6mHzPjZLjw8QZB8YPHGqDdXHPWkgh/4oOgfq6xDz92y+3odAlBJpAAZ4knM27SwmFiD
11poWrteTXKDrszUNCYRjfrXdlXIKQK80ngTEVU1sykFI2c4qTFSR5o3/YyxEOZOOaMvjsafvWXF
/d4pDUoztc2bwj0K7z1k7MjzVR50WuR7PyeLkZEeNTY9b7EgUPSgZqXaUT9qig3Lz6vPtTNG1OrB
uP/9cVe7LxQLM3NJRLfO3DbnJPoXrkhU2CPp51hfd+lUX1GGWIcLCxWyEV1nQaJIRH3gJnOS0P1t
4SJW/uM69pkGAsHQYeuxJJThYL6V/zcv5gv38qtVncTBFkTpHmWWD4KaTF+qy7tL8U9yQzosEExF
JfvVVXnYbWasOF8F+94kDpayHPyuomrdnqht3kAGhiwj1e6NClZ2B+YB7mtoK6NBp8clz4m1WEmG
pNwx+WZ8UotNRh6nnnmpjLZ42MUDhJfRtGl6kuuDyAtw/PZg48LDl3gC3ZDyY7AxGaz/y0tyw3CI
trZLKS9xYsa3xO/sAeajsBLTuw2Cjh6Shu1hSm1j3fMVK5Jn7ZTPqmRJklz5vKcGOvgxnVpdnJvZ
4VCYsZrMykiXjwHfj0y/vNREFUtcxChSrfStcnEWAmnCwuuHHujNfEJdblIcZl6iKjszh+Co+rxf
7udfAWaSAalOl2O2nUOzrCO6+3XSq/YOjBte14+telAb/hGlQS+xD7y5OTxmNMM3lFlkOk561Ma4
t1Gh1QTvLrDJPONxtInyNDw63mNcsryR5IN/HSPOOH6A50bY6VhRM2RblHR215MZkfFWO7F2oKF9
ZflH25foRd1h7saESm6zziOlVo8Z+Gh3wPCqpSJQzhIjVzeOchLKd7hRAt2sYNujxKxLjcO37ep+
+77XVvMd7DiJpQmMsMCX7UM+ZT67BEbbaMrtoJ52BCwPi9ZQpAPhALDmc9XDOR4OCPYM5PG8BuX/
4+7PdG+zyt/joHFWhb/032lVqsw1WJVkX/0nddIPC6WZKdb6riOFPL4zdUDOBiHW5CxH2T1rQx9F
DmG4vy7S7bh2gVwQW1aorxFwoGfRoh9+7gQZkfjxDZ93ygkmi90sDydNYk0Nm9h5z66ypCXnKod6
1KzsZ9Y/SHPyN1coqINmrcTndlo/whUJY+VOTs+5/Ke5WraIP+SxrbmyZp+Yxhymc2F4Z69mFDXU
I0CIKIGbSZ/KmG//LmpMt+YxulVaWNmhgsz3H9Jgoj8nw7dYsfu/zKK2pcgF6KikhRtoZIZA5nxX
AOo0NsRSlIxtbvx0esulY7C7Sunt/pUpaHjAQoymrcCRbTyHpbPbh45UXPJSXB/wZNGHouAgveZg
Mw9JCYbqRudpHP+WpScB7A5rr3+K6ykJY/OZWtfyo+63qidFFy/eGx/FsPYJYSeXrywH86nWCkE2
cL1jROI7Aej2YJwfteRo9FAEukwrEs0Y+TjYpJZ4sQjA460ANqSjqI+VvZ+TlIvB1H3bpERHc8H5
rs7q3hoMgw/iSsYM5aoZYP77STKeqfvvAoxivM/tt9zJqdx2XV5nn+KEqTG4H8o7cCtM5J0N5i1h
+SwU717MvwSqLGecJiac3HZB0cwbZ1J8bq46s9dMucQIjQDaWmEkeYWMUEsxadZIGJy7I4CWdFtB
hoXdKBK4BwcJUG6FVXCHLGcwAwgfeFMPcCPVK6dPDKFwAahfMAqXaDxhSEig8U9Xwo7ruGL/ig24
Trsu9URwDtvwaFEaKA5CoqBGGSL4IntsDg3xtg/FmpJhBH64KjsBhJJlcgQsb1psVGOZBES6+7O+
/ZZ0J8Pxc8Kmeo7GbehDtoGA8QREE17skivOdNWl+r7ceypAU3k+gTooImdonwE06yjyqTHz0GgT
r304vbf3pFDFl4lmMNMd8xUV2dr4pjNnRl2gbtbOVipMdz+g1MEK3g0KF0bG/DuzEAv81r6zn+hX
OS9Zo/EjQmdxu9GcHBIwI0BIL4T2hfRJ79fKPBPAUIEUkXZD8a7/YJKgaz+iV42XFG2dXwvhgdO0
rlJuJ1Jrk9Db4WLZfhQ+noJMg0xayxsMP+YOYS+KHF4TXfGUQ4/7ychRqs63gyvieSjgHmNaJjSW
GhGz8/3TeFM5GJep5W2EtaP5EkAQjgDOUzTEpK9ENWiaSdznYneDFwDIYlb9uQaBQh7QlZ95ux3g
hGSdT7HufxheoFgDYPNMfOJ7/mdNeUCHDBoNMUpCeAmfMRsV/BTELpPKbbFMzPUleWYEp8dRnkJj
6TwCREcySRtMivSAa8dPzQhwYWpx5dmXl4ndYTjiI5fX1uF3jmR0mgrFcz7KVA2vOoCz3QPTcGG8
3risAOlt6JEfxy5rCUN/FE92Qxgzs517C5O0VviA+ppUcqEkqxyKOmct2IFZ+43esQoo9ja6Iivz
WXjN8GswxWF0obMw2GEt+WJsiR79FvGRnqGvHGSvFEnzSuLG5Tfc76lFbCPTmAn8IkOLYYkUVmyG
VArBRsogY2UIiwndgjr9cUKGrpPJUUQ0CCFF50HiXQ5jbWjqanrP8zawxdvbOwB1//h9ZBNbYGE9
zf8mg805LdoM5ixCAdHyfC4LSsJlpbkwj63pc0FL0OF09tSwRyoOwxLj30WATevGXtm72rYwWte1
YNBsQbaDy8VKT+m9tlLqR4A5PS30zGAx/z74iUMUigWVH7pxELg2NDf4+gx7XEtd3X8Pd8GmQ5fz
cY3Wn1EOe17jK5X2tOKZxpZJ9EOcvNa6kg4/4DMwV+aLM5Bkaz3q1T3Gd5WE/krnN/YHi+ARUUk2
4znpSJnzcyoUk67GLoutogKg7qU4bBpR9Iz+FpS0Ncqi9uKVJ2NoVEbvV1O3bOL9MoKwXxibIxqI
tFEO5kcuqy/G2N5Ir+smw8m0/plpY8DE6ZvuqYrK4peOSl73U9OTz0bRUuzoCmUX1Qvl8jBZYcW/
7qv+GP7RFiyoyXUrhyhwRXCdvc1AbojIzjgBJnp1MT4FVMU2f0hQvRTkDWsamGjuGO39lVq3qqPa
7GmSZjO1bwmAxntHAHQ2583ShQBYjB8Kr6zzXZm5c8jpjqtrGH+0ZPy9LVYuNf1fjU/xlQfJiCxb
FcK0lgZfHty+aqpppA+HiThQ8107WLXVQB9fgdbl8ey3CuN8p++fuNOG0ozN43DGMfSaYvDA1g7J
jPkXNMlSUVi1FpAkuUxHW3jWrzmz+yV2n/xxJ2YDE0KgITOTb71gPPt4XTpyoHal/ATgVGTal9bb
2LZcnlbzm3qTOMmBPn3yleu3HqbXts7fpurPkCbLdXSauMh5byFzf3DFoC0TYPuAXQGc/pMBd1mW
XIq3eAN3UtT9LLqqw58rECxBtA1iLsCIqfK5/cEXL0C1wuqIXSDKLi+PV5H9gZJyx9+lyWpGsvh/
mkFP2ejWuKsSj9f4xYcmNwiByVdHQxsRrpipoUEXtEUwAQ0laKUt9zSC8efX1mVPbEBlfJbBmJIy
nukYtU9lZR5co1B3rUgyQj01k72GAyCQqao2kUEDz9NDleCZmax/bSkxr7Z1hB2Aa7uS1eZsvQPr
PSfQ4ZI+D/4GzF/w0VpYC8jmFqgogKOXAbql4wYqlZtU2EpXhtShIhmzkLAXBK5/kdrLx8wAowGk
prgsbuCo7KtV9EK1ClzOIhRYRlZs1Pk5JOoVgyOBD6JdWqN4Zw4ep1Ckv7h8m06uSWPF878JIvfk
u0dW5rn3UDt/zs+JYr6BsKhwti34eL3xInwwHob9dbicquQvvsi+hypt8KV66tfeo+un5zJewxE3
1Y0t/EMkDIqghehBgwBVCQlCXGHmwLcpyVpik3xwJr08mpBVkgX9QtuEVcUABWNtuhdM4RwJPnfe
CYnmFsxEGSiRhsqXeY6PMaNqW8uLYwoqTUNbxerndwWG9UxSeuI6yib6MPVaZ2l88NHSS7f4I+kK
qOEo4jvOIrPhstdoeMKVJl6Ef89KCCEg8qqSiuHRZRe6XTeNtJR6fzl1XVfcoVM5f0FpY+fbYrif
a+iziClO6Fv4isAgM0BkBPqrVZurFKfslCsUF9WmlkXhGnrEnIcz2jh+73N/Yp/qMHw7XXR/KV1u
cc+gTSI2Z/adWh1GBi90cHG+jRo/pr0QRgx3Euta6SvwPsTCmdpQiLTAgHk+R0pYhuMcgpGH2H/B
jlzUkfiNqMri4A3YxuXcy9pjIWswWbaomlxorr/I2N4xUueXUJ4rIHlljKgPGVFEsElb7BtlULR0
bwgGQhYEWoaFBagjXRUjYZP212vnghDpSKjaiKRQOscdfAux2i9dk8KcDhxzP+9LMeR+AL0wZCYA
09xGsz08ZWFknB2GDSCF2piBdaJqM9CuuhgZCcMuFFOVyD8uyo7NViAGCiyiGIiCdJ2Jf0yjvSpU
rDFLByfYUEeE0qty4mgQIfr6X43fOnXnrdI98cjxfubieweNpzmQEK3oCMWmNEdm7chXp0J2mJHE
kQsdQUe08cfD5ky1aztoMe4MGngQt1PrnpZCe8HCeCXmftOJbcOTKBhfsQp8szjmwf5S4f1GBrZL
EC9n4vbQvbFaeZ8oB7QiwgRbwOU3dUmxvJTZUedLI5tUoaZvaGZGfWgYfeg+GajeZNcXql41J7HH
cjHJFTamV9OUPlIk4w1wRCKbj3ASR3N345BzpaV8iohu15I98Gvur67RiWCYcxyPdyYeQSL/Q+0n
2i2bEauL095TSi0yNNgsa5h79m1ENQ1vYkJ9iSKtRwrDlRK1ZHs6MkqQccbdX2F8rHGuxnxnsfKe
in3ENSbOy1Iz+fyNiTUkF47ae7w6eonyyM/fTmX+kPMczbsoe6r5gGojjHuoz7t84atgaa5EgECd
CkFmUFH4EaNDCLDG4qIyDxPtFKgeiBjkPKb/sC5LlwF7flX4ToWlYzJc/k9oSTKlFcL8fpMeNGch
5kTIx7QgWH7tKaeBdar/iJTcMv8JqAt+nz1IJ1TrOtyb3ToTalwwmPGm3Lne1evwHcpEebfc+MzP
w+4QczvrFm1KwtqGtDkSMCGcdth0Um8iOWzkblFbZpDlb28jF7rbYa4u7cqhTVfQFy5gb2X+Ue/8
jdEJNXauUj+ZiPKxq2iYY+iNj5ZjSD8t2V4WW/IofomCEY+wBNcQUpsYiMeoTCTJjGb0QZM2PSpD
wpmmWwyKXYuyggLWBPi3TK2e21EuvjG5dl5ntt5RvjW17yjSV7NKzDT52pYslsoOxFRx6MefOjT7
ErOb4iK22TsUtlLWfIItoRgAV7+pQ/EJd7jNTrRHsMcFCG29KSMB7cU230v+uO3z1BLIlkX5KVKv
kaGp91wVsCOEA7aEcIpPgvzquazksUHZVAL+aQLpDCO8F1X1ss25lQr8snDDrFS+o46Yc52qEWZG
by7t6IVMvvF7AcoKbsSKf0sqhQ3VWGswrY2hwXuIDPnWCpXjM0RLM3m3nlHKeVKWVGR46+qSfKXP
PW4fEQNQLlLNtZUwV8+XuEXfwvMkosHBr+8wIQI/65lXXRsYDUUlk96NYlT0awTRgjCL1L1oHAlg
P2NbjkrtkCZt2BsWb5Fo94vPwTDUben+/33/RqZ5Roz27rMJXgY4RmTKU4mmVYwYsA0wuE7a4y+1
vbIEyTH3Z2Sx1CH/TYdWnmXIGh3ZOVKN0w2HJFQZRKJSCaoWjR6P2nd4q6XN3LDWsvpkT2/MOfJP
a9fFQ9W79fzB2zDaXx+TfsqI5XQTNCcQTam6t4gsl26QczyM1GggrN/ftQipkCM3loJ1FHcK7BdB
7mrn2zl2u3Dz2osj2taNdyYLt2sxQkDLPF6/dUzbEHPROgm1H8XkflJButjQ11skkL6dg62FwEIz
nOWHZbSXlP+3E8+wSUZIg+BXSI31vViXFQjSz30MdOfta+8uTIwiuvvl/gShXM87hT/04tueNBz8
X70k7/SYIdE7pP5jqPa2z7y1O8p7GJIjhjbU24YDztVzucin/hmZYEJN2uAuzjpzVitW+YX3H6dV
j9D7e1WfMOnSGHPalP4Kk/oui9nq1JRQ0Wz3ykNvRXjpPn5F/c16n2hHqMpQqdn+JD6NKrr3yjmS
8utbxeog4okCKzm1QsryTrBVsLK6dfDmMS9SOyNOf4GQL6sPz9y6aUCr+ztvCmDsByY17dp7XtL0
L2cE6+afS5AXk5geYQHfVXZ3bco8W3itwV1Tr/QZapoIhIXKlFXR5e8t74gK5+dKtlT9R1vM1hyH
H0dKG8FvXZnpVeGpqBinNKoYQ63fVKwjSgZc+V5Mgmrcr6/UWFhdHnAIb/eLOkp5dYfbqrMYzjvp
FfCW2uaSOzmacZooIrYKz76Xlm5GaLVBUDBBDQyJqdqCt3u0KZW6bDq/vK1X/cUN9qK2K5XaJDME
vJvw0XHVDSunKMwyG/pUnCRtFXrFOMLpLP4t0KiA3m/LLt8cNjd/NglUUnixWySk/koZ09dPIoo7
7AchcixiaevN5rwbetjz+kCpoX1NHx23OjbnVfSZEvRK+q+x2K2umllrik4xFqhl8Prijcg3YtDJ
5iAw1EezwYnHImVWZqE5CFYHVW1BA3ly2bZGhwMsJMxhSP24E3TGfHp+3haOmWhTohVHjPCdDZ7s
cBSVdvzhJl8sBcbx4Tgv0cJc6lyRiV7IhBLCcJ4LSRrJwSR1e4UUn5eW1Dlfx8m+ryt98ttwOYE9
A+flyqSE87fY8yJaUZD1zcanDSh4yJfpGbrFu8j+WEPc22rFfMoojs/sESDZOjmHJjx/YO0kHY+B
D9GgJapf1TyG67nmkB5L4iXuZmCoev3Z8cg70SyNESULk4xyxJ13I6TSqKqbxW4Frl4Pjqbhv0tQ
u5OqdJbRJVp3gWfP27LrD942fO41jksQtgv96gfOycmPviowzdXuPycQ553MoDjek/FZqFGP7QLZ
I/OMIdGmwt9bfDjeOPN0H88bCjuY45L+zMTq7TVCQvpsMkL2PmE48xAn7/tXy0vRSKi4n9qL3aYQ
6xq62pxZAaq9OwIEhvZ+12NgJii+fy+LF4LMgX9GQIlO4D/iw2fz0JbulJEsud/2U3O/wSNDx2Ic
OmysEJl6qQSatsFVJf5QzJkcsknJkfPaF3VLoMD6l5kUiShkPSB1UpTw0PJaPHRm/pU4hnJ6RDPF
8FX2D0BHp7Qca4FMqjIzzSSOJc3EiIi6GM4UbMsQ9A5eShiCHQZgh2ThMpMnaJr2fIw3lXmmyu4U
1AhI/17TfGXEk7BMA+kI9l8GfITVKOaAGjyfh5zKXFgRKzZVbQf9F3OfQS3QbuPdrHZiWSK8gzxN
Xdl3/x4LLGbUmwehdd07XHNnMCegTUUBCN7UVWtEU31ChrigtansLwlvqq2mE5bFsNaVEF6RDoqV
XYMY/bcVFL17GUdrKxyhlse4UuOirtn/KAw76TQg1VA7BexIsnQOPjqswtPsN2DaEyjQBcFJ78UB
tN9rRbNDSV72tI3Gu45+ilvPm9MGYAUB0R6i2ggN4cp+JoQDoRIQ53hQcjhtRT4PPqh7wciEiYSK
yZ3nVVtqWP+bRg9utNFIU4vW/VmcfkT41UkyM8cqGr9aH4kzfMKn7WgV3ZEJ/4aFvUydzR94+UNc
etGS3urhoLiStApgRtwzDePKDnuoguqpJ6bCPgSW+lovv9wRfvEw07xg2HfenOWqwS5jUW0Y033D
dHjBPI6JZw1nQTP4ARMIswdfd1O4vV5YbHNnlSWBy30sB9Qy51rzk00beJWT7sie9R33ExIBr0r2
f8Q074tNAyN8ZmJS1C0mpcvBEfbDv25zc/y+MFj9AEeHSmaDo7oaI/X4nzSh4UlfpTCOj7NSRez2
7PV5IgHTfxr+BHOW0OFv8LSXOIkgRE6c7AZfRxgSzwbduoolXejmqs8W0lbJsk0jYUWvaakqa7B8
ScXxxk8bcNPSqryR1PFNbFeQL2cv85YRF5CMkABgIcrzOf9olgxassCpLQ8SYo/qZaIlmL+bVai2
7vmyp9wTypmOTIs/p1YoGBONp5Xd05ngexaFLr+Gn88W354ptFRS3Z2i+cRPsHHvhrclkzpO3vCl
pmSRus0LfJwVU1xyC/FRHfDg4nwYtZt956/8/YUC3i8/ojEsms6a0aPOT3bi6vU7WpuMy1/x62fg
aeJ4b+RW3Ar7e3fE+dxi86K8wD+Cr5ZpUTy5kSHaKnHD0zwOPtySdfnOF9hSaD/+NW4lHseC4iIC
yPz1pmB6fZYXGrhp0u52hst3iTb0F3Ng7t0w1+/+YDKm/qd7tLguzI5RHVl+sXDAtiMSt+UVFvqJ
zxwfQOnFUXvJSKYqrqSYxAQDVq1j0U/W5znqVT+8JLWUIOLb3ixtBs2spcW+wGsrMrrBsVscOb3r
dqy8WDQeY2o9lEfTmu4tS1W3OA5VjYoExOZDau3PR1pbr+UG/D5dpcCWoSL8IBPc2w7cwAQNtrY1
9vl9s+8ygBSHVzG98NmJdnfovxYrDPjM308UNMNBjq5euH4qTm52N99z6MpM0HbTBWBZSuIU+Y7y
5XpV/NOCl7IJSSNTpIXNGd45n73potUBf0AE1u4Dr4k/fWaqMl41cgLBqqV5sEprTk1MPWglVNmn
EorQzmmrQr7A8zRZwu+7mFbRReNesXgkpCSceIKIwJNga1T/JqWCP6BevNqrVezZeDlB5VFIgnnp
96g5v6jxE2dYXaMfowhICSDIQUn58ePgloSoIXZ1LoYY23W1BXPOYG47zvc4BkpcfEwTMM3exUMr
SCp+uSOBMNuiDtht41XqsqX8eLCyX2/JOju27Kssp+1pKniDPyTQ7Z/nJtB2Sn55ckC12elS5Poh
DtFSw7bAXxP344gNU7seJ3A2Gqga7zk2LHU5ZWuohg/ocEkC6JnmhD49oxR9FMIdaxWS1Lofg/UA
DvxFKU4CmZywY3RRtbE8k/bWMQ9WIugYnb+yzq27QWim5nT+FEagD1er+Gg/K7SU032JuL3PqCkx
8C57UqYIIMgO3k+72zCA0Hq+oo8vLsEWBqDLAae4mV3gP9AAcoQ+s1I6nbpdZyQK36JuTPUdRd8C
qqFy70R2PAeacoeGBGvJ4uRu2Y7v17PPCzgwJ3M7Wv3wkc004t5SeGv7dzQMjfWD4QJWErFydR67
4tFFQoMGdZABsKLDwA7v8vNsDF2Q8WhX1cUwKY46RWTNgx8q90xhdfnSLvHyVbvPjXETQfaYjcKX
n8lqo1sQD2ToT/xnqEwWgkGx+puqRVHTr8jYfKfuzXHi3T/vUaXukuQl4D1RQfMQdLSa2HpjJSsb
d0kPm1+kScY3WAgDPTVtdpgWlDltwfP8c3XeHk2icWbJNcBEuhH37GKKkCB0A16P1eHCpmhOIkDl
ujVOtizqU0qzYA5DnYJZQ6qBHVnC9JW7JilcmUgC4Z+vgNHnVIR2EHXX2ia/bkSnT37WFzwGomO8
VQlni2eF74F2xyG079oV9hiQIN5aekMhgYO0Ij+LlbY78Bm33UmVjJM7Fo/jhd9DhMPJ4h04DLK1
vd7yV3sWDycl08gw7dvZzs3Hg/z+9p+DZx+kz18gj46xUNcYw7qsQLwvU6ybVtO3Tqf1008TJWoZ
ibxZHLn5dpQTwyI5oS+4iAjUiSumEZoImlUIIucdhORxIAu9rKRI0H+ye8TAFZVF4Eku45dCbdow
k2OfHdzY5q0q6UZ/VGnQ5ONB+I/0KFkCncPBoKFgHWcLqo2RUA3vNLjhxLXbiiCQhVyVx30ZHDSr
X3f4eKqP13bReQ9Xdg4P5veMsB49/QuIdpPPpoQ/UxI2/GQSoOlk6Ihck+gDe3RmOxNPMO+b/jGQ
xdhmkPlMLpShZg1J8dZnWvtSgkgRQW8RSbt7QQuzbn6noe1yLYJ4hY1/puezeAJatrAWkriupMrC
DNPdbXgMGYxc826yknwmD1usTodAPw9boFE7imkhzBoCwlokANIqmGQgxEIj/h7nafWIUi7lrOAw
API0BgtOQIdoIeo4QZ0WZHFGtvxyj8Yw47HxY+bCxhS/uUsQTMoD0bIcGC74n/k9lRTj7lEdCGU/
nbXnHHasYV2ajU4+xbUUchGdrR8jgagkj08LcMPOysiRIvlCDdTD/RZN6gWnWpaz1Ww8ObeFFEUR
eXJ6gs12EUDZe8/huxYLvEC3yUA4RqHfOTMgpsb4fSepv5URZHLH2h7q92w4s9NB2NFeP7EPnVdd
LBBZILGVCnZr6jCAF/602qKZTZxetubAUa80sZUqVve9N6QsvkNil5g9npm1Gm8gOZH05S5cM5XA
zcIjQwIBAOokG1zswRw0no+WUYToKnL/QbS87ANNWD1WSoqQa98xATlxAbcUoqJ6xZeOh0Cya1KH
EWZrUpmQdSBDRTAy6fLedN9e4JkHeviw1suvRRAXvhLKQs1zUo+MGO/7EFEg3S206vs1e9lKS1Dd
5ckub/GzISqk89oIjKruEK8nWx4y9ibu/BnCV8dRNHjAx7Bbh+h/S/DdLtUB9aqR83pPMXN6LNmO
xYhALYoKPnwHWlu2PP4ydi6hd7Tn50t8cFOAnr6yXM71jgexMVuCebNSsCgsDV+1tYYcnDLWbeCm
Efrj8M2g7TFkWZBBWdJWIwuPUw8b5UF4t99EGDdv0gDFGs0lOaHIqfY98+3Qbj4puJGVHTGNEbSG
Clfu/HiMWKJ82ov6fKAQLJmrCVJ5HONybiEH4Hd+AxBNIeJWnEzvb+TgjJ5Pz+FWf0vyk16e76rG
j0RNRkTRIrSkoKe4zSE84Ni46JIOEW0LJgc6et/g88zDTNjqKOEbabGmo64MHHCqHbs/9Kaq2vkh
XoFQhF7/zo6oo5xvLt2WnEOFTWP8qgPJ6LrKJBec4x1P7urOqT8GItUew94a/llrm890zniEb/oj
0g127cUJPlq4JmZGWurybmoXNNe9pM57hgRVu0ifz7Mva9YrGFiq6uWIBL9W56ZcttTwuQ1Ck5fy
wCULDjsdQPfw1gL9fxXiJEWkCl8Cga3st6b9kctdrTUfyctUxQKE6XOVd33TUXqKIXcPJQc+TDw2
9rvv2pt1N8GmQFuB8H1cfgXUCnPRqL0gjYum78CU3936rF/cfWFlzrRw54ZwpVoKKfPuXtoHvzkr
7D2pKrPXvdaL5ABD+HOKcYiU/VDrJm5B55siZ8W/VflMOjmWzaM3XL9zUMtH2q/+O2wA8tXVAyNi
lp//htYML1uNRqHOjNM7TkyZSXYK88Mq7ENva0yZgnxxDY/tx8x1l8ZotkqUFBsLvmXlOelJdsUe
qwVTVmFTqrd5gBF2lW60CKlqU372JK8tSNwEnfLfc/+mSw4hiiYP4YaV048xYqpFqDpsMVueH7I5
hmDEPicykBW9mS43f7/uQuf8MGqtwqMAMTW8QUv7L/FIluw3jt4ieL0Wf5qI0X7l+xn7KoXXDu8s
pUgSUhrAdmxMz3dRWUAvqzLAKHWYjyv6G4QuEYtqYXdrKWuVDizjWiBTpuo1oR0kjRcdoBGZTc8D
quE52NM+3p0hhuu+vXBqolU04RAS3UbfhK4CkRcXUm8DYycg64gq6IXn8EhBd+SITv122v4EJkPI
roWsv2aftGQgSeyuKGH+B7Nz9Wu5EwWKEB3lrYFp8bXMJy0QmUph9XDAaDbkeSWQ9WYygQN9mMnG
PrCt2T4MBayGlqWL3Mol09H6mCteW1gKjRm2bjTbAytr2n5YSvlIRuhCkzH0s6rw5koSRkgV50xk
zLXw3GuCSoF4HRvpn6foVotYFBaP08n7NP3kR1ME3xnzu3u0IZM9hCGLxY5wyviwH8Gt4gJnzg/G
Ng/ZHab1HJVMipk1MeSwz+yuLqLZ1qEwpEfDDqHPKnw5YXQ3tvY4EgJcHRUXvZMmGsOO/Tv3LJwG
+Xx1UCcVyqAVe6XlESFN/13/w57f8GcG0TUbmF2dLZGtDJ+zTb4qvkXY8+dT6eWWecAsZwM74PWb
JSRGUt9jtPWPOH796SXeKi8Vi6Cylpx4ChlcxygKaA3oMLXemPMy4RJwgmI0YG0vdkJi/l1+8MNU
noYNp9FVI/e7ceXdKuTpyyV59VfllKQmIb9N5jCuaOZuLLCadABDe7uCKK+Sx4YtABhSsRf0FuNZ
XPgishYnOkPuUk7Aolf5G77yCPFqAwciDL8OIAnAd0yHWy6eK5doaQfAVw6JeL4qT/xbGqXV9l2r
vwcGo81xsund/6uo60uzxiyXSP9Lj3Bd6HdUgeBJjKRH+pRxJv908n4BthZyJveLp1SjbOSJQhAV
mVQqJzt3PepTw3p5lqQ8vZaH//0Il1kEpYqZUThqqhv4mm0JEIkmUb/JmynIi6jtOIGr5rdULkcE
NJqzUTZI/QkCMalAzaOpyVNDXgG0AtXkQ+nBHbq7KHgv0soSUzWsClREnRJPmMhkUsqUzXj4ebhw
f/iyK8iB4F6xU/eoLfjs+4KA9MI+btTn/Do8CW1JQMAYCKznszyPc6jNQh6sSikm4IP1yMI1wjox
KRCkSAA+E0YpgjE2jp055cVrlQbl8K/AfinTKQRXiZ0kuslb8cvgQnat0P+GPwc+wXHaSdtILMxw
C3rAQgW/n5tiP0OsZjKtDYG1gLtkMC86VTNlFbgC2EzWBXmJjQklo31BHpMmCRFwNz5Tam/SjzUv
2kSMbZYoGIu6e/avHUrt0WZw9K9QcPM5IZ/RroLBIZlBd5waQ0dFyFFxE8oFBocNYDAg3/LcxVK3
LSbrY+KZOifx4d4bf7sGZ7NUGyWNtN6qLDtloEsVZBQPuUYpMzihljiVUQEPH/6CVkrADDKhaegq
ybmHyAtTS0mbvFcnfDM29nrLF89YvLIob06s7viWWXL4cEOHgI84/KD0A9BhHK1JPNBcf5ekmy5i
y1xqkJ6tub1tiGU0GuZG3s62VMvNC47dp5IvICr9wJsj1PHJ6V5CKmQl95mjEcJbJSb2U7s35m8X
VMh76h7yL1wTgBctpkJOW1lGnzNttENJwzXwIC9TXjgVW3nTAn7WrE7T710nLc+boZZnii9cHtMf
4CpnT2B2+fP6j8Un5791xvvksvo2AZlmJnkOaJwpbkAgBoxpAAmqwcpaEnlgaPQj9f0p1PkUSofd
oNn1nLtbW8r2TPyKcjvmI/IZKJrsusu5gXlQhvb3gUjXR4QyegxX2mQudJG1Bt8brFjit2RAD+rU
DU9AuS+UHIHMZqD7YicG/T710LirXzQ6RnTuNALpjtNAqwa+Zlb6KGZQtndvF1SUIHOiVyqeLzFQ
AKQ6X53SkuaxP1O8QvgFYoXoxu4oN1sEg/lzoM6Siyvu/Xd+y0rTdFJ75si2EQtwnZGaoxz9Lkoj
W7GMlPMd+hYnphyoHAjUnwpbnCrNq61d3QVq//qgelX3gi3sDmtpKrZiFt83R59+J6QQMn6bQMib
KfXSfSRtxsBHroz2oROSioOIX+ZqDMKNNBF+ZPea2B/qyvqZB8s05e25QIP7a37kIgNHabU9VcuF
Odhn/gpxPlsNOPlmWnid6lkmRh/I6jTBryykVWhnAx6FAqpU7lRCIh2pwna6T42ALX09rxmkLYte
sFXCgxDampPgxjPaINYQQcXLRL1DMWFoc250/obYqSla14FZ4mWuPwVigtDWmYiKRlhYUg+ID8df
9OLHfp8BP48h+EoqdBYDX7px+SF+IFzVvR/E5TVfd1mcv3jR55vdIraRCCMO2J15aCiKdmGOBuuW
iThUFB023Ja4mHNxIvQeVqrmYKU7vltjKsdmXe2DfxR0yO9faWH1whvrtKSZcegkYjGuJKMiA4uF
bJXHAccObCOBJCb1gosgwXI5S5DTHHCKRUWGepcQ5DHhrReTY82DCiwo9fgNeLJC5glvCJsd6tWJ
nkaAKqA/mGRRH7ADatUz/PIPrdn+lO9ycIVDg2crwtbQokAGVexl7WELEL2pgN4JfOqeZG9ruE6+
kQglQP3BjLXSg6EFVMsl5kZaGFgkZorTdOtprEt0RH2tBwfkMyJIL/Z+e8AYur6DqxytwN0CnX4P
mHuRBrfwusHELhUJ77rCaIbXAxqIWKTpyTgLW8XQCIGF4WDz26ICAx807OY4kkk4e3BbMkk/9Vn/
+KE9uKZBzf6alkgq/3cb78a+1EqaFDbv/dr4J3gH94aOh+2vIT5Lu1UJMuTbPgQ6KG8y0dOXWDjP
0SKuYkxb6jTmAHIXdws3Rk+tLqKkxA+9PQQZr8ZvtWpdpI6CjbioWieARCnPBasbEQLgirRIrU+Q
IcEFZn3YxVqCDvW/z2kjvPVZj7WcYJYcwRrqjS3DXTWf0EY92ZSayT2FAh2fNRxscZysSgg5Ij0B
bSZZ2b649ja3zqoysR/EV66mw1X6cvIFcnjDuhHUnYn5Eq3LA8hhJ1kg95CGidyZBZ7gskA+eINk
o45UvYf5zv292aRCbKJnvLdD07SPgqx+KKMz2KA/nwaN2T3uv5RE4agT7OjoFIQ0oeAlztZiWohc
VIZQWUz9O9IqhMXhAIxYN5bsoCkAZ1haWwcMMOP7vo98BofWnIGMbk04mgc89LSmpHuVzqDvmSsd
eIqcbCeXuVGinz79KR+nmNkahBoYVNcPt6DL4PuFNap9x21oyx++TIb+pTz52KIVyos77ji3MQKd
SGRrbVOOLF836gu8R58dtYwHWq1uxgD3OmP0zkmEd9yNNfJPI8wiPezgJVmYiA2H34tpYXxpa7Na
aHBoBXZBqbbErJIp2ULYtXWT90rtGVZRud+tSO18nZNL36DKEJbzhMMRk7spflrE53VkcBGoexoA
cWHm6gA+mvpQbL4hSDzOgOZRVYuwLLIZrDzhisUfGfEZVX5MWD4nAXnhbM9YdmafQO7Sqr2zq7lT
gf5UHgdhM5MLLWY2TWbc7VnEPaswh/Zqq769VoNyn3wbXlyHZQ7vcxSph3rd3pLDeCK25cJmjERX
wdBFjR8O1Mzpd0f9ml0aMY4xOQ4UyXH01e6Kk2G3fJWUckmiPZSVDsCgbg9/aXTLckKYE9T59bai
pTUV0+ibVVrr2hxK2f6Xf4LFBopV0tDMDLe2lrDSVhOttMHK3K+GYPJqzdXJYQiuNMzgkmAsDVk4
9q/nPXMtA/XwHrsMQHCpWCtSA8JrdBIi0ZlQivraCo61qSiqNAghs3vQXvayeoOk1u9JSJX5Z6iX
Fg15mFaJlYBdBXwU48a4TxQcTad8aPAa3aHNUekkDlOv1jDiFXgHTchTvdblMFSebFtx9Blk/0wL
BmnNA+XCQC+oX3LDGWLGPTnOPRBUYdHbV2S3uBT/Pbt/e16KcYiUYuJMr9BFL0lJSxkGdgUXzVxc
TzWpRKFn/d3zwRCLAMUyaNGw28s6fKCERFsyI8uadMeGi+u9zHd0rhy1J0Usa4FAypfEA2ZJYfWZ
O79WHWqk+Hpwb+HNZFSwWQhFO8PJWiHW2mwfBJK+MKice1IN0dU5YZt3+bmRoQ3r1yMKunG9LMs6
pJ56tJ1bdt1r+e9kr1vZ2zyoj96ETJbw8yLKzr9BTZ9gS/B3+6hQYI4IfKyldzXpzxOaKP8UI76y
99VqPmStwvuc7OyBxLcKntK0iivN3xdEnRg7cI+Hn9sLs4hzsrV3KzDXGEaGmc67Eg/SXpRkH2UM
RDMBw8PCzH9FQHiD8e0/jfx1pkF8jKKcOkDVk99Zqgvgv3yFvGYYDV0dZhJSmk3g0nJFTVbMHdGH
vGLoctCa4h1K9UHD+sRnVQuXtoXFkXJW3iD224Nd6MXwb6qiPO+lzxRcWfcaUxHVdzpgjZfgWv0L
UG6jx9Fyr+BOLJbs7UAQUMQ/m+y6pVZ2TsKUxsMvGCNXRRjljyUvMDlWNFt+hFrZSWIIy/Q0NnnZ
QwWq+FGNI9lSdAOeOxxUvJDfmLHTiG1RUnNHrZvvZEyjbMuj3k4C8zWWFkqjFFbxsVidCdUsp+Uk
ApnnkxRs0X3Tn+6DQ5pygkVDIHb8hX1ePCXZOcI8TrnhS8QPRlxldQuN+SoQsqszXu65CxLTh0ZL
tA6oXubIdGAHq22/ITzcYOYeVxLLlUez1TuSvU6iJf8mGxOCFZFnN4fVzfW0iUtd1DQRQJCZkhnu
tTblfM8jJI9jWlS5cFTujt8AOeCZ6v+UZbFu6RBZ2CSGoaVkpDSsuhwfJ7sv4avaShsAxrGKH/j8
yePfTYLYQruBiNK7NLSAbGoqzu4A6Yci6Tn9G8IrXhhFk5RSn0kr28NNlZShoPhgtsVc9UYxcM5A
DAsve7qDGrpqA3Mx9zJL5zYJKx0uU7GBnhERxidNutKtVto7V9xRKmv0LGmICFQB6yt/fWp96+mo
C/r2wxA927WsiDlbiHNQku8HRGMeZkvKWquQ2LA5OH8D6uAQtW8zN1+xLS94bcc43YWVy3oXzvKd
/5T/VjNZ9ejOKD4QjR7NhsoxjLOwnz4GyYkwxAN9Gqn5TUyVigWcFV/1V6QFKt9a5CpOzyLzB5+E
KUTyFIIGaeD/R9TDIsuogFfHnzIQDV5zrXstfQAU9eUVcW0yer1aQN4drn080eYsyg8xKcxv8x2g
sjcwB/1xBMCE9q5c6+nADdR1qLdwhdbKZajh8AvL2k7jTuAdRjWREG+nPZT/shobhpoM9mqqzXrP
BkMfVxsoYlsXAkO1fSsiczWb7VM6fKZV36OwjQVDecQz7k1AFa4JgCaP15DDQ4OortsvsNl+y6nD
ULkRf1t7VsD9uMgTfj1qVsXXd9AIA8j188c/BRDaY6eOqzw4RTFLA3gs2+rNhScFZrjnz/hSag06
WYzBN8kFLNYQ+uQt8QVmztuvP2m8mrortsaeb8mVJbTrOK5Efr4tttiX/q0C9WF8TfF7dXSX+SDf
5pQMTGG3ZpoTK+6+NDCcKew9C3LpOc5/tXV+5UnXAHCS3Fxn2ND3UT0CROpJcJu/n5oHHfDJs9oh
uZa0Xzd2ScpADWYCy1S/8orpzwSQDW7Nu8e/V3Zbn3lqO4CNZefGteS3UiwGQkekJp44IB33RJDr
oRHBxOKu1fHdl+SmTm2kqpdBENSEYTzU77G6FBmbWtdNPaAgP+uauYBUdscWBOcKHvoQHPm6a0ig
XcQAyMxTtyhwdnYF1c8fbw2G0pER7VXOA3a0vR52q/0D241LAmUB/lFF0TDg5GTLpfuNyC4flDJu
DkXlZG4HWK1vVoYD2JPuRpZQgUyO2vPMIwj9qFZ1ua0hw0SCmFG01vJQla3tE7mStQaYC89EXLCL
nsSdl0WkOeNGIxuqEPZh2BXuWTEW9l+6QCF3Ua5B3cDvJyZFLYzOgbRIq+s35efF/XqkXK2uKe7E
IzosMImsKZL3e4P3OnxESHqw3yS2F8JkAXTJbpXlrE5zi6uIDgjo0JJ8XeopS8Nvj++BmRybrl9u
Z3xnM+OwwhAL3uivfl9w/icZ/b7Ak22qA43YJpZiSfxn3G8xA1GBmLOHpu2coZ8tua/ptnjvc9kO
9364FW8octZzYDwkUc2KrgI0zyjHTT+k/7S7F+jPNk1DRSFR7+PTwIzXuD7lFUIzMe1y9e16okBP
Uh9Fj7yefpv1KUgAFs+7h6yxQFme88jyEz9awRRhzpFkq4aSN+w/+e6xTeZR6tmnFC7MyQ2qVSp8
fOWjnxQ2K8Ci8gKiTa8sxY00GFA3e5L9L0ykD16hCsvT7UgghzHNys+RfBcBHvDs7upxc291fJ2v
SPwokivjtpbG5JYbP8oq7oJhVfH83aWGLIlKPb20yo3Qp4fgCIX8vIfgUKWSjK6KwdAeV4+DaA65
RRhncEcfYxfk7S+t2dlDHw5dC2pgPtUPgU4MqFSd9eDOuIkwEmWn25FAxOFCMd2HUpKv5FKsWhrG
1y0fjqH3+ToL/FrRr7YU/SEazl9GWqGCoFvqsdGU8WdSvC1d/HE6cVMxbBCyNiPIF13ReF3BBvo3
sCW8pSkfK5R3vDEtJY6zrrOJFPfgg9JFp2HtlB3RFQyE+rOytHqTYI+Ax+4d+yencGJ/llThLE8x
WvCxNDOHlSmiv/f2k69cmbcH9IiMrF8F5VmsFjOtPgbKQ/z3hEcT0jp22qWLm9zaGJRbCJUcLPD6
tdRDXaGlRW54KjJFLa8gCECv9mCwn7Sn4QvyUKMYC0YzxFSKK/z72+XfkLA3E8iTZOU3LFaMbUTP
WKukXlTaGkll3RYOnYJjAMFCHweFMFeJz/TgxsYNyxd5cOBqvtFKEEXDcTkIUrX8iWU4/LQLQtfX
6XH3B1eaXayvw7HyxvToAKG+ZKF534tdZaOtlLBQw1Eal4sj3parM+RNoLyoTRpWrzSzu+ocOxrW
9fEjYhruWmIwAB+m4Ehwp/K/kDQFloMrvXhbiP50XBupNGw7yjNLJO67C8877eN6q3wTljKhE4xV
I+I/MNMFKOq/c/TOcpotK00c3YY226U0aaL4XEQPraqUWXyfC7dQEDKOs+tYVHc36cwNoRI6XAxO
hWnDlFRvbOEuT0MIRvcY+5HEbCJyvi3YtWg/EZxZhdco6NQhR/UfBzrdsTfuRVcegMofk0LDxGUf
OEJa1JjE2huJAK6f0N05jhFF41e4jOukSewCcsdx0NW4zDMtsKDIuahQzW25b+XTc+MfTsLL8877
YqQcJNoe/qM3Hu9uc8Qq0k7iPTzqq+U+stL5Ny1njRZP6SfgkfhJqkml65RhOroKEb14PgXqxrXQ
cJbJyKaIVEjv4wEOo5R5Vo24XG01DP2q4B+vN5zYpFgMwbxxXbWfNidgWT0lQzFSD1Yg9ofR02mu
HkJJr6BEZXqDY4NXGQ1fueviCJktV4uh8JFO4OjpfD/oRjUXDCkiNNxlUG9aB+7w4h3bLGrARVWY
h1OtcojVo6DhJrSONCqnMqOGL9++BAqVBBsxHw3gbrtB+IbzCJLFHfkEpA6rnTSzwUsfOPVp3Nzk
+OBdeO1z63b1g+T+RUwwRt6NtHD8xMQ6QMs61EOgGlSN7zz+nXg/0hYNRMhLPMxJ0moe9YykDO34
umyi36R/nEVIVPFyQd/PsGS/NuNLoGcL+b07zIHUofDG7gp43desvvpmpYmwsId1ui40n7UjglCo
ksE4TS9EeIDIuD0sdhpBdPsip1Ga9kPmuGbAILdARMGcyGJKv+Byw8yMpa5hyXCVuF8NDtSP498N
faiuyDO/QQc1W01nnTuHsdQuvF7wkoZu1tfc49aepcjQcsbugvFVRLTOeMLXV/w2Z415k+Y+ozok
8H7+ErjLKTETLr2Hwgfo3Dfwtq6mEOJSSrOqm5v+drHun6YOQwpgVDhxUhRnY8QnFPilJ6YD+OJo
gAE2llZnPkrOAPwSzlKRfaYceo9hPOnvZk7/Sn66Ap5DH40XHBZqH8ZbHTso9SUFd+SUHMIB2kON
kjrd4Mzm2iP3qFEftS2peRfmmuyDIvsdM7N/Y58STce5TCZPPPBTlOG0Jcz7rrzJhDEuPSXXY0Ba
F4Z6gfyps6Z30fHEItd/QrWEHvUf9Y3MEFEd5dz4PrShoKIp3Y7osQ9TXdXekDhfcXxeTqWZ8LVg
49cwoTMSQ0/WJkT1+vaZzKEHQpXVtMYj6S5WnrWpeyfS050tBkECnxnLTDC+4nZQ8HHAfAFvt54S
KEEYL21SlOYHzAb+pkeO3cAmJsqOoEgHGr+YC/vRqB5qqXFwD/lQ2c0KUW9TasoEVerkBtjkdlpd
2CdDV4Vwr6bVCk83DIJElVX2OL84jeUHRbIJpNKMSar2dsz1IU9jgJ5sONmIS4+AZUK4EGPq9TTh
xUotzWtlbpFKRrwAvOs/zZCKw0YTmW2E0xJew+ZcxvZeksCRTt+5BcLxBjHaR+UugzykHC33vnXJ
IH5fd60A2F27kuP3tn6ysBftly9rmMB5ryuSsE1C5uEBj2kjvSoy05NADNQ/0QU0MQa19XS8KpZi
EZOFIdf35Y9G0VTnWjTCo2ES2t1219cFzri45IRNoC4K0dDRj3pdEpw760VSt/7+OW+JI4MD7J+E
n7nbEnPZshp9JZhKsksvnyy6OL55BCfIju/tL4AO+1V8pltoLiYYuTafv47REOshp83jawcKQo+7
4gurtjTy1IPHElzOUlI+V/YAvLNNDmvjj0Ez1vfRA9QftZ/R7pYMkA5wRhq2JE7LrQJHgAV9PIad
ZrMbYvLSWIhQT4vUypGbLLSA9bmc8olEw2M+9wgxDnjjTUADzcyxGzhr3zls/n0q84KYnIZSE3bQ
q8rnfpZzBVQM6B1vwEp0vfxcx349RNwQ0UjUqj66YbpJe+IVIEGrhDrPIDd3AlrSQ6i+Jkz9JsXy
2TXrnMFswwg19GxQpncmX3FEZ//GCt8pFZXLe5EtoJcvvTBl6JFeR5jMAv7eXQ/dN8+D8Sh82RJK
VeQck3vPyrKgcWotkpc5QmQXTM1XN4fDtHocN/p3PN9IZZCywsM/vPaRPxgN3Bo4hRmnxCLSXsd2
h0POnp935aoa8Q0h+kHWYjYuv89Z3v4EZ5o1b/JHloa9bkurdkPoYRnrg/h9IIDkhnMKriGR54JR
O03vzLP/1y/aqBvDaeI9IlkDRXjhHJM613Gc99nvAypf6mBe3/u75k4riUZcC1jGjKe6NWFKDl6U
wquwJshnWws4Y5KGx5rSkIJnsPnvK5/JiuglmvzXlHoalXGNTrPc4lhKlDagGbAPjjehNU3YMhYs
PRjcr6Ftwxr+NR90dJpl3klzdrHDnu/UNv+Ir3RTCHjcREIS7/1UyjH3wyIqqQ4oOctG7lP5+azQ
V1Nr0zMlRBdLvtoGUjWoX4TGa0BG5rQXLR9hTEpA0ZpYCoPStCVEO1UlEg4938rOypSNaXPInQP1
ZNmlgBRj/uOeSNZxUi7emSbHy7dWIhV8T8fydbZEM4jgbntsJsCJTfI+IRUfKhRi5wW+qiUpFMIX
wXX7zaegpbwtjO5oDfG2sQtO09qinaxesS2E60g0LA+JZ8tPeuiHHsusLcn/3W1hDa5t4xIiHs7q
cpqL1UONqtaKNyvhKzKaXAWeTeETdTfCgkT1RQxFPCdTVgn4TkGT7eoizKX3HNjAr7ZeoWluB3jx
nMvLuxCqQDGGlZANFgLNN8gf5uudZtta4rXzrKdbCrA94mZlAExHGiIY5SF/EiYX9rSl5t0V/Un5
7WjyOF79a0lOx+BcZtAz5xyGPZJR4nStykTenVZ7ri4BXOCWhyYgxfD8RYjQP8q8TYgHOZNZ766d
ovbj35bk8/4RRtFmrzyD3ZtFTIC/S+OWC4DnIAZDLjUv8pNzv4F5wPD49/oqMItjg9obGtHCUkbv
IrnkuDnw6pYhJVSF73LTAy9L4iSkHua3GXtBbq1HubtEuMN1aG1n0u8mNw6DhHTdiLMos5mxr4wm
KIodm0+W5hyzhxoTTRXrJzpS5kcKVonsL39h7RX3ivnGqFWbCfAP7TWbDCYxELy7ljD/Cm/W7r7E
x25FzYRBw2xQnOFxL8Jk36FMwKqVqMzjsuebdGJepw2p2QkTonotG6ek5IZKifHsEZjDgITKDuUM
MmgoTtloYMlDQBWAdjy4G1zs9nDqFtcxShuZd9+Wyr/ftEGZd/aiyvLYLIk6L34yRphrlozr3FdT
4bY1yogZN9JFCKihNtK9dnUo92x9N4/uXk3oAhkiXPj3JxD0MRWyWXv2I67dghowxEsE6lCSyKB2
0wwTaDhIXmbnpbZp2S19tFlQ50LRnvKaPYrx8fCHDwDaVUj9jqb/b4O+IlaR4z7Ezw20BCsyDkK2
00JYlV7KN+J79Ht1NFKwdt92t/YRnRwx9/9doSZMi+DlTaOkR8vTcyGVNPKtMq8xS5iBJAbILepB
gWblHVi4UzUomKCPZQxejhZ2Trnfs1ozo2SvbnWUCWA5ZVnVIaXfnJkS3KyvXtDSz0zin+CSI9wG
/8qY1+XICQ7pk6eOJEEgHQ4ocpgQCeUL5+cdWBaieMQInvg63fchR5jMUupa6whCce/L/KUQptMD
R9jPiJnvN/lGFA/4MKQH+jXxW7JaIUXrez2NJD0h+c7SDf9Dq/96xjaGjl5Ud1LifC1o7e3N4c0w
1a6bFX2x4JRNdUEkbcLWof3ZuAqrawBYw06y2sEHruMWjjJYn33Xgs6SCRgPf5dgUYRcxJgSQqH8
G1c3kezFvJcn66eAaqirpEM0IB1NsfWreka+2tjTDNBRdqRI2RlYKWYBC3U8d9qoQUlpCDG0+aDN
MQLMoDNXlJzv7OZNejH55edUMYkxJ1XZ38yeIdnhlKiSUoyVq4OHkznot1sccWf7R8OVdHzLIKBT
vrWpk20MaZaoac0ZP3AZx1NNGWHBeKDFhOKXPhZepKxgb0eWe1w7k0g7bKlpLN0SkJdbmUS8MDp8
jCkr2jPDYbP0faPApb4jyccBTwU0I9H22m0fRtvqRQqNPxK8ON211bl9Cq4AN1hxXq827MGw0c9f
C0cKqOWsTpCPBSieyvQ2w40dIyJjJzpnYqv9nwHKa6CLURUjc5bdp0bAYMDw8lEq9ajuUpE2K4Ni
Rg3pDm6dJxrhmVsY1BKWcrIdU0GUIiDZL2/0a0G9W3TXB6Xl9Kd7pd6zdCFfAM0s/xt1nHXwI/lx
21Tl0fKyjKAFahZ9YB17LxS3X0ZxM9NpXH3T9TKglJVzb2mN0EYdd6yix1cx+bgsTG3R6RyPATAE
KxtVvxWvhiIvtDMV0WquaS4g3p2b18T0dhofUu3+eztWrtpXRjQxOTrDz0wLScNw0zaCXzVn5bBV
S1qCWTzz4a2kq1tl93PYcz8wHwe8rbR1mXFW/NVzFdW/0LFm7cEPvXVZD97ZPvVzf1PXjogBVZUM
ReVsBUBjQSNeI6D/SC0CYRiYjQIST461jjmrepBBZZ+95GZwEkGVDkB6RxIHpuPlAt49vi5i0pp5
EXoCLuhJ01p5SDXWVKr99n77ti99+7ry/zUxBWEhZN9i3MhDvIcAkVjuh4kg/qUnuZib3oxTiojk
7qkkwCL/rWkmuOJ1IPkacYSE4qz4MJjeQogiHtP8Jy2xIuv485p878x3wsjNf5EYuokVc6SwIUgg
6voK+/noB7QVypBUQdiIlk3AJfqBOUEsrQW8TEgo/EcNVdh9Y0NHXjbMp3/7+xvjiDubIE6ph7Ec
rEEDoIyp4IaJZYYjYwhscL2T6aIwWZGOViTVzAjcU00JmC4FUfV54P0iihvmkRGIUyIUFYpEh52J
nP8aMv3S6b+llneC8LhXUfhzowUDUIfr6TJovrVsSN+YcdyvIu9GQE1XWiMP8b+5fc3iGgGSNdjq
MH9u8SKEjTFu2FNOdOWC8xzL5g9Q7ygwaA5rnTm4F5uXsPOh4JeWxU/GmjJK6BRvRkBHznkopxa7
jo3A4jY8tzLqXbPQ4q/nqSgWelYeC65lHv6xqAxhEJcM7zo97wKIdtBiR6hANQgw5S4YNzaEqED/
WdhKVYOpwr4Mx/j760D/Xnkn97xtiK6X2UAp310CWiIwH7k55CO1Wak2Vn5M4Vkld51brCdHwjjm
rj2k5uq69M/jkQ0nBE01Bx8HqRrI+Gnm/rDRH3FppZ3sfI77pPY9/N6e/TwvHDTlgRD2jejrMbnk
BZsnm/JMkeU7HVgkAqSdoLZoHf25J/PXdRL+n/5pSvDUHeT/yNdnVqCJYvYxNPtCp/uAFuCk74nI
e/Rjj3uoTe39/uhVbOBRVsCpn2/fZ39TPEVDOiywJ7ksnWXnGBqOMo4EyYQVXZwRyLPPMJ6JH2S5
c+6v0XANrmnIuynxfNMknXlr3WL2RZlZeo0+N62+rGezbS/1pL5wt38i5ynjPiMFMzeTneRxW5s7
3Tq1VPee9J95X+mnOHZRolwKeeXMm9RmmMmnpThmltiRrP2apW+3ctFCOqnE6SYoNvYAeO51XCwD
Fm4h4rhWcvfaMWYGP+d5kViPv+Svh7+21QL0sfIh3XY15fpGCA60nn3c8p5ScNFn/p4jhaFpQZ3V
ViMl8KlhWnv1hKmdtFlpE5Gyikf1PoAMG5k6RLc6OCvPf37veeSBHKri78PECTnDrCS+hlWLvlx1
EKdOQrfAkDeskFWGAj4ECDaE6fQXHKcPcSRQzWRv42WTBtIsAsEfmxyH8/jbZLwjeDxTk3EQaZDo
nvmlIyMkXuysOLZzZbe3N4ijNxcJa7g9NnVKjoBlXoUMX7j6H/OtXd2LG/rjgqNlK2JkIkyqRdFY
BKyJv9hw6aKMlF3iqk7TxJZag8pHQwIg3PL6aDFxBMX3nkCyOgTR/SbK19PoZHQ3v+IbOFVBAjYS
PMLn5Hp0WfJcNB8KBoddNS2ZC2upDhium3oB8vG7Y7HQF5VTbIhmoBRTXcLEFD56fMpYTfKRRihj
f5Bsh5HcF8afoF+EU5yF2Qu3MQkD9b4QiQUE4d5Ch3uAkKDtLsgXV8Ws8akkSyhJ7Wx0A74JKalD
7el6gi87xHdiohHUworexNGoXUmEXDLpzsxkZOmnkALjG5jD/xVnDcbd29JK1ujJJFNtEue6KI7h
yFlBtYHzJgadNJd5wuHv72WsffjfgLNPMVXbd9bC+5h3jMF5hi2VBrFAapT3N35QNlF6NV9RL1zl
zp1T4QCnhwDBoiPQDrQiKJL+ooWhOK1n2/6FjOZ3h/3GU+cxeBM9KUGWyK87Dk8sBtPLl5BYx83q
nDB42ZpaGtDUIqJxdGC9yuNNByMGpUvHP++dia6F0d9liott2qpQeE/YrlagYcHfjvz37MWf/xMh
xoa8q9gD0KtMJ+v16QErJAP1fDK7WUR5eYSlLsTBIz779hg07kWqmJ6GeAm0z3xqvQ1V3WXC/FfY
gYA7c0Pukv2Lx3nvUG7IDzkhTcQzOtlyE6uQkTtX3VtMvTglC7quHc3nLQcfndonpXbtPALjNfcI
ROb+zCLiUioGjyQ4o9I71rkyvwKX6V2YcvBHiYX95Ia2QunzyHT81I6qV/mOK9aquuLQ1qhdmWCA
uvpaLz2m8TniqLIfJuo+0xjU6+DO1X8ZNFgN4dKdxlmew0I2Y9jmT3LZnwYmLx06+flRrmwiGdf4
hct/PFeEkgRBy4iIbhaMYW9K7UqBsr7a3tKmWyRtOZWjamFYOdrwpMfYflyvkfvQFlr9Nw8TxXHd
aSWbC280vHdbBmpQET2Ust4x56pbjfoRdvZOncQEHUbID3gwYja5hxeq5fODhFXjc9EHxLDWvZhP
37Qd43df5GtWB+yMvoKZB+/kfKLwdHJsmagXxPU+ICAndDsAopC1M5zatAK19XKm+aNJtNtmSVx9
mRsKmkMYjbftnU2ERCBqmjchL48Rj/v7UmNruGZ/NXG2rdLVEoed58wVwAKz/M2N1JT09tikrSbG
oMOJemIoudmr5gp+cWjSwg71bfXXSBlsB/lZ+riENxQGsg2Ob0ME9MpnMwt24Zi/L5M45+R7fPQ7
hZTUQjiXzBNy4DE7HEhR5PeIiL+zgdZKAIRf+c8+8R+V1745d1oAV9VsdoasmW8GqUO1OVczJlen
okkWQGs3LWkH5WADpjnfezlTbFLl/VcxkbeHJD+stl+i/TrOlAUx5/BzlNpay6bj3lsUlQHKKOsU
H+sXPRkNaq5JYkRxR3JGSgnMxX49VncFZY57dtkxOq7eTsfzyncu6uvektgI1GSeF1xZWUKcVBH5
48ngNh4Pvh6+bBct/FmtpZlJ/3PIo5nnjFep9dYFfZ41QpyMHIhLDcTxEzMDf9Y22R9Yh3I4Mp/U
+7RXm4q09D/CanRMPShsAaSFY85Vqmf4DPmzOCwnOKxevSo/NrjJjD1zs3GMJl17iyq1od3kBNrs
pIAw2hdWfj1rd+/QRpQrF44oA0KsIxCyqnGULtfbXxEBhiKIvgqkB/5YVfTL79Jrqt+fcTtXuSr5
N8sMLQqeyJVLcuEXhI464MS6i9oEKUMLUDO6NSFb3sfP4mYKRmnVCUG1/abWQ1CWFwcKoy2vWEcZ
ZcSfL/r4vfLzmQGnA8jQUoaoNHb1MOg/eI3LSirZHNzXAZ4/uD4LHsuZDgkOCPuUiJhvTCggwwhZ
MrHREikr7A4I5CKZJk/zTNtE/7vF2ni185vucEsHkUSZ3ebhORevXJafycfGiFxL6a494cep97G6
DF00rJrMRSv98k+E6vGmk/nVCcD4vAchzE5kC6BYCkbGSEYgPTkZDdPKMv7ddi4TLZ2oVXTQ76kt
5Ce8G87pPedvKpDSfAoD5mLqDW0xOxre0o5IUlyF+Cd3695jFTb106z8ulRbAX2SvY1NDQl9f+l4
RqN9Y9c6xYe94u6g/HqKzfpru3A3i0Fkgke6k+zCSke6idi1sfrcCa1Rkcmy9D1FyyY1HFLuqQ0k
JpxsVIwufvcEDVI6MbtEnEZlHqJaujg4l42zWlMN3SJEGNpnm8w7ctGV7xgaoJwVkRj0YmESyVO4
nJLPShnsli5v5r7L6bcLZFjbA1JrE6ZoupTkCOxk6km8oHIQNX9uHbjGniY3arvMqtZfw/3z/NKU
x0q9Rl4LuTkBxK/U1p0BfdO5+xf9tKIwcsqABPQDtGwyo5p7QAIrQeXVC0GDfPGYrqtUrHaBDfqc
TN1ZZJSLVz1ow0mghBgC0UXP3bfcLve40aye6Tmvh12PTfcRYKiqoMfK1qkm73KC98scHK3Ismy+
0wOdBSmmREPO2SiozdVKdbO+o4Y5cjzpG/d0g7vZR4oH6lfv3iQmUWuD8dV9xHmmWpV95lv+8K2k
5nIZ8Sf7ur7+MbWS9SgKezhKc0uMKwjvgc8f8SlQEjt6+v4oCw+9dhzscu7/Ow4JFa3ajKlvJCFI
WF3+ADIN8NcSfWozNpQqnpDknoydPPlFUQlGqIDN8PAsBCYQvYCg+NYbnTWcEQ6z1cNlqZmegO5O
bKU5JDoMSydLahG/iA7UzqMYFA5PrOkuPn1ANfzbNJDDmA4fG2M6qjauet4B8e69W06UkLc26beY
6an8GQ75/luUOGE55RUrcucNBl2Rd7MP9NOk+m4Lx26Qf7q5gno7vkmuxDSfvvv5yKgUgeQrxuVq
iPey8btGWacqa/oM4xTB3uLxUMqllwIqATsKimpvXo2pVgL66LAVzL5bAQAs5TWXfIWUOn10tw6E
r0jSWVhU/BZgthVYJzuASPBgDft4vSjttwXdMf6RVofgwiTpxvAkOI2QrLqn8VkPNDJBgWL5QTUR
c5iyJs5Qxo2C8mfYEY0BKmA3nSsfBTiPRKNvVQR1WufK0ZrUqn8Gr+pPSdPAtlyIr3l7pcpdatN1
q71ckA4Kviau7A5oT2tVr941yROOgP6hj957SaULC+kB2mSVpxy+I+wC1XUGbUI8BAt2WoYRJSEI
/Mm8dF2YIfYmVP80bEnYNAtTzd8hQmWZgYC01rP06rOHxMPy7t1fzO16ZfNV34h6Y1G0kk3JPmSW
YeykzzUkOYv/IuStVbbIbqfPZexIDfLerM/euJc68d+iSzxg3lZ61O4pQvTljkFHTS1WGKLEP3oy
7c38jhAfabH1aNsDIBK+94Of6RKaB3DtyxAJCKCk2Nb/qO/utr741wI0mZROrqtzj4/F0aHWYgF4
c3oMJUZkRK+n+Ftg0sZ9iylN3wC5q2GAJ8A7z8f9J4N2Qg4RUGReLvllZ+pdukU+B0Nv44Rgaz2t
AiV7lh1s1MOJ0b88zqeR4qnpYh512XFKfRRqSYVYExHDMD+ds/3QNoEtZaqaXfOt2G/lZMvplgip
rbkSyvg60z0DXtrt6JrK2Rr9L2LK0Q3ubzeHOpxi/E8guVLQ5d4X6UfLEAn+rfd7SllsnQkZiluM
1XC6AX7r512m4jo3+Nri0iWlEpJfHpbHyQ35/3GbzsWZnOkAsstbdoSUr5S2JKvaYQ2b8PbUZuUJ
t+gj40p4mtY//WXYJS0AsR1iD0cUViHmdyyJmrhHbuewNlUMrCWFEMUCd/cBfH27HV6F4PcNorOo
vk7qwSPTnIJ+KDjO4Li76AqRyRhBP9PnvutOeF64ZPxINy0CAVIS+uGKZTcv+SoS/5+RYdibTHBQ
bP6Nw6qW47O9SzTYNKxBfViHhTdf3WRHi4Q+uAfc+FGxZGPnsP1rrihsyTHgNAZvdjlzr+pbZRNI
YzT0km8ASLeoUbN6jS0SHWEeh05hKmDzkXMdyMkIHiXfCH1xKPLEfz1ZF3VhTClqEabjRGRvA6/e
fnL8uTu6psF3Nf7CW75ugUkQlr6IwFhR3Le1ib7Q0fwwHQdBNjY1zd8RzQZQB+lH1sxj8Ohm34Wt
kxcrGhnK/UyWsz4dUDmymePvBN8CFhMNM5fGsLHPh4DzIvZlOxLjZC4VpFCVQpitD0ZpKWeOk3/C
UoKKRkrK8gpEXF0pw12CuqNzHxWxivLnDUsVqG2C6ebwsTHudeGRG4Dg0dE891nKq7hmrYjJn53J
Nlcp97gVQ7GxiUqLmAoul1Qt0OrhRX7DXNeEy6M1zjGCH/Vr2JKuMiCuXI5c31n4YIIcUnDxJGLJ
pLibqKBwzvwHVyjz+R6GLHJ0oPXGi4GJUfVSqMzLcgysYOztixRt5N3LNjWe4LPG1p0wt/439aly
29Wy3sDAwt+/fm7QuS3PVKU4OQ3aKd1cplwq7gB7psAU97dIurAXQfGZrpmNM0Q3MzY8Pqg4Ub62
oKuTGD/DqPrUsrkd5G525ikzokD1V7zS33xn4SpbpPm4qg9gjofKFxaZN+SZDyuG685w4OXJwKpT
rbBIoth8flNgNcvWt3PhV2vv9XpZ8rUEU9Gh4wzn5L2hQEfMDvQfNr3xc1NvVG4zJHiZC1q0l2/F
8JlRahFOsOrv97v1b89GFLtFleokLD80vqYD3q+WMFE4jKZU4azDebd0/rvRTiF+1kM6vqxQKkbf
Kg7TUYZKt72NWNeBWc5FROQpgHlWdJqgAZMkLBoulm+S6jcQqvrls4i/7xY6aCevupLd7W4tD3AU
qqh9atEheDgPJYQOo1cKvmU1SK3Hsd0kddNcnO+dOXsKXBmDJ1nptK1B+ftd48YiRE5Qjoou5NzN
p6pJNPCT8s2LDJuT7ezEBSDCF3yUFnqgdKl1fmzBf32b0FkcM+Zq7PJEOVTuUchatknEvvN0Cllm
U1I4LAhflaPjKnNKr5kyIAvXF1DkRPkYiX8gBFRKmUbNlmWh7tfp21iZvLq4EH9mraehywacW75Q
UZelE66s8hBjrPAoYeUZywBNkCYzCLzkVq8r+BYGNS5ltcNh9PSevILUckwtAS+EwrDi5qaiRnLE
7crgv4fjlIphSuDDhFxlRbBA2Lc6fWlZ5ew2URRw/JlfvRIbaNbwXg/HWjTwinqVrodI3sugAVSu
AbtFTEPNP1IV6c3M7MTCYHTXTrKJfWfGdk/KQeWZyVMtoj9gfzDqW3lbf6sfMKdl7QBSBHTJv5k8
7M9Cel8V+lHddc77iLCi0Mx2EzA9KaU8ClRYrntuFhm0YiLv2YfNrIhc1UTTaHjsntQ3EuCh3k82
1ebKMTu35qgnfwRcgmvUTdzukjF38YMBqjhDCtWWn75AOxNoGt3NGPnWWhL1gQzPR5lKHB0gRIDJ
pz0QFfFXxJgQ+jxsq7F/1fqDi8TdE6pjyXM9juxySr4lIf74/1x41n0ZXOVLRI2BouYnAfNAEtPA
hH2Zq/k3yL6LeYwJXPjNYnwQJ1KgrMs6ri7asnYuBQuv4V2GL83kLal9IpTKS3TtLWMdi+xDWZJA
WYcq46ypgwyafHxlBJ6olzyaufkfZ4euQ0B+Wpmwvza4cuZEAFZoVt/yXJZyrM+n73i6gQ7qEUlB
1TilkysnYOxvYdMC0xRhFKkHmrrJ9hLx6ByJdBOjfgef/to/YvPl2Qz1UB4ZLP2yD3YLIVpYyoch
DuTCUnaqqmv8Ys+m6WgpXhrdGC81GhlJOg4cuKgDFGB7bFbjRfXTBG1pGjUmhuBRyD2ONHcqjBgU
sIYHtrl5Myscv+PdC/wqWoGOkyDVwxkT72NJX4TrfjOt/ikGCuxchdxyZAFvOOPffn5SxDat9GfI
x8/GxtV7nP3UmWnPo7pvv9YGpC2sa60PyaN2Jbbs0uJULW7CvxzubwkMb/5wOV/iwFIw8qMbQVj9
3TLUHrAxM8H3pH6WIMeq2au7tkj8iBQ5nrLqvqyEceNu+jHgDycOqV56a7yXliH+0xrcNtSVL9TR
Bi93nRkmHvRaScafF+YsfUU1be+lxRGZynCM5zF0u1iHN2I2QkQ+5w5bMmmheb2HsybFCBIDVFw8
382qKaNePVNTnxwwK3qSZQfm74Hp04t6+EUOTs5M6BBnn0762EXuBvqk7IYynPTCHFsBuvPKA4Lc
QEyKyY60n9FqH09lfwR3xRauuxaOOPuP9oUB07PUTvSZ+siUQD1B+TGumEDKza+1k6MZm9QbifXc
IVyczaALCWdQKk7bwN0tO+DYGWRc+GuoFAhTSMK+XWtt0gYzfsfND8/F5++JJrDouLlDLDA5fw/d
QU99jmTjLeEEBUM3PjkjTyULlYFiAb4IhTocAV01Qspc0pSvpwr/ADfTu5RqCrn8MBXmMCkuUwVg
xKls3pq3JEcbOyukLIDsBphqpqSPTw4m+fzba6rc4CeJA+/e2XVnTa8vYbgy7vFOCoeo9JtU3roi
178m8awEF4fEC/85Y3RYPQ6Ngbklhwm3IZjVU9voYFgzQz3Y+UWPqTqHbU2z7Ld1k0X9c/19rCIw
DLYdZWmALVQyqWKVtKOG/CBkpZLykd7Njvwmf06y6ftR9cZEizc3ECN0jepXklnhemBERiIVf62Q
ghTXmUfULvFX2BUAN7ixyf6zZmvnGujqS0mgIjoJzjJ6BvQHN0rOFGX1QgXTdM8+7H9+yRqcKGlj
d7H2Y92hoKLtLJDX6W/prelLfWD1XS+P08/dGhW93Egs7FHXyIHhlWnF7l8TYi/6n0h9PrD+1CtB
dV/dzjLlBNzBfp3Vqe/BDO10vsd72tALpP0x5QNqWN2hLk46SkPC6ioAB80MPX7nm6f0ACi6TcFa
+2odZgfMLEODq0b2QnpIA4wwfUTve4pkPpweioQ9yxGzc9FwwuHvsLWf78FEBLZ4x78Txl3k8Khz
oK82MHxLwAL5zFvRaqwu1y6ek9EXQg5DMJFXszD39Dy+em9kj6E7SJP1e7HPFdVdgfZqpL1mVnyG
Sy+AeUuwHzrr1Qw/Cx0wGiAgmqrDHAVeND1+vg+WZqBvU3P+yyhUnZYoaU+2LaBYhNDWmxtn7wKu
GrgzR7xG6TRde70lLUH5BU1ydWTwTeBJTbWkInHrTUnEFsndKNJgvWz1QU9XCK6HM3hcmO9eRqpq
N7AvLtt8a4PnHl+N9j/e8U05HFeFuiXhnrScBQu/+avr8XOoJCA6F4fKoTNxcKuZ5ArcTZGnbPyV
eWBVJZr7FM7wa4CLN8+182LXrKsMZp8HqTZa44yyw69YOJt9LyG2yx2cJJewd8t2Co4LlZYhAjzf
g5MbxKX1NyIm+IwxCWH/hHhw1evSPKrzW2FX0J7SNpHV1E1dSPEF4xU9JT9maF7TpH1WVSDzVQng
a/2a/z6RgjPAoX1iGOyO6g7jvPwKdNH0ovX6foX2JBD4qmyjhwptyvS3aGHzhvym4lwoJgem4Qdg
3/sqyBrgy1D9/+I/HU/h3xDLuVVnpTUVPL6Ff7G/Tx5pGUm+zwurnXInP0ttVN+zvAGKZ6+X4MqT
P7nx/47Huy00d76+12leVvtc8lbXyqAGN09CeUqNwubWjIqIGLU8dvvJl9xZrTu+BRAOd42ROiYm
0MfKgmQpvGVeel8mw02Xcb4ST8JVFXaG9TnebZoL9RaXnnYGv2zWgf+8q74k0WutIPEhO/JYyOEb
CX4n6MWKu54bd97a4cQm8e517sbwWF9eh7IjIdylaUiEKgB3q0szee/jgGTEbS5zZIuJn+uZKeUm
gLFq7VXXQS5ekhbXLJSu5t98YX/qHjHZwCovkRlS4ScQX+Rcf7BWvG0IFK9Wti1wVwbwj6XvTLdq
91/ufZvtMYxmAdGzQfgY3PUOvTDp0PKql7lLcK7qQPo7Oj/ftD2qkcbVIP6S63QI+OaRBXbsXvGg
fFUO+Uc17IFQqQyU44I8iTvXeEPQZ4jE8A15E9O2X5r/zGkOyNRg4/P05Ef+Jdv+Ma/SpIXEmTTI
kpeg97pPxpNKTc1giVnS9RHRaKBcgTlPzoFuE9wPFA6giXYWDREY1kNnI9VH4j5OG7Sqq9Y1Uqzl
xQ9OwXwhoIjtRKgP/oVuNym08bd++n4a6N2WRRLsc9B6Q9mjybpla1KrLYVmNKKIOye+zn47dhO+
y6M9Qr5JyIMBt30mMjYN0KiXifVZTjGvEMY6+d8utxiy9qA/2XtZZx/TJSf5k32deYywDOmF5kxd
+CcB1DBUVRugTPUO+3coqjpp2acByGM6eB1/SkNk338QadK44VreM2Bqof7RIJ62kEuy3IGlFS+L
HGSFUx2xcqb0265UO6BhlfsUb7sf5dB04jUZzaGLpJ3rm1uW1Mhf2W4h5isFcCEhPqN1kPUcjCZc
xQhZrPkXWy0eEzHOwGNHWOrt3KBdWWs6r7Wt1mkmrPNiUeFMOnsbNhp6apZ5hK+odyREegVXwz6r
m4iGgpNa9aHTEldsSodroh3TzjJ8AE+J78uemsit1KgAI2dPpAoH85M8UIpM6xbZ/AKQNDYjSu7q
ojTcQ8q6OaDq3n+k8Bfh7mZxUo2JA5Z4+p7q8Mns/T52R+hVw783Ou987Z6UGb1dfCNcceBjqPix
mFNA1BNA5ZS/JCpdnVd5yZP/mVeWMZ8VbVSc1GIhC/RYlwOl5NffAZw51xv2M9bVD5n6l72rJ+PA
AcJLPivwqOwcsX2KQh8b3UXpTNaWjru70AmUtLr4a0Vt2kkO/hPCM6qybr6L23gFY3VtmhTth9NC
Wwt4gdyXXT2qmbbQrm40ZO5wY8h8C076spVmmBJeN65G3Cx9ZB3elTajjQYwzl6I7X5g6w3xFCmF
Eqj0kPYaGFe2RLm0tVxSk6Fd9PSsZ7keZi+rJXIsIHLLRtoA17aNOIuNnBjcFrfQfrI+OnlZOdDq
HwnB1A2Kur432jkAjTrVKeA+JpY9wud/YadBqG/xWvTrTqNghndoaoenRiq/4ieh3ebl25nAHK9m
mQC3J4+TuacOblCK8Dhdulkr0PGvTQXdAQSSmhepb7WjaOMicpRxDPvt+B2pynZ0rdyyRBabfuFq
mjNhc/efYhWjtlienuJVOxojoU2nVSDIQQ/2nge2sUbkW/+haalAWhkMiQh+RdpgMmphvteFJx6U
f4rMCvV3AkJBRTcdEKQkPMi1LwlJPxZ77NB14TqNKFTZvmqFuNXbqH/lsl9DXJ+kBHGA27w4OKDF
2V7TfLUXeLX5ZupAxAWh/UxRZNF4KTXBSLVvocVWNbyYHconNilldR1EcYJC8H4l0TYhNcy1olnZ
YSvizaiX6HexsWN3n/eNCvYypbqVXttUk4PJ7sBNc2iILOothHgwjtq940VTEYV/Bw5l0YD63QT6
cNUeVNl0qmUCfd14xvpCiS2mJ6DOH/9ZN4/AJKdUljx71m8aHbV+LWAoqr2fMfFfPVmyFS3ztXNj
xoR9ijuHuVWSLB6HQe8lCWY6dNtyiGFXU8cUCIjNzivK2fw6g4/z6qWqkwgHR5Z6ZGARFEyzcwX1
6nz9oXemOCuAG3lVrKH8UipRhi7sXVqAIzACPebsjpgrb49x4gCmR70xBvpXG7Ldi1DT9oBbXHK5
i6uAnZYW44+MsgGnvw8sBZaqQv1y4SWSk+wl/+8awVXWVN97eyAqFjSfR7JwJ/gJO6Ods4pFPRG3
cbG+DWCjpXuIoI7IhJOuDZsq8fZzgXAL6MiqF0P5yfKX7DPrpul4ncrP/HJqIW+EykAZCXLcv2Ee
69k5qPZe9QG+MnUWDIvsj+tp+9FwLDnBzKbAZiz6p2VmXy1WE8Cyct6W71knIzo4vK223yaGZIcl
ReoM99/xkGbf7GDGbXJqlMd6EJ3KJS0Kt3iruAwjtpvScPIL/fwLIk83TRKxSOVw45FQcaFcni4R
GMDvJFvj5cGsn1QQcOggTdxxmR1HKdvltRz4Viy0L6cLdWrNydtJsEdyOHWIYgSiPuT4+Gf56Yxq
zJx2CzYU2R5gZ41fAIgsec2ddPu5uLXSAT/wbMS4hR+3zjovNCa+0r6rub0o0N1THOJQAbu9cx5E
4g9HgSZL0HDLyd0KjaxQph1O70dABz3N2Ph3DCKaHFehjsUwWBUylcGH2y/isNNl3ju4YTd9c7fB
Be7heZgwkuk/Z9Y8wyV4NzMJHlG9e+as1Hg9LiHiKp9o4h0vXyhKk9qGPXoTdT3HC4LJmE1YIDnG
UaOxSqCm2lC8ShdmfIWtaVjd9iEv6Dn//r7bFlQLls/L1EgRhdsDSYo79YPnN+/J0Q1ytiaIaRIE
qBHs1yo/YtLdeCNxi+CM8GruhKRKxdjatG461Tyfy7x2IX6nhs6cD8IW6Jdufu1S6sckQMWRmX3t
dFANhSao+TGvA1dVOhFBOB8y2MBCBRbmh0z6GJMxbm3D1wrTJ3O0PGyNskmrHCR4QHLf9zqwTde5
lAWQNCMlS90osc4C+1vFbB8KnWwErdZMQh2XtxkMF4WGF86dcC1r+QnSn1bp7I64EVe65isM9S+L
GPuqQRv2ypyiaGvJPsp2qhaQhtUtCehVWAhZRoAekzK9JzHBZMRNsIRZOQX9ZUa9YGB85Siclg2L
OHy2FU/Z9Zy4tVBhr9RKbw03dDGwWe/I0wOR5OWGP9vAvHwqCSD97gegPbzRJn7kdf0PbVYDZvD2
p9tsGp0CQG8gMOaep10yNXh2p04+znJ31/FADnMtlNNsWPimdHbzZ5CtEptY+liM0ZtZp5Y9iQFT
MVFR44mywp+v54U8lmd/TwplYxs6N1Dz9Dla/eGtx4JfAfJPjVyicPcTHSn+b5yopV5MPFdnZyOv
LViurTyslsxNUOnYtX8GQsjoIc42jOfJBqYMhSfJJ3KC8188EzL1CPJjWBLuLlj9+SvekKm0XYwJ
zlSh70QhEIOz1aLDqCf/A5vdtA1uCLkGdtt8zKkPZQKFmDhjfqJfL3u5k8tlbCNJome1JSUpZhy0
kVOYRfCw1pA9+eI5eVPbHwYnUboxr/e7w7K8Es5jf6GPLeyh6f0ITq8/K73s+IdrntM8ewnVAFg0
gEUw6NLdrO4v9XOMdqt1lSApDZm20V62EBVLKnRErwdP1leVxquchQiE5vO6FT3mdO5pNAAJbu2P
HJsGTKSodCIwcMyXnAkXps4gLunzRvl5QRRsHa13n4YOGzrrkVyWQF/G4lo7EiVWOmO90o8OOxat
/f6yoPZDtT4rEI+zXIS+Kr7I4rSTutMzv7CQisDZi8zs1CFJKy5Yv5JBA5MmsfCKT3ynRSxwTCNT
eDpPCq7oB1uQneE1ajlL/3LMl8rLX3R3uXJWvdbfRlfgUrW4+Rj3MTKaUYtNbtftbtHOK4QKHIeJ
uE6XrlqqWKvIIM/I0qAb/6z7nWHq0NRNEcs6xa22dZ6bfgwKSE9VY44wp7ovJ4vBDuCmU+v4lMMn
akChflXIWj9xM6zOAhptvY+O2GChKdpPbBuGxS0VrVQbNqYVWz/Xia38uNHOjET3O9PwyOlhkQk3
FjMcRe4ZJP/Qut+fBdI9GUVf1neV5BjWgc8Z2vJStN/RbAbQWR3DIn2BPhEcft5zUXG/S9yT4q5g
sX8afAE4Lovjy/+46OkBf/G5q6PRXwSMAfVOXpZaP5x3T9N1LMsjZMdDbY1MAaEneRefi7RAavA7
l2barNC0f6ded8OAXJbGFTNZ+m1km3ODv2RUiM8N8xjZDJJMVLif7D3YV7YArjCvNzMJJBctRyh6
vfdIWkMYQuhKlpwrdRnaU9qJQpnQvy2HiCokJ7JwntEOpkni03Pj+/ldOY6Z35AxlR5TvcAZtPGS
zMORe0om57pK+oFu5Tl6aW0weoqpb2HxW+dkmiVDXGdqOirshZ2yfS6NxjhhZv8RBypClGeaEFcS
FicbtO2rw6Cx+WTe7qns39k/XzmazLtWRWAg9W0kDM87QpY0srcsXNCZLjvX9b7TQWEFgmWDuuCX
oOTEWNiN1emTDm3WMHlAOoRyiz1DEnpWQebsb6q4iR/fY164o3ivccEM1PipptNB950JHoW8St8a
zO5f0pQZyJGsO+UkzDXy9vmXRKiPVTuoWlFBDaNKcTRUdF8rV1qUDzKXCFnEPEhtor5ys+wKtrbw
bAg2xoXHcUCpIWIKiPEw2CwfWPAJMpfoKDY3Gv85K/OeniWW71URveYXUck/txjCyFnbqv7UVxGf
4iJ2y44CgiMxQCaupcA9TeOtzvlEtp97SolSWRcQF7wJsG2fkz9O77nZ5fSGpR56LwR8DddVI+uP
CKgUfJUow+pZnrw1GPQQE3ifIvmsCcaH7TzESy3lwGvJdPsM+kCqSfzP6ggeG+0YqyY1FQnWwBzm
AhVISlSJwF+cpAdzeGGCxpuG5yPu1a4AFCigSUBMjB7z37as3uXwM1CjdDvDfOXyzehfEfhVXrYh
TqqFViZVs3/qhryro4O683w3geiqhgP1KJphExA1hYunRHC3obpuzgplzyCA2as+pNMlMMf+b2r0
rAhdYlGiedarK32pB+E1XlHGEscwsHa44FeEc5Hzno1uUQiDeRMv5ehYLqM+ZqEXL0+p+gKY2gtx
pqWy5Ro3sXs3tfnE1sGKP6d0St+ZjD3nrx6FALZ1toh+pfJ3S8ybCjPleIWrf+BdWQ4XzgYHKznB
8YG3PHKXB8K/x1u7QoskXiX/WbSB4QrkdaswmY1dr6R3Uya6Clb/0blJxAa2cuY4Fah15j4OIxXI
96/B8MbBmgUmI83a9R6REZeFbCpcfPqVpEwg/04bsfs2MNjOmSVeYvg9mJOPNLKBQ15rdebPXZtK
7z8RI07K1STaJNfKrIxnLPrdsR2+Kjy0R1vA/3nmk+tpc894vvMCa1djd+iWEaF3L1fGmChLxV4y
MvKB4dY3zozNpDHHXd1UOD05ZH1PaniijyDz77O09UQwIMuikxEP+NEpKx5dyBhZZ7qOyqtu48Ou
07hqYZDI28qmOZOmN8yIyri9fvh1ziW8PfMTf4Qxp8dDcS/63mX6FuZTMmxFQcnujgjoJuI8Qn1k
+nTQtzSeeppy2ZoXXD4XTAZ//XsgXpswfKLz86ogrDvP7LivZh/rfmOULoFpYr7ZXNkEtDg1H/RS
p1o/zKf1YnhTN3tijkydOa+JpJeFrIQtEoml9fU9gy+pkJ+S2lcPIpcgw/aFJNSjkukoCe/HnSW0
nHNXjMNrL+KR2y+ihwB4dbHd/tu4mVqrPPRT30D3Skd1FMBupFlS92L9QEdSgc9f/WR5zseqgdyB
aNS9rHyEdJa8hRRTubUPXdmHdfp6f66MpYYZ/DF7oeysXVwgRqJoj/HR7lJzHikM8tSHMm1R6BYS
BFNFVbT4EFhjuHfdniDzay/cdoJcmSDov3de5csoros4PeHb1jhTLGCO6Ht9RwOL/MMg09dg2xDZ
/8SJwiX7jiVqS2u4t6ntpBGGJuniLsFxqtYyNGJSolYrZFlyu3U1gku1hdPdfF0kcK4uZu4P+xSQ
MNeW9e3UJNz4uhP1XEoys+uwEDiE3GY3x1GGtvy/DWhiq2ZJEy5fkLYXJgetpaCus6MheRFOW9VW
QWzE/uPXOpAW8gF/jPSsjPA8B6rt5HmiQez2LPRRLMmS5BkDtWSVC797Zjc8lkWkqxU4G/D+Z0so
S6hkFVUmuKjQCOtunXtUPLdAdf+gl1gEmGdp65sE5K4hRLftrv02LghKgsNCQ09SvkxnkbmHsg75
D9utIAuAHAOV3GUi+OYV2lk1rzaFTX4pXF+r0p+3uId8Dt0RbMrk5GjmdUyv7mbA2L+PixWWmELa
XRQOiAtHUzTsSmMrVoY0Ve4481IstQlJuhNUC7g89r3DHE/Qf5PKX/1SzH1emTZ3vuyIJ0U/OLf2
O6tyjFqQFujM0v58hv/JsyPQRGdAu6fnYAE3s1zVsjIfxAfzx5UUzEEDunAphp78l9tTaIi5GVT4
Q9P6yQ5A82hNqcKjnScb6vvByDF5tpzzssxvyb6gOCem05ZukRgSFpNtMNap9QiP6Q9AC3IQvo99
l3QfzAPq+1dXi78Loh6pTMihefkgQWJy7DEKYU/+iec5NAN+XVaG0KAk4nIipEG46guo41MwERph
vd12wogaFqiTlGwrbCGIMYuD42zzHRIBAqS7FEKkplnValcF0LsIH8XM+0PSz2irbyEMDpHDyhyR
0gwQ2d+cMSaS3pYK4Vu42Be6kkehz3t7rKBde5IcrqwRt1mgP80Awv3KURNjXyrHtOft4B6DyaNm
o98V/NWx//w18tlpmh0sGUbDJSazxRYAkT1J4z4eah98q+WpqsK5xlTiDy14MNR4vIfJsNqGeJBO
/sR0Muvy1H5NADjDjNcgb9FRx5qpYaK4R1YEjjLhFR8MiKaRnBAr/+1Vf2dg5Ckn8BY++8qVpTHs
oIRaXWAbPaPH25MT/sMx1LSJr5CDITwYyN1cO0R6Nfva+bi2Z8hOi2CEokL6lkfVZYtljB75eq+v
mUGRhldKUzse0lI7km2LzY1G5+ffbmSj2EMVD/dSSpVNT8CbVJatkXAn5wKeT+xrC+pjWA1E4muy
LDudKoGTCalKQoHgnrSJ1riSYkEUCKjsOWkkmBI7uzc0qB860rmQDWQEMlc5WsWYVdBHlXXi9IXe
iv5uOusF/P0SptET7aFclvXbfbHTq/TkHG65suyyH1G2wArKvStDuZXmkeDJ1g9eEpdmiCXxSkF3
WwHtLwyzfp3OeYgzLmYStH7Ac1Mu2FNaSMqcDYvjpujAF0XKWZUOvHGE0b1QXo5mNaJb7G+4Jdm/
u9X5fE5Y4bu/IzorVDe1VXrFvMeC7zhbUACfWdqgCSiT1Neews/t76TErIgBlucLKZz8PpgxpFZF
Czh/CoZ/uZ/O9yO8MqDz/tyoH1hL0CyxHq9UgByQLWano7UHZyaVnC9YrMWF7OiKy0ZHTOAIXQ0r
fvSKSiyLafrrfy+E7alk89enBLlm0Nlk1vMGxXnl6U6FpxGCFKQowGMQ19w7N1hgseAnmo6Ql3PY
vEmfs/p/We32X8BRM0IIJKjkztxUfmN7SbS7YK6g7DwkGY4QDo1injIvoMUUXr/jQQfl/tFbXhZp
ziMDBJK9ZR9EkGBk+qdCU7gPdjYvH3g7nqMFfYuSaDaOJkdAidUEGW1KuUYvQYfUDnjUW0rUrGwQ
s+iI7o/bil+yZ+0DHM39kAPY0axB/XNWw6mFz8EqBvEZVLKCX3We+/FIvWt4vFApVRsEUQzPpJQ3
UWCiuT3qcGhy+5ypNjEDjg3vwk7maMjiVgAOu8zkxkB7e79rDlSPoe0egXwzJqROKNGVouQx6tYM
55mSO0mxEfh4/uWb4Pfo3qlucBFiad0PACMDC2v2ZWlqVcBPLNaw3wrwlMy0qVL3uWoh4YFzhnWL
/i78S513lSK0hhXvg/JmWt+0+Ur15qFMdxFPjwLVp/B0Np4SmryzpgutAY0E3/ldUe4wJRHjSb8Y
zsjLyfGrDEA4uLjKviJX93c/6IAuTbjJ57iBQkjU1Aq8rixentpn5hA+6h64ueffAZXi8iLZ8gnk
nm6nFwobfR99yOCE8rP7SGRR9odfM1zTsI1UyzSLXQFC+2l4QSzzQquC+BeW92MYfK9WMt76ZQbZ
hQEpNKuy7sZqyuPhTLKk+NyVObRbS0zmdp5BXoKoeN2+WsJ+dM4VB//RBpUoDnphfJT6Uw5vFjAz
kEpftsxLn2C13ZRSFgGeclD6ww1NRjWH6RTsNbJ3jTWocB/7RNPtpzjGz6l2uRZtb2fN6VssZ26M
twa6Z5tn5nUsDXDDS7Gj5Dozl8rri4bpmWXMO2fvjFOqCStJOmk1hryKfeSoc3mxw9MrH0N/Ysq7
pUTuj0cn7daHV8qWdaR1kpyVLuw92FDYyKtvlqmNjNTYoZk3/f4OWHLpjqgwaKe37MR4CNVx6foI
YoRe8QXA7NrFoFdWLs7TBxzNf4yrvqB8ajaE4N3/D1RLLOdZ3i5WOTiAGDI7VT6J9xxrgJWQgaHe
G5WZeIfxeUKfOLfnGNjIK5ATNEaNPL1ACWVCEZ3MfoF19FCGcshPoFeeE5qisG7gtLpzdcTv9+Uf
fvklr1v/JRPqBj+M2N7NY5D4M7M+T3/lidZCtcBmOYc3e2J1CDKIQQLZG9HcrNCN3yFN9YOJQNqM
PVAVI3fwqx1hKQ8rs5ue4clww6nPgQIGMloCBnnyvM+7bl5lmxq+RarbhrwwIhhLXMI5GAYWJJYb
ZOEgha6qqjhS5cxzqGEzVqqD/nzG88zjz4UkOL8nc/UsvUO6IPLWzaMXGqZmmubNIxSr5k/Ued+W
3ccfNPeu8FY49fGCc3LPP0TFnn0HpMtrrp9XmXd6kcFOVJSE5R7yqkj0XfHANexgfJgLzrJOSr8F
MxE24bOLftLlUrvAenLwHr3+27XYOnyyqZpOT1Ig+xkykwuCN1jXfN6y3aQjgUhF3onHF8qKxwwB
PRSWmwzjyAqY9vFnIw4Q7YVOuiFxRM5K44xrEQ0KgnI6CuN9JfLtgK/AVk5EjcS5LF9K2qMNy7LJ
orGLwnZoTWg4rSeHVACEtiHwCXgLSVpZhnbfH+kDCaMcRUUtFjcOEc/oHKzdxkq261iLiwMpwTuy
9m+X4K0EoOESIOfpZQaqobVcDT1/4KjfpaAXDZdOEsLnCWqEsuQaobAuMR8HGbB/jGbdTLerJuUL
VW2CYgLKLc7lQZCKv+F2IzvlaC+P7cwdkDEgivEZc3zNICWnaPTWYMzHsSXFFHQ9afk/Vyr/HOlF
L6//DuPMpo/qDaO6Id8J4fMTC1+42hh46Q7poHRx8MfpFyx7OVzFixp6t8iRzxG1ZlkPFhhEQs/j
p4VgUnVfyC8wMsvLbaqVEYcyinJLvKyUKXy0giQgKP+RSPBZrfYsHojKGxpAcHdOUYM3WhV32zhp
Ziqmzc2ADFpaKKUYJdHCMTYV3wRi2ngsKYUSniRGbDGLbsid1J7p2UZJ0NFYC0wORl4eN5OXaBiD
HJwi6yThEVygvZdZagt9dPktSGc5oyYakBhWmPt3p83v2DbzHoV7LKCd0hxHIvnJLheNCL2IDRi0
/xhpXznIAuMSzxGq0K9hz6BE9b3f7mtKI9xcpxHAiHntKMAqaXWgLGl9eND5/PBwjqjpxcGregPK
H1paifaIIm3THC9MMWSdnluaiy2U/ChNSlewVcNV1OgIto33/LJljp2l9ETUnvRvXXVl394Vtb7b
EUlHRm7HmuVP/h66IFlV3wvS4IdTMr30dY/LkOrNH3MBXtM5n3YikYyW/Kw8Hc/hvb3vWMKDX5UT
TdImZnv+KwadbTmgB7qOTmo51gfnSwDdKzHWhRofMuVZ7Jm/Dawcpx/5QWQSshiov6JmAdmJCPFf
TC5UXJNAIHzIKJ/r/dc2g2kCi6CyZzb4beWk9e061vRu15Eo/H/IAWymzYENhzRXu37/NkHA8wcl
brz1bgC+AoBgAQ+dRZUWaJb3OQQEvh3oM//9JeY7c1gmkxzOpQ7j86/U3MY8qjRUYNZG1QrscAe6
gXfkh7X6kAbDijYM7Df1JLMz3qZ1lsF/++evdtGNKcSEcfrFl27ybDTcuj2imRMJHcute96dsedO
245YzMtBhEOsvXFchyPEHYcgJAuWJhKwNS4v97meKm3sES8pLVNRGN8E1u6WteG+Gcgocc+2H5Eo
hu+yaZ+gUuwHIktQ/aozVXuTyEj04SHJyBNeebvo0iUs0rGmiTo0lAbugxsEkLTYe6FcfTk+yAO7
rJsbq0B2erjjcXCLVZWrMmhikDwXwJDPxBm+4BvI32a7O5+R72qk2UIXBp9m012n+uFZVfACBSpe
WaRZqbMupY4Ezp65UIjCSlCuLxJO3rNX2Qbu8BnIPJWzbbKIp+BqrlSfjNbdPNu/v4pyAlhE2Rk/
LLSKE1+2Jy1C8ANWoGSxCRBf4P34pKUDkJlXGzLkGjbyDJaC39ZfIzWZ7Pzr6GqmjT4vbOLmlETY
PLMmZ67iIgWtbWWxcihGDlmdJXa/I7KjB7/ivkNgFt+Ts/uepHieUDUyN1sCHx1ihdMd9ifqfwui
E//+TVzk/RyduhSrvTeI40yH/8H5kcbM6cJhjKo+j6chgmKjOrpagp7e46CVTS6W3WNTpA4YKpky
F5ACyDFQ74YpBUkwasRxZCDhdQ0hEPXQaoS0V+RdfGF0cRI7KRtN30UesZKw04fvMyceuTpbqILJ
xmdjhg5yIdOv0krabI7Va+N53ZXFrCEeNaNOujTd5nQAwEf6dzkpY+Y1/nAv0p6ebkD1owcShZzj
YcmPiDeZXzFcWMYs6FnLNwoSTn+ToLUuPqj5okVBIviI6N/+CTsctFh8lVQCk7MTqpttEw9lsyIj
x3Wu76qh+VfJlZr0/MHoyhmY++D48lECxvlNdh5/mnvJSX/nplk0FUY3vOCxu2m2LKSjw6EnYly6
huzv3KHB0vU/WvNUIbitHQ+UQRFYiqdle9xrAoj5PLsoyvm28uKQg7/Omp+qskDqB55kljmNIFMJ
VSH5fF+gz8MCsMBUlsN/NqpQQe0xMqyPg/0KwDDBFkN6YBgOEJhx6BB+3cXNWdWZoRCqcgqcHYwY
GrbL/G7ewY6PY2pXFfVptEcnIyb5dx+y5QLEefwXtITP171RYqfCtw2q27VHPQSUQrG1UsCcgwe5
C6MIPN2Z2chcuujpQsIn7M5XATaGuuNcy9Y+0RUAFX7VYiFWQjQWhBQTBAlaDBbigNljgTwqSXZX
N6qIRH5vHzPoeG43gooDJ6IElREQgMKe7tun24UqZ/EA6PvmPM2jg8D7Qx4fxrbNPH5nNgFAGDj/
sELe2mjtXPlK7X4MsrY0d5rVSNHLZfEev47oLezt4mEubDMMxXc8KZ15DJNPrZG/e0SMYL+vAUcT
AFZ5YOAJ1CaFEbJ93T/rceAsDqrVv0OjrvhQn13Qmmco6J1pg1BhKjXlGo5Nk+77HUhOndKzeEHS
vT/qn6XH38mALk0hXrUnYw1hdSDtCwA8hW5YLzRC35QK4m4s5CZKUfgIW4ckZ3feGlG0FZa6GtkM
CSgsPgeUHCRvP5t9TCDfBi2JztWU2vdyhdx4PP4S6WPmOzpHFR5pNFmv75um/+7VNqccXWwCncfu
ubREqCBkxIoN0aAR5sToIGztLfBEJbO9FFauPI7XUFA1rzb/OH441vi66yFtbSw0LOheEcnaT9E2
OH5ECCSHXzuisOk3JMKcYcR04WmgNGh+hZXqW0zak7jMP+qiLLnE+sZsBHC2TyZ12kM11nE8uG1V
z/L4szKb7YFteo3Sdjy16/EAtIHLV8myFK4HsNsoacDzfJ8cdaQUMoQQUtVOXR8U1cnouPcfaDLI
kedMrlHImZci0qJEp8jjxOqIwUcHWAfXOPJEA4QIiNsv2CE9osobHWBYUEUr46iJ+jgEmFviEMCl
bCKeNq+Tjzjh39QiL4kUA70BZLbhby0XqxfepS14O6ewKU2WPtXvkswOkO1xObhoLqDrO72cunw1
U0plUoNclH3/NVBsVtsv9WD9sQu2Mq4exx+uBNuqxBDB4KWedGYjucXy/0tw2Wdbdd6g4dar189F
PniEhCG+mQ5CCulRX/tTkQm2dsiMO/XuSxZObNawdzi0jwl7UUG5daFeIk/Lh05QBQdoRM8xxMGc
R37LUajGov5SO0L6A1xltEGzHP8dykATBFZm/gXvVidKJ3eTz0uhpMiI5B82md2UH3ilIdZO35lC
iWXG8WKV7bzWtnxGclTDkV045dmsxqxryMQXDpS1POS3aqPHwJbZpq2PWM0Axxd9Gy2aHCzs2Kpg
Fh1+fJaSZ7fRMbkjg6bHckX9wsPgnWOQjUPFWTyz4NBdv+qjck1YKXG6TCvSy+cfERLlBhZPpldL
4Yvrx7IIBTxHSBZBaD0WmuFyMORP2+2rSqltikjaPJd5a0jkyMeb9rrJpdSjyaow/N/cB+Q52ZRf
0OYtSEi1hkDe8TWMHLe8SJRCbnwIT8B8LawMLtbppmsMEQxEBVIRq/hZ0KxKkkP3Z0wykETp10YG
BNLJDZ5PoBr7l54N5WZ3igznpGLXghiVA1wdWa4C6yvqMLccYJmpsWai3bk4VW8+qEu3OackuPp9
3grnOGGNAjEpcmDVnmYoKUOS5C+RiM5MnrIXsCndNY6feXBogc3NPaSL3CW66B7ym1jI9l1tmvuy
Zll7SgZC3uDFuKwtGIDNW/mw0vCRlfrq53tpodEQ1UOUL/vlPzAgFoEuPm49KN8+F6Q1ebL+ixvC
vMusZL2k0WWx0Qj3TXheDTnH/cCnoHCpAKfTWUQgrHChGIc47LB5JmL9BSF/IC5v4B+eVGA0epsc
vhQ7Ar7armNRQBNOqJQeDPuBDk7VuFYgmJ4pvC2Zc2bcDJZ7OLzl9N37FSiL1WdAJ5hJg23qDaHz
LsqnlV1/tiLTxFsyeTaCXiL03ENnq2J2uVGLi8UdqFSdunbksTx3rthUpz5M2celNo6pTEW/TIgM
zaBooF5rhs72vXNCfSwZcnEntzwMiszgPkLIhbTyzlOVdaqd0PbyQ+S2DzznXPAZvLx9STvF863I
FxZ5DUfgg873TPzfei42Dkf1iSIOshWTS+hO5PytqD9jfKFO8ER0aLiKDuECH3vBXh7NVcP7YEkq
R6DHjefXDtar7R54KbBFmfIBYH+0P4yJ1K9T6tjNB8VdJuGdcXIfNz3CCI1QhRQKu6RxTLkYTr4g
NG6b0XO7Ktz6u1GmDbArr+x0uSePKHe1jV7ttODGwmfK4HrZB8s58L2zYELMejePw3tdJvgqEi0l
Vii9S5ak23Ly5+8X4H/7L2i6yTtclh66NnM51lsV848Z/wowwhCOUu3tADTqaU8sQWzRpxTIl/tr
lFdfBjKN7oePrzOCbL7a2VfZavqroTmtjl0MHZvooW/Jp2StNh/i1V9vssys+/FM05hQvZN8Ll7S
HxwYiCNMmxVbh70decPAqFnIwB5/dFITGh/j5cGEYPtfIpRCpBHgcRT6vpogc0O/w96GXMJ08N1r
C6OK1vqhOnu3v1nWr/fJPxabNCmXXuADDY3d3JUiSKYI2Db+XvmF1tw4hMQZnzc8d1rlv8CR1vIe
HUL6AMyxCKooBKbv+Sd288Fn9PeZUIgrDTAYmPvehHR1CiodNnlhYSlwYgFPyY3zWrgjy8T+vOwB
8qv0pRDrSTRjOWxOagP0KeLLKvt95+UXG7a2aEBoU6x4/s1d1s5uWxSvaXy/RmEpIof+6vwZTfcp
5h16nsgHi/skWbmf6/tN9tTjSiQw4nGHIM+HFxpXAMXJZqlvly0QBE7B99CGy3xQWxNIx/Irl8nP
RFW1A4UosamU0PaGCwtZ9HZaIAvBdpDsjgAu8W7o7fIRyNfNQvMqa4Vzd4eCVBO6IbzJF+8lpS3w
/Hmvgz2tbtoBKFMGDbl3K5cerAv/QiEKI4Bnq2MYlaETBnT0ElkE2/0dUGHp8omnpYP4G/pwqDm+
LQVeaGebxDYPVw8+SCqbkRVXXBdQdIMs9Sww+1zSQgA4dZUzM7JcnhdCHWy8NvnFbS6+p5a7K3E7
hdh5IofVbrk2EAr+VdPO5zbDXeJspyYBNItcUqYqK8ifCIU5lqMm7W315d4HfuZHASYPNZngF22Q
E0k60rCBssoW/+6F98zatFz15zSf3+J47mGlnvCdJvmeJCPI+XVUBVfT+oH4imIV/dgSB2LeJz1X
sHZkjDwVzz8irMN1hvAZ3zOqwI5VUYAlbk9VtBInYkIYC6XNLBQ4gpNnjNTeMpb+05fnRPC0yjHC
iRz/vh9n1IUK9GvhQt0aiL/4s1Rwjcm7J75szMwEIYdAxyLt9YskOdSE2qWmdAKIsLcbqEcM+f3j
LBi+/bIMcAbspBNsSHfnZGrHD8eaf3TXqWK6wpbVcPR5w7QyN9siLoWTo4NMr9VGa9W25KdaRR79
YMQyUQ1Ah+jHgpW7gLzKJBvKJkF9T0TEWZM3F8dKGGU9gw/MpiXc3iLL8XTxdmq8VbwQxgmaJCZj
iIOx9Vymk9CLxodi9ETgVT/56DJwmXCIPyJckogkjFpCzvFPrZbfmOC5HBc5VG0alLDNhoVnN+sX
3J/hG+3ZgxxJHILAeE7lu/i8tgbWr5brHJsSH22nW1BTWOVij5SX9UGEAxTqa4r2gSXyBJfTcPLr
0lsCknqNEPd5jYUoOXytM6gT535XV3AiLDpHfqZ2rIRhN57fQOYbc7yvoRqlBwKU0aqBX+kiXDiC
XXEKdKuFWKul3LCSIsrX0kEdyuK7wNEBa421OKRieyUGzoPRmd9YyuGQNloQrwuzWGCNqNW/W+Sj
6/QbsG9KEBg9cMYqFBMUOgm1adyXVIP+O+vdn4LztA2HyKzEDgAQysIEfvB0KfY2+xhtW+G0HKJu
dBlgZRz+gW94pVOEZwBIZE4v+xT95XXk5U8ru+BetlpaGXDDoK8x+qfVQdBZxfTyR1oFGHm6PLVE
xAeVnP7PoBuoFUAGRubA6Ae5+iSbKAIp3opz1aOsatW99sTZI/5t9OEWtFjZRC5/XzfVOCCBplLT
dOsbUnpI65a/Y9WIzI/xFYhxPA1OCEQjfJOO4tBGw/Dx5pMTAP9xJskC88QHRSkzwtgiGAPj7Xm9
J9T12ganSXSpHqVT3B7E/fIi9zRueg9Z1qN3wqBMEgUNLvdsEIrHCi8sZhzzVL8jBTSbvHDvDs7I
Z1Q3p0FOnSPVIK9LKl1/6Q1MDx2elFHeuI4Vko7NGmudmvd/H/5p//DVL0rL2Kdq26pJFu5SsJwL
WJtjAyU1w9BHaV4VOeJoVqTqFSqtGcD1BKN1rCE+TDBKQx3JMW7snqCZ8fnFYqRVkNgjCy/6anGq
3kgkc6WyjaOF6XlYMSnvWI788kQo3mCBGlMTcsGl3akdJADiO/ME8M4l/KoiU2KuCQcTtbbYe2px
Nh9lvMbPuokXehpQHn9grHv4nt1bMWAE0WD1d/VxJ0O2wRDoUrChACh7gptlBvggWjj0ELyD9etZ
6izri89tCK0DAbHLqldQsDn9LnsardtnrOOHlh+oKnsN/nvoMR/nOmsT8wzFjxT4yMjwsx2ixEIb
bBeOEkITHsRqhIgPNf0ELcoalvQN1erXDBybQqNgQDwFWcWyQgyRwVySc8jtPjbcpgLbIkjMUP9D
b2HiRkZ+0DjR2f6Wra7Ti1vFWdXq98HVO/ziaPlDhi+tB5LlB4bytbcfxjShXUVuwhIWwZdtPfgN
CrS3qzzlsmIRu9KGZawR60EacESlf0caZcae95iP5/b38NZH7U0mB6uKHt8LlJtIFa58d4gE+ZJ2
7DqsdItaiV/zhiWjYcnLgMef5e2KUyxCEUo9ykAktwVJy4FVmexJqal7/ZB6j9Gbuov2xzu8fXK/
+/LjYKWQFFvf+j/jBt5ijh8cyLe/3Ukv6v8haKWhJdlmNFHVqDNGHLsJJaZeLGe0ueO2Ktw//R4K
aHQfn1YV6Aw8W6dpCk+/nWL6B0GiFndfFq5T2hKeDUcylM7GYc/TU2AbwhycDAsPCuTlkAgNa27i
ZsgGT0zJBzj9qysMGaAQrCXKksFuwCbClNS4c9Fs6tO/yPGg1tEasPx5yamrWelg74OJvlouW0iZ
t1dWZpy+AqQPlC1aMxewIkQLOrI4WirDMWiARmLedTlEalwwrzPKqs9VKlk662GG5xppfcGeJ0on
nGDOORc9ONsUkNrvStLiTINmvrTVgQJj7IHkijiTtRWD+F12pm935FWXVn+e6z4YeK6yN97k9aB3
vRJ9vdYyVMoJ6r8o8XZy4cG7zUVy3W9VUVAfby7yvjGAxILKPZvHt1QDRvpzHytOdQ9fAXU+CK6a
exh/918014aJy7W0LnuYFslhZ6+Gju3PvJ6GBpYcmlEmUqol25PGCSVd33cZ9nv0nrMHWz+jgyjo
hqU+7MPhSlGMe31IAHcl7Kt+WlOZX0BqqTynkG6SZ6GJWoxABHLnh2UepXliaf0BS54KfnvRK0om
P7Ez4fOY6ODel99VEfelWEKbhl45YxridD7BBihZ30j07KxdE6Gg27EvhlXvVHG6kjdkRxvpy4S6
HhiYjwVLG5ZEwrTBM2wNS36EWNg4VAbGcRZCQi/NVCeT7QcravpO7yq1+uXeMK/fD1LspoQXD8zS
uB3vzSt/6EnRmKm9SjDf75C1wuARLjP2d9hIBeu0cPx9Ke7RNctQ5/H91fxGypqH6fNEHnaJJa3M
z5eHefNGTbST7A1op/NTcu25Yt1G4XGYEj3woDNGrNDyojqL4GKThSjhp6Pi7S7hzwfDjzq9CLMC
j28jHFKPjINc1HBauF+gPfoeiBnTqaQrb9C20orZwQ3J9J4C12QL5uClWLXIWbAC6NEDDvF2mcMr
ZCKQk4qNuXPXYQYl7qWWSl4DFQLGCir6COse9TtvFzp+i1iZzzle/HCLPRdng/WGD1vAKN1Jr9Qm
jAnMP7FeBqTewNIEo58rWV1m/CnovYTExRK8gdqv7g9v7HeaBHbxOBPnU+lgmQVlAGaM0HMHbNAG
N06ZbjEbxKYAgKw8P8g8AqwSPC4l+86yfa4pgazIw4r5/cbFyKonPdUK3ANKLiQFav3AyoBL09zB
o3yMlb/BTUyON6Pd9k4RDaMJbJFyxGbujg32HkFYKc5VXzWO5TpQ71U1xsoFr6lMiFsO9kPIGXa+
yhcVVhix+QPzBbCOt2LKxchIfwE9b1XechabbU5SlKBQVOB/vSNMfo6Hat+QUA2gx+1Tu0ZQbfE2
UMedWzen3B8WMqNgeUAN/i1UWZi31J20M++iCssIqM+BeBJR8MHPzeLd0Shcw3LvWGrBJtnMi6yU
EnIwF3sg+6/NK0qvio2ZHPYLgWerq5+jP6FI7O5KOrOv8zqlY0UDgYF0LWg6yU2ZB3xTnWAw70bA
rt7LHtHP2zvCuQZZ1KnsFMFAq1fiEN5JAAGqbBfW137dtRl3sfSE/tKKWa+aB9WS9cdzECz/GLdm
b0+72FEi5wtr/q14iXj8tROm1caeyzaVYwmX5N6l3sVjW9PDeZaCi/oz1+uk0rkuK9OGIWFN12sD
UI60hgPTjfv7LIR5utiy3E/dT8luF+eIXIA7uFr3Cifn73jaWV1yqA2EQDHg9XIMceyDypcINfn1
jIfsRmVFHNSTFZbWfrcPLtz1LbpZHpXL6W9BZCYqBY+Of3q23puy8xRuS+9L5AeSeASBmQvK7mfR
3LgCkMMFUSS25H9TMy5wQDkg8gIG1r1hoaNOGfYYYrWIPulEULDv18zmhfWB8TdfjHmmD6wgQOZm
IvymjvkEFiaZnOQ66qQr0GBQoubT6qQ9gyOvk6el2HxCeT8oDI0ASQhQBFzQMrV6qIi65CTLxM2C
uD7QSpdMr0UTQaoVBnge1T2dmaunT0nEeWT4XThc4AFdXXsCi/MEfNTNUoFv+cF8di0edfP/tVPf
cyp58M2T6Yh9H4Qex147PKTzYxU72P6dppYdR2H6kSqSS8sSnwGwY+Jc/XSYAayYh+W1MNnyf8Ms
vprRYYBQLXgQxrffAt1c3lzwsyxZumbAoaV4RHfsuH1HF08bCoUHTJC38EgzElvlw9e7meU3rnyE
rFXdClz/iRD8StoDc6DdIq7LNMpKC3ygL9JIVOy9V1Q+K7QjTEezEQT+YY4nkc1vEgHLy8FwIAB3
80YOLXE8wJUUcXcaPYgny615nD5XLlcTAHCZscsp0g4zrKmEQLG2qIc0lc6WTeU1iXnEsDtUGfZm
qDsKhmIpdTioOuT9n9PF/4gFRAJMgP15st46cZIJGEeLUjITz305VSpo4hHDoO4KDhiytxAUzrC6
DTXe4fmmXscN5zpvO7NCdiBpXuh3wMxXYJ2QU26rxF96ncJYdU1su/DHay04tVFus7NgRk+yVcqH
EEqvJzatcCiBMQgKy/gAq+Ge45Fq07tRk8C63XtOy6Fof3JIwoGCIKiWTrHPLCTgM/I1TTkXJKot
RguyMI9CSIhF0mCYxVRf5F4xQ9UvBBzuVvHQekBd369zgpVYnS4FZwqBF49bz1A3ZgEWZU8hvpMy
CGZ2b8L0K5rYnMf+E0bpYH0R5g+8C/8eD0e/ymbL0ABIs7ngMD4Ly3qfAxOj3pUUeE8D4BC0hCbv
1cec58hYJBZj0yVOZoJJN4fPjYnmffogsDaxpXw0KBNrNw0cV2PFunpIcjpU930rJIhN/Y3c7WLa
S8My1cFU4VmPWxQBhaliNMxF0anKFYpgcTZqfzkUjq6qmJjDEpGJ1NNPtmWlRUg1HrJ6GIRqaS93
CrfRBuGrRq/tAEz+jbC4fHrtkr6hBB+Hir72FSux2u85qR40fHntKFD08Ara5aEwDT59Hy8NEu+a
KDBLUjQrFr6JtVZ5AroRgHiM/A4/x5Ox+w6eCqAUTbEPUL6h7Kpey2IaQY4zF6Y/63KMYfUFcQtU
F+GjgDb7jk29V9LPet6vTBLvtmPXGhvCQrjZMDIQy+TP485Tc2DLOpJOQEymR3/RnfkWALJY6LA0
qVzLCrrkha1Hp6E0+LSmb7Zhfubh8Mew5pRHm07Lv6ZO3pnrSIjvoz2/rrGnLYRY2Dhg+hMvhrxh
5d/UfY3AGlrqY8AUjvqz0qHtLdl2SW3N4x7mjH2/AZa/h/CoSY6Dk1MAf4Oj9XgX5uE4JNunbRc1
PLzz1TZgqhsRgVQlyuWrrEZzPrMS47LLkkLcEMTS4xdAQgUUz4t2eNNcSNS0JjKkv51io+aADo9t
dDaN4cdrlWWsz6Q/MRy2QyLMKN2kX5agstl1052g8J42oxOliWLAsELr9BOEMG7pRXgTDTWXvJxo
szNaXmWDvf39vqBG1/sXR3BYUN4c0vXVTwoPcypJlP3NfkwijX7ijgq7ypwJLIbNn1o1oNj2cfpq
KG8e2iNfhMezP6WKpfRajfw19sIKKHYgtj4otK+m0u4g4kk3qUDLmMidd9bFh4pWD2JrIUIDaLH3
R4KDRxFbc/zBf07M5rs9Kh16UeJjRw0h33OzCi/DiB+3R+wwael2qGy9BAYpnUi42zgd0nTfVXEu
3+83/6zSvQhIIoL/oZ8uJvD3atsGyvp2Ehpt10n59FnwlOgWBC37L79CQfuIKnTBtlpYBA6M0ika
ShjQL4xYDmfW4zn0gL978uyr371kHGHdZgxlCxvWvfOC72AZ1FM2i51TMPZKK2ppQwoSQztLUD+e
DVPlPe6kQSv1nKyRFOIv+xmPSnLfMvl3mYMDfKBLoHtNK7ezZldcs1VhiS6+0zpLE+ZzF2QvQmK2
Iv8gD/yJZi8GD03TpzjnH0hFodS/DLaYgt2PzaLTlrGEZhXA6BjEBI/I448dhnpr35rq5goAHEj2
M7prloiWXSSTnM832zvm5/cXloAyrHvVaiIX/q/i7EF9bFRABdsDcGZqDCfOwLGjooD38hvqkfXe
JscuTZAU/nLhywY2iYkWNNw8YEXeb6uWyAc+qhOZRyurRuzW9ogcBRYvQTafo2bPpqakVuMLHJ2n
c0YnWYq55OeaAKNzPbUgRB6/EP6L0Zgt3jn1ADKBFIOwgCO3Yo5FEirDpHYJcp1WZSHoPuC9f5/3
AC60kyy8i8ajs80D658fhmqxi4XYiYmFS70WRgAJb/VlpPeKJmtpYnLRERfFmjVJ1dCPHZJwimn4
XD1mbwB3iWzA/3RLgUDUbok9kRzFvs30qT8c0yjTTep1txIq/SgCsxntZ+yz0wviZ/fu2tdUqyEM
SLeAnKGAF5aL01IihQmmBRQlOoWniDyfy9NWuF2CjOKpUkRxIpE6CRBXAs1o1gH+tbBymmx0rmCz
m5wB/Shrqo5khF3X7XiuWGGaPTx2nC4U9UjsVGlE79LKU/d8gYFauul2hGWU4R1JCZyxbHHiX1aL
PMiP+ulwo7RJqNEw6s/wzKa3Cc2geen8RRuzJUsqRa6vLJiwpJLniSAut+aLlccBwWW4mBJmD1MG
dup8CnDv44J9hEKh6ki9Zg+FXV/W97/3pR07w92w2ZD3BNKPBz1VnM0HTF2m6mPVe9yacSLQiZmP
EmBYUpZ+5+wDLbxe5ftvvVmTAbae8eLlFGRyFCKrp5D0aHUchtffzTw1d9uKDpf6M1dWSGz6yCPn
h+FgcYOzHxSt1oWnp7Yo0PM4k8hN/qQ4nXp5U0zOCS/OGUNUOWNc7sBsUhd8RInosHEuIQABTM6/
psHKWldYXH57ScmVofm2e/JHvpOmpIpBmpPCeJEHZ5NzTNJGtf1O2MfHSPVetppXFqdFGWZEcolX
xmI1fXEq53tyc7wIhIqq1XIKISjlwaOe9Vw8zUwGGkxcbHPc6xVp/OMMrPeIUjjqRpcXTkBkbm0X
LHTmyxeqh8EKuKh9fNrb/uQUtFn67doNDxWOAMBeH3BsTwRysl92LyciaLldp8AnMAhLBCTvM+n1
wrODavP7tg5x2Dg9CijzdN3Gp2W4iJ5cDrHF5HbfnfUAnrdE++Rhh1KK5NDlx6eiTmmv961r9scA
0sYjSdIA1d+BRaGBsCEhlHSb+Z62U/3f1WfWf1dDzZ4QY+Qd1d2Atqq9xuJmkzKDO0OcVcp39QTt
gxYws29VSUCAhKIudz+vahfw9XHi50CK2/1cYJEbs6xlsV7wrF1ouk8/LU+o641TIu0syOyi+pz+
vY5pqT7g3ixfJ76X/a7/brKrkwo27eKso7O+SQE7BxVl/JSj6u8MdSC5hIv561xHB04XAgQueoKv
/AqyOt3WXyISw9kUcL+zEdN7/ka6DaGc2C1cd0sTj5QAolEFciXfIbCObNY/CO0fbf6JNTcXpzaC
elSBPOhAmf9Cf0eHuHk779dx4tayyv3ZC7bT1itoUzPsqvnjH8MmH09z755Tc+Cxn0M4VmF3SPCN
F9Uq9BA1edoxT1Wae0p2RXWihXC8S7+IFAfzCJv7MIdR2Er7n5ykqd0MAVFZ1EPyAPX3m0edax6+
iF0NJ1rhsKDkz1nvVIZL/QQTJcuCpSuUHbSiRToOpo6sCVWj3auRI537iKd/BA8ZfTbBm1xoQVkj
UOKoOJ5slii41Gm0myR+zEp2djtFty1QorFVT8myvuWceGxp2ZSkjQsKU9Eii3RA40qR8K5QLX/3
HUSIcasRpVt5arcKGLEpzd9sQNpWYzt7S7iX5LVlGAGkVWgbq4UQmt1zyeBbe5XLUSWASNQ5WWQD
RS0VkQ8V/ugbIdE22xZ+JakJHuCayWyWZSdJwZWJa1Gb4VuFarWBU/YZqHZgaC4DWJsSxqtjTDY4
PXp457VNAXt43MryC+Q4RDOt5gPU2I3e/ToCVTLn64WhdDp4fzuz5lRNI5UAp0+VpGMRjaUl9Qa3
YT+8PY7WLRNj4JILDgroeVL8U1Yjoe35/8/kvBfkrgGy67zoCnX/neX7vG7HMVoIJqQmssychj5m
2PBW2lHqbv/AUPpSt2CqVIV4DSd4UkifKA12gV0bGq5lmNC2d1rX4rHLG15wxEsReRLaAIbN3wza
vyCbwGhQFNO8KpeC16MY2Fynec3IRNZcbqRNqbh480u/eaHTikiCBHTivRyHf7K1Ij+NGcaIFRsj
D8H6vFwBHFR+mxd23D1KuOHdV9MMKhGvUjPav50T6WwUS1MP8n3CNtgKRcPHB6J6se2Fw/3noN3z
nUUqumo8L3fe4F7HbPVyuyExQWmOERgwsgza5Uhw9p1gBFHM8ZzyoqikgqvnAuK7WPrJeVvrPoz4
2Kb8Fula83Coq2HpqF5CLhQ8jYJcNRcY/jc06FC3OVBuzTeUk/d1lEps3VWlxQnhcLAa6FqorKX2
IQ2LoXHhqW90PkaXY3gv3NAGtTubVrBC+w65pNmHaqcGHkmoD8mw1aAeGGZ3LP6n+SktACyQ6Alh
pQ9OFqd8PQ5CTK29hZcjyBqcrbQX9mGcOndkYjSdUn2jTgX0DTyvh2PfoZgm4jnoXtxjpNKVdSPx
4Yq9+f8aK1LUVgE0PclgggXjdmnFwssKErqUUUbfI04Hx0BQnYDMy8O9xv7oOTHcJjBxUmhEmz6u
GW5qO73dqRSU2tp0bYi6pduqod+23i1yaUHwLnVMiN+23n+wCLZwBtkta+62iNBpAQzikpayltQe
RCVezC7QgjJhibiQqXNiIefa7iOxoIJwnltztcWXZE1TwJUabMDpeZj8dJyV/t3nHD5tgoWAGY3y
icvAZu5BAkLI5vP4okANs9NkVGgCxMA9urCedZT/Bq0ohfw6E9YvBdKRBFqS03vKd18geY6ZI7qQ
0qOIc3Be61mSyS59COYgQIZz9rhB688yv8kNCwz+x5CmnTvMDGQIzaBRX1R8e6NGWLtHXMgp0vjx
s/gZwfP0mXqoyghsn2DAd+8auRTuqO8cK01vQWzlYip7zvOVJ1fVdyxomxFQggHjxv/523C0tIIn
utacP4H6yR67okA9F6avITAu6zBv4Ecx/cZlsOVFlOW0my+L8QEOn5lUOWpYeP5scXNPZ6cNa/BX
XhspglRqLQzeJunE4xT/D9RZ5hmzh58lxdug+0QHz7bUS/zAsK2hZw3yzfM51OZtOMtXJuyzVVlz
HWZjK42s57slUXw7dT/TtldKexT6zf9QYlH6xp2PT2KumU5xhhT0TFjopEh+89AHhPGiBnulBQ1F
Ho0ohFZsUYgX7Dz55qD6arKjm8Blvm+nsOo4e9KClwqHrY4kpYIfQCUaTaT2YGhL37HgTAqzYZSo
D/oABkzWmy+5E6Olo8QWnVsuu17k3wZDTjutBHoCVVHUeipzrHnpUdWxKf/1+zAoO6nC8VZ3gBfr
1AWoEQZTpc6ZrZE00u6WMDNshEd4+lnC/5HwsGgEcw7nAVTOfFZq3wH/kWZ4sDM8+RAaA36/SD3n
qgzUV4oBx0fQZ1LbBiI5VZFNDjSzvtvvyW9+Nd/kjFv5ZoJv67EpNFiI9P7AhXjTfILmFgfuWExJ
NhLynVIj0nEfdjpXMqPyjG5msS/Y2wWnlmNujoEFbVGCAi5S51S42frgn0rqhjzk/QuSx2pMmHIn
9i0PiGijMAi4Fs8mtMN7Lq9bBajdoug7z7Max2neNaS37x8lpdmARTZp1WoUMWfCeK6YFMSDMO2r
3YASGQ1zWgBmz0THOo9I+z7sxo5HYozuurD3wMg15IuEChJq77s3djo23ItjqvPGeQiTQEF4nQrc
RtBckrZ/0Plu490Evg739zsGyWJXwADYpVf5z/7JkMd7m5seSvlZCXfu8WXbdTz/S/YoHySEEhTx
2azxtG6qKDlyTfDFJlZqTJyJEFSmPEsGZvt/P+m7AOLZbikZNtx4KAd/UOFfSKo/vR89MtA0gSL2
Bt7RtwblmYi8SY9zgJrvcIi6aJSPz5hFh2WUXkB8GhrT2ZUjITHLqpRDynLfzSsNE4OjktSsM3vj
Lnylc3ksEFwMVRlp0pyzkEEA+zg58iuN7BfVB2eOwBpYkMcbLMa9bjW6PqXG3pvvvKvv17evVNbz
gFrm8Q0U9T4waKlpxkkEejWEYZMJrLbfsRFyydCnLMgVYEo80CJC5sBjZsPlIQVuo4GjxRcJpNee
mwfkz+r8ThkEQAGnK4DOI/H9MJEUpdHHiEKWmXsZxu9FrZYbSdAvdFx9YxzEJuqiPWNxODkv+w+O
V5rtbEc//LlwsD/SdxShMbMIHYl0u8Kshv13wwZqRNZNRJxkdnotCn3PSvk31XYk/vkqQL324LDK
GcLLRkSH8SY+BA1xUmTixVBA2ct2R4cCX9nwQLtWovGH+GupTWX9YnNhmEaLeBZG0oCpU5JKNGeA
80nj8JPdzNNs/mPmhh9TcMhLN8sbCwVMzx5eb6tgOXShHLfjaHoX3Z52aGTmr2NoUw3s+TvfpSBp
q9S5odDHyfjO601DFSvQAoYF0XZjkJ3l20vf2vHCYdapNTuLTUaI7ZmO7oowWFlq6LuR6qTW1vSs
mF4IK3+w/TRLJ4wY9xM/RRbM42DN6Mh9l5BmBhNePxr1YW1cIX6gY0/5GdQXbqFdkSHKgY0XE+Pd
RCwxb8lW5QisOwyABkmyBOrMAd8NtapSIaBk2AFpSOVo42XjeiywSIQYxesQb7AxFzwCxF8OzUiz
6h6F/5UXxuDnA78mcnc4+3IZ/lcaoA6vzSDOm5c6u+Qi9xLbM/x4OAF/PTW4I4BhFNWN/8PL+OsC
ZXk1tNel+16hJNtpnqrFiFP4m+nu0tk9kwqk2Q9Xsnz8ewJAL25pmlCI2CxCeQwRBPpDdhR7S1WP
6DbTDN8gQljIjJZ6+BFV1W6WxyrlBFE8zCvhTY/dwLifF5fRSMT8yHdFCectKf8gGmqWyIxd/Dsc
KXzf9FpWH5xBAAHV1AaJ35qKWoh3MmNWxcEkQbEsSfwcYgglQSInuqPjFblvf4yLDCRLx+3A30JI
60bG90IAFOstXcrukb8+ZPJuVWrZSAH2DuJAe8GLmWGP7tsmq8eTS7/wf98ucUtDJzG7r/UPIf5y
U1EUa+Y9SKmNlhQiuUHxO2v7vyCd+vmqTYZU77KV2oYurGLtP3fHB6XfhisL00ClsRP6P9omLNig
bxHki2ceytpciySHvFmCuBIQwmpboD5kdL2z7cJrRFRU4SOLWJD3RDqsiLA0A1HQd8+jAv8M8hYs
z2gZ1WQAg/eEeQWJsr6g/qSKZBe0t7IHZUnqm8W+lRgWc7ucvXssj4wLAF/66pMomFUQ2GA97Y3t
OkBjmYiCyMZBkWdSLcRntOSZbtFc0zIhw5m86SRt20uuJPFGfKnjOsHbSuzGBLJxHFKUt7FjmbCi
CGep9kfYfLJUSa/C0KcqAMq+usHYqYdImRgXt/kwX18FhRes4fMYKnabdT3MDtDcvfVyCXGJrP2y
R0dZln1fZdzEJ7oCSTLIsJdMSnKv2doIl9ZenFIpLM042UeUcE2Y/axNgq2bheulGS65uQaDdhap
1d+BLBkM6YjzwTBGIh9HORNb5eEfref7/xikRJz4y9NSCHjJrcVVvTXa1s1PaFhSzHX+10imdrFs
StjY9jNu+BDwBGz2A0vzGSAVCcjXvgJnpRKpKPozErcxdd0iOQynC8KaolSPvqWaQA2O5V0R6vCa
I+I15jAq4a7hEgKrOqvrPb/qg80yJji3jXSATmF1mZe9Cc19N7fZUjQ7bnNzQ5VvsvBCBUTZR9MQ
c6bEPPaeypv5tHo8d44LGAjp7VGkhgNdtKWHD4KhBtonbTGay3AtG8nvPfh3aLqUFiionH3fH6oH
FRJCZV0F0KTBAqvXZvU/qllcowoOA6a1iD3ICK+TKfZ2X0e22lOrOPU7g9J4Xq8UysrncGdnk9o0
/rlTviy9Q0Km/ByPgBYTvWSSgYHiaS92ZNi2xfCn9z+yX0bV2wFeu1pLNcDqPjsckZX/5pc4EiNo
22jEsJAEfPONb82NcApMrtyNZzl0UqFrQPsI1ZarRdtRtks7qckF70eJAyKO4erFk/Ox0S9dn0vO
DzKi1noWmC9xX/7K9lNbODFVRG7/AuQHIFGPpFL2ZWhWGgFw37UXENMenWs2VoXLz0mlymVXPvfj
WTxV7SqVo1oArlS5OB8YnsyKWaHq3UrsXL9oh72mNXY7SfUBvkfzpguWLeUjzogH9ClwZxbOGheL
Rg5krDiP3U5joikNNj7moOFSW3dKEyrTJkH+qir+/675MN1BrYmvSJj1eqedsUM37gTKBHmw2pMc
6p5zUn+C1v7NjzQNYeqxb55vb8AXIo4od1KKN8U6NA2T5u9Xj8DtLfWYk1BMxfITgJL3It+N4Ntq
lvOkuhXx1Xq9vyRuQQkm9LEdaDkpRmhGSWtvW6hX+HAOKlp5P2oRqgsTpBYDFJN4x6hEypZjyljX
vj4ibwKAjnZgfPp1Jy8xT9Pc8xGxDTCTSZgGioZt+NuSkpOkQNDYSs8DfjmGQSh+2SE3+3PrPgF5
XwFyluaPMmxeaPCQ3LZoRlL4RXGvK2NLX6YRPeRtdHzqi01BO3E5Kzs4mzhWwl0Wc4s81+oB7MIA
+v+VYlnyhWfkglgSVp1aS6l7LJR7oYCazK7jg06/KDHTnOVI0Kt8+jxlU+6K4+k87tUhHCHqCLhc
PocHRddtskDHVY+JV33/57LVoAolYHjlddkB9phfc7y6F8rhmgPDO9LSs6y+uStNWNOxar6e4lyo
4qe9ifS+zyGH+nIdaww3aAxSwI+YoilwyFi1IJXy4Yel8nS/HZ9j276Ri1e6XadkT6cT7ZiNQWub
kQbCjY/+L7HUJSnKBv3ppd+XppyEEjumhEho1CYlyfwdxy7EwCiaB2XB7M/rJLHNppWFoucsJaJe
4/jOAXz+yeFr3A3BrxRg1a5A00q879d+MMaer6oDHILp9mITFsCaQhd5NLBn9y3WhwNk5/B5LkhV
XDJlDctZAZughAl4LV8pdE2x9mXQ4Nfs3NdHg7KstoP/31E55FBqt7yaE8dRU+yo3700qkVJFlq7
LEUPNCfQg0CJ357XKPqHSF6vC/yYMVL5z9BK9hevj1SFbcvd453JR1dNd++cIgxcMXm6Xl8ZDJpQ
udtsheaXGmG0pIAsAf9RvxKsgfvgNTMcaZXUAxz8lreBPHLaAylNOV33wEj2rZpAaWWoVG8/bY1q
QRWv+ROPeRhD7807391L/nhr+ZHFsHn0pBhEb+rjI2nxDS2XGBq0bsI4cknNedeetQYLigH8JaPh
zvnzdMdRHiibz/4amsuEK6J7M692GkpfWKJFEetZNMVj+Td6nHHumRmVoTgXbvnMlNPp4DCP8Ya7
fxFIR65E6ANHYeoCr8YclNAylZ3ycCkST8rwuUOO1yExgPARcS0ipax60kTev6KgNyNn9i8p8GLf
73wB7vQ8ywDQJtcaHFQOUBsfHqHptBIWjTjMihAzbCyrF8SompGjB6GGcXP9fSSkoqAd1gkLIDzV
0C4zaQ9o0egwKMAahsMS6C2yvq5+cYqWFfeaHfxZL7x0JlIYXucjs8OHVchB1VxPHX8Hp8yu2EY4
bRkqBohBhPmelYvv22W7EN1jOisBnmxTu6wtFD24+lhZjY+j9iOInY0vdvdhCGkiFw2w0KZV8dzR
K+klQkLdwJTIoAu3KGvIiRCW/zBhIojhPAW5MnqtQmTlzvknKmh4crUIJTMlsdBIuMW0Z+1ed5b2
gO2G6s9j7DJ0qQNsOx0oQ0aCzqENC8ks3LRJL4xXcKwUcDrgkFrdDkoL2EL/lGUoBeMSBiv8h/1h
AoFJx7sr3fWmRDWXqsr4gGnqX05PW9BDi3MMYCDUC8hmr/LdEGh4J5m+AvqfZEcYokUiZS9C3CQ+
BlPzeKv76WIuzjyqozDU1hgKqG2vM7CqJwEdIY4dD0emWubuCaUmOdXQEwu5qQUnJOCb7rzAScba
tZIDWsgw6WKaVEWjFWHphtLI1p89MkEtotLdpHD0ny1Wn8pfixUxZIAmXkr5353JzKeKH169FjKC
lA81GLELA+k2UemTQLgI4Lb9h70Pwvc/fWkc4Ki5MbCWpr9B3yJu/jrUC1P4Oz3QffiVbAtyz/cs
2WdlJ1M/2v4Vll+qlMaFXIqN6GBggO5ODDSIqsC2gohz2QBBFi7m2AvtTkLgY5JvkVisDaGxgUkO
qY3X1uPZ2iC/K1K7hQ4RQpNf5VFZrtIoOK63OwlBXhJkvmDd31ZX/H0UTj5IWGnzJlRB4+SsTt9b
tfOHgI2EcAcPK+it8004H+CiLMGoqGkQ++3YdVCf1cS2t5LGZshH2PzPs7mO2FGXfXjXLN5Uk0T2
8Y7ZHhcE3phZYxNAxifaMpS7zkLzDA8hVgkPKOWDsTSl+CNpBecZTc1oOeakQmG7NREds38jvQ6z
HeEGVMwFaEPM1aMx4QytBYLK24Qq8Rr9EnzRLxAyFr/s31rW28uN6qMCfBdMW98n3AWJM/tbL+tu
jGaHQKjBIoVMJwdCB9c5fzDz0a/yLP98T/y6qvWi6mUdHLcYgAu03Ysxj3Ao4A0MzJvxU1A8tuOx
iJYoeVToqirBbDt6Dp96C4xBgkWM53DaS5mFKcTvaCVdL+P3Wf60945j25yWv8XscuBWWyx/nLtx
pqIA8lXHPxX58YBCCmPu3ssZKmV/UpHcJ5csPbVboEnWBc1fi0Wu1Dp0lG3N3B+xDjFNPNNRIJLj
vW3WbmYaS9Avn5kUGS6e3BIj64ThllP1K2QBL6tMHDL55E/V+fXCkZOYKwu9o5XuBi22qY44Y3YZ
3AYKGBVomDs6+KoZG+R9EKprjQtVec4BoVGm4sI15u2GBzkbHULZiIUxEwo9BfxYmVbl32+GApIg
uX+rpS4YhL3sbnRqY3IaEYhMKe0ytg/1XebGnXnwxFdw6iwLP7pLPUY9Ynwb0YafuCTYCZlUmu1T
g015niSexKum6+IAYjBKWcsFfV+SKSGXhAlI8kaKk078Bwi0QxB4XQgMHJ9IQ0IjVUgtqMTgO/A6
l5Ytf+O8t4QJwRbtCkSGGmlxFKt/tCvApo/+aYCyBjaOfCnRSy8X8UUvUBzieExtgC9FR6oC6WRC
+ypEgq3z/WXJPdULEi2Kx7y821kBKz2xPCcU8bgqXdMPsI1oEtpjfcqHMok0MCsgz21e0CHK7GhR
g5baDCIXIgOVgbGSV81VTHPwj8WjPwypeuJWOJcVz8NoEJcZdx7wyAsWpwaHwAjhazOaJyXwmOTL
sEEuqd04BoOdnf/kPALhJIlrxNyGI3m3zrhWUHidiuBI6rZtP43OTwSo7Xz0A5OTlOqMfEmgJLaQ
qLYH4NEef5m2V1/lPdMhCmuXbF6avSpJ+2pQ9E1Bkhk8B1WyWaOyX2VzHPI4o8xQsS/jqO8ZqydV
mulZaFojlQptTy+sExzvw04vwYIuma3mubFLNcXv463es79efkxmSg5/8t2pRMELRsB1S3XpV63V
Esz30lKabyWAtn5ugxbQKLKxMAXu0q3/9wDv0AadiMJ1vmsS+QizEYV9e9OZ2E5N8N4fAgDgmPzP
d73mn+J80YQxLMFpNIC6UdAuTz7pnRhwyfbI/5g672RP6gzAXC9CtzJmRuosV8eAK/eO0Y/uzhJr
CysXqr3PIx4QIEITSzaZhqTsknvcXZxhwHVWz8Wo14sZz8xVup7Y4a++dlii6nLEsOdPWkOL+08v
jzEOLHf1h+/omDVOwPz7FIywQDKNw6+WLUt3/9Bo7RDfGLH8MKS1GZVOpDLF0yFN2ISiv8SeOWY8
erPMFVfv/JqSPzmHbHhnUplAq4zOVELOLmaIQp2KXFKeCco0RaaE0qz17c3j4TYgmP7/nx5TfSfz
H2kptspYI9nx97P0ocumqUggXnaYjLAPU/+RZrksKTJpwxBUdq+YSEFcOa5aaYOhlwtOa4TSUgWS
J4+OBFhdjVCu6I1w5ueElBAu/H0k2cuD3+3ZNiF7HqmzxH16s7Bjjwcbe1cflMEmPGOqQafdAQgY
95OAF2CiowfD320FbBs9wZfkxFVRtMJb1G6QHSmRADkQ+JGVn/yG5nEQGoyjIxxmR899cdZOTf/z
mxNYVsXcZ9+RZ9aLmjwmE4tWGQTZ6tOJ15dJG5ir4bH63BfKNqseCzyOVAVCCmvtTHmsteoYobJN
2bwaAHQ3DIZmdAjvRyhH0H7eoYUjGYQNAIWC0Eba2Itr5yMnYh9eyeZhfV3lq0+9ELIdwyydsViv
tFevWkCL519glXzsYkJxl18Fyk7y2pb/7eQkaPWSkGSB+u7qNsx05/NxDppK+70FuSx63xSMs7rk
lVuD/nckWqcU9Yy4tT47T/v7yyW1VtQ4zHqIAVSk6rW5hDZS+DdjLF8Dl+6M+CU33EZcOWyq1VIQ
upsAKgwaigs7sWtBhNoKmqaPcj6kQWJzowPtxpOVhS4HyKPr/egYAlzH+A5GBdWTv3ls0nJeiYQ2
RHvASBxr8ZfueyDTD0KfumsjCwbx4xTA7uGCcXwb2QWh3I6EnebHuMdiSzKIlinmgNcOB+/laBzw
zSnA4ZmIt8Kh9k62gkWSgnTBZtA+HoUTO3XZJ92mf1GExKBGLgKxTMYVv3bc89WdlRfZw2W7ONN1
LsuGaXRtkLr45EONSUgGGg2d3/HaFrgSTG5lOLcV961Xpfn/q3d8EroB3491HLCe5ncr3QGjmRIK
jubt0Rjfs4UuzeJ1g23uhgluzWbrL6bmXl/tc+wSFqzzyLfHHw5nE1+E5u+Z95D+iq5WiTLmKEgW
eOda8JQ028NaJQzL9kPfutPbVjq92vZ9r5dKX9fw+xTWi2XzaIexcEs50t3WaECHghmOqs9aLSIu
FLf6DTfW4NmVoCD/KGFxWJ9q2X1BrUcUbgxlh1Gog8CW8t7Srmr52m7dJoxbQY11sI41b/bWGNFa
GPaUPQR/LXcDcxFabUgld7L/RIuMx6GdTtX0NKY8eWUNKxGei6jxJLbxe1XjMApOJ2X4x3ZTyF9+
6Wy4amfOP9TR2TU/21zuMJrwwmOlh4cViGI2lEPgHW4mYPe326mZGM5Ws0THFYNV5Z74YU/ayl0Q
hUfsA/bWFQVNb9on+KyDXz0gue6Bt9vNooxJX3JnI+e0/waRNAEJDmN05IoJ26lkeSsg5jac7Mu/
V34EorIecIXLQWibTeQdoXHcIWwr7R2XbHM0MeBN3TN71r5D1wDq3Ehx2M0JN/165MAkSpdjTc4W
dcwLOZovmc2Defll+2XP3mq13s8QZrVgxuOuiiFOrAUV8IqqA6fPuwlgna0oyjCSiBHUD4/o/0lt
K87+3U7ZozorUinW3DDqgcPQhjAhNTdonP2XWZn/Pw9ghSIGSrWtM4hle42bowcl6pDjvy8VYA9+
90xCCQG2ZNHVijceaBo0aqfWAT88IxXC+cEsB6N6lnVgeSI9WJXRTDf2G5jp9ow0zRx5Xhi5cIv+
nwPkVj9h7X7ASzZMg4cC4JVViK3QbrI15PN+1zwN3qhnhP0oHE+KRb+n6SdL7RmfUsrEWteiLYpy
RYL9wPhthVM39JMHJKvKOIz3gc6GKPKwRyMJWOWLIuEcNVu6fAr2KpESKNhJ3vHGAwdJ2FIw/Upr
60ZeIZTF/2slT0Fg4m0BZNCdWGbgb5NBrO4FJsIQ6whBTNJ2kyOpWBPHqj3UQ0SJ+ATbOWlDWmYT
5T0K7LKj9cEGbctzp+cYl4DHkOqEjlay3UbY4lNeL8/Afn/dVVQ5XwjfV3j9RYKcjbkoyxidbDWk
kMlsn2l93eyAvLuenlz+3vx6EOnBOLP2BWUxdnBBBlb8Bx8bX4aAZOSpWIMz9WUHBhpLOXviaNKL
oAHgoCwfDEfX0FpKvpRRxpcMf51MkT2m+UMoDm3aWHehXhNij/nlYgOaxM4+9Wh/pgQVVqqABg/S
/aUvHoxlsoS2SCQlDe5TMipqMX2vR4jYw/rxUumEPuK1w5JI01jJsEMOeVy4B5zEmjZ079Q8dc+A
6lCStPKSRMjoWyvleB5VLDWtnQx6+FdR8s9dj54Oi/4NqMRxRI8o6qDC/d+jBSwYgS9r9UDGfy+7
4vP34BhcvabPJgdgZF7qkoiANphBFQZUIo28Q6NvbHnWdHmeup58PmZGTWEtA97w8ZK0T84LLJsM
v/akLPAtcWENBFUTc6pvf719sYIgAPYSoPfxg1GabyB+9e6v4vDtYzUiu3MY10cCroWV4MpSD4Lk
Ylvh3Y/tgaRphEsZws/6HEobdmnnTzVus0SKl9lBiG4F1EvquhO6bli18AXHEPdgDkjb9sY7NbLW
n1Ih8EIfZ/rTZT4NnNQIGi7OOtN/P+JNEtw7KK9QtvuW2MPklpNNUA0ttSLyfI0v1eJqcImq+t3N
GU4gV3ytFEokYSq4dT7HjCffl9dM+ev/ERU2kokJGYGc1aRJyICdsLzT8IOWMp7VWqxNghaRg457
qopX30d2Jw5PIKrQ8/1xJPy3JOp8mLSyyx1AA5bCYTKgH5AORU2mCbc5r4CcgJHdC517tazK2vDH
GlH1RSL3U2eLPq4HE9XtdlkHvbbwv7SeuXtduJIJCvcHHvhgt7EoO00Y+nYdILeLf7E75EvdE7eL
befhqPA3pife+R4E5pcA5tr57lG88L3z5UjgkXfVsFZhOUGyIcGG+cZRXpKuuy5AnGByXSRBR+0o
UBKVvdr0D6QTebUhbO2aDhAjCBjnbH8bo05kBkFfOLVNusv1cKvLBiTXVGk4z6tieLyWNYSCEmcO
Uew5o8GANJ7FiPbKolWbQhTTiHlSFkALzpRJDmhdFbGM2dUnG+KGTG/KWs3au52Xq1VlEOBZuIGP
HgSUPKufEQ0bIAWlhtR1Fqv7gvQuQZwV953mJfozqUJpxP+bD3+7/Wy2/ynXbn4BWlri6f6PeYLW
241NC3p5646gS6WiFbVNbTqNja0VxeUVcUPHK/I49z/foEKpPP2gf+F+4G6iXMMOXTQKU0bloH8q
jQ8K6N8GG+zCvC5kNiGlZQyelCgM0jzaALdsdgBshRmGblZ1XJZolzFYOSyUjcoGytYyWsn9sfiY
F0O5tWNbY3YIGRDaj5z23QU+oIuSrodmrZTt6Kz9Vw1iJymcVw5GiP9jGp+CI16QY4zJzdXL8Eyh
4aGxrrEszCSxQkztIN3krSFjiN+rID8Y259R0kR0oVtloguUL29OYIEN/S7ck175fE7SkhumiiLB
XaGroeRiLToYCohPGmSRgMzyE7bUQCDcNbe4bFzQM0ymvxFV91oK/SfkAY4PO1byBbHVaDAUzRGt
HO5PPjCbzZVl+oHVjXIMcsbt2Fqe/Ko+cJK38szNSwg+2dDvzEHg1ye/GcFeMH3oQz5QLhCGP+Du
OJ5CdpNuXHR2Lokagc4fTRInCjpNpBJt50ejj36LiPITkCco/6J/vQiByBU26H3juOMI1kDn90ny
B30fACco97MGxhgffDlX71eiVW/TmKrUufyf2eI/F1nMgkjfGB9H4NvUdky2dHjxqEl0jzqR55AL
kysktm75hNcdM1uZWb6vbqsqZj6f3/xK9b3aXol0HEHfbytzkx7u3GXVNRQSn+8SKUY3COJvjaPl
BdjQWFBLXFsKEWWrY24KzUOKt3JWZhwIM56A2Ve9+VCbLpYwH66xON55jb98F6DMe8V7R1n+OVqR
Ms8wg3gd4TdWCCfWX7KoR1HSQ96CN+bd9/jBlktxsMYtaHwAW8YQmKgEEv4+LKB1BgHKyYHD9QZk
/5GS9mA8LLWWXsiGau+mOVUPrW6yzarr2BX3kw9a+97ktSP/50XdxCRIrP5ZrBXLfF1P1ZUmC6sk
zdmHsZE1q9dY6SB6i2/Bt0a8jyk1DNkhq6ovOp+U4IlcLVyMczgSkjMjlVx5uMz6PUwO9sWFt8aW
GwBYBOapQ3AsyuEqwwYYmA1wTPEIa0vtgctl1gPH5LSZ4vA+6pEcCLi0yY9ucy2aiUFPGreromHj
9ubPXpGEZl/+eSzjEaNwMvyOuItvvCLM8FA0VATET2xGqVrXHPFYYD1u2aWdwKDD//SA4u1H6/xm
B5qGXC509iPXKBW+4uMeJMhDi2iykv7GJzQGcGqwrofkDzzozQwuGclOpraTHrz6WUnF/sLrAd1j
iBEyAD3FBntEV2d75bfZrRkjoTsusBSHlT1VPWIBsh9ozsYUYSuL+IhNW4DL0mbkPpAEBniPKzsi
2y/B89uHLW470YvyRLI7l0fqHDxoqQPiIf8/RdLnRGD9eMqXV2L5rQngFu/jUSKcbYXbAp3khhw2
KTretowHeIos2REwQ4cGuYb5siFL9hFQP6sJlCAeH0tgAnGDR5iF8VcF174892Zxpvpqj46IpcBm
9/tozkrAmBeHBrHKpAeLqIIx0WquuzTaFnQkn+LUt2u/AgjiK5HnuLLKIg72Mawi0axkHPZIh0+S
sR7oa9N4sgGQEUjFiHXiNWodfhz2z+Wsu3lW9O9HDmcFzn7zNFW6fcgiAj8dePLL4NuJRCNsz73z
mcFYoPEOB4puUVVhLmupyRxC3uta/s+GcvW6XOYkN1xnyhOGyoQzdZ93iVxaGhUXMvGcVWrpV/qx
naKcabQxVCAKF7CjhjnBme+SW0Nm1OBu6N8K92m1eufxWxuRgZaqfm5k/1pl35W5cJZU68g0soH1
+MPKE1GuXSHd24SZKt5Nf5+K+5Otcr4LhnbV3d24bl7zJfNvoYobeOA94zK04Ofef+m2QZJbTulU
FUdWKrxxXYfpf5OpyOXtefAj2ojYuj/vL2ksWobcLHt0S/35OG7NuQ+WZav+4Ij66ThHt7uGpG7N
oGi52/TcxdDppykK9zr2uWo1zdgjJL4c37rWPKBNzT3Az5SV/qrglUo1CI/InODyLLAbjTPj6t+E
D5l9gcZwzPqWJm24yuJGN4b3lhvnzDqjHg+UHh/QPf4QWl1lGxqmOll8Vcc6uiRyP5rBFH0yzCB9
PZwlQIwsthZHEksZ8XGPloBVb7UgAiSrlhn52F+xZud1Ty7fjWnYIwoDxQk7c0159qIsctopIGoz
nC4Ebd0Orm/sC4qZxjpq8MdajpXBzHWqBBHy/wfBnlpBa7moWosNTkln2GsilYra6h71ZS/cJxXr
G5+Jro1chx3DnbMHBNoCxSk5lAZXuzaxgl8VQpuVtE7GPMxJhwqXhUJFB5/cyNVjcz7ytTur8gxq
TtMx4e65oTFeE8mTI+VUHCTVKLJw5iuH/D2lgPsP9mhgHPwe5MmZNGFC2sY8y9AYJalrgorL/MSo
CP74HrPUnsckV5lRCSqySkVcJedLT1JnO3nuiTa/V3YXTyOxyX669TsEkEURTWQ/FvMGfFB89L+R
yoNZvGoOgZWSnS+yO3n2LyZZtQsbjbYJJz3xNoJL7KB+M1vfOsuCJTGbxPTEBlWBBbogzHWro7ga
FST7TrT5lMPukGkd49jJV7o4Q4SS082hFB5KVFMPXaBqhCKO3SFr0iBjqIOI1iPP5rI0AESChYka
betP2H7w0deY6+PMFOGsfzJ6JE8d16FRX6mSSc5QFejQtsQEaEAz0TD328PwuqvA8qPGgdlrIQwt
OXH/uHQl/rtp5MR7uynnZeylDmxHyHCCqewPSDt6vT/W81opRWYQ6fNjFvAbXv2OsVuniKlUBagE
JbAWz/BKuy8Dl67Mf5CwmNjnZ5IRYO1jrgWpRogp60dnZEVLXQTC5mszX83H2BUt7QzPcKfclITz
O1JNhi6VPbxM9zbxS6YWOyvIlj33cszXTkkbbFXYcEU2rEjkuIA6gnttxw5sO1KXPLM1RTEPBktV
F/E4NhrbQ+ecBAOEbIfzbS8m21lnFvwlkL4E90HwCVKVrz23NP8J+okNpgh+ONbejh5zBSP+qJ5k
VgdckWn8EVAhDbE12vtOXT/eahhVkQkO1JjKQK8Dyqd8r0/NKOYvfj/p5dkW275BB7MHanxxsXlo
mkzg2iHOw/1MpRAZKjtrICO56jags3cKdz0duH0HWdZJRnw8m8XOVH/Re9UNWQURJyJeGPf4cBxf
61xdmXr9uG4vNXBnYHDgPl0b+GJuiIvatUvkzRDQB2jmjiqjUN/2qFZwCWa29QAcdwUXaFCnTcpo
3rT1UXSEv6ZjzZmAd62YzXuFyShF4k7bijdME2TuEucRf1hNiwtpS51GNlVWFiw5la7NW7dRZgIV
XAsbljpUc4vjrF5viV0b5xmYpMgJL+wDWTaYN3WaT6OMK1NT7ZYK8u2zD8/yKVrMb9owea+ZDYrG
W1nSd4Ux1vxQzRnw44/sOhGvP0bbWA22VCh9TA/R0xNHOEErnhXOpAieSlEA9euWPElgWk2/qvCB
QKOspx/k2Dq6jjNizwIswzkkjndH7VqL3zSEhXsjbQainY5+FFMOsyOqJd2XsvkFq7rEzemu/4sP
svnHpHk5QYTbeNYwhByY5ZPugN4rm8uQud+atrdALskHe5Zj0vdDoCpDyvrSo0m75UGPf2Da0ABk
8w0DXEj+MPdU1mckDut1wAKYmHXPGArBh2VTih8lSvvCAmvncTiA2I51Rmkn+GvTGNy1zcBSsIDk
43OvjviYWg2sBRrNYtB3usq/qD1aK4u7oeNR4zrQvO2J3JigyEcIT+7l876X6Nz3EqiI4kJVp4+X
mvnMJmpkdQ+XeyczcD9/cMX2X56QGjiWkQ+EXYUDSZoTNufdP5jZwuOlxUzf+jZQ7bRMtTioJec8
Wsnln4Y13RmjQ4dtkbAqc9QJcu+Xe9tkfgdbJUtxxW1e36uIKyEKOn1gY6eVhIRIy5nTLv7mDXC5
l0AyxJe1Dk7AWB6ysSfq6EYzgQOhOXRHpAgDQG2aXuaSNY4TwAojZPmbdkYz3JHZR7VIdGUmSng1
Ij4T3wTOkol2+eg3av+CmIrqaqndPWe/kyv0EBT+YUWS647SXh06D/PpGyHtPBGKwsBMRSAgLkGj
jRtmoaUEjdsCAhCZjcezt1cMXYh9BD/7dRcM9uYhkmmusvci0eoHo/ejU0uiQ+pCvK4zUOeNm4JS
tfoOnZnOgBoM2jJNr8hevam1W8PXBBYEQ6uHKVmPXBwnBMQVen+AuCNTZ2UO/F2oOeHYM+W74AYv
m1Y1LMflVBbJZmxrAHgDQq62XXjVG3GymGE+T2LFd1/uSPdVTXXfyHP4fhrg26bMnQwGmd/wyWIa
YOxMy7HUvM202KAs4WYyYeb9maAWTU6Rulc4aG2E9HEfSqk8rxsIjZIQdl/FdsrpEGWnf+VvUbn5
mM+YyTtENR0JgBoBp4Gc+fntaab/QI3N/+UDnXledaqHfzGGKEMx+cSAq+NpOUPf24fOft4kp723
C9dLvUF17tnmhiKhxifyLntyGkIVTjE5AEsgBYUdoNQkyHGzpZKxokXA7zSELki67UapgzbQASJx
440E1uUEI1U+Ifzp0XGCoyGedItzESEhsrYz25YMp/2I1XMUC2P4PKyzDwLwJ0Zr+xXtK3uLLF2/
WWamwWO1tDTDsdy6/+mTZSybv1UzRN0lypQTzwEfKqQs2Fz8fLXAQDjN5jqubmih9Li0ttyUyB24
aS65YG40qfE3/P26Bn46449GE1AbE8gq2Myv2ipfONxatCNftqKKBmzZcT3b8Dw0F0QN2XA9wmmz
vRWY7KZwFLAG8SIHpUuQaleugUrZbQ4VAojGU77FBnBTSsyAoWG7wfL9W++XAxj/+DDD3QpgHPMs
6zK8DmarEMiPYMOAcMN15WvaNkKK/pK2lnr4nvDOC8yG1y4yl4l5epXWPgsBCt9TtkeitAOkxXQF
yekhtMGDtnP5BY3nLjTKgHr665ViTcNt44+73iAe91MaYTYRY9uYPomNHGKnP9Xr87cxyARzUk4/
TF4P6qMfg/GoS2ELKa0CxfwVkE1NPeQ1YSdB1UH3QNSGGIUbir/3CZB0ubGoWOmRnPYOndl5sACM
9pwJkmjDp1qyWA5D4/z1imt6Yw49LXtjyWl0hxEQZQiuU/PBcgwQ6NJiSW7N+WKlfUqEvy4QTEIC
qHfpQrbn/qAhGdyBX0htBuoiK1+8fBtZNQ0U53y8q18dNJVkVJl3OsK6V5IfkzPSjGWOQsJacY1V
RFyItuPRtox44qe9ctdj7b8=
`pragma protect end_protected
