`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XDzlgmL0qhW89igS+AHsxvglNgZ9izd7IvdTrd/yPbvMHtGtBRVc/ZROmwjbDM8rUZOoc2Rs7jEP
F5l6klP5/2dt45U42K6706CXizEE57p53yX0zp8wvTU4L9whWop6P7ABvgQq/UlMZd0ubJDK3W5R
lT8DoVILNKrTUpdIJ45SWlZVk8yoa8cROU9V7JvEG6SWUTmmIe/pZPyZHGV7gt/ykZll5iS9EegV
6DvEleh0u6Vj8tLAFmDJkZ+drHwPGTPbEnWLf/pXYBaKudaLABWkOXGymjFP4rjMcRTzr4VW1JKq
XH4yqgoII9ZNGbxGN9fAdn0JTT4oYkNI4Yd1Lg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="4xSu8Fq7x8+Q1wvp9eYDbO6Dm1FJ/jeHnd9IIsC2a+w="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4256)
`pragma protect data_block
kCj+UB6jllZwlaLVCfeybsAnbmxmEju8+WB9U0m8x6E8vC5H972PNyyU8TD0eZqLVHbO71IWMtMt
lXn++1OiEGpkk9CGx1ulv3Z5PYsMJbpWG15D7ZxY01HkND3Gi/If32YFcujn9FWRhWGgUhEynbUR
1URVwEhJnktcbgWO7mWrJ23yJXrTnk6x1De4GE7RA3enkY0pk8J3MzGa4D2Ikk6nFBIvGIYy0Kq7
xasPgpm6B5L/O2MCSd4oU8lXzze9Iv6Mgt+xIjJv5z8nCdKWi3tngENJ5gsKSw2yHdLvWp6NtocS
M6lCW1f5vCEHYjtF8eEPh/t2yR41Z3e02Acxi5RFxPpLvfjeosYIhQrIIUoeBEuidiyM1Bi1IXYx
D+PeJyh+voZxGzvOv8RUEqYl5MpcWgAsCSlg/erkRZANgK+vmYfw9ow7daEs+M6wh9+89spL1R9Z
r8IV0/E7EPp9YYn9TmF7vJq1YctxtiYM2Psqs8Hi7GR7hIx43UPt9gxmGwidJv+S/mzi5OmW+J13
hfWIOrwRPhzsXpdOTSYZAp8TJc/NPmwKh7GXI7orB/JsxBUmzBJCzKvjoAQOmMVsgZEDFKt7jNR8
he6m+7Df53xaA8e6/n6xsfqsqvKaikwT58vSd6J+Szmg0pMzs1DXz4cPrClyyOEo7Az+mUO2V3QN
j78b7NxULszCUrWpweIOPSaAIxtq4yXEgmrGThX7lSbk/KQHBwXFORB0uVf/592H5Fvhjpa266M/
IV3UfCEDUNzJ/iYJqybqLmZhFvGxGW4etKrt+CWR18Ef4aKlqQHC0zTx+qx07lOEmQOUC++/lY8r
8rsbyMt3hhYoWZLdYsyXK5YYcjB7oZ+rTK2Lj8HmTXKyYrkJJIHmOa0YWJZMDnCgPHC13iuz2a6r
3CHnDVlJm2SC+rKErPiNlT2oZHIBT39VZmjcoE0MDjFmEVZRECwMN4wFxU2qAvtoF6yN9EyYl0SZ
0qQYB4jwfOsr+0bREJz+zX9IvQN8KQwjsHz8zVLt2mjCh0VTnBY7VSyffgARX6u/X+zIFKvrbFbu
2yzagCMufscFmMWGupQ4vLqSHnxz/vezB4lR2JRkjrA5We62X7+zHFPd1Oe10Rx9JUmGL7DxiBgC
XmUNguZIyjR7dW9mRv9G4AFaLinxvXFYrsow2Gj2u/OMM6pg/2Fv1dVoKO1XwgS2K1qUvoHYAfQF
ot+isMH0s0kg8dP9qvqpCHld1jNUUL9eCfAdW0zYsNxOEHsHiPxJSPYQ9iiKYiZoaXXjUp/RI8c4
8e69yCCvugbk/MaFnn1WjnlH2la8BegPJwSZUQfA33rQzJWw/wJgKPKyXowz/fRzoyUIAJnhWfMM
4/kYZOK2oePJSHqIAHrC2awnu4EBfDaM+QV6F6atOIK01UbfjK6yGSW9cOAmDYPUGfsb1mPEqlmP
A8jMctPq3GZPVTcKQTGKCkkrmiKrGW7IdGrVf/HkzL33sxLqS0HUvtgQfURp5b9ZgdjCkw1NTXCH
VS4N3PZv1cS+Jx3i2x6h6f4Q7zRunO9xVmnztgX4OH7o+SwiFe+gUZ9qaVd++7H6IIA1fIg0vXE6
Dd60REWXy2oxGjdaHd64GLJ8dMRiNQAWtScKOXhzSmpCRdWSXXtE79ZoQiQhEe+S9PKsT3lgi8B3
3auhMEAxowtduo21A+Whz5rioJsfVnl7ysGuYBjg8ZQsl+kw+w+jdNkP8VK7Ut0NTSBNpUgf9kwG
z8ghoFcc04Wnl2Fv+i74CFPwupOKZWkAJ3h2YQvzTawjLBkGQE7SpEUakuL6/5Alf+qzXwxSvChj
upwDh3tjZHo5Nj7+3JI4C2QILC9W+rFrUVSYZbndFRzvpbhDua4dAmhQomke2m7YEBzY6QEDnkBI
bE0CgE0K4j9E4AhndCi5r/tI0K1vO6y2Nx7ko3Db1q/Be4WrQKZWokzJE4QP5DS0dvXRUcDRQzIE
kfD8Ql11HRmW3BqaCPo4+5Ro2HmaIewVyrCkiAJNRF9rVkZi+z2cIcSNU8RucbOl68SksuXa3ohw
+J5cd/hcJwaGugBwrxtgSOeqKrqmRuu5st4do5lbOMn+Ee4komE4EabvlOQctA6uo6gPYxZUCoX/
/jGVsFcEVXm1gBH+C/cMb8PvoFCTkoK4kBOpyE791WXtfPJoPstTGxdh3Ky5P/e4FEBQUeBWVmdS
nMEh1dKQDAnBgLOCkBAP2BDv50PnDYcr/L5hWqDS/chhWXSKqK9wegFD/D5BISooC2UVN7dr3jr3
i68NzIhFnVNSZYvnNDdFejZR87D8O71MtWcXd1Z7f4YXT2pB6v52BImN0dVmi4Fg4B4B+50nGK63
RU80PZbRGq3XfTMDqecT0VayUouhwRrBcIko/BKzVfVt1nzyeU+1JQCrWRoNz7iZ6uf6hWElhK/Q
F0jeXQKcxK302qWazLIjs2JBl5clpZmi4Sw8P7xRILLtZ2dJww1LhW7yNDsAT3B/BMWulWNEeESG
DBYPGACXDtJyzxlW4XQ2y7kwkEmTFLxEi3NZVJIpAF3AgrIkw1RKba+pbU2Oi8hA1jOvsQtscNVk
gThZ/TI+oGHKBdPM6pxzf8agz2ImsiOccEKUpX/UzWFkmDcCyLH5DxoP1+LD2GcOO1y6xUIWBxEd
QewzIJrSKJgBnt0m4fCpXga5ZFKAk2PCjZEtR7XnQ/7ewknsXbd8qawWscQkI3P8meBaEaTFSPF3
Tcp+zVeiuF2lnDtCuxcktFVR2JehPDRkdU7Y9+tnqBUZXfIWB39VcdHCNSBpm++2EwuCcF+Fg85x
ZafVIGsTA52nfmI9e5eRT4JIr0xVQPNNEy+E5xk7i3lTND7HjaeTA6Nm51vSky39/t38tVW3aavM
ZTR3tcpHq7H3f1mXfqRfzXNXHpXvvggGihKpDF2EJ9gqyeG8bckmcfQ+cNFpmF9ENfuvnNy8FBsu
OQIdg6xx3P/CDeUD3f4DAapw23+yUL7byBUW4lbS12S+kO36ND1r2u6JI5eyIdf7koTkw0l6bh+P
6DwKtIIpwSLtbG3dkbmg267Ur8kYFYRAc/66XrvOxLGN7JdxZJg4a+riEKJHUj3CbttqkXYTzHc4
mUYXSF8GeTBLNu6o82wSe/lif4KxQuLf4X+tBdbkZj6a+8184GqQl5GRZvs1s+L4WRxG+WjWNcu7
tBMmmwmJqGz9MkI6ANjkNCCb8crpsdwSAFE1bKcUDjYFbZuCJ+PZBKRW9rBHRmFj3bJMSVx45VRn
P7ed7+o4lf9sSsI7SOzNr4NJZVczjc6HGLmjLYwhxeBU/dSEW9L7h++FXVKu9Btq+QTjVPBeFNq/
atJWqf3rtUj22fuhonHi5DdXPW9ta3aeb6yE/jpJpb+MCYFZR+PJrQvOHB/do9U3mVjTk98dtPFm
GmSfG05MJVIwfx7ZFDVchF8igxmiMIc+WaTF7TgqxBFiPhta8VKTan+RpUwVVF5ATILmagYU5v5b
nTaNFIeE1U1bov1KJURpqv8GamVJHeSla5dWoZTc8EiEQbHnfXwXypfngjpNDDrIgDj1UUqI33E4
ATG3YSbv1uj+lKYlejzmrQxoKhIzOisOZfdYJ3Sd4h1xDGkHWK8WY7S3TVFPjDr7qcWVKi1dG+sW
nc8CMOLO7ICU3AKFq7/O1+iry+aFs+hPckLxqFb66Hakwn1S726tuei0zeDgdCJgiH/CjqasJqOn
R77XfHzWSPfIVJZbxCh2bHTErpHuaOYoWg2Y4rULxZpMzTmFC5If/gxCDBYclHs6PfY6ss5DM7q8
8MswHj0NeehXLa1zLdzGQfPHwOKetn5VBkRntBIdLJeQRpnYyT+ju3sHXNwoDxIpaF9eMknFxxq9
O9AIwZO3r4RUtulfsfAvaq6RyuGunzi3S6GX9SJHBQOBNzto5UEsL8+DmAMoKFb1mItaRp790JP6
CTLIBouTVxd8rCazru1gObjQIZlcVj9NOVum0jl61Harj+FIs+/qyFbnVytTtPo8WJvUhiQGDo3Q
76wvsXIl2Hzkk5KV3VnjsdkO4xrSAuOHpsHZtJsHOl8GwYDXjPuA1wvCss0X67q/e0T1A+4buxdr
4nVswN3GevXFPlCfrUUIFkybx3UhICZ2snXarETEsnuaM6QBTr4KOJSAGDmRyUQHTYXK3YNsu9A0
V7YSqda3ogM/NK0aN9xRMz/r4JgFAtJxrKN7reIg4+LZzQUr+q5DI+RVop1OnUOBaudMS4JMGjOy
PGQEAatPRbx5y05+5RI8Tq1sBnn/l/eVTY8nJRmtX84jm5U6tpqEyFjxI/Ev28MO0xOojk/qBopf
mRxlWAkrhEBlYZiPyg2I4rXlAKT+WovPVrE3rwyPlE732EVIcG6zukC4aWsgB79pu/GY+KjLp03X
kVmD6zwd+qYKqWo2W/rR8yWoAAspqmW8cv19cpOSk0V/Mfq5U3Wob2k7PFPBmGClBD+mL2JQFAs5
raRvevq32M4ACQHhpbTAKYwM2KiDT30II/kV65yBaWszud+TWppiZ9PU/1CeTOa2YuYD6NlQnD7K
9IAdvvsqA9SjAmcSLBEYiT7cn+3OKQMjUikaErfVC2nssTc3n2u5wi42/1J2lqDbq9KgaUcblokO
OnkqLV97p84brizUf8ipOTwQ1N1ZxU9PYpB1wrwDg8K6hXYQeJyW6UyhTsBoqz/QtpR1ufY2QXDi
THazHvOdZP7dPZCyb0DlEudTVeJvf7fnYnfK6Xock+7vICeHaddJ8xaSTp60WRDHuR4NYk5813kV
3YetVe2mgoCcaJx9QueSzEEp4+JyL5PmQ5bTijMOFcc45Aws+5mg/Rl/tOh0DY75hqedM8pWVL1l
sgwwZeoplz2eICCG7+TMgR8D4MzkY+3VMx+r7sJSL+GTPu+JyvFGe46EqIv3tbEQwqXdcNarUJ7F
88mxD3G7n4zFACmfI6I0TOK8DpYOYVzFIkfky9iJ9xvrC7BS2otNjy84Kar2kxiEOInOOs+4qkhU
wVtpIdGmk8N4I5cvwtPMUSFqANLt4NlArqPTz850ZEJerqV3m44yZZNQeW6INNhC7O7lNWGMuN0o
zFqKfEeOWI3Z/41OD7GXYME8c3qBEwdpDwbr2pPqZfm4Ib3hB787bLTcDxuxw7/PUS8yoyPLvHN9
rYiFiWZueJGwu7osDhy+edZf7b5XfUmsedOiN2OG2uXxGTVFTVdC5LtnzqZq31MfJwG4MgJVhQn8
wCHRmEIm7CPDvHXbHvq6Mq53ua7k43lOJ6hcGIyyZC/GwMXwyapJeTnCh7vOUqZqYSF6/i3rwCAq
vB9HzOpevTGdZr/+n/kjGJ7PIc3ZmTlgVU+eTtLcmGSqHO2dK0HN2dluAJE6+d2woIe1FdcRIMMH
ghoV9xMU40YgWyMPp7qqVTv3H6UgYIPSmXmUCKswpUbQJKGmPB8fXDsyPSEhcygNPPY8R4eR3SA7
J0DJCz4pCx+lvm44rGnYTp6NeqhKZoMPuU7qgV+ctdXqh4a7umIbXijDTiThJgtefE43RZ4XUX6u
3LmnuM7u1/lbKHmx5sb2I/BFUjRw6NPSEnPCQqBYwz+NEU9Sa28pgOmyAVsrYI8jL92n5qYiEp9z
WxKq2AJ4bzH+jITo4TLNAtoVQXwfuU+/12A9ezIdRgWX0vKrLTk=
`pragma protect end_protected
