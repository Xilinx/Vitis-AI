/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
CR8vN7aeY7nINHWPNvDhzNAFV3POF2m+Umve/RSJdDqbu2DD1qCR0b7tuobi5FAPK8vfUyAJUYu3
l+3ZWDR23JET9/rBZPLwkripeRbhSFx7V7Ay+DfHaFILsLqukoBS3vJkccQgKvRWLLfEyBnXH6VQ
ASSrGa9RoA8qyZY/WyjpDo+bZYsNB7LibB9NVDWOfoxMbxWHmhgbErQgcylB4CVTW6woyBagUfvn
V8iVobc29wSDami3N8wLtEFc3B6nU/jZGDk2aBW3I9BBlp1JFda/WszLSW3u6fRFmQUrHPlf3J5g
S3ZgcJXb03QC/4pEQz8tP/OHwJYEkRJEXy6bTg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="iPWB71lZBSBUV8roxtJFE+uCtSOVKBCX+U4s9IB1WWY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2928)
`pragma protect data_block
bypxQuzwSTFsYu3dZ6Zw2tTxSLju/PDgzFs/sPY4DVEqNewGTBIHpBU40YVaF3Tn3mv3fTZEV0Om
pGClLm5+TKNvHrHcyCXhhc3OQ1QoCc3Lxdi4Yls+HB162ujNFSj2RvvwsgKPRZDi8OMW89a/SnXM
vZwX6gWffwRGJQKNVy0K6v7KC5mNM7HxlXhE+d9/UzMePIKpM/qZcm7jzkvsuprSe1SWbC+euPkO
nWtCX8fMbVfCc0XhvM2JEejSoBkPS9DzGoxje8SGNiU/DfUTGYTZuw1lelyIIidkH56RKPLA0IRP
RoL2tWd1DBbUHZyOa2UxG8DCqiNVXVu34Q7vTAADx4nbUr091YchKY+K2+DUcSDZhMoAJwpw0SVP
TjnM8/0fi6J+LA2nqKnG9Rlx0Omn0a7EdUzv5rIlNlm1DiaDaL8Xwy3ngVv3FNo4TYWbD8xMr2gr
LyCF0dfyK23J/D6VtaWZTVElYS/BF7MdwvQ7ysNjmk49Qn0Vzdhb0XKcQ68vPsBIE/CBx9aoBRRj
3XWTOMlgLuJ1gzS6gv5tKm5atePazVSIRl1WoWrkAg1jN3tPjB3B/Kzq09E3+JnO83XN5OJfgPY6
yDlUrzSc+jQtSh34fAG9EMtxQrw1uMp6xJkNpDXQaVRoxaekT9wU6J8E5t8rPWki7SEsrOoGndcj
rKQWCBRveYW2752Ffi98L+crxpvRcs9YpTTiBfU3dq4Ij1OUeZfN6Xf66pzFh4bb1OmRtZdnQ4+/
hyy4hp+3X++SsKUPOriAP6nh15KQVhKeqGEvIja+bMc4JUC+iePUXT+sgf1ql5cpwx1pT18O1RS2
xwgMgLzrp2NyKt/vSwZkWly4ROCRyTk1k5Ij4iobloI9SjGgX6+IAg0s93NL15CeBmF4k/5ZJdBb
i+id9lfqmYgUvEKkPc+44pvblB3uv4xFgVM7nLEZ/T/Iarph/5iSvFGBueMqgl1r3rPAW34lDcG2
EjQ8XqSNqFdUmDU2yGkIUWnJrODsy4m8v/MPuJgIBHMLEcW03NK6RxuhDEuXnOC8lgC+gh7Wr/8z
6lEPZt68Dg4rXvohuS3tzehEJaD2uaWQ7j6lwWhyQLgNw/TmgkETJeQ3lg285NErSJljhPvIImk3
RA4/D1fq9+izA7rqL8aejxvY6Y/K5b4Uv4Qhv6incLhSTrYen+5ySSEkptVxXWb6c/dd7PvuRX1J
lkq9suMg22FhKMHyLy2Fg5zxCTstuXHrK5feT+8cBPPri7UHoQgiukai8pV+CDMRYPrRPOsun5Wy
vZzhDCtVDTKBvbG+Kvw1/iRlCL7+e2TuHs67zBU93g1jGIMCPCXvv/um9mGRgRxljm04z97GtK5y
JN3Gf5LBh6opKO+BzfZXGxuh9C7fkj6uRJ65bD09tdfLZPQZv1d3/1Vxmike5Y5t0rmsiMpI5eoD
l7kTvdiO+CA1dYBdRI03oZvo4MSxxe9kINMrksh44GMY61/OyxYHE2ZvdHn0c41G24Vw7oj2hxkN
SE7avilZRpWK0l2vGjW22p3cIOTdvso1aariWu4DVneKlEZUM3MZ+uKyAWDGGIUpR7uk/h2MEal9
kNWpB+lJ0MIN0gCt+/7ncpmORBeQw1RBMyW3rt7nD0Y3eS6lo6t3QfyB6KjSZXiWl3BsxTQATSyM
RkwFjtUEpki4a+6wwbZytedBlrpEKrsqR62fFcaxHK3EXr67o0P5CvbjeWIQrBWuv3u0AVHX8gzQ
F2K6qm1FOn0C/wPE/nlROGzNT2G66f/rDJRkDqWEFDZIeLr6j3otgEkAn1Va8VhFHL7hS44rxKIc
zcNedB1XrW7n4FXlnhj9fiW/0gbk6YsEnGxc1BfPLv3Kr+kuD5Rh4yw0zXkhZ4+Ieocp6F/7aFkE
4iVd2/gVfoK4T2OdLkLkUC5fNqur56EIWt8DZAAkBnHxRn/lAKVCBHQG2q23b82AHSaTgR89mQKl
ZrxsTU49m9UYROKZm65vde1VQD9NkTUiPeBS02sEo9i3STrs9PnZkYYjxVWaXqV03/Nu4GC825tm
BO6YQFUsNWyhdQZms8UB0phB94JY/HqCLfofp3S/zuT0h2/6wD+hOtPiz6KyYZgSgI/A4nmy3xI3
J3cZnL5itO1uf+TFCZmn27aZ65jZqW1VeUfOLmmJvGPkyLexSzo7QDF5GVtT5CjJo5vzLzFmwnHd
dcZf80AY/ZyGH0nFve82wqXHIEm0JmThk7UNY38GE7xxIIaUhluf5thBdUOErQV2/+BLQz+5Lyvp
gO4Hk2kYdtnCJrD4Qz0SjBGOBuzsQ+iTBqZc2T74rAJyBWAUxcWknDK2Nbxyo3qSY28aTSFMPgWS
km2g5i/0XAVa6uR/0QzrvdZvhIdhCRssB5vVv1JnDmo4x4wmDcfTWnqxlIGwSuACG6usPbvVyB3a
atuWkx8bw7DICEbBtmlpragkMP5YvS+8yNpp299ms+YRp3AVzd73feZjJuFbvpZd87+rFJvzqVoM
R9NP7MwiV1rFnRjr+fkLHc9Uq0qiFZLhNZzr+9pUiYKEqTRvssoyuOmjvu0XReCa22StWmLfbY9k
LlexXgLFAYNpUexMNh8oBXvPTWA1QNzryrWSywOVPct7AUDnO2MrVGdz8hsMPqIiL7NT5NdEGZYA
8bE+5qg/CtdDIuAICa5caGD9iJaACbMpbyp+ajr5EfQnAN6sME5vVP8VODrvB7t3kGoE5JDE8Ifi
rqrosujAkDMyjXCY/4RPhQIjf8k+rrCm0S4LzVFYoi/MK7/I6iBvALzJco7tpnrdISZ4CCcMsvdO
ML0aH5Ey4p9X77pPtdoq7jW/L/ahqLSTBpdy7Yd3bxAZEvXgKmBBofebg3AX+mSbZXBQL5IbmvoX
hnwcMSbZEmfqzKpw5JNTA3L7mYnOrY510scKjPA6g9nNAVQixMW/phGGWnZq/a0CwrIybFFt/mj7
IB3srSh+5o3RCZsf8BO18jidD5UVYl7queJPVMciK/pGtI790D3W8AEJu/aJhefLLNE+B2KHR/ai
Ux8DHk+WpwuO3YI8itGTT5GxW9pDtJEdY5AZCCPUrr8Bfb8FQHu/c7x+VLHKjC7ZZDwh3SKd0wbA
Vo26hlsaA0QxzIRm+HBi2SDZ+B8S239JwB+HTVNpgxlp2C3RHfFHfR3lYxPaWRATRceEyFNDy5wG
JD6fI/udnfqoBKnsy3QAi3Fu7uZrl3ZE+ic9bTOIOGdqxQDSdhoZr60IeFD1Kw8M1xIquMhD73Nk
tmMGwKPtcrb6B89GaW34Iu9KG+oszgq/VhLoq49ggnt2rm6PNlah6mcHmYaY21iGXu/okRwHreep
9F/FL6JkUs38u5KBDAVYetQjDtwTEzK+XUTeCRFWlaC18JB1MVqQgQQa9pnPruNTjPDlK2nHdyKB
wC2mPs3pV0aHiVGPTogs5J6/93wiBlrfGg6YVvyJB0jy2cKl2zzyEBfUmBORxj2PaMBRehRYr/WF
U+xFgngxcc1MYvToVgpDyjIlX+Z0glD7RcWxNwQW9yfjYZ1J92SdEuIg1km+2RT+rxM6JE90375R
8Wbp6z0pLH98UuzA8CJjmUPCh4MSxWT5ytbkUYn+9O4BZb8u62FD5a4W8TYDKNzX98DTGPgC8T4R
0Rmk3v1K8ep1UgoG90sdKiEt4PbZI1tz21fJrQyWKyy1uBpg9pT+fbgusXwpGX9jycAHfyRPm8J9
ZxwejMHRtSXT9CruaxYlsms3serhLX14RjTCrJawXE8pNPbvMqw9wOnxDF09AqFH7ikGz1Vz5wg2
6TdHjG3P/JrR8bqddqt05Jd3UU7N5E4bh9dYyiLx8V0iJuVXbIsfvmGwfWLK/TIJkPK+/nzYWBKI
4BancZfAB0i+uEOOocFI3HQXT21T
`pragma protect end_protected

// 
