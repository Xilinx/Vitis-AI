/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
ws7Tr62s+jmqXtZ7WpRps02BAr8CNmW71yxPY/spk0bwb3dgSEEeyEDpltfbPzRxaNm5DG37+UKX
Wo6Z9oV4BwR6c+NkxkmgiNmwrYkq0hO+WcJLg2NkYTp8WeQVWNe5zz5N0bx8f9noSAw8hZYuIK62
z6rpqkeXI+EDBqHSstXchSHINm+3S/wVFLz8WOd4R5OcVlRId4QnGA/xf4cZBoDJEdh4rQj5vVaI
OeOkAAfO52w54GYS2HYK5Ymeu6O+kzpzioPSdAfXz8aGYMwkkvyMLKkxOgxQ4GDiyV9d51JkZ8hK
W4LcykTQ4ViDfZIZ9yqR9KlJNjJdTS10ByiusA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="CRYOiOB7u9yx/qgZa5JlS2BibZMz8rnfGDW7VrD+VzI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2352)
`pragma protect data_block
VroEqLLwJ1noFwm3Z27B6z5xh5wSHf+NVyI7773KsgkK+jWTL4uJlzgJaKnbbho1IxAuqc5/Yh7J
8VYY7TDs5n1SOBfkYJIHhmeVZaZ2FCeH9kBRifo2K9ObiwA+m7fwIklkKEZFOVmURtMqns6xHlj4
bWH42vahkTKM6U8x6Yv4mF0kXGh8SnDz2tcfDBelq9HcQy03QARrrngnkPGigZAIc0R+YxpTQjdP
Q5tGHswXOHnMsJoSHA8a45fKa6/OUE2EeTnGMPoXGdygecNcNE0mlR4wTlEoSuTt9hkmmZMD4KCS
EQ4vSHIixfbaWFkjAkuu1I933b4ahgrTbXX+DiJ2dFcr7M0YuAqICLRyJRRsdv6lA8s0RQXahQTm
DV2D+heAW5diTBo4dg/FCyxmzIFzVY3cKJ5HrR79ezotgCLUufyZV9xEyco5ea2cXjh7g+6dPsbk
ELJN+joNjP+GkQ8cK/PLheaBYWQPYmevZ3CSQW5TlbRCJzZRQMQBjtn4Ym83KOtdQlWX6+TUN0Mc
CmAMJlrlL+/1vSdLEORjyKKsK4JdHk3y1ZjGvn5kUT5KmJX35RYxPX3Xweok0iqw2S1of6JF1bLB
h/76WiQpnuLi+HM5WoVKUaSeMgNMtvPtIA/jqPmmvpQ+p0T8kDbIOnzOSHhKYNQvTpQv8ay6GjsO
uvxFvF+/yIt8RpGUUHnLkH0OkKy6sDMfdEEYVuZUH92/4htExu5mS1XFmxhnTrRmS24ACmzbRWqZ
bFbGg70DlLnA0ggTz8IBGQgY7A88uZUA1HRgOK5M8lCnBVXgC0ZJ1uks6XGsrbeIUZW+KCWqVr0i
rKlBw32MJNJqMvYG8JbJ8XZhrKSsq8cf9zpm8JTuG6BNj/idoDYeh9UGuivcKxQfPU2BPWJ+1Rsj
j7rUZlDVj6FkfY6Zrc6iAzG0joVcTO9x0lmSQHoexnqM4XZqUlA6k11x87t4UpUTyhYI2lVMEBvh
QzvEObdS0gG4zUDjChImVjK642OwrBSlJwn1Zu11QU3lKZxR2MjYYt32OPpuMUxjvi6gccxrxMiL
MejGCbtvpze6Fj9tJ+cVqHwDvUHFy3kBx1XszUASj/zPAe3UdYuc/m04yAoiiR50ngoe7zf8AwL5
XZ24J0tLchVBOmqe8CRnyBhZgkcScP9xfNJzbGNs2z5nRhpDKbbJT8wUXdgFmBtHK8yPFSdIX+Cz
3Y7Y46e8Pl+CIWt1UEUHn8DHATeT1U3yPvDBcvvYneIbbjQIMQM0aOuMyl3KsLMzh/O8JJHb/IKz
AK/86NbxdIKd9IgthLhwjT2W9yG80ZFp9YMTWAeMZ3g/pHUC4aslaMQRduQQVLjswD8wtXHZKFZ4
/AczFQpJCWcesV5L/lnAmtQh0R+AvOseDaZmYURvC1u09epIkY8dovl8B60+no0pNq9l4AyqURMI
NKicocZ8Tx3B5qqhl4TO4AkSiWXRaBoOfEIOrFqJuO7ScuqtzhgtFye7UmGYQ3TIl/SVRcRl9AjU
36R1vOiyQ5/+YApIQTtSskvQk4lW4BS5ZgROdNyUeRr3bVsLM/gtt6qbAbE31stEQlRSl6KHRA//
2RMhZYGiS/mi6ihsRyv7siEcjfS+eZGOmsRhvMXOsQhn6ZdQ5oUgBHKx9JlfYwHbQ4aIV2WyYRDh
RD1GvjestugY//uMQeD2vR9/O2jb/iea1xX8KUs7sD+aEjvYBpL9vSDlqt3CuA1VHl1tYdN7TC0R
yf19ZdWRGpl1gmK7oD77ugHxBOGopBVz4NRcE45bxiIw5BloxB2Nl1LmLU55vLDpWdq16p49Cdk7
9qxPTeX3PvDJJkn9VceGMCinYg97ST6AccVVZvFJX0PIzn+k8yfmTm/JBmEyUiz/6D9QOSpGWEtg
qHgld6XoODNT4adNugnVv+dXGIhgdhqkHNCCNTG21CmUKqemq8d553kwSMo1STCWUDS/eD/0iRSG
loOAU1106m8TofIbziFQ1BvG9foCqpKNbtZYH3DwCX/4bXWZdEvOt8ZznpML65dfKcGYQN8aFJG2
Bx7qbP6kheFX1EgDfW1OoMOCFM4zqBL8FPoDf+2ePzJoHThfBxuv6g1d9pqRpQ+aCUAolMauYPN7
EtRWl9TQ2STIVql2XZC0m04vzmZ79wf2pi6JJYsX/n/xIkhdLeS3guR5rPuY3PdLeo3H+8Vnbt4H
2ul7Z8inf3rn+bXACwv73dhL5DiDZTXS8r/odXRhXduZhRPy8hiirzq2RvBDuPY5KPHrnFTq7YWk
k4trgtFxtdRrf9403dFhWQZ4I+FQDzOc6tz0cuRY9BXOmMBsGTaTU286plyOGk5/f0swh6aShMYK
ye1yDpQNzZgsKfx4vUzcZ+LPJdlPxKqt8EAsWPbnu3lTU5dlt0QirzngdMtusyy28mcUN8FdNfNb
NVDOrCG6PafytJKFkpNlDC8/9W1R/+xjqKhBmi27zLWlkPuroWwh/5RIs/ELnEX5WnljnmYCvT49
KkE7ByXWhqFKZUjOAz9Ko0o9fZH3yonksLuibdBfL2z9g6GI9i1DW7tOoWc1QBPyM3BfISdl4fu8
dGeqlJdilMcqWUwwVwA5+79EEHaDiLCW/FOTBp12dQ9tGfI07qkMLtEZ9sksbCAU9kiavbRCQ2hr
zMtPjTxnEotXpr9fO7vR8jlIAQAZcorJB2HVjBUMQk9rHCLPWQHYyNItGz8a7BjUdkKaPb4iJZ3G
vxarCnL1/CuXj+Z/tfBQljemzOj4YIRDCd3D/Gi5T+KIJMNNjCa+Vx9hF1kVjjvfU5qONimfWNHY
COL5+P4Lr9Bz+8tl8RVc9azLlocK/uMCWFqTPt2QwfCnvvH7QwsdawMLDR3D9s7cA3EU6L8CNIzD
BgmGV3eVxgrHTLEx1t4lbNg3IFxvPxnlgrvtoD6WBi957r4iZNDldFgkO4mqU3yn52ZZH44ckLnK
cgIEZt/0UdmeUSE1C0WK97cN95MXHKgcgmdjtT2xVSygXoMn3Oy++0Mso9QwbR0FHZgIzEl3IWka
wDMBHdUslcCiT0l+oShhw586dDaqaobQnGkfcEBJutNeZSO7P2Yvle1NL59olIGK8yT3WFxJmoOh
7J08YwA91HMNbeMKNbmP
`pragma protect end_protected

// 
