`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
XOU04p1U8l7ZkPUhVYYigTFU6V3JKL+kZai7mUv6H2C9REWImXn6gldznG1KEWVMEpOOQamYdo/x
0+V8pVt2ZPG2Gs/W/4exSUXyIIrB4KgsyLZ5BjkCURDY87ZRHd0CQZ0e6i9DTF3ZhK6lGpiV5ghq
UGj7iGJC3rO6jJxGJayuzr3X2k4Ygrcxl3Yk3p2QPOiL3l5uaJLaWUMVqroGLx88aMhnNFKc0f3Y
eFRXZoxhIHH0874rNEDR5R7COHS+b/ie5J0Sf2QUX3Qn8j1vOp0e0LPmvmCAz8afL7IwL3m3Xq9f
NnkTaPo905svfuq1DpK4791inHMfwdsk2KE1Gg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="197x3mb6unpRkR4TRW/K4O6DSKiiyVWMnQVxcafkC2U="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3712)
`pragma protect data_block
giGA109OWTgnmloyaK8oOG3UMqGwnUSjVhbhe1UgDXDlKruOCs0g3Aynmpxa8mp6E8yQe7RyNgab
16/g8Sosz91BSsTjEYEntnTFhKQjy3hZil/LAxPZQVZ8+KC3hNB1ty1J3nLCMZ+YE/fyxrSYxwi6
A8Law9lVnzoe3WuHFDpmuWzsHTOxacazNjb+JviQW1EPIS+VCGsFRWgtRMl8lgAuvVwi6ZN/qVg/
B0JUp7wpOq0WtyD9pvR1q7g6fbmQq/E8hjqitvuHUMrBx5FkpbLJCeI0Yf6N9kqP/3FrTI9O83+h
9LAAO+BPSm43hmlj0FGHd/xnfWZ2nhlYc02V+FD+A1TpEQArNgTn9hyeOV0aUmELZZTeqD/Ahflk
ejdbdAGSfTlIIU0tC90XaczJtp8MvfPQlPYQLUnvk6mtCCpWtGBSnMAYCLSkRMd2RRBwZJtsE2Nx
6okIEi5OCJFCZGrxU30t1lPOFcUt0WYT0B/4pPHt8PV8yZ/JfNHuBrQ0NBc9FnW+4QpVtaKpZmPr
TM6sg/+Dk6HAGW/s9nROFztwx0GCUKfSDuyM184nQqPOON0ZIImtZ6x6avoWGaYEq4Z9VwhSIWRg
FWRmbuseicPdAQ51xzqtmOYLox8zCE0qI8EJV7+JJcMqWSdp0BIbaIkb157Ip/7PSBlGVjtAQCGE
Fkrc6b8IKlDEOt67vEr6Xex9rbS8fZXfy/EjQf7cfGoHq+OtGCEFaGS9Td1Q5Vf4XXBaMoV6Qy9/
vsZ43KwtqLVNGpOe0wqpopovluhcALNh57YHVxMynAChEAse2UONHfpMv9TeB9LGM3Mfygl4N1/f
xsHeOMtuHw7LnwP9kottkmZHLtA7i8auf0VMf44X2opVEddR3542bs7kbrbZ8wXHULiG1Jr6hAJb
3hs7NbOSmHEGgzkNpNkJZIgke1zydw4GpYQ1GF1j0bJBSw8yIjSXNIUA5wtpN9tglJ8KrR3mZdLK
V6bTL56l+1p9tLACZJ/AZgXRBnUv8Hd9wKPSgJUGs/oud7I6sJu2zBAfVLsnWi6j9OKYfxABmccX
So6TxpSByq9C2L5CB2BSinsI+JABUNg8YpjdbPgmtrXmxWFg4htjIddvaI4Um8mpfkjaXOVATdVz
XuW4p9a8Roq/pmQKEJcdAyrIze6DZAsHA1BRt0xlWczCDrFV8+5IwJZ4SfR9kA72k3EQOKikTyE8
AV47G8NrnyNUaAGiE4fauDz3VrZKgKhm600hw3V7uG9frZ62gP6y1XaLllcbiD0ogXkIwCNZmCy2
5tHQf8Ti0J8WJmj6Mynea/b0oR/z8+J29GphkSAqqI3yPuiFPbC9eEVvbd65ckKsWi8ao5Mws3BS
6xTJKkeCSOwsw3WFZcdMEhjso9OcsnPyR8g87S1i3WU1Q9GWxM51dG0iQNmwQmD+Mj51hJEFrTIu
evJPZvAkQfwdAF1+6v8myBncxvEzBbOGpx63USXUarqskhwa7moEcsduztKMTSiYRtDqNa1fOBaG
B7E+bozo6KgYPh1H/UkctbZnh81LGN1QCwDus5mxmneBUUmigfSADSSeN5xfXSvaI+LRATjR06dJ
+XDVdzQugi6Hj1AJo7d/wJT6SjYDbcRwREgbhpa6DSPednchJ8Ej7srO3joxh4A9Ko2Rf+99AMve
otFqa39XYLdKI3Ndma3svx60a+EBIUJZcDXV6EUgzvvarPOMz/E3Mu4ugulLCDnZwxKIkqVDLUXi
A1G3Paf+RhmE9vRnRNXWsHlJlEZSqXHEXhhFezYzK602KD/S4KoZRsny5st3lyN71wf7K/3++jF0
gwjoU38wGMyShd57+ShDtlZzFWJV64FlAAOxvv1fPnhp44vcloWNJzgZ3yw+T+v5z3dIO12ZXVtA
PxOuBZX+9jYMMjRTqhI5Iusw3Zfd1vf9JcRr3JW9YPylFMcHPSmwKz7oZ4m6q5YJh7tCDgGghblQ
FTbbIQ3DSYgsXcWgCuEKGNbY1POmP793ZGoOePYlj1+spu1ApzjO2PYY8shkfZHETRSs8JVNcljx
FTdllx9DiRYecASNw4ScYTBobfvIkgdL/JvkwRUO+4Q6XRY31pfYp+5Xz9memBVKcRd4h3MWCDed
SQ/iViEMnAnTnCB/is92jzESXbfipC0mhyQznZGnFG0a81LVQ32GAqVhuW8ec+e5olbdJO0nmATI
QJpkqTdTLGcDfDUdHb6hJNm0f5gr3S4855VEt7or7/6tSP6RXBNpflH/SzserB3a+MVdOYo8ZDYH
Fzj2RhwurdYJfLUfnXB5/u6obioVGxyTD368+tM198yBiR5laAexjYBcna359v8uCYHfZ750TIs3
cJxY0ARzd9GvTgHQc7Zef3gaDwDqrmSQOoWb+EO7IpMmHinWKlHZZPA8DeEST00oot69Kbo47Joe
IsdjcaaJr1MN+Ub/81w+EiEBJjrZZzR7Qhw/iD4/4dGmjLW15J1mK1Tn6aoNNfLJK5OqksGYuVk8
sbj+wzug9N2T5QDuegKh2CYGd3wMZiHDkqZpF01+wSq+PViYR+dAaWUXsAroROaNI4Z4MBCAbrwQ
zModU/9+E/vRiL7p4i414Rr40vC+V0XaeNJePAdQXfv43ZH7a08MxNYhlMiUsGUl60rgEl02JeF7
93EBYDVKZZQdu8X0tSaqapceSXrw01lbB96rnqNHOxmvIMwZfqLLyCSVtNb53jnXIgrEn5Jeg7Hi
qHt6eXk8euJ++9rorcK6Ua3V4qhnXUzsm334gmcsrAYeoLWW4dalQib0hbm6oPCn/Aex+OjA5dHD
HbIpI11X0MV5yTa1ULuL2vrcadXws2TYa9qlEqbyqfMAgFLPXK1NNtCBnC7HYXhNa+8zFNaXEYH2
u0HwL3AZuLPTqnR07Z4sfqz1V1peVvCVQsFZMqpG9gahCg6TBmPkt+g/U0RfkRgYg9kkD1wwZiLP
I+UjYSax/M0DHvUI7Ih5cQUxqtvz66htxZIznxrN5vFyqUGyTSg5mDRuOJkAVr+xUGu7mQc7lzpd
gwjKYznzhp0x1JFuvgzKPjjm5FZC55read8CBEWLcsdlfA0HARtDOAUz0+nJmGlqP6llX5OTtYdw
b60DTvXv0E21zqGeZ20tB3IypCmX3gtvklvqXJaSN+sNzHjfxeMISe+Vnvs4ZuuvPNDHI7PZYs2k
b8TqWTtB3XLkS2bBNqibrHFgt1YQbn6efZCZIButPKgtMu3g/9SQLI/MPx0QK6flXxafK2m6fLYU
Jp+SCbs0aWvYnpsQp+Biw3k7j0qu1FaoOUr0+epjtwn/W/3VR9El88zgZ8faEay7tkw3QHkeP3L2
TV/QQuWQVQuq7U8SKTz28Atzlp4n38dsro73F9z6PbwKiunyheQUoCxRBlrTVdJrJRdvKAyPMsVg
DJXj12edhSGIblXMCmUC4J9uOUwx3i1U5lJP6cvoxzXumjgZszMrrEyZbmPrW/2DGxocFEkOjXlM
/PtymaOA7t3ho7thSmG3Ia9TzFoOYDdF2fPf2mgvm31+4jwR3DitQtYvPQGXrg307E7Vyiex7goQ
YD5M792PIQXrDDl5rHL3w82OZ3JapIxr4agfpwbfaSyzSfC3wuUk7XcLvvjagHe7AX/Wi+DJT108
J/wB2qL9JaO6I0lh+oc1nFkOXEvKA1kSyrMXHcqR0NIRrAaFxqNs5G0vZyr6cymz21bo0dTwNrjY
1FQ0Jq5xNkw3mSt3Am+ZvY/6hNy6Wpu0AfvjlR7GxCuth1hax+hNow0w9W2EjSGxp22Jsr8sB3yv
Fo/KS4jXfayC/6RQpfgRxffnlQLvZ2Ar3swLo20RhUJq+EVFW1XOhQxOr1vuNvf6Eax++8lkYfst
bZEDCLomrWsfI9SLfz4JEbcX/9VhWO3RbS/Og1VYEQgFgyx/RaC3HOnvrocKwCupAh+ZoXZ1i/BC
ABYxHk6wJCzfVFd35DOOF8f0wP9g8ibZtsucHkkKoRMcVcjmIZvNslhBaTYO6UAHWSJXbJJlpiIv
MwLKpOQw/8OBaoumqBhN5srGykuhCyRpjcyCUOxKawHyE7DBakFeL4C4mNYw/UZQTGARzD1dP2yD
1ezG7539fsOav2p/qQmQutkn9Clkj7jFSAt41FF2D521wV5fqy/WPwCb/NjU4yR++vqKWfonWv60
/2aRoqvz+azWVHi1xdAiqfl5zsBU4DUeCzZCqBFMia2YLA6E0SiaCBN5RcAqLY7E/a2CmEyvjgqi
hKOZcuREYz2gmu5cToxM5c4CVvLYFWZHipQh8waSRIXjh2IA2Iv6G0Q86qfO0Y/lxx9SFMVvTVPO
3Yp0PvPWHDVtv1shTIbNzhvvYc4mGOYEOd8NO3HyymTUQCOaz6OeHKEcSb6ZQ4VNJk5dRH69c8+7
uZYpD9N0eApQ3nQAmfYXSaw1cLcb2ftj8Mnu8qXV8048j6MYSKhZb6gkRRUumSLK05h8vESmyUnD
mzkv5ny1OPuSR7ooZPb/DUj2uLeE/YN2B3w+/RTIrcb4jyNXc+TCAdHgINFsHiziEgeLdFeqVta2
G4O2gs5JB2rwlGpKsBsMJKdT58Kw3CRQhy3AyZLnfIVlvv3lAm6wdRIzjJ29j/OLz6Qi5IOWn6JC
fOpr+WTBvh3ZH0fwcilhOcbQq2Zfhgo2wwBXqgnTwiu3A2xeStPy6/1EXUsHhQv9J1s8RKIKJ41H
vCesCmQ5D2gFotkJc0a5QByN5pec0M0S4/a+I5LSn9iTFnhLSvzdaqDO+Tysoh2miR9Q74tntoYK
rhgn3J+6HBNyDykc6UX8qtVc13yNlVsSeUhLpzonDhJCcodg4AMbreOaGCYBA7yyFRmQHgyR1L3b
P9CVF7ji3Z4hpdM1jx5agFD2Do4luYIC7eDzjt5wNb95BeXQTQRwSgCu0nH7JgXdo7VOxgj/L4Ie
yYOIqZIUCQ==
`pragma protect end_protected
