`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
rZRIM71CojWnh2+YhHA3Ibo7IcBWp3x6+XW1+0GSk4YcB9UIwjKZR0Vett+7Z4R31VUv3QqDYgOy
PVYduIo7y7o/UREOIaMeDigSfkygmRn3U2Jq9M6D/01e0Q0Ee2nQwEpEYgBpbTr0a6WxnDaB0YUg
AuTTNS2mVgviZLn9rLNkigEjWHtqJMdyfjzgOrylPurtKoPz7PNC6lwYwMrowsWs9owONfsf0nB6
dNIFizHMbipzAxGIltQmovqgQLUb+sNZw6VKtZdDRdBopAlfZI7TchYvIlBkLkAhGiJB3KQ9CQIA
Qx4Jd7rmhhf3a1wtn3Az6nqUJ8YLSRhwlb974g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="qKkmiaDm0UObDf3Nq4vhpMILlKKd6gpFCUH8FWN4ueA="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56304)
`pragma protect data_block
BYC1CN+VtqmfMzlnggKhea49A21J+44bxO5fzxNcM85eShYU+tHwvKVkenUtQYI235Eb7sBubEiX
NnpsFofZHpVCxgz8TUR5SGUkfjMhY8z5zhMmKoxNdETo0CIbBXo3aVlb9loTHTR0N0vj9Df0wBYM
BKw6VEk+5X6X7VeoPvqWZgqXlshHDLYqGC2/DbBd43FvlkeMzR6ZA+ue9X6aOU96BD+mfCP0/Ypk
18p/sf6XqnBUQHqDA6EE/c5CDXBLqq9u6ERXeI9c/+smmlkN22fUlLqcFcEhO0iJk2hvT7yHxkeQ
L3pR4VN+tD1A5/sgOE2NmdWXqZf3mn8FnUdFotqMkWSuCrhwKn97u/mmIMh4zGiblk3iix7MLTwz
ruRfuIqDd3cA/VQ6aQZE1NMHYftYsiF8z6ZqkpyiwJbu95xEQSZDDk74o4LSk0DIu7XkB1mFMGSl
58d3axOroM3Djb7Fhcr1tMKfiFcMAIA5RnPPMHozZa8rhN6Og1ddu/fFKp7+rzweL32Aowvs+HI+
YbJU99NvgRNCC/rWikm8DwnnzDVaXXTkYH0otTbphTtl8yMtnuVsM1ALDThEYkztgjIBWY/EGdbH
RpD/jUXYgTbhXKY7xQci9HadnAYRprxpB9V9QfW7Xd3s9vyKKqwVHgIDy9/UrMF3sEUI8aeBeYRC
yMakGeAoeyFTDKUpFqOT+ZEvZH1rMqbNplug90qk2K8g93jIVlcOIfheQtRnPTenHtBBn/zYEYPj
vu7bEAp1Ypfyuvc9ldnEgLb6y9dW0FoZVzSEr9cvy3JPcIO+sRkcajQVnMQxKjPBaLZIaR7/J7zs
kEF1+54ixDuIyNX+QBxUIanAUk7iqIQDed2hUG0kfoXoL3vuow/GsZ8M3G4iHfWrH7YjpZpxAU7u
+39ASljNjmhxyj7sp43zFjND7KB7yDk1EnS5RQNQKgSwY3fvRC0feceeFHyy9eiKM0+E3KW82xi5
RDh2XoenLekPW3PgKxqpPoG+gCC21CBlAB1jv2k6OVsb0sJjvmBbm0nN4wPphhhkwJPqYyPtdgZc
CE4B7f6+9YX7gFBCcgjzQVF2uUE8CawBOCPpR/Fwpn8AjQmRUi/jdffkvL+Mp7c2hiuOwOEy8CKO
/k3CrWI5eK3oZ9H4S0YVWsxKV2vSS81+g3WlUet5CAIguF+VS+SD5tY9WBAwxZQE7u6EQYtbM4nF
dSzrGuH9TqRgcRaYrqUXqK2n1/c6FSw5xSW6tedxEgIidnvmN9orDKJCvyomtkZF3iJEMaj06dd0
QvYKstibDHg+CT31ZlhQ0w+wVkvLRL6TqedtJ6VgNxaZ4pAxG8XkZpDZL4FAeJRgEL3+K0aDVlYX
T0fUHeRYb4FRGoE7CI5jD5zLk9gz1z/JOYSbkEVn2Eozb/X3igov2OHiOwxkjAmHhMGFiaPaG1bB
v6mOiGTeh06Rj1rs7iDfo32XtJ0OcZDXSQ2gMiaPiShXMREz5RsoPHEk6P8xdvF+weok88iEkhbw
WaenA8YisOhteAeUs6DG7smvKjJcTpnXsuN0I5ZlONwMsamvGF5RSzrd48tQfugGE9mKHGeWOHqA
bVP16DFTPjgMHF0Tts22AgE9SUPG5ti6ClVclzdbt33mRpW4/Vyl2eH2MYChl1Zghk6PjCyR80YF
Cuy7H0aDmyQHWXhH/j3/47vHsvOfSdUEwEiK+tlJ8LoDVplJb4LKl+oOBkjojIDm0TKZZuDRWd6l
46+aKRLZoKfXBVPln13lFmzp2KQFQLOWuLhvn1VODtij2DAOzJj9WkBphaV6DCKLzwu4vWLXHwsV
upWUqqUnRJqyXEA10MyGBQYZ6ntMVbpNFmzC7pbPvWrN7O2NXHYR69QYsAjhV21rANryfkhegq93
+8uN7thXEI2EeJmuIK8KlYoqpKFznocGmdrRWrZNxDZr6Hn+188+uZuXnMzOFaYw7cmWyzmioRl4
c/Er0SrlqmePM/AU5YHRgo2DWNRnBZ6p9gFKB5ITSbKprfqmiysz334+pzQfvqpZbmYd+SHZ9aTp
4ML8pvazY1cR++i7/J4fz5sq/zE8wXeAAQkv+G81q6vJrQdsCEzA5C+eOLVVgEgmqelAvaP8UdMm
cb5mwj0bTcSo99ynoTlPiawMVbhKKN1y4PW+d0T7fuAphYSXaWVoXMctw2ZScia9BXX0dcRsaQ97
Feld2F7fKgnexs/7qpcMx190WgYLZP0QVz08pDpTS7IK5XK8dhXZopdv72E0SgeuLRDezMe7gsOm
rsISdWR/rCgiBuERlZhl7TpmRw4TopFOBbe4A0mE03bQukc1ld7TWmAHhqR8Ia4P2HZUAy3ODLPC
Yk82Ts+015JZ9jIwkGtnCWAmeoZV7ZmPYHOsITGKAaM3npERr7zoVlXdtto2TciFk0A18Y4hYB66
9WEBoLuQf36pqc8Gr96GcUONndsWMoJ3IEbC9mQfq75DFekno8p8iO9qS7+kFUWUEE6eZ3SsMaOR
SciltY5MZZS/2g9J7fVTY+bTyAnyYeOBpTztweCJoZL8WddUnDQdtPaOYZkJDqZ08oLL7yJrQgWP
C7iFmTNTX6IadXVnXpTGkT7xK5lBQnfCq5TCcGf0apStQ9O2POnghE1sS56TYsvZiZyr5QIwrG9w
Xwafzv8QpLdp9HCN25CntkTWo1fhaapomO71FiHwhICecnli0emXaDvxRcz8YAYYCdzTFgS0p/NP
0os77ADfm2EaFOcgMyVx/aiEn4GbN/fgn6fmoOUed0k3yi3IKSVYB/uRG19Z6HuZP/juJ+SG88RG
G8HT23cgMhF5fiAakw20opvGfzji2lCtPYyZ2EJFA/N12ziPTLSXqyELjc1HMpbKN/AXGK9wkRhi
Spl7rtcTDbxYkUR3WtdyIWQ17fHUqyxFCBYk6kcmIAx6ZsGm6ZLEE5HSJPtzw2ZjxrrwW4ErwQKF
IbxrWLOi2/HjfH2YZ0MJ7Qt41mwEu9bT0O/MMixj1XAP+CA2xYF82zKBoAoJ7zs0Y72/LTXkG5P8
e9RZxjPLEz/mcvuwPtZdtj+AgYYAQ5MGgfizwJZDEQgDAVZ590t41KuvlZtFX+WW4k+5y5keHVeQ
g+atwy1zi4XZrYd7YxKCAWmjVuy8kg3irWYpTkr9BSsX17uePKyXiqgicV/yUPXCKPk7RFDRE4GP
Pm1rYnC9G7fTrBA/Msvb2uoPEzV5PlCkDOkYsK8/W5+GVcL4W+KZrA+mk2w42nIsc9oPXCDs4+UI
aD9eyHvxrHF4YmbWObCoOPP6eY/VTrnNBSjqvezELECosUC/wfnbbVB4Z/eZAF5wL6JshglzUp6R
wDB1rxQMtIoqQWvmradFlBQevdBH/bfyQ/ZfS3asB0LKHMArFbyk/YACCya+d1Vk6rb+U+OLc0EN
uMnmCkeH0tPsXtYQ10TkxdVp/sNBAuI0AUjA0SLV1bgaFncWgobjPn0yufObRPOD4zXtmOj931Vm
6e+hZtvYyAkMF1xZGgO576rdAMPWyeiLvsFlXcM2Gr/GlVyB9m7VZqSqAUNYQIDSVpTcl95eAE0S
Jx8aH/YlJIzxzih+M0CIjzPRkkXF2JkZ3E/5gQtQGQ6NU9tTE0tJ+fT+vrP4P+1IKYazbVMEYz8q
ChP9+xCe7EZdA8jFHp0fupiRJJkaWhkdBU5oFbHiyap7R1Ugk2Qdy2IMMeHQg5M/xoof/4vXsedv
CF8dLjjtcetRkRHP71uUZ1FbjVgKwy4ofeVSMSfffKi9gPg0hlKnTipd5tCIXqI5PbOYo1h8YnfN
r2mmDcXFKVPApab9z1ns8FpLben1hF3WsCP2h7vbSsYz20/HkYw3D229gFJ7azeD5Kyt8a/x/AL5
MqBlthDXNbR/7HTcd/qxzXBQzcvJ6Q7hlKrEa25Vzz7eeFHfgyO7R+olGTFYmhwFJnCK3HKoOuQb
bU4ABmUILScFRrtaMccNePXf9G9Ofn4T2wuNjoBM6tspCeOilTo1T2B/ETa7oTHb/VaTwE3GNLW3
EpKnOFbIdzWcgAv/0zDErDroCZcpYuzTpsFUkXmCuIYRWEgK/pxGTBXi7JaxjYdLk9D6h5PaTTSL
Fm+fAxUQrUTYCXfDSNQi/1+WluxW5QCuJx4lrCJLEaYr77DgTIrhMB4z43iO5kuH9WHrqkWx9GG/
z0p3j/3VIVj3Xhtfc6vs7Fj3ko4FjxR6pdYqvJqeqLonO7rr7nUz0tMZk1sR8myHHYEzJS8q6drX
SMb8J5DsjzQsD8HOpvFMe8hCReD6npuV2nM87pGJjTlYaIrNTNOl3A4DVGswYhPK/qem+Rg4Ynli
uRrKZ5B0ToEOBU916XAyq1kR/74pI/RfORw2MczwEyUaME1KAc+SYjEiUK0XBxXEj3BhjTobdR1Z
rZ+Df51MqxgsxyGGSEwiKiGz5Z4kBO5wr7DC/BC7I/zmkbu8v0bU7pTK9zo5dx4dHWc77zLz13xi
cdgiiPVGsqtYvuVIp7vdc2A1Xy0Vp+UR3Arg5cptmvo81KRtGvhZq1RRWxam5pJDo9bulE0fzRGY
ACkhOg0fT3g4d/6d8kWtZcWNu8o5cD6ZKXdZNQ2GgZPvLMoKj3AC/QM3mMOh/02si+07L2zgFgha
G6CTWRbGibfAuy1Qboy3CZ/Yett6rQYdSJ4JV0QZ3Bbd1WRUlPhspgD26vlXXTDqyfDMvauDAyzZ
mYxVzSKFYUOcNrCrXq/jTkmiOxjMGTw1l6cEFxjxiTCpiTfYZ/EXs9H0do7LlDZr/NuFpE2Vxdxb
niMR/KPnBs4zPPOZVtV9n5G+MQxIPpJN2InUUO5RYRpRZkdb60lNglzi6Ujq7e/ZGWzgMFcu/Qb/
ePhIijc090dGHa4mYr4rOAnSzTs1RsMy/zfcDc2NZb5JqUJO0+kPYR1/cX5/qL9CjkYEyLCeTy0P
QmTIROOY95YEaVXM5YZecjOcpJ3Gg6jKzRv2CGpL/f1TJeTUbLLunzorgsgvJGDE7LcvkHkjrgo/
a5IQEZfDRlt6gfTth7hvhzdaydTH6fmaL3rtVCA51Luu9dO1YxT4F1VcU/xr1GfNn4sTf87IL3Km
0Ewbia91RumhfnjcZSALFddliDsp3IQP08inQBKcvsXhfL6kf7bVoIieRJJu86WiRhKbu8/w5YX/
6uo95p/0XrCCNQP89pDcVUhYpmLSHZCERngah+46hDaTAT1BayWHIytVpT3M4MLZ8HBRpbIz/7qM
sWfIV1txjA0WIDqA5FqikdcXMeUofzC8nIQuh8LbPuxnz5H5hZOJidNsYQ+uKR+J8EGAM764YQqA
bnLXGFs1Mcos71JFGuzPIrjfhtjuftMcEK+6WEkkTGnJ0piHlALoNqoKH2YzeE/Kx6HkTzIVNsZ7
v9MzMZHTvP4DQZKtQkbi2e5MO22lbdF8CGQixFw8rhnYo13w8Hllqp+ytZ+4hnwkpOVofvXrujOE
KMofa2g+3uFDj57DKoT9plYLbqfmbkoWNH81YGSmzzhgE8ltE0+F6MRylAjsPgtluuL6gjds43lu
XUyj3rr8qtWBswguCDeBGcrSpJEF5nFfp6kDWE6ED8mJjvcYmgarHQgqgI8OZQa+2eZNOP1g+0U6
pE/f2Hr+KrUV5wHv4hXx6CnKYvwZMS+K7PG6kdQBLD/FWY09uOnhUjHp6CeHNx4WD4wgv7Q4fXBV
xrCfaRk8t2ffJsziOKY5B+I7tWOJXRPV9E9Q5Em0m5ufYXtW+RyRY0fCE8juOkWHuWH4GaJ1Y4+d
oHQoRfM9FlRjixV4PoA0hb2VgZc6hDi1oGIRfQ4WG51yfIwExwYvQolO0yG4ZCVyMAIXhUHbsFnF
0RwZRU+glkvuoe2PaeKJVBn+SRtWJxBvQ5H2NEqCvJfuhePlxvIm86geuVHrCBTLFpqfhPL7nAny
fZnqUgi9lT8BLun4qTFMsk3N2hnZouC8fUBACf5Eoe1AsYUsifozD/tTOPXXDoSYPTy2SjbSfP8S
wK/gD8bAIfLHWH8KljS1pXnpJKZQTi6zi3+2EQ+vQ4GZZKtc8P0Hj4B4hUDa9lcz39CzwxhY4AN0
iHy0gWUs9LD/sEasnI/TTTsfiDRV0QjwbkE2Bg4VdtJusqbLi3NUGfZ47kYsFnXevwlBssej6GFR
KxY3A/c4Vul6RVQ8iaahWlCpYn9kn6Mior1aHpwIejMmjRsiaQaQpjvGE43eBYW+6+1037x+UFP1
5PNnPEJ0JaRZWXuvzBVZfG8a3JWtovRAYpgbUVKoZgrYgZzCTzJZFuJMZMfvqTF1laCQH7wDLJC8
gu8THIJYe5GJ0YyyX8QXR8bda3UxlbQ2qp09e8ob7Jnibdg/oGJpgJXZe1hjRcVyqm8DVrvvvUcl
mV0J5WC+iFUqY95WW22JuTMY/3sT9A/INUJl5cuUDprzZ+QQ8DWZ8LrtMnxOle/pqma0WKlWFPR2
miW80R0Q22xqvAZJz+itE2p/QqdmTIfnXIyP+s/LDx0z2FeD7o1ntCxY6S36/rnxosVxWZWIYAOY
10fkOxjraWNXAOVZzpkcXyxTziu5pcGPYfiN9xGH1cdYRGUzquyxVt8INP2PY+TpIvWR3pG2iUGf
Hr0LKiL7UpUOc0F4p2st66758X2syR0wED6HhaPr6KFqn24mVfWmRcTocM/0ZbY4zvmD9NxswSJe
6FIqqy7VjKnJf3ew/SAd1gEDqVvUtP8NcP19kchUMJjST+RbmaBCU37B/WnallMlfnhz8o5PHW5r
tI+7VNLfm006pZM5EikXVy9TkJnUqqemz7O5RGBs3/qDNdgPWpx3a92UlfWOJMRAJA4EMv3EkxIi
UMo7Rr/HkpimiNqZMzQv30PEsYiyCLYbzPFKpVofASjZYnFclPzpxvifLOm+coeyZEXnQDsdda1r
D9Zg+lyssF1YHBz+akTGz0J7BkFNrQ5fGjb3piI3qqNR8sHWqCQRyesWD3fbHkj3ViUjmSx4CQXv
S2eNjiK56zIABA9u93tLRe5ax1cK21bbPlANHj0Dej6uDC2TOTY/d+kw0huTBN2I591vxVt9jVg9
0i6i5KcD1ekVDM/h8W/jdeGUaW3Xln7s8WiciGfYPNU/GJbk0+pnKe2aJlfXw8RcBEp34r2IuJN0
qjGoLrM2RzE/Dp1h2oZuJHUa41YdVEP3t6PX6eNkxETXOGXquE1zHRKEam9IUPdbfaufhv+ueZ9V
JygiqrfsTsvAZ93u7X1qOy7tsoKCPToHaK22UDJ71WLPkF+W8W6V0hyhIFV4mPkbNHO2R/PhEhvC
OyGFzW8tL3MLoMP2ezrcdDIs8SCcVOtBcIw42RWuInYZDzGgCJtcfeXbA4nrFwJIEYozKHQtWynf
2Orkqvz27qRXl14DnJPZOyfwZE9XzQsy/yIkSEPz9VD7K5mVCh8di+h3VHPCZglwcIXnM9EvhUta
ijVNaekZhTN5kDsiQ5tH+oHlcvQK9HmLZtfICmGWBEW+8e7axh9nWtd0FsjA6Abh75YFU/MEQxki
VfEacajfGhCUfA7GmSoTIetWjN0wQ4Y2WER8WGSWTUfqwtYHqE3a5QyUjS71MXpQ4mKB+19WffgP
35ZZ22Vmm6QiJf7nLWBG1H3FQfKdcBu7L58q/7t6U0IgERRMwlUGms+SP+b0NwslwC4x/NsE8d7I
3/jQrIpO/GOOL6KHftvHu2qs+yxP+Q12bWwYLTWg5eu6bSAOsc6b3G0wp1/U6NCbFZvM8WiPA2Pt
/txTkkRNYDpagOIsGRFXbnNKxR+oaokY4VuR+rFcYp1ufPeBwmJXVu3d7GC7hnLbCiemh+JtSCqe
vgkh4fdsgg4Oh6wbpgGcTcqlFnjw7/d0HKGgCNFlZyIwUxpXv1neowNWyFWJVKXsYqo+/tsQRXUU
z5IoENuCms9mSzD7fgTtSPOdG2WUJxreC/4CeAHLcM6JPjxqOL7m+70miEp5scHC8UL7J0amZTBN
eEjdKFrCBpWvuUh10Tz3qWB4GBnmjDkAzcpZPmlFPJ7oh4lXUnHEOSZZhK7nN5Z3JlpSyzvCqJzo
xrKJutXRjumQz042j3jVFaFtyD/MpvDD4FtPeR2Sb3YpDWNlqFlypAGMVI7BGyAGmqhs4hk7no6a
VSZaC2g0lZR8JDwvh/RA2iyQk6u6uYPIXEwLJXBDrisDSBwDr0kgs1Iva5PLzXeWs+Yj63CFnpOU
qHz2KAQRl3zuQ8jztjaVFjt8QRkWFVxILcikvm+IOSDc09x50qiqXBe+aM7nXA85UbvbCv5HrQp8
vpQkuDKx3q5/Zx6UFxWCMNG6KMLg6bfSAk76LIEhMiKY8agiXf1+NaFSAKPSzBgEQJQmJL1ChsPc
7ovGfyEVUor5ioaQLS3q8TA4e3TKUKshmooYd9pnEFPFOL7zvQdtdDD6mwhbl4I/O+VfE092Ic4J
u/i/eX5cdVzqPjwCTS/LT60TjRHogbxXoQEki5p1MmVq79ZZo0+PIdDP1Xv/+bT7vd/iceXUpFK1
3U28k8935sOzAdHWF762AgZSYOXVYhac09ExpJOQxW9RoHugpd4+dRIN+JJVtmaX2oL49dfPQoYu
SiYc0GFwUrSbugvXnJfWIC8sB3UawkoMCJAkEZ5FmPmeW5SspA1WFAL9GCkpenTfJIDPC/XciGUa
2PSOmp0VF/v3HEACnQx51HnIgMuWNbm/1E18our6I3GQs9Du9bpJDX5y4HzEDbqbE3dk4anAXzMc
2rD70Hp0+73F8sa6WHkcGwFALZnhnHR6FuynEP5vXIB9xjIgyenZ0XTq9Cz2qqg6DQXVKjmgypTv
u7WbeIqox/amMUZdKzs8Q6cQiB+0MHvLJ2dN3Cho9fnWZAWj9hVy6tJ4Y0IshbbE1M0rH+E5tssQ
lBGL3I9HyVPbqJUAHaxMMLKBMhCVwUU4Sq8UX53d1YFMVsxgjeiJoaAKGAeIy+/W8hjh6/k9T17c
LagZreMeuAQ88DJmcN6bfkaqGmjXCD74wmfSDxELvGoM/uov20UuF4boRl/WavPSbUn7KYzwRxPm
gst5rXKhhJmvZ2B4WDk7Sv02sIDWbrM7KWQYVTlZq9HeggFpmzDLWBgS7Ce0Ub1s3THdYIv5gvmj
iAYcQV3dUcSIlHuM81/DwlhSBHasSFi/govWjUYwxo/tlShrN6F/8Pj3VsYRG12NxCupahbDsMEP
r1td084ubAcPEbKpsUSw306w+Q6GB8AywKyQhxoHWAssut+AsRKq1oRlxCY29ef6gQlxjZehzpGe
eiTmJN+mV/PCvnRIBeY/0ZvjjOUilgV2VVOLO1BreCMCTNAIaM3LKWhGm/nAVsHIWSYsaOE97KdT
1+yewDiNUWEUCHdMxPINRsVDZC5Q3aGc2YUPTQNHTLjP4ZHEbPFTpKl5TsM82WkQUwdJvrr8MQe0
5rg6DzvPFSE2JUErMQbkySdC3i7n1JDEzLt84MQy+0Mgf6YcuijCb92PK45c+9d+qida1Zg9ZuV0
W6svkkPSnWKgefi6oUrluCWD3gowl4AKmhn13RRB1Rv+CUcyJMA7ZTblqH/rXUoYY9G6vHVy03BU
MGgpoFmR/T49mbQ2dc8CDPOVK6hQaF47my8BM8UeaxSk+DiEd3PjQelVkBJ1iTOhTe+Af9swHpEI
fw6O0PjxIWsUSN2c1leoIq56PrUsCj7/7wJKNGxXJuiO9SamKGJsPSY6MMieqRifD3376bOz98kM
CDqgNvQtsE55a6xi2QTqBlZWnnXLR7rsOpNugyXucAm2oHAnXMqsxgu25FGPHNlDodCw0kC7cQKV
ZMV45QvbdwSzhHDC5gBoOo9OW2vOIsKbNKGfKYjjZJZJ+S2uEe5W9H32a7ye47rvbE44ZV/8SjeN
/bifg+8cofR4K608/1CmiguZh8y27J4pY2uy2roG1KzhmA8tYlBNjvFxNNRNdGCQ5z1iYdu7VQVh
uARUmJJpNF11ZEiWokPI9bbvZCZBtgs3/lMyZMud1Xsl61Do46pJnDN4mtKrkC6ZKfoIQ0eRvq3T
zhQ4faWmgFtfA/KPX/KlEynjo3A+wuNZQAQyR8Z7zl0e9ZJdtQ1wOW6gp4OtnDqUeeltYT+KypE2
deMrq3C4WD6op3WSOp1eE2wB+Y5sv74YUn24geDvDAUW7yawufx/VfmT8Q3FPKfTiLAG6+5o+vzb
IM1651ACP+hn7T959yYR5OMRBWBdJUNUS4Dw+Hgwnr4VdniGEfS31PdMnxAklqk/scfeFRca3L7X
ba6GKJ/z1uzXs4gCWYnQSYfjNiwCmkpOLH4qfEBjXD12pLNLfg0ORh8jLiyaBgi7SziK1zWPu5BR
CGKxImQfiemVG5+hSD3S0mwyjbxrBTwE/eknQWBuL8PAkmhLzL6C8IXla79slAbxdNa32Qxnu/cA
xrnropvmZErsD57jdy5oWdK3ofglL03cz1Sv/HBobmryGhV+4VpGPEl1FsM5gBaQOrsvi6OUi29x
ASYlLaVVpb2H0UULbZBFqzrEiS3ZtVMHaPktq0d4FtCi85N1U3/e2HUwSiQ1zdlYtYrXSTPuLc1x
vfSlvv9ROnnSBkmO1qzCCo9vIXpkdYq8rXgomDRyArvBo7E6Nlj2AQf2Lt2jgSE5Bn9HzAgndC7a
S/9GTaLRsTklz/C+JBSpHPFUEnpTy/8tx89nMZO+fWHY6fMIjD3QyOqL9Cg6SazsSWh5xa6ajgT7
Lt2hIrRt1zV+F7OYAb4BLNabADtWmaeNIlmKC2jIk4GX0z+Q19TICHI+krwAgX5lYyjXNdkI6/vX
BAw2Bt2gkk9w1UT04q+WX/ybFfE3/SCDAVdmlAS5gU39HmgaPcYz9vw0cXpo7ff3S+KtVe6oayn/
0pOfqS/jvjWnqb6vyJDLHrC5fDL6GeAlQqytN/xWssVjPuf/Y1A0+BNNlN2u+6BmSD9tfPShIB9g
+LvmrqecbypDftymOPfnNdi4h+CXeqW5foyS1O7lh52QeJCtQS5IRdrjXn0e8cAcBaAQc/HpgCsL
TiscckCQOcgqQmoAJSIFGpS7vAVwNzOySgOk6rKVWKTHnoXBMJir2Ri4JLJZn/pYFfcZlbkTNsnu
fSyGSr6gA6oPA673CjewOZoEABdtUyrtqyaYUak4LHQgloL8Uohm9PbEpCPK6A6Q1m1PPYcFIgEM
OfYPa0Cpy0T5nYtOabT+iBZu9kKwl3rZl17f2ONgkSUTomwlh8z4hJEBZDpGTrU6LWMexjuSEGVx
03HL0HP96czUGpGmWJX+itMq3y2dxBqX2N0+VBaEENpPq/KfBa/wejtbTAMBqi+qxE4dxMszFKNG
ymZgBSLjLqIy5+G7m4S2cPNE/ni6NC85Rv4oV1JcGVIixRpHmExr8X9g7iBVjLxK1q4XN77js2wv
wPcnQ8/AUrl9LmF+u+erVm34mqT1mxwo6YXTb5h7RE96P57qBG/Ikh840wMCUpHIFw6rcXt/Gvow
vLqj2WNMUrqJ6gRN1DrwcFdy6D6wqECYeTGHU1Pn12ckp7AjlA4THkSwZO05DXwiAybD0pXIhLRP
ek3cuIKTfRdN8LdR11rn8133+I3ZjEoQ3eJX50hiPjYaoitzx3r50HjKQToe6fuTRFqBNQwCr0z5
+WD3oNSFWd8JxlcnYc5QZk0gXb7Omuao8KmspZNzvRbLE3GsF4VmrJjCiY2TRts3S0yFJfuund9r
g02X1oEVqrq/3M7X5/q+sWXEvQULlkwmJ2nS2Yyf49kFGOPah1jTXNJpr91VHDV4gKyKMceaXMBN
aRTtBej7dE3oieg4tsb5+CsWrKp84dK99Z1bbepD0hWBFzbFOTDTGGSppSty5nFi3+QM2FCErV1a
2TufK3GMK9QoX3axBMYZCuGOH8DnsXnsznfuys/+b43YBexrafP2R7UfVutHAwwxbapY++5eOVJ5
rkWOmTnr5UJOobS3NvG999iGbXonv0COpTKttDPmbiu3DW8rvOnkVtj1eyeqxW32KJtJAH+kqHs8
zE72eh933UxZZ7uxo+nlEOGGuFMZRa6UnkFihxLd9jGRo1BbPGGLHcQbukKMVO6lkEtySVObOcR2
7Aa2gFDW0VjPI/2+SyZUIm9uHk6esA6ydrop5EbVxMNpC840JIBz1iM/9LLDp++v1RBWqMQuatJ0
leZYljDI0SIedphKIz3U283+DX+iMHroUuaJJEQph2dCc9K+fj5OIl6Xiqf00VsWerRldKUAhGBG
ObwoT4IKg1vjQTZbM5Ve2ml/p2q/E96vcIgtwH45NbApwOSVrzgEsNAZhDpmjD/Aa7ayHxnXWyfP
UgYlpsu0xhqpnSHyptRzAQEm92l42hoTkSe9Qhce4vs5HgzN1xJLq2Sw9gRJ3uLbna+9tyKdACUb
0c70qRwUNPP5BOZQ7flScB0F2TraVxRjFNhBfvdbOwGlwOaSNT/DfMi5lPvUtBdeKMMPXqCKGAH9
VG45gnpyEsDMlYUff0Wcdo5B4rJXYscoQLMZnOxx+bbboPIk2sI5/tC9MKNNo3MWTYku+Wcjg6D2
ZunuQicyiYoSI2jXuJUmI5jHflOw+nU/4HnFVF9Atmh5bPkhAAbp4lDGBLflFMsCcnIHwHzgGSOn
bkgW99j1h1MrJ+eUiO845Tjr0iIGHXkvOnFA6HQCejz7epExqmC6TVcF8a9VqriqDC9yvhCIAA04
igU/TIx2LIDwtQNbJ6cREQSPmOU88kCXhzrtUC8AqPUcY05dMmiXJn3BVHx+mJIb0+7BLia3tumY
gyM9+TZt7uqGR/ktpUPH1teOYMYOVjNmnQY1IVxV2aB86plHfLtxbXHKJyLFi84xwTsHnHmRWP5P
a8u+ciEVBjdtwcbtJ1xu2NQ41IJmIPxF0bc2f+WovUzeixHCfaQn/OpabrJU3lVWrGAf85RpIfyv
xPesS5CGg5kWxiO8SoLzCFdXKuSHzkM4xOjF5rrKByvXJykbZB6x4Rd+JeSZI2WkGog4++e3c+XO
8Prruyq64f4Yfi1ixJOkYaeHt0zWeWYhcz+arMiXyJV1k+luCKrq3SkvBNQ7mvz1gdkgu1r+MNCr
37fkJs32OsBy0d1yC1j2HI9EulmnznFWFcC52bHz85+PJ+U9Tgl2QXmllk7IwWDn3/RI9YTB804+
GGBA0ZfdBZKv0+ii35RKEponqKR/rosoQzcNN4PMZTN7s0HWgzpjnLgiQWRKPN3kUgwPvcABNKnP
26mpeO2rD3ZENOP81DCtzbwehFWhhAocJdBh5NK7hN90Wgrhv4j4zTmm24320mrcKAREpwPfqegX
fjdn1h2lStu1fJShyUmzg+7IJ0fox0yFGepuK+33mrcLGRJxSsO7h1hPdORIRtzkbY5mgEid/sAB
iubhplAUVRFqWfjXoCoHr4sLUaTYayoA1vnInJ/IVmjAA+Q8g87FliE9nyi1s1QozDlKQ+WyBMHR
RnNGxc2qwim9FwvXNniwfCAq0B8GveJwobB5b9YR/h64lFfuy6ZOctYhr3d93cZidp0AzdcyCIZZ
VjefTzitXKA1GwItWLrdGMBnHJ3nGyy3A/sBGVz17RAU88JN4lD46ruQ1CrTcw2cIxoydj6kJ7IC
bmIegS1z71j8FojjWtSuafeygR44vaBf5R/A7VUrHxlkP+l4IewwavrSVF90qC7m2EVFTGwp5ff0
fQVSkVkltCEoZgJvGzJ+6zEJk2r7+7RZshXHWMNKIYNFQASNQBX/n0RiPYxbayCXd5kRwm9axohw
/6/xKUYM9ZcHtGQdEqnn0P+ggxoAmiUwuumcwtY6LndMgFEyI+/RYDKc/VFD8bABPjOYQ7K7z3ee
29p3kTY7gXKemwZ5OIZvzBCOfQ/oeMN2bxP/+69rK705snlvHPgbUuPoOE4ltvpjlV62omXrNls/
3vYi3e+Cl8xuvXbtK7mdXzJ3zjTvekC6UiGbvoqy2ubqKr97tb6iwiAOpKA9HOictK87k1FOZsMP
oKUYKhXdh4yCj68Zo+nJK1Yz3xQ3kVqtQT4SVrqYD/Xq5i0RyMlxTYnIub68aFVBImG4blr1Trsa
GOOxMVQcnzAlKP8qt+KK9V/xqrGvPdnH8POJJ93y5n+xmc920u45wDcm9d3dJA/NHO+uuYViGUTF
BTAAlSOOZSkAEgJIqDePixdE42JeP1SW515OKikYcFyvvklkBfPDjnsU59GrTBxkflK8UlL2Z9CE
cPxIYCgvg63N3ZqkgzlfSxPaislakRHA4JEhH7NwOOZFdWJOVEHbnoLNSHtXrFHm+IETqU+xScw0
hrVoNBGge0UQ8whh5oKylW7rmxcwoALWqjr8aUI7w1tmmmIvM3JZJ9s2ZWp+oGTdyEKs/XpwQxW1
mqyUxsPtTBYTFT2J6APwP9HOK8GIkaxSqidzuF8StYlcmYzPmB2zmbJrVxYgfv51WeJFzB58hXeG
1D7I0GAogLKRefOjCV9axkldndf97lDOHkEJKz1orjav1ERoaqQF6OnLQffYBJ9t/qEfHpN0F5jT
rV9kTnq58XX1QX1gL0yG2R1Pvy/fINtlEqc9fbR0vltSGd7DopmPOgq9rbsdsQt09cI/HCB/7cYw
AKecNr+eLZLdAunPIAPpN/L+Koz6wATH7sHyXvk4ANID2UoR1dfhP1+NrNISwbggFc0GyX2hY8l2
HkfHnaaxszTtOS6e5cr2nCQk3FMxYyBBQsz2ub4/EVg9v9RMciMebUvFFxv3Z2h6DfA1zXkj7hiP
Q4Nc4clPf3t3W7EhqDqSGN1CXCfjAOT1lPEjQET6lJkGazooic7X0j2VlDSev08nZSxcHQhcdlFl
bKdNZ+HIrzPcGx6pKbBGZts8CHFkiFPcTaLU3z0EAup+5xK6aleM2tMWy022MmfcAIGngq+C8Jnz
gQPUDmeE7Ed14ew7HLLtNdyydPK0MQDSrHEmi4W/d9zip0ksAQORy2c6460hjxePI9aPF+mrhxi9
0u+po56T6nNxER/b0eEVqpul4tJtpUz7rLdtpbXqWWs/LulfFgSKGR8Q2cb5vDgci9LbdFuaGa5L
bBdRslHC3kMT7Evq99qrMLreeur4UfqvcT8ISET38dxY0pyf+wgOJqEKXHgljpTdCSpPmoNrykxD
4zqfzi9eKZemZaqphwPoKr82OZPwbj0xn5UKl4YJqXkYuu+1rRZ3q/76fqZ+8rTgb0sYfggR+/51
09NM8n+9nYYx5Bi4ejvTsAtSnrcigPmYnTowud/65rdV7mkrDkjTgZGA60gVfUQYycj+rEwpJJu+
XqOl23K6t7n5u60ojI6UBFf3CNHvXc2RIS7tcVbghTB4qIjnsA8PRRcNIoRaUxrG2ktuBAE/jTCQ
ZUgm2SBChGAEpz8xrFXx4lI7yzYWkRoV/FhlbyIItmsVzkV7s9agoYkhwls2oVe1s3XmEBgvDu0A
Q+2gRnBceO57jR9aeZbXIf6kKHEbPuGvtl9JWUO6fwLC/7/c7VrE5HP2Osgeq6X5M7rhwt5SjMdb
NP8jA+uGt2+qyi2/fGgTMqCxCK+IqIuygtLUflyBAxKpzkbb2HsHmPGEI+VDiflDns6alCPkQn9l
ULWE5KPoFTloToV/8SnfzC9BxR7JuFrjjUOGsmCZhM8KtVNKHghZwWT7bYljlGaicAZddT+KzrfC
tJv8QKYmlPJRfxcy+8iH4ky1UYrLXCeMUy1ahrjpjgvnsFyh8tLgYCL1fk4+TytCBNXGnUWddbDf
PjS0G70mOf9EPDX+BRSVLI6eCArYZbqxiUyeet37srAZJjGJpwaxrcabm4t1QcVDkUn0iviBTKZB
kFRsANH7WoMx0moytKL46OyvASWZ18+gdGC+bbPzEv0y/xud81ZtFlcNUHtARV7REiWsTDEk0RQQ
+CBmFwJzzvJqB7M/OWIrIn7ZCAZXp/riYi1HDKhTkeG7RJZB6UoVtdY4nF0jCS/8Lly26pV7MZN8
bNVTJNnRGvXN8e1NcEIOb8txCKd9MRdEuUXGBQB/Rq21PRIyKtI3XxNB6GpD99DTJsU1Z78ARVW9
eC54dqsxuxIMa/p6/Blhu71MDbMOkXaDPN8mYdfk7tjIEJqZ7b5IcLcaUmh+DYyaOz4llDzo2FgG
deG7DUcypU6cY977jp81bDUkxNwCQ9uPQaQzT7kSyDACwcvFt3uaLOM2C1y01RHGcygquO4RfUe8
XqvJEr2kRZm28df3loHSEOxa1mj62M2Z8pMzCY7Br3NSqXzBLUbWwc36GaWNQRgvYw0FqmzSu7Xa
m6iiZRLSbw84/qziZeh9jTAbU6Sq6aHiFStk7BlVX7xJQF/MTpilX6TTogf09oGtCeDRnCPyuIBF
Os/66RTrKXS6DS5/0Sy5N6ESQMHoya1Qdnp3e3xEwAEoTDh3ETLTTk+izIopJ4WhEatK6AfgfpvT
fFWBohOKzBUH3XQLMcUYBavOUsU65WxpzQqMwZSOL3Z0RiMeVDQGTouVQ6CpddThJolex6faCfjv
YihS+Y0SnV6TPrbRFTZM6G4skyrrPIhfg6UkDwCMmx9ckm2qGF3ot8KiG33Q+rPAOx3mO1ZT/vak
A+2iYQtyOjYDG3+sCYra0lgaXvMW/cQg2QSC6LBS72mQ4TSD2E774X+m2HD/dNavQ4ncwpm0hu/J
W/Jvs5eXxQRvCV3kpNdJ1JfATdOwKjyDuqbQkAX6spbC/tTVq+gyGTctMQ/N2x9S79nYqlwcoxPS
j/vGPcs6e9y+ZZl4dToMubteTfEHIKDPt1twjpH0jhnVA1d91gNBm+cOOnwy++KGGeSH2GUtVFfz
e25ArSKL8RQPvUTiFDwEzmcyNBMcjk4/vN/mnqsHCoZUesWf7WdukANCt9tnUYxi9YQTtHGyc1bP
gf+8GCzaFL+9zn0cj4n9Kf5adctB9Zjd1WkYzLk0Xa7TuyYEIrBtFA0yQPhx1p/Jd86jO68emtSk
ZRXJO9991MCpsZq0oD5GEZtON/QoLW5ix+vZsu3WEywwnWHF7PUatsltSrf3GcsSZtAnaqHVKlV2
WvWl0ON7f/APDH4HCKORozp/m8vXP9mTWoi2zj4QGb3iOHvHblPFf+Y6HppdooEoPk30K63VCKll
ttrrBqVG66kBYde5ZHby6BjTJ2/xHSBZTl6UNJz/3q5w+gDBEzHXcGQd07tpHfZ5cLLEnHF1FM+l
G3A+Q/4dk0HJdrziPxfrbKgS9LirLUec1GRlSGOzXm0AEN/ZoblFs843cGpl8OMnoVqBm0bq+7s9
1dPHR/Z7fzYJyVgy9YcdlVYNx2vV202zPdZxFypv+Nm+Vdyulpt3XXUE7vWb6lH06JSCbxntjhq+
PEV0a2ILJkBABEtxLJguq1VQucozogNMkze159FuG0NK6Zuld7zU5dFrDzf/8RXODzmbeZfzjQpC
ZFiJ9vooqJa2I5BSEW5fcVMyd2WMjo1j4kHu8npxdDmyINKvPsMvy2Hp0+4pD8PZS0EmW4nB0TnB
ztlLT84m66WWDxBw8lAO8KwRAe8YCfvH9Eu7cJ9MjFQ6TYCfcSDKqxOam3GCiymez39lCYQv7zuK
vtJOCBRcGhIZ6M0s9BcSzQuraJsL3VOs6MCjt93qKZ7RyRzQmV08hwoKGJDzRKgO7ipLzrLifqiT
H4LPPevUY1myyxGEm2I8jpmi3BN69yPA9QbUe2G5/BDfOMMzaYai433b/sYy/dGyblfVm+qrfil5
0cCrfHP82QU99enY60t8d9eXvsbDDNjwIb29pAM516QRSiM2VFF+0kolypcQNr34r5VueEe4wuQY
Be1lxCDGCSaRI0pi4bQOHdi5qif5jzPKGgpv9CdxtrU7wPY1rhfu4zoU9oxFMkwxop7c3FRGn0bo
nuX/D7qqN5KG7jImLhnhk57/nGGuCLFiXKZZPF97KUh8ejPeDl3JSjgTMFKBfVwFWQx4ZRPAf8HH
yW/eNDe5WrG0MVcJfnlQ6vbAklXjEMyJv1/rutFKToF5f0anvr5rt/4NhwhYfpjLQnuceQpioBFD
9S3UOdXcb4qRnFXWfxYQJ4MzhjBMkA0aouPmxcy/UUGLL89rIp2ABMctxX4Qen9ni8IY4xz7ToWx
SU2Xvk+gFize1/1h83+b5HpEJ6NrqICo541O4rZwhvwqIlj83ZnlnZQ5QPWA7W6+jeFkA/txLwTZ
YSbHtzWprM57Ray2Y68h919nf6Jsyho+bfmIOx60F6zfq4WbDQPoGh/7USIMna2MmLnXYU9pErDH
B2BRGyurpIpy1OPmna0p92maKo2gP1zeqBKPW9A6u4wxod3PnQy83fpNB3+vlnH10FBXHZjzhX3d
VkcA1qHc8cdmAWEpRFcjBCpmhBt0VZsIZl0+46TQF3BeqeqysS4KAkAK7vEuTtMeenBwd2/y53Rx
k2X9EzHUP598+0k2VSMZpxYXUruxqmOq0Z035il9zh7fohukNhvBQc2wKN2pGh96yQbVqk0Kl3vO
c9TXT0RMSiH4ta761CyxSXojClxJb8SJfkiUtkF4fdI+GJOwQpN4JjQtl8dQzHaX+mhXHCKzeDlk
aub3Qt9D87aVt3mcgh7C496UyphEvny908N4UfqdRczwoW/OcG0XQGson9jVdru2dZ6USEOHyF8R
JkUJxvFwAMwxO3V3CGKl1lX2UlwXuijoKuJ9EDNEP3sosSrFDwbDQoGnCnSbYykKcsCLsUQ7CRkP
OZGy3pf+r6JJIsCTGcdiuByoa1ReqylAs4VVooaPLT7psuuVzVAIKHDXDOmYlpQuNCuOmAJDe82J
Gpcm2IaY2n9YvKW+HyQGsuY4Qh38mmiB+V8aDH3coZugwJms0b0qtQePPw3LLOZ34WkPwWBF+Go3
gdrxbjXqDBf/HHsZPPgHFpPHGAuIao3nR9HozPgk8EFVm8PwlEZsgokfHfTSv6Xuy4SRcAKEIAxU
9dP9V8euyf8h9VH/SdnDVnKZfn70yw0rxoeBwJOoO1oi+2UdOSa5PD9+jzF951i6+CE8sTc03xQ8
0zG16bYf0hWsUKwc6NIRhrFuF9XwOrwjZUue5MQgI4LH4pG3kr8I+KJMk6zIeQ3Jw+5n3X2joeyO
dJgWbQI1IjovdjXbLsZ7V0nwr2LkXjg2Ibf/z4Cey9UeL3j+X11TXJ2fjqYpPvAvdq3Vmhdlr6Sm
6JstsgvgeUZ/YoseKhKciSaCcyaLCHZwJaWHhHul89ApI8YoIIXU2/SwBGW2+YHwv3Lb9g8Jq/lT
85UsHBokilQRVDkVO7Kt9QDsq59FtERanlFVoD+6RarknCXCm3CSL1y0qxIwfzPRioGVSkspDsLp
XlN0bTVVa/yU4ZliKccXNoK1GsV1a+zXTGlmJwTckpLVfDpkYw+LvyWxT3E+YD5vlPdiNlis9uVP
QsjOqPfvxWikg17WwxO9rZsLj8kJ+6aG3JHC4rCkpdgiSAe41h65Q4HrCHNhIXqJj5qebjrCSqdQ
Pn1oZy/hFDdAoyMJOh7+Vr0fc+f1a9ZmqlVF9039M9FgzaFVSjU5FbbhRkMnkE/kIZb8Fl105vU9
Ef1wBKraoZ6uby4UpBKQwnXRsjnkSkj05Dn8H7radXDDKCetD8MHVKBmAFbsuZP7uCdJfmTHeYm4
EkGpPghSyUmTOIDJ0IvD+2Ek5ZBBjyLiKkeu9yR2jWuFqks2pGf65UdvkjI0mC61FVZst8guf/gv
0B+Knj7JyZ4o/+uKYIW9zjNhll9DpVYsCqK8T+eqk73dxEwpixw2mZXBrTndCl4pL/VUG68X7cWB
jOjxpGLAV6Bk37KCLQ/I46zYg8w5hV7oPjnbRrcmh161uMxOZu6yUfYPecC3ZhwMXSTuHEaDCzIS
3+WQMEBnOWw1vGLoUhbnAJIFjz6CmXQaoGRyl8BpDqt2tv3IkWPl2zyMlCeDw4gViHGHY8N6+0oo
CZROwlM1lo3RgYF7KxQhx7qV92biSUq70aAxfftrhbbMGljvf0jftefUp2SniaYlqf7XzAqJDjoT
RZnxofV6DzBi6L72EKM34SfP1vG4vV7WWD/VucQ+uKBlLb99ZTQXULOpoXx1lrnusINGwQrDd9nx
0EGL+4tZZTLF/7yoNXykVlTD0WODdqGhykEQX3h7oEmUwxMmHs/GFMciogXIaVBuhBIecbnjiSwG
uguMUBrgzjH97KOpcqfEq/inE10uVuUOhMNC+TCzTvYQf7HVpupfWCCBYzlOXAN0DFDkmKQvrj/Y
MQ9lP8xzQRgwdIiBNHFZBH5vWpA/kKFuUe9je+q9kG6tk1w0b2uhIIiwpcRzwisLzZR7nmA0bDMS
2E5LM9ZpmT8jHSalnxZBqMij4GbrTExcA5En91OkyIttAQq2cZGupdpyTN6D9tYIEpZINlrjOirI
PAo+1hyULSKIQb0lqsQ4Ajq/OU1/qE9nscdhZf4fY07qe2LNcw8EVLG23OEbJ7xkX9vsJ6WpLDyz
uUsVq5Vd4Z03+2ZQaX7b4RzND3y/CDnrVnBgT+RoFODZGbPQO80YTvXG83C2cwve9xvWepxLkdpF
TR+/wqWmP+YJ8xsGohZuqcd3NgQq5y4thHEWWKoCNpXh/Iw4VnoXVviB8X1CxtPn3tjlD40k1oI6
gGLxnPKJ3+u9vGuRtxRxoV2B/PYM3LdyaQUOfEIJ38i35vWretV7awuJarWtwjQKFa0f6wERuKCa
frh4s+vBsjbTEBTWpCK6bmUmmZOL6bS5zYvFlahVDfljYIpHx67l+B374rJ4hX2DqPw3ab/hfNJw
qq4/dqUZRh3W9Ne3Wa6gWtQzoErBap8BmOpJ8b9NZXxLozkhNIf5ugXMrbDHVx6X7a0gSIrWEe/T
zDylmuxSjtjSHdQiWxo6kAJuVHdLQhEB/UJYO59pF/VVKWOpIw/oKt3P3762BYp2vo15j8RX+n9t
dTGst75TEmjrjkoUb3z7OTSnBY5zQ2VClB05SWmCFuAzPiaXE52HirUUxGctOh2qAleJA7aM/rK2
B0qTiOfKuboONUPGipK9yOCuABtg6y6i2yRbKV4umKi4hewfosWC8qiWzuxlDLJhEhRbE0TWNZ36
O4a3KgNJAzS+MBrytRSrXbXc2s5q/2j5x4Rb5Izv4AF0Xl8bHP8c4FPm6WAuwLxyvR6cy5jfj91J
wFrmI5Da2nZTy1f8kSrlShB6W+kaBAu/sdTqhalqqQP7dedLLcrg57zQ5u+lPWOHk3LqVYxr072l
3qAVwNQDtCPomKJWhz0yOTRMHVhACqSLerXMpUhCP4Wt4YzSFZxsfwh4kcM/qqnIES5thVEf7aa+
vpjhQpO60DF2lUFfhxrhkcPg4j+9WVnqc5agL5Al3pT1aWwchm+W3PsHLiixOddSscQX4tMOycTw
7JY/yaMmejutjadH8kPhq2975qDwLiu9nhvtA182qU3f1tgBpFBfkuGT1RusB7JiLi8EJwrfEGgo
q1XbTUGiZJkhL5ikGcFNJzHuOPoO6dGu48ZpVa7CXW3kloVH0k2aiq2r9J1URWvfTQpe8Cczq8Ck
mxP303R03j0twOdmh9TDvrn7V5aKiHpyxddpDY28PcolYh/FCeuMWwbjgBlABrrAg6ce8UBm9FXc
J3exldfM9XMEvry4JSN5EMuYOfD0zXrN42J3U/5rZOY27RvQItGEOBUiOWiPcKssDI5gTLE7eUNn
DVpQDxcHNOMcCuPZhXmzdQJPyczknTRGiH8pORlcXvpJlQXElXPKqertZRXpFsoJOXal5KMY74T3
XWxSPAVrRIMLsKYdGiX6VZXJoHV42TNft5Iqa12MH9YLLi0pIiCky0LnCrZuc7cI9C6/GbAEW88q
YynQwrCSNphl7ukQdERGDq5M/Ce0WpQsET3LmFPGVzeT2fEecKYkUM3OWtwPCRGAcUSDoSMsQfdc
nTwyf79JaONhFW2gA/cm765O2F+ArQfZWu/qohYvjBHRhrCB9C/Ky3uWYJUc2qvHa49KVXFMuKCV
IQz/YrLfcwZUAfYtE3r5gc6VsyGSJ972ElACoqd70RXIKAVbEiuGICTdt2iCdGqke7FH24pBQp2k
D5Cu4HRUVbJ/BCE+DSGQS3fzZFTte1jvr/KiVDZeW+o8gglcKdBDVRS7UCpDN7fBzIt+yy9pOk88
CctfAsVjse1HY02IEQdLRiohjCeaf6XcJECcZwF9RkIB/XQlurF//8xQ/vfG3EVcFD1S9JdBaKz1
LLmKRW3a9ekd3Bxu9F8VIEwYdHF8zJQb5Rlio4uoP8d9r2Znk+kqo3gGpK885KIWemiOq7nLLf8s
2nhL11DKdv3GEqavKT1Q+MJ9i+ykEY9fanckzItIyw505xNJVtHPsCpMvsT0L1QMGUFl7lKKiMNl
zhYULMRqn4VwR/336N6HC+Nt/CekcUD4gZyq4iQlfGMfllxQ5rWwNQAAJEIsovWG5iF+nXSfBCPi
4nxOjlj4E4uJKkZBkK7LgJVUDK3eWfGffV+IyVK/RGbO1Hw+gFejviiWwjzUE+c+JMkgEhk4UvgW
ZbkXETZf1cSJ+dglaBC2BB652H+glsrUpgOECjwDjLeDLQSzboDO5LBmR5fR/EVNn94W0LfzzBwh
c35pNLLgCR2rUQKdS7yUx70Vujel2XIHCrtPZxDsDfeS+mY3TQ3wBjmKhQDvxCbqncoNY8NQchOc
uEKe84iu5Etc2YEIGfj8ix+btJZ1Rp/9iV2lVvMz2czy3AKEIJtenLoaXc7cwaxflnys5p5XJ9Iv
NDo9HBH7UUMSAlkNUnxaInHIACpgj8x6ZQ6x3B8aJ6eT6eba0SRRjUc52e1tVxTJO1QLppcP0AjA
KLHjyVrZ9Nsr46e54X6EuWEGi2qT0mPrOZYsrI96qW8Hed2oHs92qoW/rKqDsZHkY3MtKpTeuoz9
FRK4iQ95mS9NZy7rfjZfasUmafPie1AqhNx+Rqq9U4u27ZLTqShD2yjHS5uVm5OOn0BconW0Vmuc
d21crJ8QiQI7TfvHjGw1w7koNoLmJM43qTqlHteyZXRG7q/9spqd6jLFOCTKG5BzJOuGweyhL6IU
vKsckDlxSz0ukF4TUKMsh85lCSkAc6aG9RVhqYNreqU84zMoOlxSQ9/4UwOaUHfmo19xE00ST3kP
9sQUlfVstej53vac8lpzNsg47X2XKsaEcU9ij9xeIrMh41YGitf3Q0GAgif9az9vUcmogmTm2f9k
IQXijs7/XnddIlEtIyEid0JWKKNeD4PXdLUlzvOSWU/bqIuyGUHosLhFh/dexvnRIt+JBMjw0Gij
ypM2OHXiXt/mqPyDrkfY7Jjla4YrvgjknGsZ7hi5UODQeGcfrF4uMqCEGWUb8EcEK8pD/WLmgagY
tkKAQWcNjSrHaXQqZ20bHvzR320qso23/90WGlQ2p2lRR9ZdPzjzhybsrOI/RT5SWaQ3xCxF87Kk
PYNj02bwAD/goGoHcaQD7d49WAys/fh3HEa/VEBgqLjsEb/1aBhnuURsLT7SoBWLVogJaUxJoeyl
xELbt/miUKpQ7S3+ZgkEzCoJYjD1rpWrU5o48ixawW7pTQIEqwA2o7TUdJ9f67CUW+Y5jMeP7cXM
DAbkXOMSSlYy3xaS32bAs3d/sUypv7hCGNAQXBaYVCzY+3YWshouOl3jGRj1squXEIaT7lObx8tI
gKKfHu+6j8dmCF6+kjwQ0UNmHEgj8r2i4hHGO4/Uf3z4BfDD3b96VSzHyAb17+7k+9XO9kGwcVT9
K/qU4daia9jaTUFw7tUxil8aTAG40O4AoHs+Uf/bdIwxcEt68ZJS6f4Z26dPsvUtenmQM/Mo6IQD
6XlGOtPVj+Ge9T8u78GBvkGydwBeWtGrBbUzSnSGgxTZNNBQWw1slA201hzsg5DQLJu9SHCxdmal
N5d8Y8ijrAv6OYmQNtmFlU3T4k9iQQXCz88TUywS7p3PjBX/Iackh9VT25XnhfKr4Gc9/LOlnvFB
B7xWbCD+YHLSJd+6F7+hUbwkxcX24xGv9u+1/HL4eLJLJKDhr/71MHbgklofCGrcPh9AmjiCPq1k
GEaTIM+SqNUKmxe9wVSApQJsxIB6qffb/8a8/PD1Tx5mAE3+1aAPOSivlf7nlo50aZSbhoS16z50
vSXu4a7IWrWdezeLBzdgv1BFjcI3RD+EnNFqfOWaRjj7YVsB5RpqmGm2TbXQlUhTQhmrxnXEBfzT
jei5kZzlLRV0BA40XiD3mohVlx9f6m4rPQwmSnz5lROAnZs8q6qxqFIlGN7pyi4FPuJl08dMDIR/
VG9MHFKE9flxbEQ9RDGBSzqeDLJxFiDCWgpFROdRJCHl3U6rbc72VMKfKOJV8PoZk4KyV3h8uuhc
Exmrp0ocqXau+BCp8AWKUpWxAhFApFThtfTF92KPyVG0t82kiDqAQEjGkyll3bQwq/xZVZ0/NpgQ
wVvZ322dGts/b4AlB5ubW3BqXdJrNvMhCJB+TgD/suAtDbNl/dzAmUccTTuw5/hVq4mDsHQ6lWmt
+yA0+4GKvq/gLCZ8waxm/Xr8FxwMro44eo+JwnM0y+1Dc3ZSyS7CatIR40cNc36od4unayPOJ0hn
MUX2HbWI2XnirFAqfBJ8+mA7ibEvdIMIBAZcdy02KJArsZKYA9yJxcD5wd9iFs9BmNC0/6/nRbbV
KUMEFOy9JXukWva+ozVLmpUkTNRAZB/Fj5gHrJXPoxtxn6XE3KqWP8rSxKcrNYcVFviKnTBxNUI+
uM5VE6lpOIi1xHhSxiI+2CtYj1O0gwuQzZ107t4ODu8iDDUAg83ayYOcvFO3WweM2Y+ac1+g04H7
BKU/CExAsE+9Zm0p5pWIOx/bpvD9Cb+mRWBKoXIjONQsx7TH8tXznrlsfeP/owrqzD1H4VkOhvtI
0spQ0M3HvVKbAbHGj6532VZ8vInlr10CQyglkyZIdUN3mWd/CVyQmQyDngZpdpie0PGDUwGlnLIe
CRCezd4TsL2vecbJRkHAkUqVs0XwJWFhF4aYl0nyla7zXY4sWmC3a+/8uK9xmvSdHd6CzH6zrxu3
83WQVcxmP7SQLc24NC7eqZ06HUwx18ITBgy2AbZPh4PDg1eK2usVERZw3Ms+9FVLZFGu1qBwi4HX
RsJOV2ujtKp8pU1Dd8w46gQPvQWW0AO9vz1RTY2E6UJeyzVlkBP3QKrKpwCCh/3EMNAHa+rNe/4d
7sli4VSv1qS091ru+ajHSiY9OvbzVidmV2+NVsnfce8QlX1UeIjSecSI9TYwVkXg+ATA1ZrOHbOc
0qx9t111YrNoK2ok10FA0/MlukEVccQx4qxFPBqLNnLSAYrdGMK6lYnlFGoL4r5H56wjaq6524jW
UNEN5dg6VS1jvtZtqS9WtV49RHfToEh3InF7rtk+XbtvlrXYhjmrTiCOoIeAGAolTsxgAZWUWA0C
4Vuz81t12oiPL1pI/tnAZFhA2fPxZTh7gN72FdNFrA+yPvVXhRnG1dyjrHMgPDKocm/ORTsxhZV1
JR5pQR6jzC2BdIAkZwxT4nO/3U8KjGp66SS+E29ox0kgarJbWp56NtauGi9D/xqGOkRhhTMrOM91
kKlyZmPkUqtBmFZ5gBxc5OHlj8i8BQh15+SeeWnhmo7HAFCCRFeqY48aoK8hkBIoeBq97Ymk7AvZ
IsA2wX2LxnxHfcGJpb2bu8lG2lRp+DQmXwMx6L7WBMfLqJp+NYTe+v9olPTvbtk5rM88AB9Mp3EK
Yb8hmxUqT68nVCp4hWVhADjRb2rEBJ7kPui6nzu3QIq6YIkj2nmFQCV7HNTshjR52ggtSGkewbSc
U3SydCcdy/znAUDLqAnTr0ktBOd+jl2462NeVRSk3Sr/00bswdUJou+wjXmQmBTIcLhd3M7RNJlE
9OkK/SWaKee7o1+4hLsQnpmK1pAuqyZKgb8vriqT96lejZ8Edn/rnQu38nimGT/rSYhAMWe1rIsZ
c1nIXAGv9T+s8q8Is0oASxjCpZVUCMtKfpcgWZdt6QDE3C0PkVJ7gF1l6VuzSLVNHqB1WTUcHnTK
Fl2PIdZPMx9BhTMeb6neH1jREuH+9zd/PUHFeiIRYYUIP16PVfDQ/yYIKZ6zLjt6Jc0Q+Q90yyCe
dkRKlDgRmw+cvBttDEG0OkvmSYP0FIN7NeRS5CWfB0CZUzA0sRrgn1JKPDrgS8f7DNVU9HMLuUw8
WWyfPi74aBsAj+oARKIk9L4u5My2v2lRZbOIGIDqbLxlx9UpkqVOFiHQKjJiK0k8MVkcnAmAwmRQ
/vNBOZVq3HxubOOEkFPUKOXpGtzKwyIxsLGmzc5dpZ80QiBcclt4KUiOUr8lRT5zoydKWPJ43HUa
1ggajNQGF5cwKVyT/GENIXdj1TUWk5V5oVIhtqLAGUNtwJ+vi4wycwfKb1Ue3Eflin1C5K1iu29j
akaJQ0yCGTeU+OIPgWibRgKIV7UgrICY/5vMJObgUvG3X+SVeRClsIs6z5duoj8TL1Om21qZLw3Y
6v64TN/bQiZ2+DwuLaf7RhktEKBKPUKaILD0ExokuOEBOR08X2HJ2bg1pX6ak5hFXapZZeEyHyKn
I6xmebWSCMEjtEU/wfjZ/W0d7gJVWCKjegtv4aDf4is9Pk713nyzT89sc1u2hGqjKI6b7HKLP0ih
lkguepMQtfOEpp7br4qfzihsZ9DnJSBxD5eBx3XmW3SN1owqvL/DipV4FEm8tVr2PbGYC5SIqg1N
u2jSOozkPAYRHdUw0lNwTK7xVmyYDhYfPL1p5lR+ghP6BGWux42ofpfBL0j7vnC7sIW2BC46dVwx
OzZ77wVmZGBmcX/4e2N8Grq7mHujDd/E/Qcpn2Mgs0miSUmcJRnNepc9lNzUD3oxqigkZjiLU9MN
7lzLznxKHK8oXEIg4DfZAzGCx1gr+EBNQPBUil/jQgL5IkwvmRdR6nHrLY+3V4mkcb+yczIETMc2
59jGKYNenF4qWlotwFv+1gKBw3fIl3exPI2uAUyRPopK93dmDdo8KNT3xP++w+P30Ddzhu1rsVT4
NThVSL/UHpL6pa1eb7E4hsd3SyMR8UcG1Q9PTLb/7SMwcBru47B65EgtyV6D85da4AC7Jf7NeO0f
2ufBAcumZ8EaZEoFU6VLM2NJiZJlsXtdMWPZRwA62Gom5n0YxXGsh1fBm9aCsmezrED1APCIUwDK
Di126Fu+Y9uT8Hyup067T5Kkk/fqITx92bpKaKDGV+C6KomqlDAvG29+A7k9ZtQyHQCkGewO7Efx
uaFHtKlTnw9pivAICFa72dgWILsPFCe68AiSQ+h1VvDtuKHXTiP+T5+XLVRiYQUcAmSXeMC7GH4x
nWcCnb/Tohee8ICawNBUBSXDbmrGeTOYwl8ERtPQohZiug0nnYbodXUS0qDG61c11FuztrIP5Dcf
/ZUZukpUpHawt045j3+OqvmtHsfaKFPCcxg745AQONZmq/NxuX4brKsS3aqZKmM5FVk6VNdC5fgx
6xVjifuLVD6x+VprUmtXOVS2b9hSanS1jmddO0oECubsfvGheEGmHF4I7QvHrmCAyJw/PInH908g
0s05ueM/Gavde55tyI8F8/KQjZZE5vIIxStUVSQDziZ/TCq3IkilV+hzc3tSz86bNJdnj+xPM6xC
LPYXEkjQ+ezSMtXSTdwTtm/J1TcqMGMG8uqBWd2I+XK9/l9UIUxuAySuiizRQSdtSd6W6T4FqYUL
hnRqh1cvTByxxh3fhZTXn9kpTvQFoyI28jcT1pqMSwMkRV+mrKO5Ds2kSiNNIjD8lZppxk7xw0ZC
5pHyKnfovHSxxBnAN13Qb72vBZgEP8diK9UYugtBEYzOIguHcRMoYr83ilfmdCQCe8S4I8UEaxEV
gxz+pUGOZolV5jxni5PDJIfzxa9BTksLCQNpeq6DqlyjkXJkLAYniVP9wj88YS93cTHOO0rvrkqp
lh/QTWOCjfLNWkpb3P+UeicoP+ejk8+dmpMxNaGifeCv9zqbDpyZwRrzEKb+VjaZ4hNx1OLNLwGi
tC3S9K/XCaIpWaS/vnv60tLMBdGqDBYVgvIwL/tulVKCjQW9apHAfNNDlTHoL+Fv7xAr9qe7/7XO
WK/o7ZW8Wr9FMwGV3/C2bXh/wZCuD4vhxOh0IGgg9vPjRxPnH0+Dh517lastRoV2E+F/3ruShQr/
Zs0sdsOpnaV3Qnym+gSgUjBB6oOOjte3KB3YIq8AZIAxhv9BgFhftPLRFYFYqMtpH5aCyGRuHBRi
yWclatjbWcV83mp57oidYGUyXfeYP3Z3DOSrrvpy3Gv6V5zxoIhWekl9+mNCXPChV/fVV9CA7N/w
OP4h6IfznlUvMAN9AInlJLZMLCFrOV70cinwEYjtrYBF7YN55JthIEe3E2AdvakHtdgo9PVysaCC
q/KsxvGUgBgD9s/+yhyjyXhXRppU/51yLOQJglbEIwtJ3lEWoIBXkMDpE8FhhxlmNSQyqfI9PvVD
KPeNPJ5DSXe+ZCJVeP3HB00hvL8f8wxCrV2TrgW3mwFspQ+3YbfPzCdjIUGoBAnvos93k0fAZxZO
EqbpeQ0FBJa4XEdI9RDVdYtZhgkYvBw7K2ZWbkvS7hr3qGUerhzulH1/SQ5Tfz8H1zXukd1/SZwx
Ora0tNzvsjhe2gF6P2hp+ylafky8+0hsW0R4rKTZKJsal37bOAa1Wrw/Mq+kU5qFPE6a/b/Kx7Fv
TMnlSdQJSBJpKc9O6wSTtDY6owE7yquCcUKeiC3hHfv0AneDutGALV88u3hX5kaD5PkfIfRg7SWa
STb7ZQUbxWs7R6fftsv2mGMwBEhl8+KeRoXQIOP89wXx73rpw85RgsDQtklNWO+EGiSoYusQ8mH/
sl1C3Bzntnt2eFK5oWxL+lR2oIMGJsFzZoMlMsv1cV8AdllnzJFjxKbssHUYSCNuqd8m4AJsrU9U
yJR4DuxGf7CUGULudLXxRFRYdBXbq7Btr5Lqad6MlNcyOb5vcpcKoUWV/k+Pes5gaKwkg+LZfNis
UAhe01j278AJGtT6HK6b7tfF76+X/dnw9sZdI3ye8g3GE79nUAgfSr1l+EO1kMkoAtnb1Jmj3+tG
odScKo0ocZ/pOgVSavZwFKpFNLrp7nMXHhxa4CfHIEpD61HEh1sbMCX4EJmmckk8dGdc7p2YKhoN
Xf/6esvi/adVfUt8OwO3iWpnuffGu7Tq12uij8pmRgm8a/V5Ek9CVzcnKG1hk/YyvoV1EVgm6DR4
NwIhKf4SrLf1+fkEbmQIHDO6HQ6jvTbpL0EVVdQWa7TL+xtiRikRRN9XPQXqBGDsEJvdDmRNjnhQ
ZeIXvNZsjesDUUBnq/vIi1Rqo8Xh9bDsuLkwj2th3tMzby5ZPqLz7rvsJu8wNy2IRV+5j4wc1ZOt
a7UUi33VOJTvhcd87lKYOJQhONj+wCbWStQz3HeeFlbDHqwOxQLI5MlXgv7hKNF6z9crijXERp6D
h/vD1aL/h0OKpZjTOLHNL58fa1fMEX36benu7cLeXCYUkTpHg9Q05PNHzZW2hBgvK2yRwIfcwylZ
zXYeB6RMfLkMqZudhgeQOUOS2sihES8+f8PrgalbzI4lz0d1ju91WGdgQ5hsElUMcMZJ9hjY3lwB
IGgKZakMcb/H7iYfk55TMIheS1BelRXNJPT7SQehfKu8XWaHerhHdWClyHf5kZhw0/Y2DW3GSDBk
tRTDKQGzZcmiDm8eBQ2vrO6t0m9rLG/SpZ68BW+AAhAbRqLpaIStuCDydi1LlGt9KLwkidLMaHML
lDCqTTLm5XkZlAGfv7cSrvglsTol8BkSH2vSQegBK3E8WfD6tDO5tuaEj2lor6WXuyB0zxjRcAad
waQ9ngPd7Ne9UTh5n/AKxN350AlMp3CIV+ToENZXPpGDHRDnbSOT8/m2txhlqsC4JPdTwkbc4QTE
NLEWIuXJqHhVDodLzFR8Xxt2BYnYcuhvXY4oLs5kd7VQyL3oBm5gJDp7Gz4fO8Zcwnw/C9ciaEFV
2rhh78U0d+zsACGASipDr1ZrfH5sWRcEXxh7/kNgrvI/RH1Jym4vIosbZV0koRtqZjT446qRa/Vo
GHFjbZIWvS0VhqkQ7E7S0eNVR1xQ9qfUqlg4FaZpuLoMN97pzzoIRYFd3QH31SZgza+q1Xl+r9eA
0VF/kuO4iPj7Aho5JyP6zqo5OCTnUPbeTAvINO/inxvhE1A2eVqbAmtJxpUfnyhYoRWuj83JRujY
Beu81W6r5wrCRjx+UG7zMePZMTiYN0ZuUOXmKE5C5MqnhOHJWws+OCJf5B33cXgeE+0mBenVxIzh
mcR5vQe4/tzpNLyRBH7NF0+a0ISXycFp6OtzRrNa3Uas91qW+Q2i5o9FYD9kBz98ZDGL+1wyv/aj
SMyAsavDWMSEz4jkwCxgonYddq/beteQcJq77Bty1DMID5uLYlTmf4FN+QyQTfzvfI+tI3Bq1s2i
hI2jcB2WEcw2Pwy2RY4MaY6mm8MA/IwWWwaoSxZEQ4I0w7tnVf2du0583wlydMiCoc6qkAz/hUml
b6IZLqc5YCWL/hzELYZjA+UGl6yjZRymcxjackTJawni/A6VHL5duumz88C5ZajuFL2obCw3Tx12
s8Bv22rxy/aLY9tlaJD93A5Zi/wObOEIozCsrSadf/ALld3tuG0x8Gg67DCiSeaK1tn8vgOAraJx
chfpU2Beqj0Er/e1vLxMF9rSSg75Z+VFgRALwXbUfP0W2UbhxpRouNBjFwu1RMAk0UvPDHW6Amr5
DWPr+8TZfVrJ8uvju/cXKGn929zUFrZOD7uld2HRUD5xrmTsufVN6f8LwlNpW9nKG0LciXCGkB5H
FqIdyYj3sOdol7EgrICH9JyAJEDSAFW+PjgUpITU0Cx8cUNXX/vb93yUKcdEjJFobTljnL7Ql12C
NKNxgmhfIcvZ8K1/QAj3RMczpzF63U0H9dmcYq1wsEabI3EdhgU8w+VqogsdtMHuu8F3+guE7dj2
WzOgmtJBVRwcpyoJ21DGRN/9XC76euyrUKLRZGnmsDQIZqnWLwXvRIeyjwP2KN1VLouyqyiYiKNx
4wL1db9Cl9S8SFw5MMdKQ1tyVizhRLMkmSIA5Q7/Eij1vs2uBGN6gUwRKwGGc0W5kPEyBJzgyHMu
8Tsoo0C7JBM+V+rpWf1wGHm/XuQcOYAK0HsvNCsLzUJcghZvcEwieJ/Bb/YgBMjXjrGQNf6szD59
b4pJLfzE6PcNkXiYS6nXK+qwzCSB1I1+M0tW9eobt8HS+EBMci7uTwExN+0T8kJDOZxCPB3gPHv7
2Q5zupVdERnDtMFj+T/2/pI4Z0uCcnPG9MeVUr8FlvLrrM4gfO8WKXJyVpNS2uL+z4oI7c75M02V
ez/VFf9iVrHzXrS1+n95O5r1aaFfwvyxyHP8FoUkkdAUqUk5pSXIXNsawFNyVc2AaY15px3y4QYt
POn6KiTte2bTCsBNEEbDiHNPPjPem6EMkPHp8kOtgSUVpC8sISOmSyIREuzURR/masnYzqLUtAFO
bZ6u/rE+R2R1NsJiIZ16CAjObq2PwUaSZWj15w5KwWuiFOuBBya2pRs2BkLO1FNFbtXjVkl4pt9A
lXOPe41hDR5s1zTxjh9cpi9ITd9meriSL8KYdOcia9HhJ6muR4kvUNBnOSEfE/zp2uFKdWipyG4C
CQKmy3AH8Q8cE2GSVxc+nKn7kIMiuo/HDpcuMGdQG6pqX6l2/IoyRYY7Z8ez+ZbPr/uyT/FX9gBE
/dvF1aIsdDpyDGwewtlzmpGywJ/o4QTxrN796BCKCkdJbqURdgNfGyyVv361RmXD1rAPgZYO+OWG
aUT7zQGyyt4kZN7zoInsldjYlJc9oRdLenbI75l2+Km6y1iZLSiSEd1JsR+y/YxWY6rF4LFwMfnp
QKZlWXTJlSaVEqxVQUtduASUvwtiP0caVraiPzSaQGdmpagTu7qqq0icqfn/O+2FVXpcfM/O72Jw
fme7z+Ye/wUNuHlmqNB9bUOi1d/HJVRRC8m/sHRdhK4JXsSD0Xu54WQPcSXAYao7ujxY/dRNwkym
dM80OAQlvMdx1YuEKrGe8TuojtAGiZbbIb90RSViROirzpNsZw7heN5vnCktVNTCum2T+h37sJ8h
GCQJ5CcDtj/aBX0tHpyjUFffw3QRvELCm/jCOvO3dBEmRRrphPFxP//iMFRe2o7grs5OEJ3Jg9zG
ftI0fftByE79XOG5EcDnxRU0mGQazs17BP9Xwfsp4m6ccheA7ThpIX3AOZHhqRSdyDqQ5VDraGWm
AS6r1hWWBGiJLV8RNIZnRrTKt+Qw88EyODsaPIOtbht+KpYzrtCpiWZceimdpaTxTK5UZf8ORccF
9ec9+G5bbWZLk9ccWzDepefproLlWAn6p/eqDQhX8st7tfLuAWltePO4/DbmEw+5dxNdd0UanWzB
wq+gM8uBVW8lDU6z7Vsn6w3AzlTMk8Jj4sK53zoBquPX5slrYDawS7kA6W5qxMvdYN2/Gk0EXOA4
RaElzz044BihOPqX1s+pjsiR9qY02uBHCBSBdJOir4Ar2XeU0VxtYx6AbfF2/UagNJ94avrYLRn7
ZWPzMLyNI3Xu4ZK9eiB2HYTManX+D+cSNhGJKKWZA4oJ7pY+lkLh/0Y3pGPipwsQQ1lksS+OgxkP
lMIfRaQa9DCoDgvDXiXdZAAlsZvXnKmlF+hZFEkXkxU5OwM+GN0Lfm1h2+9vOLW92wnFzUEvIlVq
qz7zH0WjHPbQi1XTNR2xZWbs3b0tzxv/9soQK9Do9tW6pGgHaStcWIW9xBz9Omxt49KoTtfH57vX
/O3SFjosvBfTJ2S9IsYraTchRH5qgm+Ow0bkO1YVtKd+WueW3j0t1oZ3fproXoj/hyp3DYsK+ab7
KUUkypa5SxM6YhMn3NAfslcBvCetLuF20t8vehSosvtyeGt+PvoBvEcNqxcYFzlruAp4/vHdIv/l
2HXNqkyDWZNb+Wf1fg2brsGcENYeW8xvtuUaukvbAhh2om2RyenVvOcuCnd64lTPgIeeaqE0Jb+e
fTDawJJhG9l9WS2VNjwXhGq3a7B45DmvLu0kzUp4lnn4sW1E0ja8c+47XJ4psKC3pCiNUAduBpGi
eveel8PuT41ehUVclkwV8DhpyV7zj40LOd2ImvjfLoAjW3tX8WnUbclT+y7pV+EGiKY1zF2YMJ5w
i5VGwMwsNPnVi8qgqnEiMjp/H0q5Zk5PwnDx487NWDVdLIfb2dW0kFvTUp0rj2uYRLxCZiFIO1js
9/AWCh1K7X+OmiEc6Uhx0eOufh97rXGCLS7x+qGdgk0y44q9w7Fy8ngty6pHvt/g6cvlO1y6mKBq
d6iZjyYZkqmkvMbLAXlR+oM056Th8GqHn3zLXgx7eBuVVDF5JanJp7w6dCo3dsRYfoEaJTf85T1k
BZUKxmAA533iexARTI3f/A71VmJGUVUKik0sNtnB5ekbyB84aorfhqIvmBXWQotl+U+FhSJBSyo6
EabIgZifDBk/0lvbECqCkvOjQl7gkdeowStkVM7JGsE8LI2gvwcir4jOKbsnjeU1cxJYrwGGUJza
L5h7/PShXCYR6cH/bmw9Cai7AwU+HMsZ4nUJ7111dupWyVqfmCGAPKnb/oXB/zDYzHX9tzretpr1
w+txR3DvOmEzGD3atdGSPzWzIJWBjtRyY5MprKbDPBzjLDNtXFjVAFa8OOulLiIvVXcDLpzmaDtC
oUmhtAFbOCxU5oA7zIa1/tkjNSwAKHrBaThSvT5uUKNpoOyf95+gEk4p08Cx2aFbLbQDihWp4HxN
A6WJ/zyzMG/9x3ATgKjtgoZ2O2+fUTY6iP2W2bELeGfp4ttsQAsRTpmbWiv6R9dmUe57VdVnAWTW
9BQhsXgaHUB2GXLVPYs6slRvT+1/4yc5DaPwqJk6SBfchpEY9skVw3ZOozhK3uHu/JKYIFOlJO1i
Kk+wWtYLYtVZSPp4/dD7tPMBPZQskZS53GwSvcOmSa6zZ8440lqfn9K4ZeDzFzaF1muFeq5qXr7x
HqBdAtd7cbu2OCHBnIjC8vs6PdX/KPfIPbZcD5lQxOT9cIq75hEiwJIi973HteXltgOy8yF514Bb
zZSkX7fkBh04yiegJ332RoG35B+4L/iH23tQtg1xmhNdH5siimSQWxweDbp1e7rXUm6gKFyAOS3Y
+Gbp2yFigfPW5gGGiBycjld2T+SexMVebHNyuirMoCehBwmvwxHGE8UDBPP1KO0PK4NLZunjtO3L
l/Ad96ghZwa91gufwaSNkszyY4RaTqZZtfc8CaNTVJIUP4kpEXug1HVrKT3YKHLaHa69xrzq/h0Q
ostNKPCMCkS4ks6YGZnmLxfDF0bGY1MEsNXq2I95IKXf8pYZNtahXS/7VfvoQsJD6w4bRBxVFBzT
M01CNX7ha7rymfsSaO+QXGWTHAf13gG/d/R1cB4WEcde+UMgNMZall7XG09ZtgcUCo2UeJh9Li+V
r3C29TbXWBM9/I0TwBqxxXDl3xkIxFY+0oYGqUlp+bxal4I60an3gxtGBVVCDknS3GEoWUiiF5mx
fQZXVKTs5Ej5OX4Ai9WXU18WITPxGU8pnRC6xS+nBnN6dea63k8VlyUPkXTfK6csPBz5UVC2lHml
ji43XietTUS+pK3llV/mX7qUEU58xo3xN7cbeLaocwqcOr4qyUT9uCqKZwGduPZtiZEVVVPea0hv
aH/l6i+xMPTQmbVbVhROMCkgqYdRmEOVv0dtjaBqk6LGKA+Dc51PJqxJTb9+Z4xa1Ev5ocolhdah
yjyWMwGbEBKByVSKgrZzPtPmQhfcMo+zf6RSe0Srf7nam//7d74I/taonAm8sgvs+uIo9tD+rbqC
kwR/DlaQWZSdJCd+w569Ku7b9qH6Lazh8zPU4DERbNhFJYm6QZ+yzRzCBoMocuSA22yaw/95o+kL
lIAez7722YPayEaWfp3EucpMl1/wT5f6soGvpsE+XhhgfHT/FKwnRGHhVK/SebW/efpXAmSR8kKL
trEwjAA0bK5HDtXrhnkzaj4XBEEgDBf2HxtEX516LvnBGp3EXjZWtvmqLgV03czGvFPg3Pgkumw+
ebPfK8JpSDwUigw6BWio3A27d6bNAEfTLEl1HWxSKaomHAIrhUHf8dxoYlyCoCTZPrI76DsCiFUE
FejyU/zDE0VHs8vYn1qHAbdRTYvK0gIQ7MW2HMIHeFFzMf5RYiFNjwxzU4XU1rbhJlLwFJ30rpgR
pLklt1FwWXFEDXCA3Z8zhvGhH47PGs9xAiYNRcx299IgRpeOdzXf9552XGdLQL0/SH/5KBNYIMQW
ExXcCcRFlIUXltFpCAryQvw6TybZplZXXL3vv/ab8jlzAFG4GSbNxgwcYQWl6GhXRqkSVnAeWEvN
scDj7tRWwigSFZKsD+Oo2arYRJ7zWDI72vdcPCsbAJiv9k25H8HKagGCbD+7aWlONzQJimqeQrkZ
/DUH1RvKaSehwpPORING1c/WT+VqX2GucJ5fbUfa1VHq17kVc/P2mUCeHueJHelA8gsp4xx/KAQw
l5KsmbFAKl8ttucrRxFNH4sa1jD9pH+DAjfD4L+c3ljfv9TtQlKGR5QSYjUFSbT5tUnlJijlC9zy
oHUXgwGrnNsTpFEQPSQRi+7bfecgIL8COyeRYIcd2uGvtx2sUV4mOcBArgVB1e+uc7WAZxWN5ZVp
Tg1X/S2EqGquE8A+7Yu0GFLlYv/FmhM7SvEHcrMR1Dz8ASmtmupkmcOvoY7Qf9dtykO2a36GyQ5K
Lz3dQF5mcx3VtcCyXjrhz9LinngZO/pgVVuUM/VdO2gqEI3114g2Uc4ON7DfeH+8eKx2sb2++NIN
kdVLQ6SsAp5yAoNbZnV5dkxzLIO5oG1yfrVKwZTI2gXd0oXH83Yk+40cTejkH1Eju0La5np/nBRV
RnJHMefOUaTIzIRfqzIvZUoVtPcyLwxqsLAx+JVBQq8Zg8bBY5GmVhD4oD3ZgJ/liYwv3TYh+ZeG
mEdE/aRfh4A5sUK2H6cHUb8pbFjxaOjTjjDW+QzWWHdc8p5bj+ZdhTDCYtDhuX+5v9lNcYrZx2zF
fVQxDvta17RwwTkNGNI3aHEjT5JkzNYfvIeZll5Un1RhCAZ6qTkx98S8bCchFtjSoAKwO7/8eQVN
9gcNZqWFqSoI3ZI7BG2CT4jXVg4HtQcFp8u7GLIDq5K7bEawNVgTkLJHRasE0LfIMUXSi9qZrSqT
UDxaFJKbfy/k1DL6zQJLMFzMBScjg4DTgM6q1tQSgr5F9YuaDP+5XzxyU5QL5VG1LZXoGJK/ELYB
rC3LOexvOja0ZwergPOOfa8lfgCd9Hqkc4wYO8dc4FB9ci1UruNe6QBzwEo3ddnhA0l9HplcB4qL
oPtQ6qXS8Iy8HbJy0sWpjMkm6LDyfA80ccBpIEqYZMJb8OYyfiMTywJtd7wEmBvHrXlpMesl/Io8
Zh6IK/lNqI10OZd2mD39G5Emk0Yon13UIogBlF1sKy6tKeQuCxYYTBbpw4nIzSMnkSrZ3jiJkPFN
XhQdYMHjdu38UAVXixK47tW+s8MoFdhi6mQnEfaPVJ4PfzhF9fKVqmLxXnB4vP6inXkjPB5r3Ad7
ZfwdeeGV6+8sgF3CWF21d802bCLYv6fvIQqvBNY0hb9fclbmscMTrpJ49jUrVbE4fDjB/DLiceE5
Gc3vX1TPVGZm0qi9sczgokYcAz2BIlfukN8qIhV1Yd9RDC8gpWw2OVKMpQrMO2TrAdsv19VjqQXO
sA9byjbPB1q8KT+ed1OC+K39D6mj2SSIyaT8fQXCFxHmOHvhN7qvlK7PwCabiTbElTBTD2BrxoEv
prdy8zxnagkUU0EGWvFimTlsBLj9MtuE/3YgI2eyDcmW0m1nhsOHHGF/oeMpBw4QibWLotmBuSrP
oPT9chW8fARpV2JfCakluOGqiRcbkefucGYhjY3rpIiVSs9SJBFIXtJJHrU/EV8SZNSmjRSBnitl
bgCz0lxkCS9QzXSDuxMZT11BshxgO+boPYadlA4Hqtk6Ld2TX7JGDa66aYYtw8L9wAZPdUr8e+7y
toIJ5lz/HTTxtdBFX/LQkKmuHLjE5oUhmAmmIcZlbe9pmw/FaBfFdHJ7ntVIe3F2Dx3d4qKdLZoO
ZuHAIrQAlQcl0oSWc5gmaXMIVSySU4e2knChTFilqQNT4PM0a/i5x1gOIpb+UigmbLuYn1BDVk2g
i4pqzj13WJtf5z1pV1sB0QsKbX7EcAZuZLnGODRlorFKnMX/IzCzpwBIgXPMSz0/AnZQah6rIUOi
VhaPPnkRs/aBV5a3geRb7IURgNqOCjTB4tfFEvt2NtJy4BnNUPSVe1QmNPOw7bj75G1YBdlCUv6s
sRibcQpV6nStaM4WVjvVNbrc5y6ww6WQpkxdmOVGyQGBVYmd6kj7/UP8MzSDd5TphaiQ0PrIEjte
cTRip3R7ECSwYrIx/x65tvxEXbofBpuacyV/npRr1576hE2t4UWE646IOG/sg6q5z0J1prsm4aar
TyTIQ+93TGiLlmIDcZVAR5E6T0GY3/nhNFJbeX6OzrLEz0agsI814cZ5Ht3mC3dW28H1GV7dhxcI
C9bjaUhDrmYeUjWZmRdlftrMQ2vgkLBLDbcIrM/h9p02pI+NqEuAvZ925xCImCdGLvJLSsoN7qP+
XfloVWxYSoTNxpGuEsyYXe22tCufGBqN5R0OVE5ABS1AZsgNa9HdNkjwNLrDwt4pRPHZgwMVn49D
m7YZrpRiNF+C0+fmr6nJJ33HhaUTaSv12Cb81W7yeQSEyOXNDomLtS4YH5CwdPds9kcB3uk/ZDfe
Dhf5I6f1VUgPVtiDxE/lO8UF8TkK3q7kh9nF8gU/nkYYfLlieWPrNaExih+GK552d1eeDRLoTdKv
zxTGOw2piMsA6ZRNcEYFkogAv7B1M6+A44VWyAijriafaooQpaNHP3AY6mvWEAxDhcT2odDGslax
6Gy9NUOvjqjbDqWsMizMdTI6M58geB/w6gIu6JkxGNCOyZAYR1C5ASsVtnnsFUPhZAGhWxj4TXFn
9FMsO3jpSn4QRAa1L3tUfgSoA+5eZ/uYqzC4fCWwIYHumAihubsfqUgrfDWzW1ay+lVFnln92xO7
kAwJHrEvNQkxGVcanq+YVz1Y4jPqetZIlPP3LYbpWGY6KQntMIeFGCOrlaQJdGd9s4luk+X9W7yW
ZnNUB2kMtAXhPS+eXKE9zgkGikC2C7Z/6rsosxiCqP8AvPMrhJR9NtvJFtOY9of3SneF2svvdUdN
kciy2PUkSPvwcLP3PnZp3NKjhPbYNqlAuj4AEbCrWTbymDwaN20pULnbTi3qn/vMSjvO8gPPl73c
unbMrtAuTInh8vjoZP1w0nxX6/FCsBAJ4Dtk/5HGnmx5jo5ln96CCq8tnaRieXqz7PxGVepExUUN
wT+78JMwxgpdgehWDtyZ8ckNjBreZ/LWvkSCD5EQF3/cWq4/fnLdfI8i7wg09ocV8kCswdZN9Dqd
jTqp/dh5vyIeJwSHREs50BoN1DpQeIFRJrvXYipK3VV/rXbOtC6U8BGBQ0YlD5Cb9x08mJFDTQMf
TZ7Auk8YF+AkoRnRBlYlFAmLnt25fU3IE34TGHHJFW53vT2LT8Ci59rZdo+6x/YM/CV9diKGpJS8
YhtbnmbiD26C3xjwsqnV4q4aChQ5M4sNg2iDiq+1wa7Snvw3R47sXQp0Op9kMbsV42+F1AlqyxQG
l4azQFrtikpfBGr2DW3Yw/PD7xPc8Wrsfk3wkTIQ8PTnNlM1thUVl4pU5qFCvtOqB/KyRYi9fAkC
HCM9OFVwTpeWX3XeOLdO9xvbYqUd3nRz3K/TyTfAYX/RsjLZwJZbOcWBIouDWIOKbQoIKOhLbi+5
znzFDaSe5YsKYHDygO9ZBvqg2VwHnJHKDEv7el3V7JuvFTJVfMk0wX+T+3CksHFbS3xoh/JaLsqg
tnJbHvy8wN27zxygCGYxar3orthyMA0PdQuz6qYhmZrTuF8bCtX40fv2pgaBO3OEpiS3LIMhfn3h
U+R1cHg+yQrdTJRiwDLISMRvR8eqHbg/xo0f/ioagTiB31xiSlJcoaVY/rXA/XOX2XK9d8xWexih
dwCAZjH6UQ1WuMr0UGvInersOuaU7wvvVPgfnVWT14TtI+g6eV+V4GGlpQWes62+C+rOmYgK6Gbs
luqjtIPDuvSv/8LXv+M2V+h/uNjhcfkApW5MK0ifTupBOEsEhGxKgjomcY0lbsCBIwjFAmsopxnO
e+f9+u4JycthJGN61OPLY3C6t2RzBtHzSjFcCVjjInBsyElV6aF6nUW1h8FCABEaGc6cEhSCQG6M
H3oit5mXImIMlI96CG3vZ7n4l2UiW5d4OpHrZsx1IYxpllLVIRhqrYqrODePvZWrdbCzKS33hiFc
JJU+lwvG6s3CP0wdvvlyPZa5qc7yWnFcTGi8LDcLv8UEfiJjKkZw/ILWNjpD9udOBwJLW2EqA2TB
aCOI02ctrAj95i+2sxnf42YW2vXZmGVxx/sUpnvT83dLmK02Cw5sGfpknLc5kkKYEw0XyVQi2cN+
HqNSYwNz6ReA+j/rU3K4FvLclKjKf5S8afzX+PFs/Z3HqcYY7eEZaJkvMSayiZXmcW6z6U1o31zM
ez6TqaithnF8AKiP/2/FITIbj8TqleGeErVGbLWQc/TsilPLCVG0/txY0XYipi4Y/XdaznEOk9ao
fzt8hg/Nc6g9GB11JPGD+/m24Ah9Ri/N9aYin2TAwSDhrrM78m+tvoovqoktS4G2Uqbr1GzAno/s
ka4puQaNM9QSgK7Ul6EOtje5rNSUFqtE+8QttsvT4C+pTBpl4fzkpPrlNgqOCkuPPxRBrIytOOGt
EahaEmFc2QbbcJlwD7u8XDHYJpOzJ7fjShtDPjhnBSG9JS71tCoZq312J+auHQZE/ps+2MCvaP9V
QgBg7Lnu89b5DCE0wqPoOiNN8vfMCxkoz5Q85+8bNKeuqJ5zO1YPhxackDPfjeTfRIsfIr6y5f8U
4kZAaq1CBY6LPH7w+P36YnhjJ2o+eQczVePYnPRyM+SdO1ZzZA3xH1XYao50Q3KpStXT9BC5CEir
tRf1Xb/63SaC3s8Ox1b6oQwI8USDrIXrKHd6tDphJS5mpSQDIx5U8I1PndTvs0pANe7yU1rK2bdS
5mbYodQdWdMXn2KCyRvs/eiWQO9icAFdPDkZcIlGXhA8Q2uhwJfKnEKq8niJHSZcVF/sWqYrnuPH
34ZPjhfYp772UfsXlbFAHyQLIFqlnrluMPhIzgwlLBU/+PuWElV9qBRTUZUM+C0vK+piKDM6WdMK
LHcUtN6wPL/CHCjMYSfOVB3J8TzHvT1Kvqe2aD7ueqaufttAXCMdLpmbusCuiA2ATscz/rROMh11
riDd/poZik5H9S4nLiklUkTrQNrzHYtV+9XtqaK7Q+TwZxmvqHiQLLE42G9v93oDWurRyU1IGtem
+rzW1LJFKgAsO89H7gZBMMPuiyEukQz81vYCzekqzUVcgVU9iSTn/IPFPvfEOClVQe7h4ezVkwx+
0oBjZkF46RZggcsyEx/6LMqSDPf+02xi6gKJP9Wh1bxtKtL4ZGD5n3lwqsyM8BpDoYYKpTxg9h1i
gxChLqGQiIpZMKOdLJ8fKp1K9qOTDxVPqMFjwge3hzh9NOXgYVqulPcygA5Dlx0RPlX/G/j+tXFw
n/OudT4HRH26luFISiDbdjP3HYsJccnm28Umnjbvs4KqzpkVHWSx3knMSAbcsyCV9+Jgy+QyPq+t
3/cIIeQ+ul+CR/BnlFpNeJlaRF6Mg/jINfV3zdHLiXXAKTUfRiFoQVd2i1NBPKNyrNM7BSPB+pdI
G2dVuV/1Kw+rrAtAjeR2ccC68Yg9nDq8u8Ezwx44GAncDCC+XHcOzrPsdQSoOt3cbCz1bQ4htOx6
WzRVVJchTTvQIZXF9XIMd1KBgJzD9D+9GZG1A3zqNSJCtsLizqYMl+QmLbPn2mMA4t+SjpJi4xi4
56IMI9oglJ8yvmiTuXskDXkZjC+vhXXrq3FMF+dwFYKN7XvfFqpyK0iOdYHNWl/9eUbqr7dluged
h+NlUqlV3bwiF6p/JPEDPaReeBIEMRizP6WkhC44rADJe4z4hK+Yg3lWPGluB3WkZ73a+LK9AnzG
m6azM5EyxGt8/F9Y2ziad6P+KzK+j3366j5GFBSvfhak9Uas5hU7T/veRAkh/ZXFSaQrI3sdccmA
ScwI4ZNzIo/8pmGYeNIp3CpD4B/nK0+XkoZc8GUiB00WkxRabtY9lBU6MBofEqXe7wR16+blGRYl
9mBTQA4T7qNeulo7SZLh2ZfKMKQd+zGbVNFFIh1QjxktFUVlUan7Bziluv71FcI5kBN2nyxmk6cq
nLqMQz8St6PRS+Bl2K8SJQOB1O52nyFMxWchH+aTF/iKfE0giLyL1/7Q4t9otwtK+Dh5iUfevPBt
IMo0oMLhOlQg8/64eMlH7S87KDjqLIpdxrmc7uYAIdexL1g7ceha+CrytKX7MaEsnitx2eVwyyPQ
xA+PuCVCP1AQ6aE9goiVBNi9IncS5X9Bg+p07DMaS8NFWaxEEgw/YdR5U+wsO8TeVOTq5be+sPOs
nxKtEiz54wL/aNB5YRwyYBGjJ67+fkT36m19tJ4Mr/ads/eTBMFZ6skIKJZFyiwCxnXGKAlT1jIH
sWIt7MA/+k46SP60m390XOl79sUhiZPoFhWNSeIWZ5yqJekzLi5ntwMkydeuT4awBp62b5ZTZARz
XqbmX4AwYkRWSiYlT8hmpAAjoiuR0zpZBDV1vTfg1dkroYBuR4uTpGGNlBEjo3yS8KBYr1gLnmxS
dXhBRe4WwZxIM42x55NALvc5iYXmC2XA/LRMCe3agpj8xNJzOtbC5fg1aA9mTy/Rja4OCYONmBHj
j4FWdFFA4xpUhW3YZ5826+euLKZSLV1I89laLN5LJ0PvmTwumgf/vSpMUtWgtHRAZPeObuyFMOv1
XaJ3CCUqd+yRo5VEGHYfbewOVCQqo4iE0zUh5p4hLAgyMPtYb6cj2oAVlZEgboM1qSZ8Hz4Nvv10
LN7QS/v/yLK8SlzfulB4+1zWddjYBFQV/G5ax56TrVBEg+P2F/if7u7uGZ7Uq9zLr8xBsyE3ILZP
14Ys4XVAsYBoWpDCojfpVTmk/AYhfMK8q1QEYXsoYFjXYc5mSCvwNz6U3ot5KIquiGICtD5NNcjZ
q8RjIEmXZOLOIPsydc1NR6u44zTCzOWGS9jNcxb5W6soXwxizpDw4vIYVLGRXfLI6bUGd1YzHzzv
qMRNn6XeNolOluyMpV6Lk1RZJRgWCv0bcOeDgeLmtLP+4RQLrt1CS1FHMNlyWZl2k6b7STVQYVDe
38GN/5jz8qzzm1hIcZmelHrv3Tf3ssnqenF9OwAYeVZpEtQAf+L9B6X7OLJvc5zr9UIfk2UDLfSt
RSdtnVpRCjETSRfclBzWC8sOGmP3BcmkVd4RqDBdv5C2H9YYmSulloGQPlqiX1LauH7Km6VT0EFI
c7llz6QaVWJ/om5IM+x2hkybULMlM3PvTV3Pne2+ZVPnJtT0NlQl4uEw3EIumHGa4+6otnVC6Rvx
O6d+BtcnSZx8JZMm/x4dTmZjDEE03uUB8Vnz9sxtn7tj7SEfqR8RjgmqobdlLAYM45ef4F4qmEbi
UooC0ZvNFTTvdIif50lY0v3TFXtSySh6Eei5wjacVKof/iD4lHr9OzOXuoxY3aVQrvNT/Juo08SN
5CUx/fDxDpEnAuxqR2Unu6U7Sqr8h24p5zBLMBuJiWJPBFgX7xMSTYu/GsksoTaDFvL03lxzP7F7
MEQmZ2YymjsLj+PozHA0fnH/mLIKh2v+kWO1QXYTEZGA4vDao3qtGF8rf8PGc7ccETKRAr7/MXN6
HD1cUAkAiwx5il50QleOxQG6Cxo6CiJANevIf0vExFp9M5TLbq8wzEaEaFauxxG1jnr5UI/wS52v
a3mEDKG2tJzfvHNRkE06A4yTJDhKzp3mEN7najd/4AsR7R+7I7QGB63mgNgy/A2iHoRqobgoiBxs
rZi1UrjErRf8fP6dDmwGg5kUYFVaVwM4PmtKKoOgQ/2lOHEOq50LY/TfSqddpSRX+Jft5XjxDb/X
0EbvJBYoK1T+zl/u0CTXMW9qRkvKkMlEZoe6P+vC3zdu8S28PDVEguLJzU3RNB+I7+butrcONZbD
luG5xkjs5t41bTPqjlYi0QV1uyutxZLYzMz10o/89g9CCvQtL9SNEBQvpPHt38PwAVRX4Jh3AmUt
oBhtbD41kt7g1tL+U4ttFzY9bHL3tEw9jlFp5dSwAsS07qu5Xx/BqjGfympzKHfHIEHFFX5G77OH
cjB83i7R8TAHG7q1Dmz+91VbHO7MXXZmAKaBgwLh3azY5/Z9MisIfPf/si5Y50QXBrRq84eNuThW
d5XEuIHfJlr8q5giCkAtCu/K1d1MnwnZB1awKUZwHMi/vZwKNNTnMdtqUoVIndhyVa+dxmCE83Dr
Q+L4AoOljc89leVWrTnPCoKsMfeK8RgG+Kkntkx9ke+qxMBgmYLsPRcyd6LzaRpCukzj0lMDQV4e
xs5MeiFu8Q7amGqPXDA+lCSZfERoLjcZs7uFFQWAN2WOnEDx1xoc0LrVJshVJR5QcwtwKP06801O
04VAMj9BCysg97jFn27MxtxaE62n3ItT/NbsrIxHiE7vHl9s+n7fFAcBlUM7KnzAaaPOUmr2Lz8f
AvWZkk6G5cBFYunKTZSFFzWP2deI5mGJWKvZUOYJ6d41Ursitz5WjmFhyVcNco3gQUY4oXy4ciVJ
Zd+wiqBbpCdu8Rj4EVVUQW7a24owUJ58LuXg6ie9jCwSXR8/rEsgWDJTsMHZ4wLH56hfvusxSXlJ
mN9QeO44iOP7MbVDUdkGtv7hBfho3oQMNSPadyaSnokhcBxW6uZtx6g2ejnjbPN8nenDrye5sWf/
GPeD7qrGIDhiXV7odmFNR9mP+8ExMHezVtTrZBUml1ELhnroNLHoFrtfmuuNNigRYLJwb96yRpPX
HTcPs6370TNUjlQ8MvbneJ5gr4ryhA5j17CXRyYtuGL02+XxLg76yB5Cexhk7fNUb1AsvNROm8a8
sFTO3P+BUj5bM+aB2gmWfwUozSe7r+9LmWX49c885T9OO7loDWdfGdCdkFuoyyaWU1Q8UTwy9/nQ
kOIH3WM+RyDBysVoB96EMfQsz/0cWDPzGy1FHjOcIHiTkcQWqC6hRk1AcDb8yqjDDLnwys/E+eSK
T6pp4+6aH0nO5FxlhysCANLsDwIgQ0rX3lwSqfJZJTwfC1hmcmUYR6VkCUjbsFVR4yZsoeBbeaNt
/2hgJAp120MgFHDrauTRGzj+EDAMZOOA95PTDt85yOIkL6k8sK308sB1ghevmTU5XeHkXte6FaSO
t7hCc1nGpIDiL/nnx3LKADwAIfnT6wOy8VRJBPwZNkvlPYMqB9BkV1XqIovZMODKSx8ucMrkZ1EU
YmvW1OIBaIwik/7S0mgtnQJXp0PieJYNN8cxtawjYYYy7ASH7VjBx0IlXznMhsoLx05k0Reiwgzm
+kmhs6tsao/bNhplbAcv4aJTXAGIGCEEMCwJyMsE+YA9Of1KxJK4MdKI7Mj3BUqfFg5cSAYYztQ5
koOB/18tQvnyIcuOC1nGwvmemwP8G7pIjO8RTgvqOOz+TzTKLB1eSWGI86DyUjGFI4dMDVsua4wN
YvG8mjeu5zmVD0o5kCDxskPvbA2ZdEoFqUDN0WtVVzU1U0v9irPu500GEbyuKXmVYVSzXwxAI/8b
L/bmgZ5IwbCErPigEfswl98ePWmbmmNwNORfGuFV7Bac0QX0vEVi/hc34l+BhqSHyYO7JPi/pngl
doyOXDRGTwcfTseOmNl1t64lEscm1LYaE6P2F/Ogv3rVUrdK8tgv/NicTJ6/9q3nmlwaB8hhn/Mc
TpZSKiEYQEvTDIKPiOrg5XkYiOXXIPhanzAjQVcImCZ3tI/4tL8aSXD9HBtVq/0rfhGdMsCHqZfT
EQYZhNfm12r++CJ9b8kMOKhGawb73VGDnMLUm4xdZKTSjRFeh88QL9uPHF/nyw8oBfC5c2QQQTy8
oRe9zHpaaTIjDsWayXuPPbfGxRRazBHI7Z/7PyjuJd1fA7wg7HMNmWB1Wai2vSRJCq4aGr2zRtU1
X7yLj7POEEuP7/91WsbtGAGzxKGroxKxHRLelEM+oOuRzySgqxglKpHHYfgSBsKqkseQQvyfQ1p6
b9yetIkPO7TeqUdDlJmbm4VspqLBFTOpt8TyJeVDPZYYHifJ13Hr7MjPAWuxUYtzZKRe1ubNY6O5
x2vaQ3Ql+5G9rIt/NgcFTj+vDb3BN9jc0YWnMN9jO6Uuq+7P24BEQj5Irzx1jzlgCqxDNorIzPNT
/nlSqNlgZrg+SURIDrIHcGXfLbHk2EgBTdKO8Lw5QnSgGYJwZZTLODVrqGa2v9LHfKzNazB8ZaOe
pqYEV7yVecfadTkOWJMZkTKzYd4BSBOKgjZ1oTPy8V8XxAjDIn9avtlOWjOMwbB7L7JzdLZ7s5lF
9AjRRlFlpHD5+C1QwE7j5aM+yzmy3aCe/fIjwRLzyrIHdLhmW8FhFMIa20qaJXDwRz8CriNukVBP
4whHJyl6r1vnwV+BNmzRECs3aIgtZtUGhXpy2Nio1CzvWLctvDR8wo21oPsLNb5odUCraazjoevO
LcmsX3tmXKJH2Xso8oJQOCslbUKYdQylNQIYmzdT0gbjcLeQ8axBmX30S3kPu7/ZN1c8zPwmdGqR
0s7NOFrffDVnCbdxTBfIzA1XRDLxwDLCPz16N3zTDnW3PCT1wrXJzGotqC/WZhYTqtxzky6h/THZ
+5HhAzLicTbp/Y9JDhiCw8Rjyl/PGGwECRaAHQwhdcr7gXzrSTDSNHrtFmMxxd7Sk3vkP4dPnI1Y
KV/OCNR1Z0khSPCeR88aE74cwq3DpjemZ4fP9xWhcLEMLNmk8yBi5ND4YyKUFAF/961tzMFBY8FC
/zSCyX9jIiKOZJ9AyqYrwXw39zRqvKi6rxdA12g1+ym2UQPT8mLxqeLKp+deV6BJiC3zT12L00uf
sR56wM/WtK3gBUFcpFXKEcMsibIKzqn49RDe2En8IDyvQzsDVT0Sna5PGGCC7quiTuJNomMCC+SA
oBmVwFAOXDOmNlruDdXW72FnGcDHl976hcDFejN6I0bmut3FY+foSVUIwLq0b7V4N+6rPXTD1TuQ
F/z2KvVQgZsZQS+58hTVZfY1WAna/p0LNiAHGyYltbVDANGYdC3GIM8mb80iELwoHrTBf+PX+pkd
OzL59qG8YsEbRchHm6ecy+sVv2qEoQEa2Uy6WNxxiUTdl0+UCiwJ0fnlTn53/EghVPp9sW0b9JXh
iUE9fbE1R1HsUbd4Zh8FVKO79N8wfqKRmYQ7k8QUUpEr1Umk6BCZk4jX83bHO60U+uejrmFSQnbn
RDY4SvnzeIHfoXJW9BT/2Mh2AAIM2sQFggL+DnDeFgImETxgfHrqbdPUx5YLI938KIDYEoStIdIQ
DgOnsgF+sp04US1jXHOa4gy5Q1hZzys3es3vcVrZ7LV5xAEd/B3VkdB9fyeJ4ApgSw0c80Tc3BPR
OKMS2UOc6gwb6Cqmaq+WdSoN0TQm2wDgyBVfsvZ4Kz7wq5Ii/W+rpFngF+EEz3eb0jpXbMeTKyX3
/MpV4jAgTE1we/H5CXkVoZoSuu4JBcxa4Orhq6ldzyJsMqNjrdpxKx90TioxKL6c9XNFiIVCYJ9B
0Uub0uxX2tHpmSX7AEj7MEbx3SJ0ctdyAITRQpIxDSR+VkRsm/FSwVHbu9PtaFbJhjREFJA6mbQ0
7hPnleCZwW7O3LWmBf8Zmjc3vqDL8WG/s04VSYa6+IXVjAojCDMMWH5Qs4uV1+99kElSHCM+t0O+
w8NQNI8PdScXCVa4CBDPQhWigGrVZ/MKQvi9LzEHLZzgXPNbj7s+M2lvcV0hXRk4jNY+hoE2AKXc
k+dTwOzlCddLCnkg7T5bmTFVaXEvhJo7PnAJzrDiVt9E3uYPkBhRvmY65fSNzyFJ4dhk24heQGCD
aqLFSeF+xG2je+QyHKB0gAEuFv1Bg6/ZCNi4ruqzHQvx47Ii3CeCpqb3BE88uvyrr1m+AC2qgQZs
lWC4m4GBw7UlDo+d7Y6h2uuS6oN+8ADwOa7ekOtPOUlyC3o3B7iGReNlKbjY4eALBTGl/6wiaVZJ
dJVU7SAKzmjzj6LUl8biA23MWhEs525d+L0T5ixuR+PCSfDkDOeVNB5YmmpbFdL2sKwjkSrC/Ta0
xF6jVOZckD87FIJKn363OzL6UckkN96CA4x2W4l8i0KJUdgWvL14AB7d5SD5gERxiZ/zWVVzdLgF
+KeFt6sAu08dWHi5agDQ5sihxWULICe7/RrXYK5HXOWDz9RlbLSkIkn3/ueITYah5G9S3cS5+ZLf
1tWdSEnYjZCqUS+/DJNsmwOX3JxiHV9U9NedA2BTlmZcaqkE4Mj3mfuYCbycpeoCijw4wxcUBE6o
IP70JwUg72UToqvWwMpg2M2kzVdfRnER8E89RnY5Mqq9JQwwaGrz9xBO1Fg/L1aak8np5QqW9VhH
tg7FPBZAyu3vUl4jCBT4ARdnYAr6BGyeRx37wf8deHY7anNRiwc92FKCatKanzCctW3Gu2ZOpD9I
nRA4v63/J+1E8M2DVI+3DDZr621HR04oOUvml//Exq7gEH8l4sJDYQPF0hMFggc3EwMlrYtNOTn4
hEkT6FcM3nnaRIvuzyWtMc5o+1jWmLOTTgSn5x5tLbbHpcWjZ/YEuy72oyr6sisQ1e/cF2hPC9GD
PL3v3j7OuzSjL1goEfiUWB4UgcVJ9YMhIjcIHt9S62yWbqREn6EqE5Ib5wjkkWZDQ7mwRbGqGs3+
JcpEhN1Emy8Fz1txWdjcfg1pDMfCdnjDOCMjDCt0Q+ts2cSEeSm3QiFrq2torNfxQdoU01ZY/mb8
22EduVggDdLhrmEIoWuwDD4oCg1p/KG52B2/yO7zsSahspt5S3GgDvr4Z5GGLaU7w/wi23NOTn4o
jy9x/8qReQsBA3evzcqsf2Jx/LFm8jb0wiMsL9vAaeL8qtIvDjEbNmP6dD8o5zKElDY/AUCW/1ie
m+7kK+owoJSknEfx6VQmkoBpl/UPUhY6QCV9o92MR9iNc/rM2XROKaEf5KXjpZ6CqSccCA44XfKX
slweicZxGX8ypVcRASb2nMpFAcwIdyZKcuJxNfKnSCQ5x5s5ZKAWdM1H/ds9cy6TIVvvakhIC7I5
lq51lrBzIrBgSdpeSmtRfuHknyyjba/yHazlevHtDKxaPhdvVL+SYma1t2ZWREPOAMlHeJ1jSWH9
6w1HCDqbGrOtDahKFhSenObcaIdFXAUW5cLy5S/nHSZwEGrn0K9JjkTnw/YJaI+NeuYXSwfjvbWT
+GRyDfniBC/PN0+/jhM2a/doFaRPB/9y3TXhepB3SAby65qioTtqL5lDV2LxlX56H+5d0XMJqqb2
FISB/NlqeWInEc0uJxdyOLtmJepMkadiukHvZ7YfjdErB15t/aK+JtPuie5k3sFDsYFh+HmthsWe
kKtlViYKlu3+DTr4WAjbdsKWLe/53c6RAy7Xr/ctMXHUvjDJmzjxSqPCJjhzMyPetSf540A6peOF
nPDktnQnj5TuOfTXEbcACzCbr3BAjC5IYjzPEoP201reyK3EcL4y2P1ZdkF7E8rapulfw2h7bVBG
H2PYmEgILaJFt83NR4avqXBc3evDljrEO42eVpH2mfFOz0Iq4CVBYrhmz3CNFsGP4uJwhM+w158T
a+3OmURO0I13Tn2Q5hwnbr4aN+5mu0JcEza6u2GtnyeRBUNMHPB/dKtsFixEHs8EibBYRJrEumvv
pBVlvLxoJZU6/2n2UaTyDaoAK9UE1kRgYDS1PPJa8S6NFhUWp7+MIgBfsuuHuURuVbPSSFNYGLna
e1gZrA0zQc1Rg9irJbM5ObXuwSIom2uQRif2UGrATzrwaxfhDATy3YBYU6adfp3ZejT1oIGGO7c6
UTl3H0JfbLZXOFsdExmvmbbiVI5tic+SV6EAWfpngTHZO8fcIdyP2bxqk90uu7yaZVcEjo54MQRL
VFJA62AQbZ0mRv5QumJfL4fbn17SPMnBbJaQJmxJ/ec3oG8IMpUE3Uq8L7l+8YLTiKUWOpPpkX5L
vx6SoW4YbiN+FrU45cJIHFJYCxZ0ZR5On/+T60dbvom7Npv+hXbDl/UkuZ/yeQ+llWUe46v7q2Vl
kb+8J14FsC/BWCZaQJKrWiGBJqy/pqAFTdDQ8E14tbsS4GDFbuXxibFROuRAaSVdVpjkx6QA9aex
E0cnyvj+uCRSi6/cCq3w2JwodqzZ6p/8M9Okgk62IUEtSGgBT2BGrt5q6o/wiQI8OZQyZk3KqsVG
sbD53jt38osnj2iPCwftMJSXxw4JfvQEzc0POLKs0AKibGc8cGJSbM1J5EUxwviVxStvHkAbC+4M
f9L1vt5KYyyg7CpXDSQ7jfIV254bnY8mZALaud5GHx8nJkcsiU4c1kHdE13fguxirMJZ4Vv7y6sZ
b8nTB5ob3EI+iHXBpgnNsjXE8LTk2wMVjFPoLaAGCh1iBItAlQjS1Ti4PPF9AG4rYn90uBD8I6Kp
Mg4qVjJGMq7vHa1WwS3iFgzXzILvTkZDMoyUjwE1YBMpFqmQFmiNlbSUmsW5v7OPemWwi2stPM0V
UtMZDynj/aZ8bOYEzEis4iDDoYCSmy88CDmbWYKDT++9zNfQgXLJyKy0/er3JG5+OAJ9Ezx2T9Ta
EgL+CesE/crCua+je+7Ko/hNt+W6sEsmGOqyB4KTfN4Jt4TD4BSjneIwJp/8bhECV8s79rASIUnQ
Al5d/8/hyh+0CCBMjocDfooI7AB3jpMeY5lO9wxabVJ4HwPyT96JB4L8j1pPN5wbAHDaC5xRxLoQ
09g8AW0jH+gn4X4UoAF21AWa1Ej4LO6bE6T2x3xkhik4LD+JCTz2rmIej6Q8Xm+1InDWx33+sm87
t6V3kraUI+JScs9hoit3VVcLpLbFadZR4pz5wz+4t0xuzrIvbUm3eYm2baqQAZ52RA2rtAnldNxQ
4FeqHvKKKDcHJItvOnyZstKySOouGNZTjgAmggGmtf0L+OIA6e7yBic7JUk0jg8za768f14exLkj
Q2BcA1Bs/vtlN886/TT4+QksZzqrNpeykaHaTzppcK1erVICJoUlCywAp3y0c0WueVIZ/72nYk5A
q8EEKH+EeVmVLZABt8qg67ooKqY3FrCWvC5a9fNI14c9J+nVKOL1U1KySI1iVSb3/MgXC+sl6Cvj
UDrXkR5RR84V/zQjsNaY3pIx4UnF+b286v7LrqsZ6y1vMfNte6iN4iFOA+8pydcixj0GQ2pCOhwE
fQ54W/CkUPaPPUYQmU9SJpeOrUMEshGRUsa2ITpwXelxIUb0UTfIvsAeWUyScwhkZJRBZotSt2kS
NHG1GUBFbI35EiRQDzlIzCfrszAxblAAQjXDRkApBbCNZTgsaWYM+khFMthkt2AAejt3oinYHw7G
bBQLxL3VZr6B2h9b+M/zd0GaenpOunymAFR/0i31AOalo/8azpLLgGNQ99MgdrOhOZWdmeMI+mBF
EcSFIjxsE8Scq6f0FhGitthsJNtVPf/M9hTFTHE7XdDTW/4LKFhj5WRT4fpQJMPSeo4uQTZyyxeT
PwK+prkrGFot263Uaw1ljA6Rz8uc+KazAOlyikn4lTNrq4a7lIS26kKbg+kMLDFIkhAmQMb5Zsnt
DSxokNHY4Dwvn5/7di5vLsHleY50ICo+YS44j1sPMSbi9g0M4PSjnVx1+9A4o4Vy/qW8FFC53x6B
uDW8FSWnJgiITN62K/C3WNo74Ip4lAoUlRMa62xpAsiscw8VlvehI5RoocFvhyafRs3YcmIvoxF5
Jg/vvANyJ9q1fRowvlxqM2HhabmKX+cxXGEK1+yZOlDpaxKvrzMOaXknYA3fYUbsGcO8nikU75Ze
F0dG+IxcxhaZTEGZHC0p+ZUvdwGaPg+q4VqMiv7ZkO6rPEQUU86tPPuFDyF98Bk+W1WNi3qH+gqN
keLH4MZtlcwHBl8XFwYjf0vO0hCfTzo5r2R4xOYZpgU4OK8xS15ggY/rX51wRSMi9mjCdf3HMNE8
mDLVg0aVkL/wTskG190Pjb//fMoCafCb8oOIzWPkntcH1CoXNOd9py7zKSh3K4+Z8v332gcocDY7
nmYcVvvtvzOTljfylfenwnDZS91SVukaoD3n+QjvKmNFLPBvvAJ5sc11MuFaLp9G0f3IncS8jDR4
EpD3tNfwJb9Yz5GfKoQAeQEvrRbPFYvN/KANAu08h77AC7zQuyUm8aMt5diT3Oq5NG/iVsW5kVqg
6GA/JGL1LkF1lAiMS0wX9cnAC0fuDons3fNpqOuXN4GLpMIBxxX/wiT7dvoki/OX3bisE2MA0Lfs
t+bEtA4DeK2o5ouBMtQbefOElUgpI1LDOoAT7uM5BC+SF3wgaO4p+aq/TcA4nPFvESXDhUCqIv1v
2A8BnCEMGpDXlW35RZUjAtOr1w3XrPwEPaS7a7FS0TZQNG8KfVbcbEQ4PY6JDMAgrFjSxPo2+apC
4z1j7G/Y+MbClfkUMddbgTUCko1lcONXqrNxcE1EV4BYrhyMVHNJSOynIAhVpjc6JCZcIKXpp9Ly
h0F++oD/jwVP0pmyYc/bKnIFsZEhE00M3xcKfXPqLonU+khRYP0bdvgSGXWuQkPwNvHoNQ5YYQ5D
XECNmqJJj2JuaaFUhFr92c7UkZqBGYOjPSYswUxxDcpGt9bqYuBWoVGR0b+TjmlSmdBsDg+AXJT2
ZUHEOZIo97b2dA91mw++aOnRlT9h8KD2rpsLevYEf3Ei6lVh85z6C3KvjLZyQsUY9Igrn7U5WRzF
aV4cENYzeGKmtEkOFB5UgPQ7tv6asU5s3jd5/iNO3uQxIz9oO4b2Ug43YeYaj9SjVA+BVLQMEPpE
VBUfIxy5k3Vju2KauOAFEmicmadr1TpSrKa6WHc/4+Ky1Gsz7MtrakGbTsal7c7N0tIq21meP25O
VlGIdFXk/E0bA8V5s1cfplpriiJvY8REVaISXrl4IzbIpUuTSfFTHo9eJCNvAfPy1ceVMoZkhw3E
Uyu+TrlLpSRscLA29+CeqFU7kXl+oJv3SqRufKpVDsmGQwCXEyvW1D2EVSnDEXDEtwus0dDx3D1V
vOEucLla+HdLMozBAq+Bd1rQ1HpEJ4AXs8yJthgoa8sZ4xpMexWa4YAN65Zc8y+PlL4IW/P5bC7V
8NojlzH053L6aBv3WF5MYXmlrXVCAlhp3q/eKwr32L9jYs0tff4yR0WoPNK462kLSj65iZjrZl2Q
xoNCDsrO8xUTw3pdcaTNYYY5YgV8iTkwOLf3+19nbmzXBQuCfC2qxs5zF/7DSd8+lb1cX7uHg2im
o9vCkunbPR5OLMwW4lIljFr08JYGYRJhrAXhRlH4pQZJ60ezpgPEU9XxqlNvvytQKIF7lT8/y/5y
AOB7UCER3Whk1bDLdx1FxFbO4ev3ZecFPw9IVXaZ/+r0gsPGIHfUONWDcCI4IOZYpl3em0y2o4YF
hF+4YZyUUs8SnRdj2jhHGH8FswvbmqTprsRtP1PkZ+Pri95CHJfiuMWsgR0QOrnCGi4h8edSskCA
EJRoCjOHYsYsAio+Q5WSHw8s5+bPdZwJRLKOvyvSCCzz8i5tgE7xIH7J6ojZAddGhx/OLnrA5QxD
2Gf/aF7/NGycssbV/fab5ISQe1U+kbSaC78RAWTOXyyfNBkpeCaeE0fqJNrN6hXya14awmqRxeXn
d6vd/hK2DP+YhtKjxKzQPmMQn9pO5EHGN7IOyrY1FGA/4lTOymt8FKqWY0dw8sovisYaxzaGLJGO
bE0zUCaf87vk7mjYqH+F9RQ/95vjyrJitguQlmTfsECc6IYKiYajNjiSXdurbtbDWKXl1uAbbb07
M72sMl2byEGtVrnmSY29B6IkwvSmnvEwK5+Dn3lSQk9MjLlkgTkKguvz+89asA7TpxCMCVtLojxX
siC1PrBw0sFkdRl8hrjJP3KlZCyGiX2toQLA6BDm3S3j1aMk3XGXZIpo2lMgx5fHSImOkAhCWGZN
HwsKGvJ2Pt1F1xzZ9sPVXxnq4n/77rTkTRErX87SRjkSSXDdDoQ/fldEgoyKe1v8HKo3OXX/hR2A
hnX2ZX5WZahsvYQkYe0tZAYdle5X9gFfDO/xUE+OybwEbDrl4MJHiNFin/0EQ5GaFxl0l9G5OcR2
DZbwKAM8xlOXE+SO5NCZGL7CAqGKVp6Hir4jq5/ydru9CXGblT4VW9gnwUwONplkt8Y790jXB2K3
4QjbqRB/wjN64SVvIRDnkk2Mg7DIgf8c8sE5t+HkDLbgenVLASB6N7avAcopx6CwKRghu3ulz7Ll
nGLzmr45Qu/0QThy3B2sviyZY104Umh9cmjuWW880x9LCwWe/4zXHHZJfL9ccBr8lHlKRiQG7d52
HgaidneJtZDR1Ud3v/wNjem8DxBsKjwlYD0cVj+RrM2f3keaz2FZjEMrbC4LyCS/d61nEq+lfuTn
NYpOY93CkxXb7woIs37nl6eeMty/5n/jCLfLCQYzN0wAszEWlZxt/JA/PdRnrEbLIJ9jBo6ctQWr
ZGFc88+9hw5rGvvqtpvEQO4fT1wnZfzL8R0iJ9r244mqw1wR/TZRG2jYRstyzLqimrdUzjSGAEyH
zPXTY97J/mpSxgm8cPz+vli7QMkdv//TaXtVZZvABngHitMbIePmUkectbmGufy7IXTR6pvhvt+r
6zkuslpraMhJogYMARQnpJ02uGnSuy0rV8XPK91e74M/pOwJSSNYwHcepANyJwwUQROa8k4QyLre
2GE4FTkzO191lXYlIyPm5WGu9bqtf7tlyohhoGioKz+rD43NtJP93S6PBgYkYCb19lJV2npkUsJo
9fTGGUoOmV13DO6CnXmZRnzoeosk24FyTciubMlhX18JMlWMZC79XBcoASYHUX7hiOq8BP5EPPk0
C1Ff/nGZFb1/GbVPP8S5jyONNMCadsHpZo6xcEp+CseqUW1oEo1cbwJje5gsLnFcb0N1ensE/xG8
qr7vyfNFmUUcWzOQmJrHskgHKt2iH9OLrwPbTPko5JvwbQ0HqzZCampTVtB5ae78liZaCVAzuNnC
JzIt/Rw/ZSs95h27eKbfus5a3ineKagGI4O1f9ebRRERs1+l64guOQNptexAIsuoDjAld+K01rvS
lAfU1wQbINODZXM4EgbbJVykXCn8l514U5rx9SsLLmv0TsTTV4JxaCy3ZFGLfTsatglBrdawkoqQ
oT1+5FMdUynVQcaAn4GqCU3/Ved8LkVQZ3SIVcOdEGsXjiC/1XQNFVJm/5Wnn1V0IvEsLI8xwivq
MoKJF8pF48cSK/1mVo4tvph9lsJfMIVUi+d/ZP+uHUiiVeNIz2e+vBCTQRYE+EmgdBC2CZLuvItQ
7g4RoRb66/LkXXamQaVh36pafTAKS3khtFqK4vOTzg0HEHhVjOdLEXXrDpxnS6u8rGtuxKsiQHsg
JU23ENWE7eX7q0HYlo0qwtDpRc9ZpmLSWR2tNfTHkKgfGQ9f+Ft16jMEmmk2gaxL+BzMLQZbg2Kx
HONjNIJLUYdIHtC5QKePgVg7eBsos7s/0YopludOvgoW6lgtTMVYeWCwpnB6fijyL2dtqFj20Oyr
XLztC6oKf4UN2BgH6MxGiLp6d4ObjAXIUUjh8rkLyfhQT7XK2NBsTMw8SzzcOtSEO7VWeBcAPA85
45Rdl6zrvPYEZvtwuuUHNwO3kWJL6BIE+/lv/5TVBlbqxYrysk/dG9MViZd0xDnI+SD+POkN0V3I
GQBG/ZDbIQudxAbj/EdL8Pj7SsI5hu8RRzTIC3tlWkm5o58DY2ps0/UAyPY0sQ4kCQ92yIz2X3kW
e/47RIz4F2hdUJ9Ma4ihrF+3RkK+F1KrO095ZiAdYlWOsEgj1zmkwns5yBdbYwCWSbZjQJYpL+Fr
E7pw6hYHh+U2EVYDq5UamyuSS5bWtb8gBHCg4BVLAjBV0Y+hq0VOiv5kHmYBuT2ROo/JIkKBHctW
JYbmC57bjWxDBm0nM8qn0iMIDdUGmQDaRzeWld9ZuFrcQcW+cERzWn+8IIrSScwCKzGGko4F65Q3
0A92BpsO9AjEdptaYemIJ6+NC9EwvqtzPUyhEBxJvHxKvM9SJMHe2HF6npL/UPg2eKwVeCUj5UX+
nJECIOT+0oix3TOqYnGn1E4rUh32cqZ1iSeE6+AeXZPD6KRQa9WXxGlNmpgT/5dtPlCehEA6eVA/
4erheYTI5s5FyKHVQu2d0dRRgTpjeLlxnI/08Pf84jRO8L+V9TbOROrsEJGCACqyo+JjkksfHsdA
UzoBWvgD0vOufJqXN/YN+8yUh9S8pSG0k2ZDzrEW6gXwNw6oWyopi7e6casNydrIWOOPDVjFUlCY
IbzgZAgTzxkZybeyAx22LFP6UchLwP7cZkqx/zEMi8fBqg78occnYkG/A4VGufdiEtwNhh0bL7KO
MimT2eTsMrG/t3idm7mZ7/PESRrKyPXBmc741OK3Yi5Ul6PLV+bWHon/4toAQAz0yI69aAPp8NuG
P3Lfj7ObQWvCKxHRYDcDFoJYJkeGCPQaoemorjR/kNZ/NB5BMg8G7PXhDH7G9uKwd5wgQ29A7qWe
Zsg3LUHv2CW6O/qMeHGvT4LkJhNaDn4TJ2Uk6dFQ23/ED1TKWj77fDECA/gJrWMCznw7prbIIDLP
pXdN3SUgkUALBhiuRi8kNVzJl3JWAdhBTTuxZNCoZXae2Sb9ZWTmX1juE1kDbfAs+ls9+6NQY26g
pqmVbdZAISsXxeL8SdcH77gieVy9Ni0BU6EvYEh//0dPrbHRGKq7R/ugQTk8Q5ZIr/Ld43N595fT
tYV/9HW59D4HnK1CDqutwEIKX/fuLaKjqgQ3PAALcARuh/gbxAJgsZljOa/JrJhdYJW6ehfLj+OU
QdhWdh/rN+AXGRlVsWatTPmOrg5PFsER1Nk4/rJyPorfT9OprxSoGuro0DdbGkShl0Kp2+4oRP9I
/mDlwN7dfd1voQ7OyfKL54W9gOkFZnMgmBs3Nkry205L2f7QZpKD2CrgfQLvVQQ0+5Z/wDBVXz+O
/T76uGZslczLKZGPQ6aMkvxDZQw+KVI/HQnDTcj6RU9YEicCrRbdQtjUO0JRhdJnGSal4APYhVFd
GGm07bQm12No6kqyI6jVuI/i53HUN5qfo428JzVa7wRM8kXf7haunSHWwORA+ZEVKB9auhkSBB1z
iIDTcrRW9YN1QRPvzlApFm347BXx62jjmJ0Lp1jvrlw0qOv4/EYRcBnOD3P5/KAA6ZBkhF22TWtC
cXPe8gOyusRoUBS3hRUoWNhoMGUyoFA8/rpGk9LoPV5QFuLCQmGnt/Q7GBZYVMDwCjQMZel7VsO6
pNt3kOHzcV7RtSTqzYAuAECko6jzHR1GJFeLBUqx+JrH9+3uCa8BpuHuUa/9z9btyJTHSVHyVYxH
teFWqBrbaUCLlQ+j/v7MgRB25Hu7LVzjoQlNNJh/gU91a05hiOwAxGERdW7VVu76BXUd5r7DBFHl
3QBVYwTSg23ZsM9DydpCsz4CXMUtMOUlDd68aKXST/AbCy2LMD4xhq4c2KndbC5BPdMp+e7uJXqT
HYLG2gv+RxvyN8lhkliO8UC7ogCluQn5Tbl6QwqVHMqN0onVWSe2ihL8lEopqY04/ZSZ6a7RwUBE
ilhh69YWNWl8tt3EBv+uGd28Xn5+0AXJ7iog4nJCni9LfqHyIPCTPj8JQHuDIPSk7+p0/p5Xekjs
bl/oPfVE5MV1QUXPuy97eyUY0yds71B94Z6ZvR9GCZYmck0/6btub9nYHvpGGeKpk+ugR2JXtf1x
vdRGg1u6qCIEBh55sclyeH5ALZVgSa4npzFPcQOo+hHBTgt2hQ49zCiuM4JI9nFMHS7GLFrRcLCw
GGCxv6ETKrXzI3tYo1f4kQdAxjkmkjY5WENeqRwemqtLaG8r9y5sQ4Ik7eIZ0HiWER1W5lxmlOJK
GAa1srBaNbD/w6tnha6mDmP+5ZkjyaRUwBsILAWUO7UmwYY8kZOA7Y7bLdcWLSSbIcksmh3DYgqy
y000/oQQgelqpqkpeRY2rzRO+F1oAPZTpJb2T0s0F2daiLZBQD+eYhtLA0VyM+pW07rkYJUfw3+Q
x+DVUTohHS+skDxjH2KwN+mgMGBZ/EO8jeRDD+sXKF0SJFm0+o26vu2ddsvX4g5lM1jX+PBcGwd6
F1AOsVYowdtFbSy7NvG5SOiWLX/baJa+yxLXXBZKDdtrnj02dxFoZ9y7wvrdfPpU0iRirC+y9usB
c/LntD/Rxpe5L0XO5QTT8JxWEvKx6oSHuSPhJb/1JIn5rsjueGALDoPPt+heDG0GL8C8A/cstrVW
FkCaBlohkjPnBGb4hAkcxO87Ih98pqJvuYi5MgEZZHg0JP1jS0TW4hk7juSrFQ64LFhnQGBtQuBT
sA5PFGouDLw87Fd4J/NxcyeoAavdO2vtU7nDlwD8PNni9sSfY1mpTStg4JOeZHCwQh9YOb9+Gu5o
LrkloHaTbVH+DIr7k5UNbvu5YQ4K6Lj2LMESRxL2Q5NM2La1c4uypkekcEgKMDFnfeiVH3VDnaNZ
m1wiFlTn7HmtAYSknsBBYgw/fRI2c87rrXqEp5V6k3cbQdTk9BoB7aVmaP9Wssnmpc0S8n2GuQPo
EiRVTZzuFz5ufPG7k7yh4pkPGlF+KrPPfNdifIZbeXtPCCkqO+q2kHnT5jkprkTan+mGe+1cgqmj
I26Z6kw5Fzgih0DrL6hSTO9+a6R/z+09mUjv3+jgw2v+h2S0AaGdEWi16Q3nMLPSXnSITC/FVY6s
SZtedvLUEFtkS+8x4ITBF+V9tEfgiB4dtcw0nGqOr27oudwqiJPKglceADxbF3xzzeo8uIYvVeNi
T/maCVVok9suXCNTsv1VFfkznW1RJUd1ieS+jUKoH6cQPqkYNHTOALwFB+V6kdEtVi2Fldg5g7Qc
WixgZQafvqSTxW1Wql2grxR5m4y8INX9ibKfsQf1Pw5tWexG3279iYQYnIOaDg0OepHTFeiDqD22
ogGqK7ZL+SWUi/zrpUdytTuV/DwPXFPSV25nPFD9JoL23Ry6JsKZu7aJJ4tlWLdE/km/YrJN7V4H
zTtUJt+58qJTpxQVTPM5HycEubEczWko+sSvZBTv950Ybs6Oowv0z87RnnVYq7Y0cLPP5GH80mJ5
EGyZhvcEbrKopH0ylQvMJAE7T023f8eoHsoLbsKJNf1tUX4sInqvmK07lAFc+d3azKARRaKiQTdQ
kVb0gVrkg4ogHHRfveDCYGae4EmggqXnLpzp3calgyMeQ3ZLOIxXTyTTQe+hTGVm8A3hh0ma40De
hKggf4S+zNUSJEOK/5qHEvlnCGrUvGXQejy4KrQqfqDLQDo62R/x0mc+gJaZoVMUX46srHfwA9R/
yTrAtKBzwAzXTG3uSVOkE6IG3bYdc/PNXKfrzc7CLs3OzTVy5Mk8KAQdy97hlmFv19Y5UA+jIE34
WBw9hvbF9fby3OimtDeUm7gj6i5IKC0VeYLGZL3D5RvGbOnjfdXP0qYqLzXPz9joW2OfEV8LrI9A
lh1bn62gwlEVLPiOCEVw7l5BIPSGLcXvsbIBkO+tk3JFd6Whpe5T+UmjVvwgLqlVRXCl5IlEZGwk
z1KI0CE1Xbl45rAttIxZLDIUgZWWdmpnmj1jZcx1rJ4bmC5v8Xe0UIrPdrjA9Sdxttxn3enMxbH+
xCqIPhY2LVnpMasUdPkpL0nYtb+kpBXQMGlylKct2hDTfvpKx9InnCV1lH5WZWlKyTX2YWlt4WUv
f9UsVq+6DknQxthcqDCn9w8RiQlT2ZzgBERnQu8C+K8HC3mtnsk2c+eMkz0Znr8tn51gbcvzoQoy
3KwTy8pPmqqi4eRP3PkwjN4Uh+Yq23gy1m1LHD/SxDSbBW7VIHfTEzD5pin84CpPrlYi14J6bAPv
kaFu4mWBogQT7Bd9DZeCaWsqXAZZ+UB0aLagnmu/u54XLhexTFMm6zaDipT/1OYm9/SxS0fpGZpd
QrMUPgul1WOJxi30SDiO9vSzBlRSLoIifw10pYNg9c2CSRa75EHJ0tlRFl/lQkh9+aQ0ZWgSEtvA
qhlK9dbXK8kYaWlzCdDkiyDQN6tMb+WAGryX9tFyhLKDLusEug0sqYcB3/CjelXx1x3Pxr1ihBw0
yPR3InWOL8nEOtEhJxuDQPN3dgwCkXBrqxYXDnQZdLEnpAkLISDMjAJWVUEiaa+cTjMg8DRzC0cl
UDHSAXdff2BF3EoNAO6XezDmdVbF6S7hLdV7a749qkggXmqliDhLGBZNEzZ5VNnv+YlWSYgVYrXz
Mtb5JhMPy+uhpRQJyAVSN8T/J+OhB1smmtPuQd5dImG6g8R3jK6qbeclN+ySPKb1BH/vQbwt3+vT
zMmqG8mDdcAoIS+/t9Gi7yQ1ehBdlbVj9oCEgtna/wnPnulKoFiTlwFwNQNp7HT6mVj+esQ9mRzD
DMS+ydYkBvCskxnjMHnLjRFVGuS0VQOXwsQ4KeXt+HnrF5Sbe2j2Da4e1n9kz1EIt7wpV70Y/HSV
IJqZN+48wu9TtR2btQ/AQgkwPYsLb9fiUne0e2WbNmbo8Srj48k5bZYIKbizASzSQx2WHPM+YEnk
pNa9yjDZNASdtYazillvm4W1BCnVvbfKTMTRbsdg3wQ1mNNkAfyyZVodEaUTzEqIV8fdXkXYzcEs
dL8qbGtqI3oE2NraR7rlOtaetVgzrI0p2haSSZWlJjSqY/AXJH+4ZmJi1iZLJFtfs/9t3lwarJGq
ROdKLODqH+AO0zZCBjzTid7mMswrECTnO7UfOUgwdnzcza30gt5ATvgps03e7sP9/nwwiXr5gZWi
+L23tseHtRNyLWqOM9leCawDCjxT7EsfsMkBogNm61vrhuqmZ5i4lJRg9PjM9FiW4fwo8wFDL5xf
1k/i6t1VGGQDmLV054nzz8nHEOPNrugh344kAeOMxjGiCk2lVSkOBZQYmExbvgXXpQmuF5msamfO
UJOb1mepVWFW4gHLMWL3O9A1cKNBNWWBPH5eVJ2Wp9gC62GqekvP1yj5NpL5JGZi0s/pYsfEvtQe
6JOoUdyNMLuQrO9EyuWlqOeZCdPA2SNlJSZ0dWOEjmOrML5O0xlzt/dWPBWZe6g/eyPKjJzDdoeS
FowyEpoiL3iWbhLuuq3TFbg6QjAH/Y0iSy4tvaDJC85SWt80bqf6I6ZNixd6R15LEa8VBf78827T
xUbomJia7Xp7qAz3GNvnQ5MAPzFk9oNuRePkALsR9NnArUogKQIG3rrGkdC6B6/TDTu5iCa7hsZC
XQ5Pys99crBWPYRCvh6Zt52pJy16YhW27yeJ7D1jDawjwGz3rffe2mnFZ9qpy8DVhmdt6sjkQ3JM
J+x0+OP/rh7tr/+9QJeK1p8GtFwVV3WhDVAaXoZtUfLFFBYGxofDso9LIiq/IDLDKaZthP7F7m5L
zN8ee9bO0hunKwHthN+OkLKZB2IZjboL2+O/i8U7l7b5pmwqEeoJONv8QPvN7sWv8kUSHB1RJhAv
JS3PrYr5t6hajb8wXGMmuuhXrXddVxVP22kVZZzoBAuC9//2C/PuKeRs/F4LMznw3MpqeHlntltV
LrJJvzkwDHbnXOCl/bB5FIkZ7NtF0A4k/U9nk6yaFfLqECR0b2CMJqJ0tFWGxrv9brSp8idfiRLk
Hp1ViCg6ctIu/3ibURxrrl7q8lGmVkMCzAjsJCySMBRQ37+dSZkLLAHhNBJhccleekEfnTk/0Mur
Z+AgaNuluQ3GQvtErL6tBMir3YRuCfe4LWzLJHyjAAWmO8VdDeKrInYMOCFVaFGzuC0CLh9daXb1
7Yp7gWDGng547Lta4mv+CoKdyc+qrZZisytdVzuBN1CWceRoMXKknoHEppRnXnqsPJ2OMlff/H24
Njh3ZgC+rGYUQaUFkc8+ziDWDOURaB0I1AW4irC77uQe8mmrGQBveWBRjhOAVd9btcsx1NujUhpS
dHT2AmBMuHZaVWUESvzs791/2zO1L1KUM6CLe+li3qjl8HD1X5HKnxhwMvsU/2RffSlwDjBMcR2j
hArnKWdRPXftz3hsJsUwWeR6CKdH2BiJTnnACewC8T4LZjOePjVMrFHI8kbfq6c2gvrzPGCmuEnx
VcRhiHsQUIf6EueUL5aSH1Z9tOEuHd/e2hcpCfdR6EUQbX72vLrISEeo9HY60vm7gzmkCmii7Svh
F1JCZri4hKaK6YITnV0QAk6IHAoZJWXEmhvATFdbX3o+Za8gMfAKDg9VNjFPKd+IP8s38H/bkkfj
lP9LmwSB7ajpm60cUHG4nJ/jma31Cx9B7Rh1Oj4BjeN7oqLJi/m+RkmApv8KOHY0KUr6Jah5vhUP
p+IqjP+mhmSqsIg65CtyoHhlpt4VjPJ2dPtDQylmFgenkgylGfVEFbnrmYJPfjEwM77JOEXQNH5R
jXekwfr8bf9N2ecIVeygmV1G6VFnFLlY9tpM6/vhSiSC94H2U/DJ/H/Yu7iTvP92r1pjhr2AeC6W
CggTSAnoGp+rzzF4IPrt8+JHqzQjS7EX6i4pn18UmYuBNqPynbDAOoiMVfLtu3CabS2rRLLgpjHr
9Yulirqb2piVxKo0YYYbz/xCSnYCBcEC/Vka+yE+9ZoObC6yDoqTbrIwIX1oXPG9TdbSTfaZpyL1
sivpM3HvVNsITMIdsC0+Bo7dvcHZULBhIW8Whw4mGjVb6RRp3I5Q7fJBd2oEj6IE/SXy2ToGVnxC
9ub4Mh5X2bCrY7/OghQ+8aumrFrgcnUp1kW9bOWr4aS0ap6zwLf6fxCCHU2zSjTbwelgVe130JSf
vrSDeoj4SqtiGiKYIN4N7W5TxEG4iPUI4/+DWCQvl98IvpwM2I+0GM2CgfJugz/i7TNccoXmZzuU
Ku1b32XpRgtFCKDYIygRN5LrdPz17npC2urSMh7R3q0vulN1K7oPj2M1T6bjxtgIP64FPt9nxhCx
JnulM7sGsZHa10zQOSGEHXYy5ZDXKDZpykM3auPQK8gXd0QHY/X3fL1sMSZRIX1dxnVk1J3onWO1
A1J2t/uVhrpsDYOPdBelU8vWv7NRcmaMwqSBdTVFPkZXrIgTa7KhW8S3rF29M1afeDye83GpVba4
zGtsfcxZoEH/KZaNGxRQxhYI4upvzOuUeozzr1Miy21+gA5k2IGyLpMUxDwy0HbIbvMUnI18qgDm
GFyAuC2FqheebSiXd88Gn50Bcj9bHwByi7bc3lSOI2nsbkorcT5w6moxzRRxKbawe4eF1+6J7U5/
aurR3jn926OuLetoDndHIwwF/CCH7NosFWi744TNS7YT68MMioGGlgvZXcoAf5U8AJoAt2toIp0A
CbVFG4+RqEy/8dGPGMAzEmoJscCaSdlVtjaNv+HGXsOxz7G5gVYpIFr03cL/p99t2iC21Qta/OUX
+yLZ+ZXuqB/qX2dgHbs4qL5OIatMVNi5NO3pUpHjoWVriuN6lx0y5FYu8o6NtDvjoDvWAtwwCUxu
ew32nFekkvo02zSO1CuImEZ9TEG3Fme8rzWQj7ucopCyXRfwHzcYKOU2tOo6SOxwD7qmaEYrgFZ/
5b1u+9oxLTqJqmsADWdysPjWmFG9ZrH0vRVDnPm9VCOh3Z71Q7tew7NBWv0aioANB8a7N+2a9DuD
5mKBM5zEQ+zuuykSmTqivhlDndvFLb+Q4Ar1WzVGvID0hEWnRq8lmS8RenBw5eBEXVxVwlyIEkqB
NDfDxuonxrQode6DCu3BKrluXVZA5HRuDtDeJxdNyyEYVD4WVo4rZbN0Q3y8hN0nrgO6DpG+2ppM
kCC70n+4c6s/2udAIpMr5GV8TkD4/NUcjwVx2bWwpcfjKu5qf6HpcpiTjfgon3pJH/MZFhOtveE4
fPvsevH4Qx6wFyTEJMTrYEWk+lDdzoxdDuyMaAgKeO/t0CltnnjiQMw1fhq+jPVD1eoi97SoQARB
1stZiXEaHlJpi5UNeNVcCNnxf08M4dtDHext8Ghvtl1g5ovuSjVax8hE1WWiE09ItucqcJpDFo/3
4bjeZfiDF9fR4HMs1anKXmS36feW48u22HIzIz3A3NnCF1KaP0nnP/Ym26RF+vLowroQW31kZDQy
AWLSymDSL05KEUfEnxW80vBPMFZrHDyJ0VFMwvk6pu51CvbvU+HY/VR1Uc0vXAgPITnGE2566c65
3v074Z5WCCbOXcTdlzdp+RxrNoRRmk96CcwZegAdhCE3BViI0nhH20uh6Gcfto8UBsHUdvXZXFcU
JUUiFQqOFoIdQlkWkLzAbVYCn4QvNIMjPngaqc2fI+LGnUyzi8dLXq2qACdQwvGZzYVlrLNniDlG
Ej5dn3UW7gzQTv8C+TLzQIfh9xRmZVflbvszj1VSP36WOBsJLz0M2GC6oJ/KsfTVEPvHntRONBLV
guMyMqWZjuhIOw2qXa/ho0mGj/BLqaTo1jDtdGGZGxOCXfklIRCRRZlFcFEC4Zvmn7y27BoHXgf5
dqgZ0ppr4lZPwgMsrZ1HiJX5NVmSh09jonVUp+Qtdy+zWco/lAVXk9ASRgXMVBEJKePn8nSKsTWS
yQqbF6P1+zLCTghZaVjs95bhLLUnqb0ti+Xz2SkS+VlOePUogeUf5lv0oVlWvXvWoNy9SCAwLKQS
ioM3lDc0e9Jkd++0WTsBlqJDCWzR1lJPuKkF08/GrcEB0b44fa/j28CwO95ImpR2WdLZOxe4A39f
kZmB3RvWUzZTaemUUZeYJtqjSa0zcujBNRAx1PcMIX3Fl2YdjGh88/r3JocJnc8KXK5ZrC5RjiEJ
z07vC5h4QQvywYjPyMLnr+yohUhzQEHPYgRZ1FD7bYKIxxapr+4dl4WUj0Kq1GTI+x3ugTYJBCtY
mG4n9yb6uwrkzAkREFlXvo3HW1ESY9UGYUZnTVQ/Z5UvjAHnKz+uuPHudpxQD2anSQURc0ikqeun
cFJacncuw41mds1pp/JOgECy3CitHn6wkC4BbdAJ9GdDkPa9Ru13Rbgfx3pNbMM3dYI0WdB3T5F+
/sfRd0FyMKwMor0gt/OL4V5i/mIJ3LSSO8wkqHOmVuA7RfOmiUiDuLems3+BHIm/HTLPslEMkIRA
dXT6HAIoZOdiFwFeizPZ8io48eFfvRyiBqQzHWJyhnm9+7WwCYRhY/SiTW4R4uy1R5lonXkw6AL3
/lMt2GFWUBQm9dWnBnjJWfR+Q4OmM5eh5/173Hw3XgIDUgMQ16RV9GI9zuG3FM4o4qQEm3aKkInW
20H6tvyxRbOHT1j/IcNckvhf084K4tDrjhesr8+wvQdDk9UhVuBBYtdvTkAnbtNI89GFsvemuolr
QxWABzhVcEeZnVQm83KurxXidSmHzfUDsckLM2MNxXdXCdCJ2TFmB9yURty/F1c118gPgN9XkeXr
O5nPINxJUGHmb1efL6HkwiykadspkeXy61CZHJsCE5WwaHxwSBTGRWU8VgTVMpWRE5+N1z7zfavV
BKLq9nffEto5mqVVZO3zdA4LsmA6JONOMWMk5gbBmVUhCNbhO0H0MJFEjPa4mgG4O6ofZDPDN2hZ
HIwOsZry9SI0WvlOv8H7V6cjMM/nTRN9fwpzmomdcIOpIKSxcuavTI7Dfcl8CFG1wlBN2eECS8Ij
m1/FNKo2+QaG//ISwE/4aP6aDra7jIdNWgcyRgXxZPzFOYi9zF5NMWbreOuMhExjV1dXfk7V+xOx
NzySxHT/OGcPC4N1KvY2A3iRKFUvnhicZerJuK9kRcGECZeJ/7PAmg4zxtZPIlQF/p7gxWES64kl
XMgm0gSR1UPAsa21+zjmHD5L1ziWKrfV6P2XHmmu2Z1y9zFFJTsC5XvYdNzaPNWqJFn9s6Bvu/zT
/wn28l+3Ruty9xbo3mqe/2M8/5GKIKTfs3zVtWLdmNQ7YLA08rC6WqjDpbGVYQC246T70cJDBEEQ
5Lz1vAOgqnilsw18z6Ki8QvKfyyVPw0lXC411pbF47hb46rVkiH4Ws+S5flUaZOboeqVHAPkWfky
e1ixSDtNQDydvPuz68b1de+2BUR0djDXXTWx2NkjoWGp8MUkEejyPRbmCDZOz/tN2IO7/62cvqSI
QCSnascmf1lYK4Pp/A1xwG/z+OAoN4tvuiqkrkTyqgF2E4vAyjHjlE3FL4WOGSD5DGYZF2fGgt/I
PNN3Ni9Ep0wVALqpKOCyt9QsTMkKEUokdRjNAVXc/1mKFTsS8wIM8F0RPP5u18atJeMYoaQiu0+g
lc8Uja1BvPzQ3abFU51O7+4Ra+GFeWmvcBIbt/7cBJ6tmrdx51+ptYHpgFMH3HxVseMC33xIG5mW
ZCSkWjRZKm4XPSxzuMSqBAHrLnbmPIkgjWEMjYhhSe/UWCzQWDC690sLrTTWzaIlSphtsO9hlAWa
VssaHLTP2NV97eY7wPpprtfJ+ONTGq1X63+qpAKROhGjEYShuTq5R6AjMWzHucDNP9VNjGbsyni4
zhqGwpObpbj5PQ92ydsNPGE3i6tl7ewrE9UoIcM8C6Nd8JoCos8juk2TtkGYfYkNPS+BuMdE6iIv
jLFI30TowfNG1Vg8yBaz/A6VthSZOWhSyY0FMZf7w8QF4DfnreaktUyLSdjvOEDmF+psHN5ERJNa
Gl4qe2dhaf8mJL8yQGVzIVKdQZKsq0H67Jv2Cj1eDn6R5j+QOrVxhTLVkLW+JpVbYldE3ITBu6MF
V+PR54M80uNy8dDQhQd7MBX8CW6J6i/7DnRI3zSOe4PbsVrcpgciVwBVYTX8ZmL2Dp7DFWh7RBXn
YUG+MovdsoEF+EfxLWHLKyjD8aM3v8Tym/odGkqaD10QV+S0avKcFR0BE5UVoIhUKygh+71CTuX3
uuOP5K/5WLnsjWJwxdddgpgpzxVSwdeo90b2Ywt67tI/3+5mjELFI4YrfOHTti2j3Fu/DnztJVCq
6Pp5iIaeoQ/M1HuVOmHEHPDsDflSwzkJ/XfYl17KVSW1iDq5jSzPaFH1KN03nE7GOGIviIwXH4yV
M4V9fVhrYgKIhHXsAs4ck6PKSnDQD+blRHuix017Vb4zAJR7M/vlu6Auw495WNZ1qCGWYJV8i8hJ
LclIZIDMMQeLNvQjJu0rWhXpFtBo8XtWpZYI3gx1E5d+gAIPNsnR0w3OiwvMg5CVbfEwWMmp+MK/
ci53V5fvwqW+2buv/SA6qCPK8ZD33zM8eO7ngHYUEklXB0P7sq3m4rpC4c7LmMmIom2ChZBrWiJ6
dyCP3F+O8iM1EXVl3YsbCM2vsr6RcyDGR26b7obuNs7GEIkAkUE1DTnzLX0i8CBrxsQhXd69o0qk
/l5479izYLNGIJNJGfRD+bnoVKC7Jiii5MSj2Vl9wpOXSWUv8BCtRehKUeRec25d9GKqgm+nzmE6
Yn6iMdgyM/R197T1ikljyxuQOSbV+gDl8mJ0VZcLiv/BKZhpdhlKrBRadEvbb6tUAckdX/UDjcxH
Gt+7lgQ32rKAu/4nm34SJXAE/2zPVYa+BUSCev3qPj9j9sIq+7LFcK9Ea+1bsEirrVX0T062qCDS
POutFkb7C/Rnu/UH+ynL6vFASyChjTwpEgXFS275yzBtxnJ7Kao/0e9Ubov+Nsar/lwSJQTzrIlh
Cj8xFGkgQBAO3cUBDhqOJplbeE7chtuilF42nbSxvWpF3qmVt4O33vqwTshWc7b7htSsdygvWNwJ
SUDfBIGmykgYjZKwk5+GrUo+q2sPWHFnexHRpfb0WQYBG3v9omnynCddKYEC46ReqTHbrVZK5jyv
zNKGlTjyPPm/MIQPoFGDb1NT2QnndKmSe6LljmRqfSlLFmPR2OtlorkJk5Z9nGNdxHZ9asmtl83t
lBzhaOrJZ78T87Sh5TlE9NTS+e/hdYJmC0sgOrB3a76vuFNZv77O4puJPDavAxu75PNAZlA5hv7P
fiqYF5YmZstk+LY9ebKO8BhQHJUCgwAsSHNnyN5GXQgT1W3hcm91TSxd/XlnC400LLUS6NbHidiu
5mSKh3k8DsOjmNMCg6rhCUjRW/aVES1qi0RcCGS/rkxCt8aby3qnEXmIEt7WRsuwPIo3zx1ej9Ig
6mQ4AZYMxFKAUPrRezOSV3ZheCw+r9i9VpRnKCV9JYZtAvnMiU4wMiL3u8hxfOSXT3vVK8h3fj2E
HPD0u41T89slOBFcypJtUD4ooohjlTN6UdUkl01EqFw1yUaV7wy1xISCeGxK3sE8h1J2iv9j0+cb
1qklLN76QqZ6jkh5X3x2Lomi33XYgr9NW/7ZeLarIWtUlv3effZP7b0fCe8VpwnDtOSMPq1SeGIK
8Ki8de/v/ZTDDKZgXdyDoIykyM6Rd1/ueqxWoQmZ3KrNZ1NqxpzrBM9VwyfAij7VHbKDhvl7SZ8a
gWYr53ce73dd9ZmMf3n5mei+DcqvXeebosKv4pm9QQZ2zW97ov83+cXsowlCWbYGy+TESjrSfIat
9SK9zqL4+C+3bX2f+5XZpPQYaC7I+MhsufdmrOeHh5HN2ZjxDCtG6fAMJHa1zTUc66LttN9kjZAw
huiHImKbULKkscfn0DaHSOoJEIaEILCKIfALPrsq2sbNxtrbuzswE5fD8FfZZQ9d2h6uVG6stTpx
I0q91cCZW7rb5VK/lHCO3NjUP41bWkirhDJnJIvQDmmx/3VaTMejPuw+O8ccGj5SBO5C3VlWzKKT
7Fq7/hydvx7ep3nTL5Xkgi+DZtKg3xshHGXi2m8+Ws9YHmTrK9MiVi3B3VojWGkwouE031bpJBj7
+sm63ibbzF9hVXUbtLgDHJZPzfOln7TYkshch+2qNOBwqzjNLAY+tDjkgDS/S+RkLpwKJ7zV03/W
qddAKZz7DaK9Z5POPcuuOSbYYXqtjuiiC7PddgzP01abhu8uGyI3SGBONwHM2ygyiRoxVLVyGThA
FpH1UCQmu1riP+Bw+zrKJKtHLohBu7sZpIX/1G6cHQmeS88t2IC+ctirjV5Hv7Q9e08kMbkXOuE1
Ef6qRoe/Xdd1deXVA7zyROpQy7+79tq0uCMxyme3pjpZ+Hx2xc9U5z5bb+CdHqyCV1mSKraUcs5n
qKoB3cYw9UHe/ApN7bGw0AwNPXkOtXbj56pFpPL4k54jnvdSLimSzktp8bYjS4D3rdPNM3Jt0s7T
FlT1sTakU+PeXdsh14Rope7BMzY5GhxFol/sPIZmh30baOYCutevarqfRBz/1Jxu6p0re/HwIAOp
Z47Um9Z4DcjLZmUii1RfRJ0tNfC/ZXu/ER9kkWS3EOo7NK/1drZQSpzmEprbCLjKD1FTZrSu4Rsr
Igek3DhTjLPtWBecc9rLUFDw8+Les6z4/19JRAyYX1eLMjx/kpjo7+ZwnzqWVd0LBTQv5WdkIfDK
fRXB7BvfuNIrBwHv6TaWgR5X11lM1P7HRGEmexrn+5w4ho7rUIRWlrMLOhKN42WhVgWoV+rTF7Du
XBnV+aKFGKxAx/7jvQhc7YTUtd8or/Aj7H22AANIoyiFzPtt6g3CgUkMfpfdP7BwCqNMR6b5BK8x
41bNJEsu5k8p6xfYDTTd2hG6xzYV0LrHY57f5m4z/VcP2+Wd7AeQ1sxdWUgvi063itq6b5KckLp1
SahavLzC8yacmfso3jMnybjakssSBNgkmHdzswQFtvexBxNtIMxe6IxHvEbFVUIxDLEH/glo9ADW
qrR4W9ISlrmhIJPpOGyJ1W+gtp2uzABoGzP5v9XGzhWgrX3b/CLlIHTqqbc+4l1AgaN2d9y6V1YY
tfiZxd9R9HTM6FDOeSODVCmlYM095xVj2Na6aPE873VYwHqZhFieadUZJ236B7NB3HyabFUeBjia
TUOyD4otb70+6OZRolMqkVGgVkR2SmLv341qOQisJ20BMNl+2yXfBDmB+gmaFj2o76Fhjd2QWRqs
aeXUtcYXZL5VP6AsruL22CqspXjsYsSL00XwcZPiDx22LuGsiUUrys6z+UDy0aueNPTr8MjmgJuU
5a+QiSFe0a5YSAz4r70LMQlCNyYkxe9uMgOUrK5QJCK22XzrnaaHi73LYE0eWiPA+ZNwDtW2E+XS
7eU5St7NIzys9RCfyhBsV/RSGmD0lyWPJmRUXouNWc4oLms+MvgPzImFYPDyVu5Sx+y74Ik8KUFJ
FutPsANQbG4ACNPrw1d6UfAWR6j12WQvfutFMNQkljfQU1sml3IsTnef1/T+1c2Yk541GqDQguoD
2j8Hu1UNttZwuJBjXsR9H3YWAWM7e/5xTo3IrBlspRYanlI8J0SFARseulI6irT/sfG7tpKo5xvT
tPIagGiOVCoW/1YoxsKfCPX+AKg73awwoDn36uZwy51t9BNQ65x+3TSXNqiblcqYvF7vsmW8YWqX
MQBrCBESU8axtc4PHJHbnWaPK7ri6JDMmarTyGC0dU3y77FYR22RGjtzpBuHnIqLpltzpStBDBUN
MrKMI+Iuar5m7qYBMnL9fH5T1hHCNTACzY/363WZn+s/qohRrSw9zBxFcEHlYzJumOEfM3/tPg9c
lfPluJ15oTuLQW5EldVnm0LlErgZeC0rWcQ8h4DW5o8inN0TQiYtn3ww0zhsptxZEjso5csrHEN/
7yFlbBFW42haegRPtc/ty0o/pa/ghDSXcd/4bnmIISJXO/quqRNBMyyxtVFLOfYUQxCg6JtpEYHR
qPQUBa0ZDZoQIblJq7tbgwMISALYu30YBXjvy9uEOSCE/oncRwWSZ6GBpT4nLv4tYFFVIuXwIQ8/
2hIt5y9hJMZc3NJbkvMkD3t9eGm0GgS69ZD7SH6kSQYzaFS7/tXM1SDVGyTTXkAUUjumTkwrBh+j
kfxmBixf6VQFdoAdFfBH4ROP5p580BL5Kyg9eftsFTHhywqU0Inc+1cx0EJZJjydFhzpWhf9ryzh
2omoEQO8iry7Vr75arkaNIyGItiD5NxZMXtgQ7ZvdbZ6kVrBmaXY05FuYRxWIj4mNE9Mcq8HvUmn
bXdQyupZEZ1ySmPCdfPFZ5iuUtUyGzEi4jgztPNSIYmr82CEBfysM+xe4FWobt1oWFwT6vt+GyKB
WrPaYF1A/2/8rEw7trhCp2O+ZESLSRcR2LyqheXpl8DsVhXWve7bCJujtVsaT5oT5E9AvCxb20Qm
t51qMygBOZKUHcuDWUlsv+ZHTMuw+ohYYP721fkUiUWK8BU3+CJGGpMj4y+TNlOgwXZEz9bhjtCy
N6JmnhncXznuZICbt+QhIGove72UW88BcP9KJGOvSm+dz6OA5Ks8ES0Nzm1lZp4TyLM8IUpXW77y
BoKGCoSeKostEJJgWUqVLezbCGE55ggoAlP8tqArcjF4Y0c5l/7ylpvC3IA9WPx/X7wo93FG6a9o
d+DnqGXor66v8+E0SssNDBDON//SDegXC2f8LYSxSKz8E5sq8/xThYFup3IB1GkNPjKuDxMZA516
rm9Fp0fo4KC1lf+LxuxVe+FFeWnSSxJK6Z3PI2PNxjeDr8x0a2pWsV8gYSVsLISdNN8FJCj+Ha5W
r37NeZ0yL5zjSk5Qphk50NxRR0uTB1EzSV2T3Higd8uknZ0Bvcg5DYmK6T4i23PkzMcHVY1SRKRP
D4vU3LtMLhP/qwWv2xpEvU3wIuXO8gifA7VdguIdMWK5oq8EtZy0pnSCAirDIcO6OS7c2CH7stO/
N3U1BUQ9jFu3P6YsmADdPuRNockt5p0ZWiUUIHcDmyQJWqi8o5m0BD2Oejrs0wE4UM1bkpb6r4iu
SoUYcNHjCie5/sTlMZb1zM8LU9R1TsRoWgtW1+KgAvD2ntumcPReeJQpxqIWtnvePjusnnFGpvt7
utbbpF7rnpdXUpzV6bY9ksENeZvPWsyL+h33O+Rhw6SBJjO1VdetBBKqlCtQhHXVO+d/CCYGCekh
O+DQOOq3he1Su4j6b71VqqJBeG6M5N2RfdcTI0AZQ+AZUYsh/uqtnGZZX0GTcq22wOo9ik1COavG
ZzWN6yj7Qd/FdnnMHhy0OIyZpFKT2rao2BZxZnY1t07YWC/3YGpcx9tVWnodpoFb/5XLaM64q0vQ
VF6eFe3deibuH7Svj5JI8SJ1RqHtVwIDMnEKfXHwQH8IAcAhK8z7YDdfDn24NyxQmBGl+zVTQo8y
wldci9dN+9otwJA9bzD6rJdcSGYe1bxEsS7ccYbd26ayKiSmCSYlWJzIWHoZhda2OzZvxzop5UFC
LP8p4xW8SpyXF1IcP5wo8b/9z1YuH9hst8OCuOByq/KauVrPsPwdQxj67b8lpgtIso/gWqnctmFV
x5WQTg9k161APWI2mjCESJWmxU24Co61NCtJFPgLmKkJsab9pLj6v+fAWZ6KroacotBwMlAIScy9
VY1pBdVw4gAGALZ+vQJcep/6d5+xKZGCQtYw35tSxa7/I5Lj7D6RqY6lYxMoG9a6SyqYBuVUv1zY
EjwJqjAFB6NsUjzWOvBqLhDr9OB8+99TyJWDy+d2X1ByU/zEMedleg7w3j9SOaT8BWqWk+C8Rlbd
xjLVnhiTfkC7rMlUMrqkpJukDwLFTUjjUP8rUQChatzJxoAba8y417m8HrOZd60PdVCPg6qSHbop
miQ7FtMwf38Ckcyqw7sM66D87KxN49L75P3LpCVsZ4SxjNW8c1Zvd/m6Mvi5Cv9azkkRLEidVg3T
cEY2PXJ9w7yDmQ/eXQxCbcXO9i9bLrtwRwKfrxKKjH0BXkFmqO+Z/FSYk9yxXRjW2TVfkoAvW4p2
/aaURA1Cx9zExM4zcnhLCE9vHZ5sHfZKF6pFFPl2/CObL8aVt2JULxEPP+WsD99C/3h2qOIl7AlO
EdAUGAvMDMBBQqkuyGznNjMkPu5MDtTyefDkddrFlCdnwy73DQ4OErp3nuRlEW41vMrKVmKAcykT
xvxxEZjf/EB8869z3+HzUPtqhK8M5i9CtKB6qHk7J138rDWBb2WGzgFq0IQ1A/79GCGRQY0hsgks
YyOpPZSsdZTNzbyHk94Oc1dKFLJXjME6j1B+uD3DkRWczWyWIyXlxNA75fj96qYstPT86mlaPjLe
45PpLiSsoarJ5oRHPHIH+x+CMXZ1o4dSiK3B/BZc78pKDnV7caa0KkHYsyZaQR8YJ4ID4VfYyGMp
xmDtg/jYLScIVbv7oYu/4gXMqWN5CWtjOBn+j/ajcH/lUZXLPIvuJNQD57szFiKCm9OK6enNfpO8
eHdFo55XVk2QdCgDNykOos8K01+TWFNc2WiHNuRasqiO6891uQXkJx/bqFsJPC4omAix2imlRjjV
pN/FNciDNajhjOkwgBCXZFb+bwUZSJiggXamj335IgYMspsUkMAZeXkQ9WkgZDP8SiTdW8nGMFyw
fbgiwc1wb9OvD5/EqglVMaq8V/J5GIRvcS6tznaL7Es+BvusA1MqfsvdhHhuwUZO7kxE3tMJIiJJ
ot6i0PMQs7BGTerPpmB3XqLkwjSyGVSO3C7DSH31pxZK3uoAB0/eCbtxkqs+bsyfDdMhURuwUP7y
cBthPgu9pR0l1XVnYbXSzxanC42uSAN1JnXfwONyUcLzPaFd7/r0SDZ3R2Qxe5b4ViZo/KCSCDZ4
pi1kgm0Zc4ByyU1zfnJ5LxbbiVET/XGAh0aWbzoKaRtQnf0/mt28SPEGX5iOZONTJ4dVTdAvq1Br
Ad1DlzoRjo4R+jDKNM4a3lhbJtmfFj0IGb9sGCOlxpqRhH6Tqya9IWRJVzR1kGxGMJK4pWo2Cx/B
XDuSFHwlMaxN8KpFCp+Z9soj6sfDHwdQfGKlu7HOnl7Unpd6OqVjvGay4dEdSKVSVNhaxYQWxZY5
+DXW9Syz7Q0hOePwv+gALlHbrLu5CY5JKsYY884l/1SfJz1kzvEgGtWJafJmEhBXK4husTHvW5a6
cgrICEqUlAbsLi2MKNdL3JUEApqePrDDmvU0m0mr7/apnkYFlflX4eA33eFN5XNWQ/g8h7REIYib
yrSEa0tIexupAStDHw6wlaneQBSGEqAcOx/yKGOBQoNb9z1t6Yl+Jh7EdVmFyJDn9uYsFjt7T0g3
q6Ez6cT+XgYpXFE+vqpm6C1RISY2d+X3fPYhfXqqpcQMt2uaSGC9KLxtYGbDMRbveziOxO4gwYw6
BH+WzAZ1gw3RNH6yu1eE8oeOcD10gxgsTolhQ0pZwUfXKh1jUbLTr1qIyvKSP/Fmek/TWsNF3GJw
RRaqJr1zHyasDizKh2Q+02K4hIOqPDXBoYbcSoNjVmJNmSSdXaNn7Le7QQl/dti23BuYCUV3/pyb
5+3hVGfbFUAg94Q35lgdDzEkaYa/W8ZNGUukbkwG5CjgtHKGkpRdF61SuRaVa0uDhKhRE6v5cI8K
p5WRZDRiS8LJhhjEkCAIYnHVXKk0N1RwDVFoJgRNNB55ahtUf7+pUEa0Jm9ZxxIeDyyt/C11BRxB
TVymaLzYUevBl6/t+hTHhwb8zsjP1yK6N8e/5+H6qXoiwhX/MEPOcUN5M1LvPltbVAbfjb942TAT
Xk4oLbXHDyMw0/OmlGV4rRWGXtN+EXBjnvNxRNa1lCLR4S1qpghZ5+Wx+YlH95IEO4msioCJHTWI
ciaexsceSUg5rLh5rRykPhxeOtVYuFUTa6BKVP3iElQW3lJM20qleJLpekbjYpKTmaQassV3KeJO
v9MWWIg9pCxFWDuluXCnF279iG7D9A9hEZz+Q9t0Y2G0KwgpPrammjqGA0H4fEJdIIqbFsCpXJvy
M30SPooSFENzgAztx9YpnfrtA1kuNKSeL4z0sUrHjGDZNXplz3NvJKbMyv+g53KGZXBTyA0FT1bj
5cNa80206l5hBJABYTySQFZKa9fG9uwrB185SDFeBff7n7Sv2h2DW9TsArnjFy73x32rbkQXzuJs
LCQ4Dw2+CSsAgsWF0qp6U0mBMitfAB3/A8TG3T7L0mJ4ttwQ5BuD27gBARTQ47LZpK1863NOMXlL
WjaugQAGudtVJSmTg1lJlEyVhzl4kxtHB1o+nfl3Kl1RZG5yRFTaSnQMua70Mle63ulljcXTlnQ2
0PzPMdhPjxVSWkG5b1UvHY2R+eHrXqX3ltMLSurPYnmPHXtIn4xuep0TUwj3dm4MJ9nIjPk6OjxV
F+ZNmBrojkJMiQh8fKeAvz53MN+FFszSeJMM1Nx6t6HTrUkORhh5oRvHzbHkpqXRlB8gasJ0kMDb
0ooBfn1yUFPopgTHm1KWEcs/tVZXTpuzVGTJgz8vpMRtOvU2rLpIjuoHboIkp0sFDJORmoKd0PwF
SY5UZdn4ualFGgvufwZOhdnrUwdm90AbuUrqJe15W67UV0YZ4zhMMe8/JsiEzQM9GS993ZW4fPig
ix5NUpU1/K8/ERUEvOnrh4OYlDduFRnpcpknpEbOo4p60oXqvRTYtIGKreyvP4O+3mKCt5Iijak9
EOf7hRpjE52Lo1fOI6YXsz8apkAWzbCPc2sGSNDh9A2yTwEnWNveead0Amp4bDXtxu/XohK8gdq+
nmmzUA7KCMDjVnQfbSbIMLqY+wpPBt2bgQmltTYodOYdZbS262t/pSLWdPCHfyjld8EmuJDjXHi0
lbQ72MgYV7f/TZZiGotL2tTNzcQbjBXL4S1ZLq+tShSVvilojkqjCzILedlTIoCFurB1jDWXesht
ySvO3uVn2e1jOtAyhNXUM3OiO6BqkXk9FPAlSMNOWQNL9tH5G2OfKqGJqR9RhR89IHkhuOHfSZRK
RSlnZjNzxosp6XE66/9kyT2m2U2GooqMnmoIw+bxKWGZUSS3vnSDfRiVc7ShXMmlxf32NSFIo0sv
OU8z6vxKeI46+xGeMeH2qDSbZbiKX9XbWYuh6o/kIWjTATdl7H7tKs0yn20SLCIv/K2xNQPUsVb4
DXkK4SlBqJvOlBaGvraLA6BXiNazLqFJUageG2rysNfvqDGzwOJxkKXHMxY8+tuA6FtYHtx9K3IA
WQffwgRfj+OzymNUaTeah5NvgCEZAPN3eAD59ySYzSQOAH/BlkQByPLuHfQd
`pragma protect end_protected
