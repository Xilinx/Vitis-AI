/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56960)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvl74G/mKAQRknkxLdH3/dLn3zMAll0DTXOh7Qe7ckK3v0fT3L1gNqpE4g
acY+zs4JrrB9h307S6+CNKdL/uEHy59cpZxrFEXcezADhDOpZ9sLUKpCefYocVCvR/+vEGVAETBk
PeZM2vJm18i7gYo1BB2jkpSgJaXIN2UtcgTOeM1OmzWXpZAS1dYrASborS4dXnu2x2ChPwbww1Mz
Dqd0r89bjv+RdC1WUOnPPD4Ri0fWkp/Vg6dO6ig5oSVzkjCkUwbdFuf14ule51SMP0OUqHcmdvNX
a0OKMcPPQNCzjSwMwWhLUog4rk+oX4ZR+3G9wJw9CRYwpBJZLGCGN8CWRKHi+IdvSHFShlfifV3n
kh49lDtYrWlBAtuMIkycp4CQ26ptlEQTz7atexUitoVKrjEJ71f2HoZghfbdemnzn/qfsSyYlJ/A
G5QAHfje3gR/7uHZNIlnFAJiweK7i4qMFwwLFk3GhPVHaioToRkJh87YwMYUSWfy2alLtheKAOHo
82FAYXeDhEQfv88H6PGtSfhW2oqZmA0HSr4ZSUGEQ6aJMINkeCcemFXAz+uda+urWADIdURjnwFX
fRqlikgpKSXGT7NpjlVKxbGFCMuF3iCdHP6C4iG2tAqDhEug1ArKwIzkGTfG1ex/mgQ4UKkoyK1I
T+okz1n4s45l7PNZGqhq7A+U2pNw24BZ2jq3xIpRxRYzrdMUjffvPJBRUV6AZu6tVgKVN/RxkjxC
3UKdit8OttYLD+0H0PlbYvs+5SJNsP02UgWLVTnXUUcMmp5Rfd8F9FBkie+UTNluVcs8y6UgCUJH
mvRHlL8XEUoFi6WCUp5BFH316q8WpsqU+JpH1V5jIuKV8CAXhpHGtrJgNpAp7zYzUij8vamjZ9aK
NUsXVxsZjDtd5XJsJhQw4L2F2qXkX3dMsvoewvQWGgzC6y2yYXlvx1CA2ZY+6VnizJBn+/t3Um8s
StLMGqWlaau8QFPymhKjybseNwIqLN2Mk0CaYhhnRL2SZQRwbhqhX2+V4Tk3VaiK/uOKxq6ohNey
d8uRsLmIkBGeBORdkt3Xjhr8Fy91HB7N4eoLH8vnbGNSOnLBIQggWxESNd/wB9nKSbu1Dksamhwq
bRimm/OdkgAy6trAHEOLAWYLRBreu12pZh6nAfb5UiDZ8yef6Yrkfiv+SinnGH0ZqJWKeJta3V/1
dcKEnr6Rr0RXDMFDZasuvBPTL1e2ESN8HnP2UfyRui7nS3pVsETu9Gr1Ssf4s4g9KV9J6A6tDTOm
XF1+d6+zK1rqG1jwhTk1IlitixieCJJ776A1uZrdWAVGhoo9jwvFZkGPVTHyRfMcsVKuOjuNaeyI
3uQxGHHx9ps/2H6ffZuye34qWoanhWhCund2EumQv7+B6X9Jta1sAURW+wl3zYUZPfKGbTMsrebR
6CzulGlv5shesm9Ogs+MXFb7MIm0XWr14AmFBCY4CDsSbdIIN8WMGnXdCfI18VoZwQ73uXTzI/IX
o4vPCQBzzjciTbW0Y4C857970Jd5+c3F6sqjlSjiyFWX0WasbyaCqnmuCaObg/P88yvX9TvgN5jw
oILlASu2VrtfEHWXlFM7I2wTSCum2CYQH2ZzABiQjZ6B8d1vwn9tDvj9PFTmxeV4UpEU8bxZ3oZL
3ZgrDJ6v1KDzr1JNWBgFVeNscQrvW422FNJDc1rmgtnYS+PUD2e4nndxCphXVnS+Y0knO8E9M+3f
9haMgs3CRLXdYcU3VnFRDY+Pi3qlGaE2biUhMdrqn2dwVCXkfgSnAeS+LhQkuAn6yjPl3Wwq4/8l
ECoP/7BFzD5xE3V7MW7MxzC81pEallpIE3iczWSlzcCCyK+x+/qSr4klP+LRoLU+lrGKxeP+4mKQ
EalVV5jhuFxHrfGFu8GLvwq8Qh+fq12nN3wjKwN35kSRbIWvfkLBa649w+37lxSPfV47fec+FWpg
fiGCcC0FZJYRZjCtZ1/e9/XcpOYRSXoCWStPO/lwA7CYLa58gyXb+1lz/6XB9S3WKsjAZnM4ZyQp
rLs6Gs/uwYYNut1iLyNQe5Y6hlBqn+6GZGvCcrl1L/rARrVspM1DD17vFd10633r80iINKUfL06Y
Rb8KWpJKjM0yZsIh+GQLH7AH/KmbKei42gdLDz7ZOzDrfwbMiUOAacdHugaZBLl7Kij6O24UcjXc
pd15ccp4aCRW2+4AlKOCR2z1B895iLeg/bvZBw55tmhZINYEXDfV8pQA/SLIk8DG5z8hEUdD2VGs
hsCPH/tyutPaC3MNoz0Ji1BExSioCZ9Ovpt4QN2xHpjJ4ETTEmrUmbzardQ5L0V34uxMdKkiYIgm
DcOsih+VPDrRpNdYqp3mQAc9GL6PbHFtrzu3vlNYzw29iaJeOKKCxWSAcuP51qk/R8CLXgWNnLUx
KzCk5R5nB8t5jGOBvZcXo9h5kWr1zBNawuGS368NXfz4SfpeX042AcnmYQfn5nTd6hScPRM1Dn5b
Yfo9QK7AArnfV67CMiSRTmFXffwstr7AAhT9Y17sdyPYNjIVuUHpksY6vJryznEDBJa/tNUkLslO
jugndevsTVlSFDE5syIYJt1AXHGTo/96HnK/R8jMEeCWHePAmVE5cjU72OfXOVyz2SefxhfUWkQS
XymlNlw2VigJ4jmiIDeVtxwxCPnJsihOqB9mpTicrrPoyCAbr7kSu2HTxdEWNMOxS0/srqQggnWM
YhxXXjVS7rMsi9myCcpiRwSnOsLF99fLP7WGzTHBBwOxtAqa1Q0//BBW6NpyYVdrf+IS7CcC1D/v
Z/1RD7MGGJn4tzSS0Xv3wMFx94jUsLbUuWZdvH6yYZoqWZ0T0Jo06K3+VJ+lDm/m/qeOsFTBxNgx
SRjaYnHXjKAN6cCtRNqieKf3krYrgEP1S10aIY3IqGQ2f7gpyDOG5bgjsdWG4VpCUmFFGwwxkilz
SvkVsjV6NxK2zLk3wyf1TTK1eAo2UAlCXUEXddnz25cucIt9DdoRCBVUTJRtkYg2hxeAa4LIXdbm
cQoDJuct2t8Tje4koZuLsGAKr2drqVptKOEK4mlB6sTUB/UCJdSS6Gxsct6iHxi6TDN4lP4+uYu6
noVX7jo7YQ4MTP++J++MAZ96F3Jd3c9HlN5Da/6nLp+mUdug0WHXlsyyWge3eF8GvkdnNaErQUbp
rpK31YolZLc1PEWN6xt5fLqWqmdJ6OiTH1DRX2DjRNsQ9w+kWkstnTRleZWl4j8Bfp2lLWy2myCp
BkeXP3zKGVagjxGxOFfA+ZkSjkLaw1wMOWrq8n5CeMPThBeG9knAxWvwDGsB+VwZHNCw0N4dKdVJ
Wf1GpslKnW6LKAroYjU2AALkc1k0gRtmokBG02xqnFkv6B0djSr3WGAIttgnVJPliYe0qvUqNUJX
zYMdd7SpX7suXREaHI/8YIVnSXKrrJEK9LoXj7rqZuVyUCaZVoemzobUL8/8kqDUnGoqoZMIbz1r
Nla1+cwkV5EsRawIkQeXdcQU/Q0XvmF1C2Z6rYM3Tyy5eNo6zr40+muAuS0FKlcs6nyH5c5/TU0v
D/P7Q3mwmRqEj17FyVYWXgKHZaNF2+S4e3V49Y4IOvY06pa+eZDu+B4VifR9h1WZFBa0Ty4Bpj+1
45Opyaijxa6pHCwNZ3U9swLa9tw4xIlHMZEH9vvaMWUr01XIj4qwnQ7EZe+KY91ZUQFL/kJ17QPJ
nxDNOz90NQeiZk1dM1+dn9wTjg9QLZY+FBd3LEhk9gRrCfy/YYRV+0SEnKT6nPshZfTROMcl69eG
59Xh9TSn4K3fKGVG7hJoA4BBU1vrG8R9+BkijccFn5/M1qC46978xuzhCpLijT83pC2tZh6PUVWl
SNsAwXKOTrKguaH6+J56mNv6Pz2bEPtMV+ljFXzLNuvM2cGtNhLMaSC33eWx0vrRxkxCR1jqrkaN
5SnBW9XpYE7eLXsKNhbFzkdMvIrUfbDrWyZJY9zNF37awgtO9JPBB4GEISew+0iSqT8S+qR4dT4u
CCcpclfZ35msLDPfluQRe2umNoLZdjV+LLLrfRIk53GpjomJ0jjM3uf4wXc1OJq2q+jGoxBVDBmb
EoU8f8MfI997fo7Pz1F5QOzAMkUf2duQsxjOKWCOH+dHAZk0VUcjHFtrWFpi47tF3WlboR924zLW
Ya+2qvHtl/W5oQpMlI7jkwPvliTcnOoThJO++RyjsnSn9lXhlNQXhA+J2uMptmm5v/YcvcsE85t3
Du9W0qtzA/0cfxx0iJubRbaCMq80FS91X34ia7EFG/FhFtSZDgHCDkETTCpqqvGFEhIwuwU3U2Vh
IX4m/T1vsYb6IRre89IQPBxr6Ka0SRnIpDzSNtG2JbMinNoorhx1TT1OOr40ZO/XYTR2hkMJw4h3
i1qPK7w17rEq4fRUb9e6WS0I7EVAuOWh878LfpNEZRpzZDUv/XqrOW2IPatcZPgNWlcYSDBQSyk7
CpsMOOonHqEQULEyAPG02zTFiy8k8BwcqBHT8RS3Ng/Wl33RMoTNzNtCjPy6YNqezQia9Jcjraib
vqy1bjcpfCKURqKTbnBpwj16tVXbLKeDtzm6DOP4gdCE3JANNOkEhw44ui948oTVUuYACtVKi0Zi
qAyTL6HBHjvpJevsgzxNLoO0yqBaxq23iFKLFCCI4OcBIoyNt/GYh6XZjASh2NLazbPHKFNJuOP5
MRLvQXlLzBYrIqtd5Fj80drSI679v7v3JRqcnceoyiyDAJWWVEEN1+EZt9xkW8n0avjAHxI5tpUf
CKSVHE3XXnng8Uz5MvtW6J8g1zL3kShqu/B3PrQLwWbk3Sm1oIcEGxaUa7EYhXZJ/vJd160s4DUP
tCioIpEJY3aH6oBhxqruKcp7fZJRfdNQ8RMtQu0EQVHfV9CBC4ec3J+ZbhV8nmeAeXkMPCc/fqsv
I/8SrUlF0BjPJ7cTqmee30lhaarYckq6MWsXY0aESV4kbA06Q+WSrmIVtOplSLlrafaEJ6rFRDTj
UksHW8ILXf1p0D1HIaAmHr41o7e9xIr/9wWtJAe+5xgEHnYiuetdPusDNZ3eENdKJo7crQZ1iFCE
Wd4mO9oYdh6pi8uOQq+OWe9W76bUe3rze/lOc67DvPApsCp7NM9W4AzkW0L8D4ooyr2GnZuj/b8W
ALGVBJdsscu1P9clZ701ny4HQIPajeIk2YoxXSEF3tEMMUTskEKE0hBIAiI46988ECu4gi2CWFo0
dCqtn0uwZJLZWjaEcIMdiEKxxf34wm95P4CmlPQ+rW46+bfk9uqVwntO7hl3pDlprbSaR9AxVAYk
JuhemE5K1hyZD7S6niQV+bKgYhuotmOkKWaoCzXc6jdXWGkUIPCmALYQU53f1zopqgcD4sy1JxKQ
esJOg+jKL6T75Lo13mBqOmvYxUON9SU5aMS9lC1jxxIQtWXnmX2h6uQdBD59CIJto+PQaWHv5PwU
d+BkbqfITVucgswvboEUJbVgyIjmqcuiN5g7u2Pun3YLMEQ9T8NaQlmmcxbe67PlGGERUhgThywl
b++voH6YKIeXKqiqtsU07+GUYBJozfLwbPjtfdFy5674gCu3UiZb74IW7bHYbIVEcbphuaJho48t
8KzLDXc3aTvY/2tGae7BthP1QqDc5gk1vxqIKVILyZGCxqMsRHMSaJ/go1EuvF+A+gxAL4uyD8sT
sv6pJbgfneBIuIwSc7+QOGlbyoDrrqkZIAeYn20OefrrXtwGCiluYqC30EHUOsXxQ/Z1AF66MMQd
vC2m9Lxi19MOhYnbUKKKCq86COu+qe553UAhm8gtl/h3k5n2MLAfo6u253IFqErznQTlbSHOrF9/
t8LuEEVkUPiKrxZ7svrPxYraSb6z71ocrYwfbrMRdc6r2sXgxJou1gT1IE0a/bZoGr0OhMUsBabR
O7DC6UnXmdVwJEEoxBfJdSWS1wWJwHWyMUHnN3BApnIiYonOJQ6C/LnSgFrR8pnq825+/nxS6R1b
7dQFCKrYQKnTwQs/DIkqwaz/1iNsEcnU3EaM4nI9qDkovz/oRc/OLXcSY47KzJdCLNczoox3RaJC
NqMH3vh0Uj4654vuqmc8nakrAEimkFXlhLhVC87rC7HvnCzj0aU0LKWE1GC4NIAgAiHPPoe316ib
EukaDpHC1hbO/VODMJv+zddWcjBoTcPJCVSjTQgQ9Q82NQTl9p14nJoicwvVhPADhBYYdSZ91NnH
YL4T2URnK7gVyVHey6CFihvyKz8qtY7ZWLhLd5i2lo5xD/A/dccyyekn6V0vYekrAsNhpJmAL6ZH
YQuwXwPfybhQ/myXIFX7aDgy6kVMALLhqDUY5kHCsezJ6Ye65cRoMPq1lMYqmoQdpEKByFx0TF6n
Sv3oK1bBrDaBsS2diMexGSv/K4ii5ByAYJX66snRTFnPOoUSOCpUKxD8cqtv6GfCMcFRNgNDgUdH
YVwcRaVJZ02SiLqyPDCOgQqSg8/OYY5jlKZcebKTjbvExU3bxzDhLj+waT29vE6elof6V0irnIQD
GHVENxjS90enAU2fBogx3sPca3YZGZ1Syvnb9LYi7pgyfu2wwKdwxqEvyb5Wh6paGPGRxadg3N66
e4fHM/f3KRs44XsH+8OkDu74Ypr+4GqoWSFMVwBeSRgRX+ol0j2QSno3EZorBKHC9vR/V0hxkfUX
4rR/wy+whzhskcYl6G1XVelt8lRNhMoIdWtjPPkitiRgyXpAPyN36obkHNYpc+aO5YLNDj+HvGaA
y86pLK/+r6gdQkh6jG4JEoFpR68NZ4Hwk/Bs6CzfZt6p+EPTEivV3qe/arxF04Lvhwv+mFVHOaCZ
LAwjvktYCbyT7rZ3rWiqhE9ptg5Jn3e82w37bjDRQAkzIV+CCI6A9gKlQfWLWsWuf7DpPAlW1N4B
Lft1hy87Di+F+YFe8l8BrWEfIsVhmoa4oZ6pEQFYWDUiBCdLnFcuKS5leDPUYrnz7tr2w3/GCZpO
v+CcZLCa2kqrimAc1I202Sxck5/O7E2uadIViHiwySdi10+cJDcDPPSFKn6XIzyHZXFatt+S7+/K
apfuD6ouPad+rIsRTvq+iIr1wb5UcVoTsfONUh4mga0JDXwXbliOAx7DBgha8xDfYUJD0rFgDZhm
/MNRVejl/RNpnUPwipq7fa8qz+9TuiuwNehzkCkAbFSp68Se/FtluzG3C8o7aio+I4NWgy6x6Sa0
l+fjXtB11OlTQSVMBYlu3ZsOq9JbjTBJNj5M26UtGRy7lHVHoDigl+4mvSRRJiMPo3gKvbWp7Yl4
hhg/FbcDCnRySKOCkcIEZr0wH3LC1DY6hZVHu8zrdGKzbpGTBBFqSFa04aOIuv3C4CeVTyqgUBLE
WTeGu4GO70ogLqTHqZbSBR8erGV4TZKi42YeO5jYAH9LyCEI4gxHHNy55Gj1Vzn3IFi6e2sCCNmu
ApWXG9105z3y9stcYbc2crdvL5MQhwgEmUsX/kdBH1xeApLb8c8aVQ7uXwAjAu42yCIvdKBSf7h+
9MSVhsbNQtECDT1FH9NRsd3DcWYScbKK9hwxdyyy/fXfpjNeMul9acrrP1v+qNVxo+aoZEp24xQ0
RLejH2yDnKV5SQ1+8q20KoAn0S4SVT2gSII48OctPk+86d6P8FdgNhdkxUrbXGpN+mPMApdTHKC4
h1BwTlY8V9L4w0ihjvWOD2eNRtDtgpTo+lSY1Vxp9+ovbn1i+66mEyWFtzHHr7WLxqGvgAms7cSX
2M2ENEbqGuu3OdSoXMGwxpzJ1ccANtpc6jifvnZ1FrAmgyOfhTmxap8J5IU/BqF62DGnfWg9eQ50
z0cxpqUCL+q1drnofUfTjmVZtQdj0YJE3rwB/TkLe02FC18RCtwe1jCxVDGSvxaxrHo4Sq4pv14M
pHyoE09ab/19CkZIc1x6Xb3/4p7VD9bMM42nEMdvTyXAjvQ5Lqh41dqen4AjyGG47dSyP5IgyWfY
uQx/y0cLZCTm7jwTn0nM/ULpcKUZ+9YdLpvqg5LXEVv6r5DXPxiGWNkUC1cMJfNjFaEEUZMWxF+I
pdGNbPuYM3IshNfHsnTHOmPCN5bkxpRECTRHflqVvxEt2P8poM6N/3CHeD5iuPMnRseeAY7RUKVu
NfWn9IiMco04k8DkIH33gUJhAjmrUoKTH48axnCoU3zzO+2DxHr3ng9pbYo5uvImeL5fmdskejBn
N7m7WbNTv/u7zYkxij26LXhiw9TtOGxssJnwGT4ErTYMj/fkvBhfHI68dw5PguVHwPMO5Vhq6kiZ
YZzaSJ/EXUNZemO4Jv7F9EihXGAmRnitQ+RS8WgiZBsvDcD04hgzdy3Qm00xocXzbPg82W+fQsfo
UZ4gGkjUm2z3jeOvOPqBD+UACA0X8wqPSqJ+kVV87q1vGpaQFDuFaiPp90L4U2Ow/qB2KHDAoICN
n0ai0BGT7vLbeC+NgRImlXdFC2wZws+dDG2qxO8qQtMRoTcqQo6C5cJ0Hzr/VUnFxmC22QhgIyMs
pjjs+GoupKXd01xEAe++q02WgBE3pSQKfnWBRSV6UBMO+qMb9evJGs8x2l3XrerNvgcHiatQKIJD
YSmlQ7MVEjwkWM94//XVuXm1ogAFL/5BIv89ByjIaFg9YdTZBFXUOb+d8aGtz6XwSj3iqrb0HG/x
we/bVPd7ZhaBdtue/n0qsVyG/WCiT+TNa0nGk6A+EiJnQ3Ws8dvjzKcvGKDdAb7ho7oEjE8X2Xp+
VNF1cWDdwL4B8auuj6wkhZ5nQJg2rUey6ZlO3yvbpcxwUIGiQb6mOIQn7azrPevTrCx8iCEgGEiP
Nc03OzlggG7s/fSesn58aRwCSzFEiSP4hmLZDRk7AY1tS7pWyHWz/KBPI/RjxJjRnajWKeE6pSpo
p1SlNuYGv8/UORTt6dt7JxKYVYb4tb5N7d64GyOGlKxOP6+8gYnl6T/UQMRpBXxErUqSRdh3w9Go
Oah/5YDtYpDm91lsMPs9mNZ+qcOjjpdPPCWv/TgKfzHoXPVcn+KQiPCZZGeC1Yu7LNqnxwnepZkN
VQYxhYWm0StkaVUNO3ETnIZ/Y8nuEJGa8yz8SZg6nqNhMYfVkkrLyAWoUnY6Mrqc+ECq23j7PnW7
HGz9qNKcfv3YZAu0ybymEARKnluWXj+5DzYyxZcTRvm92KOqtIbbOoJWPct2y5uccF4yB51mbLDo
5E024iJj3G8MQyIXBSuZ+T1t/yB97HzgXCPWpzdp/td3Rwj1HSfKt0krQsyYuN3czu+EgXS6nNeg
Zm/n44mbmeLLBzI1xeAG0yUoDIavqv7TpFtTf/aXYsLb+vMUAPNjHKT8Sfa3MAwj7E5teYOyDGux
sASLqsemHyczp0qkux/TR/QybM00XOgJWVOH3gD8IavBWv5pgBEi1sij33VDtWW824HP9+C3MSTm
ROsvRFpxEbDPCoRsv0mv4DhXOM86dNc7apVyQroiQdmKA1mzMYq5+w6i6BC3gzZoQtEm85YcGVKD
lHxGv4Wsgxm4so6kBNZLJyoGK8j4vlYumb83DbbDLwGHONi/jxcJLYnR8AA/7k0pHna0ks7G30fm
ENJSsR/0KImBy+J5tXWSOd0DAWnQh5YcgMwMtZAxJn8h1rEnRtYlSTwyRhHGlWcpLXivj0v6WogP
AF4nVYVUUolmMQHAvmr8/bgdJR7L28dGJVSaGK+N7KWCA6H2sVUT5s/ech6jGOxJ6J8uDQiQnDRs
+z3eUTd16rsZSgD+VsDuewigDHmB1gYdjFTmeD+rZNN2zkLPzrxEfF3gxu+Wejx3MlOtDyYma/ov
/oqY5egMbW8UR+TD8HUEec5x53fDk5mbzZR0pROlJcTUln5zo/97RSm3WjREg0JZtuFlw1/IYo0n
weXhcrD20dMl8H+CYc6H3EZHl75XMpT5aMCMaiIGqqGGGUqtuEez+uLa7g9O30teYk2GwN737Sw2
NFfk5Ds9ehzwyhHDzxRz/ioUnYD7Jkhaxrn4zbZ4F2GdBVIekfvH33cuD9VWd00LwTEESP1ggXiY
CwwtG0HwbWV4YxXHVvR0KV/XpIz47m9+AYkNdaKuaLu0s81K/FWCXv4lL/gGHx8i6JMZHPi7Cjvy
WnjQVTkIAOsnjOVLiANKmFaADbrq9bn4RC0ml63zOBg2F055nj0PW4H3z5phDz/c58c9OctbRPn3
PPrWyuRdyOeItCFO05fzR+/i2KICoQJHl1AQ5SlD3WHcaRHy/8CZCM4TXZdAWS1h5jT0FuII8hQH
scy2CbqJ4DpyDLncza71T2qdWJ/QDhAsRTS0y9XNC9dGlDE3kTfZAqHaU0hcbQXMkgtUT1DGz9vx
IlIfPQH8IOq0PUB23mtJCHD0z7AHFAp83EfeRfrx31z+tIjJxKx2KwMRxnyqonbiUTz7Mmb0aZQM
7YwXAUfOQnevIbf6H5/rBu6cDVAl358GlbYXTGa2GX0OBXhHJevBetgP+NynAGN290meSCZwMjTz
rSBT2bpIGDHGz25ESX7ycTQNSlC1H4Q1R8T7Bv9jjbCdSCEX/rWUcHQ17TlQFNdTvUaG1ErBPfVa
j5xMppO5/ZJVAL6rkP9+hEjWCfptx2RXgYv//dNSB5Y9EX7AXCwNtkccURzcZdhKp4khuXqTvj7y
SWiy3giHZlSKZO8MjiwuG9c+WtSTeI6CTVpCy26JnJ+Whx/+vYI5LBFCpjtEAJBup0d16TwKFiIm
J9f/kOZ0Go8tEhOjBhc/iDtNScmnsQiXP4z6MQ2bu66+UNoe6iXEZ/Vj3p4NVmxyBSZBB11UXMfq
b/SZI+70rCXmUmH9LagYGgXKCy3v5U4TyJgpfS5+WgggRRL8ZJoWOpZsnuf6vXyH4IzDIOMKwz9J
KPEF/iaEDCuOjZDMCQJ3JpULyWaSedSmf+Xmmaq0jVqsqFyUeey8QgLwOfpQqltx9lfemKgnuqgq
RvR40/OZguSSba4gZVahcTx15adGX5gLZ/Nns9tlkZ9lJAR1CWuGeSygcpzqv71jP2B1NlHLJYbX
ZG6I0yqCvY5cUBu2eCyywWxR1w1lR5EnK2Kpbcv0/DXoFEutp5XQkrJzVw8k69fK6pAJsg0XlJbd
W7LRFrU6yu8K2/+Ev+ywBzZYx53OIDcFwiJuUHF3o2M273udnhiuQFjGoeInJgFlOUSp05utO8eO
03QMqUKlBK8oIU1xD9sN5qxdbM5OhBHQCKiUKJTIGrhFqqR9oDVYNdhGySmnim3ykpu5qmXqDq3/
QcNlJONNc/rYOF2iEYZUAEkMAZtKdnHMD5NIBbTHcm6tFPn0Oz8XinUl/O4484eiSjndGTQJ3ABA
uv19phx1G5yQP6tWIRLu4ZdnvplIGgLFf8hgQWK3ffKUQfGAOXGpwIqWaAgJqBUKpuuHa99SMyt3
Cpfzvg9ro+uLJw9UkqkUqYX/Lk8JDSFQTrz9z2jT/F7P0w7/V1w92qOaInlTt3lPUC6f7Qcuji4j
jRQ9NwZrgYL3JcRwZ8zFvj6Wm4v9NMeft7MpgWEjkQWeb3x2hWpInaJEp8Di1vO2nNyr1LzhVoCp
CKRJyveUgyOoxs9QSbflR96d7nbFm7RdsXZbZov+mbTw7Jx93pu/SMD/zfnLTrpfyQ345g9NZa0K
qnCm8/TwLGOwLzLEa+GHb7D7c+0jULJJe7uoU0Hz5JRcxxBApiCXNRYlBP5otvOLg4L4Iv9pPQkP
9Lb85NGtlWDS7nSXsgz0jRCVu76j6etph4C5Cpkdjs3h2GUu+Mcrt1vKMqlTiowpCvMIFKAFgODw
AQsT3wyb4+mVp7GsL9tplifdUypAsgtEuKM3FmSbdSjrIwmEmxNRmtaL8eyk0Mp6brSJHyGkjGa0
PG3Lb/oPUw6gD1NuxNbONRpZt0ug30eaIg/L41nixVZc7N1xU+DMoEglkgZOMs5csnzDjsDEMTS5
Arw/UASqyZ1LMGbDuRCW674jd3YRn4tXdLONHZsD5SJMqJIbvLmjQTPinrcCtAA27EDujz8RGMtG
77fczGFjcg+POJbcnpJn2Hy/ZFS2IX67+Ocr0QxAdZLx2XfPse1DRHZe8kcwMhV/Vt7W/d/NPjYv
3O5W9GIHweerHPrxnK5QEgADaxkJLEJgNdeOG8TJT6bWv1Ao8loWNJ7Qx8OAMZEogZacUjqa1Htr
dMQHt9K5o+lFoe7TaLCfEqsB9qTf+mC1wa+VS+fsng2W4qMmbu1DDhqltANfpiiJCaMrjcu8D/NW
bbNeQaqgBISjYMM9ELC1j+8xAPmWHouPNZSFGBMdmyhV2DIj7IZAxxGYfSQulgFKEGgRedzyxpAE
39HEBWPlOcq2GdpeLuQiDfzV+WBNKZanXkpr98nMP6pi+0sflNa1p12aIz/Ga8MM6OuQSnXuCxMz
ny7a5K5lbaGL8owEgmAkWTUBcU1Z80Cgvre4U3D5n3GUSQnONQLu/ysqbtW4/u8FM0xykuT1jVr8
qouoIYS+0HaYe5eZKFy8H2HVNY2jlcI/mkaegXVRyp191BHkR8aX8YEmJ1BX0SCPy5YZ0d/ce3lC
9zZL6jdjux27EL+VQNEqE83hqdWyLWX0oRzgBzZgEYdL2EKI6t4j1HN9Q3FOhTfFtUXrQXvaMDFX
/o608bjXXUrEYUEvq5/UfS1jE0VqVa3q8xDmpCihwvVfOpDQqO1/5JOq5W4pD20+OYfCF+5HDOXK
BoORBNK5u53yckNC6vRjDQzVYh8qIMIHZASVEP1lUWx7OEcxZ6Y+5QdtNPFqkPQjETFpnIQ3GvCJ
fEYGCHXjmSWyCWKVKpvVPdt87y3fAPM4uTK8izNHuI2z1RObpCYXUqbUudG7L+rZCpEjQjvCqoST
fxmpXpjBTqhg2QWynuyw6xGcjlYJtO4AeJtRSpKHyXcFD3UAOncAW8GALukzfJz4wb0A266MrqmR
iV/z5NkI13Sw7JwHDRpeL7gr8k/SA2uE59NEkjtR011q2T0MIw3MXtTPlLmbeapT/pQuNfsr5fqx
DEDD6fHgxCgxkMrvqjylXEiKMTfaUIcJ2blkaOOKn4m3e5iQfmkNOAVE/3NC97GBWKu8FT5SF2LO
OR5TWUI0xw6u9ch5SWPa5v8scCIoWjrfeiVkDZ0OD9d23qMLb/pyOKUCJdTanjE+GlsXjdbDCYMm
QJQfhDzf1RWjGLHTx2Umt6MR5O2qhWJLNOhI+aknX28trN5rnSt9MlYoAj03Pk90zoY/eOjGqxCC
gkiWXU2krCkefffpZAI8DJ5r5fIfLmXAmFCo5HHEdGRjqHKOG20szrQBVFEVciPBp//0zrbeyD5y
ISdlDJIuo59gnTdQHLZ5xm3VSu5caOiJRmt1wZQXYhQ0T0TzlJZQGER3WHNOAl57bnjP7DWjcsh6
6X5qagS/HhlaRXPvnt9/YQ8ZxTOGuFA5WAPzrGZbyQlVgE6/Sa+xb5uMDG+QNY75OuwrE4/ftAsL
7dWT8VoVSbcC3jHmAzrQr+ldLr8huc82GtRdrcppFyg0ywwtE+DG4kdaQOEYKw3duxW3LJKY1+kF
fpvAIIfMrbCrmr5oo1kcCh4UjbzlvsaL6SZWnKrBhPtnyRRZWD3acKnG1u9AhIzMuvkZA5XeXUfn
huCyIsFKF2vJdW4pqSWgzMk/jBjHaOzuORmZl6h+lPtJGMjQ6I5tZxIz4E0yGW8aJlmY2bIFjOhp
C5tx/2UdMK1jMwgeoKBJwyd5MzEdA6B//CmKVMxSKZVtwd/CBcb/+Qwv307j6mszrIos7Ad7iqjo
9R7Uyv5ZZZLpiIv6W/XDzYB/+bcCQUYHUO85/OZel7Wu4S6+qN4+M/GXmuUyoBR4Oqs1esnm4uJB
JmM8bK0p5G9bKC38KIWOSAxl+nrpCFQcctuNwPaTKvV6AjowfwXq+qlp1cQZOKFGsO+SG0/YPKFr
xzVL6gyoPMKR2f3BcqCspdAb38SFt8VNgxVznTP3TCmbK3y3dF3JO8961L6wOHy3LAeIfTqwtiTK
jm52DCBammtwqnskqNPtAIbivPKD0F05zItK0GqIzJ1ZCkzvSzPz0SR4y+Yp8WTuSyZ49Hi/goVG
+8Sd++DoZR+N4uNrR3hk5ywF7rW85POYTDNHq4iBb4iN4XOIMP0Gz25AQUk1BTQY3RYeAzngMp/b
g+07U99IA0JHT2nkzYji1AKykR4oLAPhqhts3Jaac31KfwVF1RRNNiS6zVYG+oJdC0kDMjNWge0y
I0fsr/0DktOiaYTYd+N6yvaloY1SudctpqUO5iptg6jYBklX3hlPyK1pB1xFYJ3ZFSMSdbfKV+2o
N2bOWJtwpIsUFvGF51h2q4X7eyiaCyJB6zRne41/LtASOUNol62OuVo4g1IrY+oRECV6LvhqazsQ
3a7qhgFVJ3xTSWUmdkgwyLsvMJuFhj5yzzGbd4Utubzus7udRFPsLIf76/WbzqK37lq72PN/he4I
4qn4F7vVmLy09ptg87pF7PmYnaKQWSBSYgPIZBLecJs4mqivVKOl8VUNe074pMzctKyCZcl/6CHG
WiVNu8t9Xk196ftny5995taOlGfMmJnJGim0k+SvmoGjT/AANCbu5ayRXGyVossQIwZA6TmA36Fp
ByHztACxqszVZrbxa7hsXNInJmntaHqMhHq3EvHDFaguWih9CSlhkO3ByxsCUA3bz378v/Ygnwpz
UcyvN6uUuIS0Jt9i0o50e0EXRzaORFWFCZfPEc0RAcBSs7kp0Ba3rQsuJJTgeS6Xm/AmlBZmwqHm
WVViECplTWs34INBXRHpnYrJB4jZbpeB/T95knM1tdxtSspjidVA+ilmW8x/H6Foj+XCupMBmHeS
+tWtwDm3ag4V3vV8Rz94KcHAnkn4JFbdFosR3ywsSYpO99r4YkNuvW3oBxSUK0OHuAr3k2t8BaqO
SS4ZLKCEPLsUBxvOyBlBSqffD0WQke5QhmyRAIj+JU9JNhAZFyHnZaTkX9vluolUOEtOVYj5wDbA
ICpNKMayEbIkEWJg0qOnGMmUkgyUopVynAK+z2LmsLZtQ0k/vaXswZTs4c/pOLp5CxPrWQ6YnLXh
TxOm6H72foyZW8PFZNg7gUKOqVoKPmQkXNhr53u+P/smdbVAFTi6DLDxrYNclYNtfteJGX2wRZuv
83PcrFKc9HtJHsl3xYcBg5ieaRdtbuiP5tKCVGU5+zyjqDbVeehYdeR0QatpOFLATKCCVvRwaU7e
qGSBKuJFGiVTA18LIHQvwVRchZ0EWdig1TH6ZrRrnv9PqMwcCsH+pbjl+skV+5TxY265c4Vt6oAj
rX/4yiAd8yNw15O3qIZNqI5nPlVBrds+tGSfUSPKW+S9dhOsdKRvEatRMVvidR3hTftqmqqifgAe
xDlvu08w2P6oxvANOYsw00LbEAoNZ2BuKhrdDXAvYI1XcfAWBHzFXDmmCCqUwIenE9oEb3KBq/O3
/tS/tqhmT1oIOipCawlQ33t14pIwwgh3xTIMimV2mljkkV5my3wgnn126KoexmJyBUCgWn/J3dXR
CQ3vgKwp+kxG7VXeH1DAB53ggNI11rP8N1xxvtZx/Xu1lBA9dJiteW1+oWuFd8Fvyr6KT2rzcBfF
XguXSujLhciRkoNlM9rKSmb+jXJZs4NL19TTLUcs/+S1SpUCikyx2skVn7Q2coB63kYDXwsKmuHZ
bM8tA25GiKN5rlZh9BpM2N9Q3mPta8fZGbFug3+rzte5W+kGPVq8c/4MxYqJDYZEmzggnXzArbTK
+DD2CpaV8CowQzjFVcPAnVCB5MJ44NH65M0wJV8O//6lbEfoMrueL1yQjfkmjk+/bs0tbrLwUbDV
Wquf6hDnZvfkBD5eWjZ3t+XfOkyYuk4nIhEOGMbZkc6RQnoceVYbp4/MuBb4r+n4HiNuMLvhScGx
CqdPsZrB0EepGo7WGAimvM3fEZwA68i4hQyaPI8f3B59/H2EzvEgSdidBcPSb03u+8hIaIEBlzcD
Mf+LCRSZZ9j5UoRPU+zxRlmPUISMkiI4t2n4g3DlCZINWSsAr4jWD6Ic9JsHeosWPzAxUys/liiL
3OOP9zJABq7u3pmWvcCENVkrE3NveuIo9Vi9ebi+7Sw/svX8eCABayulXPSZFq9+hSFwtDB8Tvmr
sZPwy8k3HRvszWaWvB15ZYW2Vb/Gj63GNL67QqL6OUfNPagOCd98z2tt9uRr4PaATeVejo1ylXU3
TkzuvLu8qld7wHVaXklnLe1SSzsuzMAqAKJY+RVBT7FwxicqppM0iYDfk9QwhXQ5bTvcc4tnqK33
UzhfBA4Wd253/LHkXcL6UQoOAxdrm77vrlnrHevuSQZ4CUO8B4REOT8vxAhAJKPgX4+2IgidXHU/
ejcMoD/b0oafca8BnWHmLUtIkBC0DZnZaqQZTsgHB9ABPlaT4hG3hjnsiuQP6yGIoWnWhWa5GjpM
FJPgbirffxOKmJvPZw62BkRfGzDRSUEg5Wz9dQC0QXy5XquK3OwAPN0Qw1cbq4rylbZOjumY6TYm
xYpsam7N14cntVP1C5u+/rrcZGEF6chUBIJ+i5JDXy3KB7Od8A86CMlXu0yf7FMNjDmkt/QvJW9p
MqwJAvkF87bZxn0bMg6klTZxxEbUn1LqetbYk5zEb1txNHKKinVAUxyEC6eLHih0TcttIktwXF9/
1edDZt8lipdFjMade5Xt+22BhoWhRDAD6CW2IgLb8yUBkyBp9PT7snS65LJVpaceuirrnS8DD3zS
60cHJr8KCKYurHvm39PdsklWxAobZ1vbBT4PNQkJ+0uj2d8JFMaj1s47DBDVfkAbCTvcsV0AMBlM
M+ynK4EfnlAgXE3jmMpf9Yfoq497036RPUChK2ndgXFGYtMTZXSbKEoSLDS86srt/EgSdAoIL6ws
waux3kh6KlvtczGvJTb/9jiZPy3Txv7oT21u2j5zKrg+/r+eA2aWYyU7u3Tkqcd0K2O0cSXCbttK
e9nQsYWJF6wARfV5y2x3CBMvSd3+ml2d4hVFlhfYnoGMR/htI5Q3OlfYyPhE0zj6GxCmINwoKBC9
MHlB69apO2mlaaCqMpRBInJ25khGCnGWb+FrG3CHeKFLciy7ev0hnh1BSCVlmeg6QgdJbIOarAWM
QL7fW6quGNSzPc7h3b0kfI34aBe3IwI0UQlRyyPKYL4+/wyvSA4gQgcbCg+/4mFLCP7z5MrygeGq
GOtPorNU+AA+yieg0HpiDcau/1roEFbzWjplUbY6aucSijpnAbMitHoptqCAnTbvsnMlf5B26Nwx
LykP5dO36fKB/2T2xKMMBwsSysraw8cFR9+BdMsNUfLf8yL/nEt/+PKM8i3tS3FOK8A+Gj+0eckZ
RMSXL2u7A+001nXiAs3kuBxjBh775Am4rUQurTS7QHTCI55B5L8Jo1XfYJTKR8ujpGtgUf2VhVvf
SxE9xgBMsNHPTdKL5WFJPMSrYuSFB9SB2hMQojoAGUrIsTC6FYRNoOFwSuLJYCY7lecIiI6tVFRJ
kMsM8dwZibTYWDvjeVKLDSaSdI37757mpLrgpPeKz3v0+LvMbKQzKG3RpInSpzpWeXTTgjK+V1zk
P5YB6DinefzLlYN0FIOH/peLRHRDmQrh/pQUCqvNzW5IhTP6JI92ckJPM5l5NzatOHen+fgma2aW
OlYp3Wn1RHHcnk12G1mUGCLoRhWVhrf7P3HIincarl1yPOOnx/sShJ1nWO5OXIWE3bLUf8Pid90c
tD4zrblaFyjGkgnRK62jGWxAZbC1iOB9vGdsqO8zcN6MQxvHbGAs2zJxEN6ctiFO6dEFdCQWwEkJ
5LhqysBqqI5u+Akqb5JiCKeYpBkMaIq8myb4Ima9yd5QhfvgYcNhk+yz5tNo6iWK8xE+jr79ZkCj
zRJCL4fOsqAd73Kmhg7pcfuw7V0SnwKY45aRRF/AFYYk4y4ob1T49IqG+Iq7k3vKufixv9zQmG80
aPLdCbLMzedCs+zwBoDbJ42Vq0/4m/5R+8O4ceTqAOdY2SLZtAGDJTS2e0B72sZtvfAiQ886xjNp
KVpjRHc1BxDkybvW/RVTRdu1ufbHh4uZsZyex1WHdxARxA7N/7f7jgHVNOvVQQMpQyxoXNIMJIUU
WJTF7LRHNyaTl8Lsb+W/bfNlD/2oo1MrYYh454MyZSpiucm9M3Uq70cB32zhjV5ZAESqBk0c6wm7
rK5/0ZA3jYAJG/Bo3zZDGNTmM2q/yuz7hCy+FsgZA2+PvOZSnGocAVZsqWibhun2awJOPoKjtsOu
xEv04CFk/VEk/UL5Q5eyho20RVKMZLonMpdPhRKQzeMyoufC8Ajgfcu2ka9PyubAaz7M4C6nclci
+6sefp75d6i08KAeYozy2TdpJhqtXcQ1g5/zZd+Lo2c4krFm6woqjUz0NBGEuYbM7vdVZLbuQ/HB
6TU7WQCH3Oz6we7fEqrgn0FCyAtOaZ70vowIJpJjPe6Sm0CGExwpswzgCHENHBLfibQUpoHVKy5Q
22xHJW7rK2vwTiWRFpgFOfX0OHXp8T1pycz+uk2Dhz2wnAt22zacCPeuBcJ2dmgoT/jbl7SDVK1S
zsutd9lq5Z5D5jvmr5W0k2CP+RXaxP1jpoLOrkp3hLvwZmf27cRbexGcR12PH3lZ9gcoNY3ArQpi
ZeG6vCELxidUBEGnNyhe1oG7PMwBtzOzArVIvZ8C3Mx477+QXe1LS3/Dpk8AZey74C58Gfeu5cW6
cBSHR0dGj07+atYErs012XSLkD+y3Nddu2t3f5jyzJ19vxONguLQPxNDeCakYzG+uy8w2b8i417c
xW5kJAd6RRo+6SKbHs4Gi6Pw2h95KaTDHUcBeeM/AGLHW96SfzuR2kD0B528B0o0vXssW5dYaEoC
zR17a1tCFwrZD7YHMXR9fzjyCQktGO2OkfrahNSs/Zy71YasZsYZzo5keYsN3Nf2f0ZcTIi12Af3
1Vzm9oSRwgA6NBmF2SGcfAHjXlj2vvEXMzJsDVdkoTBc2afI7Ae+VSz1JE3sbjI7l8oL8UA5YKvw
lLicCWE4uUwGF9evd/6ZQFrRQ7/uvLefqqSDpnXOEsjXdg9cg/0TpCTN8mkAE1t4ssOy0Js0otmz
b3+4chxyGD4CbaVo09TMMR/fRip5ju0CGpLNTz20s0tqmMtE+qYEqDrGXCYFHGSso1o2xdjHAego
l6B645DRbb7i7cLWyJEok5Og5IWb6LOpLwtT9xW2ojKPFMb12xPd2rTWGg7KODje3M/1CyKhvHYW
nGXajUcsI6Qa5+s5SpRc2paGXvupEOLSNcxHOEtFw8yuWBVn4Kl3JX2gHArVYOqtfVOJs9uVpO0z
tJV2zvpEiOnfbDBzyJfxdoWBwTk9Lnkm+zT+jHvMHmPVCeweFd9WXDVmLmfgrdSeTrFiK6jiu5rF
IpTeJHQ+qZcWzPibR8F6dQc7KjDmIlLO/tiiiDarsvQMmMKRMP6QgO6utfUpN90FNzdZPYPdYned
Ii2qm7RiZLsLZhCYAdJbD2xRijv2iJE9GqpNrhyW6R1YkvZ5EvJnZdWavzZgiSKbJTOdLgQdH6xe
NDn7ea3TiN/Kr9F/8b6Ybb7ltIY4iP3yF34IIm72ZZSc5Ul43QFMe4sag1R1AF5vbWPaw06Bv4hR
1Jd7vnKmH2yhWRYqBRnXn48Lc5m05AYQOH2L3v/n44MkSSddZ/0ryjR32jApsx8EZpAtyhE+gwgd
FHPEoAYZGjjfzeMqlFVT++3NP5bVxhBwJo4IeWxE2TG7dp1vWmjyyO66J/IT/SrZH4ddqhblgovc
pcVv7806zP6IL54UrXA8Ov56D+1kGiPJrJRh1aiKgKYapXLTj95BVkgsJdzpymCqMcHAX3jlujnB
2Ijv0SCjXgYqySt40uGcSjKaFWsQzUfwdhaImc0SJ+btqeTFQqETrf/h3l2kETNnsXh+HYS2LrmE
TysVim6P7eTHHbBkKgfrrFxoev/PBj5vS1eyADfD7XzD/T4moM0dhXnPgTikUVp8XRhjcYPkpnl1
iI9QrzUtyh0Gh14bAmOrVcaZ629uNfZ/kQdd8OJYD/HZVgHKmPJOteYBctCjZkYRKcOn5DR7rYT0
x3V4OoGkwOKQ+W/lWYnB2tyxNKq05u/4ybLEmNFSHvTENzI1v6CCdfjG/n5U6JJRvZFLdj+WxNsi
rkuKBfoqkLjWkYyHlRckeceoi6QuK9eVE6ptSEk0FNHpiesWXlPudZU5S2M+b5tbCk3uAToGVIgX
Jjq7uhix0M00zBFLQJmVf0ckClZSdXL5qEDuaLr+/l4KDic78k2lD53KKCRQjFKdVjnO0rm2GtKF
Q2JeopG9SGi4Ym8eHUo26EwSi2Og73411+EfuQhIzmN38anWa4tdwjwzbtSynnW8XrL0d3WAeigd
UNyqs8WS4uTUM5XY0CKgIyX55oz4ilYza+WCMC84SWSYfVgj7lIe3d02FKDq3mqrZ3O5OIjDHqsc
vrpc57F/pqEjlOljLy88z9xRbvclMWolCGvGzUtMuNaV2CrGyWXQzRYG6480dVJcmukwqrwDCU3y
n172ps79XZHsdozlDTSfTwrToU6mhqPaASvHOEuNNy986srCPi+6APlmdCLptgiEd+2O4B28Edct
SVTp6SpStMPK/GEWufnZ1KY1toTTaACqZs77tae42jj3Cg5qBz70wyXSAKuh3xex1CPVBCeFPyD9
SAJFOnBTGuYcd2ct9s3aRddPwJktSCHyB856R6lNPoCkp488mM6Dv/RJ4K18z23y4msLSBOvTQsH
VuE/HGCnTIZAPk2IkvdT9A/Y31ADbKvPsViCbmL9oJ/S3ZPMNfD8NiAwH1lyfsFiwEoVejOIOBaO
9WVuWHkEI3vfyc1K8K717KGJ2cCWBOy2YMaqRX/yLncwHSqNSIfF6DRx5ssY2ctasBLcUGEZkpXI
rYBc7y1GMxy/Vikk7SyOiJUDsAlnbfSdVkNUEM/50WvQB4oSHw3M4NJrYGaItMMalyYwBsRDgjU5
59tRGwVpXLP9K0715UETnCivOvfYeiBB7QM2Yaun99YScX9onph5Y0UuO/KW9ghaFyjz5FD6Mnih
4Ify/YviMVfmayMKT4VmQZZYTvOhKzwMYYYrn7ailcQaMeLmDLuJYK9jC9x6ssCXrEIKiIZ+0oJy
SI7BOmMHdrAUz6+sY2ZU+mBd9IJPNsxv4Mz1JEepONrR4L5XoPhGSpjBehL90PHfVB+QxQ/4L7Yk
/iEZZHOSOODlGwqCa+x9Cf6l4CxLL1C0MNJ2JlhgxoQL6JGYM9RBzAScuXptk79HsXG0I1uc3Cr6
rd4DfCp8Ry2Jvho8nV1iMmQ02G2Vfir6f/pTQRzrrp0tpRY/bwLApHLMSRxeR6HxCoPwHtZNR/Su
//AZJrznDqTBRTtN9Q2Y1R0ubPMriJW5O9A+PlNe1dTdOgUIkBVWietf+3VFcSMxD7T1hbW/0Tlr
b2W1j5tclIepH0oodIPHRtg60np03ThIIeRyaRRklUoE0NcnAZWlc9rmS18+WDVRQmm1gl2uBLMO
r2gp/r89BbOvnk6jq7Zt4gSjVO+SmcbOLqljGc54oFwT8nGoePhU2m98dVy5pPxvk4ccs9rXOlS5
VNuKCelCVnMPoNs0R1oWHm3Aumh15nKirUHNscIl3sRXYLIHecvjl0J+MigewuuNwmHVmPC+9dgB
aqMGop8StrFybq5IUl7hVKaBFWz3vBKcMa+PF8hU5rKwYdM65HsqaaZWQiht0MKUnfcnfVX1OGiz
6JlpwNvhARcGisHJxVKFwPqrkt2/cXzBSlDciRdBTGfAcKKcWAl/qhmNU0ZVDz2UazQf1ZJEj6u4
hoEgzMTFncvZhp5OQ58CE59IAGn4xhqu2jAY6dcJtKp1kBu2bK4YzgSB7IMrDGL36ocyK6hegQhZ
EOqO69LRWtukhK34VRw+Ahch0vAX877zl/XaxMNdJV0y9tGYjNXQ/7LeDyeevtzGz2Kaa7P89GAd
iMoECBM0wimkKnYMY40wU+j6E6NXNCF7Wf+2qtZExSq7gTqD0orReWtlBE6g14FOr/OtwYLAeU5o
ya6TcYMXLV0Zr53jQnML2bSKUjzjgmC6RyyEECevoAkzoKdi+mwlXQfQpkZ6tIV6m5QfQfsXKs7a
Jc/xgQSbBJS2KNDRpFqllIgIb4T5cMkeeyzBpUCFJiykvMnGpDfBOsOOsDsHDdNyWzYXWX5LrEoh
Fsh/l5DPsfESxp/GVbYk2WD5B/nGHG/7nXMpm5KYwH5nMlbjum0z8s9xhQpuj4jGJCHoUKtdr/vw
IAbQr8Kj5M1gVLd0sL3b/pTn+qowDivaZ9to3ubWkYXZ/aWOy1tTOFWkF9z027KQKX1PRXCRHDRc
x9UZaZMqVStXAsV+QfsmOJFWyCWEiapDseZWbYQX3fnWWbWwIcnmck4ydFl7hlGKNGepjZTOldio
E+pGKN+hOCw+57aHXW9tqeB3i5aaqluIhvinTpb1NWAMlGGvvE3PozbwnH5ODgpNIE8mE71s3Fch
Cs9iF5sw/HU52/UgHxa/7SQePw0sJvbHY5HlKoI0Vzb6F5JNFyElTLnAVjnRCUi5GoyV+oPlQXMg
CApyYyrxrN2NUT3KXnoABPStoj1LAGTak3vqZWaXCGSkCsvXhyHkRniXVkdE3hYFoycnjbR9GYrU
fU4JeBcgsKagDvPxwYspMfILw/yEPMqWuQ7I7rzVA76BoYSJO6dLRYLbBDzMbFsoDa0gt7PT4hvc
8LYigUmjJ5IzGAyZn4HoqXKToVnKtSBycZG+HvSYCEYtzWssap0jj6sIecXNILvKtlJlPJkeHcz6
rU9RJi+sjFnxtSLFIVcDGxIekebBscN1IdVjUK7QQTIHcHuSTwRFIIN01esi3BbEQHTD1TtWgHZW
/ak81THG0hdGVwsVJYpYOKdpNQfFRemoXI4xqtCxlavhfMrcW6RFKZb7U/b1GwHlAm9/xccnVRS4
TUCDUPGPUf1fj75vz9HpTV859seybHz2EyvleQ7hl2l83pDCiu3KOhYtIU67kZcc/bKDfnT8H7SL
mnVqrBj4522TaBwhed83ivnhW+1F/WyEJJcjF/hPGzv97L6sA2VtDIbZ2LX1j8UU/n78IRZkqtH3
8KmvCrDY5zcgPCh3KW7M7+a1weJeb8A2JvA9p8Psw8zVp1mke1/Elff8zAQ41YmCoKQfpjQlHlA1
2kpp0gvflF51eWoVGXB3WEOamrcew2SJLb8rgeMX6CLVHj74Q8W4zdh6Jgx+Hi0YoKlqvsVxg4LW
Tuol4fUpmDaC6kGzJqxAveq4CajFi3PAvWop+Qr05FLVxg4oYok5FjEupYiGK+f6svLqQltmBj01
wPfDqSPg4DXq6hDC7RqZiRv+i73hQreobCRD8zXWaiRpU9W78np0jevq6MelP5m2o0M0WXmWxAGA
1+eHPpk6hNonILQxePOebXUXnKdyE4+5z3EykoAM17htlFLFF+ekyfdnvbtfPn6HsSs1jfdTc8AI
O0eANbYNJdT4xb0ts/hKl0VDvanW/qjuwQUIWu/2iYqGvH/6ResdQNuF0MkGf6dY0HEulg8jIjgQ
NdMrGShgcvJKEFHkrv6mpmvLdljF9DB+9wC4r9FeMlXW4CNHoIkXNAQOGwGJqoIsvqOT6zFZoxNY
j1G3ES/LTq+eSLbn6taR5QYEFfzc9ABIblpQGblRCav7YsE7gJU8tQ6QFBILObvGmsO0cA6WDdr2
UCTeOLLct5P+7VTPzNQY87PgbZOkc8o+4QQRZ4pJOxCv8CQ5rN2GNB46hH92Z+RLbRhkmb90mm8S
REe+ddwRUnzlP1sEhIwMn2chqO2woe8sWQzH7/Ong/UXpJs5Lclg/3PprcBtfY/rRaV9X5KjiYr0
YS85GYmNeqPAU4jHiKr/FB4gASnAavoM0wQpWP7MHdacGwcKXAjEncBZ+plnGEu4ncYbz/liIRup
aji2j1Nn8JT61gl80FZTLD4lo8/mSiIvScn9Ac6L8fcfnQoWpAFmbn/crhgwd1ZlCr7eHjiHCYfo
lcrsuRpePZtZYxuKv9+DVmNuT5KJAC1FWYsMftHx6Nkne/OTbtE78ltiTKBOKlmFGTnc9owjkDBQ
puQ8DlLBsJzf732kU7Hicab84+zhgBsyw+6MWXa2ZmqTzZrfw2LFdYsG7YxCPUXPtTL2PVIBJ8Zd
+XTNeabDu1AfDxE+MD5CP3ec3VKwt6G55CPdVZ8Sh001KS+aqL/bA2lEVwl3B/6iqRqjtJV2pZpu
sTVsViB4283OoWU7fyw+XQaoHTvVT9owlVQ7bs8S5ajpj0bVy90qz1oOJqUOmTvbFhHMY5SsNUUN
P+br96PCntdDUCOqJzIIaKgOY3DCgz6UpnGQ3EPJw+wFGU3qZOGM3uS6TAcw+BBmnvNEXJD/XZd9
9BeQgUWXpGZakm67ztgaowhETd4+7ZEOVKiANr3JJnIOzzp1xlkL2+7ot35MSzNfqctAXeWbIoCU
D7QyZwMUxk22NQ6o15HMv70VvFbbj1N8GhNA6gDLcBPvYjMVyxSKpCuwHVSCpcWpBZa/8pThFyXP
NaZdrkvDKGqZERVeYjaWUecVOik+SEJW80Ys68AFMyBDL59ZUCEOzZ/yr/mO6QjYIMG0axDVA90F
CNSLmCC6jFCDSLmBSE8nk0YnI6KhaxRKIPGLJsyw1PFfXbUdtG5V2ueLTw6Uc11rkGos4ISXPoEv
zT+eEiW1HmgPMd+Bl0KMbt+OamkQ2BralBIIjLGH9gjwX7bQTQZV/Ez2L1unguAfkuugzV9T3NjV
ETyt0+PnKGjzhKhjWz/NGF/WL6G8HB28XQCoSLZUfGn0V/OLe+y7t0a0Bjjm+EoRBDPiLgxaHTqg
mDomoWvZXXtgBr7Yvtui4LfZ0QHE/3NLEpgozNiRCp6OJSfTDpV3VXPr6idRgwALlnVa57CyqKJc
dmJYkDXvOgRE34SfKVIYkAJp4NaLdp/BXte1ypPmZgQjctWmktLT9JTTraN5Z2SAae6fuqGQVWco
84uzrOlqrBbtgzJYxVEnAFLXBNhBdNVgKF51NRCrz53/nYchjLcfC+rMbR5qIUTjkxm9jKxcycQV
cJYU8RvGYAdREhPfiCj2DTXFFZ+bDwJQaOTp7ntz1yqjyOLeGuVky7S1tOIOxHlU5aFbTi2OTDjK
w6fr2VOOFFcSxJi25YxWr6pSQASRjhqoRmsfrnQg1Ghnty/n2jz7VM/uWDlQFPE8QW4GZHZGaKxZ
zL44HcNY9ln+dqCvhUeqspgfElxYVsjYjFnSJCR1pxTggOuflI8RME0I7+Q3f839L7pHaubD2XTj
D1+hQsYFTTHMFhFELbWfEnh2l2Huc4DMBfAv8zBjwi5Yz6HPLycIrE2i9i9+AXprXERLKzzvUvoT
577/y8BOkRG0qdsxgRwpTxjQqE6j8I6FB1j60nSKHFZ96SwbVrf+sk7fKmEYrqDmyKoddeDob0ZY
3XbZD1/MsZlisR7B5x1+50CP4/KJFyunVQcj6mrxTpenoHxJHV3eHL92mIDTrGHHqpxYZZCHfowL
hEySWtSLuz/TEuYmvtwF70KA/cTvK8z2dagwJunxjC2BSgcl/c3jwy6qF8Qi2M4ahPyFMkAnej3W
zSP/+GKPCRH3EczC03v8cLSHNOjroyzqvWwTICgkB7ZHAl8N/m4KyLlyqu1c4Pm6MSriuVQVsrkc
DLEU0jkPhxDYCYRwZyPojErBxgdtuzyTI4P4nD2fcMzugxd3C9TxZQrtLuaQ8eBr2SyISKAf/G8U
fPxXESeXzC6qiazFNdSTUUA67aGaGfK/AS6l5LV/DdJVbzO8b5jgCJ1ofn1N1EgLKMOQNbZMURa8
xXjEcQM9fHIB0y9TsXVzfIvfxJdBPH8u1vzZA/k8IfRmQip7fve91yCWxyWJ6znoMAdhZ/TVk/Gg
HsX0sNu9+qcCDs48QOcLhpJ1+F+j5RAXyfRXAgzoFoK3fos2roidRUWJX4euEclgbXVRZrfEvqzC
dB5LhEXiL2tWpfbTt8ARH4QBAMGmXWGQu5m+VWspjBV25/E2kchas0JuRnr0D/BR5mStV7hEbqTE
eLc7Fyxf+1i/qv4qSM0YX5hnFqSDBFq808MxLA9XzQX7bxffuAeOzNeiQlIQUFzZtIwtkA7qmD5V
5RJvKL+DXS7KTi/mVehK+LuSFnMJYNK1vnuJ08xVzhYh3ecPoahLNCAYmqUJ55yyeOPxcPYFxZU2
m/eDoasnnHlU/lm+MQNF9YQqLPlU8AxZw2QS9HFau3kov3krODU0HNdv6yMznRmzHi7bAyPfNq5I
d0zymHyE8vwXfJVTWHP6pFtWmogJHujhDnoEvHxg+J+lkPvDC0A6yEzS2QUtZqaNeHgdOQmU6RLp
MO2J2ElD2oKmzbT5tXnWEimvdeRF3E4HAhgYH0NgIf0t6rQ44kk5p9I6V6rrkuZBsUQdZZJT4dDK
ErJmHwg1G6fTpJTK4SifqBghFF4XmoxWjaTRhLBiqfS+S3LD5nang/7g7FDLHZQG30lBurLaEtvs
U0WrX8y6AV2KVKjTgpIgeuwagJ85pctTqXgLbtn8NYZIEyLDKD1l36CoC4ALvoZAMR7k4DUiBFph
MKMsGbwFm/RBJMFrskqYah74dNXKnI8yYJZMVknUGuwM03BBM8KBt1NpEL/tsxYBEOsS3r3PKYKX
M5pu9vuq9z4RUejhYXe6Bdy8yu+NK+OwP3OJI9shr+BsVk/PX65TQc8+I5wS43adkqpPS3y/VJZg
tRosZu8kZOtxxho/G5S6nJmoEtJ4LfDtKEwpNH2DrW1W/J8yU1dMBCJOf6zOKCrunXz5k3NCufFr
ez4LZ9w6TvOu1iW6fcPGIxe6DAM+kBOL5qpwoxVmXl1i9QHFLCMHkTXB0x8+rBXhnHG/91ADJP3r
cmhf5MTPyj1Sd7bK3uUU1XX6NVzNFOTUOaMWLSq3JEwsfqKZFj/Ezz8LA8sfVamSe8t9OKAJZvfS
8A0RlChsqZKOAImmXoL7YkqxGC7J6Q+NsIhFpm1poNWkLb4z3YMwOzBF2rzOzE2gSkG3w51x8d77
a5vns+wMxiV2qDBuCvkCVnRoAorOiXxRBTS+2GJ9nqhl/JkCUEKFVXCLG0Pj6b3dLkMZDakvbg8t
HpdO8ypzsD8JkWeMgZqB0iPgbcrgx8He5K6NK4F5KhcpW7jTI/0Z+1PxqcTXb+N7NU3I9lQL1eeo
pAyjqrqX+kfIiraX18auLP35qTn8Z2PreTdYQ/n9+f3QYg/A4YXvXgRRUEAW/G7TMLLzCxnzlt1M
5fnZK0UTtD3I9Na1PuicfWRa0YiqELyQd40m/BeYgRAc3lHnYY200HD7Ob18CGpwr5Ht6MhV6xUZ
G2VU8gzwsVJ4tn9lMDycTJjKUGFywYtKdW3uU3Zxal1q1ZrloVHAENtZjSPBAnJt1+zBJ5ZoaW32
tDDtMy1O538wxM6i8DDRFVfk6ZY9wMVzCh3hO+czG+79yNlxPAbJY9FNFuGC4bShtcKdvZtd/bPX
xo++eNC14ZEhTMxV/3vpPxaLis95d3tXGR5816FjyBVbU4fOiBy87dwesWMEo8njeC6mfweYK4hw
YtVpTC2naggxp9EKr9arAU4TJMY3qqQ8X3Lvnxg9ZPuaS4DK3yaOBruZMC1EBG+EKBIkNa0HH4nA
2vWwhH+v1M6ih1RlXndFqiQi4jdg3B0XAxKV2PFJ1F/OlZUXpIWqc025UbMsm2pYw/9dYWAtgoqg
oisxonYZfMUzAkKeKokHy64zVKEgbFmFuTbt/AeSUbPq1UGtBB7PV2/9Y+N3B+loocP8OdKtd3Hw
Tq/Lzj9F/yqz+lZefwXg6Iqwn8cVjSYsLRsIhCiowhhLaJ/Dh9HLMqKwM+q/JR4oBqgFGVpNA/O0
vAxai01erk9B32aWU40fSNtoOSqlOmmLaIU7GcY/F82I9zhOZBrmrPqmSfxJR7lGAuC3FnHGy2ZC
IZNjFKpbsCSlofopO8lqhpyxaR2zwCHOsZ6L/pdimojU537tRDZoc4zMnr1+ChflETwOYkjKPGB6
6T99+mok46+J0d6oeCqaJvYGIgJu5BqMfsmt6NK8SGV7OAqdODanqjqTECDdXWygnU2k2rwByO2N
Pqlf7t1rfMnEpC7P0VseyQoHveXsTzQaQ02l25m1ZMQGgRk99ksCXFsn9wd9hP/nzFu69ESvVRkq
8UD0Dwqqoy4UmWjOaSXRZGR4IJ6ASYY9TMGGPmYuYlXG5yAWk9fAB86A78x4ABWHPc+JoiBtmfxD
rPcaUTYsFlXMR6ADkEMUa0wc9TnrU2UEkGlBJFMpMlnH2bhclNeLBzDk8Cpmj4G8JDAXK8FmHuYW
HZdEZqZpe9tgF4YvpQOW3aUtflF8yeJxFaaq+IdJ2UBtnBsl8ItphOMLqeBKcP4HlU3rkXz3zJ2T
LTArnZZiPdy1TdYyoxFVZJw3Nv7KC8Onp8fUYLZ3izUzi8xIcrRrbfIxDU6DkasczzuppZPdcC8r
EUAy31ZS7fdu+OJ1ApfdVL96BiWLu/Ps/Cd6QxgafwTqyurnlCyYqlMpvCS+w6Pd7G1D6xVz4ckL
LUjom3/kUuZTCkISnA0oJ7puibfZ7+mhFWEC2qtU5ZQGijcOBQFD0Annm43IRfH689o6aitUioxo
zBX6b+maAYKNNm474vgKZqcwObMNkzbsig6awr9XiRS7bUdwgivmMhifMrxoWbJ7ABfddxZTjXo7
Cx9SSwGojtEiDB619IliMHNSEuTP/1RxmggLMazuxPOiGzhGKBbYWgMRfIhmsF6EdlZU/dqeSetw
eMsye4fnJzuhBNnMtvG1TeJ1LVphhjbuGYufnXATcgrAOFLBFKdI//qdIriCv7sJ1szjiTuyhctd
BGxYB/1BOE3qUB/UndCT6WY146R+gdwLwhcbLuoISB9ytdStkuZ/yU3XaOdnY2u5nlSWrLVG/eoG
6rNBZCiPT4n/eSsK8UaG4ElbZlayBxIH3zPZ1a/9vWWOEERETgaDEVYp2xMP4eWG+HZSJqElOc0k
Wm97GHFGbZxKdsNnVdp1M2mPklYz0ExTanAl9cJxy0kLcQ2W0ZJZ25vD4xSM9zMpotugAyDi+/Mm
Hs8NHdb23teNXsc00RO9oLRGfSAkY7xG/J+Bl5z4cvQEUc9UcpTDPSLEHZIMxy4wbrfvu7UMv2Qu
UWLH4dx94xDaNgIku4v9wfu6ftk9NKyta22SCvj8msqMK6EEdj7Zd4EVjd8rI2C7vmJNGNmWklia
HJ+n9LEU/EOzqPqRYLusEbaMdzttQfCPnIQjFPhugXM0w7CXT3jO9u4SZ2D4j+O+NPi5gs6Scjfh
Zz6965SU3CdQ6GvYYfiEMpIFOiLd4QB//26GdcOT1KqoVDEA+TzhVN0nh7+qSfOJPjdWBy2rjbku
Yi+NePLyhLAUzauJt9/Gn8TVsP189wnaCbAVWqY+pr81YRJYwMp6psxJh9ya4lMZnytLPVWlKGXk
tStJCR4XNjh2U9+7pXRiSWH8BcxOx6NHzcj7KcGZOKFhPUpnVFFsVmPW2ohrx1jJXUenI/km/ZoG
FUhYZAr0jbZ8Fw8JlIwQx0KWJvkzv3m1vY+BRV/hVNcnD6pVgtdIyMru5vgGqm/eXwiCCw+eIvEi
RSQNvA3AJZPUQJiDBSSq5zsBTqv3+wrR/H22Vh1Qm5fbT5FqBbR2ZewEy5nX+QWJHCowencekRZ2
Y2D7KkPKS94arQ3v5bCYuUnzGci5vggoEz4OOsVVSs1T+AbRIzKKrO3BD1tc5/IOUuXikE3hLVh9
RvANnXgI6sdrsIoqMnJBMOWlkXiNrLq4Ip1+rFRjHtOG4zVGpyhYH/vqrlLDcZvosqe3GeUJt8eC
Zp4gJBV4FobKCKqttHr3hacHEA9YU/no6eePU23RgT8hfxyaRghLrc3W/auGYRKQeXBkKMd4T7Zn
ywxzAKqH16xny5TSyolR0I/eg5n9APUurZXYimBYdptPLzF+QzenRIC0XeLlkLhZBTbRo8IrQMiC
oinBABAD9uUIoasi6HEpNK/jNme/e6NPGdi6JvHg+oKKOeWaeU8AktOLeG3gmcnvm37YWk6HWFV1
M5g3e9DbpdHM4jpXUTL3UbYzqfnbYWDG0EP+NNMKb1uydZDEmzG9CnAj0xSRx+1RoLxcIzElaJDi
js/9Z/DdoNkp+aGr2o7C7tjtDVMuFus81PdKI/Eog3NY/xpz6nK4OAhJKA5f9bWJfhNIyDfnTflc
IgESqryl5sMf9a3ONjN0pFQEnRla1+uvH2SmNQHM+xhgaQVerUCjkQDedbKE7kosBcq2S2+CSQ10
iLWkh2gu9R9ire/3FTnfDCwlP5XeL3BCuaA5BxV2RexE1yDH1/7Geez5H2E/2IF7MajFWHcK19KA
HYb79fKHYt/Z5wnSGFf2ffVGewp3rCEbC9/80Ch4uK5CIWY46Gm25aXL5hlNtSneV/nCKmPJYVEE
ESrtIJW8T7f5tziucasScQu4WDHlTY7XTJYHngGlr8wqz0dyHKa6KP6v/uB+PYbGCTP/kMF/Tt2O
9wn7LIK8SxpvQ+tTw1IA+98XFo1eU5gmkjQfNoUaPSBKHnCas6V1285zYFzHDRuoOecFVCL/aVOK
q82fTPg3OLpm2Zyg0udWP/neKUNwxot6iBLAW2QCv4yDKuWNHsDFikS+lu5Wujg30Bh+kwJNcyfh
RKkxpLzG/Pf6Ac3lj6BZKdDJfi1G4A7cdSaAVH61JNdjDO0MKd1M2ySwu/Zv8y4aXYbjBj1kmea+
HGFub84HxOThfIBRoDu7uiTKZI93YLjFoGztF18efT4d12oUvKvjq5cZFGdH1GsiBA/5aX3cxXDX
q2gjkGQXOinqDG+cJGmU+Lp8CeVcG2bdCcGzRLdK6VUEzvlUjYROFRgQsIUjZo47vD6i6NTAjuJ6
vQQPtMl/zqZX1Et7+L03wX+cDnWClL6OViqdQTpFSQbOgNqyMah89lYxSrldxjHZpf/M3mFOYlzl
c5Q2M3SQZpTk0mwYpkAIbYx+4TKBeXLD62zPPNOkPSLF8QsBy7wxpf/2tP5a+BI8XkM1zmMOtUmh
7yp/rZ2fjztZsbCrW9Ddw8SGwVP6ozeXlGemA24t5onorc25g0X0FRi06uF/Qbrjt9zLmQ7wMqne
XxaNt6TZvvlpzAA4CRZ0EdyjoDqfSaJV89Ftk0V9QthqQ6JAKGeEzwYxpkpZI6L5QLoX3yBd6PVA
QNjvCD7EeZrRSgtOi716d97a+Xc8kub0BynC/dGz7Za7ngqlDtyF7QS4aYC1yiLmojTNBdT8pu9t
5wb14a63jE0cEQaIxOHRC2iK702pjt8gFNaHo5yeVIjF10NFlz7U9Owt6mP1W98LQM9JHHSlMnLU
mU3g9gZCX3O/Xb726nXSusAb2mRf4rIwx7j7JtA+6Pd3dNdTUwOgGVOE9f2KPmCVJvylfyE/bClf
DDa+ubS3XwipXnW0WbKeRajoB1Ce2z78PgH8W+8VLYFZS/6JqEO2DAvPVYHsUm7Zq3HEkVJ0pkkY
qvRRGhQUQqw/Ir7SOpLJ/biTZsWAeI2PTI8XaKWUZI9L7TiJZ5QMYlGukb+WFTgCn+AwgyWYKKXz
TklTuoYlX+jIkvyqRKoOCCMfuvYqc+NxUmIqcTUQjcpFsNzfPNUVS7CoxDo9hmbLbCzk8qVVIANx
uD8kND0Rary7wXVeIPd6KxKoGpRk5LGjTyb1XhDZGw6hZ0khRA5H28bjw3NO+2f6bzjzgHXhNpns
jj27dH/TSKFyJxw05JOdr/JMZrt0iSp0d8asF4kITGKFCEYBwCamb0gFL+39ylnBV20lx7d9YISe
vmJ/g578pmtZ6zfBjOoKsvKIFEL0dMJ5c9aAwlHazJAj8IrHNp/w8wZUAZ9KXAfv50Ug8w8ZvLxb
SlLhSZKqGuMggDVLKDzTQMop/PqK3cEazk7H+hKcQ5POjElGhJhk5Pr9IoEVZE5x71/zzIZkFli0
FcntpLMG1zhu+VzrgErg8ANJnlrEmpwKO96uPdYsu6L27I0dIlLFf6Ex3ip9UHnAy3KMGN6iq7Bo
3NYN+meCTK5EqL/EGv6pQezqoLdCKQBWWEUxhiVuC1FneRtEsn0vlxORPInV/CjnWTfmMZ4rlL61
q6df94B1NYNW0pNlSMZDjO1I9q5jUcX8N4ln0/B+zWuETzoASLuBHCMlkmCt1zwMYiMC1YXynk09
+vK2mq8mRUvCRiRyoBAQoc8j70zt6Uc6H3WMHSsAS7lnNKC7ewyAtXYFXIkEmho7oF/jfkkGGpHz
E1ysw1/jeNzoPK1/7ZUjSMt9Fk10qQGj5BZbLxFQekniCwAh0nB9w5mmnJonDZn2mPeqSB4VrH5P
4y+Fvzp5IQnr299MyuJI99MEZzyBfa6xQ8h2xsfxMFGGDlVgNCZtZiJWj3435O3dXnqemWiv90HZ
WUFZnb3hiC6//gb9QBeZYQhXm1JkpprfKt8ibkz4/0TIzn3aUnF+cwGddQr4JNC8ul00qhKHZg7f
uFgoaBD0cdkzw9TXscLt6SoEWxReOrqInimzUlk1w2wRUfsXc6N8XpBpMOuFD6hsJa7e3yyV2X0H
8LhNRP6RHjVMWmHK6o24pdiQy8v4DHlJfcwTTiLB2sHKsbnRNkBFVrmeeWkramr0TO/WzFzQgZ8x
fMljsAab1OJhtGMGXxn6T1mGuzPEugZnqRFimN4BH0nkzDX45OqeKQbu10LBrrepqX63Kr95aMdf
7xS1dOukdcdc330MwnDy8qiqMc6Tx/9tQP1VeGepO8dncDH6o1gczKZ+QeBB0x01UZOM54q0ZlM+
dpuIlFPimp5u3NQMzUCG56KwDaLsluxMQUG9arhRizBL6IE+8GLThQBs04BbIBDQpMyEg/rLp/r+
LYNT3mfLBTRpN1OxYsXph94hr3Q44t/88ZsTA+gtEtgdrcglDh9RaY8H1vED/0jO5jJ409ntz0sf
u0vGiJ0LZ08etWSQHBR3rsMXmxf2riLcKglfUNCcp/8Kpr93VoI3i8MTw7xBt6iA4+AhFTz/WUQm
WY1+MCMRJjPN6rU7Av0kuXMPmSv2QSdo9UFPm5a0IIFTWn7TT+IfMNpNFtE7XcUGivbP2oM+2mQa
950kpcTNIqFfK3/FAO5NyouNixUj8CRXP/726DA87ezu2L9HfSmrosXMhEtgDGTp3LystlSox79i
K3pnMbF7tU6ozn8MLzeYqN12MjstMxsmWmQ+T8CDPJfdqYfw6IMxI2P9gLDhPs4TR9AfhbsgLaix
p3117C3B7DXMr0rMchoUQWHoSwy5dw19Zw0lwAlvMquauFdx78Ap7+3cKOzEoeOLh5Pdwex/Bj9r
1b7CWec3A08ICN+OcolZpXtQzEGJeZej73R9wWN6Wjs11tvBXRiW9aUdqYaZpMJby0GMlL+Nzbzq
KN1icpkZPmcwb046ZUQSgyGQ0JDlrxyiLx/63668Itu5DYehn0fBZt6pQrqVO+ESqhEE5M6Xerkc
JFwDg9n6LiU9jxWjANOmVhzdDjgawml18W5P6+jk1NWA2yehiNq8ioRLa+eaiJCXXQPXkWkg97DH
Y0wdV8e8Pp2mWsYODb/8/+xzSdXYQNuVJD3VWJ+3QCdRWlzZZz8p1ciT3SzXAXYxh9tdGYNwZHEJ
/I4opP5o/D0XfL/jS3BFJf05hLtjIu6erFbazkHKWjsvHcVRLcWY0MVl84/Xt29Y3GqUoFPcKPiy
IbhV5caLoECjaiejjyVYtuX2SzPmygyQGgrWxYH9e0vtx62DPE0V58o5xzdm9qZ/cZ5Rj5p9l2zw
/l4Gyt70chA8KogaHW1iqaucuHCKI5l/AazNEs0Mbq7gnpvDnLz7Da5ywb1k6l8N3E/12bmRAXJD
FDCuhZWhDPg+w06/xRnKaHC6BE9FH8cVFZ3h3C6oK0VU8TZwlTwIJqkAUdrCKaLbQYsf7mgjjYkj
6MiW06Jth/BZlwTyBFcBI7wmDTlkyK1Ue0gK5P2aR+W8AmWb6XHcFTvwMAYieng7jUE8N8h/u2LH
6UTZdKaURsFv8EIkPdO6m/fUWnR0PT8u5BsjE/nDI73Eni/sr500XGo7+w2Vg9SRxXKbZW6pJyuC
tCNCJ5BihgFroTgLqDfhyi04VIIPIsY/O82HP6cFm0oJvSV8hx1br4vZTiYGX+lCz9KkEwDJkzaA
+M1P1MTghcionSr/JN7AZ0LXyxhAZU8mWgDJc+KTukunEOasX0l3ZA9bwubD0qf/0tgW5RBKFBlk
DZ+b3Shz1Pk7XIlMclGhqovXqSpgGGayuKR2aUuBJsEkkkyyD2IODnoRKR7RLUIIUng6/7XvDqYB
SfyrWPP3YfcrhErjAKpl1++W+nU2JL3u5UftqikUJma+2q/7JIlfC2axR7rq18vQrGcNGg4MYM1R
+QnFfB7jcttCG9nZ1QWfXqnXN3EHg44z/MQB3fQpqT4j8Lt3bKQ6qNc4VwfgHTsUK6JVfbz7+/os
uMJb2BRmYjujt045jvnSkGPtqVUGG8eyDrBzrPPemadMp5msYo8DBN2dEd40lRk8mCt0HVQrHKNt
fLuC4YILAibi5LIf+oOuZD+It4Rjzl9HNlV1zAcVMFWOyZozvs29Ubdnv1pIfxCniONHoasRhQGm
xqy/d3hhD1TuLt0uTafYGvRrFEu8L9+vytALnMKRLeqrKcRJKKFvsoUSr+wDpEUAgL/CbZ9o9x/4
vm0zGCJPdYFRDXO7Tsb8JeoymwLqbm6EdKB5BVfLQv4cX6HE46ReuDnEjKxKVvHHR1bVLvsTT5VG
1kFC/hh/Squ3U23KiRoqv2D8nGG8AnvH51oA8CDhc4gG4tTL7zt7NEcCSd5wiGX0fJTatbsrtlLG
++LrVDhmjpyoCHZ4+aSb6i3ypXC5J+CYRIaO5iXCwMj/40pt2Wb3oXlv9mnT41Ve7jYt+mCO8WIE
+dOntJJmRyYqFHurKZHIdz2FlY3Hu5I6mPwNiUtz7wD5i8irjlvmiXB7LgLc9/Ur5GeMYjyYF6by
+J1EzAP8rtknQ9C0UJejDD9yWGhHiZIgTAJEuRP/yI+/nlbA7sso7dr3vCI6phqb8lyTlI704Rn/
pkqzf+Ahy/lqfoJmkzFmVYSbW4qKztmhpiUTChtJhefyQO0cBVrIBWHG0FYX+AmfVY+ZQHYSka89
fr0TohprZPnSYtajZZmUJZHj9Tn+MYSXrYSS+3+OLO6JHdOSrx98Gfmf29B5VqbhbA2/kqFo8YSj
WQU+AzE/JGy6nN2V9VmcqVKhFyvdeiTzLmJ16N+8Dt6vwAkKoX11uVfF4uoUCwyTFQll2SLxsSEW
Gjh2wY3wOxjbOBiVNGwBcapVjO7rblZl41fnUmIMd8hRccK1hJyj3HKfThbDw7aCJQYyjcr/VK7+
QzEdCJgXpJQ+apfXzC6Xu4b75WnfJZxP4z3xmcQyHKDhhLGzGbIzlu71Kee2KUlQgD5j0xr48974
aueVS0Z1/BAXxAoHz5PZSZqQc5zDyt8haPf5rWP7E9qeRw6L6vHkDQIVXqNS28CVClS/nucHqE5w
pRt8XCu5X2XV3fXwsUPkU6FFp+42z1RFNwi9snP1Uu4daEFiae4Z13a7uV4Sj3LEI/D895DzzISJ
37BaELBeI+LSR06lzF5GX/SbHllEcZ2C91Y1ZziOPG77M+hx9CaaJj93M7l8lN8fvNpVy3Pp7NMc
s5WNdDagEZwRAfKQRdOmPqAhr5n19chKiHlLc4NaxKflB11pqFwvbVZ2bTBJ4tgzaysXisWI6qHe
vf0iSkxyo+KAKDXmlRMODUdNFhbqXtMCidaML8qyVZKE3/aeEQKuz8oWPe87TUVocFw5/J0qpWpD
C6GmP6B56hYuLTZ09TjnuxCgfR+OBezaQKb2/lb0hsPLly6vaba5avduJOFLjJuui9/D+j0Jmh9j
2VrjH8Rp22LrcTFNZmmOv8Fohcq+FT0QnQd4LtckQUoepjqirtmLgv3gNpegiI8eayW9oHdWCU/q
KUVgXG3APU3lj2oPPX4nRr6rXEkxoZ6SGiWkbFvMPAfv3p/+I9HBM0nzlGnKsmDyRV1MDmTeToJ4
H6nlRyz0pejc4WN0r4ISeTqFaDbX2wRURoi8a/E5Cq3WTZrMnHlSUUaV5yD99OVwHlDIBX05yHSU
BEN/zxa1xrweC5IHljWXT5a/z7t0AM6sr5IYH/W3crtLjQuO9ZkaDuz50vAzttgVBO2chNqc2zJA
qt/+p++pbsKXq0ZgR+JoKB4RESnBXmePsPMRqtsw+QzKbCeTR34kGmoxaFymoWLqT5hQKeBd/lcb
9i4OpdPLDLYRDLX63YKVSmban7jsCdmQunei3itQPziHVdcJu6uqHxVYRrCU3gsz8y27bBoYwjqk
2AwpN0ltg04gRQ0F3q72JtfFF1a4DP8vT5set28zYvwyG3leynlwQ1d/Xzn+Lz5APCmAnqw2QwMy
4k9ItIFaAjCN1cminr373mfOoIT5lnEUi6JWPuJ18dICrctdenfR6EfuhYR2rJwvt7qM+8lcRP4r
247g+S4vCDCW1WxymAAQ76TSpkmO3q56WJa10GZJEIeZpdlo3slNf8IgUE3rXgmPZxlLWVzTKc2q
sF9np5U95EURhBykAPFlOeOJn9ZsgKx1cqrFNK0i7p4DC7jH/33JRtP8dlYX0Jcdg55b1u7vxTsM
0DGrQ8QU/Fj584xu6pYHniNjNms0tvNBXRxEc1LcZpghf5Xy44GaFF5UM+w2ZtGI810JR2fr1+Mj
SXDUWDLLnU81685D5aVdqOISbncF6PzCHWz0hVPDlDCIS7cQzQPMdb5pd2enKZCUsXlUBAYaqLrb
CXBLQv0yl/qdYb5nsk5W3GwgGAGgenvtV9ahusHENsHm8ziv7pNo3ur82/TVDCyQKPm/n3MZz+eP
Qr25dTZuXLCIIew07YxV+XPjfjEC6tePKmf7Pg7/yd9afqSVmvXbgUn/Deg/OpH7TlJC+qmeTGwT
QSBuDwxUiX5z7D6/1bKDr47s/Dz/UHij25aO0f0iIKtqJkAdB7PIcXyCmn0rcAYJKbkR6m5P8sD1
7vxZcWMDO2YKmsAWxS7j9s82Bp3dTG3xAgKEictA4T8mTXZW9yqyBEUXMaZ2Y92+ihutX+zWiPyA
yJRqEXxIqj1a3yejbzpLHf2MgrywkeNp7sYPWWc737EN9ujvJ8DhDZ52Auc+Iwd+ReWs/p3XJ+6C
7v1yYq5JbX6aBEQxoSdaYdm3AlhDwXIN2YbQUe20DL8F8HGP4310I5Cj/t63JqIYI6rZUgt83Cw0
ZXhBsPeZHNav6l3LBhC1+VViV3ZvJhXUtd2Z1U+nWnPUIHBKM4fbYMRFjMcss5Dyo4qyU4mPy1I6
0JARWTiQWVLct3L3V5QXbxQc+dkfntllwOcaGgL+8INiQhDiLW+fAIJUJaLt+zfgEPoIakP/OfVY
21V71WvGV8ahd9XICjWG+mURwgKVy+LkMQmx/+6UK8cFhoFVmA6NN6rJ1AU//9fl9bGI7j0d5jvt
Iw6VdJqhsmCTqNs3qG+yurJZbI6/wh3hiTwO1e/KgzaYJ7Jli1rUA+wzymWoa08GbF04tcDlvmwD
K8aFTjUBUREGczx/Qa0yALPXZHivmofSYVsm7iaH40Jfjqt+kteFnQekGz5nHtavoynrFwqI02D9
QA4+zzJvLbA3enBSMeJx1/BD2dxYpliT3Wph8KlPkOrG5S7fFw0WF262N/hgv+WCkdemzX4PeSBc
VU2SD1oMQSh2G95iPQCGy1zDkakEFzESha0WhADo17zWm+iBRhjvrlOFdItFgwML1lhMGGmA/ANp
sQPeqrC6PBXxT1ew0+R2VBiYT/n5nJwD6Pv61g0x3WqM1zTjHPGgssab1oanCvPRu5BsaGi+iNp0
9nrtyN5f9RjGG6rMqUGOnVLIFjaVif6Isd/MMXavYJDgM0QRmPtJl3f/cSkq9G8MfTlZlYsG5K5/
Rp9k0Nlg4qFGsTNgLn4ojW7hz2UzxKfwh90CtFya+wJ1CA6y2HijdB439AQf/3sJ2PkitGCw+EB7
RdLv03cMmqiJcxuXv0xGCICvXlLWUk8SnlAssIXnknKYG9XdunO6bmhU5QRPPjUVmSojOrcYWZQQ
3WdyZTw+0UJr9NcOgUhd4BamzhjzawzhwGaagU7EWQ4fWWOhW/hKC8/QEmKXmumoKbgg1d8yrorK
iPgHLo6TkSeY1rQKgRVsDagJ0jomoole8H8BJD35ZbtP3YlCt0uI43AxxIVJoDm9KfTVo+rJpcTi
0C3+JyKn06kJFdu/RwMWAjjMN6jcYQ4JA5jmXftaCMujkiomQgIsiZwVioU3hnitUeEWZiGS3DPb
UuOX+M8gx+W/25VjhfhmHPfupdHA1YUu4Qp6wjWw9DZkp/CIX8NQ+sowjVtcMm2H2V+5CsT0xth7
90Yrkcggx8q76RWtOQKid2PTzZtvLvKkqLXrX8Fbsmm7HXTmf+SEO29fx2iCOESBJZNJKUgaCdPu
sWYA+FpB/tN3Bca2J7uc8KCvixTfngZjtXpa9IA9SQal2LV+zNQXdpFUFlmQD2dQVxzslzEVyb3U
GfFenunZOkD4E5NFGA55iSl996HUKrjmdWZQSvHyWNE3TJkA3+1D4L29GYQjcWBuW1D69Jst6iEf
m+tHkcI/FtJ3s+zBY5v+0SbdRExzD+H4DrAf5AjHaYxBLUGhC/kS4CqAiVtPxEMdnvtQ/PAEluu7
3dVvIDzScfmpU3GNLQgOm3O9DO1FAcbQruxWvu0nEa9bMIvox0SEZ8vPNUehn3oQdlgYMJNhzN3t
9soh5GhXonfcF9FyKLqbItsu246n/WQMGyzp//gYw5c11uI7pAz9Tu0GPhMj3zEy4md6elNCdNwR
Xmm7665h9RO85Vlme0w7AhCmfhgYvrvBBuzA3l2AH0q1vrJ7rs+gMMuYCJuKZFnCMhaMYHCNWK8N
QU5V78eDojWbtOEwPIq1Sn21XeaXzPZg5ckj9pXSiKwiwE/R7T1ziIfOD6p+KPFgyniVK2URYaNg
ko/iuDr6/Ko9FQTqpFHmLsS5AFepZVQxamyww2ixGWaebUIS5RqCS+VlqhZLxUND1uGXJucn0/G5
fbXhtN/PTuZ/yWQuB4pDP7XTy6raG74Ab30t+0dy4kDQW0ppBzecZvqq8sfuHuHW3PFsEz/O2Me9
6zTMFjAYcqmfZ55K05wa98tPoCm+MDHuUw6Q36FKVjI0cypAkUqMHf0ZxP0uYtMTh9yFgy9iaaRG
aYLhMVRIId1p8ldMdu0AkroyIDFFwn+XHSEQWSdxs1hlf528qYh6Pv9dHoePtlbLDgG90Rsggin8
5SOl03Yo4dMYjBlCbodsynmRF2Xf8489Hv8mOq4l3dTnw8nyt14KbGgkm0cUhgE340fASclJvQtV
eEm1X2OHS7bnXkeXp1/MgxtCp33ViSLvODKVXy9T+Rr+VFrGzrfXx+foxWiVx5v9RItzvkZ5uw+D
xvhhPW1AHYOOg7mHAODJqUTzq5MvxzonznqrH93bZcNXdL9ZcXlHuutYHFabim0Gh9RZtDrfQAia
Ot/BS7EC+H7dw0Sp8r8+nP2E2B9vCHE0dwdbR5hvB96V9u0vwUavueCrhL9kzKxg+p7yVZg32gPe
PMapsp0QElIy4y80XPLtgPLD7hnd4ys9WWQUblDbRHdJB8czSMszr7wCHHIrcMpSKWdl8iy7xf+k
usP363oeWFhrnj3LAfMQTeNKzDclQF4JUhop4Mi4ohTtKu7VWYW48KgR8Np3slsQCBGL75JYLI8r
Sm2YrBRYH7L7oFcn46i35xGEKv7rBML3L5DzEB6myzUkeAtCcOYOan9IgpRNVkDvwmM9SeLVuaIS
Llwl//WpRbr4kGUKSeuRDIj4F7XseOPTDUng1pAlHfQw5mbQeLUmjDW2KzfaYmtqx9CWMSDtKRI9
kKvOpgpeCJwbuWO6SMLFn+dIjJfHw6BZyAHuzlGrdyRqJlrdMGeVi6MJ4/3nv/y7cl+dXeqojixM
p1WTBfbNHSu+24qkYEdUJXBhGjIkcBM3gBmmtN7/qdxyWS2QOLt+6qGfccvPbHXFoBuas2cmibBH
Ig2MMBswwjvZigfOHZBIH8Zs1Qop4NlMGAcel7z0rnS0EvmtvZYO4ND0aKbJirIjktu2vHfftU3e
hk0lWqIYt5HdPG7TZBpu0ONFHIHjJI4Bz49t9Deg7Pr55dnTFae92bRd7Wf68Y+RdK1RvckZKCG6
023PVOzHtjA4Pep9Xv+FluwKIPNwX6AJx82puzxn/1HPf9KOQ/lRPF/snabX4IXD9eG8wMHM3sJM
QR6aEtth0iwb8AVjxWeXJhgC5buduMq4Vi3y2whtLPMfus4OyENMz/EfgLHRm1FuJHdIS48boltd
aqd4bSjnU86D3+Id+4L8sjNuPL8C6k46hr4JKs1mj2fuggCbcVd/LSG8vDuz9J26Etea9Mw205v/
Q+fbxQueI+bJlK7oGLYvtZh4TqlLB1YNrNN6mWdi4NBfX3E+9QH0neGzoOz5HJ8g6fR3Owp3xzsX
NvmgxiUnzXnuvmfcWH1PBsa8m0okbWxUprGXERpWMz2dpzlKJ9nhCBmLC3Oe/RmgYQ8MwzzggXys
/eYcOa+WtweUzhPg0koSKgFICPR355gzAqzYCgqXiccUTJXJ15rOuTmdRFSuZXvVT7zsbDpK02sD
BbhMnkqZV/gCqXc1RLns7PYE+21I8q4siq051KN7pyHW8DkH/RMIeX/jE4HABjpP7+6h7PjMPLvq
rU5zJ+zQ23knlBHx/m2SLjI+9gbhQ4/mLFfNlCNoYRHk+A59pEZvG5FgEb3mFhr7yMBQrJlUdzHe
0f9K+RleivTLgPoQWaxAQlFLFlH/i7wu+kQ0JeeViBdsdgDoaThQj0q4v7iodukoKqVtosrC/CVo
XZ92fgpWwRh8Jhb8iXNXFS2hdSDi1rb8L+PF7a2Yt31uoNXgfM73J2TKUDaonhWq+ggNGnfh+Qu9
DAShSVY7edeFBkOuXhAmTxvQv+VIQ4VKPNT+CpxP57YtW2yMFzZgwJVMg8bXCPrKSM3RIQTBreRZ
ULg8xMHi/tL6qw4TBBQEpk/Xm9y1XLA7A35pyWT/3MfGtgvz05G+7pDjJi1tHZ3MMACXL2sGF554
cHI/xkhfHgvsrkx378tuhWO6969zishR9iaj/9D6GzjwGgWx5OuKkAGV3SWeV0DvH0jHubnLt3P4
6qOzfKAF53jehnp/fwHNK4ngjY1JY8jSMFpvegUCsZyZT4l4gwzM/gv2LYDFOkgClQzfhT7fLp2W
wTrkK8LzJGQR4ciQ0Liq3QvRtp5LWBV0vVGTvWkg5N4liCgvvKvpwczF50j9YvgMgrYVhfGl1iFs
xk2TPf3TM/SpWUwkzRz6mjgBVvaCXpfIdJdIL6oe3fRRa5/j2YoUVEuagbUMUy9rP8aoHlPIA5/6
S1tKu56l1LNxohjU8CgyURIr/AiMJtpKKYEYoFDd+p3qQ3VUDtocX9RxK2MOJqZdOQDVSNai6tfM
fmK8mMYjix91g0UQCnWY/79wTbSNaSCITV8MbtwevLFO+TjXWkjwDzRU/6ciDB8WlSZT5ogftzaq
iBgCEK3kgoPCncZWzbiLeT3Hurs69EuGAOrKhlMvbYtDod+VTkaEk4sssw7mhdg7XOp0rOFm2lNE
dH2MvD3+GlqXkg4lag2+pfr+nUUK9N+0WzhJKStlC4Uyqt3mxes2Ibi3kDO7QL63Ru7BpoObIetu
3hqYAHEgkb1+6RUmsFsgymHvRUsit1K7zHm5ifwGZ5dxdF9A/JxqNBPRUSQjEg2iiFUmMk2VJKuF
ap+Cw3cHkDPQL3aW+SYgod24TojktXe2gGEWSG/mOX+PHk4dgQilStzlngsPPRswXxBSkty6QJrn
Cqut217xCKRf4DkGiegoTZnLNkiKKm6AxOUal1vtakDAitMfQ9/SGow85iIMPBJeNXJgkrjklOXa
Nyp/STIGcOrV4r1AT+9jBP/PMfaxZg0pY/B4DhWJEwiSMIhWjaMvFRcMB67iiBFv42/n5Rk1TfoH
s+RXf14KVnJsfQeGbN4crctt+Rd3escjbqJGHgjh0PtY5rAM8EB4HI4CTYU1WTktGh6hSRGJwE78
fCBttvpNzZFqQBR6NqZQCdVlYWtrWTtLyJYok0Fchy9xK6an6ZPMHPGfqUxslvmY3vAUcfX2C/qk
lIpJorhRI/UvPfcAcHtciHdqzod47D/Cm9nvSQH0ALl3r0u4F8BuT6jc83F1Z4gEOqQdvZl9ePFz
VZWmFJVDRUhKumwks8+j2p4/GPuOU+GT67vmTei5fGR/MeV6erFhUz3h3BDSmBT8oPd9+FNunFYd
2o6+1ea5w2+eakhqVIz1SjmAUo1U2lf6JweQQeo0K09skgsBsEBc8jcRMvXTdCGWJhzRn2uGBCPs
5rjFb/soG69PanvRoozbpMrFgJbApao2UFwg+vRru/nLlly2092T4s+ANugdBAScriIloT3b1/5m
L3oClbqZtZZpk8JUnPMyWuU3CbnjDGQ/zOWQed0848zs+1d8UEYIMHLi/3TAdriRqBI5Zq4UF6pP
VDp7qmJHopFUX4xzdULVjV+A9+ClyUES3ate1KUYe5nYHG06dN2avFuJ2sUPk84cWRfjc4/XZcB+
YWD6tjHKTBKyFA5I61aqwnYksPzlBqew/PC/5XW1PULw2e81lOgOV6181XTE+rCqSQFlo9w39ALM
0HndXtYYz6bdmbaIrVt4+3Af7LRYM8ouwVY7Z57RAeH1aZsnIdhsJ75EysqCYoVRN1PG+mdNFs7O
IBe6BTPaHIGo4jSp5S48g63M1Oi8DaMsxpKPU6kn8oGB/WlGbvS8z6fTh+4yBW9qTTFgrM7f/+Tt
ZJDfG6BAhEiZqw/tvOxNv22y7mCwFLoYC0W/NAsDnsAaDQMg75JXdfkzStgutDxtNFq6btJoac82
6cvCsdI4OXfcuSN0c1XcKywTp/kbVqMUxQo16/vgtGqV96lO8WTnqza09OWi/vRoXVr4uPtnPK0r
5/9qLt7dRHAM7CGO4odpGzlAl+WUvHdUMGd/TWmE5FUnzhujbJudiFGQduHpOiU8SB+pQkWKjJlg
8dFpdwg+RW3qOZsOQaTpOLctDSgDJcbJ2NFTbeTH+UVzZGjrjCdHGK2NnFjJX7nQ/GVc/5K6DMT9
WUBn6wnMAGrC6f7aZ+9oR04kZ18QdJSLOsiNKQ+KBMSy17EnpHtXnbrEsg0mtB0WvW+vwL6QGoH1
G7BIyqCSNJkbrV/q0mELPTAjwfFXR4DrYfpL/us2ExR+E+joA8dvI5xB+6nSg9+8J72QHpV4xcyV
p9RlwqaZlaoY6k8F4KcR7LI5ZiK61Tp7fYvC0h65+dlck0cme4tja3AQCyFGuiogKdnYx4vnYA0o
Azczucms7Mq2ZHQq4ES5pg5cE40tBy3WBo8ijpkRH9YXSSGcHIRUByCRnHZjFdmz4plTRpNVOOmW
EckChDYQXMr8+s004d/NrhgLz6cKHoDuP7DtMWNC2ZuyEHp17hCJ8SWxU3aKru96+IIy3fy5+h1H
TJvLDhsuto7+sNCL96x+Mc9e4Ru+6Qv9OSCbEZd0oQgYADPook22di25Oe7/ojrdTKYXtLlu1Tha
nwjt0Av0clrrOQNXk8tFdD90w6a2/SVfLhD5qAttJMW+bxACaml3rJvNTKY4XFNnEsbpS5nJBMyz
iOtjOlCiI4Bekonen1+VRWa2x1GDTig1bjFq/Y4rFSTGSPZgkxNAZDWg2VeNJ/cpD6Hd9v3pYj5O
yBM0JEYOte4ve3w7o2Ecu0RP37U4kTXMQGrtgHw/BmpaE4XNt4aP9u/PAA6dy9Ttw+Qx2zFK5sre
w8HkCIW8IHpVsaG2wa4a75lr9xIv4TrvJiPNDjt6HdjZm4I3rZulAqyKnpU+WWCYsW1KdO5Xw4Mf
w+XpZYRKhg1JaOrr1MdEAaJLQRR7ZedyiqaN/plqGf2ovdDcrTUfJg+TsmPEqEoVXm8HE2v3nIeJ
vwqm/gtXaHnazx8g/rmwXj/RCFGZvgCracytJ9AC3gyeZ4cLg7kY2yEO56KbONBGFTRU837JxkW0
fTArvuuYlH3UVgYZpBag4qBo4aDB0pzKSy8bDogKTT1pd/ZqQNpsMJxFaB97i4P9Yycya9GuMGr4
QgxLn+74gCFJj8OmCA8EEw3u7UsnpLTVp9xX72kcFmFR7ZQGW68k6zoXor2SBxl5uQzMdVR4tnwR
Z+oO842SNiFE+W0rsWLq/nAO7vQnU7lbv9Bdf6w731RTpYdxjI9NjKdy1QfZBEoxt7kMAZ/fJv3g
zHA52cK156+WtnP7TJTu0svUK2ERoRypbcPUDe+/SL9fO+LNza/TTcMgBlB6LOI67LEttkFcht3t
wJH8byZ0Fim19tMahJOcbvTuLD6W+FSzQO3UVmJw2xdoKuXipXm/ssoBgDSIMfF0F8pDTb0CZ1T9
4YZTjODJHDOqqN4CKDTP9eohALQWxtfeoA7hA3jsyFaEtNqQxIp11AeG/haiYgx+8XBRK+hwtAIr
LBj1Y/S/0HnEdn+VByg4FAcOyw5LX3vZ3KdzHa4MxqjHW9t0gmLRq5hSSt4Lz/rrZ8B2DGz9dyHb
sQWll5F2DPqSZLs/RBt8v4m3ekfhVY2nVxRbJcqoZtPaC25irqo/qjlXY3GDK9CeunppqFtetO6m
JYyyb15g86lvdrb9P1KYDfok7CDm7b9v/iPCTqAqU7dF4uarjP/fgEDcZLgSccRyhgMW8Zs3NESS
A40vdOfm9DFLF8O3WfrFTPFxAdby5E+2zrcYuFhl+KIaNa/DGmUo1DkjM2MBSsRYjjySCTK5aIyb
8FQ10SHWJ/khy5Bbnk02gm0AhehkNTlrgn86l3WboTFn+Dyp5QvooCVZs9055DoTserDIj+Rfc92
YvYvzTjHry9vw5Tz1GTwiVF007ih3jWcBX+vtoedyIMxo2C29t3OdCbt6gztQ2FxAGdtV1GcH2dU
e/94kmaAgRt4y6v8nkjTDLvokNu4zFYFXZ9AIMNHr/Ds2zl5nRgFJIHAVe5k2SdlMSSrRZFNiMB7
luvil5AnIGGCRPqswpFJip4GjwNaQubP0XSnl6borsh1VAELrxJR5xV/sDSVRvLZpYF8CB+QZXFW
l3GBHkxKPTyvWCsHyH7s3hmhhE2LXARo7QDtdwfKTrIDav9F2AYvob2QNLhlK9/VNbWRTg5zJ5sJ
Bib6sP/aORP0wPaIuxrXrcVZWObsf2+7qT7MMCymB6Q3U4NhFYG/BzuB+qM9bHk5PBMWqPz5oE8S
eHkIdLzyeMY2LjgHcDUF9ND6+BidvPP+wdkRlPU9yxLlGTYYG+7pYotKvpJyWJk1iaLnEvTF2FyP
xrMzMzb0ptmRqQIRaAkutp1P1HTBkhAu/i0UbgnYmixTWOzyT8FlOh4AEdyx1GDn/5y8I42pERAw
oBMneb9qbHrYx6/A0TF/1wbgrxB7NxHkHB9Bl+D4Axh27YGUHHH6oT1I8vMaVkU7pNRf22eK8vT8
wbXQV1/t/Xlde4M2d65fbC6M+rjxeAL44++ojvVpj0aeuzsnjEovfm/0qHyXSSBxyzS15nZPKssV
1kkJik5bAJCf7q+i+4xdhtdYjhBxm/NmWzgdhfv9M3XnUsbUENZDIsyF8dnUUeTepTuxDPhQc9To
A60ie3dKwY3vTy4nWhVwBoYDbi+CZGSCGr6nBK7+ZdIpJV0rhsREOdLPY6jON0udb42rNZghpqPh
tuZdFEHXXrk9HMOwqSQdp8i9Ihmcf6BnobKP0wuC/SWChxXKpK9FB4o6AXEqXxxgym4c+cdhjPAZ
L+48vXrOtaIHIeUlkwCpJeFfKSbCyaEqGjcxMq7tyGfkaaqjZIgB4VuP/YN0NxHew/+9cirMrJ7h
eN0XISCDv65yJx/LnKq78VuAwGLqgpYp8QbYq91GaxdzbOIG97zTglxNstZi51x1rdlTeuj9Aqj7
WYwmMxhcHZKL5mlT13BAQm57G5ydcs159yKURwOlc75TpKWeXSQsUk2Fgxvf7jKl3ftrljgRbIqP
rsC5yiGGNsAUJu1T75SpKjov+kVZI+gAC1Jt/eVvLFJ/02805ZVurJVU70WEkwlJLBAZXSp9o7Ge
gxOKIlU1a6MssVuSQvE2gNf8vNvlVfWz+bq+2XLAGGNlSaXYKbxmK33IKUrQoqyVMTtjHH97YOC6
oY2fuHL6EzN8MYkIvpQ82n0PhAuIBZw+cbeQs1vjq9zt9+vwb/IRwPNfD89kpv1AnBlzL4UoPscS
VEULge6YcNnlVxSKuxpWQ6x+NIedOCfgNMn5olVFBGD1GlArNJQTGR/5DDlaEDBAetyAmCmwvIta
LHjJVgYP6QfenLMVZ7g7tXB35ooo1YCxOnXg2NOJ7/IWXdHGzfOzhY/tJvFgj0Cq/nxkWZe32imK
kLIbD5BO/ZwiTfU9wOLpmltJyNj8UlqvLluXsu8szardBXwqTZ1yAIVqYiTvCFf3wOGOweBwJnfo
m64e87M3VUKweYOONPu/FqhVU6+gdKkaG6gKAqrBie4LEnNi6eXTmdBvfYyeRYgs2H8NYiAvCmG7
4rRB9QiiYXScE0Cv/8NQFzv2qwmKUbXODEfKXJYGYGYcm15HxF8sSsq60J49mYBKmTUpfleCtyr0
JM4iBBXQCb1QtT6S3uUPIUOE5kgIzFLd8MgwXmUonrNFQcp8o6AWP3Qm9fgmbzzlOShVHwJL2oDr
TkIrssiRpWxTmk7t+iZgLTVTUJHCD4MmkkDgIB/++S6d/XDsniTEvwDh08VGb+j2vNEj7LyYsrLM
7dddj33/Wsg8i6kEYXxXoaRGlrQLoLpzOf/9HZdHEeqk0gIV2TTCTCoBIStbtI/YlssXqWtDRaL/
LTuUXwkjjihQhcbTZQved2sJAzavXyb91i2U1Pd46+a0M8OK63eLCDzYASYVeNC3fWUDwkwxD+vp
obdKVjrWCMYHtKWzCkdLl+qoQd4Jk9B+ciuPWpsUE9Zpn8bGt8lYANEEpcNmn87hstW4eGPgYA+w
OCU1KJvCpC8YsEim8ktOatu007G8aYuCeMLbk2frsS+d1Buyx6Ep4oWSQ1SMhQ9Rzp7aqXNuUzZa
+BzMdxayrFUN8AEw0b4VrROsE4dIrUH8zvA0/QJcA7nO7J91DnPvtJntzo18wd0fx+dFeAmSA3Qj
zFQAY2RMqep/Eg8u4Oxao55LIbDNaCxZWmDM6c7TcRdZW+ZnPKrx5HBFd0eDIzewlfLMZGa1XM5Y
Dmmy26Ryq4pxwoOHcBD+OdlCgx9M0fcpf1RXJQzeYzbLGFHq2/RpDzgZGyBFsA33M9yEbnOGRxQl
2zyC9+Q945N36j72sISi2itIhItdtG0V39OPEm3VdPFhp7900r7dajMyGDk14QHW+Qlhb1Mtgulr
S7xDx9rxTkACaqF2fuh5bMhIFuKqGxkYy4lMP56ahfHPvx80ePePBrvjp9OggdfanyuguwFUJE69
2905a2ea4kF3B8Ls6mM7sSdGL4+MU4JPL54HLcIH0vIDiO/LDNmshHOaMiZ74xcNPKWcIJrDmX1D
1CKFgIz5SrTsgwZYqoXX0A2mzcsdMl9yLSB3LhW4ohCtp33n00e97iaFLN98NPDygHTxSkyaTwb2
BbowEoI8KmFBQb7eT29hfYN6ete15ay2RXGNfzNT+cQ3McuYRQ6IBR51mouhEBg8wVYc8BdwhoCh
kSVNi/iSWW+tkWuF9zbSsulLLvLX5V2SveJLPEMdAuM5mo+jbehBtjTMTdkBaCOxpvCbyT7cNO58
0YThcUz6bPAd/+kUKlojnhkX2/mMLSvcHTAxD6d5bprU0e2zcIa4NoEtcLMXokEJ++r/yHGx6yGC
UCkRRMVrpG58f82v1MmjNcXyfe19VduCOjITHRLvl5KD2/dw3U7KaVbGCfi8CYJSesDU1gsnZKsl
pWWzm6kjfqYmIVGgKd8PUlRKZh/1+9gRHvxce73H24E46kc+98eTz9+fyVhPBJ3Z5RZKUhtRUGkd
h0qVSlU0wMt7oSbu7z00BC6a/69MVzW8juAaL0q6CSc7EholMj+7ZaxNMWsjOVKLZbvQg3MfGHlY
EE8U/6ibslM+UJhb6O26PU5IDivXSwy8lRbPEbhhULACEh0DG4FCDcLD44axUVcaAwdLz5hAG9C+
eZMU0QswPkvnBHkKxLpvWxtxHrABeAJUS9Brv4nUoHf0inLJn22lj0CwSYLW4azDOo/xjFMMCTG7
OCH1aaV8ycGyrmGCgn0Dp18Vjb4oTjDI+3uXFBdWFb6U0H1Iv4Klzmu5qbSJuTObw1Xa7Sk/Si1g
A1yHrhsNnjQQvkGUrU7T3OHuZCiWrMMyVT76leoS/0T/vO88TQRs+yhuqcr/HHSZ5VuFYttyXIXs
mJH91orEK/qZfVeiLzzcz9aKXbnoHLklr2RckvZV92GI1c5eeE4JXDIo63P8XTkXXZsIbjR1DWjq
FnMOkNn4fZrdMN9XKb075fG1ll87lW8W3EaMOOUnkK7MWtV2CH0tDbXZgDN7GKvs/+R+k3J2dGsc
aOX6i3gzJ7GWuOCavvO2f6c8l39d+KMo99Mn3FX703gE0avgBR+dGZ+YDlrVaeWepCC2IMg+kAee
XZdxbtdwsPSg76G9Rn9XFBqA4BuZ8gYPC1eWI/JyuRZ7yqCjdZJnnv4tCC6S0m6YAdqZ986FGrPz
LcRbIfn6iZ7PhsToVDrVadp1OacVi+TKs1o1GeIWcb8NItOJBE0QrKUk6EjZynPNGfVRsieKzdQj
gUk1L8Xd1UAGH2JiG4vjlq3msgTk8SB5YzpDzCncCG2EwZjbT14w/MkMwrrivv0olyd8uT/XVh6m
0n9zxxVu5dwUHwc97AqbhpLqYo++cHoBNfPk2HHDMoBIPTHHWxsRFBGyd0EJjU1ESM80mcsfr9Ln
x7wfIrZnTdoNv2n2IzP7MPHczVUTF4Coiq9cfKLq6vviPUUhea/fxxy+DCVtRjMFoUzycgD2PijZ
5pu2eQuOKJecdY0YGYpSc/vAO6Df0SZu4ypxjwj9z3kUJhGGsSScirkUplW4ZYvhUDbu6dUrUl5/
Mu6EPa9DZquZUilACHrgdAsB6+f89NAE3Iz+esAddaE/hLODoUziD7ZukRaNXKOHUDtgesYM8mkX
euj3GYZX6UQHW0rTx6sKz2CJ+L3hNOCfkKIiekN/Sou/IgH/xXX/CITHh+t9kmlYBe+DUU0iEWaE
Iy/X7RNE9FvR19Atn1e/ILHOLKZ+MBB5bybLL+3OhrxB5yun31DRbna4942MdQvr6MgB9eEHYr0D
77GLFj5E4/r/JGQ1oWFO2tpLP5ZIi4y17thWX7/Yx9Kv8ulwk4v4XRNL5MkhV7ERxDPSLNRAbEqf
AIVp91zbizOgc41IpuOBvfnw7+kPtRQCmaQbf8UH8rhoKizUuUmkmPszB7BcAZudwyJ+4oKcV1q9
fLv8t3MGR0WphGoVKenpCRd0Kb4embQa8v8RpuhCjZ1vhCV2Pf6DdalAvhNscN6WgOYqkATYE+3O
795CH5M55rmEG8meae5k7nNroLugaFvVjPf3Ot6bSpGpYj/IVRJ4rEUs/YP9RiuiKbVUAAkq84t3
7S+He/4SjzowkDV48GLm0jFGTeVIrP5irJzqINuCsInD0suQhIT34j45BjNwJjb5v6IsmwoAlmXD
913dCcCx7lwZD4OsDxwMiBJFeJ3UpIM1K+mqWqd6BJbtteLpMk+uPEFFgmjMv/U330UGob97Sg2m
FPcNmt8/+o3FwFp3YqQySHURngI06PAzi433pT1YWKC9fymxd8JnnBiuEG3Vmm9P8bIby/fjQcX5
rOjG5LrA7iFwvn1bKhJg8LeIFuslu271YtrpJjZ8w8hrTIDSygub6NqOA2uJHh1nOkcazcR/UwoT
OrCgAUIvltxpM8tXP/ELgv1Fc/6rmIUGyN61LKUCr8lqWF4O+fZO4RVLWU/k03VN8TqPIaUQ2kvr
E0HrmwHCFighOBrj+ekf63aossqXstNaiBytkSz47CyR2EjcHQc0wnUGnz4LTzSokyZlRrT9PMOq
XcpSc2S9XdLEjRLmDBge6SGh1VKn+HcHYwgT97CBj4UsvCtw28xkr56XiLab2dB1CUPx4URt4X0r
5u1vd3p08HixdIyPumBcJzvNnty74+irt3Oh+KssdOHTaxj/RSG2yM8LxwZINBgXrRtTaK68tlFS
/WRasprJ124L0ZF8qlvn9JP2jdrJvsRA77YQsRGTbT8pVV3EsCZRQkkmo2tEOOAr58+jYdm6PM7f
p2u/bmNXG6QNrzIIZ2mExQOaY58jugQoQyNeApIxrtSKwejz5M6Sv52r4D6uugbM4nMjp8Jq3Zd8
crvNjnvs5W9EW5vww8DcBuwW/EWaNkeIDdxFRSKlWkUaHuTfy0Vf9mOUQwJ0LcgYic+Jx4ghszAN
BkxJnaaMDI3eZ5yuzvWWPiN4Fi1eaR2pjqryIW8NbdOwFN80pxtym4uU4NMNl7SGudUqx68mh+RM
eq8Gy8Twdes5uf2laKVsrl/WThlVPjZSXOnHkZC4plODBPwmEuABzr2/4LsPDglAvBxUcDfFwYK4
iYgIgiIcU5c+Ner5fva7pBWJ8UmUAAjn9q0wEJcT4+hDe7Ulau661jCv28gLl2z5ycnnTRFGU1vl
WrSQ2LypqbFm/8FizwNGb5DGry9b205MP4VkngOLPhyKbppjFwrB2VgQ2fzxt09wlJ2BMdCCR2lX
oVWbSjSXLYxUm7/WYR22Wy9OQmnYgmMl2C4Zr0HhuvF5Ekl/8k9Zoijxkjz366p8GFi20WpUTy+z
HndsqxXcO9tvmebJfIokCpJtuv7rpYi8WcO6nMchn221jbCtzaCK+fG00Y4LyIZ6MJQN+syWA4NU
k9ewxDzoZWwz8nIOPulXUmRKhQl1Abu7ogh59xvnxd7J1uPFroGj+I16bezIUYA/mB9Um2pEkLXf
H+adDHfchpjlCRjN2P2rdNDBMKVrLwcw2DlnBrWA+JHrcGJNR/zKwzK3nBMvtsoDUKbO6OK0gde1
QEZA0gHoeOu6sKAvAG1yGqSKJTpLfB2umML7OLf+mFDGikaWdxcRiww8JnGonuRMoTohqkWJtESR
nZzbG9mLADZJdAPpt1kdoaDReVVItpbaKk+P56PGDzxLZcqFAugm8DIQeJRGJttqjpIpVcxb824d
BlvpvYr3PK3pDwjNxKKpdhLAsUaIAmLfKDwEvjRonOctL46kVrc4VmduU8h5tJpxTsy9ytWZAT72
34T+0oBSWd+rYcMtsS1MIgAMQYpTO7BJkGJMCVh7fqFkAMONr/wxu1lOmCpp6wbCVCOlXfclN6he
V5COz8KJ9Jv60NcE5hhol+cK0W2y1RxBkkJEe1L31+RCKICFZWC1V/A0Ya+3MZwN+QmoIrsrwsmV
y+mhE47UitimTz3Aj/Qwspg+0D1cPdsZkMkOnxeRY2dEo+o+wTNRBpxykUIwM1PsR+24RUwH+BzF
zZytzlXB+ZEKq8u1d/j7IPrcD6fF+mQ6XQUbwbcfRMgwZtrRGRrR+YMyu+mhH4noU7Znl9IThL3u
rxGA1xnCOQZBavIw2Ru7dzLzHYlpj+gwTGbo2oTs10nnNIPgRssf0lTb4JY/NdE95FnXf0HSkXr5
HkHJfFtj9fqwKabwa7SqhTqqB9dtKEo4XzCMkWMe1+iTHaCag2JrZYv46NMQYYKrXQRNLxVaL4qs
2lRVNeQqFuBV7cOymyZyt6hZGCh1yxtX9KenreXfCFnKYfoxDcBhRVhER/ZPoUR5EFYOSQD/MQqn
+pPbpNTSeh6lrK1ULOCMazIkvg2TJO8+Mmo9/tTYdQVZRg/JgJnk8YPY8on7z5taBDjHe3qdeal2
0fMnz/0dM3NZwCbn0XEjLUYA4gZTmsJgV0OFqhqBx/aYBVOO0a3lN/KD0xFs8D/9dNJpVnwyox4S
wfmdpu+8oBJRd+k3d9NInMTH2a0Yw7mrhMp3KUrf1JZCw6LT980cRCtg/cwejmEpM02iYtBu4CjI
bZA1q3mC/5XPgmws/fVgnRPHbJCI4AxgWyi+4kvwYxVHdANs5qhGq+t2+QBhuXnLC/s8WdqEEGg0
WN5JqBsEw1WFhu/jFjsFKTNrqfVxAi7eoCv84RdhUKvIyKgP4lkpRDhRIV3AuBy9vuq+kzSakzTW
xRNAhjbCTN/jixg52LTLAu3x47R9tUiuNLqjllOccV1BYfL3BksyHvIoo5zRlKw/gyqREqyqpe59
xnaIEqTrBgUm/G6HFqyvPzF8E5UMe2HX9XHk7eiPuzgbzuqfqKJOJbMD9u2bATBYGn/Qsiq7WPzp
cPIwkiy4W958hK85EzUm9FbepXMDoiJMnb1V3eYUjFpeDIlOVRVZZr0ebPAxHftXi3wh7nbStVVG
a83isf3jYMOG7UopJQzT7t0wLGG99sbmyNaAS/w0Mtoqxd7tYbf7/prhgL13G5tGGA499+8hSZnS
KWj1/3WVW/ai0HvxJ9/wqT6DZeEU7kOXQ4Pg84sSjKcqfK2c/2aFIfzmDolJxwZHe98KjMH1f5WB
ktfN+99NMGFP+bPYdtdmgnhJ0V2vmVQUpiuFecJULjFW6f0Ejtr4Sl03ehtIrXiw/c09e00GlOfA
86PYJpCloKhr62dRbkJjiAVjx/iS7QL8auge3V/G97lfnaL99OjkwCuwVgRXEAO4iOdZ9tww9TJz
NICaFywSeCQY4wOmtLV6yuiCdmaODm/Qsx+bpCtwK3XA8AETWQlQLmyRgIXSoqW+vkd7gMePvLJI
iBa2utF+JXHDmiNGymYS7n7tKAvkkByUlXr8b3e54r4iFQVwlH8CIsXhYXmLcYUqkxypFLqPX2eI
0UrQOJD04STFz1iCYkCbVaNi2Lkkbee302N5AQDKQJ8I/mFG9+sCp0KJ6B/g1Yz7VuseVWoVjOtX
7x4GYQ/+ARuqTDkPzhZp9E6MMTyUVHTozmFVI7f3kAKkk34ySDi2BpvOpBFsfi/eABUjaqX5himm
xIUZZqWI1XpHq4gdlD1Ya/8wqoGO03593fXiynQvhNlm2PTtKOUSxBPc4cjFNx0V8/MURxtL43wE
lrs9m6G5SIi/zlML30udsRaPbpegxBih8s3Zul8yDCVHSgXE6UgI0vMnL0gHoyedYGcijNqt5jwz
rA2mGYuDo+x6zPD79lZJsEbW8n9Vr35fsqD8KW8MeIh6xQsG/Aax9FcWBR25rTgI6b0yrDwd8ngH
5aDZ2iRE+GkAj16HlsA/Qn2YMJTA/AGRLDRSHnUnMDxsTx3VL6CXohsx9QN8BcGW6tBch0vdaJ9O
OVaiGGVicfcSyvj5IRjZbpc0s9bmQ9LbIN+2cscw54DwpiXp3cIx6D2ftFaW9pn7t7QczP03uGnI
xc3ZhQEo2rBDEgigxGFswFTGDELYGSc36UkNPwuTfYS9ryALo6sg8FQfFpQbRakk4flzeW28VksM
Fsyu7L5U0iN2XtpOR7xquzTxKN3oxREbnccyRBBLQnWrCGT+U1uukn7NjMiVLfBdelnIbN+gkZHP
9w73eCx/ucZKtTDy7SAiKTINM5WWSPNULJtYbS8w/ElChBysSDRJ0o1PdpzcXGXaRCceS/T2lRMQ
gy0C7qxZeNBtDEjS7RRk2EdsLsgMAKH0ndAK2dsvq5agK40kaHEH8BIG1bKV/ZhejT3kRzBTK8PQ
obkgeFTC+CI6L4JtQFTon0xmjXi+IlwUxfl7+OAysRn9kH4yphFYxHRcrmOHM8u2tpDl+7Z5iNld
zmJnGS3q9YxDW2B7gkE8hKuY3FdgSimWhnW9rlYuxSlZwQyiXPus6UKkoEksJIfZ0yfsml5mTmJI
OREUNWajDMyPGo5+vZBFvisH2WspOyOiz1BLuMUQD8DYN4GryPmcs03VxBhYe4cLrufJCN2cDUDM
jQhAZK5foe2IAU1TNDCCGOuK1GeS2rtkjN6tZ+5AnXFntSzTODf0JmOeuVGSxOoeA9r8wsdKzpJP
jiGNjifYxLuBNH6w1raOYbPAUvVy0Yggh7sNqPbIO2tRW5kTYNnBFBWYVZFGvEsJ3PUBEQA4CEXh
2c4PHUWgoco/kynLEiNyfP57gKHyXUUewknbJFy28bRB3pGTHo4YjMHVyOLbp6MPYBh2stTo/ygj
YNVuAbUgVW/wBEuCl2KkTGF/T/RMN+ekBGBZtHbNgzeVnKNhmj4zkuBI50UdhF+RVpbS+MwHdiwp
VGdevFg87Pj6gAWoSS8tvGqO41fcPhAXMKRwcxn0+nc0Zld4GZIanl0jE7PLoRpLalK9R4pvEHZ2
MSVmZbzi/ULPKzv7VQ1hpNbxz5p0LIqNDnZazKvCvQb5JF2hy/Yz1WEEbMvL/BHYoJfBTuuMaaHW
J/3yIxu/ePR4PkD5dDhyIKlkWHQgh04x1JhJ7nb0r23WI4Q641vfbGS2+yekFnV9YArHr1IKXc/6
8UILrSzWqjttTQeFjLLQuz4tI7zqkjaDbq1Zh5Gkykzrgs6hDIcPk4M7ccIRTH3ANxx3dLpyZ5qi
is2qKK1v6cn5aAELO1MVYn0b+1GSVUbnx7Kt6IGeJMu6jKTMPpJ5J4wzZ5YqYf8++DE2DrfuL8eh
LkNcZ5B44sF0DYIEat501/oIeblCr7BIYP4YO7JDc6q+ES2SJ7e8j9yKLNBCt9uP2Ubf5BJ8cfXl
w7FDLsI8lfYtXFhQ0OA53QHV+miV37SJ0Gxzf4N0ItlPLOh1fzjMubvPFvklwA04ilvtV9V2YBvI
eD4/c1QhVNBA+6yxuzrwebgGMkQSNusAtLJ/mkuTZ8ZpywJhqI0RV5Bzn0pGjgBiHqTJjdDd3qGp
BnA9hc/BDAZskL9Sbhg0CEfX+N2Og+aw41RyUj5nQ+XzgGrrdyQ+Q9iAKfH1t6Y1W8T4II3KBv/R
hpo47p0XePK/sx9vwW/8mK1WYT+0J9yIl/CIFqMHPHyyTjvfNhe4h3EIK1iQYUDx5yRK65Or5DFW
DDMjThDInf3gwaBxwtUB8gfHtdJWoItG9UpNtNm4GF3syuoxih8L7CNSfsmTFaTQlvNRcejlFA57
rlrEya2xdHrNpTqvRAu12Cjm8ILYd1WxtGw7jo4kCbgINx0laTs+B9SypTZ5vFh6m202DZgV0Xdy
lapWKLiY0wFf2cYT5TDZJc9fD+Pj9QhkEtM/EovAPqKX5eLgWNdBRDObt4tYX1eR0GF9tgQjFbV4
lVxcuDc4Vv4pco7NFEzxXxZoqhit+YvTk1KiQ/Dyrw+m0wgKPgxBmW89gxpSr+Tj5PIVXMMOPRvF
W754ugn2dqOJSwDHEixnxXjmDmj80nkS1LEqYrbqCV5i9nj168YP5VO0JurEPORNVn2YChnf0Nf5
5HJzAmlEtPiBSzHSFUt90kEl52ohltYXGs2mixKDci8g0apsp4BhAtWUJXBUpHyXvvP1s2UMZhPP
BXngNXRXHLJitAY3xc95dECuqBuuwaVHY0B4KWdUH1aeYvpJYL3sC7rj4zRPz+JdH+J/5TK7TUrt
ncxrvZIrShwelfsmrmS5AGdGcZFUkFG2QFPMgXVJcSNIhGzoA1+JL5IvM6wIhNu2B9blKhCz3B7z
UTdkLO2Fr10qz+ojlP5iHglRrOkxMWUbV0ePsItqMqAXW8LZMEH7SYgm2AP1DY1KhfKbB+ZAtvER
JGI6DsOPlaO1aKMdS6aAL9OBe8/DhIUigKrzHQ5RoablnDpJhV/mFwGc1ywjOqkpho7Jboaohfk7
AJA4iw2lCIUgeFkb6sr1VyjqvT+G3TLsFxrQmNifoSVTnxVqPHpGHidIDv+8zHeLuaXE7OU+htSL
4CG2aIX99DRoaalFctiHwSR30MFcYYRmE/lglZDW5XbcH9+fkNZaT+PcsLG1s5AA3AGSniOyrRgk
s+I1KE4Ivl16zTX5H81TWOgz0jFNMahsj5oFE4/NJ1ojU5o2Njuy+Brm1gSSKiphKiD+ALtXJ4A8
uNTEjYYKbRgIS3j5MGXha22vU7lZrKokEHl3GTQlLm1BMvBf+dW0z1dm/x7lmFCqFAfz4v2khYga
hvPzwX3zbUUlG4KwbunMzzGstw5QH9uFsaJK+T+qsG3bznrp5tcc7E5J80QGSQ6ls/Oi2tnPUFlf
T91/CvFoOnzakhohTcP7Z+PUrpe/AQ/7etJd3KCdJb8LTZPAIbrv52RaSeLpqt0b9PmcubfIIiGe
pKGKifNw8w41QHNAnPY5zmfbw6qV6ZSgfBCX4bxmqsC+eKvihQr3EHN2wPhxC2FQuul8LpTX1yhH
4uv30KcGNKQbDvYJ9TGEnr9eNf4AON16KBedtKrXtllkMk/FIzAqrz1at+Tv20iZnXxrjSGPFcD/
KTpUQ5HeB6czNo/nMdXSBP1vaSZxDCd0VW+XJy/iHtcMf8llDl2Uj3815nX4JiXg37sYIny16kq2
l8HskX3ojkULhGuEQjZDNsgEg6SwSUuDEzu9XqHWfbXOZb1A2GWadfcui4nADqC2rSsjJW6+kaTI
h5+v/QPdDqIZ20o3pG4s+ghbxqN/92cS/p1+Mh/rb8qR3bLLMAlbSICWWBgPpFJMsTaVcdN8+z1V
juGCge+KVcmJKILCPDILspmVmIjL7mtl2TXVxBX8nI2YufAVUTBIC1EN5es8WeFk76uz3dd+NDRj
J6JD8ZqT0woYoqqHX5EwrqiSgWTWFDq1tTw7GlAiuQD592VD1X7QUipfGVaprP3ZS0dQCiWAAE4H
58bHBwZ4s6EudMDsY4P+ah5eEPm4q1DlVkIQHDWRG+gr7WH2fcDF+FzuRyM1PeViWSgLI61OK+0k
IYKIDlmCudDJWlze5qD9SlG9prYa0UGNsxxIMUKYY04ksOW19FGh6QxHPSQ/xDrSyz2FBFg4xV88
+qbNJRrLD8nDcRPcetqAYsHOizY+hGR2eKjkx/qYkB5b12EEeUGTi9gZTTTZcZDhL91kFB5jIcWz
L8hktqrBXNWXdVw7h6v9QC/jxzXXl4HITzTvVNTdykCrMSgcq8SZaIl/hXYtSwDbHQ7Rd/waVTR9
Yc3XAOEdFqzHtH9Km2KNZKtcLxZYM4z0Lirk2s5Ei+Y2WuLJr3gLFsUCBkpWd5hlJ8uLQfYJC7rH
ulWv9D/J+SnB6Y7vDVoqmjkgaWa47lOG31nh6USI+e5gX8nrEl5QxBa6mKWF7s9nu7l7CvklHFYx
wSbsfrHnYAYjsfLH7FTewZa0tnb2gYmC+sDcLfV+nfvCYkMRcXqJv55pTiXrHqHDNOYcTyTiDWW9
+CVOy3PQwnfjpblUf/h+aweuCLJB6z8MRTOCiG9p8uRqrCKx1OV/j5zRivhRMxbLBA8gIutiRTCV
dE7nQ+eq8XFwkkeSB3SO3nO4ufjp+B9Gm2AMlmQv9NnsJIZQHPbMe5dwnHFL/KUw+jwz29PQySp5
tZQmO6UeX+vb4D8hmu0VDbmlP/PFg1SdygYjqY8T473Rdjz5BaDda+lTdlfYOjB+yQek0n8BGLZB
Xa3E7JuS1EwLRhfc/xkCZq2WrRMtFSPpo8d1xGzng900yG0125ALRs/eBF40hY//zGlTx0NEKvM4
WDzys6fmxdW7EZraKhvBQfFAO8m7d9xNT/UOQb7TWAbxGMlDuAYJWeaxm6KJwHYk7EgvVBMrPAVS
3gpAxn+1t/ZsD6g/69xHP1p5rwvV78fpxh1GCLFGuiaQsti4CxQU7xtt+QmZiVQOavE66nNZF8Qr
RoMfgOGej0lyIaOtzFuKW3dpWBMuuXgheZ8nIuZnssnbeizGW9shgHSpXcR8OlA66Q0K5d6BvKHO
JfjMMPZXV+ywBc2viETDw/zPSPrBqRl2Ve1WOE9LHQgjAupjz9WL84Cqn9h38Xln2UrHvbDBw5td
MenkjW7nHVDR21521sYuACm8cAdVKJrHBe2KuBKigSTY7VqPMT3otlHNr25qvtGHZvC0F1HY2y4O
cDS90mVakm5ahPwFKsouZqhDJxSMc3wtycctKJSnCmtNQpWG/JpLlowIvQdQOoSh1xpMqf0RPUEW
pgtBLYPxI5gKhP+DqN8SGEnJ9jhNlzC6rc6G0NN0p8cT7gVIqqR+vkrfJ3ew8dWqC4+XVq4jXJq1
SI6/R49dIiKThHPGFuyYoMvrzCRjuwEPhf14S+AjPmD1QBN3FyhDIzoSIehcijqYYQOrtzuu8r9x
BaXxY0P8Jg4Fq4V4g5uV279GnSJ2Px2O2cDun3SNQTwloweplQJFXNGcforarvBGzbSbsRz3MvPx
JzQZPziUaJHt80LCTVfUjAEBcHBQVxhuYupSwi1zkMpSHrB4/l8bIJ7dE23MnIQKBgGZNke89E19
E9eSm7VtyTM6YVyvxnizFIS3ZqbnErAwkQnNLCoBNaGEkzclpLVkjZjxCgKofPgnbq81DvRmc4KC
PI68AJTeCO14k+Frh/PfZ2fVGwCfiEqH7g3Beeu8sN9LWJaP22bZre2ztX3Bs5idgmJIfl/JmVjh
gc4lX0IxSHOZzOl+ez0t17lmlzrTt0H9NjaSYP9JrqdBK1RMgTwKD67uU1HICot0ayBgf8Xrr9U0
ThNr6pntMZWWlMKewpxcNGPkz8HooM7xxynyta7S0laYi7MBn3FjDHXh/g8ZXuWXBrO0Kpfp8N+1
t01SoGGTf5Bkh0nZpOq9mpuhlg1JfIcfkaYMTNuQeVHhkaDKgJPGNHVwH0H3cwA9at4Dc079J3Pb
pSQZwvO5diMqDwDoqtOFOmGYJQAVKOvMXGrlVgXQl9V7I+AQOecfIbuD2Brb5iu2LW7sM35XTc5B
9OSY3NYh1lS+AoFpZWp5SQo2s3j8v416q1mn28jPrYBn8W2O+q3Ive/wmpf68P+Rz9Lvv00Hp1HH
FzDP371eSW/96LQbxzG9MCOOA60r1pBe6mte0zE4Xm/Rc0KW3X/q6IwF7FpRZLJdNh8GC16IaEuv
IszOCGEXLse1jvim7QpqHU4cAZT3fIlnvTx1dqt3uCM3aFZX9vAQZNIv75/PaH9R+5UE2HdTlPJF
v/7wMAdYJALO4OHACmmc44eSYkTiDJiwCH1VcUPtK0EBmsAFTOTE8tMnYFE64FiR/XXbmoTws2kw
krjQU/qrW1hipykWzROD1SrNjsFrYfyajJSwJ6oqs0bakoQLe50foncyPmy3bOszhexmCIiDh6nd
CmX76lOuLfGYVjXVL8T0QbyD35FOeDaXZxkZUkNwdv4ax0szdHgZF76WL4HXqMLwoNbZTJbnghLy
0opS8yh4rDwIjntjBdr7ai4AwJsLGpxjWL7Zd2WMmDE/4Dy7nQqJ8NczOdNqh9QleUzFVsGsNbKX
AMaLjwcP9KF6M9ZIv45TUCdFXm1LcfE8bYEb9VneveZR9Bsiv7R7R9l3+qxVIvhgAV2swJ6VinIH
bCWeyIrERvs1VTdtDNA579xV6FxYdOp7YwuQEzK1lxN8GK2+R5BArUxL8gk6WanI03itchENEbpX
UaYl6OcsDloVbLouonNaO0eRFswXDd6+YdxXsuzL1kSd4c+gn1D/ypvFlEyF1/OXIHpNQuI2WB2/
QbZ6ZkGYCbXBJiZ2FtnbGlat9avEXYO4hwAi7ukm0Wb0V9P3jx6U0pKpOkM/F9bUm8zaSTinEcah
rGmnnZl2YUsU6NQ76yWoXl2gmMywTynYRrMgCw2QQySbOFejC6E0X9Pvt8bPloedW9H7aJfbS0Yv
oRgFER/IaPwTC+ivcc9RYZpGzUKm4dKPMqEYgcsHuux4YrKj2+12fixWGew2ex6m8jBKZZfpw/MQ
HUnSzDBbVKldp/VFRkZGJ8SjNlOc9FtRqBU8ZIlbWgB8dnKxukYpYHqkUA/UB0kW18zmGHhJFYSv
oxH+ZXjV7Q4y6gPfJ5x7rbwZJwP6M7ZDLUz9c8BxF/K1hxRIhyUTCVbNicG7Zz/6k2OdMfVuqK/D
uOjP5EasiKbZF8BdDy9u2K+4DPchQwC7R1zfARG5Ow0CU8BeIRXK2pYe+e5SEbgygya4sLqHo7FI
lRpVbOlctvKtFZvf908ZjeKOrG308F9TdruFKBkDx9SF6qbY1sU4nDcS3TCqcHyOUAPxu3hp5xvy
WF55Cwi7pCC1mOXScJ16LkdiiyDhebEzwc8hkcmkgvQ+RJteKZxeMI6Jxcx8msP50dC0Z+93Pv6J
RdPOfrXLO8oucqDOE1lxHUPyuHruIN2qaApsWJJLQajrDGQKNr5LFqnZkHSroxQKfeaKzBWIvaew
zEZbDWB8vKdvajMdh/L6kIq1s5BN9XSF6PbR3416rvV8an7DpDwCTklGWO5DqY1MutqOu4e/h22v
4eqC+rdW+dEU50KxeTn6WHx2/VD73NB+e/MlWVPM7VrjO4+IZj8BWG/qqbeI2QrolDB93h7UfLdI
XVUqllUOQQNQjg0Uwzwua6kRS1oXJnXeRNpGoIxnXfPyXZmq5uGpZw+ZZ8uY8rMn+0A17S6xX4Yk
n1HbT17n8el8abWsaVp/hNtQXUyRMEoVhmpAA3lI8YV6CFq9b84eYP6m4b/ADaKT4n3raobML9P/
zpIUh3ZeQbw2XwrdeOK+Tj9EqajptqbiYZnkbW52RoaHjvwXculWexfKwTLO6qSnN9g9a2fH7VLw
O8WaeefTiDSHn1z3HoQLwvEW0A8pYSqgwbZ2qaKhyKQgXAB+M9Ha4TiztpuWqi4f+praX+ufCQVp
CdpGu2VBjBNalQHlY6IC4gfnUakfD3OntN0vaVdYhBexHVGSc1H60pneqkFuSIQnj/KQUNpEwx9P
MPzQKtgtkZyIURxLGmJihbeFWb1K192JZh/5iUzS73mDJfLdkXvKVXqoVNbIhRcH1vi2euljoUdK
TzCW7o+3pjB/Gbq3c/xi6FC71uJm4gBrkYRdkC2H5y1kp0e7bbLNYLhlyx8yIzNf5RD6SL4/roWU
+BR70Gqm5d7rPCAdRts3b3lVkR1yS0N4Ciex5aCUPLV6LT18E+txeNGzSLdqE6Ol04pUra3JaA0S
tYH+4UOb62N6pmb1OG/M86OpZVOgA4wd0WfQYzOVDp42I6fROuBqE7eDwo52VNrZFsGCaBI9j+N4
Q0Z2KUj9RFH1kP6YaXEoP1kt2QvGVt/e52Aw0TI9zq4sVQU/7AaGGqeAmqwfH+p7Bg7FBFD8ToAu
0LYo31sCzLBLSG5uSlhej4H3USJ6jcWvoddqXcjU5DIBC+CB2P0N/iTTC52HpQ8cxSehbIbLYC9e
X6wwX6SToDMt8O1Ll9VRxnk2cirz71x4OTnA4yGEh1tglTFxNgR2oqbvEZS+VnkRqFbE6hIfOfne
oQxwv6c3mMu3Piw6EiZQV+4OgOAC7HuPW90pYaCv2R8mY5okai3EZjq425y8ykZoHGq1y8rd2ulZ
/2cH/xL/nDIeqx/XqTRChPer6SjXPuMHp96z+dic0yZwEGORlGRDHnLomuTwcwnvhgfb89E+l6+J
38aSjf7OPKgSRDDG0A5uomiboNdETpyNp1y4f6zOth06h19W/DkQ6oHY1qM9fI+wxYO6VMyikQCw
o4ntX8T/R1oojTfiBnt4TEbmwLiRyj/tebh0/iVr58GrNpbUjBRB+ESLv00GFDPi6s/j/j9+fFDv
E2TBGqM85a4/YZmRjJLVZkRx3cTtaw7Y1GJr8XvxfEvJMgDkZdZvC56dEZBn9Fk88or6jy9/DXYl
yIK0mr98psdP9IvM5g6O8L75OPtUYH5Ep6H9nyxh0rBOD0/CECR/alRh/xO3bHTjIJUl7pObeecQ
a3D8DXVAxs2542DlulmMham8oOj+F93VxoKbgTeFjen4omSbqXhq9iZYQBKOrerRQb/LgE/W6GxQ
pfNkPF40parPHmgApcLJYGIILbU7frkwBdfsBco3I/iza7Tac0L71nxsanDc8k3HVpfrkELYEmZE
xaQoJBHwgAsVj0TW5yw0RcbPFMA+G8SBEDh/5+hngRuGtmH69MwwS/EG2KAP1SgN4Z88OfcVLlo+
l1H7/mbzhi83YkkOUgR2S2yopkkXWQy2zBvPizcejh34W9LR++Fzd36DjAQcfRFXnHmFRymsqZhD
/ALp7zNFl10MaCgpCeE8PmS7YdS0l0WWM5oE9x66VTdLDUePFL4+hQPz7FTGmRNmTGwqzMQVyXAt
2z3YwzEDVkFQgm6YcPmEnXfVPZyjMSD2p52iABteUHvpvcnfaKnv7rLMLH89r3It593KIlnuSKme
CskelReqpUqMmXx2KaDXWK4wmtWxb5wLhpyayNsgIuwYpbKBJTNw3mtlRiDNgqRxykVokGmIPUJb
ob8WiSl3YhHksq9kabTbpIbSV4w3laHlZ67LJOodl09pN6DoGeCoj5Yh4q7lMnAEV0guPCw5PTIQ
yhUfKPobtK2q+xB2BhyYM8r63/SqM64UIrxHl97UiMfWBptsScHFpBEzxWt3uXnQQs0ixZK2lx+W
7XTLEwFVs638CNPm+sqLGXZyiE6IMTOMi1v585I3lD3xrcv0KBmZu0WoStpqEAZD7TNBSoCL7BAT
T6RWcUaYAe685857IQ62oXsVT7xFreZdHeix8moSAyaSkJtUJ2xjayvnr8LkubNPl96AO0Ju+QJU
citEr8hAAxSgBSCw0+iITpL30ooO3ktDTAioiW0wYb0j7l6Wmd71RB8Ufuk9xU2Rb4INQdx1aY0I
xj0RhIFsolB2fzqtsNEvKtI7+UzvV5J+a3zW2euRL5u4eyLx7bvdxQP5q1LO8mFnqaYmQXUprC33
GsbD7mV+WCFVNVUdPeGQrpRm6W1qkp0qFE3XZzgxfx5TRiGQzVP6McCwdC3lSIgrPo9SP7pnIMJS
G6Zf+Z3p5VLzfsnCyYuHgyuXvYnXMTeV2B+0npaRdgZN+oXGe1QyPcNzIREwszkD2wI3L9ESy7S1
G/q9R6k8BLtpm42ioGydIDMrrx9zXM+JBtmr986TnRzF1FyABbkTu7Nlpis7xbjIvVxY3916C6n/
Tzq6NbG0lqwmBup8ODTR4HsKHSboe3C+nTsSZe1zePwKZ0VkNHQ+6HwX50fdZrTukST+yUj7eteT
WZFSJEI4h1ikJLCiefCh1MauxZpPnxT0TSGClGFT00EECa9UmIZNdYDKsnZcKTmMzudc/cz8KUgl
gQ3s4ti9optMXK1Um74/LOOeeDXpcVicRlMp7LzrqtVoD7SYHXfQza0Zgq1irmWC1dd83D63hCwV
bUn1+UAo0/2xwXgQPPKzMfmR+4r8mhXs/N0fFXGVOIghS0oNwBaiRbTX1bgDCl+VyPSjvZfVfxRh
KFZruNrQZgw+5nzsdEXsM6khestWVIPVVBFQ3BR3umMONvILrDU6cTeAVRVoOEsrvonjETu49hOa
xBzEWX5qSDQsKTV9q2tnl3xJJF4KUfznU1wPshrrsKAFAkYBMSQkNsPhiXaW+Vcw3UqF8T9h+M0x
9kQLkiPI1KgMoDvjfu0t9udI49PyQAnzdZSSQTX+MYus+XKpB3+Qf0ZxAEGv5qe7dJmyCDqo3LON
U0lWYMZqnMYByxeUL9vXDoOq5eTmmIDk2MCsqZNycSX8X5/0wcXRyPfSt9GWgJ9t1VVmmVuvN2ae
cNgao12K90K+/uPHogIs8OSvWccEgfeAISqKh3dESg1r/Qi1IQuRqHg+k5KF47VlRr0IY5ggZERZ
Y1OJ2h7ZSy+CMU7Z6B08XatZFchr8qj1rjGiW2cKw742LUlKB/cEUURCvmKakvjeUAF+TTx+QNty
8shvtzsGZoXAvBVyAG1O4oO4Im96n6WGDF8Fw53o0Ir60sa7GWws+VjgC79Ij5LfEvzKkHqBLsLn
iDM/0FLQGDLKprFouja5Cb0zzR7FiEdXqlCk1pLxYGKE4FRxDEhMv1sSK1++KXjcLXX4jw0QWNXW
54Hrx+lubNwoGrROFUry5kVRKZJBhD8bsS+iTiayHpnz3WM6eOlBEEGamcIigtV/PK7to7x4yOAD
jnT7Gz6FEPXzr/ACus02Pg7TpGS2x9WXvXJueiBgOzbqBoVrWdZaTuk60/c/ab62c5GFkOJYkNit
cVURt+Me+TNIGEfQWPmkjY6dHOvBrhe7vG3kufuB/xOQIGPTxq+ApT5x+GQDjubes9Qbu5g9M33Z
80N4KWMDc6EunW4V2br8sqqZ3dhIK0JEHeUnmE+mKwK/ch5rtPEUARmiEDvo6Qp00bpYM+WMFTFr
RXX6iwGUUNA3IYQ/cJJ0wMvqru1kEWt21/p0SARS8d9CXzBhVf6q6SS1vXXv2+0guMBMQFiwvuSi
NS3ZH09N+yBdq/0YW6y9cDMzMRPCF5bJKNUklCilIRdNwl7Hcw2XURYnyvHup8kC83pLZnLN0fHW
iSkOlihHJ7PRIgsHkA/I/+QfW1IINybhqpW/LipQgiWh/L93kYzIAp1DLx8nN6hNIayXZSK8MRk+
aAsMW05AIzntJN2Zqj4B4BZnz7YDGKn87YYATKx73C3ViBIkVtpnUvg0wV541cM72Q36X9juC+gV
ECY2ytO80O6BClPalBCl6aOkYOyS6PgSVuaa4XIQOPtbifumtUfdzyAehnGKiefggdbe+Oi5X92+
hecLNsvUjz78IXFQePhry5hxgflGfS0tutaeFqePlNS1/TBJEsIVnlM9KsojZHM9A6RUKKzIVWzN
JUJeHAoJ41KI7ZbeH04WBP2VV96eNEqzCjCP8sf/R6cH3wOUtW1kXs4LUWkCX5V3Nw3gsS9RdpKP
W6VMwSQEtI6pB4gRfSgrj3uKlO5vLoaLC+LVPM7EYDs73ZIChel9ZTBAhYWMx2JZBRYv8hvbfqza
kU1NTPxBoh+qKL8NM98msly1o0i4JayrsahcKtNTO6maHcg6ubgNZYRS492saIeqtd+PfernXp6O
GmJgdbdchHhFC2ZPMMlhKZ5apxrRWg0ulX3Dq/+s8qxvEpHY7vVOt3Sp+dWKY9Qsd03wkXKOeZAR
1zAaV9Ifzf13MNLMzpMhaqaShff6IPk7v9MogX4F/c5ZKVJbQOp+vGxDQun8OSPbox4AT43bM4ic
T4A0s9T06iVvKJnDG1OgQv8tqj4xlV2dfoa7iJOta5e3j3GoretmaizwntdRuEu077DjPdp/RM1p
e7cugDD6pdwis5ERopuGz4yi3koSnB/rQiSAYKXUKm6LkLyOKFf2uGgz9r9e+MAV7KvmRXgL09UM
MxXk+fK7T1fHG5jDYVXKwcvc8hNfKrTAS8oUvWQ7INNYTVP8wKqEtKBqLvQxt/32vftzoD8bknaY
4NsyL2rBBSuzZubMBiB/d7DaFlqDs5cqtu0+MkA3ND6xL1hSUoAUfGEd06k/FQbYoneuIF2gz+Ga
mmeCP6s95HjqHJLlnN27g7wnlNwkEbvT2aivgLUAqBtc7ixdj1Bixr1X5r0qI1MXFKZLLDcb8MnA
LUEd+u/+53J87OJ8QtkKeL4Daev9h/0CAXJ4qCX0oCRtCSfBn82mzvhpmFOr5rL52RMjcPcDgtag
pWZWitmHH2HxjaKuW2fqRYccaRPsqtTy2X2REK9vvI5vomDSQCCDHqitO/DbSPjY5BQEZKKc4vmH
Jp8NsHgqldJf4XaTeJaOiqXDp22UBz3tiFnNl8kWM5GhMkXRogSW/IPeL+mX3hAPxcKMqhoAFpYe
WlPlkPfW0/EGalzCQnBSnuQiBbPZiJvF9xc+sVnpDpDqufPogsupFFQh8QTQpsg4h6DwBYyM9CrE
nlbfjZSmuf38FicS0nD9m1Ujq3/h9gxkz09NJ5sYzB/ru7Obn2TGdnGxJlV0QmasevHUkXnrvRgx
cuv80P0bjQqVYjt+n7dy5qQ8MS1uW4bGuWEUMYEqx5FukFGL1W3Hec/boshPO9deW3TPYtmLe25g
L30UiSvBw+dre9CCQarM16TZ3e5qXfY7GOVCBP/33YSa2y0lN+AURL6Wz5eP2uza7zvvLCetNHfD
ecRF3Hs4Ur4yp+FbLh1BnEwfJImY/LU1FDvKtG1Qn23mX6i5Cvy8gj1Vc+nxKF9HCIdu3cAI5Ehl
Z96j9CXZi97RTc0U9Ae+6K57oNmDPqhtwr9+MiNMGRRMa9cnGyjA5Qs2Pw2j5RDFtYLyq06D4x7L
pKgvkbj4/dL8/t7bTjKVVFwjVnKzNejFEJBbu8eEIFkb6r/34rojXhZmyxI3ijGbrRbGJZtqWZQ7
amC47kcpvSsGrIzXKfKa6In+MfiGis2REIU4G2J9ScNzUTME6YaC7PC6jwDvmSq9kN/+FeSIZWWn
zoQCuYCNrqHL2FvdNsgemJvNLB0M79U/uCQfAUshXZf3wGPOS9Jg18JDV9VIRauX2xhYylPwz+ks
4S84wqDwpMdC/K9yIufy5D8GL96zHOXVT8T6NY2MmOap/YWqFA1WhGrzC+yp62JqKxTqHaJhY4AB
dJnu3/iGLgOBpGCpk11KWIzzLHHYWjO/ZuDBNle1pmIdN0a6sYAoD5DtkVil2CrAcXqgzAX1KQi/
iT6b8QbZd9dU9FruX45R/azFWZejZYMAGei6Jn4jJ44pMVMar1OCl9XmulhDzYbFZmUKUbMS4Ohl
7oFwegHBx/8cQLXzCBJ+VioKqCDK/aIsk9YDvfQK6L1aEowO+yICO+qjhIZ2DSqvp6g8H9NOdV59
zn15yKB0W2cgVzAJKKglzY7ENuBn333ymKUxwmwCNMHHZfGp0KjDEwjZDaryLlEByxXSeoxwJEH7
nX418N7Ct4/Qy2qWwnC2BL77mDu1EIaKONIK9NfckQQ4xGsu5d9RwRwaQu347waK3lcO3k04qSHz
/abxTH1/xtjJecMBWe8U6dVrSkJvqCltJKiF2ja6UIgMI8XVE8NlnvXtzYnrAY5gIBn52Yj4H8dJ
HVqsJhzWrLLOvnFl+UGtgSro8NYclGL8Q1HBWChm2oGpEUcLq6q1WW5r5709lwl5yqEJx0YSYtgs
5p1/mhDkmyF9Mmw77USVScKbbgv3+vrti3xetLniW0KtpGzFbCx8cEW1t3yalS5eDj2eau0yyE/b
o+EbIbBWNqo4dBrWPNuBQc6Ui6pd2Z5jrhkb73Yh5aHwlNmiz0tUf4x2tHWLFgYZgmh6r18jHHpY
4jHvr0D+c3T3Ocl0fVRdwv9ZJjn6vl/jTBzHvxKJF2WBzr1TZBFEIAdDl/h1xydpoG34SM+ml72O
MmY2SundPHB4V+SdVy0bMkEym5GxiPC6ComaYUyiP/uaPXJBQmmum+O63idpxLSWZ4lM1gcFsfe+
TMn0kLWvpS8KwvwkEvXMYy69S08U+nMo10ozOokpD4bSM6PaJig2E0r07L4tN9INwQnCIeFcCnGh
WTOsTTpAeZDiFdiiwQT+n9eMpk4dVKeZ9ugGYOrcJwxOlR4qRb6aWXhn5tn6VE2ZGU6VuPqIs45A
ahThdkDUBpD6pQOD93C5Qrdpp78r+GQcKWYWBakdu7Lv2vwSZvj038d3hrVvNbKuA0WdfzISZUBg
Yj10n6XGfg+nbf1pt+x5bTsilKRNevBNhfjGEdfGXL/MgywWzvim889GSlwujNDIokntHWER4hiK
ZQEjMLnggXjaywFed7Ep9gtNbHZ4gdC3ReheaDxXP5sjdCjM7/Dzz326o0B0Tb2J++QnGdkypMem
p2niYWHESb/2oFNXVCA8E05azozxaaWuoRLPLYZmx9KY279EYvwnFAYfxpfc6XrA3PFsyhc1hXOY
/TpaZX+VF4/WBJKT/23EAOUHUiTVUSsQ5PC/xrvJt0qDsoHpCfGEK4r2bBprbKXh3BQVLr4SkAl2
xgC13p1rPTPRh6sNZsm8aZqVPHOiwekCFXRZpaPNyO5yIcqYDa9384VExAK79W3skeYjrZxqPgpL
1O+sQWxNlcPOHWGY1z9zgnV6AL8Yvtlhbsc8ieWcp8NqSyh5LcCRaGWPf9pHYAqpAIpxlvbn90BF
0epcQQjf5G9rps9079h19i5KacIz3uBzrwoUSDR79Puki697nQbfIy3gUsomMixHbjxfZ1QZPSoQ
ug/8O1Nq0pf/KdawJsiICG482eAqkeHpGRVenvdov7XVEdjrVhH51wjnAhk676PNlePj2fEuWcEw
7eDs4C1dqEmfSY59ZRHJ+JHh7AuIIMr6DThDvB5zn8wyITYwKfvQojdVn3bk/EsBXFYOW6mmRx9G
T2E1T7sYBJ00SKMXfsmPctr3vtjhvJc0XzR6OyKwbQ9phf34o6esJ4HXE25hSy0tG+0kcZUdq735
MkatIfr4QO27rxNClXKfhp6wg7XY74In8ZnvpKjXOzRvFaVTaTqFQ73j5Bx6OiTv8iOryXinfz4+
1X+13VkMAfN456hyVBPtWide3jX+rYaKyOZY+POPn6c52sospNOepjGuI7kSt8nsAwJMcqutV6Gf
ha4Mm5k1xPYIXwBYxHOGuPQv+/J/xrnC27KS6//zZlD7gUP5xq+cUJSslfKuKVoXPDbngwNKascs
lXxZRYGj85Bzlwy+ahjDeZHwe25teki+CLWMyjOGgd2JwjY9gRKylTV2N8sof09PUcNkiFBxgdLA
PLpmL/FSLtaRkx6RN6PMbsl3t/XWvpD1DZsBzDXF08uKHG+WSxx7WnGMOqIZ0oqdVlW2/f4aruP/
vA4c0efDOdSuqZrjdhH3e0qPDE6TsYd9+lX1iOEhIJt+/s5vWHvGPmkr9k0qspDUZ/MPX10gGZNh
D9pEPw6wYZvy46jg+Ne58jwkQns2dh8e0Jj43VAlIpjaRzqmACDXKwncQzXhTFgQdac4iu6tsAee
PdijpKqsZSnvgjKL4UCij282ffpYMeoXX7Rp+9L3R5HaH2CrH4SE9ov1EN/qrAgKXI4hdc0uZkt4
mj6G7OpD24lVwny4xfDfK1/wP25h/kGVw9jQ2CrplK70gqKmMGx+k5RMlfFGLUZYv/1WjDenQYhe
MUjfEf7uVVw1vQUCZV+XtLqBefIFDEPdh9Z8kCMFCi+3aXlojmx2PxGdWjvU1WLPyuHtJAZx6pMy
UnvZOb+8oasjGfYkVLndgRaqvuR3QqLyXkEVv/ruNJdR+AKKMf/2i4FMe3hWIZdPy7ppWrM+I5BR
l7Rjn/whdXY0FT07WQInJN1viWQ3kHGiSQxIsPpnp3xSqkGY+DOyWENUbWuEeK803XA26x8Rw6vy
J53vPepo0w0EdLARzmZowVzkQmdVcI1dx8lOncAoticSSP6eq8D8EzgX8nFY/NHphLfZPP2gVkie
dRTiARFWGQhMSh7mCSDdW9y1MzcrNZrcmvIiyZQ1RLM3EW6K6FjkkBHIqoBN924W/hTSg+O9eAjN
lXceS8qejYdmMPUUPRX5gaXqv9fs0oaXe+r9xdUNMbQvf1yZMJwIadQVm2n6Dq/byfur1PYjopD/
r1F6PFoRKNOQgYBB6CrdMFkdE+3Mco3fxVKHAid6dhMqxPLcxr5XP7O6LS8g2Clep9JzWi9pbiZY
o3rTX6ZxsunTWE7amn7FdWr9KHX7ngYn8kQbkyDzVKGx7s5JxC+ivSpo4Ez2e+za7n1lZ+Lr1hl/
5oH2TACwCu46NHEwrMmDtFdbQKAWA6IPKR8BdMFNwoLpUcoYPTkJprfsIf5P7jvK301P1BC/ZG82
hDryZO0FIYFrUFUvnmu+Ezv0nf6lc4VJm5SyDD5XElARAi8wbysepgP/JhyZjaX997ukOWsiCeQH
tlSfTR9YKTQlrryDzrzBZJ9nL34BoVF8yTcvRpQHjYlmvNncP3uW5tqzJfpStsOKRBkum2ET98l1
wXMoSydsqv8ufJCgikdHUSxi0zCe5iDpTAVcC64CHoIYb8L/s25Hyjetpx9vM9VchMBEh98ONQ21
y3z5uqAVY2ALGeVGTTZxejk0roVgxfYp62bbAYko/7z8WfnqcIK1o4aZsSCGJ3eJhGRJF6AqgGfa
6uzd9qGMUpkUAd1XNK4CyY2rr0b4L4f6z8cJGoONb1d+mxvoQqkQZKcY5BbFmdWDpkR3b3SItYc8
G8wLjfOlctbyXUkfAxheSX5VkcbI43XBaH8+ZJ8db/e8WnWHLaLfOgIw6eacdC+yM/jVG53S5CMN
Y6sTckw7deiAlOiH+rvAQMp+WLEbB7l81UNxlPdx9LA13cG0FXHzcSkAaxB06GPvGhtwYuE71CI/
71iPz+V/qFrN/wBKyNGJR23DyNisdyTwTUaCrET3D5msAsYwmQo6ZU2nD5oCXKdCAoQyRXtvDQJ2
W5ex15axMddkowCAhmz4ldNs8oLF9t9wsMTI1mG73Td5+xhcK3O7smuJYL9THMPPbNdh4y2xcPuc
YPKV7LQ+0qy+oYDgJeq6yXqSpWcNMLIwkZHXkchufIjExzCR2CcKBVyBrIozpQdVfCQbBUbidudx
b6rLMax3N2c1tL5RoXwFPCUUqTHHqXvTgyvZgl/mQNm8ONpv2EOTvLy/1OBRvceaBW1F+S8oa1L7
xt85Q2f0neHf+foFZoTTzs3kDlgh1ia+Gvboe9j9vib5aThbFtBgeyTzFn/K+v97AkfZpVz0rbc2
7k3cU+S6CHS+K6NJjG7wxbzxcImhIvmaadJh3/9I+23AGgG31XzI71cezefA0qptcB3yRdgPNPfV
lwQD+LBV6KqtaspvRgBK+R/qvfwFdGIzZpv/twyRDvlbbQGCgv7QUJjCF3K72sf7/DuwrM7TfuEZ
49mYNarrojV3wN4RgtiLyhbIVFHTuHL73Pxb7hIVA0AVY2E+Pa7YSmKmPwy9hMvSDjpPUH3oobHh
uSEarCJC+oTm4WR1bIXXw4fiMGKoxKX/ygizUT43gLtkUbuQl+ZbPR/vs8VfLyZycLUvIduXBx45
fZgG3j/AEz++1ewi86tJWrSaY6g2/7cvKF/NuN67AN2lSYSdRPbNQFPJaxM5Z6fU1cMmavpeuSfu
iE9yK6mE1CovNHxi+Z62bxWMhTvNE4I/5sZGz5sB5+/dyVF6gvD7Sc/koxEsg8N7hhp1DRPhVOCd
goNvPPZSex8WKpWKgzpQaCxWlD8f74LqL5EO1LxzsSigCfQqWuj9O10dsBjwb59fLvYcP82qw4/w
G0a8cFGRcuJMQUr91zTa52TSg6bX1S4QKQj8ghUreoiws8P2TqjkCf9goEyCJDXmvIuSB43bo/eD
lk2aeu9Yq/e6QjQ6eZ7/yOcWjUJfEN3YM5zSlV3q4jAntv/XwSynNRdsjiKw4VF7Rs8BNhsXOcM9
rcZ12/XOHUf/yIcme7Ua9i1z6M+91kBOi4pSkyFXO4QzQDi4ESokYdkzFBnbC0LJ6/D4UfwaQLTC
dWFVyAKKYFvNQ6UEyP86QWSH78C5w3eXqReGZ1PmeqrCYh2xqMy67D6Gl8aE/7RNKzYhnANYCuEp
qvaH/JH2bMu2ENKIbrkBwL29xKDUKfNHndzgAxvSp4Wk1HsSq97e3qpkziEqN9KvPn2qJ8z0MMKu
hbpZQQpyGby2b37OdqiLIGGAvG0zRT4uBvsYZmU2E/xRoE/8mmasnLRMYg+KjjRkdDJJJa75x1Yi
q6cUtrg/ovxW24s7Qnbnsqf7L846QRqqdRos8G/GZQg5U8G0VD/aP5V08twfGAuhOCmKOclX2NT1
IR4Dl50T9wT0DfF8QCDX5ne4Ls4JvRDsObdoGk9MNjSaVdmiDuIaSUNoby5kAxOK+IpzpiM/h3sp
7kmAnUyoDV9t6eDZY1qbG7estwls8ZNc+YqTbRLLPBGwOB7Lu+r3mvyTOhKnCruJkL/5+TfHz8mU
05jPSE6Ea+TVKzTMBlmXaYN2GT8woetxlI77HIlLYZiAA+6M1OhXrR3a8MUGmNV6GrPTBBJnAtIn
H2vsYnRTibo3ERR3J816SQNoXc7Zy0C9LDUhvjvVI4pBD96bx2X3b8rg8CpzZOecGYewj4xEuowb
F9gWnVHQ32fOrGywulxwhPN0R5jFv9etDUSYkCAc875KDydK3aWUy220KOpbccw9heV963X0GLOE
CtNmoHlH7sDuinKogfz+/1hCHBvaBCcvQ+jmNCy+dENt/m/cWNXYqMu5/SfuwnFzhK5tnKCzCuqX
cDTTR8n1FISYRonOXPrnDoMAvlejvsguUTRiEQXpFkznq61x4M3huHkLWahJ3DfQd4BOoZAx8sd4
Xsk9vQCyFDIaTXB/1+RcSsn4bcTnn42kB4n1SteIbbWjqXFmB8hx8+GeChH3OmHomX8xxh/1tJf/
3a50HOz9Fru6LgNEzIa8Z0ntJj972YSf3wOMMOckpkwgdJbGFa9kzLkchNjGhTn+OpWXkg0mskcO
uFtc8BCTNp7xV52EQLrcW1lsTXbUDZaUl1tIdsVBJK/KvR288y5D5tyHUDBkViM6DH0wX50B9oS4
MRgWc7Ei6vxIXHftlKx61vw07JfRN1/UUgjaiMqF0JGrNSkMjwhuZmfL2KAH0BeNDeMFABlR4cwt
ot5Q/Dkpt5LR/zkxvlkAj0vGq+BUc1TSlaWitxq59LydxyfOe87Y7eR9A5I0A3ZOHi52+lPdH8jB
fFnFifhfc8S8F/2JVPb4A/q53I6fNJWlgwTTIUplBIGtyUOOQpe3xYuMJI4/mAHphNidRte+da8K
1TDGv9cqbqIVkVsMQ4c7SKztgNSBeX9SGBQDT6FTlbx00sBlY8AwcUk2NUpSAqGoq+kwQpkQqJe8
IaKiBeIdGUsgJzkZU5Au3r+9AFpvV0/S/n5y5N2aCJ76CPlaDK7mSPFya39hYAtkg6OnR9+uhdHF
TMc9SczzBuBjaoifCX+yBBnCoqyIJEuO8BtGEjJyLCPpZN0+B5CeSfDuRySTjsLQswMi+jaLidBL
v94UYnxddFecv2ER3SwHJQ9MU6MhayNaR0ZuONzL/NQd6nEde3NlctS4cGfbecmkSwg1ggTgl1K8
D0YTV6cw+sabjKX3WLXItYDYHbphbedOfW0dk+2/QMvsWyWlkZ48y87KmUDqmIzs6ixwTUndldk6
ZNgjY4rRubJaewhxaj+izZ7AF9cbWCCAGFB/1h/Ily5i3Z3KpA6Mnp/5Lps1BXDp3s/5vYv/5EMf
0dWKcD6XE+mZBXPQIMV5uCqMJDYyZnr4hvbPDiw7EifEU7MNuM5CaZNL0KzJ7QDd3BNAoAzWe2HI
wHbdU2FspL2WZOEhGeZlbuJwMQhfCIY6IOZkT2xoTZGT4pUDb4tsfjYh8c6FP6i7mwp0NJhb16kK
oa/yzFPGtKuy5/S+gZsWXyNbUylflGdt3tAyGeMwlMJc/y+38wkfSjBfLy5taR5yjRjSyO0QfL51
f8TWDGkXulLb4UbLI3QLlMuuSU5NbpjzNG4wDAXeKKOR6VFVf9ibp7y2KT1KEDR7nx3nwDPaA+N7
1NQZPCmL529QwvQUPrnaU7VIyRlfhLoh1lajFeXud8Bl4vtMT+FzcqglgP+zmbHszhpxT9bkcOSv
AA5GEhbQpVUpHnHUnsa85AV6OcPWWoGmqgJN/pgfJTJWa6gTyIEB1lEdLyWchmf0MwooR/kz+Gxp
1evjCBRzeRuDofEHR7kiRJzi09bNp98OpgvxeoQedFCrdvMyaSfaTYIlpAkYQFq9EZmY6VMBQv7Z
9t2ZWpbMYm0l8v+4V+qHtAKhsYfUI007/mAcwn3kmEXYmDv9vROVhhp2tPaILA/ssvialB0JgGpH
b6X3f4BoaWBdgMKOO5dyygpruHm1gpoezkj+sw0PwuZc/42b22YSHl1kL4/vlmFrIMKkTQhnpfAW
uxJP14bjple5v6k8QTDdWHO5GVNJYuTNwJdtFW0fgmieoyUY2CACZOrbx0g5zk2I79oITmg3Fb6H
ffop6uem0TqK/gQl62OxUMg8L9ghi7Sy0WcOB8sEePwt0maL6bVtqdbjWVXZ1g1LQg+LJgz4zXTx
h2W8CXY1It4uSbzEWQ8XzhO1QRLnupRjiPyJk292FGmKQTiJyAyMdoIlpbI7Q3U2ROs33X1y/hHe
7TIH3oAhlkzf5RcVOCIPa5Sjz8ekcP4lloCmKgKApUtBpKSc9q4pwAXjkOoxxJb5Z12NV/xYjVEA
QSqU6jV7E0rtW/OHB23Wj/BWel5Iwu9TFNPbbDiCkDqKwVcfKiETijwdiKhBZA4jaIg8SjAoCAFb
HXe/unpDmpOT9LbrhYJ3geOGzhqxLIIEi9R41SEW3KDN7XNp+b6lLA/MLypypP2T5EIaEIWZnOqg
AN7tfyXgZuECusI0W+tNVI/sQyp++kqkqx8gdn5inU+VqwjUqb5CCB1gLdk1ceXBbF2fW7hKcAjW
LIC8CDR/H5337JrHeWpIqugyDlXSk18cYW1dkOsCId/65xI7kQBGbJ9fn36kXiBl69YB3epxnqYn
cD/HOMXpsXq+K2CQChj/mt2eFF8MnbxtAvZQI9MOpeNvuyC0fBZXllxSqtJmy/6SDdNkCLGWhWu6
uMOze3Zy1QQuIfWknoU9lj4e1jK+362/Z35HbtaIwIiv3wi3wzL04PbzXU4++xYvLd2U6HfTprB6
xzryM8T/oLXZGb8kMuSLtCXDD0lE/m0T52K38rFKG0QhvH0c1iizKHr5YgUxVae5UnwAqDilYkFX
X8DH1vI3DEAi0bA7ScARlfqeYFwhG2kVz9S9yCT3DxBu6imHB8w2Y6fNhCDWeHoQdUuUt9ByqAnd
//CW7Fo1Mt+mKbDBoBGVRXNWqktRTJ4SzBsVbcqak1rL9x53T3y4n3AsKl0C2LLDq+zJClf0ASV0
of2NIfFmpSSBIRCaNNmwOS2YKJSlpuGlA/Hh/pcClPLWOXLKMWuXVYx3VpCmGUAHGbumunVVcnvK
CetBCQLfTs8fydT93v5OkC2e3Jp4QpH2xWoxYSHDHVpQmgxxlLtsWS0ZcT+k1j7hjNQovkD+ylsS
Q465EEPibbqs6JDWri2V7n7mBnTMG56cxm+YrEG3H0dMlKbk7a3nEGbbimQtKiEbXDgV0R5/KPpK
pKWiT5ul/VmwfTb9mEAv+hg8MAOv0HrB4/O5dLoFiLxu2WIDoskfjJUYSpqO5St+eFRSWquaELlK
rEoOxoOAWf9Y4smYlJ+SYp9AdOfTtQAlk2rDpQH15UkMEGUa9sgoRY2BplOZIzK1nMAcDYNxfs8J
8n5QTU6d6kW9QrNQv01OOJwjndmJsmpdxU4wbHYHzScXNIRDV0MCnIJFeCNP3hWux+xPzQql3PKo
HG+2Kvz1ayzczzfWbgbWlnpoYK3JvhASchBITzHlYH5nlI7IaEXXGRRTF/NnqAFEp4aAjVc4Hw5C
YwwUhryikkDXrk5pB4JECzmIGY7LGLPruchFDC4uZf2FAA1+Nz1iK0qS8bMd81UdmeiByYaEdjnk
YeYFPi+gNGfCqGtzf2ElYQBz3npscLRGNB0+a+qwtjNtGu9d2aKXp+mC3jWooy8g8JHdujY0Nuhi
imwmE0fe3g0pxGhDt0Ak7FsmeXTz/8jFafT5DbYFRb+ZL4LmSrmnjJuKS1tDdcDc1G5sSy5Pt33a
mq+9T+JRs6rS4yNMyTB2nN6b5knrk/UYvp7QP7uEB5qI4IXxXDAx1MJZjhFzWMa3+bOAQRagwz6A
r4nfLSFVzcIJFY3mqfD5427zAtR3VwHq418js8awnUJUtEZ+Di5P2fM72/MNfJTS+2jZ97/y65yV
BzfBf9Eg59PJD63MQJ+x0SUdv/rDeo9++RJV2yV5r7FIsi5iZTnYzSF58HYcyKnwkn+pNM+k2jNf
8I/yDkS/FVn+VgciwKv+3JtZE4sXZGGebYhAPdE5ruJOhCZidXk+7eAiBy8BycjaIrrQgiQ2qXvF
pXWwNKHnZwBMYN+BBEzh6wWclQ4Usjjsm2jn0/1Zl38l6UAwz+h71WHXtlPYu3H0SuSmmqBXNlI2
8BVexV58k+20nb6FIn0zxzE=
`pragma protect end_protected

// 
