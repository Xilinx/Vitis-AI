`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
dxpBaoWYmFr4ZVs4jAlJMqCfYlNgYQOC7euOYQHWlgOXMAqRW8RhV6teROeriN3h4i8i+71w5aZx
8VECEnx5KjSytUWHnNpMTNpRlkPDFhgMe3Jz64cvpPwARDDChTk3G1MT2NZcOBmFpIVdr0IQVUxz
fpKu8jObVjWwKVjvvnM3Qf/pF/T3m8GvIhWzj85g0l0bRdAwyagl35UB2Fgws8H8UohJYvZ7AOkB
oSV8t2mKdYJIma+PIra2yUwZHnhgUaTQMxKEOQVHrOwk814SpxDzqxlj/jvR5CT0tzlYRo5K269a
V47uzyckKVEPA3g8lvqy9E3PccnJdlHT0HfgyQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="ca5u2V799fDZjOVzii9XcIKcDUahlwkBH5t7OWHjzkY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22064)
`pragma protect data_block
Oj97jVbqnpGdVTKlmdOV0kyrh5z4Jim5JhJC9Y5uh1hpNPyQGmdqAs/lyxKBGSFW3ATKDudg7NHA
WjvSa+gKOJ6Fd/mZQcQ4B+v4+JyZzx5V39ZSYQDCWEiDeINOCJYTfPhJPQBeOzrxI3ye7IA9vBS5
H2fzr2seNjgSynwJaffde1y7C9h+GfTRLGZhCNHruiAmdFWhX+jh5Ybl4R35uK/vzKuuZr+UnARI
nBJ+VT9rrfVTtnv6Z/atBuUOrnyXqzLBAxGGYaY60hwY/ffGQCarq0LNLXqwiWJ+oZC8tTy1Wdyd
DmCBoAE6DJIaubVGvB/eS9w+PBCAiuNCxV/YZB4FumvcSdOk1rRaOt84YcpJleYHRER+oTrmTVEW
tAN3xtXtNtPkmtCyHXE9R8Ig36RFIhrgRoph2DLi8cbhqWF+THcpZZIqkONYYEMmlzG+dqrAqzch
BThJxTk86Th7jjbZJwdIMFuRWbXuUlyQ7Le/qGXKdVlKsey/S1u9/Hdzyyp13ltJHJf4UgGizaC5
WGBhcV0duboanKwZGA4/kdcZ51Ajb3uC+P+LpfhILbM2SOHUV+T/BaGRVHCsc+BtlT7JWgCsX58b
q4U3Xia7CSMm8M0xAAjW/+phJSzwhP6obxo8DlPKwHz053eCC/eL3kSQY7UqOWu0C6hYLnmIyPDj
X89axYeUIlRbh0NojAkUMJMxAsJStmC4j2Swn4NWuslhYAdNUhrKJVwIhEIaqQ0gXKB0X/PCJ/7D
5JHxajmHk0NRG6oVoqLyzsZa11bdtvZ0GFp/6nZw7F3TJ652AVD9a3AlpmTApr0/WNLAuOPBCaOt
aTZ8kBB3CoIcvaJ9ZJSTqt1R8dceKcVqMbQfWBJse8vdafcm9TkOyDGxrpdxDsgjoLlqKgDWlXXM
bSEY/X1oZv0MP1SrZCvTNILZpGiJU8D57whrVlSJH7swqAbBcgz++l1OFWgj4U9QcJ7oaP8W4FOd
KWISupzpnuvwI2dKpZkF/RT4Qd3C9jGrOWL3kbtXyMkSim39We7OWLYtaiOqJkjKCl5qolkEFlmv
V7V7739Wq+mF6vXPLmyHadGnsfg+waDhirxqXoif2V/mwk/I0QQKPX7lBhgTwFv2r4UgtS/KYsdz
/cAHbBEWbLmFLQQfyhqphNnA3Gm0tScaoeTJ3nqMeJ0b68+WWb90o34p/OTD1t7Hi6+Cmh542suE
BCQByfPicYLcT6Lzj7JRTf8fWU8DA493AWMp5XbkFmyxMJDITdZ+RUWfGVgVL+SGPKYk5OIHrlWX
bXqdvRaf2a0Ftw1aZrWXnY7YrJonsJKedA95YWtAQ50WtUzaWs6txVRptaPhqkIW1Dkdy5UqXHdu
HVFLuG95LU9BcEdfzdoDoYWWhInHHBAr26xKqrWMEO5Oib0LRY0m7gS8x6M5rxAsRHplIazyovJh
MLaEFh81SjLxAkC/TLoMdc9CUipvfIOvseuB0bMYppEe208hOnJQNBE2UHA3dg0WCstVeRMg/G+e
xVcWcN7/eaQQhSOOpkqMbWuPBm5CRCXH+Zd+gPwG54/uYbfywxBeLh6FcNOabWClLfXqgQcKXvh8
zdTCgEkzLjRtYBYuS7p1vjVKdsGqwVCEkACoVerYleC/kVV4o9yN9iaNgZScef0c8lsUyS4TB78b
BI34yYn8LCvHge7WajZMgQ4UPlYKH5wUx1T64ONRSZX8yGE5SEDaucxYqVDRMe2MIWGAeHysvW8o
3HCC1S4Nv9fHEJIDgxIflP1mrfMQdq1Fy4U8P/Qk2mmGwBDn9H6l6rxShSCuF8OFH4K17PCCAvhD
h1eY7uD2xkX8hSEDcXyobQFTpkavfWkAxeGApmcjCPuxK5FFUN783ZETubslrmmt4ywsAdlFxhv1
ivRjJmG2SB8A/MCPYnQ2mwhxkGH2hcN3qR/Y7ErX92Mb4ISR8i+Yk0c9zEW8rJ9722Z1hBzGWiIW
Tk0Ug1s45rJEQpfC9bJ1vUFLQ4HCS/XNLONTq3f4ymj4CMhEPS7yIbKmbHrzWrDhwLwdMDNZJWDa
vAEzSkdMxLR3qiVbO1aZpyciaC7HzkUYgewQSZt3W9yhkyPPCY8RpRRFxH5GK7Jzp2sQmCYpcZjn
gDL8oDDJnooz1nSO4+nfIAQ9QnxMgj//1lUADIgpuQ9jGFirzYn3jN+woIXk31aDWOWNi13q9XVb
yl7vXlhWBwglRnQScH16YV9uEWiCRdkOmopPQRNci3VN4UkmiWM/2E4rq8oaisMqDPQSTcKOv14R
vyPryx9Xa8HOOmvr9AHL/5GFUMccon2vmd8MQLouE3skLTBlrAzCrlr28wFll7jxiSagJrYIzL98
zFd8dSGpa/xpX37xwsFsjOtyFXBZ6tB/juY3mk5GLzCCBV9IXZmsWwPuzsDbN1SYNWSHNJJTcORd
GBru2JNZYibz0CYkN4Sm9EyqKw8fUPn3qmu3uEpc7zUpDNcRnEj0l+org/6ha6dQKkbYcvsu5IHv
Z2uX2RmUSjIOzViF2oR5UE8mC45sbdI9MzgoqDg4lieJ4edpUOhGl3SkYC0omcQV64ep1tQfg0+C
7bJSJxwai4nkNl0xJEpUB0gQO6E/jr6hAiyz1KWHC/hIIZGLpAnw1THeTND/QaCUW7/WRLelFfph
0hBBdUEm/vwT9zH2Oc+KkhBuifjhelUVSCTGlteHknmCUw/s27lM2T5YMDad1G/LYzjgcpHBjzr/
M2tWmWW18kfUZzjLnEXuJPA8jWHOEzzSvT6HlVRAoLpsH/HTu3VjsAsYjw6gysWvu+sgbk1MsqFw
9soTr52DYvTnvrwH512qkKLEyIBPVxGqxL5KJAB0+K3fpNDSPDN3O2NsFDZ0NPLp2JkIDfWy8t9I
p6B5KPH38rJuv/B7ECIv4paA6r1YLmf7KBYAq41uMJrLLwp7Ou+wigLAm/Cs2rtLaFzew1BKN8nh
5sPbrN8X2NFiJ5aI3H4256abQh6xbaBdEaP1BdBa5YQwPixiAyW3rNQhgmNt5yyqWqFaD80Qc3ut
JC+M4gMFRV5G7LyoLYgqrjvf4XKHI9eo6AYP0w4PgVQXaSoL5He57JIG3KM5UtjmmreGw5j/i8Ce
sHIaSHdVJNJoY6N69NoqEPcYFWu6OCVB1rg3cgbSLHutS92g4Vqgx/FrMksvGaRX7Mplunb6lkh0
ZAdkAldcU4dprshhn03xXJ/ZWB74VzFZsO0wvCTINiAYdnyFn08a3JSBosuyXCIbPNU4bV1sPKS1
6sNpEm2rKYnqEjPhvQwZ0P8Gce/H82Gv6eFGXS4q5ODmOn6XTmH3BIIi1McO7O/kZ3MgJXkoNp3l
70ltCSbKrpLEd4qUFKmJGOX/FU2E2xcaHgQTNb4skgFCZpvZHNFfF9XpMpgv9VzaujliQxwLEfPT
a7IEfj2v7OClJ+gbdL+W7cQ7Psp2Ct5UhsYn6YNe6tEF9lFRI/WffNSmK3JqE+dXNfM4Ka26MMe0
+OOjW3uWvepbcJYn8thw4EeKpI8xgclpi0uocCfgB9bjMFxekZxUoFxWl9lyaCDBRMPCfD8OuiKH
9zkT2dGZ4vqQB3wOZBFqyYMiasn83ZtasF4UFd3SFhfYysNoN3CLoeoExiyPKN7OcO7hMNFD1di2
wSB0y4IwpBEZ10kx4ve6WW1kqhp1DPW7VuR1QQ0qpSb+ek2UtniESpqfgvJRKwVH/2kOohfXLRij
NlMdqrPXzRSn5dDuMr/9Ffa6HKOCbKR/izggo5JCxpcJ84JWPRsvdA7mpabi6uYmrHWRme4MMN15
WLAPG4Ajj7mVympc6svT8xJEuD5D0OqCLwAwcTwNOnnxA/NYTRbvDXUrEZN+W/sbKAoFH8KgMfP7
ejojMEoAM0EFn5JkNjypIbFOIJTvC/bK5KkWyLaZhLB4rhb5Be9IG1wqzluTPPvMLIqZxcm4ifa7
bsdtvPFpRvvNp2m4ZiuoMb2jr7/TgoRA1mUiqAMrnZ/6NRvMTTMDO5eBWrqEN5/bqMUDpSh5JVJG
WWA8/5kDf4DcWAtYTQLLvlGp8PxjwH3VnzjENpxLMjGaxn8/Kj6ndlNpBfkwrlkF1TwthdIp6BCc
JiLFtyO/R9+4iy/ySSGyf8n3lNC/lSGtNQwnfvcKsonAEe2dYqXD3MskW8vMb69FoG6QJ5BeJOLY
OcFmYsyQWfWIVYYr7fEHGpRzAyriXA62wshjXisNLvkfqINn/UMBZsOExqlCa2V/+nFWnGIQnMMQ
sThSIwjYS79kd+PYs6GCTbhQmIMjyQJPaz4POo1XaeUKP/hUq3gQyJO7qqf2NDYpQ8HKWVLo3rWJ
oWKmXTAxkYh6zcdpZlGmoTUPrgqTcTfXwILmbW2pw+ENyV5aAdqrdm+qZKFRwEfuUQKnNkUy6mm8
8Qhlp4sJ13zvm6klvlsBvRRLrw6ck0kZnFV2XEblM0qwiE3Ebo41Ij+N0SQqlchs8S93HEzIPpr4
ZFskHxZ6KTIzykXKTo7DyKWLD5momquWkoVaFUx734wOIae0jZyLumO9igQVMBDQSm/IjG+fIKeE
P7/W2j9wUjwJhlTLZ2C3J6ra6Bw/fXWKod4k9Be72e/I+GC/Dk7fzPC9j9o27HyHtcPkphsEjo8s
atmu5rPjmjPxbg8z3N/rFqhriGvc0gCgKq/H8YsPdb3W0qu6iXnWb7WROx6MTOeQBPOtuBIkv9pQ
cjDupWC6Sju49Rx82M7OyPaYH+g0RCT73LsAB7bMDnWf8DBQNmbL877EEvhUfs3VZ8en619jnZRd
nqp+Tfw8M2aa0kumKsSpM+Rpa9JicFIhxwFZ2Q49CEzW+1vl7Y6AEbmRyAZ/YQ1vgGH30nyjQ+Wj
dTIXWcfnrWRk4a1BdKTR/Mj2gsQpg8COgI8G7anTcNQ9AHc4reh5+qrK2+SlBS7v9vcDUclEirH7
0tFHX3aG/EkqePmp8e54O7NVV7On/9D3RZhM86h8rQ9b853VxWdsqZwt6BrLVvC52jy/cbC+y8sV
FfQb2OvA3dudukf+Omf74ojpycAQNk6+kr9uqCaWnvEKtY4q5dA3NnVdZe2XoxAHsQCfcRCj40a6
J2ad6cffhOVJ0spFpA32gJuP0JroQTZNLIhn7ONkibuE7AX9ab4+a8a2PWRK1Qi24T219G+ueV/I
kHzRSVZGSmHkXkQX2y15gUGGce/AcfGJQeuRPlFHT/jpp/Su0q9sKOGaefJGl74nq0D83Kk5Q0lo
jYqh5wQAIIx7Bq6Q1fXWLmgQcyMn6T0WTpdtnNbRpURf68EOpu2S/5NOxsGwZW/lOdNfvGXeAGh6
ebt9eto/IXtfQntM5FFgbLjPErdfHk5EMojCGSgoxDAnjGzAjftkNwR0J/B5dAbrnJvimZDU0DcJ
UNkQgzyewSSam+aO9JuLD/HwKszNKPo9AcVSWt+kH0c2MHKGYAdMjzLgtN6E5JA/KVmGN6KavPnX
15mQbnxBqArL7wjD4Aenl0tvnjdxf7ijE98EAHo6esNdP0iUWVnbFWTAwD1SNdntJyaKqL+HHDsJ
lWmjBOj2LrUUEZK044wnUvelAhs+n++CY+zdrS5Un7Z4Aj0hNCDgQDVHY8Yjq2HDQdfSuy+idCCu
OZKY9S+xmW2KRqv8bzif3sSfi83r3TLvV8NQWPaaLzRUmMsjm2msnnJVLPy7KBnIwvCYqjviIn5H
vbiTbqmVQZC+Bt/AuDX1q91uk+tPgQrnLtMw5puYRJTK3dHn98uF3aSB41j28e4b5/vnxWnYBawd
65QRj5OieggQ2mouiS6wzO9OsZaRmAeLN/y0FiUPVAkuKfEwbIdJowAJTV3pVUiiANKHgufFV9HK
nZazQccOJFvR3QgoImQP9YTMLiJ5/3odofNXVuUz+P7GIdKlPbRWlWl0TSWhaNXojd829aTUmiSq
ze9bK1HCVfY1jDE0yv5EY+6JmdfW6g0/uN+dgSiPfFIyeWgZpbjVmrHyh+9SB7kfPfHCBMuplvDu
345j48tyUqGOzFlGdyZ0bN1u2QxoMqfh56j9+15WOTnfUwhVVbcuU6cXyDTRIaoROjDAEMXdnKkJ
iYGqiCLz6yWOE1wZ0ueqYnQ8pciTPxB1QEBiVjcKIgNfh8JipH93TbYqw3mHjTQ1hlDvmPnqlps2
B+YIVHz7tW8I+bD4TFU4qtblTSh1ltia/ppbSeKbiKL0OgyXBVBD/Iuan5D5dds2KaM+U2ThxuQB
Br7nJ1n0Czhcfj+wvTQWD8rnaEB54txtClw1wq+FuDppRSMPYUyOQ5v9qzCQN/7O3WZf3sTaGYGv
sUuDJUxOJ0/Xh2dolXLZF06mQfoYmQvGFxXvWfQWr1CqIDftHA0HqAGjOYxnbIBbmwJvxNfmS6aH
GchckztjpJAQJQjI4+uL6P27uPMVcb/cIHoig6BbYa4rPMthGPXgd+9CQbuXhPfouTafWnU9XEeY
mk+C3rDoDGD50tCskAz+RIHy1vv5MHPTCkRiAj6sTgpiCV6iN3+a0QFfl82qHwf7M/xVNPFeembv
LEaRJ+HVPHyHECjP+Xshj768ZjXP+zTpWFVy237W7pAzLPY5r1vrTYCkZu3Zn6isRIc712nAHjIL
lrwjnh/npsSG8kSQs8eGTc509jlWT1IbXBynA2fCB7DU3R28UziD4q8rPKptj3/lbWYpjsFlQUiW
3EsLGdaBkhlSNz4fdfWBvm43y1dJ+SDs0azMpiSkzjOwojmuIxzHPc7BhLUfvAEdVC50fWcKwZHd
U4A1+QbFUD7UG1wKeUgGPjjoRB/Q2yfoyc/FN/BDmq0o9j+Dy7xXUfaeu7sEB2W1ovrcm4mfudy6
KFiHZn3bhmW1vkabhORUd4+E7AAxWulrvRNKI6H9ibmv8UKEWPeK4H2VaIE5REm+LucyFfx1R7PG
WuCNPd/7foedUn1l9t1/OBbmKZ0Bgi0vd1vk4C6yuZ37XBvAxgQBcS+WGZn1C/k1VX5ZUviYUBsg
r+qewvw+D+aXnUXOjxxfVV2T8FRww2dRGmTns2pnyGynBpTYV0DtpUts2rU8cNRcLJp2aBxfxxDa
DW2a9RDFgien2qi4ymq4tEtIRNsO3DD4S3UNQ+6B4t0GzXPNx4m8SLNvNvBKnadK2g6YL0Zgn8x4
2o1powXDnGEK1991mLpFEabYGbk2z1/ns3xFWumsD0A9CRpZ+xgNTpdNdnI3U9O5c4vwX2PngN7f
3L48jOp1mexbsJxh8HtzJi8mprTieEC2Alo5JAPXK3iVUYaiXYjA/U65P6A6h0Fe+MVOQYj/oQJM
0Y4oOyoml2XCSXp+rByqU/w3ADHLX4ULI6t4405X+jwmXc4HHSmegVFPWjquSPWEPyLKnS6Cp7Ux
vdOsRICW4nBwcTmIBBjTRk9FCibcHXREDgIZnyyQhl/NDbpQDukw+pQOdAQULOwxqhemgliKbtyQ
vGZhwa75STnpVVD6a1zSnn52mGyxTqRvOw+1/5dec+m5OqZAJz6XlRhESN3ZYStG7lhDQwkQ40C3
768Lmm2XI6BMZXcgDaO90oB8LRPz71jbfeavTAC+f7bD1PRIGuBWGL/sgZI60N3FWtf+Px8+UKIK
dmzRP8WPoWkibLoHV98IIYkhWKLtU8FfdBWOkXoIRvsW/V2yvs9G5uTtw5ByAx3j1+RVAS/wIuxg
4vd/2yTiIl70XWjxX+d0tvTnQoJyETLTY/V/1FM7Wi7r0Wq5ezfvn5Ro1w2PSf8pP4I6JkB5GayE
oaq84QwHf4p635H3u/Z/8oNyaROqVT/g+jwEvoPPUw7HEVha3YPUWJsdlgSMYFfg+3bQ+Qgf496U
oGB76hDBxt3XwxZlQY6u6xEw1FHyQ5R2siKu2Q93OY/3TAK3JZFaxfFZ6eLPrAanOAvS2EfkkE7M
MHRI1aZe5gvUhduETxrbWxfQzSNti3fzT75p9VYApomFAs4N2C+ymU5LpdDwzZYmP+sDxUAeIng6
8rroWA8FkWsI5/wJD5R4yPTcrxCDjADTRhINt5Z1vIhYBvyaCbX+hSKpw54lVBDGLPy7WVI9n6PU
lxOpB8xLnpunTPxFKT3irzsGfk8825hBWVBh/uF/CcX+ivEhyVpN3/yVreajY8zZA4Q0g+UjNYtN
PpoYiSs/ZEi0UqB6oX4A5cwT9aVynQVAK4IqOGbkXSZuO+aCkAw6cG3OapfkAM6YlfTCv5dTi/Vs
gJsplbAy/zrYh3fbswxdS/9JS2QrT1kD/9/RH6tcLPGaNEZLBG6R2HD2uxrZJhceNzsI3wgrGxv0
aJ2skZfZpprtFw6Cwx+2UDOqPYyUD5CbpOmR1wota+F4DsHh+vjBspyk47mWSfweedwWAnWfrXYj
l7VZ2T3AYWZ2oNpZD2ECzSsP8pAjW/RLV5RSA5/N03wLSsaAeWYD98rMXvUSpf3h6K8l7mIEF4+4
b/8BzV9lMVSBcBYz/3tk47giFpbZfbVnsa/vDDzYYhpy3vRDhbwyNterJ2HFIIZxc8+jlw8tH8Vy
vRTjGeiFLYe9gsYHUJ6y1Rk3CRXGBGVTPDJirRyzvWVh2iKg7eEzDUw7Gn9v+aBSU0y4MbLDLSgS
0H0d2r/CW/35z+1NPM4cqFqL8gnXZUi3N5RO7a05v/W+YTfKxxdO6uVjCiNTOOtSotqT6xgWl0k6
gKC7H6Xtx9HF13a11RicOt7YHCrUT3kMENnhNWzcTT1liTvwM2qDjSE6Wk/ozHVSmhzPji5gN8di
/E8kzZWsTkdaOWP0jsUmy+Az7BLugHJvJvNKb0IrShrv+eV8uWk4qDfOKd3uEXXvsN8OW7UWmq+K
b374xR/vhn0Tqe3QX4yZ2Kw1EppuduNovaHI4J68UAqG1VBAmMq1yWCpnk9qD9b/LJ10vnPd8GFm
pTpq/5cnBNsTnmu6EhP8RGUfsmP0k+rHHPaXQwAHo/+a2LHqNSi8m0eYZx6lSwu0grKHjf+mD1te
ZVp11HjLunXZOSdZJi6wjGDIz7MOK9vSGkTzrNRwyRkcfiGAlBRZgIdNsPsOpvNu9gswnVdswSGR
d3mJrA2ueQBqS24Q1OsAPWK4LuTvGhfywTRYTzWTxXanqBhu6CrPvWKm1YKQrcnyEXMt7DNkPCbn
OguTtzog2Fo5HUAQiIckN5cXwkQDyRzrVTBq5JQ3Sto9xNsSxGD33RaH5B1QgBHZ9k/+xSPrj1Fn
KYD85hLAmtHANEod6sXvLQwh1s+Duajpvh7hbNwJqYpVtn0WtDnCTrXS4qfVWXnDmWnLIlQDGE6m
4O5Uq6rtA/w4ZSnVuGXsPSm1v6izSXtF4w+U3b+mAmDJgg5j6IiP5+ViUrSW2F/seZxqsVQHp2c7
BS4IRB1yK60etYmVmt+LWnynpl+XEfTqL1a/opXjrfXMOGxzodViOEbunR0ujlz8yAEYI+BZrfzO
dT0JwmbL2ya58Z24OiOIlhpwDVTxHUvQlRHH6E3YM4uPA6RK/Ym14AWaaa08nGhIUVlylkx3N0I1
hzBM+i+iviG4rtZHmbzICqo8TvTaQN+aB3l8pLUfCHTs3Gumd4pxzIY61chGuJUDKk4MaAO0hq3H
AH4E4Wn++SSBsIsrVcJiwl9yvdOF3eU/BqubgbqiHji3i5OTZLbpa1xBU4iXlJxIA+IWBsrpx6V0
OyXntNmX/N87XcWSciEwmNvRx5LqUVEzAs3j2UM/IBhhOmRMuxx/NmiEmojE7ROWKvBWb2C45E9O
1Q2qqiAAIE7xxAI5QRYMgYWpLOHqVB76y1f5LSi7+mabA+9UeW1Op2qDV9lh/e/PddQ0tQg2WgWE
fqx+e1ZkD3aCSByv4nx3w4t8HBwyym/yTFZPTg/NAHh1tI8xPxfwD1LHCS3eQfyrgDdc5y7OVhF3
ePLTVmcwkGOxRB76unp81CQ1XU33z5IkELhZamQp43yTjGLD8BVZkZFpqyfoCArE6jAYwMBTlFdv
momGmnHgoA5sujkoHCbuKZX+XnENWo6FLWfBUNOXlZCm9LZ1JtloEVZbEtI5t4756qLYh35AX1w6
hlPubpfqYfKGuLKMTTgAna+9dD8zwHZYXM0FvzDEgT+2u1F1AJLloptK0fTtdxK3YjeE92cAJwna
UorHQ6HbE4sSHuNNYpLxwenggLAI4DMHwzcs0qRptLlxmtB9IrJkfY/QvA3fR5tvqGmBe5AUO7pm
Fv2Akd78hl0TvyOhhGvIPV66nVJhHkBV8ifo4R0pSEY4UZK6zMfcZTcWoH2wGGTGz+RjLEQVxm4w
DTvmp7fnumkjG8zEsH8jcbml3l0RermYtvD/4Llj6TcvqtkWltxiIB0J5m/RV4NZwzfFc7AOe9cL
E6+xH7L1hJAphnngPYZtg01lvGUnCcR0+/wNl8UdPCM+WPV0uZfc0t+k+3pLgafqaKBB4K4RtR57
KySk8jc1/uLmeN60qsyFSqgGAhyBrOum3UG12OEl5uWu9as84z4+YFCzrA2gfO9KWMS4dT61ClfQ
wadOsvygCET8c5/wP5iYMHvK6ycbPybr2qw51AXIGWN8JJ0HKI6+SOQLbLAl3/YWCK7Tj5ildCBY
neePhVjl4oUwrAn4Cqhs2Fp/zV80ckmzkFujd4W68aij8CrLuGa5r2PNaiBYBZYs8UNXD/OnOvCg
3MM3FNfx4QW2qaDw9i3/zArCnP3OiEOkt5ceoyTs3dFNF6Dy3DUG2Wd4OzL/6TPnwaKtLMnJIfLU
k2MUB0uk0sXOvk4DrxT3gSruW4lG0bToAMry5AphywHErZs9PdQWl+33xEYm6UCtPuq/CrMFtNI/
mJVW0+06xorTOG8WTdDCeJb2VcwV0dlYj+tnL95aIChQfgEdEToyDIgxOYRnndLYKCTd/fgqiHzr
M5NvTnaMaFbeZVzslMkawLcrbhnSg6UmWDf8BQddBIJZH+44mhC90HRFYvl/kqbVkd2Q2QbBSXwI
BqcI8zHJcIFoadz2RgM0+P+acmeVeMwN7osxxx/XZOBP5sI+/budd0x7HviHwkFOyyygvblC1mec
4rMu+CjWKdC2ZxyqUyI4n66uosSDv3cPlDp4fX59y8F+4Nxfv/2JiBn8Syq6MtENrVDjIm00DE96
ZmPbZSpM/af8znYHnjQ2WJKnRf0gPAlnTlx/VDtCZNmNRjGBLsF1NaPWD3DLCUeyEG8PzCQH8QgN
ExzU2H+Lh/dYbSpNosfm62nu7wBFaECpbR+iuzW0Jsfu1Qt0d1ZeurBps46O3j5juVSXVS7PPOrB
ycYFYcb4CksvQ+nuhI5Se1ztOGwdyx8s50So9r9ozwMeXyECcbTFYS97poxS1x9e/ng7qq+Pi+t5
u7/wi79mOPCSFfN+HXckPtKntfNVrq3tGgi7CNmSlxifw/uuk61dojzwCl67BFNTnVqsmhhaUhEw
ABsfPmP/q0UWS/ZTYGE+KdV30obBPzvllzC8br3YR0EdaeKV2B8+2irlBuxZVa+IUlhCHNF1x4zg
8UNo3/iTw25YvSEFWM4lZkkxTWY83OdtDuptnWze72mmOtCbfLuqhYOG6b4yUwGQt5DWE4fOGcY/
pnTwn5GIXQgjztJ9/+aP2ZqhfWYL6Di5CgzS8O8ZPPpTvYxLQ0Cj5MAUFcrIr/CxNsnv+PlyLqNi
hE787jiCQotgT7ZN0ZUTGnxYlr828/p5ulEj348GOv356hNTDLBcxRR30fryW//IxyVTiud/Hvnu
Er2EdYttC9FaaAIkwCQcnwlYK0VaX16lkaScaEcU/FKCYRKntq88Ms2eMXfHelk5EK0DjC/gNVXX
k7q1AC5kBhSRARN/Xa+sM529cTh3knLhVL04wrUAFwzuk3ddTWf7Bfp+iG+Ogu2OO7gyfMMqvjO9
8n3k1KXZKBMqAwoTqz9Y6UwAvfZXu5Nf8sejwCgm6mbjSmi6kpo16VD8IGWvbaARoS13Kq0Hi+xl
KVV4Ow1kGawnazFPAb+jwlKiyfRXFVviwK32OhDayMNJPyTuv+ciMABSE5qugjohOkdJVpK8QZbg
A38aPRnk4R1gxEIoKc0ps0OP115QK7DS23doumEHo1CPQIeYhJ9SwZo4XtQivlrisozXZk0Ia+aD
n5XUFb/za5hBc89+qLfJkWU+KlLHm/TUGuFBgLjKuNJoMS0uT5LnJsl5+bqyqC92MwJmKFaVdHdc
s/LJVHvaaehnQe6feAO/ot0zaqpqylF31xIt5aNaZhslG77AwiiX8Fm20nzhVFQU+XEXrVH0bJal
KSOZSE5CfDz3gOBLlqoNDNpL4tmMuTytFUH2VO/viVrEKZgSKK37veF/r8FFpZ66N+Bg/4Wsn99h
4Ds5V4Ux62RJjVXhr6vZm5MGQgR0FzjBWGgmgzm0jult6TXNt8PZNNiiRsH5tixk3DzCZwdG8Q+P
/iyoTV9YZNAu8WDDAMlvbiUeFBg9CAa/2y6Q9BjgWuSHHedovGpEziSv3i8lTk4aMrpU/+rLY+eg
Kuf7ixoDnEGrh8QRr95mKvByvGnmd1u/EZxF7dlHT6YxzEdDzpvPTfoaqM2GVcpTYHk68fYK3HGz
owe/xOX20bnRPcrmEmJ07IQJM9dNO61iYi8byzwkfPrVktqr+W10z6/DRw7B2CFLM3tUEafHOi3e
JtJahaBeMtzpyz2e4DciC0FA4PG2v5ETi3qPhQy7jroTjyx3bS7+T9Cm0MwejiEWJukWyIz8snfe
m9K0a/ddP9V4+D7OVlH0tYDkqtEN2oVQvSkglkROC0IX8m17ahWbuGrUdgLbi2VrgaBIFsx4+akf
GdP9PWlze26/GDRHQm4Uc23zKUcdpsDfO9mdPEw6FVul1YuzYIRoKKHf9DgDneBIAgikl3/Br+1U
L32sEyMbSY65wwE1wL7r/fr2Z01XItaJHDh9qTnfbWWAvOHb1AR53pf/9ZR6/HsI9cVtLN55+db+
7XH3WB1hI9ef3z7Qoa7ampZoBV0awX4jAZfHKYddxLdGeU2T+Wwx7l5cgl/ozgzgWlz5j+kVH1kg
Ja3vsgSMB4ee/o3fLEOjL/gUoMMW3n+/QMw38zWWeEfvAXf40HscAe9re5exq/Z/qwd5oLXeAyWg
8fcpFE0q+R2vCa+MrixqdqNfvLtCxCZ13SpytyLtrN1ivGZ6aqI7yN6RBVXU+dzY7m/EYkzcj2gt
WjDzOFUSF3zPRt3liFOCeoGnA+D7D+RvqsSdUolfMGsGP86CgXfGoRL02pRm/Uhr4/1ShL4RNV73
Fu+IpJY+efMDbx3K2CMtXr9NWjo1OcQO5AJ+6m09JdAu8CsZVhZiZFEWrn7yB0Nn/tLg3XC5grex
xIECWcn6sbPOUFX72T81K38uir8IZnX3ujXZC41R8d/CByYY/uDSkbmbIRFNDE5tiDb9kJ7csBwe
qGN4M+x9P3CRIS4zA+vvO6pBbq4K9qXuM6U5/mMmnCacEUfx0Fe/2O90wCyS3YxGopYN4cB/fpOf
ZxJJpBJE31uKFWM+N1/P8SBZrql5MhHf+o74yi/uc/jg0vAaKeuRw4/H3Kv+v1xmeck3QmXS/PcM
39yE80ya7ZpoIczIfi+17e126jdljtkH2W8YsrdxQjVieP2FTRui/sA4RAYQnVY2MtFJNTc+vvjv
bqTiSTBMYorTKpRfief/ffgIG+1rsrf6BqfGGrhQ3Oz7qiDh+DHySY07o02154HzNmAEBCIfnrcD
rkhkHyL0lZ1K+mspXk2h1FQRlhGonAyZ46eDJduBT+7C44jG3CZ3JvCKs+UrvnU6r1BZMG5wmwI0
snp+CbvlX8rUY1qCynPn+bUqYKSN0QFaRSnzAt4XdE9B1pt19pYAU3G+Ft6h85Yy9kc7WLG3drmw
BHCEhrEKHalpxyqtLdvx7EXxgpHJiBe5isC2e+puEooA43yKd1mJhmb3vAj/zpXMycPEg8Ej/cvl
7pOch7y2xlMJG9EmnsVXfUHkQGl0jtsrfrrZwGtRVev322+EB6UhCVkKbEoeRQqaTaOHuk4AFgNF
vo3qGbtSl5pPh+UajYRdRvmuXRK+q2tRnLGXlt39zYUb217xbJtORcSVJEyIUDjMZFcJO4SSjGrs
g4q0IBqOVCRyCC7dR9ONZaOpqqsEDsOjcbtJITaghheb64lAtjmfl6FYjhgMMch3MuQJTzXzMk5J
/21r8GJ+EepKX5ZAe76VxLxWVgs2lmSfelq9O1tAFalNvlQVRU6GYrs4cdPGkYlAtn+COf530sVf
hIkQw+Fhkq7YYtBIiy4kcrn3xG6N5y40cRQxVGHQuoLOvWesd0oMXT+zNIiaEbnX9CXv2VCvyXHj
woF9Wwb88aFCFJygQ9Rpq59GBNUYTkJtn2RSj0svR6JqcMhPgCMLmlA2Xt4oNkiOcB9l8qfCpJ6+
yWy+Fv7YG/lKt8Flzb+Dj/3kRAnyKM7z/ULokC5IMsgflPvT1k70Jf81ybVHu8EnoKSsdpw9PJyh
FcCrKOiFE/9QbhrjMeL7EbX4ojB4bwGBwi6IgRwuDv+Z7AZlly522ySbZNWJTY1JXQipuMsNbz59
TZ6Z1TNmoQ5cG1tfJKSJt2PTAkLgbTQ/+d+mP7V3jlxkJADYgXqY/WLj6OFGr2mml1qDk1/feEHg
SCZ08+FaRT90gHUfZhS+WoJii4UhJDfSXnBvrpY/xHccgVT+0fw9FXQoJNCwKP1XCguFdDXWifIv
WtZ9KvdIFk3JaYfKaVnOEa3OXe5wLJgTwptfKbVF9Ccbdn2L6vV7Y3okDpUARuGiKAZ2Or14+W+e
lemih4JJQKhKgrg+ElTg/xedgh5FAZzm5pk3kLWRjYrr41igX8edJdXKJwOVkcFrbbsk6ffLz7c4
lQqxZ9Bve2Pg6oBtmFuosRfi5rR4AbdfVfWLk6zWkUkaLTcYlrERVC+0voxmrjGlU258NC3KCVof
e1htRY3PZJcGKNz2eeIX4GgqXkOajjDUOFKx+Y+y3P1F1OIXkutBdzIHk1EPE7VEztmfn0EO12Dq
DoSx8skW3piXernDHd+ZjxMz+SJqJ3ql3DZyF7cgzco1IBlPT+Rom20r0eVTxfWsHWGNBVoPx86u
8Q0vJdHfxCPt2jU+J9hdRyaA8s7LN28asEiFNEvQIuH/m1vaRigVEG9nD3l2kNg3sUn2ofWZZD0F
Ez0MgjJRc5XBYlVWpVaybRdVvFrBZFriz1obwM0Gwd/ChPX457jA/GH/j7bxHsGv8ThG48fiYvrt
1cYeyOj12D1CJejm1UtTV5p57yPnqPiHLTqWu/qpysfwFRVpqokV2RiLGC825iGZvDxuvytnDKWp
gQ0Z48u8nDxzBEGdHfePx9s3yYeJvyjER5NHJ+hGol3wO45DLho7bn6G2s43Ot/9NvyLcIyUS23L
q+uvFsNtlz03Jv7sqpgDPGso0otWtjlSP31IUXq3QsGY56H02USllbZ7Vrm5O5GoeOz7Tyo/Ielc
kvs4aH0HoUw2XJCd1OgiEXAZbBp8HBDsB1GR4p86sR2+Y6foP83pUBO0LU3FiIewIAgrJIpBy/jI
gEA8DpThkDWCAO3x95pm/T9WHW9GV1iM/CSCUAGwPgWN9vwK2LVEcbySxhyQ221NE4Li4Jr7w29B
KPwkFjodyBESL8T6g2FbErJWn4XEtTZiurgdhsP2xwikcKTrYdv7Q2kkI4HmxOBY48o5i+2VpOQY
990NHkhqPAdvCVOnTwy7oGo2O6MHOxe5Sg208i48Rvk7K+/3+kSASMj0juu7PS8kv+K3l9aPybXY
XVCvPZ6gvgmJSqO0lep7JLxHdpapdfW2O7DG0Obfa+K5WdFHAG8BG3+zw5qpkReI+j7ZIhqiZ1Za
nH8QtlAJ4rB+NYkBbGdaIKYiuYMrRv82uvkMIElAMNOgIevtJVtw87FolL64uaMGqEbVINqz657y
YKoU8h7M6ZzlBTjOToFlkUxIz+khR9Qjcr9pbpgG7s1wx3mA6kg9nPfFg1QBpq1aAzUsjXBkYdj/
iaNP8WqM/hsZK3LT2ctdtN2w5zLbo6WyF+RCRJu6QWSWUWKSn03g6jSyeYK/+xHCaohMifqpC5oa
ilqTegaWhcV7S6Sk3tlqhmYS0ON0tLOB2otUuBzIJFWwuwbWbY377CtJIkivN/3DBaSJO5zK6ssv
E/cjWeyhlPaB0PH8Sp67qiHabtxaLsm8u0aj7YEnKDzswSoNfFAJzAj3l/8NgQpIWlo4VpjRckUB
BznTbi0hu6A7HacA1erEw+zAdzs8iZujVDdfHMhQYn2FjBGA/7UORvWFd08OT/ZUpsKvgAUzGZ37
ushFllR71sh4eMI73Mn6MexRgQizgxezhwwL11NKoMZBAqdC03J56X8f4Cxu/iEbQhmu9H5/o5kY
8CZVypRd1l26FFLEW4Mh3GH0Yk5IN1TORvgIf0DWiCEgHtTx2jA/gz/AHBdF3HvntWjKknDkdVoU
VigM7jHmL4rEHAbjJTmdc5dxzAqIoznwfOCTe+7jdfSArHpgfwyF8n7mjTFvOkvbDduG+N4pDuKb
FKth6J8cMTmcMdeDFK7n2/0K3Cv1bPt1xvkv2sec91rOIwzfYffzqPFwbQrGrr7oQf+22HEhlIAm
GHxhQoZrcQuhSXArQkSaHXKsu6mgZuczlzHiwPH17T51sl53m563WuybUcVz/EbYLilOeedwkXU2
zSNO8vBm+Z20arRrIzh88dqN9fmpjsV/U+x91n+zHx1GwgVE44N5vp8QC2n92YovECyaUA73XgzZ
UW5hr/kwKkANwk6RBYiLYts7Z3ukR0XdHIol36wMTXL0yF2Lv21yzsCFSQDDRDP77MCREUgU4hTD
XkyQ1FxOEuDRC0/0a3O1W5tA1wB5KRl3Bh4ANnUA/ggkxtxP14iEX5oY7Hi9IfP7onaVd602p0dq
wp8JOhvY/utu+la2bpiaQl3iSXNBwrCDZRcLkpHNOFcfpy0rR0DksuIXrzJA6iw/5B/32jmC89rW
PyVPxKtxBNdbCp79NiKqoQm7H8sdo5Aq3Hd0BdsC99xzBVohzEp5nhirGnI72ZS4by4OcR5I0D3v
wz6aQnFve+WKKF6oqTob6/d3HX+xctdAp45FsB/wmjSv12Q/QasAW8l4Rjpqi/Dr87mr5KOpimUj
n5GVi5O7JKlBEGVXGbcIskSpxAS54T1xI+/KodJv0i2dgBt3QeqJH2c2GPLU3M3EYi55to8/6hfx
1hfw1B6PHDaZJXjPo7nhDqSN8ctZqYVDUTNYmsvv/OqVtSOeEPSdRs2kdpCnurrtm/awyyC0HP0W
I29XXoFFI4bbE3Uehbu0CB30eEiDmHp6+yXUyLEtEtMNMElodHgS8h+AeGkyTmhw9Efr5Tqd1V6H
LdHa0xVbVVtaOr8JN6PJKOL6XodMeyoVG8qCq7ZCWq/yOTpKrw0sUYK8qsaarXXdoz1KaJk0wpvo
H2BjmK1q17GV4xFEAYZcO6RdsUAE3ulx94Vvx6L3C1Uhstof1xXwCaub3BD0jGpEQJMWLZ8K8Her
prtuVowQY86EyiHjS9hsPIIk3twf9ctGsG0UFDisZVXhLdtYoEHtakwrgjcbyG4bh0rp85QB4NON
P8aPoiK8G/9Kh86bShxvpeu7ED385uue1amjfxz8xOk6PnddG46c4mDH7zXgkHZG7IYn7L1qeMTB
TU2tAijUOZQpsuzpY2r2eX9tlTTc1ctTtGi8u1kEkufZCUCRqwsBw+mRrxSHsxsk4WAWWnPTepTb
PxPy/Ky4bqLXePjM1AyFKT7BjLKDQvUHuA04AQKKsQM25pzTmRs6v6QWV1oggJgFgb5cQOMU+3Ig
HwuLOR+97TRVHcvdbzow5WSLPUQac/BMHlBcxQXvhDT4ahAlS1ilrDY6NAFRbZJoMazLNXeI/HtL
5L5nFTGcXv1VzAufLVDsT+XyxFyHRlFqjyrmRWICm+NivG+OfRkZM7y9b593QtV1PI0SDzl5aeW7
xc5S1keWeZc2e3JlmkDV21u+XzWIVLFm5ooyfufw5g5osUk2SA4q2xnk0rFnIbTMld/VgGTUrI8b
Gf4KV6ODWbVsNUS/pWGAWAp3nTZmeCouHgxD+XW26gBjSlU4mj1uyVblWkP50gTzkL8jnmNWTvFn
DvzGgTdso8NsgZcp+4HEbW207xiB7zyJWwqsyLVav4M6MzqooWvQ8bOc7dHlIW0Am731AETGQzmb
ZtfIBjmb/0SOrRzSsB2B1DG90x0TCuX6uPreft+VZqz9Fq+/MoDThaOsAfCNwqJ4uXCvqvJRii2q
JTEcYOFnsHWEpL2ySx5/LUFxA6dyt/aUt7h0hsjInMRyRf8duV/+DavLS+SQf5Ft6bKNpCUVU9KE
oBoSW3H+/KhJGIkYbY+xse+swIS3dPJsS2r6uJS6Kk32r0aIPjs6O7oYXQh8t+4GiBRTtDvhMJL3
lKd02cwxEOK4Oor+XbZza3mgeNxFxL/1FyYFTXoSzJz65/S8vTQBFbuImxD8U6tALa5wujk13d+f
CoC+abArx4Qs7OctMckN6CxXzRcBfClJkBBVo96HOcVR2/5ZrUnUFkm//GNzJnnHvarK63ME4I+L
iG9kLiw2utbwCqxlfWd9HaiRyngsyC6ZPkHkdhZ/xYdiru1chuHpNv4uX7MTW3CgzyGo9gEVFO2t
Zsy2ZoSpTmCbZYZErw/IgK3WFCml4+Jl2jBV5AocYHeOCQIwRzoQu5GIiUhhnL/cw4FzALxFc0Zf
bLscoiwaQ+UyykcuYY3ASiEyUtN+n1c64CPw0ZNMeEFrJvYbEeOUfBw80big1TL5CjiyxBqDQzt2
Yxq26t9pCDj3J87nrh3aFv/8GDAlRKxCzG9mdGzNq4N0WHpSBgnUJKTF8egd6ZO6Xc8s4/mTw76B
d6Xu3YfciKtlHiHFOWhZrZkEY7kXCncONHQYa1he1J+kakh7N38kiomz5jo1j1TTgKD0GndSvdKr
TTwCmJZohO17AjiPJRSvG3kNHEVK6bojteeTCRlRwFDhFv3HtP4+a/x/799BiJdk1kggN90euSjn
bZpa3iXIRlmz29cOViwMEe6bSE5O6xp4eQi4NqMq5iqJOlw+2ONZfMuwxaM4EWUwJmPc0zQxX6qG
OThLni66LyuYWIEZeVOdL7LMHY42LFHrS7z+mNFlRKqbsHAoJHlW8j8NxZ+VijYKu60jozlu3VQr
1/JC7IzEiOSiIfbksssj0V6LWn3pnnOxyVm+4SiqxxaQpvF4tV+M8vXGqd6fzkRFFcSRJdlB/ZUj
7zS91X0tf0He0TQVksxBEXNb+hJxwHRBc2gxT56C6rClBLk9Pgrl/+859CdCS1bl6JxXQOOPmg7a
8Aj6G1ZglaNWXCbIHEpBCFzodkvWAlKTpcHnhic0zAMyr+7IXZBIwSMHFEswbnj5M8GWMQ9fE7my
pz6XEvG9PFFoGRZci3SBv2JYszDSGU3Q9gk1Haul1h/VkP/rNsZBYScKAPaiHe8+32qbDB4EggbN
ESZ7kn5CY3tifwukP1FILleS7K1YjAtUcxKqsiLsc9R2N0fxhOmDlCe44WnPRpaw/cOYi38NeBYG
yg9zDAEuFFtkauSTLuQls4uanuE7nuXR+gAHlcAShiLkiZHwCGsZQLWXUG0tEJZlyj5ibcA0HI1G
TIxAMt68gHGOnTgGIaUj3pIi1Vd61/LUm0+24CaGVrPibVXSrHWRwDnPmHHdw78Wso8Iwp1eRgJy
zJDtixCSnuxt7KBNKbkQ+KfMt/i/4P7NKqd1rJ/aWeosgj6qyba6Xd+HepmaUwqwhBIE7sH2PPE6
QA90+Sv4vbjLgGJMS9twqlLV9tWfoHRgSygF6TSsCWBzE8c12H2+VMJJv0Sm6lveZnaKJcipB+z3
4uLQO81lHMIlX9LKfWriNGi5MEzUkimHFsT593pMh0a1/P7H5YQveH8tJnZwJSclkCNM7//cbmyq
1DyJmHibgF0kv1LPj+bxQLVYnE4zDlpYBiCUhIHguDM7VC3vBEojU4I3TF3T4azLY8gu/MYBqmO5
JZD387K3Y0IRMDf8FA2d/Ym00PvvfEdlTsMg90OlXP3DlorRwx6JnF0Bl495YUp8Woxvq8Xal2Y6
L8TDI5JkCRk23Y5GQQVfZyQ9XkeEqe+vky+kK+ojDlp5m7Z4XLpXF/iZMOWevcBsj6559eaX5//E
payNtLgHjOFGt40vT3oI4Vlne42SUMUglr1T35nm1QmR4v8e747T82y0Nv7XjZpMffDzYW+KByoG
f1Sa1TmR0NcwH8EeM0BSWqGY4M/CA+xQmFrWtWLD11X17OVmkHUO1OXJCDjrX4wZtxdned9RNfDh
uVBfy+YudnphMr/URXbuXKTblVtfClV9TJjhgq75+nDUh4yhU5JKkHZ77k3LIRcIVAg1LXWCX8OQ
ji1KGTwfLmhqksO64yZ0BbpatKSSSgAWS8C15EMo23ra1FReNS17eZ+l99J7B9EHQhhyLqN4IWYW
qB/1iL1F9xcD7K7ZbC+kWwO4bGEO+V0s0Ozzm9lLFQpoC7BLuoVCEZoL3N8gPGx4JoGPLdY1F5af
hwUQyfs1oW62S7D2YM2guhLsb1Fiz1hHsTdmYGZ7Df049CrEZwq6xGxexRCeGywrkEZFW3CMMLPG
svvotYd6kjKS78VnWa3KYXbeinOMJI+lqPmr2LbawVjRz/7P5Wq20BVNHO9UIoOBpM2Fmqh9xALZ
oGgFdS0+9DmC7EdJ0o/k3iZBVmzKDKrF4nLmtUT+NEJ+EundJOyMKftmNlTj6BmSXvYpDVPeaZLi
J4nsCQ1kCVBH4SpAtMFUzdku8AwI1WqjUwsZ9w9gc7K9ukpzMC4zF1P7Nprji96IQUbiU6QwyX4n
CkaU6F5FOoiZCL9RHoEy+lGoETJX8LwE1ybZXTuQ1o54qEuIhu86if/D7xsw4jUu5f+rexTvRNUt
pUyQ+l2YXPfK1M1mZ/VlbUUWLSoHz6KYz07gzP0NApM+KcMLW6ABg/ViLc20JxjTRthK9okWht59
WroEL9kMWVNRNHQTyRfxzwhGuzwZzI2UnucgFREWNqapoDCcSYbYQeznINvUWUUjcIHO1CA6GQRv
WRR0J1lomk5a2dY3AajpjAxtBTSi0rzVV7T7pcgc+57zU1nsw+8lOdroeZ/wyUyU21EQwS9ZzoHx
g2EicBi27KOYOGeaZQSoh5Tb8JJuwvilP/KWQPdeobXOmaBWOnSFophWEdcUOZ6YnKv4YHZ25F/q
4jESW0/crnVkh0sRvgOq9vXop4WpcyHJNP+941JUw2bB9xUW76QGuYgc69RM1f7HGHqnKBkrPNGz
eXCVR/AuUY9KCHqn2JyxuCy7NoZKSSy9SrS61i/8vb6EyT3OYim2pPOZjxuYiUtIcZmIlrHFIMdJ
SYx9MzkKwDrjxS7hPkg8QtSYAwE0NwAMUrfhVUfSBqLxHxqxKKTI3CExqmmWhy3JVu6V93vNvgQe
e36qvYDVgM/GPI6W4Rq2a8ILAkb4RzXniiHl99cQe+srAowuHnJRG3vTyY93M8HPK13h/CjfzdbG
nwD4juV/dZix+xjS8W3AZFaLH7vGcTgGkUP9ZTY1pdkdx/DiDfOS/KIrVOFKF2ZgKSgnUPjzWbNa
bPHd+Az0hCvMxAiqH08pEM1CAJcrIWnOSLS2NOM5scVSJAEZbZZg+CuaVjFdFjrq3wIs2ay0PbCZ
I+1l6R9yXc2KYo5r/PlOCYPsz/EFKFheTQrC1ZvZ/ZxuDHegS2bvR27TY74hIHcrrvIveSUzFgYT
CHjquGRVLDR6VrIvJ5LMpKP/RNcG6bWYs7qVRy9faFPOwUh/cNpW7uAL+Kj+ELxjo9y5SLD8GNIi
VfJngLSXzSHmumi0JiBFzCUzBL2fIKx4nNv6/Xp6dT7h4UBtwGkSA4NXwPULoE4H76k4qjxLjjwH
9nn2U8ECo+5lzNMh08aVxlu8jieUklxZWHu97qRz86AMvjOTa3qXmmhtZffN1M1veOh8jCzQPoV/
ceWzs3797TyJSulmlMxrXlWUcdhsIueaZN2GLnNK9KRwcWxdFE6rq0Kba1hDVlFWJhZOiVjM+7NM
jyWNH4Kxtz+qrDqleux5bqUhwBZeKUnzHt066B+e97YCTtrYJlXldiNZPETzvx3/0gmZTDUvlKao
nLRqApIYgYpowk/8PAt4SeDPT2hrRw7kiTHSQDCBAElOa7dDHiC+CI8qtkf9sY7aP6OGVBCDltBf
N5LD1tAAwPakULdbGq1OhVdQvDh/FLOPTvGlaRiK5FMpHyt6s4om1Fmcrs86R362rwRfitOHRIHk
p4dBSYggHbWqANOsj3MOKjjPAV6YTkCtR9WZj0EbyBnK/3KiCXT2AVKZxY7QsQTUx/QZa0aEl5Ln
x435LQgdlcAUwa5d1Wckawhz6GznDXmlDVrdm+JBOfAfzO7GJiAl8wrySFzZWVpCcjh26H7AZEnM
0D+KXO6FuHctMKQD82TxJL6LjWPAanRsS+2wx16w3tnkn2Zig/Hn/6HFvXlvrl33sw477GahOO3U
rx0xlpbrIM+RBXJbM8ZzT5gf+HWAqtXIChieL+3qDXfkjK2Dy1mKLvBPuqT1mvECFsll3SneeSkG
4Ij4yXCtoHN/+8t9TT6PEMzAV3HhlN/BrJl+Zh9Dvg4w7immh3dSZzID/OZjCFyRSTTUz4A8ZGDL
KsRgUnylKKgZIA9BBOvTmkrvN3fDU/gsE8sVhBzDNqy1i7gSHb7rQsyCrJKfq9QVlu4FAZP0dxx5
JLEzd9XWvzJiNoxmFWKvkt7hbjrv49ZaAL4fQEbZ3+FRcAOUQbRO08FULxdlirlNzh3vWJJXtf5G
pw3N1nV8H/c3tqoyCxv8AMXLZQh3KcwraHvUi+qh9sDf6jVrCuwn0k7yTaJfZo4kI2YD86ja4fAV
tBSIqwwUur+9sqjr+bdp1Wz55Oldl/F7C1w0kFC7JX/kWSTC8rBwbKdjmwKBIGoRTQG1xALAr56W
2fR0n2vM6JWD8uyvxmyW1do68lHiVE2EfYWF+u6lfTYVuL3aMF/chXoFKcW4sBEu9zTeOdhsBFNG
V09CwB/Wek5sVy6ieA5/dfR+BctEVzNtj5jyKtEVwpbOYNWPTnGkNKwOvBTDpkABFYnfz3PO1dW9
i2+1dhLJZOPknnyxqaUqBdL7Jor5WZTwjJh0CYVP8hIdJCrlFH9MGmIxWOlcwYt9fwqs+89r7+1C
9m29BDIlcxbrv+hhCBkpWobusTmEnhZpS43df1Y/qpz3Os2y3QtaNIIEqbmLyNbDONObeTi+cxfJ
0bsHiIewgx9qxRFXS2HOPI6bK95htYggfiHzTF6GSSiU3amv34RstP3N8FVUXqNJ0fwPgOhd8iaq
F1CU1csyMOWeQGtdrzn7SvpboOOzMuUS5JjV0zj0cSZtcbmxFxOwzIYKnaXpSsWwPayaxKelX4Ym
/BFcf+tImD8l0QZLKAQUH4EwN3DovnFWLtuESVwYf3vCyEjzGjRmvA+YUCLAN7sCI2Cov6PehAK5
FFHlcootRIX0PDPuf8mIyL0ZLRBBtMUcLa+1bHWjr6jSup0FFnzHub+GfRTvUGRlJTzO6ksiYhr0
49LLpU03/91cEdfGpLumaItQJL1pGaUHTryODfNVVOl4r5VYDuw9gKb+VnB8yYaaUJrLNOs0eWcs
ZwEhaUHGdOtJeepv1fa5EQW36oqIiLarjObXsIMCkBJqVJfya1JMefXqGfZOb+UGDAPnNKQmAbNR
u/Wf0sDMy0nH+ilnVhvt7NSFh9RJrrbXUVA64Bho1gcLHVhpnxzyyhZq+sdaoWCPFRq1tCkPL5wx
LZ8KFimsNLAEVXmdA5isrsyC2sjcT3o2TgStC2vUX0I1XMZ7lv14LUnEuV75uuWpsrdW2zsQoRWV
NFXcPSgef+TXGJtRvxIVCSmlEQ2MBxyr3vpHbuBOi6RqNA9BTWMGWg2EY1fpaXOFub+3Nbtz05lB
ENZW/iZxClFarAqfGGuF/9rGq2IP0++wJkhgqhxIdxZT54BfQO9KCmIsOoT9rnBBzfCQB9bIVC7a
NZQm07JPZy6ONyFI2XJHSpfTy0zgjmeUmjiSITz4tck1ThUAx6YwjKOih3427k4xDjU9DrfDIbbI
Kpc4L8MZVmD4bpt8qa2qNkN6o2F7pZQM3LN+DwqZCr3Lr4qt+0se31SwK19aegzDHu6tVDvfz2gO
Ks7TrCkK6zqEhTKClUKlFlNkLPPt/MIMOswMgOm2XnxaQZFmQ93nbFFAE2EwuWf/LfcuVfHo8TOc
nsqUtFww7p2rObzSbLdNe/n14cEcZfoWJ+BLKgSahbMWfWd482NCpDBC/Soo65c5uys7qN/LTH2s
hibcl1O/G0KsQtDr4eyQFUTW5VYGDBKtD/QHoJedH6rFIkv9S7FXETBBIqoRgcE1nkQ6iXCRlPtt
PNEM4aJfhtxaV7c/3zlgjYmw2lH3akmIJVQTotBCYPx7Ssca2S/IXmQiGJmK8aXQjDmyd3X5McIl
J8Qs6M/EMmxL3f8YYVW5t88NTicROhmkcvqf4SzPEtQ/JIyhc8VHOsN3jLvUtK/7+2Evwy+Ikhjp
RySbOuu2uQyxHwiZHdLHjR2DMZnR6yZn4iqEnLc7BmBNE72DRvYnkt7vhDwDpGDEPsVYgsvlMn9K
DV7q4ILL4beV3jVumxHg5H8uLEX4XTKHooCiNKP2jnjtawJAqriAqJa9lXLWja1jB5EOmmiTrOPm
ACG47QynrtVm1XmTaV6bSOE86s1xrwDdemBJ3EMyQUzNoX18YacpD2I+Arxai/WJA23QXMElFJrb
wSW5B9+x4pCx2mQQq289UTgrvjW5ncLgE2tPAmrQKRpRwbs1Rs0sqAYdUfxXxzE8CAUb+F9hlIpO
qBiKXEGuTmBSp6zTrZqZP52EYPWd4gZhb64kG+y027W09qErjwqlG0BlVUuUKC35NjfJOr9LAG+o
0r7Cb/HezR66F+tYVxWOVp0dvprVYcuCvzYJ6rwTawHD6QDTADhh+vgtX31cVRXedynqmwFwVJdq
peYo28oto0qwKJSqr5uP98CPS75xKZ1oVcOyXYs1r/d+/IjfyxJBrHeiFlHBsl5qbnAWhuGaAf5p
Ql++4fSZG3Z24j6tQdNOsqMJS+u6U1ZdWuLT87uvIJAMhxH3jvRxbd7nItHZFckOIXJq6W72pa7h
BzsrRG1KuvVALqLF2xbUiwE4rGHAdjeNzIxqMmZ4esJh6MGXQQxtKxssgmJKO+riZ4kEoFF13HvN
vG6oDnkGg60N34LproHOmHhuz1vhnjYMRsjWyKrFHS+9rjSui5kkNEXplLi609BiREq87AeTPd4T
rHgLm+k2ixuwaP/hUF9khsjAjMbKKiryeWyKZceT7CJcAzO38keFCxkRgGjhUJDxE7uwWC82vZkI
qyX0pgqNrXWLhvvshR/Jt8/Gb49vAV0iNsaeQLtTys0V73V9d4/00TnL9KRKRb8EvttCcvTgCbUU
dbuAL842n0oS6lbdU2CXFNBUViWVnkJ6gbGwevWomBtR09Qf7dwDXuvTj5v2hJ3Gj8VQqGKOzAps
M4vnFeLtj5KpX0JgNlBehL3ny1cHCcdCZeqcfJmbEZA2+IX29Cwky5nhZx9nnEcKfsniXgdun/98
hVtEo0U4IhvfeDCpm6ZY+dHdH/H+zqMI9uR1RxltOnBrn0icMXJHMV2UEAABmcu4OSog6Odr8X+y
PPjBpw1V3KUAd7VTLE5m9Wkc9A5rtvGWRiNJrTwNyXv3lUeITZk+4UpZ08M1mHceJ0Lz0ObX+/4I
SCn/rrQJLLKjXFa5WPuyZBzzqpKzJXcrBNNlT83Nq/uSB4cV3w+DXI6tULITA5CGCK+cQpIddy8f
meV4KANYtIR+2PGLdfFNQfrnCmXbcMlNHIjMWX7+C1kVJLf0YjSAB6M4KgVf8DtegHAylLbqjt/Z
bpJm4iO7tAaOZl/tQXFhjh02X7v7nIz6Ky8w/pisQWoJ/dQb5Rf/pZ1FkO/PcxjZTldkjXeQi3IS
nRuTNmNFCYTmFMg+GIgMZIf7I8jBL9ua2h8ohNqpbUvGSnIaHWrvwK7vdkp/zHu6/kF+YUHcENB5
gYKOLNlY5LEsjYTetX+SpnyhuFeXznKr8Lu0n3437ReO82zq4gmz0rkAbnFMlfiYpa4aR99UVfBk
5yHl4OZqHwN6e4ETy/GrbodIaMwRzZXvDM+YQmhS5A03gMaXmVj2+lvH2YyAnA0CXOTLi9VDt61F
nF9D0Whg/eOBDD/vKjyGSrZP4aeg3HrMTlz5GAxS5TctTUia6r9tcdMnKvzs78Gf/Hcqt4RIq6Ch
ZkgTHokDSr3ojKFjg3mfC4526MWoKuhsWw5snABqeI+3LExOMzhAloxHqfTbIwD/HLYMo62eb/eo
BzDnEz8fMS0OzUevKe6GcdrB6vJPsy4TqpcDYn+YKZ6t+zcLc4mirx7+ikPV2HOm5ICTdn6/gb/c
tEmy9KHRk//jFT2ZSdS13TIyaodmZ2bDN3y1dlDrzexHrqNwEqKB3V/gKr9adD4RFuIyPc6GwXNR
Ggum+SOeZGfQ8nyonbZh2XoYiT4aRjpV3WAbU6tZZQVcRR7OwG4fdDtwfO9ZBFpALieucqM6WGS9
ziTj7PMDhP+kKRItYiL2TBHaixVmc+27RFYkqr+xmlIMIL4GX+MpMvpo//t+16dktHQO4K3pcRZg
pkJ51zkCFK+CtOxnA66taaQnTsIQmHCa0/Q2QoYc8r1t28OZW8qSonnqlgbK5SFKFnRsYKhCIPya
9GpgCH6sJKgtVBufIg9VQ3Y67A165bN0RZ86Tol2LXM6v62wvp3gxpPf9AI65/jNVkLqx0g4EBOm
y6lbWqJWH4RgPzoAiF7OmoUFZvr6SQIHOIo8PBbvAkzb7m+isGf+BW78e5G9NCJk273dICoIBtsr
ZK+UHwSMkmd1i7/JEVXI1V/hJvcNnWxGT9vVw1XHp4EvxV2xVPcqrmBtn2zm7BFJcJPgIs55P4zx
+I+Rj34A+0Oeytrytb/XJkFgOyWZQZqFWoXRf8bZsiOcQrjmJ1mzFdev1WXtvw/omTGBpnzmIH0l
AlzmFzqQ+sbn/kvo4H0eaP/k3OSIOnnCuluZhHZvmTQf4+aoUE0R4GIq2Rb3ZHPLLxf8BXFDPHi5
zNMpqUcQMTA8fzzOxsN1dzmEPCHH9+pAHjyjEPykCkk/MJoL+EAZPDAw4OgCxFA7isuJSdw8C2NY
e6ly+4c54lN2xPYUQyHkEeaNL8IaXI8JEgGDKe+sz+8pyToIOCPmw9/1umTMtwGPYxWDwVFwHYu2
FYA+U+HJVhhx5NKiPjAqHKIXGbVHRLOPltFl6+49emLloiZ/U56eBKcx1h70ImC79ygYLv8H/ibK
RWIT4LVw4iVF6Xof3tdNFz3sX7RqHnWoQMwbL88sQcNIrphDxZva27KPfO2jkZMBTf5N3YZabGey
E8M/MiIe1GBOyy4zOSDDbF2TeSA23NiF4/E8RlsXNvQxdQ3JR+PeIqnsWqtCuhoxI4AiewxYuAUt
gPmju0QuVgD6f+wM/JBAo97RtLTU8+QbA/cPCsHTkpp7M43Fb+kjdTGubWbCLX3jqB7afEvMxlC2
P7aIFaj+h0is98JTg7HQswLvZRkw0AyH6D2S1BRUB9MliHpAqpLXO+qXYNG3K/uXfcVpwQCANVVL
l6MTplWPHahoDT84hDQ7Kwf7Jaj4hGmXNERy0ZdTcqpm5KKctmQqiTg5AcrByl0DgpdeCfCPN0uN
5y27O3LtkWlwZ0skV1XZ9Bwhj7KFM+t0Qs7xbWyGlrFpwXN19FFQ+g0/1ITY4NIE4HgG+EJWd3/l
DsOgKVj+jEPagWz/PBgyBJGGMcBOUkCs//erfgK9uZbppI8Hd+0xopImeo7WVpILfly0Y6s+jgMd
ipCX1c82lijRRPxP6197sBYneBsJ40miEuky7oDghOpXmJPuEmLFvnkykgsfoQE5FY97fNOnm+jq
YuZ1jHEiNR5/zE1vX2jnzjIrE+XAvleh58YHTFCNFRAIIUMqF0T9o18fHxkMx3cFNXl0VrRAlEZh
xhYPBCk0rPUTeOSQiqp84A5/rj8OcqMl1a+UIJcshRnBm+B1cGHEO5mQkI4KIpllopJXPR7Hpmkq
uQcGNEBcLEqi7+Ltbczt5zCwC1wvnW4NTj++eBa+OSK+jQD4+XJqAC5WPULfzRKaBNrrGn4HF9Zu
AESjwkrn3L8es0q3zB2oY5oIz3yAnG1QvN4nywZ7dYgNUQLMA60CAU0L37lC1HqG95P97zktvlrD
TXXOt+JEh/vrxWYLDl/ZJBbk55ZUiz9aFNQ8Gs2SwWW3P55sWB5VcXpCCYcNYROu5wsHES+do2GJ
+/kLMYOpdygs6RjmonnVBeFBfT7LmWmXmfxIaNOoh1z3+S4uTMLa57nvK3KRDm7GqGRpn3ufVFiy
BsR8o7BBqGyGp48Sb7SR7tBXLnjxmtmwD+qBsntnlr+qjXXukPdy6MQmk53f0shYxhcerx5zXd64
etBPdpc1/O3a9ogpwke2hOsuiwX8vrojjCG2ATRTVTAwoYjjIwrdd2coMth3JP0rM8A1jCynDHBX
eEcPuCSFGeaMLMacRniQCQwQ9hQojaqcushqyD1JktZpoBHrZvgIlvKtGdIThhqU3S5RHqbgGV6v
RhteCf45uk5w3UL4zAND24MRG7SsxF2lM0PIrqYPzqHRkqpRR9nrEa1epstbLuYsF3FCO7lK9DH1
s0D3JTfRiXPp6EcKY10I++VvSL3UpnyuifeuvHn7ZDvIEUX3r/1rE96tfmCdIeQ2BGBYXNR4P779
cj8zeuRlQAX/wLas/OvJuROHJdj0W95x8FDE+ipAQaFOzN8nR+cL1sPTIidR0AeYc78C+xQGavvu
0DA8HFkj/pLTvEhZoCvfuAS3GeZgeGeFp1BzsknfPjHMox+0Bjed/8RoslSYOigyHLJz6hGOLcpk
wa8XgIzbv++aZYOaBgyNKilDZUX6+tGx2J6KDuA+Vejjw+vS+cKpumUM4DiagwFlsV3EKi7W/31r
x5mrRtHnPAmEVtjoXyVPR4VIZSdbm80uCEt0SoOLAIq3mBmTh6iElysE7wt3D6ewAew/15T1SQ6U
79hLNeKtOFyKDrTNoXI4k48tIoAq4FEyMs5kn34/8J5YIb0Rlt9/JOhxzo1J7TS8YsHdhRkGNo9t
/2iX6qfBao0JECQUoWCtHbTP+cxnBbDlDPwodD9+JlJvsQAo9Qj1B5/Ga+O/kEsmbcuIbRiU1OOi
PRz0P+U75JZ4q66a1nb8V/FUugbduI6jO5PSsTjRXZlPJdr6tL5uolF3wzhLkLqz0qjOvdQ0kCIi
T0t0RkX3WgAlh61ZF7j0pqwbNVJ/FU1Dxu7AYcNHP7THjN20C/A8wGw4lIC+lZkrFAqNq/ZRZ4oo
t+Qm02w=
`pragma protect end_protected
