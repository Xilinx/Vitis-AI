/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
FPGLUMyFuaQ37LtKrDJDcJpFRmyXtiM0yOz5IxJEKKib4meURYWjLX4hbkXcV8f8MTkZUzMghGHT
emzXur2r8fXKWmXKiRbUjv3OjVpIiK63kvrAPl0PMfuYEJeqFAG5Hw2ZIa9i8Pyu8r1T819Rw5jI
oxuicHf4hlMUVzbKknNhMaH8I+6xrEynMd1q2t1X2v0dxIzQr8atJR6pZjy9mLf6eYEUnpJbJK2/
jA39SsW0f6K2pkGCqQO+HrXORF1ae4lLRgGl7LwPM34gyUvh4FyYMGx71i7mleiB34JMmmrAF5FX
q4BYdTVjRdq4n4ff5GKSh7F6qa9KztRheMUC7A==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="EaCzIzKb6KBxAMRTaQERKgv0xZapdaUBSOUcJxrfh1k="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 880)
`pragma protect data_block
B5WbXoRsjRJSt5Da1QGvlxx5dP3KrOCAd9Ls+Bq3VsPLLbY6LNUGcYGNCPBnwSLBg/66tizTkexR
oDoxgt5Ffpb0w8mYnzngaf9VDX8oPj/GQhjyh4xxPyVliau5kgg8SvEw4GILQF03kl9tt0Pa9HFH
ep2xWME5ID4M1S5rZmNt/yTUT8z/dopvrgHc7fa14NGjpds2wC2Mg2E18TxTZMNB+G2pNMsKhi1x
EKfcaniV7TPO3X7B8aPWOe1o+5eIqGQ+EmIb26SfTsEziD+X3qA/npxVcfdjny/05dgPfrMHwI1p
rVHw8MayaVKYBEbX14ickJgp3Odn0xZyJxbY+VN+RuCt0GW39ffUuNA1YPkE69KVZdyIfppaGKUI
TJkXGE5/2gKkTFDJ32O0CQtCvPOcLOLaIBMYuBIzSxx4G+JjFRjkIhnF2ZQl9L0Rtdgi3xeVrO9V
9ZMNXuHjBH5HIqYddIdEPD0MOKNvO4BdnkxOctuHa8vS89QrKN6CYrAllkH8BJFdbWR90+pWNYeu
ExcWt0hDbHoOdxiKwhxtMvIrkvFQlcaW6l6LV/IhvzJRZ+ac0Ye/c+5ihmbGIYgUmn6yJMWIoeo3
8wQEsQ9uLZ9v8WY0ovgXL70BQxcvb0U/Xmg6GQrF7eJu2Ou5CSTZvr3ust1SAc6tvMvhQxVfdHJQ
K+kmYhLEK66yHH4TbpxuWWAWtsvw5+EzvR4mIStJ705JsYPSZignVM3dj1pTNFuPP+cKkPJW0CYD
dh2WDOdXP1/jVa6vgItvGZUN6D3ngoNMs3PgkX7Ggbw3PKKgAfTBr52m0I9efdsektd7LNgumeei
e/mgfT+waqFayQd+7kNi637wRNQHmniUJ3rMieSOvwmS4DqAwvdmuZAQF8DqfSvtWpMv0ixla0ZG
T5X95Qwfc1M1VwoewDVR6PT4EehKp3+c/Y7WmT+mLyiSseEwYvpkXZnafHA+DDRgTiFiao6oLQjA
zbqn3GdZxWlKLftr+UnKHcsIBbewAncFWAqeCuQ9BzUINbJ8cvhNYFLvzelf9xImPS3AAPSZcw/D
jok8amGOnuCCi6pf7cqFOwxB2quXuu5Ybi9lVCTo7xNE9kJ6X9EbXeDGhrIilWHIvHZd3lj/aYYa
O9FOzuwCa7Yr7PSpvNKQDF5QDSFvRxW0gQ==
`pragma protect end_protected

// 
