`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control decryption = (activity==simulation)? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
mBd155yWwopSxgsq7gzhjaF8ibJoBh+3IavZCa8IPzxj80vq9wOF1kEXu89uyrgWsmVUaVNrNJ99
wu9nKmCkIByDuSkDRxdEF6tJ9v+SqGmaL4gl/1mYoVE6mvDkwmNpTq4VJZxqmsKS6XbCi0c5Ft8A
tMf9TJgKZZ1BX70r1Owoqk+Su2T8oQw3qq9FReHf5XhlXmuv3qNKWNkc3ZkGGYSxdzr5MfC22xrU
nmcNqb3QLKFS3tIDNRA24ZaLs04Z5J8IRy3bSDVD9cGNHecGLg+PJ9qlm000aqL3LwZRjyjTp6T8
YPAn3mt/jXCsqKjeTd9oWByhMyRAigDp22qQZw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control decryption = (xilinx_activity==simulation)? "false" : "true"
`pragma protect end_toolblock="EltejxOFv4gyeNdq1t45PBJ/MNJoZvvwX91CO5JCzGw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 47616)
`pragma protect data_block
lNQQTMNGMp00jL/edOGdF2sVG0GXNsqZ8L2TmE9kuexEiiZX0v5eJdD+TlG680CXj9CZfhKT6W6+
IE/GK4YYgDx5aEaYVm3BBp/UCAVzzZk/HseLjQlmNnNM+ShMgOpoeKWzAWI/I+7TlWGoKhNOOMwI
A+XwQTsN/0xLnZ1pAsA8w/A8CqgmuV45/z25dJ8a3pHZnLWNzj26mFDor88xA905h1BMjzFYXVQu
mj3XhLazz02sLxF3cH8eEGV7EMaWZFGu2VvjyYadwf88XU0TkDk3VQ4HdGar7mRwQA/+/bKq+oyL
ZjSzGuypbstskbMo8f5qMAo+ONGlmwOIB+wrAuG93nF85Dx7qYpq3dYR4WKt4Nns4KRh0AtsRZtj
5Iez64J4AiNcf4SpdLidx+gbCifdc5jZwkBfM+SYUL2RoJp7Q8JSCqiRvNCxw5E717X+8RpzhAmQ
ldcV6m158TcUJtouqR9wrkEErmzYUzG+Xvx0rf8TPDKXxtB4YTbNK1k5mLIAZDICRD3pGtHdwtlX
LTTD5QYwBdezSk7+5D+V5WUrO+Ov/EBWgUdqwHdg8GBKNKjOYUmYreu9KLhLVJDQjDfnB2UdT6KX
3HSMpSCzIkXinHCGil8bcf7/Poa0jaMpB7Tei7ciDlzitW3lyewfoyf9qGvzxO4wsWyLCn7q73fX
t04WxxYcO36GkdYkuA5WNURB5WcLcEMz5CoexQfAjjVDywStxIqPIK50Aduy/fDwySG4JAvw+tLL
cA9592aIVcC3b0rUdLnq3v6gJu1YYG6Ex1ot4UuxS0fuExGQEQGDi5+1T0zt/Jw20/MosUf/BG/H
bU1FHIdsAm6uft+7I5naFNkYDFv6fsxdnfu/MX95XWwn1vRNirzvgSpKb5hcd4QOYknPGL4xojGp
sZ/5G0qZehfOcSBTUwqBYwtM4gmLkZgrLiUWeW/+FNXWDn0NY2ltMbohM50vnoaoynLxGMkjWGST
+ShwzZPpZgxAGOV07TAjXi7/AwOrnFMZ42eEcNsk4cV/EWOJETvBK4Qlx5qPY9o0o6lB5GCXTCjc
GpUq9Vi/wS4HEv7p4La2Iy5ASpUbNMYEsYTWZMktcrmykrT4NgrdzYqkEHknZckgfCRGierywkEF
ffRmYNfmSUx4KJP/YU/cGJsbeobPmiKZQEwR5v+xrb9sE+uAhmOujqFQrqe+CRGr/pWjpDaAyyHz
LDwuJmsbQYX4VypaPZ7NnaLUf+MRSnS21BPhtzjoF6/ggxNB5IPGA00RUSfaKCMqfd307h0No9j8
m1+KHbqcOfKaDHoEQC1qF2XgfMP3WqT6Q8NFC6mYpk4+Gt48loiVHxPmMvh4pJ1M1d1HaeEpzIk7
MAlQNt5dzEA8NpZ1UG9NHfzbDxckXU1kXeyXNl0KSVmLRt8xz1VTvexGiyBXRNd4tNs0+Lz+JJRn
c6sEGMgIuERz1/QSA8Rfy8KE7uUyTaHkGwL8sCbJUHoON64QEv+KGEims3bbq1hGj+Cuex6/orFe
X8Kvbq2NWQWOdsGYZbV3M1+OufEsYub6GoVEdr3VyC8hpnEBTtZNDYssB76NMYdegDpJKgCkq/Gv
kxA0Ty1xFbHRg7Q9B3Q6sTvkFdw9zzLTv9sTFJHJ52tQ++lsPZR14o7zUvipea/uQhyVA0zqdKCv
51quvipox+y/jsidDJuzXMf9MIbk0DHxQfXCo3CTV7+Vksfg70bgsdMuQjof4m++lDmbjJ3NPrrM
VOCSwYxLVJYL91MxvFH+ViTAdsHhnk9sdOnGXEDtFX6D6XGY0rGARbAXBtwN9LQSpiAbhW91Fg5f
XKpovZgTVnJ6eThuGrNf+ZWJBU26Q7I0p3UEOYuNUvDqOzVRGgFjaSUtoUk81n0Bf1QJES7d7H+w
jO1G0xSnIw2PtPiPRMMIrIKhqHKOvo8VGahaarTZLJYC5kSGRzNH3q/0kXvh7GL7mjCw1u2Xwlbc
mjCTwqANijKOT2nbNXg9Mv1V9nuqwdgqAZMpR74O/iA7GqBTKWic0UHosw1KHvDRIDmKyhfP/osm
Xtu+eZgRDxLWpWbe6wQycEGRGdxk1BD8AUpGKdT0XRQ9OnMAMl9tgG1gXy/rrqekFFkOt3kFZYjH
Fh/XTjIoavPG5S5yvGZFGZ8D+g6DYTVb7tAhir59cFL1jYQsn8rT2qTEjglIO0ALCAiJYwrUpX92
nqnnoUpQtYvsivHTEYBdFZ6Njd5HwaZQkeedAeCT9BLOja/2oft7Jqr0tWAzKb+TYaEnywCUWkel
R82evT7m5N6vPcZl6rfiYhaSchm40nOYFMVr7s2/Poia9b6C1MHxazn+OtbuicybA1s3zjJ87FCE
1RjjMg3ZhIjKwI04tI1C9GArMuZgfxTYu4VQuBqOF7HpFo93f0tZKSSL5LHtO2gl4j+P/FoK4Cp7
EihEV/Iifx0ICjzazuRyndIKC921q3i4g0qeFZOt4WFBg4dbmNjfp08V2/slWTrBazcBh0eIMwd1
4pwtdyPgqhvsT0gc5LEdag3r0fMxXhKblQAgMOa/jQ3Y2pWKh+opBNyCjfzSOwYl+EbLDrvus6Sz
DBzwKgHDEvO1huMgTI0jfb5AuOTrk0NwQaLR2UaySe1qgo7PQNophl9/pes0dVTJZzL11IIulz18
fhg9LcIs2bRA5Q5T1PExEERJ+LVtoDRk4lkc3kryMLZITLmVSiXAgjfwAGveR80C7DdFFpZEN6K6
H6fF/v/RDi4ByE22B3Yywvs0fJE4Z6FsYryxeMUrdQ5tMOXdITQCCMoV8JAB2yX7eRM5uJY+oVMa
uI+b+YHCiKp5u8OPEFG6gPKpS8SkxmkQtHQvJGFFBkpJ2JALZBkGBx4oGEezAYL1WMIuPnkKc85n
t5J/qUrIURMlVk0i1rhG3EW/0YuOiLp7djXHwmb8FS9L7ZisC1EAqIUXRte7ad2h4pe9m82nsfuB
w4Wvdp4LY0qP9Ef7n7ycinw7dfeQ4RUOuYjhbqCMHRLBt3ZQQmlsqrGLOwXVE6r/puJ9PqAYfW8y
SpvOh/rUKDbGDWQSrAxuY5F+7Bv1pHx41WtZTrFrSgpso7pcRLSp9jQw+pHrsoJ8lzcbcTSZAf3L
WtqWJdtWfcrETPmtlmt4zrjJLbbkthqa6B9r+Vq/k/IWlNvuR5ZzWQHa3rBMqfqVyITLZNfKZ+KU
7k6yVhrn+6I/bmmpqmeAIKGrs7QMiv3YLtTfB+oc+AFih5xP/eA4DPn8Tavjq4kakwYIZWZjjViw
Mq2uebf+IcjwueuqGKmWyylM3cNdZd3p1Rgak+lXT/SK6XkKbU9KG/Y5M9/wPsaEbli4mHdqciTL
PZAhtah57938QUkKikWofUDMgEA+XL0eaRXIeP6m2Fzrwew7vvH2xbAoBkgds9l+OnBentvOPUP8
XwXejsBBxBSW3pk1z8uuPpmy0ocT/rvV1ZXjMqRXF2XOEoBoIn0eoQlqAK9jBnOwK0sIG2Roeu61
Pk2kYs6XdLN7U+Y+WK3QvkC1Fz9RzYCKsvRgkhEhRV2NfqhQ8tX++uY+nitKUvsAY3vMNrNqJQEu
8JVcpNpFlXmFER+AtqRsg2aopfhfHgd3iFHL4mlwE8v5Nlvu36fBowyAaULAvf1BXSgAL137343b
nl8cvJunnfyp2dHj7HpcZjbw07X0dkoiovixR1CAqXl6c/iEPxshuG0tzSgiVPdJFbTke6KZM+A5
oHC9fDNIdxaHU8d6HplkPKK4lUlU5hBzFl81fTbaaIOGnvf5CEunyLiHjdQkH/MDx4/GWfCso4Ol
eX3NCLe5+ZW2AkwszPqg6ow7sGiJ8MdwF8u6Q49XH/7jmVXY4kCox5Jzn1uiL0mUB3GBcZuTU3AD
t8DoEOyzTpQfHrkV2LF0IF4lGIjnAriNQBWxFsZmiraXHVFrlptHZCfAPGEpqRjrH5x4TNxBKqt7
obeDZiXg14VqtDEZUjoo2r8PFAiygvtxB36uyTWD9AWBvZqyydteogAodfsUbXfzSlOI56Dax/hZ
qCr833nM7afHaMtPsYOOaQydYdYk8Kz9ko2qwBjCPjw9WTCBjK0TtOdlAyUDEnucx1P/MFNc7Z1Y
P2u8/W6KOIMII9+jn/jOKvWqImW9gNO0GQALz0vi+lPrWxyxAqIUDAIWSjD+hoAoToo7SGQm90m4
od7+v9US/RkF2rt7x/zQlqlpql0XCtRU/CJZ9YGOE6mQEntxQbcpJjBJIbOh8i984zb9GPKee7g3
rZtdGC8BdPDjTXqpUB9YiEQyf0EP1+DnWy3ZPrUfFHWBysTezOIKhphcVmiwrm+0wW+LA0G6peES
q8nxWOo6S3xDSwyWFSLqnfYd1nU9Jc9cQfMCS9Q9+pzkxCIQhIxEhtcF7yRLz1YNayRrnudSNHr3
6fR12ZhwqKW2tN+m9GqBFeu2WgnFX9YZ9Y9OAIRL1PiDPtUXe9YmKv5yXDaWiLwx8O8aMcJlvSv6
IQySJmSkVdNj0UkcqyIpigsapr4q/GTq7WzqLkxjsRtXNxYWkua9FFXfBdWNUiAA20P8JQkCDjth
0jnsagRhVqaWlzyaEeJLieLlLhlagz2mBBI7Fzijirb31IVaS5xOLv8BTVmn+epefs5y1KsbEFZF
U0xwFUhqAqEmhBBw+F1sJsHEjbd7kekUevud6tvsRZxv7Np8iFscz/MUOf6r/+wQL7xRSbZOoQ+r
PI6iVI8aGW9nRJmkGcoFLRGvLPNh27m8HstqpjzMB1+9BFYy5Sa02ckfSu7i62TLAGk/B1bhny8C
1B07QJGOI7+d5REVrToDT0UDbwi1m82gGzEnlx6Zi46EfOd243Sg4dByWakHutsXuF8jTl1dYkno
hPJh89RGXz/PDjOhPSrpzWvNtdnvmrXsr7JjGg8STGLGe4hIZ4/UgDWnSKzqIomoWBPpx8gcW1v0
ua+03ZA1ky+KNE06KczkgQ/Roam1oXKWv6p119v4Ypxq/tKdyxHH22yMdfHyhx5axXowgje+kmKZ
ZAmfw9OZ8SgGQUiIMAWllqmjskTgIxGSJbqLHV93JJAhef6q1xM6yNvzqCKF0k/ChNJ2ZmD+ebjz
UJcJcVTWU8K5XZVtuH4vEcvOKZ6tXNrPpkllk/ZVupb+yIr7oDBFAEN5guanQ6AUyCl6EF+1xaJk
btWxq8w6N2oLoMzk7A1bx8eu059xNvSj3MkGk9QSMQFjAXjkcRnjmo6wWZo5krNuGptPqtrJOnfB
FzsZY0yreb8AW4eZOnWSgQm5QgbY30AmR3d+bvOmNZwNKuWk7Cv5dIPyJl1fl4wuRIFUoXBE50OC
13n5PiJ8vGVXrEokTvAw+DTJe2Wgo7/yW5Jo26G8sn35fpV++ywKxlC1vMSR6/BMZjPSVBV9Vl6R
NXVNV8JDckdYMQCH/y+CQDLQOSF6hFsnhCod+vpHmspZks00A63goy1HKxvixHn+G19PVYmMsP/F
vHMC1MsKFMvT7cO11yJXgQqiIjFVCNpM0kjDvO/XOHJFI6r4WejrCJI2EbpGHTzwOcZ4P4ma6vk2
Rp4JdA3UZA/tkTg9U+R60PkPvRtbSEo5Ih5XImditGKUagxf1OEtB7RRqRuktIsSAEyEz969+SEg
9OmhO8CTYELE/7eYaQuvNKFQ1PrnZVG8keVgJdMt+gugPuUxbSIhg+x5ZqD3fyy30P1HhgpcpmAR
DrpjSoI+ZPFULoygoP3lpevacM0qY+PDqZ334KgduZy5ihAPzHnBwrOXptWIMWH/J0vxxll1BIR3
hsPFtF9km8WVna2W3HAx27ESXVV242aeKOY7UM797s9Pdbs39oxowI+jcIU8CKqtLTVGU3OW+X3P
ks9gRSzLVGErHDQfl6kpJ646Wak957Cp8gNS6y4soiwNNj7hi/Xf4x4fnzPQ+a9TteKXtB8MKLIS
3HYVqjznT+siB3OOvao6OHvRqIDhUS9ykBoBQX1iioMctnbllmRNLmPMiwwCTQ3DQOq8ewNQ6gUZ
eT6DJlmuZlnMYdBwBYvMGTM0oQelj59VIAFCsC+Gn5PVNg38fyzeAR14QDyLQYPGXQfSIRl0W2lY
VoJs/SuF5VdfqvwZmmGSl4o2DrDzIti+F3wICcP4b4uGmFJXBzUL1x7iqWKk4f0FZkoARSKKWmE/
O3nSQFZmk10W09pLKRuaDQtQLwMXmMwLgaUaUXFzfQSC/GVUiJg8+ob+dtwQzADqNF8EC9k9RYbW
PWtKNNVm4/AE7CGIehB+M5cC1EN5dNM/LMFsDWfACP1aCa8KdEx2amkA0Pvp0MKwrJqlI+qdSRCw
EQHTgMP+dMBgYs73Abv970pTckr0Wgs0yKGHdSsff6R3Y0JJGjDhJmLa4y9izZRAJRVGHAdqkN/e
zghS3i0fULB0LXdAhjb/1BLF04SsGS6hdZYp+sdjuYriAAfrKx0AxofSzL5q8LtOLea1cMb51tEi
nksSqMusxPul4ejD4LIM3eLtN/x+pYY/BMDEbz/t7eWZTA8msS30AjpRgqcSk4cRIB7IDWFdoz4E
jNugpc6dVztI2srs34PjXghH3N0K4yWafKZGNvq5XscdyRAYyDaHqVz5dEWm5LIXFs2zMtzTmL84
NlSuQSKAyCwR++KEpM2LRR/MR/KGQpBUZ8JMTGmgYTc1tnEwZdwNhsGT7KvwOUQkZ8xceOszQIdF
e2jV4T88VBMvlELiQ3Ql3aTKYi/rMYN90sC5e3UA+SjOwalfM/KSwphphcSBVPCdngfE+rYA0byl
ulV1eUK2TUaVaucXkPnDpcP4CCeoLWExSo0JGzs/gAtLkleJk5bzph4RIgaLC/RK4ql/kdjqa24t
tyGJ2XtLprGZM5kdtAKh2FLdVsntEAxmM8gmiBYMMYOKvelpqbiCK4LDseYgSVUHhR75E8Tj/B7m
K5QBu9wQDM8/f8UIQYWRwd1ifL0zZ9jTHBjZe7y4vFrvja/N5kjsn7FrPTeCY7mYDOOZeTbJ1CIr
8bB3QK4R9QINaNv+zE3AozpHYwC9BBA7ryPndrq089eUdeRxPRKq6rQLJE60UahuHnTrISHgwTt8
DoCZoUrPIIFflJwP+3Xo23eknigmu7gmZRwBGBC9qcE87z9c0pFkRzc6boeVDyOvuJWhSMMXTfb0
iVTP/qR7YxkkPTvulqt/eTL7H9QLngCZD2cyn4v1wwvRyPuRvwQHux5kfAkcX5tBxHE3nm8x37+H
ErQu7zaTM4R+yWauC+FlkHNCyhILSJ4MCgqP9B0Jc+N+IBrZAk+jaPBpCeBku6WbzEsDi5R7/clv
4Qys6NC9BoU9mPLur7L9a/aqlbG+lTB6Ck5ouyQ4IRk4TJRx8qFENyvQQ24xnnVmg6JYHhGUAVLb
99Nhz4hj6Ewddn04hvZ2e2r1Dg86MU47F8EveCgqA4vQVoHUrDHVYHzVdPtRZhHn3elL5ptc43nS
oqzGcB8PPFtc5tGdVQN5nrQtr6wzB4y/fgilic7NoziYCKgsudDjjelZ2sM/yz/nk0sPwk2Qf+zR
0H7ByBSRzx1e5FBp2siLg13Rh9FD/EXWz3QoLl0B7nF4m5NAxT70A26eT3CnjSxe4cLuFpg3LBGu
NP5HJBzdNXtPghBnbEa+02dIpviX4VgQw2vHGUQS5wYP6PESXLiJDGEPVKUKOyMazhIYRNVa6TjL
KrA7IAQD9h8cxPv2SpIJL+5jAW8SS8ajo1xtuZzy5Mj3gPo9sSQBOu0S6KJGTKUvDvBnE+FAfFRk
mknHi++2yMYcid41EcxwwmS+QTYQusRjpvzmJrtwLl1nIm4yWKIRLYmEJ05uA9lhpgduOYuKpxkB
Fkjr5iv2xS4d25/6i2UaDunnkL65ZpPZmFCRTDwElB4WW5d84/OIIbVt8bSTXILS/EX3gOu2VUe3
tFrxSboWN/FCtFnOFsL1A8hEMu3dYpahwKMzYzsqE4xyi22jVAMg/fkbDCngBBtJPxT92lF6KyNA
R9KLPIPfFHa99eWe1+FIawSFkkJK9w7M+TjaG5Gx/QvWQO8NSJxq91158x24nnTOcyIVWbsmiFYy
C408vwbEUAVqpBO/r6gN/gZEXEZBshTC43qSBLEYS7uWAo+5ngnc6q7UgelAjpJ8MyXDoO/4jDFP
Jz9xq32aCXnAMK2vcPS72dTBrrkgYhmsywLzKXWN4FRO5ujXPJyHgzX8RxEk2jKEahmkbdvXxrIb
vbJ//bNJxf6n5+vzazkUT8k7mhjMCLMYxQ+n8ZUIChvxN/b6qGew/IkgIc0tOJ9ik4JVAGzY808/
vQLhctUILBgVdcnD27a/pLJ+MIlgjfbnD+WqS3tKeka3dWeyPmZ9slB6gEInxSXfBjfiTFBHeoAM
p5LjgarQal+AGZ0yKySAeAW7M1BPef4NQpTGWIt2mebQpeKtsXqvnuCsE4iQ18Awna8eNDtWZ/13
AciDH4kGZ+WcMrhIL2bJMk8J/NVePaWu/onusGVSI/jhGmMXTpc4VCf6vKVwjk1k4zU+ga6oTsbs
qbSgQ8RVxNLQLfSwsdmU/ryWnnsA2rffVxPtCWTn4Id1P01xfLh4Mlb/0pbkx4+VjZ6mXs8rCP6/
pzmUzrcOnQN0W1FEBem4hA07TfeeI4s4BfyHzGicGB7q8bg+N2w1QjOPsy0Z5O0qRJrhA/aYHp6A
Lce22A4hjIHBGSHCmDzegqSAZAcN9Uah/JjPLaoJH6+LO8uSpJU5PRD+kVVmy4OqYOu7ow6Dg/3n
V+wKn7Ei96GUD5Jpovgs4NtD2gu3ZRzWO5SZonCWEpKnlthA42zyptDDmKjUmUhf3l+mPjZ89Jlr
Hl3vFco95YC7Lqg1rTWudHKWSY9d3KmFw/N/HZSapWjVJXILjqDck4MVG6ZOBXB1SKxmClKBqfM6
2mtH8igRtkC3Wo7GhOnmKizdN1nEuNXJJ/2oatsgtdCdQNHFhIblPB+ppGHASrfCWNp4j8WTlc50
leSGMk1I39Vh8SYWRjI3TX63ev1DiyKzqBuMbrXRrKobTCSM9IqvGBILU0boM0RoaLTnTHxo0JNs
GnVpgjxiSGskrqjJSB8LqZ2UhiqF5qB94x4/jPjYrAF6iwXGjnQ2EZ5r+WIy/9q3ZE/SCDhBbxwK
I1eo5IZSkoZndawTfkGeXDdnCsUmjmG/sY0pjActNFbZh3s/OYooJqjSjwSmm8kgBMEQa4I5K7eE
E9AneTRyPJ80klCWNoQbEaZBR5HyY+MrWZ/2dt+D4H71tbDgqFEKAnoQAnPbRl+mG73oYcxh6Bfq
JPPiub4Ra5hlNgp+LqQ5OxakVEskXWV5ZAbSGgR02z56A6T/nWmWG/pwqiBcx8aA3twpFWbtvl0m
6zxl7HWXBrtSiiD0a+2bKF8O8mipgGrnRMZXyz+co4oRUfoncFqn1o15DtiPT5KhdBu7XYgIgtdd
P+W2OAt7E9WCyqBZxT2u1Zguat3cfI267ud6Z0dosy+YuFCBHSMXLCQNO03vtB8hP6G2XGxORIsM
OVU/n9wh7mRCtP+Tk0QSQpmrmN2I9vLabs/rz1YaASXEG3mL8kBTvDohdaR6wz1PFjAkIKkBGgAs
0of6HeE2HWzGKHG0W2xAQwLT/M/a6GpxTfVrubT/t8DTF5RcFAH+bTJCM4WNPSqelPDyIPQGyVCY
gOjXLiAHvs/ZraB2vTV7VioQZjIo/1LHd6vkHMB4Y2a3DHxgOk1I1rpXjztkkbwW2pPV+plxlPQv
EOm9yKpAldcLH2tVSV2mrZWU+KGTBLDJPvGK6JjJ8vvgrztoC8j4QSdAHJlzG3OSRBI9vcsk53jU
g9yVtHvi1CkyMoK3X2zEZXUObzjNcYjFZtz1julWsR+cuofwwoCfJoAM1yX+lvrtHMz6kQ2RT33Y
hjaPJ9eePQGG3XHDp87s/md4G0ikNRxr7zG2Q1gtxWaq5mLpIUCom4OM3vjmpDWZuxrdgXVDWzT2
zuXA26nyICp9n76PXIGsav80YwIoqzTcWXsG6yqYNtjQQ8B2Wfi8imIgdm4TwFhAHSbXv4hMtOHx
NeV1154vsxjG61pgPHYBO867LkfYRRyiwHPbD9idH9jan0rSedj7P+Yi6cEwV7bJ1TilETnDjKxr
qSWNi+38VZOng6Xv4wSdndKcjis2wdG1PBLM1P55WX2PDOR6OR906P7mab1jcZD9lHKwhFhwP/Dq
qLfecNJMHvv8YWwWkzoftDgb2WH3FddCFz2eaTMmlSWVNg0FCUMOS1h4xcW+ZgscqtJgRjzSWzf6
trMOnasb02JfahRBoU7k3NA/fG8jJX/+NOpq9EkOvyK9b8opSumw/a5FWaVlHF46t2F2YAusbivr
3AMQvcbVnD7/J/xvCzJDfLcSBmWQgL7YVimTqElBkrPRzk6zoSQbU+x2N/4OC9Dt92SLjHzuJmII
xAelJdUvP6mTiL27vXtZXtUMs07Hetj6O6mm5U7VsZXy90qcS4uhtqi83oNIU4E1+2MUfPV6wQGA
jIJp2R3svmnNbMeTD/bjKyUMda4Pap16pdpiI54lwj8rrxLHPi6OnFSCK6x5bCB3vYcIbm8pLIns
PRxnVdEfRjTFrtZmmuja/wIGLFTewGpgfg0LXd9nPUVoIxN9T0y9bMvNSTFrQyKX8PhiNJRZ2OJX
YMl+xAzOOJZ8n3M+oBTVDt1REcc/PobxDjGbwkCG06++BdoGEN96OmuRnYmdvDG1RI7aG2e/htql
P0wTTBVFw4PbrxUat7OW4c8L+GEbO5EDkgAHUvHC6StC6DMiQ62cqXUCnos4M0E7YoHxQO+JEJu5
tV5Kg0aWyucRvly0XWku5ZSJlS7+jSgJyUsKlVcOwkRPxBg2EsyMpzItxUT7D/qcNd8Kwm3Cr9db
bwLH7Dmtqn1ovPfi3IdVo3RBX9g+B3mv5vv+H9MLxVqt56sCfT5r8EGY/3NB2B8rE0NF856pVWLS
X8+76sM1cJPNdgznnpH+GV0ir5CFYkZOjnWm+veKPywC5CUtEX12QncqWTEyE+MTULqfRjKXKhS3
wCmzNOj/YlqPjPfXtMYstgkFLOaeUxlPNcs+2RQIqU3jD+nwgV7e6sjww5kRRL+yT3wtOyxHeXFz
Akhn0cdgfVsca9KOje/rSD7ANDUrnfOcgBSmZmZwl+cHDpCRRsrdOvORTYmxQfk8he7+JDeZSCD0
sE0N0cu85C07TtROBWS479anHd32MTdONVZMDuXr+iD9+VjZwlDfpfoTb/6hIpdA8J59l+TbHEi0
akMjLq/aAOX2f/zt+4xeCIFub0nvA/CF2nsd27a86abB9Vd4AOWzWO/2nQj8xzH5xIZ7iPcJUDr/
phjeSueTT3MpbQFf1gLVQ0OIRCIrwJlFdGH2zP5G+N4ZLA5p1zB5KONDNvYQomHuYkFVYF+zRolq
LNPjBcf5UOOMdvsMunxgRj2N3pLJ3g0wuZmrPiUIlmQyoX/l6LqvhTQe0b2wa48OrK/T7kQVY4Yq
/AW9NhvK10JXwKgA1GPOQf8YLuPXM58dhdz7Ra4cqv6R+OjvPSGGRe5nf9KEcfVLeLYjAifsCLG2
MBeLEaiSQBxnnNtbwXySaXffO5/PskEgoJBpT7YblMAN7yLKnexUwL3uoVS+UUSa4Mmpeop7D/JY
vy4YRD9insGYBhV/FQsqx+V03ULgy1FJbxqPGiHYQyDFYKBW8Bc3NZWq4YyI0SFnEyc+r57tL+BK
UCL+oX9JmLir1QZXZIakJLg25asuUJArIbGeZr7xe/TL/Z6A1pm3bbUwFaDwzsffXfy8nR6onvi+
mSoAGeQA00MZjO+fQFhf/7MXj6NkFxAitBYJzti5fOQHEpfg7LouLHEXSAYfKd6z4FredX0hssBo
+EK6fcV8lRM9p2VKXrpDmIaMJi6J9YCmfb5hIon532EHdjdDBc/GbP0s0Z6VPh7Hmoz7rLGyl3HM
kadtEa/J7+2RtJpoOgtXE5MiEuG2pn1Q3eQZ4UoSlzhRikaHU/uoFlDCTY4OyO943baqw1NeR+Xy
VhIZF34t8742/KSKLrz1a87qYQd1nccGIDYOfqPQ/kAYNrbwZ7I4+YlSjzSWd7i9mWCY4vu8yQpc
MpYJYlnqk5+c7E0N57+Ut+HzPP4zZG+9hHdwAxH+l3u6pLAsiM0uXZgE7DRbmrnCmPtJHiOyr1V4
z5o7IcbrR16Et6I50KWcVMR29yRYGuavDiSHvw1maUjcTdFJFap0by8GVI/RfbsGxi88sirpqt+Y
HmBMEY4za6obYXo/TweTypTZkhJI93Lu6adfFz+kzK3Nw+HyeYkb7AC8Q6gdkvNgeWi184NQGzoV
ivAtzJ+Vc/Oq4SCycasgsrqD/7Fhq6pwv7Fe7B6hhUalpRGbhPxMLtqyDIJlNqcotJjLuSW9wgzO
cmtNS6SP+Jbi955zDMpERrPlYV1hSw0PCTd2joFcRcYUwMl6cp6RcjDjcY1/Ls+8htUHezHyhnmv
DPex/8fLcVu0GOKlFUEAn9avHsZdVELj/z3SktFhzzKc0PR3T78fngRAK/nxQ7h8YJG82YAFWLNw
HnRaDqEmofJxe/U7jrx9NuBmepgJDjTiYuiuO9/LcYN39CKNPTlPaLfJwBV47U6U157NGkob+nIY
bYM9swRxyZpqDx4Zshaw6+rjXRcQWGgP4+oRC+IqQi0+fA+ChPMIAUn0lmc+9f1IfBabDVIyNhB5
On/3Lt6RMqaw/SjshFRNXww7SiIVHSyAMuNNMLWPhhHdd48kLFv85Ve67RQiyKCaOQbpzd8tTJ08
KVB+kqoaOs5cWl/PafFjqcQZK/mU+1Z8iCj+4givn534oOt0d+IRZ6zQvbii3ZbUkiLAy0zgJvLG
j2+mhJ1Cu33vstPTvodX0K2yX3PiRDO4rv41IszQf/y6obhoJHW4N/+K3yn4GNIJ/1GawUY54Uvc
/AD1kiWzpV4y66kgWfHCxayeKC5WOSS9lPFoYM4TA+Vlr2CM+m36ewI+xzqU2YBdE/0pS7pMwZ9q
CAopsKmZYBuK8jX0QVPEQwpyvcawXUu9NuLMdWymkyMPJhd+6e0pyBpUvGxdtRNEu/4O4OXqNFeL
b4xQzqD8IaVwhf2wYitQIbPX06DQje2j0PhBKtGvUSoYYmiwgdl1bU4Vzx0c/R3VqMjfBcIsu/32
NLTYaA3u5ZqX5YIAER7z+cSqmEnnGPK49xmUvy1MdX1YCUQCMUGUbs64liFeyCDHeVash1h7rnYs
KPY63pRcSO8qkluys9kl1soB4wdto77QlTo57VykOE32JUdZS7ay58NJvIA/tZG8MH577AfYNolE
zHhN14V7p89W6WPcfYf6CdT7One6EB78uohX6AXQM2F3n5xmGo4zzUoqZvVY1UjaOaDN7CENPabt
L7mT1VfqrnRPsEj1w6AHKhYoKIcvcQv+cr8hfj554IeNxqvCZo2oYwuKM3xHVmwxsBiVXMoBiPPm
9/36e4NijjGB1uGEqA1mgeD1cgMoJMMz0F8KbhXOKCsZf9cyeTAJssSr0Y4Pj2kFgm4dfBF3dSUS
NBiawUH3wUWjuWvqr9R85Z8r0dov+qc3nOLLzA1UVVv4DkZhUD5wA9kJKZV8ObjJyMaxjXqTbIlH
EzzLUkV55NckknWoYUyA5SB10HbdpnSlPhc9Cvb/Ch5xHVBtVS+SjPPD+rVlheDtd6o+36xlXGw8
PFW1DIRsac+Dwkr0LZpAQG+paBNbN4jc2lBHYU10FYTWFmTlbT8uA+7mc4iDbodxt26h13sR8Xja
ZcIJKgqskDqKjJb9UdpaHJ6DEUQXBscaE/awKBRNpqY21+btbkooeMO1grinC3lr7l9olhTkrGn+
FN4zflBkW2SrIi71lihhJAF/fhXLZNlI420inmlYJN3NkBQajx1D1EOiw7HzNCvUj5kYhryIddob
O/A3VdYPMJ+BAZHvG3qfVNw1WgDJlkdzs6vjUg08HVDfcIMyiDLqQE9LIfbd+q5KLfg/1jqgVyPV
Rf/dgrUeRL6F2T+DPWr/wMaBD1bp9RLrQOWBFrhLYabx8qpeSJSzGEDTEgJAxOA7Oj2Dd7DPvEbe
cbwhBtTARcnRFTvI6zTcy33Pb7TMhNSpJ2Pp+RRqovIQJqgoLJfxvSG1dET9luamvps87wCEiyvF
BsZpIxrfoeHAa3cBFXUUZutunR5t5/UTA/ahv7vQQ6q/B2Z6e8BW+sHrSu815BC6+OAuK0jk0H2/
0AU1L20Sh4VIYje3LiWEwxlDgW8uEIUc2CzPfoaEB1Qi4q7yh5f+cvhW75XWhx2XgFtZGXKaAxkc
6J8NweSlT7WQekNH2ZRY5jWJ/4ed6fLyqjUPq5pC7pIUgE7uLD8fdm3SmouKZwBtL/+DoAiBtCN0
I9u70wVHXBeGOuvi9HAZL85B8UenjzBNkDPQZJTVAq0GQma5M6/pIEDK26/QmGNAHaF3ZY0LlJQW
CthhjFuXaUN7ZCDzb9MDvPlys1FoH+XWfTBaS5KF22wBcIowzSNB7OdVaWCIWnEUdN0975yOFBVM
ZjfTKoYTs/j9h9RXFxMvYpkcTncSnOTwDWcX62Vs5c2rBZjdrX5hLEfCM8NwmQtsY95hwdi7NRDn
xXSxRBawaHKoFLXwmOzAJHA7ZoOYIc2IHb/liKfvhMKCIPh4PemaEiV/nsmb2RqxmfU99tZUcVQf
rWbw/UKudQ1uO2iGf60ZWmCyENgvCS7avz6Bb12JgV/+KbMzlBadHdsvCi9eO/10qaAU8VhJr50v
gcWrOmjXd0EuNJVzcW8oOHr6g8abEQ+6vjymlflXeX+axmy3Z+jtGvxNZrsmAlzUxJVdk/+hx64B
2WjpwpXdSpkaobiVmiCfkwys3GqCBBErZMYFCaw3N1yBL2yootElhDqkMkCwQYmEjncb306YGzXf
Gt9ylq4QUspZkoaoD4Xnf1IS9iWAPcUnssTV5wmLRVujOqTheT3dgrBBxY2zKb/lHFxR6j5Ux81N
RwvnvjC2K86TniwU8RxPpbDiyxSuZ1iBgY73JJ6e5NIG+G0VISZ8mgi0b+g2LEEVkRYS1A2aHgwn
0htIbbC4qyN+QsrHbmYYyqA6t6M5xcoyP4bjgW5F4vLlsX0MX3QxIKbK3JQxX4CfAZO01W/VOgaL
g7Megxtk8pqzDx76AssBxudzLEAgJuDKZVAPcM+F1Xw4xAv62moSBpU+68LaU1B14uLvuDuZFut1
wR3cYVXcUxEtKs35ARbNrVLa6FYZ26US62CtFkD7iRGO2AjP5Bdrqsnc7c2xsZxshzmn9IBvEmhA
zTSzVqtGVmOQwgMujbxctYt9cRWaxwRzeTZxekaYzOBrSuOymUdInLealWo2LnNlVia1xof8aOvd
K00WUdURSLIIUaxY/vYU2YoQKclujlr08GVeQqnDgVuQDQ2bdDx6Q9tWAkowPYbym7yOq23nkRdP
NVbkqmrjd4Y9T2WpVm7asPJArX7Uk8Z2uTBSrMX9ZftKI92Y3yHYVw7uqB6zolEDORcRshXKRJRR
+Ch4NFKhDzzJccIMLkEPleZkb0PQwOEdBqkn5UG1uL8cz8VdHoMqnin23yAj7rPh7d8IBXsdRGMx
cJ8yXIBBQ8QA3roly1zlXhgpBvf7NhR/W8Rlyl09MCj7l/l9T4+9szotLIatTOxH158gqyaTv18h
ferepu2l+4wYEdNFyJ9RAjdAbZphelKd/qPj1as7Xw7AwVCXm9BXbop1XDStHV0bmGCNb+2dXh4s
D4jfvFe4mvgd6CHyMEyPxKjdKS/olQP1P4lDVx42o2R9oR00y/Yf/HJT/Leatsrw2QaYRNGieHyw
a+oAyRyX0pBw1IuE7Yr1QsM+XnIdq3jYU+xYtyfd72cTDTr5pyCidUYB+XrdDMPljds0DNk24DYr
5QCDZ/S4XOq4qH6GLNhwDbTCvdU/fdOg3ss5B0BllLsmdyeBs2Wrj7f1QogwsTxTAtspteW31BKg
gT6B3sr0p/bhFO7h7GQmbkNFtVtKJVNZ0RSAxPa1XU4Dh8AA27zFdq6/KWDVKInEpgk5qDI/ydJp
4JdsMWR/y7CKZMXvowUIUhNTXt/HAevKpzYwVZyIHlD2niMSv1ghY/7p7LzoDs837mZYIaOSBCTi
lBNqfEnryIT7Bf39CwUBujZ8GFbssEP/oCkwhj+ETVbb4Yc1NFSWBLWzL2RoAoiQ1zFpvUxEv0ld
jurNSXtsW/QC2jyQZ3l+j/pMTI8gqnmXIWYwQz6X42YxsYwnfjD+cH4J0iuhScwQZLGYOKj9X3Nw
wXxso0RiL1KJtUK3vOkSPK+a72493aoWLGTXrp6dK877pFgBHe03ei8wdqln+sJVMNRUH3ARK9r8
pSMOAZPxKrzyi+uGHDPCa+wTy62ClkPh5WuUlWQDzwP9XLDTjKGg4+Uz0AhUvSXW18i4cnReftSw
kKEglKx91FAFq30YNw/lYqLtGxT7Yw199qh3AVnzEI0gqRxnWvKM2mwatvAlDZFABSOWaIlgj4i5
yXQ+Dy7vQUzDdKyGw9tHsc5b/pIBCQumXO0/+dtDkzvNrOau2UgdNuFvA+a2Kqh+jPyJggvosyV0
E6ZzOS9GMKkxTRHvtvOJgqp6qoZWKl8/tsTN2NNWCb9K2PkRMDp8f/3JLIxQMHllHhxFUpANzFvu
HM6VFndtpzBzd3V7GmJihmTXxyzAaYmbeVcL/wW9KsA8Z8dIZLdw5yAbEIt6VAoCg5Cb/Zff/YuM
/K8SuRrxtYVDoItI9hFXClb+xlv7G/I5GNEbvcMH3e2ma3OsNIkOJ1lE5xwI7YKaJczMnlM/dG9/
ggf8NAAEz0bP/Xn26pzK3WRyl3e1yaaZ97S6UDmSPJphHHMCM0jMBTTMY3nL9rJhl3GSSsAf84RK
fg3bslOjVK79DOJBoGZen5qFMdT/+UYsIm7Lzm3OtlxydPEt6v1BX7aQU7nf9RQl4qBepssOJy6Y
od0eldR6q/Jx52x6p+0oOaDluGVn0ldRPHeUfaWQWZyKm9i9TDCqR1dB4ksiTPK+iQELhDb2vkC9
BgITZsZoBQ2loGpu5Dsh9AossKm4C69iFpZPo3xAYilSqdaHUK+SddYPWIQ4DUYz4C1hvIS5ro4Z
C08OKKpJ3SNCeYw2eT2slqyXoPNj9VwMHAwxaRU5VJkkfbl/w1MHwKItW8zsX5AZuSqBPOoRo62t
GnivCIL9VWOfy+051+TkVkVuc74wB9iCdyrHZepqVEQ7Fe5xF7m13yBmopwFEJTynfDJ/6V4DQra
5sfEAUDGb0XU0VCcs6S3fpL3+RJ3Rp1VLVZRoJsuyJqj+mTHBgK4IrtieyPjFyNeCqgXyApbQRuy
PYqn7Yrg9Xtkox6q0S2EYm3b8B7YgQSntbMLmITYtnRjuBXcBE7H5UsFl/nDYbglaA4gpOThCzJe
YQKVkqZ5rQMFZoSycRWka7ZiB/J6nA41cLlPH2J264bNkb0yRAGiMvfZgo/5E/GT5j7JSE1qQcPs
OKXorg9SXAFk5vUJrXnsfH+Z9rpitBKTNy22F4rq7Hek99bU6Z6Gq5siJP2XJ6TX8dGRwmY2yWci
aFR1W7P2dIWzcuPFqmTOe4b+dcUtwQcqlHPXqz3vomxg2/ENg1NtplXVkpEdveiYwDz+MWU6R9JF
OlY1vGTDGWtFLs4MQ3GwUEu9acZe6tun0oXx29IpX3fGiwh/QGHp3/Ia1UaltldGsXKSFZHQFT+e
Rq3wYR/OftAOAviCzrQPaUw6CWDkAxu/sP00tZ0gHyLcnrXYm9B6o4+06kDjbzIkbtVJuo8yGzNl
9DmHebdnsG3FbMsc3Qx7GZXGeMJ4IK6i+FwZKPbJFDRuiuqrQRUzOYUngjpF5CQIk62dEof1wev0
a3GnaSKHQhpdaFwyoOGJ1a9GSe1+y088IzEOKhfNpTnC80cNVtBkkHgRkwWPcwrA7Mzm9MPrfkBM
Fif5ktLtHaUdMphbZ5JiE2BNpHgbQWZXEy9nKHm454ooZ87lb6rqFDkjLF2IjKuDUpwy41k2QZ0n
nEGkN6/oC+qgvn6hdgIKtLrHdCXdqlZAGcA+jN/D2oQvWIh5kiwioqSr5gNl0AZjxfZT6l3dva8p
Tp455WZL9kqgyMu+xl7ysgC1DJYOo+Zhfpq+Quly1fX3JymjXQoHZWkkOE6WiYvNpv81njA6vN1g
SyoXGROIx7+V/AJ/ANl9NNnEwKFYbPH1/XbBXn7kGtHJ41avL8njFjCPMNS+K+/M6nEN5E4uRAVY
5zofopuVwRkKF2ex9STLrjiOgmClFYDruwzEjOJk3L4uIKdLUF0zLfqpuaHcHj+yW/ytZL+4WnIi
lF5B8TNXoWtyPKYB7G8spfXMdEEpy1TxlEdGbBEL5EjtaSG0XuI4cLGyFEIB6Qm8JF9/CKDVQSMI
b+hdVrvByP+Hh6kjuIWUHnozZ3FlrELoz4TiRy3rAJNJkVe9l+Ue5DntNLMcrrXyVugaYtXloIOW
7CF8GHcN/88BqK62/lhTVkiEuk9KaMHTvwdleh8cPr+nYLxh415Ek9lQAIVAiW6S6AgPBMe54Paq
Ehctql9XNPhESyw4HEaZLmmjTXe7/XanNS7/ItHuLlI3r3kzB83BK1nGia9lvV6kREbXcx/CJwgM
6DaMuhszwDWqMXBlDN1bs/Dwx6C8C7M9f0WPr8israSYlcOJp0plPparXLECZWKxpXN9k0TKMaLK
qUkVWK1HAg6bRPnooj7AgFXsF9eUzrbwOJSSKpwr9L6J5YwR6GMlzl4dMNNXkyGhTeYZ3F8nVX8u
GZfD9CqdV+YFLEjSdEEhpyuyYafM9dk5hJTbJlK5jVvluUURsGmh/Mon3DRepRBkhkw8UhTQ/hEv
vvhJWDVB1OpnYPCCPJ9iaMzrwSM8qg/4pPOJP3Xsci4fo2/xI96Qr0lYsWaBPFsSYo/TIMA7DuII
CJ6ug/QaQp5I143tWS+mRh8DWirWw8K00rpmgV3Uq5E/Ll/75C24P8A76idpvB/CRlR5nhvYxkvR
n1ATix0vXqvjkDnYaiCyfV1bWU5dccXDs3/W0O12E39CS1gAKeUp0MClRDi2nEwy3lP14G6H5mVI
g7/85st0wnNosevCV6NFxuxX9N76woJ6IJ6zO6ARRHLncc1QaOkSjmp9yk9meviFjOCvcfVM8876
88f6y9VqISkScTWaXGBSINLFwvovJg2EJt3SsD6WKN+CbAMWcZIN3xjuEEgRCUMbxxW2P6a/08S+
QCoX4WkBZr+mMrEktdw5vVB1e9UF/mNud1oYqds/KWst3wN6irFR17wpUSogos33YFTOQI0SeTNs
ullvlT/nwexkT/M/79Jlpe2txenKo0P/3mkL+rZNi86gBF2idYiBHoxNyke6cuDpDGgSpjHGrjLI
uz71QCqyZOaBry4LR/HwzaBeE+YWtSs/FCjT1pr1aDMsp2MZU9bQ+QNs3+Em40p39SWmcyXi8MY3
GVUojE/S+e8+sf8QtWrN8WrZqUtGpxAWPs7jMoi4pJkUfIHqkr3ne9rkzA/pERUyzKTYdakSvtZQ
d5Sm+xr3cXdPYpg1Wcy+Kpgr3rDzk4IhE/9HTLfdcz6VR0byDSKHnmJLNnQYtF1hUnDmlKFQPfFX
isg5oRfsXIdLtGEHfLxkuc3TWCljdazsbq5dGPQks5tS7chshGPKKk0a4awLybibaB7bLPw+MYnP
IVt4SAQJ/q09IJe4jHWdjLMkrsY+8TsaPuc8zXDTTQejgoCN8TC3jWGpX7b432c2ZBc+q6w1mx1B
1puxhWike1lo3bHtCif6KBO1R+jlRnzZe17ME+hQIDxhlT51wfEieu4/I9uLzKEf5sYIpjj/1vQY
1Q3XnidJb4nJgrjQu+vorxZa0uJY+mtMAw28spYl9/S4xAtEoWdR0Pk7FPU2YR0sTa3h8OzV9Xz7
fFhgr0f2rN+GLp63xJmk8QEgneNotCLnU62GayaURlgSAjlTvEJzfdfxZ3i6DxbB8PSZR3b7hr53
j+Xahti1HK18gkFcJjOoyikC61RFLKVkKp+Ypu1qNumJNdElO97ts5bho0h7aj6GmbU2Nw1cwbAE
GC9icI6qxy1pCmHVb1tLjYNJUc5s+HKFppXlR5KzaxwNhxzdhqylXVmRYTcHnY916G+QdxDXFyxJ
N5CjQUd1Xk9kF6hkfDnjhZUAehyz+OLEl98TGAYZ7JmGGNYK2rqrp6fjQIHigZ1ruf2xIhkhT27X
MNw8z8e4kEv2p+cC3qntZ7Nku7vRxTfBEnq0hDOVjrdA2qt0bF0Zuv8/B9xftnHdKT7XWEBP8apM
bsQbv9FoKH3oo6lNaKjrpkumx1Ik4cL4NpydDhYs1WzKw8+GhiqV++9fBCFCplfg7VefTrz/kr2D
IWZun7fMy/YinLe30McgamJflwgTHgk/WqBGlZ91r+HlXRDvMdymrmgVyATPAZPj5uT2FpjqlEUL
IJVT4+x93PJ4V96ZkXLgyaE/qH2s4Ct4PkM9Z+klhAu8yWI+IWltBU7xZd/+mSg7G0Xk8LPQWijg
h+HShwQSwEJNM26zr+rSydx47F22R12VH2qDYOWktzNC4Dm3masIdXDlluyubUURjbkuwNx3Vrmg
Yo0D+G5T8qQV949izm6aEsIdI3GWavrshkMukZSJ9UnTw1t7aYCP3AFxGWuRD/v6BhjhxobRxwcc
kP5yGhX5Ak5bzn4Yyfh2UnNp+3E3kAjtsx3abHBb1UwBFLbN8YlIQPZhj0sdDeEkjUPRZlgbuhR8
3pawDLYf4Bas8IYo+IS1ptGGD+lGzGMC/ATXFhw1vonPBJsl7pWe2txwzjD2T5rUhCxkzXqjqM4b
RcQjDHr5mNA7zxIVVu9L/75H8UVk5urReZC1+C/s64XEYmk3ln0K7ox5pEeGW7feDeRGaStWW3UO
GgPgBmCyN9Kpxgto6ZbEp/dnarns0+4rMFLgKGRsOG3kr9XZPSTuEBKFCU1/5sn9wuojQ8S4GX0C
Odb1Z1T003PNVnXUlRVHZCApYHtEF5pZP2Flzq1HoTLmWWYUfPX0LpbcGVQfhwS0nsMgnJzwSfdO
KUzZkXtCbZBO4wDW4PuO/IsHPS0KtmSt5K4L2cjcZCRSrRvIZNOm3le0kfgbVrNrH5H4/gyXbtjN
5YBfkyOO0Uv92XZAgBijZrJ2hMyVRldiuTjBasIsf7Ldx2qO5wKgCkHuoObVlQ6AYp56xNVb+6bg
kANcs2nW0CfC81jx4xP47oseceL1745dQfSuJLL3d9COyPS7SlNHHPlZEYQU0DQyefmZzVqkDe+z
BomvSJNHdkO4DkWzjBf5ESFOn59X02WKktzq2vuc2EK1KhuwnlcPVStCKerE+AqzQxJFy9q//TwY
EsGrM6h4TiDOQx4vjawZp8TA3EMOHcX+c8Xmhc7odQcbgzRoCGbg5IQqyd5DIMiKT/i5tiytG3Q6
nvhyo5jv8DvU3SiIaH4ukQNnuPkFb/o8lnGbsY0y5IlpVv02/cm/ofy1Wyw4L5W5mLJXtwJqhOS9
9+gemxDp95gjaVQ007EpCnhUHY2PCUddkpwPpQ/BEFriYSVJrpwVkYoWXM9LAvi9Nkr11c9v2rxp
qKsrTC0bLL9opL8rhE8dKezWwRypKbrGUioMQpF+ZZj04jJeeSNYlev06YouxPeNoNmJ8JEJBsJJ
GgHnDBmntPgAlyRuqyDipe2aN6M6nm95GJ30iwKjqZc3I3G3JJyKeaLdAxOm9/Kgxoc0TjNQnOom
XNUkJ5M9Js2h36Jc7wWwLylU2NCOaYSgxD8FV9CcFDxspkoKyuBAVMBlT8hdj8ukip+rXDrRh7mh
6AlbAgJX5le3APmTDxEwAlYmkc2zukDBOjD9pJ3vNsPo2679XeCd/0MuI/DqV1yehP7UFHqWOl1d
xVC6PdU/1yfEUrX57ZnFUD2ih1GFfBJWYmnnbvC1+lR9mkSvFjoEuic9Bo0QtYIaC0RCKpbAAeAJ
WtpSnxS/U1Ieg3klLZVtU86DGfcWHex8sB0hrL8RF6jSmxZD/mROZ0W6RN+/YDP7Ku0IruhZX82l
e0JeAZo5rZK5K05Y/sucTUuE5V7mlFy/ejM0+pAfyBU1W37AgXC2GYGhPoV+tcoLJhW3PC3Of4An
NWoor8pD7y/h7dIk62iwffIXNrhfPYtWn8T5r8TK955fhTsbEqGX+pbWI12xEgU/9bnGIDv3Mfuy
V7u4uQd6bHRlCx4P1ZwOAPZ9k5m00Gv6ZH50bUSe4hXr+SqfVfKgFtI8MXDqbciQ8Ls1+0lCyD7v
E8iMPnTb00V6cBQ7raAmtx5xP4MT+31giYEkkltu2WSbK8jOD70hEsZ0GHkuyIy+7YN9iRSHIsmK
S8sHFz+eN4BIJk5lHo3pBXSoOhAcFA+rwjmuDcQ7/qmXV6SxXZWwR4CmD4JWu4XOYDRJapYynqDz
76IvfEJjiAldyyfAU+ipHiTpoeI7iCLTvz9xP63zGO6WatEHvSI52Q2ItsltVZ+wiIzNUQgb1Ife
gkCsAcdB8/UEY9G/BSGHO2ZcsSRM9Zmno8XlYSMOFbshzYeGVGjemvBbon/t4ngtWAPQcOh4WSNR
bSma+4c708yDmC3+HhLfGD48jbks3frrdyeh5h/SiA3uCSkwYWjOm8QnPzzCw1ipxEAv9QuHFIbg
5wcDFJPM7W/uOEmgVRhEh5biztzi12H00PRwTq3uK6SoQLm4aQgpwGGt2drIv39euZoVza7TeUvx
4349GgbFp1vk2JesT0NQe1MSwV6JyX/Ppu45XOqr3JdmFzFdrUWunyDcoIEU0iVeJIsSiytvsk2a
gw3DjzOwjTnQvYigR9m7DyUXnHcNrhCYNornr74TAUiBWOmwbcxjicz3LIEVfQsvKX+AeBhwwOUF
GoRSwHs7G6WgcD0UdSbzcHKvXsW3T8R7E6InsRL5cQgQMCEelJqcT8DbwFmM9pld0J2+KP1f8rSc
HONHPpNrs0xn+XqLbymgPfZto+lrQeWvDMNeaK5lF/DlZn1ssm9C3TlnUlInE3e/eJy97Gg2WL8/
CoaI7kY+AwZE607NIUqe6Mpuf+7WwnYOV/imCtKbnneGD+2Hxj+SL3FnRlIFrl3STZKCxX2kg+2S
nuT3/MUooKWCk8yW3GKu5vWrrlp9FihyfZ9epF/QjVuAX6XE7+JJsmwOQNm86xhID3bFZtzyGRUG
e0rrRHJ/V3MRW1dCdT4fhr7ftX9D9DPY32n36VES9eySr2FBTeXdXs2aXXkKm/PhGDO6blpdjUu/
ajO6wN/JlPzGeDSYumQYyvx4Zp2uSHQSETBpC01uS7M8d2EAFn4s/4jNegy4HqZaiLYE/GvYQpln
P5gsT1hShKA6fsf5EYXMADt0pQe72I1ONq5MaRh6N33Z1PHGdWHYh01hOgXt6ea1Hg+NP+XsW7v+
sauzJ+6tOUts6JMZmMsDzesVp50edUoInilGvHuyk6pb/BTJM3HLnEYjG0xBZqP0/0J4G7jPLz+u
Qm1ccfQfEGegpjwzlj/tiYn1OLednN3a6vdjb3dGbBxNiZrarbt+47hwOCP8NrwboHavUquNTN7z
jbHA4sosxTkpGfrzsi6t4Ngy8q8IFOle47Z8DFWalOXripRePUzD4ZkgzQv5XExfKmzrfHRNr0eC
bb+4wG946yhcpFHC9tyZl+XJQ/gf5LpKQZ0sPGsJaPGrqEZcT4xQUMEBhwlTJVg063VTD8n1134U
PnQWq8x4+8R07SWfNxhuJoCyS9yqrecvWDMVUAzzier9pP9deWIXnrurJBbHOGi8R/70MbIJuR06
csrgHWu4zwIiuMN9KVbdNwBUta8r8mgz4/JOdKDkmRGt4p/H53WsHikDKPzeJGt3zIpnTPiUYeD6
OJ1KEepUDZYK2jV24SipZakdbykMquS//M/vbD9nNyH4ZPZoS1z+0Ui8Jl/9Q0PfbT+OsLw0hVnQ
5QgY+njax67M22jfsh/1Kj5g7PsTewINdP4pVRRRHg7WDHwZe4CsJd5F+9DVUuing217rgyW2k6v
ft6p8TDeeKsjtdvWOetZMNprTrwqEF2vf17Hrxc5VoEEsFEVnROfu5j2ICTMq7MZ4PND3xsVIAUY
8yIScwYK6QnVo9M11efGLpr6z4aJ+Pbvmox0zBqfzSEZrsDVM8OBoTzp7DqY7+XfULVevGOP4GHh
zeuFfpMU/z9q6jeAfauXonjlG2cmoOjXP5IKRls1LI3EkLA7zATMWk/dJqVPlxchkg2izaYvfB7W
mM18/AHJO3L7YoqGT9tu5GtwR3OCn9OcTwjj0zwwXLLpjnAPxDEtIvN0oKLW0jHrzOMXA1Q0Eccx
GvdhsY1JjzeletsIw7BWQ0uK9Cy3Rjt+PbaLRB+bGfbBk7E6G0Zugbceoh+1NVLM+bbUBfyb4X0f
/9EoXQAOBJf4jgrvH3lJzqZCNwgQdRfF0mR2BY9KTSW6dbnfrLX9w8uvosWizpVuOa5P1E3ZXwBQ
RfDzUv2vP2V5VTj692dYzCCKpQAEs20Hb9LibPTIAim2sbztxt8tdPrBM7QSdJLqcSgD7s4dRlVr
dJKzznwt+qtv2VGrVYfAPULFgj4eU4ILRJK5yYkPjnMEoMZ0bTtEVUKficCrmF5GvJVuDahDEwX7
ywRDeGv6ujLVWoJAhLa83rC2Oy4kBt+e3Fkndix64uhwWlJ3mPuAAJwWC3UVG3Kei7NbCYLfnmSw
EndMlyUHbvgvGat2vlBUJPY2EMnRZYRiB19LkmXJkYq2Xbwcd6+7TZ9nKwq22zrUuBH/ewwWwO++
DnhSsPZSUB8t6Dn5exjVCzT9W9eIYqAoXz8x8vZqLA1SQFw2Qk6Uv32bzEE8k0LcjVdVwsHsol12
YXH82a9ptRDNDueICsaPGyvwXDII9N/oKlZV+wfcRawVrVje0kibLjT39x2lbuwKnZMNBgDga5az
SPrxOr3iytTunuUNiNYHxP1xYsxaG1hKP6eCHUZors/PG4hatwodmDprEQdME76PFpdiRHGhUqbk
8/CVpu2I5+ssPc7U41Ze4EyH2NSqGHBWXUE14yD+/UiObiIxv4sXg/TsX/c57oU1EXi/eJ4nEPFL
tSQGeWHPacPZEGog2xYhVMCQxFo0aZo5Sk0fG06PXGm4TTDxOiXM5XLjvgHpMi0aNEptxFWcMh0B
aU1hCo04INtvHzG/f7nZpR0nFA5dx29TK6gqJdLn5KUv+P1FM9JcZLsdCiW0LAy2M2MHgDHWXQF0
z4lLFJ1108uYxcqf/lwt0cHA6UGmMQNEA76imd84qS63R5CzTIK/jcUzIbFLlfFWjbeTlLDi/ISZ
znc/TPf9pjA9SjhwHYHn8w/P62i+Csoxi2m9YML433PglL5dq4NuMQR9IGcilnEIUYYYd4MPSlCi
qjdieJ9hWUz9ipK8wgsujICLw+JADExWsRTo9na05Z85QVXBDy4BQs3XD+IWba/gkYR36El7mFmv
QTJNQswtyHXNxjHqSwlzzbg4v+DIjV31p51D+LkqcmCLnbv3OYA8QbppjwH6NURoILtlb8xaCdmd
XKVSdbXGdsAcsosZ6DCwQ9/wc1/4J/zeanG/EILbCBQOhRt1I3wChU0UFEZhpJdIpE9bgBzBJm42
01ooaj66508inh9ok/ix1VpTMfFe4pnNxjUs/HAar/ln4u+a//AH/FBhXaA7aPvFuleIOFDDneDF
KKR4gyQbtVp0e8OPe6ZXO6ff5DHMxAHo4PpQYyt7uv40IJ9Z4oWHSAmLsHHecDwiRElvZGVroxkX
8iuWnBqjvhFTpptyA3MTHM5ygYlOdIL/V2I6hi23q4ocGosSdkpVTd4YKqCZUBYZQI6h+nOtyFDA
oQNr9tdSdWxS2bNXjXBZUJes2Y65Ftc1VrvORoD21mTn+nEybXV5iuD2I+ZkJApLt/AScpgw7WnZ
mMcvnO09ogRMQq0ZFEGXKarrI0hiYIgFWpp67zSoTdwuPk/PCnDwzeLSp2G/Djmbx/RTmO6iA4qm
33ROkkeJi19iiloBnJa8Z+sXNQ5thoSUtioB4ym0cRwHVlAoULGJCfUO30CIvwwKgsqYGQzOZQmD
btTmKUg0CshaIcyxiWSegEC2PoXxtOOPPjIGnkdKKTFQMUMOfHzCSxJoQUP2jpE6qXxhePzRX8M2
9BtJALHDGZN/Bm9h1pSez4DF+W5FcP7cHNhg2Zv4iMT/AHpK4P2g8+MQXxT28c8FVclCzZSNybOL
mE7sfNHuZ0ZPj88trOKTmSlM2mB1038YNhAgD3f70p7HQTEa7N0rHgXjfEjL+syoWYR2XVBPsxDb
hSPkLcn0NNlIkeU/jBepFIUaT2IRdsxWNs03to/5emqr6n2GOEQaWoy8Oi8dasfgaauxEq49GsRQ
7/JLC3wRqfSvUQEomi7DUaddy0ig1z5eTBuYxNDthw+M/YnDc9Ukxqqlp8EXtsSMzO3zbLAvlIPW
c6SczTG/IMpeJ1JBai+P8s64dvW70NJ7y8CEot/wisrd2mj3XQhINTuECiga95W3YFIF5Xfvl0EP
UkeNUpc6PKK7eJy6qiko9u4blzkPeRaErZKadDE+i6DMMvj1hTC1S2e8rPAULKjZsrYjwbin4nej
n8lSJK/zpoasnqjmHqJs4Q3E9svoXqLjzGgEPutQhp6tA2Yexa3sJ6K8MASOTsFyBfEQuPso5fg+
EIQYaE8Q8a43HlAphnfD/F8hMf1qFBHWE/uNjFNqswCt4WyRE3igQWrNGHRhOea+/yVlQv8J8ve5
hhROn4ZuGkLpW5dvNRTluPGcR5szTfMBkuZQ47/NbiTyHA3fpZE2nMCMVqijbtj4jjqKR8wVGp59
yjl+4lOAtMF45Ka6hqAcY5qVKiCIgrGXzyDik6mJYSGOjqfqKRbMgeJKw0Dh8pXtHXLj9Ld5DTYA
mqkoW4Udd5FJ+0Cn8wq3WQCydEGbkc6cPWXFUrq5C9OEIH8P4JrQqJgDxoK4IkSyn3CsoeUR0QIS
+GzOG2H5s1zmt/tECMITf4w6gqTqjkGy8iwIwiMOb9MWhgP8cdTcJPhS3rs0qInMrCc4WgYL4L6j
pij1VqkXZHzGzuVCH/oonp5iIpkWviYQC/jHxlVhOgY4qWeRIQSgOXT5c9XQHe0qT27xM9ql8fTu
25u5RCnRKPTLIaguMYBy6WqF4EQtwNVEjphy2owNYHWix/R8qnIqa2mFwsLwQWbt1pKMpMDEg19l
egHYwCs+apZ6geGBOsQzDwXMywKv2ZC0LtkZ+0w6DjgPCWyna9NFMbF+FQweqUpG+wWOICuml+bX
PIywWKq8gVjYJmuUMCIZwotVZ9JThT5w+6i3tKX1R+6vkKSzYgupzY8dUdgv9A+gXGbk/kIaoFJC
9rvbnI+1EwMLGUfMtxTjr+eRkDUiTkv5D4iYSvSLdWNgfVuzf0uZrZfoLuDBqvAadmHGIfnXfXtK
6dSKYikwL/wRzjIl9853a1bFHv9d2RwuRd0p9vJsP3IzZ8iiDTn+0OGGLfI70G8/ELxDNnmo0glp
e0q+R4j3qYKpunhdcDy5DtX3S9JSsoCWtPevgdFFt/7Qs+YEOH4+62pB9OTg1aQ6+kD4OphgAFJv
x9EOkvJeMA7CfoRe98wTtZEdr6Ikodxuq5Xi+7vkCCeFChgATU3rn/YFfdollLKAFep+meAAEIFk
DySEgnqwp4K+4FFwRNQEZafw7BdpxWLohQi5tD0CsuR+jBqgmlnEwzP4orNFaGFL5Y7HtzM37165
TU1zZH+w1zTps3VkPox5sg/S77EVU563NsScNHVuwf4GE7pQDluOgNF/SCdryI1W5pNR+s+Du4Nw
4M6atllcRCCqQ8L00klqX3tJZTYThJ2koQFXzaeSROYLUFdJuEj9LJhi/Wmj/SLYx7nVOZbNvMx4
6QBrSzk76vBkmIf2rzqGGawsK8sBVUZrzPfSKPJo/JOs8bjgKABWjY6LbtVM86x4yseSmrJH2y7P
kseHqzMst4UYohiKF3br6PYAVJ4KbtLdDzmQnEJgcX2xmBFvi9+Y8KgM1YNqEpaisV9VfIVXRDy7
aO4Qd0iu0FKm5yLG4VQxdu/hnmLPwlHo7s8O/re/I080xrQkhNW9SRt3XB+5lFmw6iAcVEO53z5T
Xrrl4ebYSlgfGqYV9kqOpdcM7ppYm7pbvSGmlyoJyGUlTmBivVw9z0wuFl/z9p6+LzG/4Jeg/eQn
RKyu4StOwewobhnwJrkiQVYLKPKve+90OCFtcbhC5FHHQVJEWQ4TA8sXXJxY5Ovsvch8t55QEtvp
JFkaG3PTWnZRNWjz7FUP9M3ExWLG0CDmMrJchI9HgK0Ijqt/tJVThPO6JndZlzzi3aH+GOb1oSwe
qqVYc0bmJDKWzNs+Tw/p+5QKzXeHIhg6vs8D8KWs5UnxKN0bOg6EvtpBzHEcN6Usex/L4DzVP0kX
wRU9Eh5urLrpfhoHiJGP0vhw0p01hlI0uElfugMEeXY0XGZ6pTXxj/kuy+fUXuxTr20tY5ru+0OR
NhqxyIJTH6FA5eNb8DBCdPAFXCymGwdHNXb0bLNwxDZDCH50Z5l1Z2431OnOWW1jG1u4vPA/8qT2
+NHIjoW/syUtHhSlisRz462376RalC+/SuXNB4BEzqspDQYqgzNOmSq71VEaJiO30lXbw/b0zftU
B9n4fXDIdIUkjKq9nMPj3J2rAg2h28hlWAZh/4uPv6Xsid//KgOrwA6wFF4EvTN5B2oLgq37UX27
zlsJmHn1Bqr2461QcEMn/DyBWuWdNDYcJdaQv6luIDA6qyUswglslLVUHdJ0Uey30IMrcKnVvrrg
aVIDkzPaFN2vgQAGGYh/3I13HGEhZKGLrV4rFWTlMTzZQvfVsDAvkyIztGNfdNziHQKMD1L66+y8
gQB6o6A6/u7DRr+/zXCejRZSLBXgBAyZBgaQdXICHCT+IY+tewH+CGKwuitMX6CsRUgkxMamVdQO
a0BXYidQoAZIbj7ZGtOv0JVzCEuwFzFvjYvfsBnS/WghkQTVmLYjilInnrMPonBThN3VyFrmZkyg
EAJFMzgbugxoJn2t3/dQnM9dUWmx1ZUwm+C22k/OQWkcgtLGUJUIz869N/pu/USipXDi4wnW5IhQ
NttbTbF1tl7EORlF4h06tJfUAGJlTTh8EJlfh/DE5qdfI2Af2uswTJJmdQjHVNWNvdLyyjud2XVc
0k/ZhSXCpVy1WoQqwjwx9BvhKqLpJQsA28qU1F4PxnO6APXDdeY3jGY8QEwB++hE1gtNy3eU8MgW
EPb0m2WvJhp0ctxg6kgE1LH4tf6iQjQ1fT6uA3TNcr0PzbESlyZBkvxfLITP93G/O4A1qvQ0/Dv7
FJn+TuE7GktXKtPRUXCQx5Pp9mywZzJsCaIbAkKT5rXpg3+T9DGJwQ9YNnwa+MeRHJK0I3nW6Tvj
6XYRRbNvqc4LSZETJ48u60TUfxevIqhaIiA8FleZ+Es3fJc9DLl1Zzvz1t8c7IkDmoSBp0aYMciE
Rx+e6ij3opxh3GQSP0BOZ+yesEqDNjPN/8S00eOwh014iKxfBQVUfmx14gbqna/Q4tghJHxNEwPO
Uv0Z6T4BGZaut5z6OkV+pep8apP0DJfMdN6dBpTgn5N5o83+xAp+m0Z6z9WkuQmFy2YhgYp4Uk9N
+5KN1mZkLl1/Ijjqu+6JAgv/M60M2jCLdjcRoMJTxblBXXOkId2PflSzb9G/7uJoKqoMZ9OGA8pB
3dGOW2H8zU+xWDY5xsh5DkMkDNZgO0NrgNeVaqRJRVqH4jUFj6eNb/cXo2bLwGdK73FBvA8Kbrm6
7+UgDRxD734KqTIkictvO3mGmqOxU39M9TeqkhYLq7cvu1TlQyjT80rIpL/kkY5uNmivXUUD9srb
75PmiQqaNL8Oeazz3EyZEjy481RHwk+4yvc8sFL8y69MgzULiDIEdVZmQuAfUdidWMp7IXe7ZVkk
rCI+3hXUv4RMJ7GjoEy3TBjC+n9LMlZO567Yw2liAnXYO0bPfOrohS4lIUMisK8BnnLXJleFfwrO
uo+D5eOWZRn8egwgsL+xxaffTcAPQHdz1NEQnKC5XRhsmBu7J5dOSa8giMLReuk4dHkZo+vP6Smu
pAmwnWnG79h/V32ijqOnhj4Kl0x8f61pKVv2GBmwPGRYdzrzzb9ZaWFgeXQXdKzMxGkmukQmXOaH
3TXnEVY0LQqgWhfxSM3z/4a3LtbIZuSLisfqRkbU8oDob+LHDKtwaSHmZGidCkiIJ+8SveY23+Bg
6kHhXfQZn7i92vGWsfMJHImUW2ZMLJPE+mobYCKH17+aK5iQfzw0xVm0EK1ZFFw6yCUXLxXmnP+0
R6LtSnENY0WJWMz+wVFpZS8CJPUcId31LqfBaxNGV6D4XRbpd4ikSnlZDoQe3P0vgnS/ZiZyvO9x
DN3+4Lg3gjUr8p1oi3tdM/oyjI/NwJv6vw18ncPLqhYXfMN/fYKKlsOBGSVYppAWlpge8RTSox7q
xIXCXSMnb6u5WeFab7UFJJzbY25Km8vUIeA0TDFYWOTUNooocr2jd52u5tQBzkKc/X7ujBMIYxM+
+tK/+3/ZBbxN0lmut/rd/XJ6vWovDUBndxTqvR9pSyxgJIBDXnyBMD7RhkfDLsyxQuf19yqwJaPE
7nZOL3GDxwgA78LJE1z9ipvPBSbbmzK6b+ZFChvECX4jUkf0Wylq0GqBcJbTpFIJ1dUx9uaMJlWz
PAYdbu6XVZneAtOD8r5jmhUJp8tfg86F29PVxWkTlxT5ycIEE/m1VNTQ+nXkIxok4HLpsJBfuzvw
Rqk4i2P9GJ5jW+BzJLS89hBOOd+/yItsp+W0/1Cna/dSXCwJh6pF9TZoNYCBpvQF55VIos7ODxFf
aPEPyfEuCDySPWTrJa4rDJG4jY2CMPmwgD5jURAgRVwQIB+BA3/uO8yp25zLPsd3LLXreQewNUBr
PucOp6/c/QAiwMNaT/6oAm5xJU+jFmaNPgg7liOi8FXq/lypzlMI3mWp7lUTR+nS10XybxOZdR6x
CQGKn3uh1BBvBGhF6bIIEdJSlcV921FkigYVFtZIB4Wl11Hrfwq3Yy9Exmf6RGJRgmViktP4KeZx
C6GPXW0Iq2IONn8WL3kYT/Efx5AWX8JX0HMLAqaq0YTtVo05YyAQHpvmzXWNP6nlRRIP6bzurneo
W3GRtfXNImwe6y+68tVyNayMz8/yXDqOxkuMH37fKzEcxpI9tAxpbpiT6/IhOSFCiFcoTrg6t8xa
LnoNp/fEZyUlwHP1+xIJIlYbAQhCy3/WIBSnpwu54HkOgM3lSsMAE2TiXiIJLj1XtewzcpEL5aAl
4TTrJ6Uq/YvrjYIgEjkVXrpeFv5/czk7V8a3v2K6rGaqfwB3oHsiDCnXgUeumtnjuUSdrStEZ2MM
r5eCLTh56Fjy2l3MewR/NWCH3U2sbNsiOhm3nT5n7fiF1nM+SNV9Bl3fyekISUH2CI7OaBFdRgPN
ugFTKpGbD6zBDM+SE+hidchldprJGBvjoIKZobofNOCOCSWgvMoOI4jyQJG/jJUNSC3scww+XgxH
DdawuqaIs9H1YZwcxII9R18AnthabNzl40Axyn+cFG5EZTWvXwEbdQgzqMvwk35PDcIXEKx+cgTg
YkE4NRISIEN1aCKhRyfjsgexuZIOqhLmJP8lQO9UmATuwn4dB8cSbbIEhmMYEnHWtlt83xsD0ZLk
np4AzxiTu5fZmNDaR2lmt3Kkt/T2oh0S2EDjIoAh+5hniAbNnRWARz5NmeaRfb7W2m7nBrwJhYmf
4Qj7JiCYVEt+t6ctTfqqBVcQcXKRyjnrMUul8XrrGZ4e840ZuLche/T2MoDb9PocDyDqOuuXXPig
Rk5Cq1gfd8ujIpQUJsdAq/viGdAw3jpZcrmqCzVytLQsEovs0J4pBKtiY+PED13WIpvR1a/lxPt7
jxhZKM40betqvonichnmg2+QJ8F+V8EayhAHjmkmTVlZ0Tu0ykAGB7tY263cicmfefB5V+5coaqs
rKi/w1rVnQBzyf991xAjjXFl878yBvVa5BhPaescfoUEuIsLQAbMMRBh4EQAfOCu2NP/HcRZ0VNu
v5OYF19+Y1j6WFfQkqt1G8UDN9TGQWQdRP3NdBQeN+Eom2sc79eWyduaA6za8e+2fwUDr87msctl
P/PrMZlTyYOauKxDA9RKt3EQHe9F9s1sNmMPbzoLffvC6WiUKcjdNYQRLAEoSjlninN3S2jhH79v
9ycJuOLhs8kFF2EwQpdq20p4vWtg+y0qVnd3swHXAYSpPmct9ApuE7CFCwGgy8Eu29vt1yeoNMq+
b8zns5MwOrh61JWaM8oz4BdU2jpmI+py4Hb/m6S9J0ELhX8jl5ib57CwPNCBGASj9dl9qlzHnhyC
x4TfMvjwKEsTPuh/wCYbO8gQdo+VHRw+ZOPIfUiAJN0ynLq1gX0HSO7HErMFD/4E1yEJ6RbSIjpF
8SCFpR7SJ9+AqjfXdS1oBkfxiQ7UByYkM4QoHsOtnOSveGZGou9ni2uU5C51Y46UXHDn7dMDGfMc
FbC/YLW/z261U/n9f6B0Wry8uHFMe4RWB1CZ8r44A68Y/SASohAgV44onvaL1VUuhYCXBTyE0F11
s5fxJ8euFFuFAYtDLy3u5/p6weTF23HbL97YJZEj6EKaBi83bgqJRfMBe3+whGnDKQs5fAh3aXUb
sCnb/CYgELYZTLSv32Ci4EFkaHbNLB15FLGiEiDcmnxs9A1840ptIHjzTxnAaetcT6gX7baK1fRk
x+DM6AFkKwBBRba6pK16YvyOtEqpl0egLCn9kZmTCxMEX2oWO1sugFpuIZKpURGhlVp5t1/7F611
8z1Nq04UU8eR32jsLaJmIcK5yAKg5o94m0clH7uFBJIJATgRfl6p8nCpXYNw+7ZvfQQ6C5mT8CDq
RnHZAqFpp3H+OeW2YVhmY/skJRAtOF/MtXu5+rjo9zs8uIZTiB0oFKbbiRN1R2tcr7kquWwI+wMs
er1LnQ0gHhrdV8ZkYQIZ4Z9AyafRBye9Nzgh6cM87hI6p4Wty0b7d9yYbmMNgSxE9Ulk7UenQE65
lKfDhIVw8vbsXB2ZJXwpLSkw5Nlrg5ZQ0N2ifGoxji6ooP02tP6q+hGkqcMt+8WdPU8zCFOCIShz
zSK7vAnHGN8olnOjRqHA7qAV9lRHhV5AUuslU4UaT2bSnhlGIdknFgJRkePfQEqpnbyTwNziKLB9
Pp1nUJZAYpaKzq6r2/3PARhPykaeLLpvgZEMP3PURfYgcoksQsTsV2jXk88jZui+AfVEivwqdTNF
kOfnnPZEgU1jgZ7tEpvUPs28f2ysH6ODNWuOlRmtI2R3oKir8cdeHU7/lzHUGbXUUYnxQK3+hXTb
X3fUR4cfmGu0Bxx1W5Mhmp4Tfyb6tnzNcYAuOYLnYgKQZkuv71Z3dgS5SDA49LdnTna+NTXR/E0l
axsz97qT59oJUZgU7KnnEZPfFmXi8hA2o9tsUjUnoHcWsOCXr3fXykYq6J8Rt8Uasn33Kebu4PDf
yCqiTpQ2tAiU1xO8HNzENZPtteZfSeGCNbxryXiyYmf5aJ3miR+JnrW1iUGavQdzpr7Stg/qhRqB
SkvgIY29Fa8ANzmPQNgpT+dclqg//yEgTj+PJvR1/JDctYgQY+CKaJZ5PdHBqr1e0OQCO3geBW7e
qtX+UPp7dBQpIQr+biuLalBJ2eB8Ewz2B7beUxFatG9oOZiAeAq5+tXE9J2v7peFeXbXbEsHXNvp
TZ2F5uz7RO/awUuEFDpHQ/6Hirxh+gCKJsNdl4jfwG38XO6WbAyYQ7aEU6hLfmZwrubc3r/qTEM8
1MDPIbbaXbBcaixkYjn87d2+JYfAg5uJ6RP0dks7bHus+kq9UyXxgA9U6Z0p+qHCgbQd6+cIF6JM
T/2ApGwd2E40Wauzcbtk39lZ9qUc0cn2ARD4WwHyadMKfpeLqixQSoE8ed6mg+mo41k0BoBYKQZU
fkLU0bL8La5r8AP0IikwT971Un3C5jtsakjT/rhusFIjv6rWkUF/8aTmB7VyM1NnUxzmselHfY4M
7myz1yfgjEKsCH2jsMBLr3v+MSm2hqm3xqJnmTCD4P3PtvoMp4KwpmdlH/VUIxySHcw7ET2p2zva
TIsIcjv0ma0iD+l+Nn5MSOMgZJCLG4F4qendDGQUJvPWhASTKbvsuPGNLl5lMdSlGPNX64mZ7Fub
sjw6SJDrS8aYB954//rUsThHz35talWU2xoBpS9n9JWQ9HMWdjGWvaBHUx9N8iuevzHB6284EC9x
A/iTakexhX0T1Gcn7Ac+++c5NNj7FtEutAcV4hTxjbDMl4xivSJfdMaZMTpKE1u7v+CzOLTeiZ5Q
CIiC5WkGm1XK+0NFKoCCYwTtx0vQ/cfdejPXQ2KlsP3YQuHGa+oc8d8HHBg1/XyVU7ITHe/EEN86
NoQ3VydOKU+LV1AU+INUNckscmgIfSj2xiiyreSOiJOLHeq/8mIcrNhk4kIDUpwRbFAGsMwicjbw
jG3Z+9Mc/KvheHDjXLtG5qGxDG7T/vE8qqYpq+aegf4LRPk/Rlk89GttU6U/7ieyFuHU4F03yKLq
3kavMyBlKhy9w3yKju22aDY/HtaB2UzIaLfTe77T/Ns1Y1xwxU9zLEgK/4iQz+Jg68jjXr4eKxI1
NJmeZg7P84meKoSixwFvd6Ojr5QH947dd+6O670yIGV8j3+dCN/zx6NTHIodtxh94tcP+rH62Oa3
rd3cHp7ChwM6aB6Oxaq05GR1W44iftYYfEO15fLnCvMdqNLKOsJ/KfrmKV9zyQreqqe7GvZmgLN+
OI6bC5hAV6qdEubNJTYd/9xBP0vYNTnNSP2bgMs0uaVhvEGUZq1Wq3bfnAic98bVwmvpmF9OrHiZ
y+ZNjrANs9M+dLHHrU3EJI4mgEk+OS687i8v9RAxwR750gWinBdUYmqstr3eHE3Dr+L5so4id8bg
HVvelsaRCFnYvIzINAcmEH9spM6F9wXr/wpFhm5n3XBKrepo2D2ovW6Ks3lePBlwEoNNCy2gSQoE
/JzZdM3XVqu8ZeNYaZBmACvVSpxTX9LOqFpWsl/Nf4BMYS5obecV0mxkyCc4JmUo4eXJOjXF64nS
JLLc6s4ejwJKi2m4jLrqpnbFbvzbfZBzELFuY44SL3JgObsWmkYoPiOnn0lyIxI4hQlU5TdgsEbz
F853DZy+i7kruJzraJKw7JIbx1hOS6RwSu0bZ0ZMEmdlY9LIcZd66nS63IVKEITiJopYDPXvSAYt
HQ51AROljCATeLodFTS6KWNwTsVLmx3JywNt47OlPYqjENYorvWui9z4uuQd5+iRfNA+Df2fHR2f
Dl4GJjM3FdRqBOVc4zMlsBmgTlSWgiCvEMz3bcZ1IZJTXAy2LPogFodnmh8AALklpLO1sPhMmLC9
9IJukCMaWhQ3w3akh2Ws0I+RC9kUDbPn4uqfCkfoVr1O3R7FWTHxFZ+Ja4QcrGi2lrh6XRX2HrJF
AgSQowGMRSHjZV09rPKzjfiSD3qtub/DIiRzatzZp17Qco2lIZuT3ZuTxtsob9LGTDiIdY1H+NkN
tyVquBgGedbRfaro7S+6FBQ/3RhFqs7naiRssDsW4PJUG/ihEdRcc+Q1VNf71Ss9eVx4iJrb0zl0
5wC/to5DncazqpXpJW8sbnvESv2AG3QPWjrbg2N+Hn2DaCzpfHZSV/nKl9L2dmnQHnJx0E2ZNYAy
MPJHnEYYLSfTbJI4sJqamInscI2+25FfAUfYWrM/YGqEwQ7uVVI/miSkqkvDek/Kyl69qHsxcjlk
vGBXMATszoau0CDt2/etwgN33pHoLKeluaaVUnfZ+V+bUUesuzT9anL0nUiR9TBwYrSYNizc1nkQ
ZpCEzdx61rYKU9KoHPbSz73swYZvEU7D6ANuiwyK4bkBdiSZkPmUQ8a5DOKAPtKXCk9TNt/M2Qdm
wtkvqyU2gxVki8018D7QdLjmlEU4c1Ac9V8rtLSt8ru2foqTpvrnNGwn0ZsLOtBh4q5nQweLAH1p
UkMrQpNI64obImIUWtprY3G+NBr5KXg9DHwFEyqs7des5EoZlPs4jOoC2GaLs9em7bMsvQU+lHOF
jLU+mXbeHBhFGWCxJe8juKQbHy2Q012wmn+wbYBjYA7fCEW19FY88AeI2X4Bo3Ly6fTbgdYAGtnY
GZexDc1ab9U9cmS1wvwl/iItT607NIHkWiLAoozbCwx3GNBRAhE2nCJE6T5irj4NLrYAGOmRYScH
L2eZbCI7lz70KQk1v1MAp0u/AP4BeKM34BoWBtnHSZzwpMuz7m3fXBntxb91RfPu97MjiAxEQkkz
6UhbTOPiGD1wOuEE6G4XczWFQ+66L2uOn3p5yXboG5siyQAziohzVTiKKon/ZklT59B2y+zonz17
7PVCEfLWJPcQuk9XVMekCn46V2MHiKAAIbV+trq4VA+YZNa9goiV6mMhfOvY9rHJAXjlzhNojUfM
SY7avzIKWUjaDSJYfhWBRkFb3mmXZEN2zx25ymjlC9s2w4ONrwuoZdSR3ng3geUAybx+281BkWFB
rkkYRBaLbyAMKNSDJgYQOtv548RpAmAB4bbVOMgy4sBttEPiSDweeZu6EOfzyv+sqaNm68Ys6XQF
Ij2PFFBZZPRodQkrpuO1t1msn7chiK8H6+CW00uFGIRut2TNrGJd7jZMQ3c5nniUuuK8A77TMRpi
cUMchuQzJcX2cPX6UU76JdIYn9nKCCHOHo+5GEscylmZiHBeNSNPXAwxz5B+Nge+N5pBqdWPFHRq
DbxTeYnYOWcYGH2mrHW5doFUwSSGTOqfnC7RhM19b//EZMv7QGCyCUjJN9GlrGsz6EMF4Wu66PAz
mE2l/55shZtda/NjwdUfKQn9v7qkTht07rpdy/oAjdS5V5izh/Npa/QPgH7NieMypsJcT15wzitM
YjK4E8FqKhN/a3UOoSJyM3wsFxALuPg/hhwyKaluRZ5vLPFaDNcR1HtaJf/ymfYknlp9IDS5UqfS
VxlaKnl5Nh7lp/93PBBOt6g61z6wcnhv5yKGYWPiCrvF3k2tVOp954qbrx/f02Aevey1sKBNtfjc
xj/JJSzOMTRTm5R1r69EvuvbGefn0gUH61EKrt8OKHnlLmC0x3vvilr2UCQovUS3s9pKa1XG9ys1
SdHcHssSYgi1C0pUSEviRs6ZgiuIajRTYin4xmT+fGSfhgBGs0oZqGcrmH9M0r3mNc/DIwnHbmVj
N7D9lKv0XmQtkZjJY79YlzwWMHaMkmSqwqnQlHLMaQ7ZAkA5LZaQTXyAESsPBzcH8dmlfzyyxvGO
SnHyq7/EX55M4c2TcUiyiWBpak4pvlfdwwSawd5YRi0Hfs0FPDeMKaxCC8sYdqjVlhSK7O1FoQp+
Zky3mnZgQ4JPZIbO7m3ISdARXti5s+vPWiGqpk+bM/NblNliBlK0byW3DZZurXsgCpQA3mZ+9vGy
IwhfDW16heAiIznQ0vc2O7CvQDaHyc9zYLOGXSZtHpvaNdsTAwqFgpWIXzIIGfUOGB3s1dQa0I0R
go6Zn1xYLJavps5JmeRF9+wenA3A5iZ6YAhAQ7O19bcarFif4ldTcSQpoFeAr/O1BrCTVjRELIqB
MmFOWPDHng0g/kODMRaui4QHQByWZwvUWNyjA8+5MgD0on8gm4p/dPv2fbuoW53otmuGnM807neh
L1oUISutjizXkTyZmIibn4qmcNSJkqErZuqjCuZ6i+aIK2siV7tyovngWWhTcLYt9+7BauxLz4f/
ZNoSuPxUeuM3YehCLRu09lbwmvpLn+E0Ac5Uj/Ls8j4hFa7UrJg+LSZozO777PnrJn9xfst2JpQR
tNg2F2imup397aeveHySBGI3lDhdVaQDKCYCpq/VV6mxaF+tA1ZaD/ZrbvcbfFV8MIgx9A3ZbWp1
CyYBISPO1UqyoE3h8RrJKttJ5hCf51y/17WjlotPNR+6T4b0vUWUoS3stqkJet7Qx6pBUybComhH
azfFVzj8Az/XbuGZH4fjK0iJ9Rlf1QfJM5CvA6HYC1Yu+WStRxsc6ztIdCVVlv5/eS8y230c/pO1
ygZ8OC67lY5zQUiWDLo4i4Ue6sobMQmdCgC5ucNZx1nGVAy0cUKoz9On2uLnCOb+UYcC+F9usQ6m
kiNiKNYcvn+Xs1o/ZEtUOhvlxBq7cT7YP6Difvea/N3sxIoRbtt7pmXd8/gGOGohBvMJyN4X5bVF
VgxKDPT+4R+xcjWtOuncth4jxpqIfVDVA6O5aSiPPMqS/djk0AfkqQZLueA1e5QLkU3jRzwrY0rY
u4RxQGhjSM3aQIJm+YOO5HKsFs06diEctTd0hxPtO1AJzsPG3XbM/qdzZ5351Mj+iwZxgJZsb5DC
SN/8fspkzljxOPuT2B08Pn7cGXO4AaY4TXU5S5grzbQEIi70JkrtnAISI21V+QFQYblFGbvt6ELt
1ZHmOZswVWkvudrnKdyTSOOZd1F2b5afSqqhauIU1SzOpe8U+3Moqpr+0+luTyklWZB+gQ91OJm7
XygpjElI+LUCqBhdqT37qX8+fPS32KHc9P6gNWHq1+89jt3KJiAyHpo6xZGD8XavJo3L536v8QiD
mmjbZdCVZ1R2Gu/gjO2+Zu4qp2OXj8q7KRSQ/RnDNWG+m2RU3MlvQN5Ygjg0nAr9CGt+HWPtnzlw
1NO/l4nlH5KXQ0JjkQ69AeUnDMVuTsHkM7fv57YmlaqE2hDshD6lmUEUouuMt95GhcNk2g888los
PRYe1oC8cCW+pQBmnXSKMUZUIJ3VtlKRkekAz7IPvWDI6B8i+XpBchh0dwmBIP6RlzZsbRxui6BW
PEZCEvxdZjH7c6GjzXe4H0oM5a+syhajhd0oUiolgmUu4pDYayHqLorKd6CzOuw+yoIvmtQt4SgL
CjhK3TfcGgY8KvruoFzmL64W9utdmlTwbhUT0SVV2++fg3zQTHwVBY6/8GlKbaGoh3TY1aIlYA3o
DgMBysmcDpaA5Ebxu88dzWLEj5ZshwmjPqIaaybbF5JqUOLawOUXZ50slkYF2b/xAdhgpoofg9vN
iRvDd4DmqeCE0mlz8iXuvMHs2JRhLhDU8Ue1qmH+JP7bzSSkW81vRlgis8KJX0wnQ8pwzIfKUSXf
I2OUimMwoSNEGHzFU0C+tBQCgQgCLz7J2v7yEouDTyVLo2R1DV5trzHQvKGoFI4I0mtgQZM/swy8
DNOWe9L2x+TrBUmp1d4jzI3rIJXOccjaMviy0Q+s7wQDGHsZUtK7/+NYULuNzdZ3K4qui7yoc02G
Ul5ZXSrWeaxGXcDLG+/9Fc8KE0iJnZ5MIeEMo62lOT+/5Y9DTAz/q+qDIE/qFyyM8mYjQu9b+jpY
yHgvIauEbrWigaDXvfHOWHJsgR8gOIai3tOXb5218szqAgZ7nyS+Fa2ieEZKcidTurcu7VuUP4Bx
gwlDoxblumaKyBcH6QO5sMc071UXKsihNS7XKf2VY7U5hJEUl3blGEXaIgHRN48bQvTP6N46MrhL
necEx0+YwH/XsUmUlE6NYnB50Sa8deVYn8R6TKC+8K8xBU1kfOKxYot7hCTmu6UrThTK+Nxy2kRL
wiZH16ujeK1um+k4cMJmcIkn7OtCYzbTCgBuZbw+5sJgdRgjXMcFPkuA2DbHbKb3YU4qcvdR1tD8
X8PsipYIR7Ph7wps2EFQUHvxntfZmKAlJuSJzVzMNdcqv1REok6MB1FElagsTogOfJu8CKpAxJk0
YRT9oP3ixzCNWw6O4Hue0mdSMdwBMOvGdlPUZYt8mSPbgqEaCoiQRMHZIN/qNyt3HoAKp3mHzEaQ
VvBAB/OeZe0t1rMEsYGK2z68hlA9lNFoXPC4NsX7+trA9gs34MdrqaFJCUoht7TDuZdq/CZK4aFr
53eIfhhFz9TyNW6EtwNgRRCjG1RUizVYdCr/ywjGNiSQlllPWyD+iA0q3PXtmroUave3WyZsunkY
kzWfccEP2uE5Eedd/AmbqPuE8r1k/PzdAYZ34PQ/u9wnVXzpziG8MCZs3H4cF+V3ji+Wc/19OPpG
oEJ+cYO4sWDCPbVWHiqvUba0zZvbpBH9fZpxK6sR6TDBwpdrBUHVUmBi9rwLVD2CDnL8+ltvF9Ng
pIal5/nN9CG0OpKb4Le6VAtp81SFPxbzbbVb7iEBR0mpEigWW/J1IiuSXVh86XswTBHXM8JTDqvc
OT5LlGiJdqKu7gbaeC/8U+6SwOfJC3s2Nz4BW/v1Uz+8qd6ECUL7AWYTngJFIM/mLdK8fmKZ5pts
mMIGAFIg2J/t2eJ8GqlXIUna9PVrIzaisbnp4VXBBO9X7NsTTugFWS8mJ2GNwCPtwcM8zhkXwKGe
fY0S2lvYkjYKhoe9arJO9Za4oDUfihWmmqzy/O1h17avI07Gf/x3efBYnDzXUZiAYNPdccrtoDSR
Z8XLFuVABf3pmsRqnOyaTO3rUSRyw8k+cVWB9VJjGBf54mTuJj7wVVGyDh59X2FOYezqv91QtHeW
22yQGHA261gHv+i85QWbBWWcCiXE8we3GeN+il446+dCWAMgkUD8B0uv0UHBctHe/wCSzOOlTO07
O7c9BDIqoYHLMEyTP3rRMJZ23PHuCGIei8DxN8bTUe9aPl3R+hL9ratws/WlBffB/mvnL6j8Mmus
S5tSzOd6Q9MUJON6st7GLdYnOgt7+zWYga6sUrfQATz8y6T7PK6VVry0sfhG40F57ZiJVN8xzR/5
P/RSN1bB9ao6EVbieZv9lOZ2v9CZihqNuUi3wZrsASAvt3Z4M2DxCZbIG7AZLt7a/oJDOEwkkgJy
cB3HdeWA5uxCvkIejx94iYNzW9rF//CXwzzoRYp2MdsTq66XSdCnKCdnLlTgqF61t6RU5votifA1
hxI+gmHPRKezyfk3MLbFIPELCRmObGO9ZA6CJMFRwaVuTKjwKHBem0BsYk0oWz1u6ZQWeu+kl6nC
PdPBWG1kDIYo3QT8m7Awxq2oHtaeFKUX1jO22ESd8he7BFs3X+qCr5VoDtiT83QP+sNRM8b469v+
TBBXKQVG3p3FAiB6zdp6DN+0Gp1Rd74i3FgS7t8jLX8lxRNONRLqK1xwhZxwrmcI/RQ9SSW1YJKq
mSthNvMEJLvk4iWRZrkv4QDY6qO31HuDWSZYDr4t7zcA7PzmasGJ2EarrmCpBT3gZm9yH3TmVX8X
aSplPOatHRpcUEYrEDCuMrEbumfunS2xwIcXfg+DowaaeJfIAUVrAkmVdToHD5WYNRnVb+YCAY0w
OlAw3iEELzgiFZmy6ysnx4AToRI8SRHS8sOVMTHAIstnM8WIrDFlHtUv+/fOSV+PZKiYtF2Bychl
qUSgwX77lathgGKqclyWkm5m8xzm+bhJdJMGwCHVPVCINhvNpqh7dkY/5ciyOVIjL2w5efQg3yLe
oVsEqTMbvXO4hjcibpONh0CW7vFiSuiVrJxDBv0STQB/A5o+MY63jqwem/QR1sERbmgGNjC0xgoA
D7LfsztHowyaxG3XxppCxL5rRUDbFEH+lUTXKXQF33TQgJVAYjSCuSQL5d/pRCLWXyUAMUV+uYlT
MSLEdDTAahAaGX8gyji+11EKqOUb7DHvmP9ytGGXFVdTuRN9+Fc7gAW6JBShVSvKiPqEYhLAKhXP
Zw4K57EZEGn1bx881uQ/wEnvmtdk5MQT/KLVntRFq3b2oasyPc7qiCPsLhqbjMLwn3tt/14rnUfv
BbgQnce/1w+pLaiKqbqKpyBBhUP0I6tGIyIeWElKej84UIAqf0+Di4GM7KVEODRejv5BqPXfAw15
x3yUb3F4yxPl4CKEuXegOrYNKreWZP+qQL7sS4HTkgXZur7RhZA1atImYOq1swos+jYqZeP46+AM
SdjkPj2ijJYRqGcw929onVX8KcRH+KUAKCwPVo6dn73jJA8GFrw+m0bFYKATJUvrAjs8UKjyPk0/
wDvD6OMcdRjHZ8usFy9OOdDxC4x+9Lq7W6i0aJKYrIsDdY7CqGj1nM4rWgjgZV9k1Wly6aA13Ngt
94MTG07XlC1BU28QQWq8WXtpBLwFqhCiT8tA5n31LmHk96eysdsAaLXbT5YvRwpjbz8NvAeUCKa8
rvSsYoijYlTkVgQk7H2kQRkiFr3yLGpbcM3kWkEugCGe17OzVj5eHJ4b2sU6AW7btBlcUdfMQXgy
56vGjO/aMpoeIPnp02XZ+Iojat1d3+WU2OPBsVab3IHBXQOIL8HMIcQ2CkaUo+JvYyz2zsoHuaol
biioqzhV7Ys0oMR3CwBknNhahRTewg+a6sPApWR6lhNKWA22QV4x0IqM88YKPDBCE+cO7i6BcF6h
1woi5PGh7jpFFrJC4sU7dLWns8KrEGmy1hQOW8v6uk8tNvKeBrRiUASN+svx7Oiq0aW44O1UK+wp
I4ttarxa2wZRhgRqm8dRHM6s2alf3rUNxIfxbWXnDo56oH7hcjAbKpNu/h7poN0RfJOiSt+4oQi4
iB893PbWZk4Lpwv/hqSL7jccuZ49w35kTQrwu5hWlOaoJtTFcOqfke6u4vT9agHb/Pzr97O/F0UJ
wqMLoGtjs+pic1z1RjQAWL2UbC7AZhhLcQiv4haYn7pqlSXmFoGDgefagUrE9f8OLuA08taMV7jj
cRMoyl6rJAB6sk+zcjbIzCyFNUCqMzy/Q0kSdmrr94U0iSaNGBn/oCQAeQtIoGxYisLAh6qVw/uz
Z/7GRXgtk91PLWcKI5XbHZrRLomFPTOJo2lTpULnwXcbtTDnEJqEbmzeesW9lL1mZ6LD3ilhigaz
gKC8yG49wi8NFHVMT4z2RiUL+R6uOq1f52k54R5V+UyL9iaQpSRGTRb/I3UG0ZQCSPF+2G3nAkcm
bkya/yDwZn+FmT84jMMdfhaWcr0wSjlPJJ9R22OK+TcuyaumMkL8P72NxrWNazohQ3zg51RGem/7
Ip6tb3PWO4dqpXQ3zFk0H8icoJznqUSUF8d4YNkm/J4s4EvYkESZhYFaqiGYcJ9H6Sef6thQo8AD
/RBORRz+MYwMWscP1V/TrwPfuuBNzEUFJfkFA6iKa+mAdHDoSBQAbq/ljzFs5lt4Qgf8xvnMsXXi
43X2hRigiWmhU/ZKnRKmgS5rYXJlGBe6MaeypTGNat/m6qPNxb+1C4AcaG+py4cp1RzG0Bk8ZJFS
TlGc7ucYUDQwL5zUdp0rZeonfR8GDHGZ4imyZKynkYW3P9gtRGI3Wb+mAUavdgun/aE0qeJ8r5aB
X6dlB4zft3u0JvWRIR65LmxeHS+IMH8NdTnyJ0rI5/P6QVUCBEBS9EvsuM5mmlLKfscHyXzLaSaf
AK/Vv/iQ/MK8MDgDJUFIo6ORhy7KOQLRa36YzBRmtev0YTIt4nyuWV5Kx3Hx2p1+0aUeagzpwS/u
h+WnePbuDHb9QV3hsF7bM69bgwKDsAmWidaw89zh7QPphbbJFDu5pOlT+dftq5wWJulekhs3R8VH
OlT9GCmsrHheAE0cHYsfdT2D/Y+TUurvvuIpfXL2GApoW2IABHMlufnEKAP8CON6b5dr8rbvgCMx
0Fi9YlAmv27YbozFfpdBd8CEcfiF9H3RF+K8Kw2fhAwB6+Kc3f/yxIJIVP65c2YIuq2JoyX1cZhe
lVk+OFSb4v/tZNAVcMkt+/tRw4ncf6n6qbmedlqod0fIOzf1Ki1Isf1I17mmJialAuUIokEJsZlN
fN8vz1ANNseQEvHOoFnDKiDa2l48cKXbiSbu6wBsMSbeL39QAW/FLQwUNr4qJ84yKm2VErej3oKv
1o6XFerahNfiUzcBHCgLHImPRC38dCpWKTeJxCoJP/dX+kNJWeaTcuIGpHPshYyLrlbXRg+Oafoa
nN6sjdDxLP3zS0Q+h27t7WhZKA/VHOG2mFPshwHBy2DLr2f4MgUgEQMW4epKubbKSEYE41/5sweG
DSX5d+cdHcCbc3X+pQqQpMjGbCX8lz/wUKq+Kg2IQ1Xtg1u8UbwVtbA/ZlrCdmaAKj9IJGEK9Uo7
f+gtrOTh9YkN5TcEsF4SuOeJlBeE86j80/yuxVK+TzcpICRvJRC3ccsFEm2Rsh3ThBI4b4BcEt8Q
d8HZiqfyJEkAN1C8qHDpmx28aI90FOdOVyZTMxNVZO++ew9P7pAbuSd2U7mKEUHyWNGT6YwAuhef
cAZVsiqb2lFen6wwQSgVRR6lJjSXpVW0u1N4v7h+wc1agc7UblOeQ5VXGcbjudHQh+SmFsV8+8sc
avs61J27POypswOrrSus/Uxst1KL7fOsNZlmfryeFywh005TUzt3X2Fkg+10pYv1QXVVmQTDtOFv
7jhiOmqwKXTUSw62PZiyKCbUkHeoBRocJxOlsS66E9vAZAXBoBqgmCM3lZVuCaPmp2yZyB4wuxWz
u4QYeJ3tB+WOp0jSnKiSoo2QX2HY/XG11G9xL6EtKtjdiPHZ7pvJ3Rvu0mp8pEDi+pnhkD1hmF4n
yNkZhPuwZeBNZHTYZ6TU8w069Bu7hwF/baIzbXFW4AKO7E1XB0BF9MXKu2L0deSMZ2YAkpOAzBLl
5H0CQGLMBZ5gN3EbN+l1hy/Hj08P320JzrJ9bVvcSPGLbH8d8Gf1LKh+H9BXO8XQXfREIGpRxpyf
QhanZXT2ZS1uyiZpzX90c6hCswx/7ckbrxUUlB0Kn5RHZubtbD/9pKtZIxoHEa+przKlg6gOGVqL
hcItYEvtMWLdJ20DD+sqIjB9HWwbtGTaaJfa1GK38kRmIBcdQtnBvXoDZqDc2zXNIEys/bVDaQnf
3mY+O6UyXce1uUyVNPe4Oo8s4/U91x3nrjJx+RC7SIry6VE11IU0yCnIMIP1ci5UZ62RLjWv+f+Y
axKZQKLbK8Xb4vRPy20tOaqTNLREUYJJ7qFGSubnSiBqTh9t9SVr4WySOhErj1J2Ld0fwS5h41Uz
4BrGbrzkurSASOqP4FNfV4+4SNlZn0nL6TV2A1xs7DESJ8/GVTneJChdO4BAhKgP70ox92BQ2MYY
AEZEGXsyrFHGKD66EzJa9WtR6nSQehVd1+U3P51YzFe4jNT2sw/vw/pZ5ahyWdgp8b8xZKquFwvd
AAvymrvD6JlEfDqiInu5xaga7mTlFz7WxHS/qVy8rTRCAUXv7Om3Bus6C+aT1c9e7nezggq8pQfX
cZ9w4+Wh9MdXfXi25GoeAwczkAbPkBq1CXU12D8GIARfQqZWqCC8FTp/hHUUD0txh/Ygxfz75Sza
vAWZfMAyqu7FKgJXqAnxafsJ/hiPi4V9x5VTqKiai4G02TZBapIQnMWUpiuiCFFYEEZWcwDIsp6D
FoApFaxftshUnTJktueYEP1NX7I86F5j5kvZtjokouuDQJmDppQX2YhIB+5htbdThZ4ckjOGzhTU
/ZEtC1+an1RDYGxYj2SNdlDzzwdb6lg7dVai8eXnQ5Zmnc6PO6GGEeL9HQyXTfFHZitOh9QoxQpG
6u5qpJaGvZojdZDpPBku9kCZputrAFQAim7FG5dcfEyNszaO6MzHiMsfoDk1JvxTiSrpNKJfE0QC
3AyqqPCThwBzPw5m3KuksWn5xyQPVPrZgplfJ2dPdToL6+XlGQV9t5ZSv2hxpg3Hk6gvRGuy/sMg
LiePIfpbzSGtKJFx0xH8XsFbbpCLsvEMkEr8WGFpHUMEa1UcVyqTR9ALxv1R8uhayXzuEOs0zzBI
AHrqpb36v336BwGCvl/v48Giiz0HDA7+7K+3wUNIUKgrwsYnv/opiDDIo+8nWl+49qlAY6oEu8a0
CtDPV7/34Vkrx9ZXH4E62pVOna/NMjiVEa7IYtlVVkKSpV1sD1YGWcmUb0o3lTDnFR/+ZhibP/mV
Il9Vd6GxuUdJxQdui8MCyzMjQS4kFfJGcEVrXgOeyMDY6f5ZU3Ns7fz/Oqz91elFZK1ehjJdey5u
WAdkXZrWl2wHFlmwLTHHDbJdopBHDE4giAvReniW66zYhfRUgxn6p0VmK7m7vhn2l0Net4abu2en
LgStfQlHeH8ijOtIjU3EBdxWD5Srl6UG5X87J+EnqZ31KZev5LC33KSqXfjEIoTBVy3teXLtc5Rv
zwMw5FqE78/b97/MhHRnu2T7nAuoPCYC3GDNfYnkIgD2fgD6z/7OM1vrbcTJ2+5IYSEyS5uWESvo
ZV/jDgAYohIz7tjeeTPhGOeffGH3SU6rLAYTZ+3jmt/DVXbBxs6vSp6bY9BW4RSAOn+HLnCqxEfO
Ia7SQDPjn8hO37dhqRJ81Bkxzs9Z8v47IKSMa+Bfm06D22IQC/RwbJNHF/b14i4DWyR6IR4B1sf+
pk4M0hZxAFE880jd66GirfHAlqKWuwJPw4HHQGlfmk2Mk778pZHqovtFcuNSPQ8wkkVYWJVhoIeB
inVmqPir5LxZ/UHF/hNsGXykXdANHwrmiDd4/U7j1qk9VsGAsuyIFtmrhjbbR0gUu3c5QeydjCqs
l/gYSMFcaqaism5eDRMFmEWzF0iB2qyCBNMiZAEQ8ELwbv9Xn4+n1cOegzfYewdOAm1vHUdnilN4
VfClI388IWLMy/vjWZsrB2WN8RqI/djxkL2NMIGj7FD084jaBkeTZ7nlpllw/1eN5N/l5oIGHbVg
YKHo5pgYtZdDWv9MP0NhEzFjpUkdRFf7eZw0kKK4i8IxKYiVRKazzjcmr2VZuiQJKjrx8zEzcidM
oqAjSjFzbBvAojIQ23igSjSCBj0fOFn1VRh2us/+YbH6a6vwL3OZ/hwJXFdxXvW1V0OZkFrwmdln
O0xP9Ml97noOc/Dqw2keybDqAS2Cpcjv6qdIJRRvQrs80/3mhMWXY5DDxFAbuRVH9PF4/4CEVK67
7F8J5QCGboGrc5uTV/urUAcNqTTQWR63Z1rSyS47IWmt6tYCB9yJvcbOWxANoN8cqqZMzbTreO/L
FT85W58vbx8QIwz01NDXSddb5NGckzC6zH1jLa8U7OhVRIgsT/Fpt4tJ4eQaPV59c97C3shrWM9o
AegS+k32APTA3W9HX3TKbK7YcB+nbzlR0NT30ZcOjbcbcwc/O5WZoNXhBjqj5I9zv7DX2tyEZBbS
N03CqD8XqQdZ1OEAJ1hzDTtF/Tzm2aZjksWeFVq1yB4klYSeKKkdQWeebKfNEWvDvxdMvx4T1EsD
PHIPZeTsmamSwb02lugGsnj5+vR7Oo07CrufZJy4COuvyp7eDUmUHGv98Jg75HJnfW62QTVJMEB8
aviYGsuI65a1jwI8UxFcKSKcs896fPteKTsBE/8xnV+msEskXWBDiynmMmQNUVDEC5+755bmPXpJ
juCioHH2UPAajt5qbk01IbXOT1AlVNfZEgYo8tuQflLQ5GO0/8MRyw6iRI+DKZWZGBUUtotuEArb
i+fLgzGNW2jwCNiZQ4rmSoMaB3iv7duzmorv7qSgbFIve2JPLcVIk+xQuuch4L5lrlGFCPmH5GVw
QeaIKPlM17OJCTwBcUgzI2uAKOSLuYw3+ZTouVS0vl4riLyCzCwatkrcOtepXxxG6HVxKBevq99N
zz28/pQn4+21CXbDGqIXigNdlMW6YP9oYPzDXFjGhitCyTR8tw/2rpzwYymJUOHrkKlB+Od/gOz3
cGNv5ZSyQHcQivZiEPxP1mdwaOpwF58FCORxU9VXrkAO8lsXa1FMPtK0NzK291i0UB2s6bVgZ3JU
ZR+JZGikVRzc63SmBUbd/zkrXxdWhxYF4PjxxtpVBUlX4swnERdzSON3jFceWnofqZ1vc3XzCFhW
NNKguEszjKHyIJXaK5FZ+SsHRj+N8PvqigJWEJpOEC5+VfCz+kOFuElyyahwpurLevxF2yExaDZ4
G8O8yyATJ3GIglC1czhLw/HmPg815dH5ca8dQRIeoUhstxizZVGCFY5Y6QYwemWsMNW4IUiulsLQ
7OlVCtI5yWScb17nyxL8kCxNtSa1pZ84np6BFjO3RUp4n0KKOoOQp+SRT03uShnxSh4WEf0t3Cmh
MIfPfIE4vxWEibMfKyvcsIbSNffOYw92JLg3MYEP2GC7N7HaHATvPm9KALyJlmdZ971oZWj9tPCk
ypyEUXBJv3Ge0kn/nVkhEmHNDt2+k3ZdwU9J5quotbO5bid0OEdLv0owjMgqf5A3XEQBpiJDkTdj
si6tpaLatUprFCKZG9vAdU/og+FpboPwtYnhhR6UD6eO3XK6iQRPO3156SLqGNauq/ZvW/0Ub1dc
VXW+estBDitdZgJ5Wc/SFXaLZj3gXI4SwNB6R2k52BiAonpQyNzHgsw+4EOOHAG6ibE3pP2ZILWD
htv/jt8ThqF27KaVRjF2lAYuzLXgnS3nWRZhWLqFwA1mREnLs8wBlIJlnG0WG2CfdnOUY34v+Atm
G/KH0dcGrVCX8FQTe6k5+rum2ljlRyyhSQXb4gPGr4p0p1QJip/POt9pKMBt9iDuH7KFwrubgXAU
D4nx6WCn1AT0DeuwmFauYRQeUlU4rtotogMMZlUb5Efe7dmyKZhE8OfevCLN2m7IolD1SONEQzCK
PjrVasj4N8BDAG05H8k3qr0urV59amq7O2f95b2++/EVyfieq4BSwN2vyWv3OXT1BQ57ev2EmPf5
hQktWbNQegctecwBe4tEYmb9kzjTQ6GykzLdpPFuTxmG1OnuZApFK1bLssbpu810gZ14Z1gQJ/rT
cuKHvymaUUw92n3+V1Nru2WVe64tZRys9SYY6AZYNlHZIlWySTJFi0HZ80anqCbaM+FLZvgZoS2R
UUh/qtJ2dxo4Eo0AzIp4klsKLDq9C4yl6A2HDDEe3BTFkyIyw6ueLBAXflhj0BjV+PgyCe0JppXQ
TBgLMqXGL4mcHF4zh47Ls+Uhmbg+xU6xua1UGbKBlXnSLfhKve9anXgc/NoKER5o/2Ch/TUdSiqv
cmLdGlOSoLBUMhGp4YUNDfRsnAlOybHGNRDWhq8qEcuPXKMUTFsqJ+y5c/rjcjTXfvU8vHDMJ4gC
Zsc2dpx/jgvL7tacoSgUMg5i1EOuE9eYYTM0NrwlEg0/dNv79SMqZ/10AuFJHEIg2BPRxCX4sMhp
7iika7QsAcVT1pq4e2ZkZFgtFyRPGgifauAWZpCnwh5mOgg/UGMn8kVXhAfv4KwEx+Tc3xrdE6gv
Pl7qunRcOGmqs9AsX68d4xd4d97/+xT5y520bQ28cfiYof6wDhUVtkzv+pDA2aVhrLU208PuWrrQ
6T9BgV7kQvXC53tjY4rZvsG2gqDAiHe5u/zADTe4iiAuGw1pBlAEI61OdLN4bCTUdUg76xWOfUdq
gFarppStcECxj49IlbdmYto2t6+ycVprahR+RWHE+ZmybEjlg7P3eYH98gzXloxmfrmBsIF2lu0p
0vRvxhzJ/2YcawBYuGLlBW+XZhrDS/SWVJx9ZTQFHR1fTVmg7dSqRswVDXNuqtc/Gbd0MyDAowPn
NYri8kl1j+7i04l2P/5mNBNypm5z2TLlEpdZEu+r1ISJoRTqHvFx0rsgxecz2WrOMRVYitwaxyQO
J6i9VC253JhdfGYXVtmOiRA09qyXIk66zsRH1wRUUiYiaLg2EVTycoy2YNVxe7MeIy/7LRgw5UHU
oKT/1BszRTv5rLQvg4ncbPihv6jaMGEy8BxHSc+4omHjWhN2fVqYzaYLiWIzgucaWAopAsv6WbUs
kfHgMslLYQ1euPgiWwvnoeToVGHaLbb1CH4RZF8nQCnle20gcsVN5FGpgEYG2vrigUQWMxCs9y6i
ZbT6uh9JHwZlNMtgw07jsJY0X3RT/0m6sv64hFCStJ13HDXx2uNqo5jauhWinmM5/zpMnpsI7qoP
2fA+wlMnpLK7fttlflXNt6NGTWzQV9XA+RvdZnBEexMf3tSGZmL6dLg1e2WHaof1rZPp7U41Nkg6
nhTr6fH5SSD2oI+LDbxO8vTWO+g4ssIy6CxU/qvvaPn2Z0JEBlyTpaNDsKDbskciY2AgjvOb0/+3
kEZ7uMfG9RbBY6mLfXs4PTUwQQGiOXtMTGknhcWtvKeU7EN7wsXBUsx7aRmC8TIcXgN+GtDkgfqA
6O8cG2b1kiN8lQcn+QF5VDVnvKuSM9tEX5/pcOFm7U5ibi3TQjvDwBXxforeAuVzrfB4ZNeat/6X
lZY+ynzW2qGYhyGXnSEtKMSKJn+zmumxU9G+xsHVNrxLPVBs6YmZdp0tP6LEEdtTUR62Ns+qBkQ9
Uv8UnGCx2qMZqyTUfO8P1ZK5nkkeLf7iqUg9op1yX6irCSF8mnyrOQPVY1QfqGpXIC8VwUsyUuj/
ad2G6F7s53f/gfSnuuo0AyY/bfbLo5R/B1k9Y1mi9xThAZ3hXchzn/QJHAPJyDYzOdFNKmnOJrgs
oSvT10Jp8hKz+Uiq0IgUrxAS4JxfoYlVUwp0Vq8usMP2brzPCo7NB/ZZc/pXU9Fd3gNm2Et0zEdF
n/3YE9vHFQDOXTbPfM3pGK4l0MD4ODLjLc2smTA1J/oyT02mQXkfrIivbWxg8jKFBzLt+WBU8HIP
Z0w+JiKu1an5OqUUyzRkHj2YQ9hdeb/XD7gLrvo2OCP8zVXyno/ARiYIegixcqc4ezl8dLUpCA0a
nC9hNlQ6lp1CZnhoejqj4Y7CYG3RFlFIzNzjunA0sibardYZXfgLaTl+1EmcIRLcbcb814SH/9GY
IOUQ7SvI9u4BboLXhiR/8YcOk52RbLdOSnZV0VCEA/zmAu56NKRmnyKvLjDTMqn5K9thHNQ0H4xi
v3d3ExP2u9+In3Hn+4OqTXyS9G/DncLQ5bjqli3KFviUQ7PLYjABlljdwV7Z8WfRpD4i31+7JfZ8
r5GQVB6C5TnIRfPogVhYHO0dALTAFKPtq73y8NC6rz2pDBgy3bGq/cZoDpu6QKiLCFNNTzHBLlF+
+QLKJzm747TMjvpOEOSVXO6Czuk424nHWgbiKekUHnSGl4mPH6gpFTu8UvlPMd9RjpgC9vHLmNTO
OzlVxh/Z8hUDvk2IAIuJDfLVD56hQpcRH+DWs0DM/AdI7awEpUAibqnfMyJqyFjirqxV+ErSl/gs
ALgZ/Y6lXu8iUZTomIDOa6hOIiR9rCiCMCBvejB1aAPwSxo/lXQtXPnRMkdz3efqsqCBapbAXqM4
ZyINFfHF0x8e56UaWENlpHOIh2t+uHnqztZb0nAOiruxYTXDFGDTq2HhPj+vZWojRBplOMAsest0
RId2Nzhc32WwoCnWZvhocmriAvmoSw53FUGB5gAr4AS7D94yA89AGd/n7l/8SUWbEfwTEl/xo6zE
OzDTn7jLP+K6Y5ZhXlAiKrKdtI/4ML6aqK3l/vGds07SqV1RCwCZt6Cmnv+uMRDxS0AFcva0ETfa
oP8nuBXGtNimfFu7wcn8J63n4kf97I3H/iTrFU11UjxYdJZ0HwpvbqWVh0k3oeGF6L4wolcPXrpu
Gpmkku0hofwstWKASN3GQqdEsBT9chIO3f7SKsU0QiNuAXD9KA/spfT1EGOtv6E5bZkbe7C72t8s
PXmEE9ZfQ9+NhRKOdcU8wUNTVVKnxLA+MR//CtO0K01qVN9tNM3Ttdftwen2KHfVNdUx2NbUU3+9
Im0+By4tUIVCg1RAuK2KnBnNv/L3qs5aLM7ShKAJ8BSVuFF1lVUyT5/mgLNHtiHSPXtQGKRpXXlu
Aaut4OSo5wIUKNgXPFXSuCvgmeTEiOYhoe0kj6V7Ch8p2Vo9USLW9b00/Ei82+70kfp8YiCydWg7
wE4ZQ0q2ZdQjy2SQzThkMN6d6GQ76cctHuWHoIDHx7lYCQE47YVXePN4TaaShQ5IdLWIlVfFnQw+
OedGhLt1+4G4QJKRgr4IU6YuXoiaXyzjdlgZWauaoUdRaN038qEBA2g77enw7pRzvXVWDak1CJDV
hUwF+8sAXDdnh4QNa1g1y3ks/wn46QlaXj0fz56biafBrJH2nb/BaspZZY5uoV6E7tgTLMEHV2eP
c0fGxdwB5IfnQYk+paN8hYIetM8kIybmzekJxcUgLwAlJGxdWolChTTFIahI9Ug7S54+5e67NfiF
dvY3M+uc4JA+jPjWZg9U57jETdKEx/sP+VSQitbuY/wKEjlPtoYZuNJFmQWWloYJFr8mt9ossund
0huV5CzNe5RwvSLdEAf3RoAjxs4xMD/KcHrAczwrplpsAonVr/5pC5pxEbmVi7yAGdRuG0t4oFiS
BvISAepW/DKeZ92DOoRlsIfRnne51QAy+Y8n652XEGtnLBAy3jd8GuEbFG3FyOD0Oqdrkz3Wo/qz
oh07GaTFNYMdk0jpaalQ8+uH1yEshl5qXVScZAnFNGrJrs4DE5FQQN0JtFJ/q9qOuW+dYWv5qRLs
qGjN5qBPdV5W7r4wZUok4hSg0AvUuhQp8041GhD1CZUSoKb7gH84oz7bUB/dsHAilLApd2P029ic
5DPdvMU7k4c26hlpEPrTlT3rkD+R/boNcZ+waIoBwNGxKAcc+yCpgEEqzZbCD5o2PgwabYbwD2sX
S/ckk4mwcsj1b0ebrLjiYIuhHeffex7KUW/Ddn7BYywb1N8FIxUueZpAbXGX9g0lmLDjnYajs2PN
ZhzXipIUlmzSJlT/gL2wmSxSoB3hDNBByUnegE+kMQYPR3X9x2z3WmYCsV0HtQ+dDffI2f0uz9GP
f4+aOn6QUGxiRl5C2GgxfKS3nuWS0zrXllxQAYQwMeD2UXMm7sJ4hRcM3NPEVOVIFP3CuqnVpaol
AHM0hm2nnWXZhBP54fdVNpYTRn3XAnRfksSq0shYjt4VHEjZ6lnqIlZ1b+inRlrkz699STIW8mVr
hp2sL/KjkPUGDPBdfvJj+tUxP/sTGKvpVSxtGdhQEm2/MRaFzagnMemz8iL1YjlQo7zfnZRGlGYX
6A7uXA3fR+n8gwp+s72Fvc+OGTn5MHazgEUMmvtYXpVQteRXvM8/DTBIEhTqb+pSdENGqfUh7oga
+GVNrWK3Hk+dbSf+tdVDkC5zxOylQxsN/AMLZw8I2tmcFzGar7Z4hWywolLlbS38tTdIkSO5oSFb
y8LQMY2a6e/pEqVWUKaFjr6a3xnXCttX0x3W9K4tBoFKPeKRir6xpeUKDOjZbYwv9kT9BG3CdKi6
gKjqQeMdvylkoPDYrfovDGGkV/qDDneSucleWxNYNu38HSEvfDS7+B/jGkR5mNy+fi6CixAzoNiU
uK1e5KRhN/XMVlUUWVkSdXurbpIseGSk+UjizaXQceX5Yz0/aoGbxwsUTvehKm3fBqStHbTEGkbx
8nZ+oiNSDtENG1VGpkdfUNhVVPqBFHfACIR8YzV1P/kMFYC967wHGrK9kV1zrO6krOEVSsDnORkU
N5bbtRS5VMlDvzIR1CX3PEJxbzfBi/fuDY2RGWTuT9XujsFVVfA+C/3nOxEksc2lkuJzUVvz0RSw
fQTmE/WCuwfCDSkSoj5uEE2c9Au2G6KAd3ueHvpRRmseIgq1+PXKbpBFcuDVkkBmYG8TrUdxmxWY
4CwPE17RoMsVhrXwalf7s6bZiE4ORRGHlM5qJn4zJk9XccPPE49aWz6ep5Nvuro593xNnJ5BxOMF
auBFcKWJFK3EMYHagsDk4e4MmltjNWcjX0QEG/KIn4DnZUyH1F3tBG/8z11Jzvn0dPQknmre4GV1
r5KX3i2OGp21iBlhff9KXupkLGOGkgoMw0GKkXhl0fwvcHraxgkxQwBBX29VeivAcLrozF8tM+bl
UfEBStPQcT1u4q/SHbeG19MZptrcgoV5S8xXb2sOvYdBpyRZ6f0ccVZd15Qe5NIgp6YzW//aLAcc
It8cxgPDABnq3KfAp0TMMovh+cZQRO2KhwC5YWGVa3Vt+MgpcU35sClf8tPqaJtlCnitLhS8CMVW
aRQi2LzqF3214iK8E5q1uyJHKuB781exFfw9iBWjM8z8zXM3OZcCnLUsZpfkviRrblT4wmemCezI
f0+loTZzAkX8TaogOeih7tUDYBs8GXnj7Ws3hCEmi30RLFkZywyaKLmPcRvyWH5G45BVZCXEjGJm
IpriP+adOeXxslgiOJ0b+zwr/jy947S3apUR0IB2ZgNkwxatLS8H/JuBXR364krByN7j/rntTv/e
YyKG5dK/R9HJlAZgLcJi0745zS5uaX7b3b26eqP3l0xQOAOuctNOTnRwLACtgFZFpznc9VzNvH5u
O8HfX+Rm4ufhBBw8NQbkmbtFZMZ3vAw6dbBaJBS1vkSRbYO9BrGPsZ+TYPUx5C7uiJ+C5WPbyM+C
WJmnWKsn+ow+/u4IRAtNF7A04JIM06lXEgtp2awQN1vnJPVchQ7P6iZWfRB7cvMrjM4QbJjxz2K6
8uylCCoGgFsbhK1a8uVwQDCgquN0+srDhKZ3yWlykqN9rZqdFA4b5OKNnS4fJY1VpMxI0+F6iDIJ
Pjq5HavMI501qhMBwSpYrtqHUBXOJF/4UpEFUcb+dFbIzAytwMqvECAXCDJtukkvcoZdwLmylCqJ
JFk3xJa29NmbsEsxFFiY097JyIec8VrO46D1o5sieEaGIWpwDyrPjUo1u1J6b7gOlx8GN4ueaQ3W
RWr4xlB4fs6lqR/r4JCySzZC6qxK9gxt+dn7e3Gepqo4wrvLlx+OCZJGsZorPJE2i/zsg7ajahPx
cR/76siRolJilo7mIUz5D61KMYJe2+ELAgqGzLUF5odECqhDh6Txbm0ZScmW4BuSAArz+chOgX0O
PrXOnaYFjpjLtxRnYH20CJ5Q8lOKn/F04Lg0qdwiCHTazh3G4QJYhX4nTDy9BVpYUGA+ZEHzfMq5
Mj5NQWebzr7dKk2VAVJBCFicK1vwe0TR1YvCCox1t1kJ4BkvJ9u0mcGh2u+AMZTJtJmj/TKu/MTj
BjX7q0pLSbW1d4aaPYb7HOd7lSBECFQPcz2hN/cizaFdFoMEb/vwDhcQLqrWPawG/fkD0hV7g+RN
6Dx+pfBkU/XZEuDeE+fwJMJiCHk9B+tko/BODGTX0MbQ62MjmrKeCY/y33X1pvcrT77s/GZvYYOd
7QvOD8vrMMIsh1yHTKd0pwp/0pku13SQMtE3K8/ArVYwMgLJrhNqBg8WgzbZQj50Js2LxRgpED0S
qoKj40cKxGISpW2wvmBeok9gTnQaC6kVtHdttJqmIFIFSALR0wTZHPJ0b7JIBSKP3VuMFmzx6ith
zRqqOxwT7CINqj8KSKEb6zjDAGiVV4rLmFFlJp+tcrLFDVcbKjH8JtQY+EPVn/P1MaQbqA4yI5yg
2CBiihQobWeLED9AeXQBSDTY+NQY19iqlKf6GCNE/g8S/8XBuej0f8QWexkWbFYxLLkSURYCp/TC
UdBdyjE1AlkFtK2T6PPcLWMpZKBEpfbzKyRGuH0VHBw1WwCCoaYRYuaWchOvf6e7+VdoW/OdbUAl
oedbWCsKH+1cTrRn1pHDcApjwtjXjFxiFY9fAEkw6M0vTkBe/7K6OlCS3eW/rSADazBbrWEE6OTU
B7yVaSGq11BKbCA8Urg8ac5hbQSlN7dqE2+Xxxb2+Zt3/KAqM2r+K2VZcIAODgTlk/N//Sd5uRjZ
pEKAnDqkLMdt7KjX2/FwTr3j5ahC6owkQ3bwHZnXb3u8jUR5yYYw/0xFbfXgfY6qNzmqNXBWc+fU
tT8kqx2mTwffRboUD4pDEGRYGa/GOPO6jnx+0sU6xTD1ei0joLMkjlt2DM6QKAbFGz6AZeYz7A2E
JUNjy6+ERWAHVfaXcDrAZoaNxhnXPVn2usJmqiOV+A0u73dpvKpO6bcpbV1qeHTRHIJmbFTfTnz4
ejB1OG7CwslAyNS3yHfkJWTf5XjwjSz/KdV0i9qiVuCVyQwCnYFkW3nEcR4KRaCdhfcn+qS901yv
Z+cNKXUBgLpVkkFqGKUdekgofRezAGJ47K3ws2lE0JujzmjBT2CAMO/uVi97SeuxtnEsUPUA5NO1
Hww6Nb8rSyN2M/6M4Xy1Aiik8ksbQOXJkZPTPS9WgGLj/QK5N/kvByIhKLivLl2aWdTQR4WHIvUc
MujSwr1bGSNeI6aOpECU2Co9I8MzZZRRhBY5Gs+EMhkG9Z5dxyU9hSfPNVOLtueOArtS8lfm4k/u
Zd8H+fZVet7IC4cIF6DdcrzARUOSI/vNIv4V84zy1wk+t3vhItKnfvOZvr8be/NTgv3+iCRkaWyA
VDhzSn30r9urml9NOjkr+yRiZr/yxx7vbQRpVtt0Cx/ElT8iqxw61WfnAGi5gY04QKGAO1TI1fQ9
jI71/R+FOSg1VdXtRKHOgqPXE1J1jVTJuzTr7q3pUSuxxQIhsoZTfOAF3PnwARjCWVtvv6sEAeXa
bd+A93qRS6ewbzls+dHoWvJHIrS42N8l1H84it5wX4aybNWSbbo6wNTGG+X02n/oP2PQg6SBzUN7
5HQijDWxIJj+vJsoql5IK4xnU3pg3qTfw5Esc+fAI0H3s5OX5L/Z7iWh9pt6SUQT5rX/VSOXclKW
jzxvtkba/hBPM5lel/EIoKmxod8RZ06ctA3CvJ2XlzqZGhO9xFBo+vDw5CyJcpWgbvC7UkLiwNWK
wta/Jbn19ZHtMFQQk014hElmmMfojY2xqITRNsz7GKcHzWDsTludaRqsncsaMLkmff0VT3XV58e1
EZxLw2BRcv9q53TXI+SAVMEDMKhXc2X6Oc4IU+0hYPgUBlHHLKDi8dDdJg/sjeJjAHzGHjsg0D9S
Bc18H3Qq7pjSb4nbtGPfM8j86jg/IWUUqnHfhfG0P8ZmPMU9wq28mqJUVL593vyDk/blY060HPhE
5Hc5uKF808bBltlQk06/S8Kn46HHAMoctfJmbkGT1KFV/RZxppTd2BrX6AiaafWzD7MDh+ssaBWU
ntYLlZXF2u4jKjc+TQhNw+dy6ALtIF84rcpaElJvyKO6VIIvI3S26vu2pdNOt2puEZC1DDDwkB86
c9y6RvwnuUXcW7FTxnuFnV840WLGXYv3bIfHiH4VKERKG3Lg0I9CTYC7RWyEExh4tkmTNUF1QjJi
tq1QFPzAneqpIks4QRw7ZXzsRzFr5Do0XIQex3+EMauf7j8t3XZXVIDchwH+lIaAQOJoUPZ/rc1g
dJJJy8ZLZaMUVYznkzzzw7nyQ1VRDJGkRcEQD9m1jiSWqV+uGsd4bXx4fw364Tun9JC8FGzqxIO6
ijs3419iU8gyy4bU64cPWzVBCxbqnFwbEticrrxLC031IN9ec3/YnZ3dOYa7EXaw5ifn4MCMBixX
uWMb7PVTsEtZtQsATZm+bUT/o6JqEJzhwnw0VT7EVma7qklNUkOJH1dOO8pt/ptjXXW5XwMR85pF
gU7wmG0flRT4D66WMIMlGVh+VBVpD+QdgP8q23g/PMsLG9fT95puory2MN5hpxiTSSWQH30LIFva
P5FBiTmGSxlK6l4/AaOlL1sdf+smKTmV6RulxbjRGWNYjVd1mSeRG1rYJy9qNKWR10AWu73kmRay
Iw99DEZZ2n/jSVD4MqXAVlBGzNaBCyPVpPxWp7enxJFqASSj5vg2cfRZCzrg8pQjB66eEbQARsVg
dAEooonbVbHxDJPw4m3j7a9ulED9DDbH8tYZJy091IgeFYRaGP615DqJsXSx8JVJdZOvf13feq/v
7QHDoSXx2xWrnxD2Q2e3fJYUFY6iwgIa7yerN2Vh+ih+woWvR1/ymyP5VkoozcaJMmSSvsZkuAO8
g8tGEfkemGUH14VcD93EhEB9NMNhpjQqB+Z7dfnUocyBmEkqejcJn1F6ifuyERfG6e3JlQS43LjL
97JgD/HOUIqaTve0uF5/PGn7uWj8JoMqL3aBIwybrtU0Tz9CT9LoxS5et9+euM5YuFh4qQzfPB+r
JkdBuCabr4bmkAH6sRGxrtOci9AG/p2uM9ch50WfRFvrw4m9o8RYjx/8YtMYR9DGYS/AMPfKtnle
ckttlVw6zuxV6B65PwmgTc892SaLcW9sgFhmcEz1dnm8I4WsMt1LsO7wNMv04yRXQBmtiTgBKvcf
ZPJNhZuvZ6ZtKVUsJ6oLYrxa3lP9TKuyAsFM2pgZSwGjLFk3KcEoEZcnbSOGmQozIUyAv/cMj7fi
yKRllL/xb/sqahxfAofVGtUGFFcBORgVqzU3CcpKhlnxnzAKKR/SHRez5VWMu00TJaMo1qI1OCtT
FzO8RweTt1L9yt0yAEwGUECI1uAFyyj70NtUrzeZL592xFQxfFDxgP7Dr3LzIWv194COmUmq3aOU
JsGwzsVoDX1UDvJpdk2EYfXtszC33RlAquyaHYI1kEKQZ3IIqclBZK+MwaxS0Ih7tsMizlgbzXPV
9zK+w/kTQgJDhidl5aGPGmq7Ex9AzXlZS9PIXj+eU0Esz59AQB0g0Klv/H7xYj3FQxS94x0rqbEU
ma8LVR8fLsIJ81QAEoxrzpRZ9aj7gPPuRHQg2o8MLuKKfzaQZu0SDlJCMzaeQGAUE/nmdfX6y6Fu
tIacbyP8e/WwKvuKoiu5UTKdPWWMYAU3Z3HPr8q3soH6/SuPLQ9RMOSAuIhE5d9xaVHC7PL+XfKQ
TxyPnH0Nj2tStal7Fblvpw/kW4DOUgEuPx/G4y2kd9sKq+Wqn2trnlhBmf7CgKaFsDL2XaabXRLd
4kMcOVkwSZrTFp5nK4iTcgo3nS417d4Ud+oWNf+o4JO7MwFYVlimeilVsEujI14M9Y7i11/f4mZx
oVAEmRKGAcWk/ExtuhVSr4feqeX/KbmPO3n+zUi0yOPA2/gPawbXwO9kKy+BcRJ2AvjOxPvqS9Vl
CfVzqEKQLx75JABlKR2WLEf+4ngtguDGU2Y/XcyCsjGqsoA+pvMiWdo1hnNdyIC+22jY7QwABrAA
f0N0B5l87m4ZGplXmCB9xGYiEzT+hTXCglGFZPPYuaxikWiGTYNryD5IcQYEJ1XYnv7JteqknhGh
SxSSa34UWiImNgiH8kzktN5VrBdnJYDBHczuJTCCwaYAKri7fHNbAKRHW9k1dKuXUDIEVZK/nd1E
DAxuOkMZyP2FnEGSA6D4kFIHHkvUH7XLoT3/gijvGOaPscyviNTES6vGfJsDylH1d4NFHvy3o8PS
6gAZewxNIIQai9fS1f5l2/QIJwNvjdzfgfQQDCV6cbadftO/0s9ES3gf9AiR7az0HNlkuEMIl7yP
J74L4Vl4j1uzhcrS57KSGViy0RCkLlHtOtTZ4tewBfXd7Whs7wWmeEb0AgNg8F+qauOPyQews6l1
9JJJkWbuTaOvRZURFRo8eVpHtWl2WUZzQnIwHkA97veXvqLU4eurWzbBzAq6ViyMTzabhAy7TdZa
E7nMKXJPHTxgcZHkrwhaSihSNZdsI/PaEz7hgbqXdS2kDbsYTk7Ckui38w55LyrIlbXNAxcsBbvU
Z6jo0lFLB4ns9SNDxjPj41YdpU3Lf3bSmc/vKiRrVgs+B7w4XX0V9UAFMinZVmoXC2VDf4wAmca1
+O3plQKNy7HYV3qU5IXDNrvCZU3l6bdvtCxe6MJul6NkoMWU6poE3TunOzKV+kaD4BNAMwaSGLZ+
HfCQ33VL+QOFd5HsXqzcKtNL6ecIbNt0+qeUMgHvEUJp8fANVwsfA0wFezH9/3sY34qXS/pEaqAG
J20kagKqJXJg74N+UL2hq/ylzI1ubhzys18qNNwJ5rYRWUW8RXooHYHL1rLHdeV3SF8M+zjwLMeI
OoIl9Dnsqe9dHAqnTCQNZY3UQ3ws8n0KA6yUFaQ6SG1+nliYxFsEpAYpM28QnQYNu360mOOpK+0i
y0hiaqLL3WgspG8JN3rMe9s1L2BGXadISNnM8MOx+remFlPOsXNR+snHlRspI6S2zwwlrMM3L3z7
CSLzmHzh+/YzIomv/9xH6X0hg2v65/6bWkYnSOzloe3K4jlrwrLDhqYEeVE341+4nwWJrOlelpeT
GL885AB0YIDtkuni2iVXTInRBcyVvHLE1j1Jf06+4hHEATL6ozC6DreFi/i2y09swxLyovhULcvc
C5tbFAkKfGzPzrAhMluUmjNPILRRtQnvYRMpe2549dcqWMPqjgQJQSTgCRWows236RbupYIaMUSE
2alzRHdf+XEt+Xo0DIo6o2z5na8FUOIsVZAhFrPuIyoHx1F4izWe0T2SFiKO1TwwlCgBtIts0hQZ
Bdg5ihLDb4KhF1Dy9czUtTdcdILOZlEgmhD4lJVVbSnLSQuv1M9LkaDzzq9wbFxG07jCj6/xCJhX
ukbxBQxlB/1yUJAQKMtArBxXZezeGfcxszgtswe9o4J+62sZ+QetjoOZm7rB0iKUyRB4XyUDW+ib
MIsA+OFCYHz5T1XIBGazzo5+AWUGdZdN0dg3973/Po8MFWSFGD3ZC9wshJa5QT+2t+f82wyhW8rq
+a3ZWSS1S9qaKitepkD12N99QELEb60Sn5dkXiHoFunbSsosYb/ku1ksiB6fuAPU1eXDdQg5SPo+
FlQYyMYOSVPERuE2z1itUf4/aoBN8YeF+ybIJAed53dRg3UHCYTKhB+OPIg6p91VCMaZ1G/IyXUR
Lb3S3LYNpChG8sIczPyXw3/+eYcs05C1hz5byxBbt8FcopLfwQUonSrzVj+cNffMObgjSsYoat8M
2NTN+IN2v9fSWCQIpulci4dB6wG7ddZZ7J1m3p+QDd6MCCcexOhM0A8VAynrj/jY6oHW2hB+ba1v
QIqS50wL0sH44puQwkE25p74bcbZgA4tLSRiim9LI+2ZFy9YMC52mJTXyBC6Akrlvfnl6q6+moCl
C0FsB7ScugIKvOFji24i+81IqcenTkRzDeCgpamH+QEzYfFsEc+qz7z/j/XpU28iaVeVRbGmzd9E
77DWFn8UbkPGaHf/ek3wFLSH5EUzWK9NsHBz3uXIZ/zE/MmIh8H+CiGzuww4m/aHjL+ZdEH0PsFP
p09gFqLY6a9Zzm3vNzIR6AoBNddEfuFUdLm0p24zqaMpbMdaISmLQLrZbM9eELvy3LLth8EoueGM
EnF9hv2M5AbYT4iHmRJ+gkPJjvAeVMf4TeknNxBa626ZCxBgoUvT8bteCEOWkKbJ9X/KCNDa3PKm
cG2xEFOAAF7LqVQxzNcBe9zgpajKChfyDXPvTjS50gG8E3XtDXaWYZxgncHuenCzeUtkGHATyrvR
ORbLquuUEd2uDfh9muuyhYcx7apS8VfVq2FyyPdWx273VNM7qNdhz+hFD0Kxj1FCzNVQMcUVHGwD
/YuMdNneh+S1LzD9OFwxVcgOYf2fghMiEdb/QuXC+kuUGtjAOxrHJw89c1BfGq047/NfCUfNPUWG
6UeiVn6u/nf+tPrdpz1SjLsXMxrHFqP3snj15w/coCuGR9VLARipbITU7HYEpzBqv9RtQH7/EX9S
BmumxxiAYXI2ezpay4HaKdjUw3GLo2szgpGc/habm/oec208Qp2lxaxHyBtggYrH5KR5wQXvBkhi
EKAliJPDISg4DnEXvkwKLxB/oOU9MFobMDjfHr95yOPgGPmarNHAIX3EwJPjVSy63uydc1cuuGl9
UOLUi8hEbfBR5aaay6/UrRZ8nSGHUePpOALmalEawGgOQjOpyy6i7lVGQoolEjOrDra8tCB5Qnff
BPCIxK/w9apPYbGfwZoK0AfUeycrVuHBkOfghA25vAoYHOITsGudRDvN5WKN5nr4QXjmSwVtwiqD
bJ86PYkQ1Uaij7B+x8fm4XH5N54tlQ8mOvMyhJ4RbnZz6ANkZmbfjTCEznGbPM9xKWal2edkQ9O4
k8LTidCXWbomFwSomLfk+CNVDt2ml4fvfTOcl0yPL4KZhkXhs5kJdqnPvTv5MpwwngsjP90Blo9k
vlZRYDh4oSdQRk22BOjXE7v//m0epzr0F2wEYeaJBV9MWJvR1P73P17XykCTGqrWHd7XgF+i0W8s
UHTXtn4nDCcmpF3UPrueMvqDtZGYHy07upuByAgQV3d6FkcSbgbEWg/sXKOQSkhCCgqE219t/2/V
Wo5VCw7o3PErATGcLqIjBw3wYzPdjIBQBU+OlSrP9PRru3eg+G+KMuy6Sv7PLuDk5W967vkF7iJC
mGXMZhXf/KM4Im0CPFypDGukCrt61WMIkQ8RUZI1i4432pu1SguFRDB1IheOzZ0vT0Fqd+KCl9a4
VaDlurAn97zscA0HQAAfvfGj+AIn/6uhw56xiMvOtJ2I29Q7G9rVthBtunKS/cqm++7ioEW4WQhD
V7Q3xnangEmsB6AjLcfMSetw62eD5qAsXSMSv9KKVxnZPX+/83/PS2zX0AzFs7hrgNiiddevstF+
cGoUhMVDIjzz+t9aSFbW35DxqI1crVXIMwhnKuQQ0Mq8EhMZirLvRcGvv6CA3nCDI5pZnIiczcbo
FETdhS4xkD+ElK07v+R17lH0LXGCEheBJ3/hj+RpvIE+veZb4kCO0RKhwnPEwp5hlsuSuUvCdifX
3pK8yyfcNNAzkO5YgSzkmRDZ+91aVu8rOyAUkjEgWohOT8uAdHi3I6z8X1Km0PCJhmyFJ4s8XWOU
VyAgDQ0wiJ+r5PPxZ89jcGS7kjXkZfrJETyusQnzac2Bn0Q7Y6Dibxm36f8owflzs4G7cIOvAame
Y0bbB4/zlewqMQ+2arcHCfdYLA62mZBhzcnsBvyeJD61Oyp2G90iODZOAC9U5OuSjYPICoL1rMiU
Bhxul4RQiU7ZzLI9cOPgqDn02jybKNM+6R0nnvDYT1oiAZkLDYStdsCWEZxLi6oNDEU4lHbgrZSz
PR9UjONkKRjwKey0lXODH7DaI7bnbISZ1yBktfMBorDWGoKRwLdAZJ2uzRl3fpvkX/KZrH56fQwa
yjNv3WTRWc9IrseLP12PcZI12cMugoLUiOqqnXY4Ugso4GqC0iUhVul0S2F782NIpMKKDtjb56UH
TUNO20jbQLjqk8aCNv9IzhtzvJrJ/wMwf7lnm0gJCSkvBlCeWTEZb3QSk6mTEGp+s1Xr1in071TV
RXtDzAhbNvDoJhLs+WlFEMix83jHnqWUdaKgGcg8uHwrn+o05jCykMJq8q+XIYfZjOYGATR/orX6
7bx8Na9CJo6HD/dSSD3pCOOB5+yAQrb9wOsy8jRmHD1ciJ2BK3sW5Lgcn79Na8R53P5myBWhG6nR
koRXaSZhFvC+mHinggQQjtt+4QnUyoAk6Z2v6+Y3ctl2gtqlGN6Mg1MuwpTXVhMOEuaz2bDDWtot
HJLKm1jccGjIYBoTu3e21OT/R7GYRTKWXuYCd1vEF3yhTeS/z2ijes60sC72QiYywE0GuABAxkQR
Qs22RBWNLKHKpFcNLBMlRni7lHD0FGCaHdTQhTOpdA+lzqMbhuHbff4nAa1IbC7VXX73nnLDrem8
EW+GoxUo59HiauX3cPju2Q7pVO7VSRVH950p8HlXnTbOgLLMxbBPEyeSwcJFnAzjNfHDMu3IDJai
bN2mvhxMyw5V8YA8E+20xuWMCjVZ2/FN7TpKf9Ud5vpCoGMP2IbWACuVxxAVYJsKUQm9NX3WkSg3
ap7Xj1AlR+JSS72rZwuhe7uztdhSOyI+VXWHtahIQsMtMs7961MuxU4nJ9AOblv0R4s076SG/jZ9
SvC7K2Qq4/Kg14V5th1nXPbNiTVD
`pragma protect end_protected
