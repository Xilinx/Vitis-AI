/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2021.1"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
cDbEQIXrrFOYVkt+S98zy1EZxWD0ccgWupPE+5oJq2Ca0c2em+nRfD1a7i7EuzvxQCBKk4yO8Gxa
hr/ypv/0pnnCUjBVYico4Wx6EP0toFapCWS4x+26Y1+33hIrh1Wwe0rg76NWf3AgqCLiN7oeTjY9
3AA83t6UWZFPph2rHTpL4JSUjnHIURfzF6W2AfRYpxWI1LN/0NUo5dLuBr2MDZ75boS3tIyKOkj6
cfEmuya/7yutfuyCqzt9iy/C+MmQp/MF/Hz6y/xBrKehypeGCKZ+mUXnfkzQCAK8UHeLiOPNAYvS
f5OCSn7fD5AI9Kk2WkUQHE0fQSz6UO81FVCdng==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="q3r1HqVJSVyIJpYBAvyqo50RiOsgeEHhOl3B0P8Rxf8="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1398000)
`pragma protect data_block
nRLK1g5zabzRKTTJJuUHIQs7gHPOVerHTehHzzgJQ8G65vUSR73DuqZxn6cNGRL6LfZlxWdaH7As
ay3FTC2cIUZsRbo552/hExLty9QoFOWwng9n4yhO8zpuUg7S5w8Qeo/4OJ8RW1EBZtOeW+KBP8P0
1BRmb5qiH6iW2o2TlpKd7OEMnqnFFjvzjPEnyww1XZAQStGs020lNJ8XJCKYMu8ZQ/sXLptcV3Ga
b943ttLCSgsWadEKTc5JBfSrltnxShO4MkYhXtLZBL5NHTeZsPWEGz0yHoAN0qROhPnK6eG8OerP
kJY6cjhU80LnRfH90VUW+OrHUWblF11ySDZCR6m3eDbF3d3Jfey7adMlnQEjw9EZF62D8ThCPWex
Q1UiVW6O/kVITvKd6CPQA644rQ9Scysv3yUR+SzcP3L67VgR/PzdMkBN3nWOTOSX126WmR9KvmCW
r5qZhwd9EAOwObC+ZyT+kbUNmPYTPAtTRPrQJw8l1vBTccasQVpUBYAMOUX5Ed+4yZUnIGlxP8bF
7N71gThUY3KVKonGNc3eaWDrHe858Pbkxfy9oQv1vLoAF4ODWULyCpLeCMvPbBauxImvBh1yADhv
0FgmHaCwp3inrCldOvFrkDYGNyqfVYMZvSLckDqqQsbWY+AOHztKNEc+B80Ma1RWfc+BxcIYpBaS
XvSwOfT67SNxQKGrCAxIWr2jxEEMOOFVmIWn8eAaKs8MuG4PCMHGJLlwrXHYgWdQkgepdB+Q8ySY
ApKm4W92fTnsUnHzgo50SHcF2hv/rq4zxmeLBvbb3sfewoalyqwVuj+OcHFfz/W0FOCbC6vOV1VB
nCelhHPX44Pa0W36fXzdk9LKaa/wBV1iT0BKrPT4+QpeV+zQ1DfLe4r+DnV1DwNrAZbOTh2xjr3X
bXECBs9WP3nVbwS6mBzMK80z78L+ECJJCVcjtymwqaPIqUmL/Mwc3qrxqmvnnLHjDmNPQ4q7MC0Y
N5QCwChoowHiyvIIEhSWwYRFjT/ldZGDqq23QNuKb43Uv+LqgHbHiy8Y6TkyjvzJObf9Z8mzKl2D
Hufm7s4f3GCTO/MyOejDRC7jLjs4w00UyfM9N+RhMOLE9FefFCiqV65LTUPIG9KnHHrzfPjz+9Gx
mUHRolNGV0o61CcLscMKWFNW5R9FFkZYSlFn0dyQBgrJFDLohchV3h1KPVLvVgIkzSzjnJdiYaJo
SrAH8NfSIzaH9vFGLFEzCBc9eydE75/Jo/fbp2JPqMHAPJqX4pgbb1sIjIHvTnnviOfULNsffR6H
EfIZM2PFPx5wEynkkiyf2VTMtfBYsXnw5ZGNcZJXFyc068CukQNLANYp1p6Mgv8GOWeVXrUdA4p3
te5zBgVIveyDO9JtliwKwHhAaW4da3VaX3DKo97Pi1OXSSVgxRmX3xm3i6bJVdzM5/qmg5esG9Wd
zrem++fjBaCupAwpLT8ZAuUEv7s8zY7CrjFFPGPeD2NErMAW72V9yF7LJPa46sXVLprMD6XXsSlG
dkicdFHFIz5kycYlDgOwVFktdAdSbXG2XwSeexhwfIRW1O5jGkp/SeYHj4Qxwt2vakf6HJiE1gGw
VXstG2lOAT8zApmH5Gvh1HlsHNa72GMCX3L20pVlL4QT+SpoAeBJtDWtUdSTmBftk/DYLyLt1iTx
bsxBki3prorR9GBySBorDn6fR2XhxkaNGgRLQ42LnKtsBXvx8G1sQfRAWq7wDGSLT2h/hpVQjNLx
9yk22U+nNwPCHXw/pBjTdKmj/80+5r0CI/oy9WOGLpBGM/Rh2X6eVo2IdcDfd8l/EfKSWAAXefK/
nRfR/1ETalxCYuLsNFR9h6ghUizT5oN6jaqeQ4TkbOsJQGoFGJRyLtGq8DEyqbdLmVDpQLqLdsx2
FvSNdcThkfEPMXgtHPscKbOgB9WUfldkkGflwk/5bZJlKiRuHjwUT8kLSCyAmVA1VdxE4UnIEGHO
uV1o83OqWJ+GV2GQctFsBKIxU4Enbi6UQSLbh2YXUegf6ATSEFYObW8f7oKsHKjDQYZEKtl7q/1D
A+FWmzw3IEZtLS/+JNQKnBhvZ+qC2H3Sb4Ufn7Oxs78B9RZt5i3O2X03J+rkfqEfLY40QvCY/Vdt
SRouEjASuEAeuWmPLLlbSMWUeLLrLLuDFvbcs1YvTdxb49zsaJqYRgwxSNVIMJTgBKjTGhmpSrzh
UzhEH1ZVTSCh5Gk5bzGfck2CA6oSIBrTqZfPTNWCCK70iWxNyb6WhlPW0iuTPaFGGuxnEyPORPCb
IWrJ6xCrt69i0AW99GQQWzKx21uHul7NQNGq+rmqKxLQOI3RR0Cq1sIhEW5AVifIcbXCe5Giyisj
AO2M3unzfPZsR1NMKqtiHJTfa7DuAKnDykvv8XsNO4rBR9htgbLPFvcuQZ4YUDFhIEU9xwu1KdAP
aoukWHzR+uDCKYEHFvVv1fUj870ayZs0OsKAPm83OsLg3syQiq6bEN115TqQAx63H7zbBtxb/YwF
qkUBdiZ8dlgvz6yt8vsfiG2LURS41YaNPG9XTEHrcgeUXRQhGhJZIvBLYEpAN2kZBMhxrokJixgX
Iu6NNf6vgCtx6t3tS+yo28e6zL9v5P74KFoN02TRKqK0MdRmK3bOd1i0FReCiuxcMPMNHGKiB/lg
ZhSqcVrOU6MabI0q3R3BFhWr+Qn983/vn3ZhC94q2MLln3bPwPugn4TAl3iuFS19eTe2UcTcbGpQ
MHeBm0mUY1yHfsGLw3L2D/U06Mh04c5JLNseLn/D5yBqy/J97p2m0RTqoOAVRar8F4JEVRDZdFGl
X/iqHYenIgNUoxGWos8NwctRRHboKlfiT7HSBtr7XPpjrdKfrmnETksrBR/Ugwr0kHqpDuX7OQzp
JAHRQxpIJ18kMk/QbQz1oBqdKAyg9gKB9OHlh7z93AKoJ0Mu/hrc0RY9kWPNREtYDnDJIAKRMAYw
TIqlYQ+RzG54BMcebLDXLAguzPeJkrwCtEOb2WqfuFmsJ933FaeV+kr3lWQnOP0ZPv4FWR097ThZ
XF63wHs5NYbPKQAuEmSS96/j9/7mnPNbui1Cl2LmqB+OVoa/m67PBqDrwO9R7p+qMVaxpIqsc/Lc
QkMxZC9zVTB7OBaZBPXYAZdeB4/Q21ovhUUbK51Pk9e3StgAAQw6575e9DkA84OeVFBmiEs82XwM
p0qDppfbxdwAqf0g9qyEsJu3xCAk401Pydg3MCgpcGm3d1tZcFdUD1NFdZtRLpZVxgw2yZMvi061
B7hEGeLGElorEAnsBARvOMmPQU52HV//z7D73XFBPzVHI8JohVLXTJwl9PO0/YnlDTTODJhTz4MT
CAh750x24m8iwkdEGWCsXDiO3eG6yaqppDJRGhjKDNJ2V2k1URLd2sWGWzUuh1sdOinl+Qqb3xez
vnt/CAJz+QAuDvo8YmxgNCAW3WAxGnTBlOLzvA7YX1LQn6azIAW+UppDxwQY9u+T7D54lrETX3+N
w0rpLxJCU/5e6IKTUdCD/AR0VyAsHWA4R+KiljSwWyMh87jQ5ySLm/5a+74WJi7dGFAHK3nWc2jS
EOtQhW94GFCGKNFs/NqbusxJL7iMC1sS2mTFQdOiekFPGcWgv+A4+FjVzgkTV5d4XZZNfEBlZh5k
uMBF6xHvvZYqSzsAJCr8lCCSWqgosY9yJMldjSOGcUY/TPDtyTl2U3I1okpOxZh79UNfzZGYuaCJ
l9KkYFmveDeEIGlODuu/ctXAjT3lJTIfAr69mB73RLQ5A48i23AWw6RQJn5sT/PXr0cYDMwZUUkw
JTGkvCwBaXs6nYtHyLiUPtlZlXDIm0zvnqwvJDHBtlSIcIW/LFHlidrO5P2IdsD9FP+LRTpWO12o
NcG+CrzYsCUerqeiCOlCr9veKdEzWc1pC6q6DyNregzMmW78evCbT/BBK6xPLttljafp47oAXVQH
S9gdBAkJwjxw2REkUAAsWTZmlE+fINhyFQRwcf9Otl1mdD14Iq/O+ei4PQsh0sRtXgCJefJrJztf
c1Oyd2uEoVASkCrpHIJEL6J6hqORHEfTcSc9tnWrYeSZrbqjZNhoTuxM1v8rsdHpNLQEVkAtqnHl
/Tin801gSnh6AORAehxNJ75qYib3gtB8LpppD3mYX6Ww+aL8A83sBZwgocHOpsEdbDti6M5ARXd/
Iq+SM/u5JAnmP2l2fIvOSon3wa2RGrakLg8hFwa05+/cHUTyPgxe6/U+bsv1AGFt+CbwkwtglnVd
oW8QSzrWkLTSKvk/76NZHWREk0BWLYuFMLb2zD/Bn4S0MjfXyo02QN4YYR1UcIYV7W9Q/JSV7kXE
ohDbajwXWuQDRdJ1F2wNm2W7kD8+tiFRND0KS3i+AUtsNV7LewAEKd4wwZMX0N/v1aBILeOmTzN9
pRbRn/W1KPODnGAaeYxyGLPIXRsgG6ydIbe5MbLwRnZSXIJ4RjuZbfj70JctTJTDPXPVOH/QEtym
GCsfF6jVwq/MraeLdh1NOviTG2t1uY1EcYXSXOi2selvUoObJOCGol/sqf5libFzYIENJS0D7gLg
yKJnQAWtMwdPPt4phfSKYfetKmtb5rfN32RefBPiu8+JdaAFp63ypLn70v5QCd0cpFhq+mXUUqwh
EzSH5VlkI0wTyMkeRve04zixWzJqhb4SVOeYGLP2DiewOma1LAbBKNukcHhrt/KiDkf6ccBFsZw1
MADvva6AFz4CU2FNJeCwU68TxtDYNaUiU4w1kKVjKM26q3JhorCpX/cBaJ0KdmgaMwJaHUQHve/t
6D3ZVleV2fWb77FsTAPtKz8Qm36dBcP7UnRouxkYrNW+exin9pXWUfYd5s+OCEUwOQ4y7zxveWRV
P+vNRcNgAEv77Q6bfAHGhKQ5+gXGcIu3tlhy9emhvYKyjXNBYxROZ+ycUy8nj8awYl0vA58N2I5Y
g8L8Wn4ANF/R6pNDfkmzSoV52ehxXo0u86f4zMgQGr/szCBTPDgiS3oUZGOFnNaZ5KJ69X6rxYXH
6vcPzS/3+6B+bvkfrSmg+Wb5D8Wts7TVlFycR2Abm2wkvs1K5bmWRqUBWLGTYByjrlWdtdVNmYwB
0O6HVDoAV8yphhcUj7y9s8YaSPXKHgz6cLWoTxmUQ13y+pOrL9hqNg1hl9UkAda8o7gllLj0o+cV
CgkEUYiBHlmRs0ieoyOkrgiTQQLwePrW8OYFaVTIiD9Xir67BisfyzGczh77C5X7fqYN/thKEGUb
mcWgLTSQHNvoJj9vdf+WBQdoFvAGlJk5QPe9NWP4HE13LXsQC0FslibzdgaRyJylG8HpIUHbiLbi
wjyRhRMpF562Cyi9nv8QmvYW+U+c9srIBOy1YZNwz9wYFeQr2Ugs7DBfGjYALnFKRkfxGnkjc67y
P6bWDN0AjMAsntB9qgKJFX9ghTQBle2KFCGba4BhqzajlUUoCEdONNZJoFNgB+VRkpIxkEqA57ji
cIkAgZ6goE9am6zNadej1GOeyPtetMRKb2hPig8fQIRNubJfP2S850J6XDkTVKNVzE9DHhfAAZ1t
Szk/O6ycRYEchiTifTZ4oWIFR/fwRCdYFHusvsd6Zd5xuStiLGPB0Owi0Ift2cFndUvdrgDyORaD
IAt9OLSwAssfhcqdmz/6FepiONkeJM815XJ5LmN0nMiEmQLVI31N7iTqAZccvz1LX8OcYb6u6XUf
8sUZr0MgECcln33EDOTdnH8QExi3dy0+1ogqOkgO2+C/3FqaMkxOTrbCt9fQi3sDrEuAy1DsQrpb
xTSk+pfHwaSbvH4cPRZaI2dzEBF7Um4y2nlpITGj0sEj/1KpmZxFd160WzvMppbP9QoXL4A8nvH3
SXhJMC6PWL8qNrBu2Do6WiHFj0LsT04jHL8hqUmov6CQmkXGxZXpMu4gClXXy9kD5n2O9wBhqQUI
HxW0MUfJEACtjcIqnktrFdF2Us6SFVcJop8P90KxNjtT3LH1ZvQvBmN+r/BVPtUB7uqgoZ4cCWgB
pj8j3GpFks9ESaylgYRlvB4KBN22SXjPgzBNuWHh58oWTnKwZuiMtFCQ6Q1gqfwn/R1izEjZR/ea
46TkUnwGJ9nPpdSgalFv/nboKmBl3vWNkGJkLSSypEWQ0NowS9nBmMsY4CNx1qSg6t3UvV5IN5iy
zx0j9+rffK7fXUisnfeanfibbXIT4fdoqg+1YB7N8t2cDvrDVAP3SgznxomSa2O2V7tddaz6CpFN
c+8VJ/R+FHJ4nRKhR79UBvB6USxQiUIpks6x0qU5qTPzXPomOT1WgUkL0DXbMddDzqBjMNWkIWFT
+lCuYFyAEffGXVzwUnxjlY40DT6pkJ7zlu9stjXLIuc9+ki6bzKyKFddVDvdPPlVY5T41aXY7zLd
oIsxur6FAvtjOqu0WSDC8Et2ChzDYGd3CG5gH3cBxXzP2FsUiDtJAJgKQW+zHnWQCr5H3QIcQuRf
ZLEXYn9Pytb3SydCxo5nIs5RBOm1HZQiqLfB6l/eIYTifKgVgqf9L1x4xkwIiY8fV+gMYPwxmeC1
2WFkUWrBmYiFIXiXTMClC1AgM5bnS6H2K+1zBVBWxS7hGiIeiTybLfnH6V3Yz9jrhUSQ8sbKUUqs
KFxhziPV/+IfKjy7/MPzsbURhJ6lfmdvA0whDjyoDfika+0sSTcXo68pzvzjVIdAoI82Ul7842sC
HslxiaZXSE98vXUjZOkiaq8bP6xnENnh3tCqDzbA9QDssLcqdCRy+aCTuJemIaeEFdQhxzVqp3VM
bdm+18pE4pY/r0eENXZJKf8JyN3ReUgfD3zO607TEQZq7GPiVsvvQg5drPW0ryxKkt7ZxOcg4ocn
Akue9gxnA3XxsF+h9/3mJo+lB0JimvElOcBI2YTTnVKhLcKvGTRCO/0x1Wx49DB0eLpiRNrWO1Di
4zwu3ytCRcq0lSRD3LFpbCbt2a3NYz53kci/XdqDEaDWxOWzlSqzjfAdx+k5AWp5/AyV38Ow3o5O
ZsTukb+ta/UL/xDU98fTq9bqo/2oZioNE1M/JhqpaIaGlMp7k1VqwK0C83zKlt5lqGVTcr2breGt
a+vfXEnX+B2QDX1DFBbu4A9P6H/0XWA6+plj0zCXX1Lrr0GXxatadNcSyPZJRvESs7WxsNgYR49C
8H8sGjuW03MVmAJTFnSu4TXFACR/W2FHgkTU6GcRqEObrL2GrIERDRzPeO9zYmVj43Yo9t4WIPbN
vdslkSH/5tUoTF+JOrwbbbvvKCu3wdGTmadIUNd8IlJeREisfLRnVTMCm3ByVkDMa70uaEU3NHd9
ZQ6k5WAet8/TEq9oqnb/QM7bZCa+kwI1lk5UkmXk9CY7rHr2gSDmRUceO/1SZ7YEAZto7LOzTKZT
wlOILzV2e1S7OFkgmHo63ZbWsjEuvq3P9D8rwNyA9unygK86SesnaAglwVLzzDP3YqNS5EDpGB2T
AzyTXaer2nYmKUgmfNFft+H6avsj49Rfr0r+QEMdd38+6inVPy6H0dM3gxvb1Yozh61vwoJgRYsG
GMCLb3VkKt/JG46d8O4J3GUtKCn/lgjOF2YPLirHn9OrtpgkIzgOWBY2GAAckNDvXpF1JWVsQ7aY
kMtRS1cHD0WE1x9xeEYVfwWOtDfis/2M9D7sdXHak/W/dXVNQmCUk92Xjm0lYn/Jz28MFmE1AAzX
BczVQY7cc4TbIBFbrfF0AFOwr1zzTFtRsTLQ4KEd74cYzlKj5Wj64uuPY4UISgq0Da2xYs6F7ZLV
qd+PEkXK/lCih0JeBKy2nC75L8nGYY10vFTa3hSYYj1FB2ip5kPD2ekmkGZTmm8TrYbmbStRpISW
6yFSLWu+vUqEg5AfLRokDd91KKK6Czh7dp/hfPNZlYz9JxaY9OzOr+bltwEKB/0Qf8Yivmv+d4lp
rbF6dabOKK4ineml8gyBzm5nMMGvQCIsVsIHQubjpeA2yaFCVddCbyGR3vJNZ/oNuw+XGQUad5zO
ecOo68mjZcY6kakjCD3ng3QAGTr1vXL9qNznx6oizg2wYLANEhxd9DjN1yMdVsx34L1GN3K3WFvi
3CNwzKLFb8GXdeqz9zUMcJG5Oez57HqNIi+fMYk3AF6hDXDW/B8/epFQnStgcA8pr0MOFJc2Kyln
6eRKSP3ImliTt0ffmLkcfZEbzJCuXcybRtyEBxUScQ0RMBrFuZlkpQFSiyEsx+er4YmOehIogCr4
ATKVOK1jhmZp+Ge2FAvS8b5ByOEt6Lss169NiDn27VzqSUaZWQyr2tjffhaSFXnUqUThRHZvMMP/
dg80dDdUtjimbBumtVVljG7Nr100cbuiDSymp0vnD3+ComPPpyyAQZlSH4IRrBUbvTyT1L+VdB/s
RDz6KAZ0Uk7+xCBpbKudawliHiqGjkvyShHn0jR8J5Fr+FnflDjB+o423vEJLSg0BeaQGQCZ2Pid
6SkqI1MDYhqzzFuOCGgPmap61LW+IhIcMksrSCRoT/uBD7M57vbIVb7izcfQk2PhZ/MsCnOqlHWo
3rDMh0dxjvXCcyL/FeoTCjk573+Bf0jTQp9z7aEeww9ZOcRmcJfPAOjfF7cWv421x6tBZ1ERhvUI
zxlj5rdHft+frVfU+C7t5Ccgs21JS3VYgR8LTRhLnDVv5H8JicCT1RgPPvihnpiuWGmTdy4ZKTRi
VDXkOXcZWZdg9uilTdT4VL5J1Ov6lh+WMdHqc/hYbqqkKJERBa35QSVk3IZPMjkJiYv93qXE5RPX
E0PHAsC19CiT8mkD1kUhu4z4PU2RbcNOSqJdzDWmAOXWcq9hWMGwJiJUzVsjoe6GSCW5UbQ+3Qhl
5Eg8S+PnFRcc1ClIOJW8CjwyudH6icWk3bm/OIXArGzmDlnjx/AxPEQj0v8dCuZUa8A/jCMvcjoC
0E+i1lMlONX04IEIF9l6+sVpmqNyULzcA5bHIl8r6WoQ6rCvfJyUh+xEIgKtfZRwcED6cjgAwxnh
IsI/XS6YtCRiA9n/+Mf18QDQUnyqQ9x9G59Vb5rt+6GmlkaIW+Ga3wLGskTHpcG1tsmgDA7G7xNU
KaSz++tAABsRdKflRJB6TEzpS2tQQFu68lr4PWsdglf6m1/EQ79HEm6So61Ne7nSSg343vhXy0xm
jLvMUDVhkwjNrknrVVn8qtfyRaYUrvV56+kDQ0pjZf806rtlDCJcZCFfgX7xhtnKnYZ0rsUULm1U
R/Gl4ca6bsRId/Qvqdshx29NIAXM1G/Lf/JHM3d/bpqrhcPYHgyZLiTZBasBO1ForYHNBDkSzDiT
HMmHmA43jWpgqz8p3un5K3r9PVlkQwXSJbxbnckacOk/R0l63XNGYwRphjdjGRniDmT/TMoGO1Bp
d17M9srjlEyDh/up77aGG0R+ebMpa6884/25VvteXxvTCWiZ8dt2lm+xA/gX8BZfxhN9thO8dDOk
TR3WQuH9RmZQo19U/2nyhR14NoZUQZ2DJEUX+s7aBzBPK4x28UEAzZNPkOsCQCWzjTvJ+AiT8fLW
qp3t9vGWTRX/WwrW58MWGj138lt4qHgydgLCeymK47paVK5Y4p3AbxGo3CxiN3sHPQyhhCQPLgQZ
FWn3ffH1jSzVQpfq40g1glRp4k1FCSbXRaAIWWDLir7xXoxC+37PnQw/xIwdovYCekJdQ5heQ71t
WE165gN5jUwhTU44fpLYSZqUGwF/kAVDwBSoPNxPFtLpGYS0V2q/5EWjQbFmN0tENeEyJ0oJg/PA
K8S+s2Nmcp+l+IjrKzDowKLFYKYp7njfVDvXYZTdcFUejPLRiufK+Jn6Jj4OoQBOnKeDtUZmffem
VuYSRdizNumSk9Z6UYPuaiOol0JJ+xlIElNouZmZrwgPd48CSRhO0w/4QFolsme3AOqTPOCnYefE
J2gNoJPDPlSRtKoHpJotkudNtEAWwaqbm7iFD4cT0QmDXPAeBZ43PGNKEBvDisn6eNCSaZlPg5Bd
pObgMTMl72uWjtGNys48nAmvGlAgNXqbmRgLTTfPgAyRGNlgs1qj8GRAiQt8bVyG60fFYSFNKI4q
dTWnnNmrbuNGkM1CyDtSiPoPULcfTntyD2x5YUPsZF7WhoZmmhMWoDVxd8nkGUr0tFs1gitDHeJA
1C2syc+CJwtSyZ6a5lIcWFpfp1Xh0ZPyvxbyk1CqJKHFXfik3+BFGTflVal8udeIr3FoBKkR1Qrx
ukvzvZDoLMzQtM7Z/OdhEvia+galQmJabO4e7Na0BlRD0QcEuGhEJBMfBIRIle9GwACvii6+Pk0X
klMWCzHtI334U2i1Bip1FNaadiYUhcro5QBT4w6wrpooyttpxih9nVNuvEGWivIq+nsQXTHLk3Ph
/8Iu/XJzXERyxYduFzxGYPot+Vxt71dbi4KqbmYCXAFQw7fWCGGUpUWX0FpkV6egEPIaBzy+Oba6
vZCLoqsGO/vOzlhX4f7BRzWeJ4HcTS8VkmfwYTFGPDxyJrZXf/DgfuoP/9UOqYvise9CsdgNGA4c
Jlys5pYqgBppQ9kmWwuVHDQZdM1a9Tvs8XQ83ETppem3iN8q7OWAK+fNL23DADOJJGqlz9MR06Wn
6nAsk4JYX0OEHUr2ZWEkE675zq7WbnuY56+GOT9+Xz8a84Pnr5ByKVGszcElpe8EkWFgD9AQP88L
L7fKOCAoq7FiLMbtzKNQhnIe0xoKupovc28+kyOu9VXXpySivXOo+udc3hVpNgul3bbFviUlNVBW
ZGpuN3swpKiSV2y2C0sHNn7QD+MPKWZ77iE4pv41ENd8a4Vxc8WFVzBaART9DggspdVliRUSN/DN
TR9eUGA52e6QngHNEa/BtfoUVjaJTB26DIP4SgOAGnuR1jhsI5qk7LRXXfMAa9PjmMwiEQwI82fT
j0FvF3kfhRY/dBlmm65ZhJYq9dXonb4IjQoFaTL0PYlb3pTwtRmChOwP8hw2v3NWX5rx3AlfY7rv
fOFI9Xzz76NBILoqMaChTdhVOv3iFt3Z32+lD+iR+F5WBEiCgnHU5AQ10NNrUBeb/en4JbNShoxb
Ofu497zC7dzQf7aR97V8DcRo68vVowyYmtOLthKiLvWH77o2LuBlmovsqQ+Yki48yABZU8NxKwQ7
iW8a2mQPIswpkqkOCXc9IfwaRryWdl3vKl/1r8rHv8uGDtOwmO2zEqGilUAglqnZN7MsaHX+iHnU
2Ynt4HKRDjgtEZIUQ3z0AfOeud8ThtTMeOQ79m5+pRhbablvL3wxHrts25L6t1RNkKaOScLE9QEx
XSGIxIB61VtKjKWZ1emHfJrLZLvatAbLBzBiqPkhOKrE+eGhVFePArmqUlo10NA6QaggqpBBDYPE
Is8eWZbtnpJHTr8a14blcYFS0cAs71ggUhZqEj5jRSfXfdkunLIlH1TB6xOT4t8vho0bVQUY6drN
foW0hSvu3NfLd1NAmkwJ3RY0qusVGTXTqL6wU6YtYhRgoGlmH15wlSYHFbnSUMSvE3X4pqZQ3T+e
eohGVMy1xkCVcIuPO+QQOQ4CZkjJhZZMcoMhZiazfFCk+N6DfA5MZvjbfPvhp8DBLQ1ZpRNMmIlG
7q5aLAdZ8x0uEJ0UUaVwa3eHvFOTgbolltEyUMOMfnpNv5EnQpqV68CGXjoIEuwayRwiwwDYGxpr
gKviaguD2scBkQsy7dg2rI9VlUn598tftW9QAVI20ainoMJ/1oAGxmc+WBw3PU8FxJjgModPhFKk
xuZ2EljtEvl38WFoshEr4YTyEIgWZTYCchJSIeisSolzeJ/WKOU43nUkDPvtFilG7qKYw3Q5TCzs
SuhACjYVJsb3DOJpxUD/jUnh7ZwSyMlujfTCV598rOU69J7kGAfYdAp3P4QIsjoOV6Y49dNdVKXX
WP8IDsSuCTlhLlMztsV35CA31nqOx4oPc9Ef80RQwsoJaAsBdUht232TI57T79RbQ4kOzKc+HZw9
DhoLXySP0cZOgAPwrmGLBNoPt649xvmmWiWXBpKWW4xA+zXxGfn7n3GPy8KligHCX6DD/sfs42vW
05/DeLfFWJ7ZcfLWFtmP1e20cukC91Get6mNYOU+uM/TErhIBtfL07MWE6YYwdow2HNNSeAB+aEf
dkMwzSIa31OkviovvWl4dpyn+SaPvSj/PFbxftHPaDf6V4u5oZGwrKLRPUXRnNjUDjdSih4VwVHm
0M3S95moiqpgaBRlvJvyGL36EGvq/jxGDKLwdYBOarTjjxuBCfThfN6Ld6qG+Pye3EBVpmMIsIv+
PpJyISeEDvenRAYh1X51cA4n6JjXJKxn4Btl6sN0Z6Q7rq+QcwwuQA95MswnuqLBTdHcHDj/l7El
RaykICsXEkG2paj7WPeYLDwFbXNDEinnUTaOc8Ia5gl73qSJQaMsgSboF4QGY02r/Ipsllk06fPr
xi0riui8hi/6MbJ15bjozHRrHUzep62ciT7R8tiDjIm4OAFqTntnKcd/c+0/kEJ4FhFZVFtVlAqi
dVEtpOmSLIlCQHu/2zOh+ojcQXO6q2KeicxCilho/c374zgFQPvqsOrNqREiqigsZAeAAj50Jwpt
zJVSHqD8owMT/0uKxFSYbhW/bvMmOTiUyT4p0/jSBXYO2uoUAOkHm9Lgkab8rQUvAlsRuzjNI/Q2
8sHfGg/YqJzPKdHDzaQa15l6pQYG1GZOUpxdc8L+IjxzYIWoTUX9lF2Eyks9OY2F8uSjuxhGCkXD
Mf46Ljtx/DLophBNVPTTgHG2/E1n6xd1NsVEMSo/+V5OAkSjYWEJENUowrNo0lvkO0FySabIdS/H
vN1zomGM0vWq13fDazDK4+hpYdRDVFQixYo3c8IIDwFfVlBleB2Z55wEjBMkth20XATJdX7PTIp9
wJwnYdhcjwFCwWtnoEGQql2Pc8Uu86rh9ad1ZamWxOkBrscegs1EeW9w9q2DjqmPg4WN0Z0uJgnH
2Dr5+RoDZRUgrIXAKfXaAbjHOgd1JIJGW6amcfhY2BeyroBoG5USKb9fyW9Yx7v2P1QYLIBF7oLi
90SNBmsAVNJUOxvNynE30NkvAUt4XjaVqNru2JzhJs4VZfh+Iq7kIDogzB4zEhuBFLjtc5Bbg4Bw
W6Edaqcq9xDB6oqfNt306Ez9UjQcWgnCLNXUh3stf2xGy1BCt1kOIsXN4niIoUaU+xnbtobi0gas
t7/jQeUrXkcGsHiTGOmM0a0lX5ivzdMdrbAly3Iw7m0PX3tYXdIJCcD+Y9anPJPYn8bV2xa5w4xh
pz6P37NkEwX7oo28q5sReVvQUF0y1rD1+erD9MI9SzF2e8mzMtnma3jNYuR6iFTCppv6C1tzwntF
xxG3ck4up+0pE5S9J9/RIdMfwyUSlZ+5D7Z343cyvI0ZR57J9pb+5JTPTMNmk7I+iWCZFwlLVEj3
vnghIFIU+iJFqcgYfVzK9rD0kA5r73qVnF/8mcEya7yqeT4WEK7j962NUGjrgmwHyH9HEFBtBKGS
OtwlUgJSqo03B1VZnCg9KNSnPtmw5QMuBIYNhOGPzJvrs0WcnfcjeE2eHVYvI88VQJZo4/VEr5sr
bLP+Tl6SOUanWr4dPFZExTFUaE7dz3ZAwnAzXVSWfWURhTS095/bCcgFgcCAOTOQe+MSwVjwh1Rd
68QIeY+M16zcpaPFn9SfGNA+WruO6eLGDy5wzN5rDpoohWnvXEO5o0iBCq6syf9zkIXh7CLUm8Dy
QlSTQf8cLAUAGBci2X7ZJGtwtxil7gN7Zi7epVJoM02kY8WNx3knc77m94z20uU9D5ISsBBzvTDB
MHaYuQ7ljmgdwAPCmYl8D+apVfJQMN+nnu05VwELwT4AYaafSMa01NxUG66Bl3hE82uGU2t+qKLX
AFC5iS1g3nJNGveZW/0u8eUVo1B1Z1LfrpGCoOHRUxQKvs5JoaEeTmXEgDg7BRfH8g1c+s6Q37ZH
HmlZmXDmqopHuOkOkkbLutaXQ0tPr5Fy5j/KZAUzvyWrjPw3NyMj6j9fTty4Vv66RzhnXmNRlLfz
9bQL+RksEV3mHdUlYgD9jCFgyEXjNmuJ9ZqzA18q380Ky7l9VOB1xnzQO5lNlxx3zEJKtLGu0e2e
36Au+wVrR0euUe7GjTst6Ij9lxLLzfix5z2ZAnZuZG0WcyHfPWhDyj6kKDKYITzneyMrGKpLsPa5
GjC25VxQqUY4SpW6yPYHI13AhtKhbaY0TXFs62OEFnxbxorIcDWVctkAOZ3CtoScDLCDt4M1Ymh5
Txv+q6D8ibtiE4oezSTSrDRGbKWR+PCnP/LrbBdCoT6PEcUdKnajnJe2Nynw74X9RccMnOHBDrKm
C8AdvumheZu8WtJMaUFTUWiFE7qRPSnd2QsK01cWA/jyFlAIT6fw8KCVt3YcxtXnXEjZ7RjXvl84
6lMH/AwtzB0FYU8jo17McT9eoQLHi3Qs8MCOXgYZ3P1Wcu6EFLzBQ0EI5ztqDqjTt1CcBRamvnxP
HPmjb55pV1yAisSSAe4dLtQpxiEGQTvhNQLfTfJDreFwCmdTmqBD91OrjqDCLlMAv/uTXBRUV7E/
4MIYQJ60mC1aH//oAF+szhCjN05vKwvrAnZ2e2lx41y/w2vXDVY1nK73isCSY2FaKo8MmvLHh16p
7l9U4S9mqqrSFPZ9PQrIptbLjq6gAxNZOgzW3PsHt+1mTXNTEgMxp61ljUYPd5Y2+vgckA6Lexqp
N+ClafQsDw745+qGe1r0hLp689q0vr09nT0PtmkSzq3ksn068WWOAsncQtfj7mD/HqHgLrWC4mH/
To4I1kWWlyiXnn8DrWYqLeRiWKAjGgSRet3s4YK/4wXdKG2qakDXV8L87kneoB9Ds9BYCCnj9m3I
hveRzoDp9fINqph+VXzGuMQlpydhxQTekoh/b+YwfHF3sRvWB4CjmJ5i81TRv5i7iEs2pIc43i6n
3xQeax/hpJAqbDSqx7AnresRu9qbKQRft8cCc5kvF9vEi1jRKIJaYo8K1wXRaLFRJCNOIczxsPw1
581q520cyHgbA316nQ89PvPIc3ooHEuqVdo9rkh6bjxovy2AGt4LZ+3LWjLABrwj+H9T3Imcbs7t
qy5V9UUxXnFQW/7/D6HyD/8eQOLMRG+28QefsN9AMmoXFnhk9odtIBepuGDWKMBvRz0Bt7dg+wSS
51T6LgE0svNxFf5f/NuH/msDNCsUK2FCvkknmRzVsY9ow0A+nIFnIitX3Aj5HnlCxg6fEl3iL5UR
lvrSY529cRoBIe/meh+TvHPreFB6OQ7Tc/7Ye0tu5Wtic+IQ/zzsZLfz35BJdw+KIzkEVPJIxTWx
8Ip07wUl2RWvjC9yxNZqo574+xh1mAONNcRxOjJ7p1vOzaYFMkDnhqKeEpswr0ugfkCc0t46r97U
Uv8neaa+JszP3vjx2mhxmwMSa/LTKP+HUmflxyAUu8vCrzznTIyz/MjnZvXD0IZy34rrJ0aY+Zpw
EnNoEgCdEEghon54KAO3ouEVyIXTC5+30qc1U8zELveyfB0/Reck0PWvkS4zGbzI1SXI18qrMNcz
cAoB3GpmzSdwpjnUrYBBNodAYqdvrAFcpgngFT7FF+QrsgrxR5ScPpHoxKdgmKbPGq345HWvoKsO
SbC7d+Pjq8OatIX0SrH6L8KI6m5LDmN3oiuConicutmqxyvTX4LXZnqBk1i3ShOsh77eOI5ycg0X
osD9bOwlVySi1BKL8e2qHBCCuNTMYtNvi9LUbmEdnw0nDYlFXGFZJB63SUwfJSSC38oDAeGQ116U
KIctBSVc2PADaQrcQrbDQ8H2PxZQoG0/EfCPMyIth1kDPX4oD/FqGkA4/yHTxcIuWnx8HCKrYFj4
SMgC3H85VuFctmXyVTUl6Oc0HKkMxXpk6DQB+qcKULIgMSr6Mexwil0XFZH+HGNM2gpbgcklY6mV
yDDAdW+UtWbQtNuwalPziDwmbCM+wAhJvNgPgE4/ReuTlB81NzZM88rIv3yANktaJHYdC0ZraJ21
KVIqiaMELPQDIny1Ba7kkXk/dnL8rgO1BdqkGDj+MnhyN5tb9/VIK/dgqHd9AGu8VYiR/6aDKyKY
H6vfU68ymyUQH/1R1qqrcW8G6e5Y8oJ+aEzFoE66ui6Mel275kig1jGhAeNaS4QfSod2//Dpy3cn
srTedqjpQ1xzNo0jIdnEymuz426mMQMm0X+dD65UWJSoTo13AGHOw/03soesV21tcv+OGFmD1LwL
rA+sq4e8N6OXmxAs2eowR3QM9zEqBIfDlTWX5t7OSgUJPvX22OdWGSXoALCHxMZJ/PPk7yP7/mF5
w2ytlIRe2s5Gsu0um3Xjhv9D7cWI2MiRS6BWOD+smWKBLBQvgrTuJEAub/7QBLYz5bz8gbM1NBzp
csbxi5bgZJEbC4lHVH+VMH//LxsCBhePwMKE5n23o6EMw+jld2sg3V0zbb7hBSUY7vHYYwp7kmJP
zB4tuXTMqm5+RoB5Ne6bF6tPZIS9tq6VOwjUB7M+vNO3lKKLXqdU7vEX+v1opj+5i8tW+92Rw4yQ
GW4kF4Pf40CMAOpWIGxcsaRhNrmnYYlToDxfB7AG2Yb1z0cTsmb1c9xOMhJtxLBwVVbSDVPeXHYp
c+n7KEB+Z5a/6RPzW2lZ/a7CcnCWeyW1Ad5V/Q5/eKhZ7/pRwcDF9WL5Sf03TzKHGUVw02dTIujV
IoiVllEVC5qfw06AyH5uNgq72bOSA8koIzlUNMsrquUs30cXnw/q2UO3gUuPnuRFXRa+9uXMyAcM
CM2JrML4sdxBDzxsG8bZhmFH9EOWh2uj/APicjb7ad9toi2+s6hRC/SJiHXqVL1MccxyxJDHaVD6
Ehq+X7qFnOjWrtTZTELf6GnHpbnRvhbsfffW9UiKJWQgzY/QT9o1V/WR+2qGgjlala1Z2yMh+yfQ
91vZ2C5/C8n9PRzbKhIO4kB0eZh4knNDPOKbWrNBIGTy55a1kWCnYaMdAQ2T7PuKR9Ke8hgW9qUS
PQCAnowqQ0erqdTATi1XJh4KtCdaZ9PnGJik6e1mhC23fTbSc78yYM6CNd91De/WCupwuF5HND27
EZVpc3rjzl8f7B2bQBi4m+uSWfVEOb4PymNW72DFj6NrMUY9BBLlUI/G7BcGOljaTNf8qqzH+Xeo
q22yhRvyjh9n56cpL0ZB/pUI6FL2nyVx+8td1CMn1XW3P9iIr0QLjHGo86YZ2bQfyG6ZPRC5LfDU
WRlD4f+I9uqmEG8aOFrStJLJ9rpJs6/3qXPGqDmIXkQEYTUVVxetM9+GZi4sfpBu2IPkzVttjiNd
72Qs7ACk2iDdiWBI6wHWPNwKOanMdMLvv6KzcoJhFsyLHASP3Sw4EINGcHsMa363E3uyKd+FPGDb
osu53dmhrwnzlE8sAwHfLXnOMJsS+jxbVq9nFea8t+uqpylzqk8IzXeUyAWUiafSIwHh7fEfVIfU
9KF244/Qkjgh4N+VIuV+mNJkbDtY1r3uJdIbvPBMzAQ5C2aykld5BERUjgmqHa1HDGPumism6jgw
IesmFwAz1rcw80nsnZOvOixs74n1gLim1qw2Dqi3Q+5s3bHuof8JpkhD7JnxmBjy4c5YK9r01DtI
bPMc0coqfVldpmMXEeDVRiggEweS9QCBoLbLCXaMD0nQxVBL/NPJV2gF1AJZIybt5QYwaUsw34Se
qhWq1XcONgh4clRzIldPeud2FFJOch1MXL4B9GflRY8kIzB6SVrNwJbGjM8s83p6Kb77y3vOui/g
CNzWJ5OIUNZNSlUiQdq/FhXFfwSVPzYk51slhPryyFP2ToldxBaThSMUNE4yMHTPwI3Uet0JxB1C
q9S8hqsRrfcaNH6bWAjYrc1ly0pKerSArkMch44jcUdahcYNjU9m/B9TScWpPo6/mR9gMxLUAAYp
gRdTcaPftjyLo2mPG9n5gR4ytXfBUCDZP+rTZgJSeLIt6Sy1oefCmoFAPBq/n3onHNXs6w7h6H08
fqQyIobTdgpIiOUgc1VUFLcwus2R1z3U8uWELKzp1VxUy3drQeAWad9dfGXRpB9bFjrZTc+E+UGP
6LyvkfWwMN86oEQYvbqAFOlXpL2YJhTvGQLE7HyLf+uwqZVW0l7oItfK1zCKLIuhYO1f6qy9CEXM
KBRjAsyc/6RdrQ2KtbqNeQPTxraDdQfP8GrqPhEeIze3lRRWDCU+QD1bKbLKKGG+3Y6Z4SSySaO6
CDJMiTetLkvi/GXsPCw2hcWwouXqElcOO0MFt7mV3JMKaTxJwXc0nu7Usz2uV8itj5zAAQIh8ATT
1/6mdOwjkVqDC8YEmtf95HKO2bw08AmdgMvJ6b6j22Yguc6CDQsPb/PDIVUb5hp7qFBBJMOzz3xm
PFKB+xNkys9MMu97mp3Esp7mGDa6gEB/PcE3Aq0lZB9ISOOQdf1ScyklEWASDmk7JlvjKx4icfXB
G02VO12cimYAsJPGYQZQZkwl1lMBLMczEHadwNh73Uo1/M61E+joQSp8ytqevB2b2/pGdceXjJxm
hhZdxPHF0lhek55DLsUagUWdPtNS1kq/FwsDPNxRusioQbxqYfVb0gcfQ3XQ9m9GQQgLa/jkKAkw
octjjKI8c+CdsvXxf/RRHu4nhnDirlNksmVh8ZD0Bi+RXFd+JSGENxzgv/vFNwb1BfuS0/2DFGtb
WF0sHS+ZKTCR94llbVEbCgbzJu9dpDcWZYhABpj3U7/KTv0oo1UXZpCLyERoeNbu3nCc2ecgaN2i
+SoMlo/ai6QipW4o4A3m7R5E1glFZ9vw0PyTeK8BYCZEX6rf4wcvulja4V3ISjGZGZuFYBcnJeFO
R6w4oi8+5Oz2Y0dYRS1j2CGQFiIQ9zxlfZxO00/MrlOh7FqXGU03MICOgQbCUfYuqtg2o2fiEO1p
dYOOtjR3WGEWM81+/4X7qSBl3RmKDJjLvuBSiaPebW/Js8RYOxUv/hlNZE9/sN4uUKAF33Y/E7oz
Ah7XCr0PXy3hQsOugzGkW4PvyEB0PVLu30Kaq7hl+oTmDRBNaVe6iXCAqcG+JevjGNeuHDM0ceds
FoMjwbcgxskR+nb0cbhAoNvGjFr7ljN0pFrlZggOp5XqVZAaTZXl9CEAj0O/LykEg06fLVhb4rTI
mgzC8Gx6U2i4M59/aypVTAlDSrG5PCc9KeL1aeXfScnqYaKygdoue5NQ2X9aIWjHjb24+XqrTxb5
ixBxjlMfAbiE0PiGbovMIkFqkHVN9Ged74p34/N1b31me1KwelZ83sxjfjjcQnOtWDsYGlIcGwYw
YpxXxaHhQerw5ZciDZwJKFvgAGtyUAZ1cIiHVp8HIXB1vlqeUxNgOt7mm6PZ5MTMJ1ozPYXrRMJO
nIHnfRIUqji0XdntQFq1QOeWDRauk914eCk383465B+aLWf1rqGTyLGvZ0+v1fZhFL7FUHmB2HEx
hSpUKYEfMe+HgHVvqfFuIfwbpSdWIlW8FW4giXN8Xzpfy1ZRnX7OqVlYSH9SvNRamN+BeBhuPrMC
ZaikCnpVHi6fDzQc8nZAohEHOjigbYVe4QTuwp1Di6dFN2xvkx3C5PcJgW84F09kK8Noh1nx9adS
6dWHC6cOZN56YDr6s87kYufI5nqdNn/WeYkaq0sFNE1BW0xJ4olNhei7BdqFN8DFFvMYHkfJmOHf
NJCNPatu01lKy6PdOKhJbHvWwJGOTwoy+TkST3fiFtxxF/XreD03vqi1sZGYn23wxEYu/YQH4lAA
lQDL5CHk3HmJi3mhTIJzxR2svqIt8O7vMF9TVi05J8RusCZ2LOktM8HCL30em65sXYWEUgkqB1/F
JN4MJSlcU5mEg52DZ3raOAmlEAfjR5lLAIKhuAtWmuPnarARY3OSfqGHMYlUOSw3pvFoZ81sETA4
O7SuKzbqPl89Tdl/0W352F0D+asKYtFlAZb02A9ev2Jm152EoagEZy0h9t3lW9bODNXRAeAj4VIM
IiKZv/ec6Za+CzMWcp8AGl/sTNxsy19OCPau8wl0Gx10PD1jOGSBcEho5yHxJZnX/KygT7QxRHiZ
0l5EaomW3nkMxhdcsBOUgLjKzgtVwwogjoYjNRFrF4gflcnilPnMf4YmUNdb1OrSkLEyOSdMP+AX
viGZJE2wPtNuhIoZjPmhKI5QMgiXY1UrucTAhPhKCWQX2zGqcYNYGgESj41CUnX6mV3+nIzlb+9/
L2/qThoGCkEaQhl+HYFDn3vtjamn2PpGoYnUOzNnaFJg6yu5Yts5wE8CUe69jbqwmCLXLFEbiU3E
ydVSYjJCuBEryBQ6W1P/A5M6EAhE+aFFiIOJY2OBwh6x5kTlW9zmCk5tqBaKSY5VQSHOvJ/MIC1+
qwgLSHNGIksFhATxdBiYQtayD7y3VUu2G5Pem/IXBdeip36fYvWpf0ILqLWzposuVp+FWLTzDnC7
K35hR/eOsFNCu7P3cVJzKWrGrNnYRWhvR8YK/ezzEFQXEZDZ/KsEEdYyT2t/b84ItED9t/NCAr9F
MDs/BUblmTdQFF4lkEGloboKCkUNNE8wvyN9+NkiVprFXyG0xFcnrv26z6oBaAfiKfVBBbu3NyEn
IAZ4ihNJst2EQVpYDQnZjDDeaQld5BqyXRqUoAVTFZ8UjiSSiNQBhiGLQOw3fSU/T/qSEGQoL0L5
yUgj1WDvv0U+/TnS04VRhr36jylXyz4XR1WZCasEK4Wt3VdLFgp7Lcd6dztF1SHBFZtehrYMkn3b
OTNxWwDtJ8W+816TISpqvY8+kJvAQrMCJZ8Dd5PQaUA/mVdFDnsBlXNZBi8b0BNugGK4eCzXmQ3o
1w/9xaLwzwUBs8uGVOhsw+dYcg/VrN7Z81cbnYvO0RshShPjTo0pYtbs0JLRUohhm36taDBuvktA
9ukugsOld5tiikbiwoAomMEWolRzZkIZTC0OniHG5yFzH7Wb6CAJCtm9cQvjZMBn9aljBXIgvbBl
6yeSb80mrdlbeUlNPYZ95No508DVAk3HOtTyYoansaOFdUd51pSq9YtE4h3lPSaSBFNCbLFqIOwh
6CMODSla7cXMQLrM3Awx/YWtMFKJNQwvM9YXPvwZwpeBO90GVAqpD+ZYJ1EO91lSifkBs101fRtN
nQ/vWAE6658HqN7lqCKhobBJ0Q8leZHmci5gQ5Lzob4Yeyn75IP1aijrGx3EjSVKXT6eodZDGjQb
g2pLZOl0jzDSGAgWktuBey1D6Y1Gn837qc0dIF2Cfd1R8a+rVw+hrrFqq9E/FwgiA6Xu5ZcQpIAt
Ndz7yOmiMZNEEyr1l0qCQFJfSm4/vNoF6312At+uvzlHQ8G/tjqA/dYKhWGTP0/lvhSW32/MJkrH
73Gg2sKG3StXsb0irkTGVzgE3ZZUafc7grprOozEtpsyYGAt11iNhwZT5qzppE65b2ece56Xwhr0
LZPutP4yvP6SzbWB5TtbCu5RuolpOX6RN9sR7/MYtgXteNznjJwGtFc4bV7QS5Cym9lsfrwun0gM
vMpVQI31fJixC0Sd4rbs+ZU5RJu0JTOa98lTo3vmWce7FDZdoSX7FFx1QjphBwY0DJfM6a3MXjWC
a11E98TPkdTRwWfRwjxtjuu7ffUJqtveUDSh1X3vAd0NqJRvVKCpf7vxpXCtjzwkGew8KGIfO6XN
XjWBBgKZaCHGQU/gz0zntgk54Ga9Q4vohKz8YhM+oYl7MVeCg5jyvwKZ4ifBDyuY1nhGHwvUed9U
NkbICInXtFriQj7Kmm+jpOD26wsYFnRApcvfIAWyQhXMU8Uovoj9yMDL+JeSGZH48RYd6ygLznDb
6e4xd15g+fv542Xh3rCHjcxtAAnLONSXwzkkVIV7qAfcNWRP6TKG4uQZEH50hbhlMnpWBfgc5/jm
/zYOzqKC72NbFcQONmbgFhW7ccXUIRmqCMsWfhpTKRZg0cFOaG6EylHhv1qbvTF04hSUgDJ8fkAX
F+B8ZzchlUsGg/hD+TGXjtXSs+/bj72Nyf1befT+Cfp1PGmtNywn1yfbr4V+oPunQyeIi5xd299x
wE3KQufngjxBgTsu/XptofukCrXjoo+QfEHGmMhcdMWeFVKTv2dHxMKJ8674AHldsBSkDZtG2U36
kDLT15GD7FGMUbHpvScFUFzi4uRw8YMSdc5MRSIizFTNdfhRO++C964XE2IFlW+wO1yafQQyjJyi
B5PW9tFajYNfSuWD1BAz6pnqN/enruHNbWIBAExrlD2lBdLSxUEwciJFlmbgELjAWZZvl5ChzRFP
7bnKuNKV4xOnoTjlkcTPWk6MvDM6Vj39AX7KRlCFB3wAr+pk0nWU05m0SCZ9bPwYbgzccUU8qLI0
NOQfsqJKPsMTOoz/AnX0CkHJHtOLVE1oqzAD8y3/c3en2tyIm06J4X6xtmn1Zf/690AFbPiSaBRd
Har551mLZe1YHmq+CtpHTj2I5hJFDyABRBxH6YeTa6C49F2OZytLyjLTMId34XE4wxN3Ot3+1DuH
nW7XgMsO2DVo+tyb6B0ilz8OFyIj2Xo4oVwZ/aySkU0UpNod2fsnGT3VgPToQwN3BuqcK3IHSDHw
xuz8EXPy5n79VCmRBJDzbNJgHWEyDLLBvMejvtHi0NFltXcBSL7XcaEduqd6vNuzt0NDxDhAydW9
Dx4rBO/qcUtTUOSFMOLbe1cOHIEQutBtiZR2fm1WoxD7qDersd3xCdtM20y6v0INPq6+Mun2uTNx
qNAv6+vNJPRStVFiIwkesAG2mUF+0CSU9hsgkx4Wu4pfc6EmElxhpcVpbXXOxQPFBXDUjZDV0PO0
iKE2DFIBoXLO/xofx+o+oaU/edxdbJwEmr0lA6c/llWEFGuTiCmyaNeMUkZ/uFQAxWrp+p1P+/9H
822ietBfclZX4dgvBKS1vZNqMGQAR/HpPsCg5asP+df1I58d6xxP6rzMdJAiDruTjeaw1r4SmKLg
FYTR81togRE+4ea7QTFXi/4rb++Hu43ZghEwMiMmSRPQyH7L8d+2d4BPAFvVXmmdWSUkFnFjFodo
De8mi1a45t4hi/m7bHA31H8wciWMx/btaRQNsYULHeckE4AMY0I5qvto+8aOXGde/TO5cSZhqS74
2J6rcbUqZsMfYjFxcJAMUZKwwYBlZQtIfWLiqfgsCPPlTRzh4B3Epgkd8L/aLeLaUPjfZztiGIye
e7CjWo2tpr9+fw+pj4AK44bGbsxP93GVSjUQy8Cl4H3ylG2YA63ElDgMlfpLq86z1S6Lndq+RYtz
mactVkICsaZBwx4RolrzfOi7y9sl4t7Ft3N+OC5OaYKxvUG+JhXIA1DH3yvTxoPqmW26DUHScxCm
eXuiXL6/1ADsH0hUop4PB5XfC4KttR74KaCnaVtw7ZJ5V9a/Wp0tIE9jS3hZOm6AEmqaBlhA7jzA
2CtsU8nE6dhqE8d/BqXuS4CMSl2jwPl0/mVQiiyCPCCpPQjfTsjlgt1lfYTjZI/tzQlKZh7Dg7fb
txilVX1RfgLztogvoPXf0Hikd/DPTt4cdLPEZL/nlYiMvON4unbQ5oYPWMAKVaKKuRvneme8BVYv
aRMRhv3m0cODD7HlSSxXmqv3Ac7YIjPHKbZatquE9GFP7/yHCO3feKZdh6WOdvtzyVvomVje57/3
WjerJPdJqodOGN0JJPpR6xKqIISvloAYmKPHjCcO4ZK53t6uAJlOJihYIfT/NdM4GtVCyGYmYjop
SdH+woZ/UKTis0+R1Q7M+8XrXG5tKWOqYHFTgFvF06s1VvTsBWcGOfKU1qdi5hFo2I6moWIYj/vk
ITd1yPwEg4qzqETEEYSQ5MSvZ4tByiVNf1IoLRL2dS10S99c+/bS1n7KnUkJOPdqxQydxwyibfY7
VGMEn9hSWKwdZ86Cdnvi9c+rYlUF8a9b6IWoT5sry5yfF7N8kt2RGer+qOoz45JuJQmDb1lbmsvD
nrgVqObBuYiS08wYjANXrtKud+SbCwYE8ajrt7oPcD4P6rKdPG1h109VKRME4TKsidHCM5Clj/mF
m7qdbcsBvYGlCVkrByTkP4lKsfE/zzm84bLUPOeahJyFbiFBCk0aOAfklDUJ+xCIkuPltpRv+jfz
RJE7nS806rIfCHThpuLIBJ/jlZBncavlvPpd9pySceOkf3TZkoQxBcjN0lduTl9R6SAuo7SFPMrV
jt+/qxTi5mKLar32rVGnWK7w9aMEqHPhYdERk0s19cLdU+SkhUCbCvUNy6kiYGFbwz2fj26KJ/8K
Wov3gkIAacozWXrod/4RHU7XJpDu8nf+MHRnpi6lonug+Sa6wG2Y7ESWz3+OCxfWHPUOcyrY3ymI
MRICta9pn/sUwGysFUCU/JsMf45l2eTIXAAhu9I/BVMIrtKDFCrR6Ku96DEVSimx73PEhj5HCCw7
DS2PPU1wuxChpEzqDUC+ne6EPKge3dLoMPFhqZwF2kVhuhgfbDQdnC6pMNU3soVls50yu68MGMSg
y+S+m7Y55K2CQAC1ErNC7vEiyXj9vbonHnTo2RnO54BPqnHqxbf/Ls6ySMFiTiUa3cg9fSLMt+v5
LXMV1jdtfAz/d0Kvb1M1lqsHF2Eu0FSBL1e3O78mo9xL9XZXo+/pLfIyrb8ja+YMUamgezI3D8ER
6xoeMabxM4SOwxuvzEoNoi1ILa4+q7R5BtvEvTaC2Gg9JkMs59+3v2rRlIOcg8GKRe3xRZH2qBKv
ZBd7H2+2wAjnYoqZ+UeSJl3NvvLc0NxQEEA73FVDFRDqwtFILtv00iFIJ5wL/NSLuPfpyx2dCMAW
dEdEOuEemQX1kc2vKjaiZNI+8xbALH+q0XBK4BW8ka0/5kMMmTzvHbyXrLU5ghO362KBwujDUeRh
n9pIydmZkhjQBkQGwYJVfMAmvVxXkGmgCuvM4unoL0Q5cAc1l5pEHR9RqPcTw5lJDH2etNG1aZJE
aGGYH77NEo32rzlrpMQa7XA41oG4WiarZRxbj4d1mMCnNbVQBHGpmUpZOfkV+qmXqExIiYqeEy3Z
uLmyarXsLo0nHVmT0NLMLeOUYbxYRP43PykEVOdr9DtzcJfrTDw5tt7LMmR0ESXCERDLUBbGFDTC
ZvjevJjcG4lXwTqY7fC8oJSqJyVgkIIIrp6r9RU8tiVL7LAmQaLicZg42DB1Ew4T1iOc8RGNDtZv
D3CnvqLPrdSTT0C4JQEJ3RpVyFgWGGbsi5BoPl17zn+xt8nt+Wl6InQfrtf+XNJmT1xAqXF2Y1Db
/qpeYdOmmJaIEMj7dT1GHOmSDKPiwqLcwC6Y8ykkcwnQwgvh40Onc2m+if+fZCFzGHh8qZB8LbiH
wAp2tQ0Jj82DAaD0Zsrz6wKuQGgL2geNpG9XiDza0wkT+YYXh4c6MjOt8/EqONxkHqExipdvB//D
b6jl1oR1nJOteP+uN/jR31DQv6R/x2gvX5s5D/ZKtTF8m5uXpQRdaHXoZ5UpwoPsz5VwL4cI3LEg
0sFrVv9yWvC/a9Wcu/gF8oHbpbpZYO7xM31EbRppLVVsmWqK69LIqBJgn/PnY2ELmNqiNRAO6S5G
7DWi3QqY2SYVO64Ze7AV83dwZhnVFRNrw/egMmtw8fJgbp1uioyr3Vf0rx+32BfQmODL2EazrpyP
HLdM+tueHZPzWHyJ9zvBwcgIv2SmNYOUlDmmKtGRrnVT4CwFThzbwvVXNPsITHnZ5eEIX7oGqB3j
JP0zyFAT30fT6pxZvUo5pPRK9Kgf654l5SXpzv+q+WvI1n3NGn3qBFcatMIKFD+7vZmiJhhWoy8s
CHUsFcwV3MbpFS0rErncfb6dPF31IX88AdofzYblbe6jq635drRJGSsiypFNxdMerxZ41MYRzFbK
qeO4RJliAyny9QNVimqJO2n1D4O75WsrBDLT2gZ2mo8abDlS1vRmzmuiq/vZSg9/5nDdhkYFZbUe
XupAQ61u0Vaqd85VbY3dqIVJjKmD7j5uHy+xBQjqpwDb9LPul1M1lu4xLzjl6n5O866M+Idbn1dS
EjyX8SF4wa9Lw3hI8XVx2JxbU/VduFOfi2DkKFeFyPDYEuiNgbXag+sQpP9JsEc0Nrm2zweIbVNq
K0T9wvCG6pn54A/U5/542/qXCdzntcmMSfZj5doAb7855Vap46wO1lUhEzlHnSypLy2nOa34MamC
tJu89VTbI0bDh41mF2wCmYruNJSMsJvCBBZOIqrCX2cOsYJahkI0QDmO4ZVm92dsgvM7WqQ5Za6n
zvuCpcDJ6WIQvQNjrn20bvpt9awqAWRfvY37WydOSMprYB06my76hTzxo8zIgoA9InCxQqY5OKQR
Rywc6P30u9XmFlCQTv3LvA8OD6tps7jj7rETDsWv9zuovyIAyUuC0rcnHQ27hEiUnyjr7b23b6Ox
jTgWCJkk/RJ0fZ9HFJUnI3p3yAXrsxA3QcozGerUNE8i3Q0Ui1KrlH496N+3lUR1EWwwCGTPYAYD
NweECe1oz4K53j0kczMoSkv30TrBRP24GCvx1765FEFwZvzGDiCNp/DqNF5rlwpYcVhLzgUNeAc2
n3xSm/pJxQpu8qtaOEfT0bofuuJzsipGhlaXQNBnMQ8gwRahetJ/0vQLzChoi8Y03UWpxVKpOpkd
23AmUYu4R0eKXhGPrAUuRxLSOW3qfMoC9PGWBRiVWgNlNFXT5pY7eHlRuHD2tjF8zqMXhg2T443m
res+avqwmAVkejaUaRB75jLu+5Wl4eroz8+ppnOg9eLvHsVyKTdDfWRr4VYzCiZxF7Y3GlSMvq/3
8OHIox11LUEWIl7GXkMTw2H0w8qdh7+XeVyFYRGQwJrTgiz3mgHObeD6Q4rWPiYEvDui2qwQvckS
/RqkVDfEIhkjdmUgjYBYBRB31OgMVW5HQU7HkFlIR1xpqpR3qgEnBw5pC2yzq2AlCjhIa/fT2/Zk
6uQNdGA76h0uL4R3bW++9ALsk4LEZTUY+PhI7PIF7uGuEg9mXoYcz43y7UO4DG2MEnwTvVZCqQnI
oY5ZSuNzr7XRvUV2cTJUkm29SHcx+Gu9Ulj37Z7GZLsEeFZxjfQhzgXsflPTBDVGknhs3D5vppuo
5XQLOxeai/ZaxaIyZ22lf0OpQUnPh0U0g/9hvJdTN8tspZj8NEwXwtONN1ARxAQQOB554Ad9vtwq
9/qjZcoEn/iGaBzIiZJeKhlmCALi+qYax04bH5+K/e375BjlE1Qm365SOYtdJZUFJWVfACzGZoYB
yxcIRt7JZVTG60pA0IDbE6oV++sBGj96HKr52FAaoIFog4dalV/++OaZxz+xs8f32Kq0KY6W4WpS
HWUCHkRHEjuArTZ0H5Q7RPIgA5KiPoKU/kgi143jJ/qf1qAH5L2OhPIJ4HPywcL64udZioKjvQYU
ht4fpYjI/Dbfhck0mmIXKgkbVKkJYMnXEyE7CWYupoc9HHAWDM9+MDQMn9+LztSjhTPinp9rSBaC
OTbnjQXjz3ErB6G2TI0y+wIHSGxGawqGPO0LFidCWpud46VJKKgb9AK13R4zcPHaZ4x8JYy7zITS
zqNSsdMMceKcl9+bom8lsOmOwwB9lNZ4l14lDXZPfA9kLQeBB0DpR7Oia1nHKruSR4aRtyYPHwmz
wEA5nT5bw//zhO8q4Ov7B6bHBUvOxTg9MaSW32KIQHp/2HiR2j0JdTNVoZi3Xc/EYYR0ZXxmm1Ms
4CVba4lNjkfoILYrGisBg8T248OntsLQ8LYbNWfDqcJ+8R/caN0R2AQth+yM4rAUffkk61S13Cs+
/XbH5qoS9YFk/nNrxXc69ma+vRH51H7UWxF1lsVFSAMDY3AiIgyKVRmjz6sQj/nlWk90zfs4ZTpW
BZ0uLdZTlMS/yAZe8ZBZqz7LONqOnNGdJ93yxsiBVX7HjnbHYlEEAoycTcjA//+q+DF9gnFxgLHK
/QpHMyHxi7MLNhEAv7c4YGM2x4vX1R3XWw4J58T00KoN6K6eo7R0tB1rhYxjv8ALRL2bZOSOlToY
QFDzPq7JJX++Wfaa458bxH0lESkoEpTZJvFBDsNh05GtsrS+i3AVr74X1lmJfIslgfWv8lWFRd6n
vRhIwPPg45+egfGi1RE6lsjPnTO0zQSnumLi8zyg9QdgwlkE8hn1dBw2Peno8IFIfL5lqbrGMO9z
AMHuXEXvjZtTte9YXb91u0uCCoykR9voD85kxzZRs+0OaZlQnKlo+vjyNR0HL8ZviRJ5NAeXBRDK
1eqPnx20acX31P7nOav+oQ0Kq7pX05o+vJoaKXO/CRHm29nMS72m2Hd3tieK9ulXKD+wo9yhZugW
ddDEN/GdaoSJAu2rpesE5t8uI+rxydRccyGpZsxbRU/Uotc1iMoc/xWafJkev2+mWhn0XKKk6ILl
Yio617kkWUr6IlImXAyMRAO70AUU/FZTzvGShbdecjR/W8MykqcQ3xKTndw2OhljwKV3c9SV63C1
/dMMc4qCwjVVk5F2uvM99LA8CjLDBcPapFS7xnTy7wM05b6WRb69Z1phrU/kbFuBbbu8ZEQqOnk8
QTKzGs9AgihEMdoGQ7AqiQcjxNzdtZeHvXr83J9FVYKimg9ZcwgaXrm/uLdaKZWFDcQ+UZATbcKH
VcmzXFUbehmx8NPahR+1znu2PE0z2wd2OQ3jQ2anZzKKY1uJzLEvxVITiojehovDgqtCN5VuMehp
StA/FNcqi6oSia7dEW/hLvsi8vPprcpVJJ28aING9lAa8q1jJr0Kd2lYpkrgAyyxLcbEIo+r9itv
gfCdEKVugHBEPhFMMoPU929jbcYHNMONCEjctK/zGD77fxR2Ysg5p6k2jZRc9CQuAWb3KvzZ5tUM
3XA/gFOV572yMHKSLDOk2BIAgoBktF/Qnt3VPNEzdRxarRb69mevq3w1GMQNo3O8pjZhuEDwnoIi
zzEFCQIP83XT7wuygYxN5jTAfaQPizwYDvoLP2ktiAXyW8PwBfLi/D4u+6XtsB9oK3kkYm00vwud
vujcpMth7k+bQYspRn17GbxJ6/nfIhUoaYfkRIuYwLeZotnPwaekGOIvqDRSJKEgxfaukEcG33nA
sZFbEZkEUKBJxxNJsZDeXo/lepRRnuGhn8Ml7XWKv2kMsX6nwmc+bhH+o+NOteQl7IPUYh8ygJgJ
ydwMa2WQ4b32186QcKg05AZe9sAeVoBW5s0sp4pvyx15jisRWcgxfXLR8A9zCpLMiTo/3Wo6jytu
BWm9zqANg6T9ghweiApiGuXlkFs0ij2g5ig2O17YM4pcbC277iwM0SEyeWUe9my+ePtmqIi9Xz8V
SBJ9JsSEEEi8b1OUMj+QlGykccS3xnf19OnayJhVEC3jh7rYCyBmBL4XK72BG1x2GJEOJQtvebLY
pZijBvJ8aNPyOIPLTHi/rTK8Uj2j11mPoIuzZ+Q0KtRkPm6OWLH9PWyfyNZJmOlA0tkkpx0JmpKN
BxtQQi8JH/a5LJjhDrVYTFbYN32KelmDv/4z/73rF49sQ9Z/66utNng8AhWqeXln9Sp8aCpdinR/
30gwhJf3yrRyHXHUSa7X1nMYky9yPizsA3D2JJq6mT8H56+Zg4AR80omk1rfm48Onq8b9jcpBOqD
ajHgLVL9BqKiAB7ADBmvFQ/paq7YxErnurQyDEqKoUeSSypeSyHaygTIHoxS/cBYhPmHoGYt7orO
wCm/HSithsGkipvtlzr+atHy5EVa0Cc33A3nXsU2EttI1OKjfsv9dUTKechfiJxDHJn8d/gQkYQM
eYcqpO2zPhic4it8XOlMKJnx2G/qDkbtkTLb7/2RveLO8VT9P5zCUPm9+3GaZHBIf8I2NPtwjWzV
7Ox3MXNXzAhFWrkCRIqSe056nYzvcV1VGFtcLRTpRE1L1NIMYqlnRf81uPPSul/pq9pmQ7D0xgTq
UmUDvSW/4gWWUjJQoX2pMHZdX0ogG8HEbLVBoRShPSAowx3DsuKYb8KkME/Eo0FGhNEt2Z1bk7vs
GfMqcr8k3rIlLd2a8imjhe5BIkifBSz4USq5GYcuTCMkdnpaCdcUBAWcSVto7/Q1vt4QM4UgvH+9
Qd6lWD+fz4FOdGumW279joSR8+5PWknsbiTqKkBjQMRU8lGcuy/D6C10lkj3/xcUN009XuxqafQR
vGxqxeFfGMyg9HAkTiD417/mMzUt8dPK1WcIEvFlZ6EAfo/SjBNIlmHsl6z7AhN5dicbDl8Hq2VV
SHPXwyIHAtB598ReYwogKP629qYbm2dqA9qTQJaEgCJfghpHPB8UgIzH19vAFiQnAjdqd9qGHhsH
FvZm9FI7BPc1Dsg/Vpsn5glbszYivgzuRvSbJ9HINtJvkBig1JLSErHPyGTD3n5w9rEY3nFpJD21
ukpYwwExRVW0BmJ0ha1hwaN6raY1dXWrxRm5MC07Rqb/PnKG/p6j0jtNgiucxs8rYVoDS9ZxywSU
c4RLVNtHYrplWC9nG1jczNhYYt/ETOqVJJV69SQoQXLxOEob3P4JyK0kGToQJffwvNJIuR20JrDP
TWPei3MQdIVoz5oOLf7MgLNO1Tsd8CLiqWCnlGK6cOLm8Ie1SIr102q7tNiAVJmJ/NSR8z4Ei2A5
QWxWwt3mpe0qXMiAeabN1dRasuIiWZIsuL6p545vCXlM/zrIIz4gDp2atgfcD39hUg1cWRAkGFZK
k8Ax+lAfxheNQSf4kHVCRfmV2ZNWcBa7m3wCHN0KgiWsWgDKsmBRkPW94p65eMEvBCBhicKfROdI
7j8i2c1Eybu5wik75mIX2iUKNONtQdvYmEM8Rov0C+17mGmy4YaxnSpIgxMokqFpxyWQlMv1mhGh
sj7USO1YGDKDGYU9jWLiPRroGu8wWzmU95GspX5cruvJ5uaakfMNrBL2A6hhRxItxgEo/Pqmiv/b
50RGhMChzmWINTW5MwLQgtHFjmARWU8p0rms3QwKsKLTxGW+KmH2EfM8CC9UMffweQp4O5qO1bhg
WkyB9ExfQBXxf/OZpJQqEV0TfCuPNDqHX5qdgm/h+g0XkIdl3k/HXAqZp2DCksXDjSkRWhnNilZY
QG77M8jVTaLTiAiNVHR8o83wtyk3rbMOSGa+XdUfHqwh40vr+E0o2KuNWlMYYKW+ehXKMUyqjvi6
wV6ERlIRDToY1oDAMqI6y7mqyijr3pAFFuD6zxYBXD0BCoeaPIgyAKxbLlEfwBoluYBL06CbRoC/
sDgxwgPzmOrzwUOEiiiULoQiPSQahNm1J3kFEui21qAsevo29qrt1b/BUt6AUTe7FuSVO3JkCaQH
AQ5AUSH5yXtRzGQJyEUkEwtGX1CVntF/cpfW9EKPZlawUrcCUfSO1hZA5T6pdH7UaJ62NEo3B9ES
1HFUSmboj5pVBgWVHmY+dPDJswF3MRlYEyBjw+FF2fWjEwj3BA26w5y12lVNrXkPAXwW6+Zf/UPJ
CI6z/gimx6xlAhBZkbBgoq5/gEGfEeDrJ9zsrzq0v0L2tf4bJzChLC0ZsZXeb+zgNHOilavrgL/A
SX9iL9SIPI7Z5YHGdN94sriLGopV4cSyFkOra/cvKOFfhAS6O53s+sQyA2B3SQtvpTy/zYZDKSgv
88qDVKURUj2uvBLaN1ZW+6H2plMRbPXJZovOehBD98akjAwKwfU8uSQrGQ3b0AHsapDKzzgmW9/W
inixD8XFlpXm1ZhCrUaXIu/X8dhBYWdGexJdNn/dV4Vb1gEnJMFm8v/uwvP23C1sQeSKmiYbsPkf
Z32MT5MPmkKJBSk0eDtW52BASbw2t/3Xq7qcno+5lJRqbIGoBgrowTpo8WmVF+ById15H/qzPN16
kw/1LbD+lCSbjWvqmYVSmDk7jyWGgGlYVoXFWLjAsjP/yrQ6hbECt7mu3HtucvjGdaXhsy7v6ea/
6qTiP8ms4RpjqEtmpXO2BPy0Pb4d18goFYIAqvc6Fzho+V8a6zQr62Hv4WFQbM66nHwdSn6Xxelv
x26HYkMSZb2UQyCwgyLPtZWD85DXv4/SljFRV5KEtRw3Xz728L/YYyneTURIIeY9PWOetJjySxux
hYht4NPQ4Jb46xXkdIcxWZB74XRLJy9jaylvlhioV3Le9Y4if/kKMy7l2Bl8/MFMWs83+RrV/soF
SZHCcywnr9noKbJyonHg0CjHd0PPqoOAmU4+jRTnVnt9K2DMt9EwJbghmpB4dEjyCN0Z4T+F2/gc
OE+SD0ftr84n0nNcf1d7sj7MaJhwTe15ZFc3B82NAX0BB/qxrwMWcAVQUw5f532v6ALUHzr1Cm2y
IzdlcEPePoy8H22JnAY8lNh4c4fporRJhQLPs5JeNRvg2JA0joSY4kAKVF8SeEs6OU3zUmgMDD46
AWHRqfXZSxaTwpBHY7HHOVvui0jNjbB7JXEp9uKDwBxO6Q38jBd2vlZXK92hOw5Yv4yljWZGTje6
s/syUouEwRc2zPkvM7xFY/vLUANezddQTvHeUuVcMiej5qr2Mwkd3e1/uzJzs+/2GoKRdCUPyVMB
v9ckXV436lPJZScY2Cw+dgwiVoqbSXwbmBFXLip5TWwKUBTPKlvUxRua93tR+umqgtOpc3paSV+Q
0RymTYGsRyf/sbqaTcWGh+F7vRPo8ZfEzA330+P2FXwpJ3eA4yv8moSQBcVXu+Wf9EfUd0mFGuFO
5BqM5EdqcW6NMalC9OvVeLhNwRBGhMYXKFZ2nMw6TlouJn2pSCcGK6Rb0lvImfNT6VO07BTMqvH5
dp1mBOcXiMB2kmKuPTTWeOnjVRwrlQOB7VTxyUl7UV59YvtROfuqULwKB4Exiw4daUYRjq3C3c34
i8uYwZvlHETLwuNIJ8G9pmO8qHNMoeYXR7aOu/an+jSLxJR9gSbGNlAwUYs+6gqukXQNxoGxtf22
k5upBRx7quh5olx6e4WFEAz6uhNi50cqEU/DYxU9YDi+twxA6lDP7opz9os2ya/Q3bR8irmjdxCc
ho74YDwxZO1ATqeDa6GPLTBwcevWhppwVP2m9N0XD1muhPaE0iXa6gD6nAhurKzhbR9wrJzSD2ux
1f7DLjd0IBPzifw1BchT7kpgTGSGzVZQuo+SfBiv1R+eCTqN14vcUOeQdI+oguMHJMaJpjbmtRE1
+zDxAPwIJZBXohSk/bfZIks8ADqGJdH1TWx08sV8SrF2fxSrQNDTQDmKKlXbSYnVlrqZyd8/CK7G
LIQRii4XBajfwQnBOGEZTEv5+f3xZYEmzo2jVrj9kB2VUw+AYQ3OQNLtjYS+Vb4yG9lNWF951SKY
bg2EG5in4DwxcpfmbgiLhBkQ7++h2NLCSaqd8pJ45TB8MpZdDHIvCGzVb0Ey35LuKayRftpe0i8a
wd1pyeg3Aw7O+2wlaGrSFZlOngiPdb7GMZkE/B92gsJBV9VYlzs5Sp9bEUVbn4NqJKKEhAXbh1zZ
zqfXjvNBGluT89avwAMZDRf+fyXyTgOAj87gJQh4GBwDHx17/r3CFctFDLsiSn42GbQDr/iQgKTL
6YMeRd+klzIOMHd2OYCP9aGfGJZnSbi/BHAobHNFlY2WqQoHevRe2vQ+SJNotc3f4i+BcuEpCmam
I1n/CJkINA/YTP4Z8dmSGVb1DhbRMQ0HOC3fFoZRemcmqNTd83AgxlsKytI9W6DrKbwIClBwJrPH
8j1yNdh9YkqjLLbns+IwFzPLvGIXQhRfq79f9e5UE6T3X3sAiaUDVb5xamw0hTiHj7WPcKxHFXsa
E5DzIOWM1nPlHwYn+Y+V3urVmPnoprxdaOBElOXdFjhdu3qPE18+rG1Hkhj94QpYRsLDxXmrpNBe
2zFTu8o1kRIG9tr8+63INhid+6tOUUYWWAa8K2MXdkjKRszM/H8Z63BUOer4UHdIn0vJclkLZqIa
xjwNvLaJhUX2Wl4Qs3WpUqOmGjX70ublFx5a8g3WtsP5hc+JbnR9UXCUXMwq8toCFrGLDFRtQcV6
9X91sMXaMQ2pY6bXtZKGTzTlYWS/sNvrMgbLJdlo9EYgDXmEbTLbS0BShA12yyb0fjo7IuAJgSOI
Osg0G8hUY9XKqo7BkHJJ9w3RENZv5B+dmxt2Y7bRDjaNxKB33feaTXRh7HGIDGRhJxbZqIbcosMR
YWu/HMfTPUk/5TSc7d2qwHKubGKAVT6LpjnflUA6Tsawyow6UIJ9i3hL/Kdtd65KqNr9j6M5CJjI
YABVLpTw+gCjdCPsAD59SE+Q4BM8ST7c5LS2nyJxoRc8+b7tJiHwQ3fpkPzXJbVK/yk7PZKs+XH4
zSREy6wAdsqgxrgNgMzdMGlOOWYjgKC7LJSASsKYBl9FF36oLdKcccBKQUxtQLZVhBdwsFs09UfH
FJiAtvPsg5Mtx1kvaqGNC20Y0/Ndld52EMhT5/LJ29g/ODxXDHBrx6pj1X3surH4GEXNI+v5OGMu
YcR3qIFhT5DrEI2SGQmtDUxOYMfE93/yNoGZRTQYhPWcF2/w+f/EBYCRIhzRctcpincn+xkfNigJ
ufM37mbkeu5BUfFguQfu7sf1wmxsu4Nqej/s63BwTJDEK6ncXXN5yUuNeEmpUd26WDg7dfwqLqeN
2gBy95Ne2VmL0/zdLO/GKvOoQn+iyqo8mWcABKBazIWRxfgoiklER7LgSi7GQsIzTy5AT6Ze9Opw
EQyNTIfdcza8w9k3kJRQTZCieQ69gTYG1Agj6cRRkIePuMSB1CmE7QK1N4LlTMBZVSog4yokDpMH
Sd0gKghSGOtY/lXAbcqY32RDEPX+sW9rqAJjJp7oAc/fSqp/hEt2I8wJbaJAE+S4Z5jS5zGeUruy
P5Behm92koRsU12usMiA7O8gbRhRqfjM517ikOeK5WKLsSd8q40fye5ivfku8g3YhPgja+TYcsHk
fMz31I203SAKiO7AfcTVSZiP3FluDQP717XDGEOM/KV5I/DElnZ8kfvylRbEyxCogif6GLpEI8+e
iZntuSGIrHJnF6eFcS/TzRNOSqAqWRnVD3dJjHvibxCxRiTUjvEU1hxeYwGeqhr+ofZVKVHbTK3X
qKKgC1NDEEKNXbLDEspcvIVZVUJP11JFceVSX86paGXPZXpuJiRzMFg2mtsX6Ai3Co0pY9IRT3Fx
FvUr13rWSy6NOgAcxYkOmhu89K+Qv2kg89OMrQlWAi6Xtnl/fkG1kN4gWW+gKUjtizGu22HQS5g+
eJ0V+vGuqbjn9ReOLwAGq3BdB1Lt0C8Zdeiki8iyLmQzRTjuUOPeRY8jAWQz5JnyOUfIASntgFI7
fkVaEsVNGzPHO0IWiWNK3opWP9OTyxwSYL1zDSehW2mYZkjhnmSyARJh1fDLTX6unT/GXbkLK0jm
GnQZz4Tg9U9en2c6SYC5HO65nZx58ZdgncHsmcCKpE31um9mVpM4D2EJlX16tFs6e4XpCq79y99R
eo0KaD6A35vepz67swX3+hm6PcQzdRC4O3JytINhYq1dX4X4o+WHGGF6VG/q3J1OuNnzwWAmGGSl
PJtto8CqB5nPNbNQbIPkFIRVDXbNevmWnozJW8IU4CcJS4++9f8w94iJibl2UrrQMgjWzQOpn0H3
jXBov6gZJTSBCD8uDGH0MmgrJiw6uU/DoeDWyddf11ygGzWzx9f+pKBT7Cc2wHhY5rwWXsKiS951
Hc1i+sbIA8WtWBLd8UmWFj9FTp0FvSp8rgUI9K/eCVwSNi7UQz4DAOkK/pq3w69qlWxEx00nmwsh
xnHhdrF2VT0hv2yYJ8YGHh/zFQWBqy+5RMmMuh80KgmfVSX0iMHgEkfYnybRaXsRoUbA0WyHUziH
pYk2jMmVIGpNLtXA8Y6YAw38wy3wJ9IbOobLhu5MdYmbq7IV5MW/EAnK7iaMVcCsJ6J/m3Swikby
EmOOOkRJf0bFx8SFAuTp0QNv+839ZHVXrrs1pYS73/7HNcuvpRM5tWFVufQyWTHFDPjH68/wCmMi
TkLhSH+QHEjCBf10h86ExDHWRd+pbaYp8Ja3Tu2OB6TkVVQaDGTKRmJaqh5OTsbq//UI1BW+nneV
UYzQZQeDQgEzr6fYAumEvo/CN5A30fGcvy09L9i1gUOnTzkRTpTufVNRy8Gax7/iWmsAEtTT/WZS
c1OZiDdAuvrLhbmcaVDdMIJ8/MpnYXd+OwngOySVwpkl/QsJSXTMpazpEIzcR1WVwFS6Jj/V1Evv
SzUywF14WwYTUhxFDIZTi3Cy9mNjO0/auTF/kTw71hIRpRVzFrxL6r1fDwCQBmf7U1cSD2TibnUg
sAa6T3UsDDAT7o7qXhnhIbHRCGh2VeUhhmSQzFHoYHwaHTSpLlntMw6akDpeMW721MRbBeCoGlnu
mk3i1CywSe+nScLT3J/av0K0j5ZIbEAvtBts+GCudSd1S3u1pYUbX2M1kDVQ87k0zlMwteiykwjQ
9iKJLmCt08CvRtS4Jx7KLt1aSVy9ztZpUp1xNPJyrL973mwzHArQU4/KNWs95FMEkkHsX/Z1Umug
P0lD6Lb3ZMlWFibuT8ZtTY71cCkU5wxpqEtpiZSfio7RvVYFkR6H1sxNtcA3b1mWuk6FizMiK4r6
H+MovOtCg/fC5ZJvH9NaFr6z/vM56uavk12hD4XkRVhOIegOiM7avuSi0CBiTmwZQ+EA4efhtWIG
IQXVbspF9OjoRKLehsCVfRj7qMrsmOTIhTt4VJfeaacmXJ4MQubfb4lSZ1G0z8JndIBT+5mnm+eO
sWrZI1U9Ei/cYdCz95TWKhsovmqeUmxsjGS2f1aSBBv+TMeA36ZcCBVBjKe+JeeuqB30ExBAf1gk
bcC3reiWAVoxa7U2GM2NbQcKJx034B6q5xEEYIiBuAgZN4SWTrPre4sRgxokORE3BMFsYsOwnsxd
oAnS7AIi4f2UCgpDO6bHPaqEZX2tX+msOC4+TroEP92IVWNiZkNnsYrkstzL94FUHbovfWlSyDKy
0ovgpswXkkU4JxwBwYqzxftkS32ApkWXstsvzs5mL1UGbUnKXgnw3TahuvUPIaYvL7Oi9YBgqvNR
n2GLXGT7MNF1wvOIZ0tgt4bisq+u7q+wyEQbzx105Nw7eDnUiPrdBzCoVLveED8fWAZkKEvjZem0
sB+Qqyi91GX3LPLYq6+mdiJSzAM/jwGuHths7jkTbOI8OAUdbArSWnK4ercDC03Wee7mkvTCIdRZ
uuPpQsh3rTxQpn2N3+XIOP7dpfd1R39Oo8fqLxqxi263DFaWxjUKbCdv/orsBSIbDObnK7V15pgt
ZY/xo0iQfbKLlF8fAS+r3AwpI1IlPI3n3hGM6yrCRSjm7lR1OBoDYiToG2AIMkdFAYLRKo8vc8eo
FtwVeGd4RiU9qt49lvjVb/hV3/3JSLSDGTun+ogn/lXEdckWiEAT57S7OQR1rlUPo7rZT7Z0rFPb
N780TrCr24pf5scFQmOxhZ+DS8cEbrX9VKVpP6xOSOn6C9/O4Jl5myI8xB+lgqlRlBKWcvcZGZtG
kJ7gZG/CSIw7BM6lOEol+hXrUNgImAHbx69Bw+az1RbekBZdImOe0IA3Ha2vLZm0PsfOG+tw1RYz
hXLFDUO3ZIv22Ai9psu3nrIuXgi8WqBHXagudd+8QE5H6WSp+0VnBSJMd+udJuU2l8ufC+fP5Kzu
+JMwfSPE0ShLaMJRkY9xCvSY9THwwbcOYUi2m4B3FoRoPskNa01aI4KODyNmLUoeqSAjbdxiZ1LL
LNQC2QQBX6GGlmpNLxJUsnFhfKiW8CcmpXb0I21QbzvHB+KIIwT5rm3CXsk/4/h4rVZWyOv2MXbm
g8TRcLXZ7o41deVpC/2AQ/Dkr6vc0IPnA8/By0+MihKOhn3ldp96VpOfl++pk7TQpbgl7beVvNeR
bFzZg/6rwP8O0WwNsMvhV4DN/UdDhmtG97GJMBfto4b1sohzuBcLDpGNHu8ABCMi3HuEBNAEwAI4
q9Jy4wq8YmLE9AvdpL8YurAW4yd2OoT+etitVs6fyNXtSWZ4lpfeMEBSPG3pvWpyCwoz3xT+6zJO
u3aUr4szhV3ibJJ4DXHIHa119sA+uypBX79IluZUmCbjYQPAIeI2Lgj5ptJcfTX3Xn6S6jLuHzdF
AFggDRgm6WmptWmXI1jjbG03waA7SberKyy8o9uZZro3nLOXvETDwSpfXDEHlzUPpNm+Rdajeyb5
rKGUDBIk/yLdijoPiT63meLyLOS0XsOB52jxTlTcKDSdfR5wC4bZyDXz6HpVG7hcE2qGkUtQLRuV
WDtcCrw/ahMkV6lY9freRTUNSGIH9Y+5zvPQYIGul5hLctHx/+ggaFp7XnhM7IuClG8p4Py0pNiI
8aCAEKCFxcK594VnDZDP4NPl+kUrRij39ukSyyoCAHnYaM5B5NdRGoKcaQrKd0zk1CqJ0JDgWsUK
nsFWQXFK3fdswooa+koV6QPr9szMJFDk3ru8vkJSpaju3C8SZcLTxhGQtp2+hokdchkgqd4apFVT
5USxbSPVl1VZ7HmA722kC/J7WgsjezS4wokCNZZ/6UFCnpJX+Bal580BlXoDs0m2l8sqbvam8ZRa
z6CqUiiUSAWS7ak9VGO0GXl26N2UIi5quAhPu/LWeYlNv9yCuUTnSwmdR2HGYG0B4ZKAL0jVKjkp
HlW7SRMjGQyYoCZt/lZMoz2cWmB7ohlNRijGoPAgyE75qBC2LG1kkKLGPenNKpxHScgr2w6tMeEx
cJBzbx/W1HKoLhA2DsEsF/enpau9VRFmGojGCbjFSkBtK14HMPkYkH6zulsVHfc7o0tTJ6SGCiHw
iIl5kN7jzPhY74kHHw2pfYAdCgJtGn151wlSxeYe3t3U3liNH6kjgSHN0HqX7TvzbtnO/McZfuL1
tCg8DQ9jsXTld6/Lzwenni0MOR7PCFJ6znSCfJWtamuwtvfO0tUekA9rq5LmH93LnUAsAHKJpUCv
SAuaKAlL5g7INXz2miQGaE8RGU7z0bkNOvUyghLyXieCE3T3+M8Ea8wsTFMkl+irqnblgnm3X4Rj
3Cb+s9QiPj3v+foJ5T6ja37SwL701LmO0iqtKMq93XF+mtp4xDfWFTNnllQ0erzYpYGQR/3ZQD6B
yN4KGJnFBaI/qgK7eJVZ+MQ7N/lyBxpMqGX/fweBI6WAwOdsI3EFEzYmKJkyV5JSVMPtSz7TkNab
a7Dfg6lkubTEpfwnA4mizHaxfBh25HdXWcMtWmRK/Hzw2YwQUJuS+CgXItbmU++6ubkUaBYboVr3
H0ZeVrTV7cJap08ogWJFV/LMuVhYQdXz+Kuo2efR9Z+gShPRIgMYfe5xI54C8QU7+KlV3byplBZj
jSUckfqEV35csapHLkfs1rT+fqsEgq0BhPN00WtAy6OO2Q2P9WXeauVJPD7w1U8nPrtzlwM7KrzP
G1Jvxlhuc1PaeUnnRcNRzy4D5lPiJ4N/+5EsLG+MzbQuept1dpqL4RcfwoIToYqX3DnYCGJJT8IX
B6EkidIPhlTU0JgLDoacgyjTVe2Be4ircwP0NZmebWPwjctBCkUFqTzE8s9mVl1C2LUEdthOzXoy
TZHRzuttVdOmtPSVar4ODQijewO54x6Ic8i6aO2jg3AA0LVDLCiAb0hRWGIFsJi5H8NA1uhWQ30q
quvyP7YdDb7FDwHbvV8ZXpWuoZpFf93JRj7Usz9NBXR4E1g54u1XarIxwG24NHSZuOAiAShyIGNs
1T/3H22M8r+wq2dNylSYIVSYqFV9M/lJIWmmVydf7FQlnp3TAYvXiubaOfiHdC48bhQERUoNngZs
QiMinQfw1PH48yTffEL+f/JdQeZmdQdco4fLtr8mjhYMwPbZ00diRAEUjBtLkfThxhTeYXXPHPdJ
SCgMfSQZf1l2VfTSyaL4xfdlIa++5bT0IUCaYjXXo4Mbn8nZ/4IluX4BLDzXzFHqleyHuWJS4NPr
bWOrj+0IneKObwAcAHDApWZJ3bS+Rg32fWiI1d0zg4N06coDCjgPwc/XDYOvBuOltt/eM7sI5sjG
wbWyLYbt5e3FwFEXfvXbP3KgMBpPkvC4Nuu1vEHl1cOo9WSRJ07zn/0sStcNrBbjMvzTpIGuWm9F
4N3+KTU3aO4l3XcRDFOe7G0KuAEOmiAhoZ+4NKPWtNpRZF5GrVtPJJpsWqd/dbKsrSuGyAgCGp7x
ysCNMMq8BbzRN3Qy7QOHk2YhFEvwq30ewj+CJraYs+ir0rKr6ODe9mzFGxNrpCcwXZTdYvBd4dCG
rFlNe4rREIPa23uHs7HZPDrzY36DTyvXLK7LbBhZQZKLxUv+fZ5X/iRrIsrC2O+K54bnpMY1qyVy
p27RJyrYoH24d02lhGeleSP7EueF/+OIHeP1aiLdt91uUEFjlaaYD1X585O0QtxX5Z0hFXmqRA8/
hFiHi65X8vKOe2rw6oT5WF4LV4hZXJdIegbSfQ52BHU8zatAEcMf6LIaiwfeW9FQBHwmjNL0BBEs
l50TF2OeHcrDoXedarkyBXnp76HfUFbM2sg3/XfEUtZyUy5UUMp3crzXSLQ+ecJ3o6LImPg3lprP
0xyXcD+GRBBmV5FqUz8L1yBHL6xJMMJ/IFvEx67cwkh/bVme0se4boI0/+d91kplJObmMmIOVF/6
y6hu3+acXiuRb80zD4G3Cj16LXYDw4fvb4De5a4d3rDESrh7uTGgPUBiY173vShzfJa0Tu3MVhDG
emlcxhgArqkZ2nonw/8Czhqo3OnQYah5et5G729ztVzej4hppTKQ0vGbkJU4wwqCM/SQacO5RkWl
sFL7o+10UgfWoPCH/wrCIo50aPCEDssaI9Jj2fs/Jm8U23EfIMCduN4TzquU9qMdnFpJVIYPnsxX
naMo9ALFhDA1ASdLcGYv4aZZSTipNAWCD1NhoDDXNXlSIh9mJr7wRBpAI6icIf26jRJDwfevUT/r
hAN5fVWYZGLntR3gQLCUivUo+8YIMdz/nifZrlg7sOEKVTRHMcArclBDthPEQyDL3xG1iBSRFUXY
jTtoRI6jv9Xhmz4teIRESzw2S1VnY1CxpYxCj8hELCeFM1ty1TYulAO5oiSvV1LJo7B0zn8vfIl7
XpLB9fZl7eUBlUd09KIb1n6jUxC9W0ldIGJVQRxcmARkZfefPUjGWMCXTjyXCwvSNnFfxL0fo7Ql
Z4cI3mrYpyDjP2UQk7FAH6QHQ9p1BMFCbt0GN8aeO1mvUH2EqhWUpniJJ591z7UxoHeBGW/229LJ
37qtGmnsiSNVex3hb1Wysny2yN79Wea8wvfnwMvfGncFrK+0PkOMl9AJ+VWFlkIxH+VGpDJRzWxr
e/z3k6cE1+HE3GiLGQZKY8gCUw0LFmHy2abVEx4o9I1c3fnuqNVNPswuaswSmM2GFYQU+KAXuBRv
J0uPv8Kue7xh/YGgzp9y1hg0SvCfteA33e9a5LbH7R7mIt3mcd3HKI1/UdEXk/q1WPgYL77GjaMl
tmASXAmRtuRk297CTdUsfAdQcplv4F1JcVCl0qwPHrened+3xZLQXrbEa6je3/JVFMNPBqmzeyFw
jHJ9xnYw4T4qwFf9uedx/6KSoIc4HDKcnzroEnAalNFlUJZt0zrfzrvdhkHiT2AuZAHpNI+fZnne
VEEXg6cJPRsVQyG4nCzw2sDjivUX1TkYXXYSSg2+G/xskZafVdFGqJEBd60Jzkcnly3SYzlWb+Gu
rsYzebedIzMxJBXMICO9IvdrYbum1u6tXHweL4/hxT8nVv+2ZeWKCP0pHD64UvjxoGv6k7N0oaZJ
LduyBlEDJnrlFZ6fUW4ZQwJihRTzKG55gkr256VY1VIZrLuo8aSARCXmt+Jc8Y7scvc8TgOaAuXC
r1BLUKKwIy18ry1CzzKjJTQ74ChGSu3UXJukGEkcn5UxYTv9hrYHOQgIwcs1e0cJg5A3s3kVjrjN
PeXKy66DTDwu9TRqahrY0evUTLQknPFANnBRLiDUtDkFZVaLTBLlJlBX22YrWk2/uVvdhxNQtmWf
5vI/8CT8TNYCmjWuyRu+zoSFVGXi07JrG1wZ4guojb3vAFf18F2TuiKP9ppnedB+0vNRpbqbVFpm
ichGVMUpivye5Kpb2v16f2BxHal/8H9XXDvFjZazBbs9/evvxaruKjzCt05lZ6Dt6NKqoLosHPmK
mMtPq4UfqLy4Ve7O3aEGpom+O6H7fmxYQNPwdzQBlyzYrVDmqF5ez8qw1F9Y2pWcZBrUh2xqab3p
nzIfMkTjhDDGTLfhp/Nz8SoKItQh9MmwEBxupPrpJmgsuvObNiCi4vQjtp+CQexKCMb2JuLugill
EjNe47FX5XpnxLbOOZ8wW9AVcgi1cILyO5ChUFqibvIDj8eF1vFQ8hjrc56iP6GHXfW1/aQDH10s
8/Bzdqborf0481jo3qrSPp6GtSTaSmDhzNfT/GCIiZWHok4xVLpc4Rl5OcCqeKYvTJbzjHgoy+Xw
duhB0prj9acoc0fMpfLWfKqfED2uV/AlcAPXyezLlrDbO5GlPuK7dw4gYhnVnIdLuuykzitpmdfd
nDjQ3bn3Xd0jm+os1Us8pTya+4ewADYUdjMuoDjlTpvtVpMCLixuji7dIOnCy/qCLXCNqbghWlVt
7qpA/AsLNrXSnORM9fhQgTtP4l/oVeUL/1WKCj6JeSzgK9MJE4U+NdO0sh9ajJ9py5yjRpDmeEg4
zw/8T30Pii8FbIX/RMGUYaH+585KoPF+jSok2xX8V+wQ6c5XtYHLID6Jw9GqhhV5bs3QK/jng5kr
JogwYsztwbyl/VQFuOkYplsTvBR7euM3oRYBA7Y0ifiFs29JCuamuVy/WIEgvrxAA0VCKxvmU88n
MOS1Bx3kXzVbTTFiomk4fxx8Zho9jGX66oF5qZ1O0WszwOJnDLg2RqSqWYgkDAVJ2/Oa6+XG8tzF
y5e507y8cb+WBldIUXhe+6fuws+igVJyT/c9JKwqBeyeULM1cR6NpShA5TTvA9JwmBYscLegl7nU
CYEOjHv3kVBUTOLKfH7CxOjhYn9vgYhUnjajqNoUwfhq9+NsPzOz3QFUazurCw3V/jQXaTqRtXIm
LL7Ia//mGUBerBfDZoLfdEIQoo1MCvx+bD6ZJz3O6P3lgE1U+AxnBSsPMKFJPqd/V11zUbK5Xnxl
4U9d4uW+/3GslYhPcs7dvkj9CWc3j/0Q/wbS5yv5c6XeMIqFbyuaPSRUoquJWe3szkQNAaDZZv5I
RWintmO+TObhNsqIxKu7YhkfvPCSfbH5LvXxDXotSL7DRkupDdhto8kR9QtFBC5Gnw1he6bbMXcS
JrYhpQAatRLF9y+jsWxLlfShmZ9Z2vuAgAftItSQaQtBAfPUqLxPn3E17n3mp3lBb4464V6g8OC6
/GiHoVvPFGfRBk3/hFsLAWOxbPrKCxhVVhI7gLuPZy9Ll8/KWE+awRSz341ZgmCLGjE+TLuAH4S1
pitz+92n50y72C/aILwIii7WNNsU8zdC31Yfaly3aSPzE9jqcwMwKyXg0ls8zBlvH9KV0DHDyXbS
nPRDvLlFtZZ79I95cPAvk9w0iUj7gXGrbdIsI2/5RnEB9XOqqv6+KyoVKTH9y9va3RbLJW/00na6
ec43MlYpEsT65aWeAT9pFOHkqRSBNve1M3ajea0a2eKITe4kJ/cfB7LjeJvhJrtuXiKhgFcIvJmX
ZObYT+xloMj7THp0fpXR7E3H65bevB5V0c8Oa/A3lk/rXQZBaeZKNvmlXIpw+AP6A6GOFEpojuhj
X+LIK11KozZZMU0YJKWG+Tdw/Pi2zeqxxHt4N5kZnGyMxYESz6DXchFWxXlDnl5RB6GZrk74vdNC
F/0RV5IHJi7ATwIjE3UUh6XXncXUUrQ8f8UCOgWq4c/jXiKiGN3thuV7ckhXpqxg37/5bkHTaiMM
si+3SRAqZaNONVnZuA6pOoIfYAXU010iaXAXfGttdNgrQqUXzyKp3fXHc5u2+Kf2DdVflAkDlt/d
fvDHu89Rwj8GAZjixmuV5GY/lBSaV9+h6BZz6JCnyQ3av/OxOYOYVP8bkyPvZ1uM9YwmGtDhX6Ta
/8lx5duFD4dRqVsSNlWZFthgm/ccMw6loHMa+Z0rjqIJh+tYByatqLR6HJqMAwQt1umiYhBtbzm6
RmuVw00yhg82FBF4ROxEqQG8KVNQPd/WpJnLHde5COKv3BsTjfgKrLT42wZLhi4bsqpu7oddPndr
eoVKPvC7e/ddpundCQZWfQXPmj40KHgTrNz0QCssbP7ToImqLE6j4QWFbJp9xiUFpk3jwVlF3E7q
5j814lzXaZqX1xFeHzuVP2UBFst/q8xl76vaQg6nMdP+WilItULesoc9368o/7JbQcyO7n5QOoah
JITNjb58oGHPCBo1zVnWfSLrm2ip24Jd/Byj911aiI3fIs40AkUl/7OEVzcestRW0Pkl9AZPQllm
gXbN7B/XE4FziJiTonO/5QkruYWQt/+YemRyKl5FrrPus3UN9yXct0Ft9KBdL8VHJ4uB+8HTng/v
kgNVH3PivVtJk4oev/rzZsEJeM+dikjGvk99/drQX6Nw4o+/XQ+uGariShw4rbP5Vkf2A07EmsD4
+rsYkIuZC1arJtSr+dZ6G/cUD2dA+dD9rLE/XklddEL9AP178OsXLQwbrWN06ZnoTj+3EuQz1haA
sWZ3/irnjdaob18gn3iPYMqHI028mbjwwqrdcJTw11iseCgEfzlniJT2W5SfCTvED9EFcvgpGkOx
LZ0zUOjOXqtWdHpwnVuB787dHAano3l3eEfYY9WqPIfPfyI3rd3hj5DXWszPq5Bx1GmSVPN5gT2w
HHsI/378axHPYQ7fnRz7Zc1En+bRWVtKk/0RW1B5x/mFu/SfID/KiTEor7TnUbmKUdpln3klNNZa
Sp96eXls0btK3RqiAMTGKeEbjRjPlKHlHYuQjthJ5AYlObrnqxHv+m3BpSBT1tQ6jote3K9dch6E
Hp6lbIqcOnY+dXfVwj87PRqB1kywKDm4+7j+g+qOv+YFZha7xzjkab47HRkRA0TiYrCKyb2/Hnfl
IzzOwaOIRM6DL1p1NEHNQ9J7kcb+DyMF7vOMp7r+INpF5sBKN/ayn3CQndW0lWP+cKH/3d7oR4uE
4a1VQHA1oT1yc8MN//QH2dThxxu4FziZPpSC2knu+jl8ldXEBrOtMfyXnVUUu4biYC9TaeViYSTN
QSgVHqvHL+Xlf0TC1aq6oQKOxgSQS/1dTvSZ5E8SVW2vzY8wJX+XyKvThQ/VG3JUEsi7iUbvWFuc
fk1XsZhuD2TGkDNGZw5DnI8A9iM299Akvg/z6HCa8LtpXjbX6KxDYTl2i22M1YUbab2TwMU3wrLv
7xCho4xKQogfd3B38EPoeFEd3z/5FV+66X9rzi7qxyPK5Vz0OKhcZj4NdbHL+dPFUMGY3PqodE8R
UmiKXoBSbI7JefFObVIMCQ0qn8d7nH521QgZJ/G1UQ/CDJV1wZRjsj4yARxuXd+taV5wjQhsdiui
GwtMAh+Rif4sMwlkmfAjrmqasXGXs8MBHyWz3NWYgeygdAawqxnoML1SXZh0i6yz3jmiqIKXQ1PI
J3dLYZbBcAgptq/BoVCLFJNP6y04VeGLkv/80OowsOFfyp9553w+9JMsRlLssSDAi+17zzU9ZetK
O7tAJuiVDq0rmfIJ91JVTwTfTQEpe6L5kjbk7isQaJ8SqgluAUGI44xgI1TbE1hSWonFxpa4Y2kr
M+M17Pvb/GzYqbluLcu1ERYz2AZO8Xddtc2+xGyvdO/sWmKQR/+a1bj9mar9cZ+kOiQ/q0TKNJPq
1UIverj5YzIoC+yGNiAX6Gal5ijGu14XWHWqNgjYhTWubeEFFwV9rphP1/9/qTmqWXBuXCzpuzcw
VKk3/f3EOIHjTOPauJfo4VcRApVVog/RepEmrdfYOjZX7RFlcN26Vk2FLogaoYCBISL4DWwBnbip
pWbw5CLv0IRNx42eHGXdK9WmJmK7OULMf6MK7axPRVj63n55/aj/XggX+38cPzq33it9I2PgcHnQ
e13yV4Nso9wjp0jmS2JxRfbtSVuI4okDF2WiQHlSi9ZVVfOl0qXe+UP4EVa6vjP875FbVTuTCQxz
AYKS7sDnzwSBfcGN/hJELZ+WKYkMkgdAvPSFwpj1zyTz47p1/UltLSKASz+ogC6tuX9aogAgMq/q
imVzXKZalGHmWJYsYDxvSzC/DjwNizsgGyDre6CYQgNjuEOhBzs9FAxHx9WAMZlXjiaYIzRDbQIT
szswGlNksLZt8/ilIYEZHdntBaMtsRmtQ0V0G9pSn4XxZY3GXNtuopgsP4fOY3zkQ/Sare1VNG1g
oV5D5MarcX4PL5H+Ohb9Yy3GHeX9KPT4WA38KF4avZ6iwdp5h8zK3zjZZXem4Ttw/CmWHSpYtFLt
bas1McKCiX0EXycxlC8+UXlKu/1rUVXtvzUEblCRR8nP3BU5X1ePNt439WkFhMMe9zPXfPguS57O
Bsnf+XPcq7qlBuZRbrF6ZCIkgQle4NUA+KxVYi8M1O51CMxOv/FgbK6g4wD79tpsBFugl4vKd4fy
IXuP66B5RYbdNIRetKC9/nfGKpq/K3zseQlLCwe4+vH3u45JQvrIH588giRozkEdEBOHJCsC7zQe
hi93o65ENTKuAUtwuc8ueXkgIm7wEFeIDAvBfNX1bhntW4fMV3eHTOaYvtlm1dGBm7ytvj9JNS9D
EbW+1Mu86+CNOHpvVRr+41TW2hOWxPs1hEeVuBGz4AtTVXlI4TOqHfCmxeGKkaDdAj5TlHGBMuQB
EFqg0jffudj0dRL+1FcTYhyc365/79niv9V+XVxeoPd8ASSgs4P7R0qQPoWBbD3/UQ1NdKBcgS/a
w2ZcHLNBAQMhHQ2oTIU4hAOTiFgN5NQCyHhTp1u2RQnhoZ7Fk8/i60LDsqBlsNKV8Vb/er3B6DSY
o9P52SWZaHUlqnMJuC8pT7c++vfeuuzkvhS++GxebT9E9Z9uVa2Y+HTuBgE9UQ4WVA/bzwVKVi4z
1GroHM249wHxWDKuanNokCumZ3FXYJED2r7+Nftg1e+Op5pZAd8459f2THUKoxXWrrfjnJvjZD1o
E86KHFWRzc4lNAFLSfKq5cbuDNpvJqZlrRzJV8zTUjH7aSxr7hxt2QCeVr2gxib1L0xUYUMvC2oX
Q3kxxXm7kwvLQ6VibUwaTndtL39ajqF2IT1BRJF0i+U9jL7I88jJsf9wxDr/QJ+eWs36JoGr8KHY
CtOkG/LEjpzAdSeOum54JGewgU10Q4lOlqPZZ6V39Z7EsMFI2fARAI3VHOBH6evENT1k4HZbVYKr
A67UBgBDFHDAxWpmfy2lKQnjPw7wARCENlmDex1bo+M0oZkauCFK8bNEZkRnsRvzpFGc1fODS3S+
yuekaMvWpBXIsOWTkAXWXWTjiqZRuWo2fctnvKQXfnSnWzaDjM7MHXD4kwYtiUCPqj94GhwlTY47
CuuOZaEgUvHS6LQWdZfjln4AVPAg4GFD1vtSgnSnCqTvvVJuHEMCSXZLPnvn3ok3ONcYx0VH/ikD
gXVDqJe9r6tv0GuQFMwb4wMcIfWkNtZOzov8FWHda8+CQp79vYrTXEdcwcvSWxb9uNYl7k2zyuvu
kw29B8cweXrWkPtDlz+Gb6hfSC+wQddKVJW+Ii73g3nxmJZVJYMwqxH5MBOA2XSpQI5oBGhsINxu
pTL7mQ0OYzSOSaSpbaGayRpCbnwlXR4XNoEIPiWeYPKUkWJFiWRQ9kivARXD2nyKCunOOY6rkQ7E
2435ozlRcPNfbICOpEaw6yxGfTFg4lzsB66sYmadvncDC0gX9FGf78G4NVUIlKGZCBZo+pCSfQpi
wyZR7YWDa7/0QsgVk2QbUQdFL5B7niOtwv0hRyB2uBogNPxZrk0Puxyn8CplGmrqavbKUf11w8rV
H/wou72CR7XU4HyPdewif6rISRLpXHHoAjJMrNNP2CxNYwJ384MV5ViRxzYtxcATpzn1hLnxwY/h
KdiOSMEi0H6PuqB8Xskr9JnKjK8o+54tM4Nz8jD/ZtLjJtHK7XIVK3F7col+Lz3XekkNJROgAu+n
SOBN5DelDpDo+TMcj/EFykym+RiNEoe4g91BiMkoPk/Ndq6SD3ruHPf4MyDp5uLg+R/+2y3ihdsI
5wtCETI/VKNhYaGQ1OCioCnT7RoUfxC8M+XLosvrnFofzU3alVqbA/cACBRqj3FZzdbjBeqx+IZX
PWbrBFqQRW6mLPBcFHgTUuXZCKQAApasbC6a3McFNmQUadc2OK4RRkHsJNHQfUtjH97WFCcf1W09
lJpfqJ7JjucYUKHHP9Lh3YX4ViVjlnZB7XcP3Z1u39Es5PVlJ9w47TPxNPkJDWn9dhIPAbjtfrep
H31MaW0pQK2FJAXo1IZn/cX4PSdAfPisI5y0cTSg1Z+M+cHc+yvRgqkUugN88sLugDIwUxAFR7C8
2u5YSXNYwtPuIHwIgzZTo4sBmAwcCOqxZo3AAebxclImi8sxYqW1WpJIEzIiddmQUAstkHcure7q
1RUIbXiDxd9aE0hqFQFP6oNcbnTJkuWkgJtodYoHFINWh9vsGOM89oU6mZtHv5L/yrR0ibC0bjIt
lkRAN/qXGuPpgqTG/xg5SF3ymkJc/l34RISXUJYYGZjkog38MBqe8hpxn/unm/AskZq8/q3OYUvG
Y6Ud31PkYhRQ45ilqgWZv910qLLmcsO0YGMFyPZAzgWlJykhVcfz6XImGtBTpZOXrO7DnNe3b1PA
h1QZrQUkSVFXyWEly2PZAZo2pV4jTw41o8AMbISq99k4qHLqXuLu8fzr676LpuKaO+mTqRPJCs6f
b2mIjn65y/ewKhczeGG23BRbwghzhFV0PQsevBW92w/33+niV1oHfmgh6+oIgX2TJN9v/BoIHJcO
Ap51fF3SgsePCXF1xwG7BXh37Eap3W1s8wADlsnVfkwep09uZp+xJ+LPqdRM/t5x4AesRnloIcFx
j9uOVPHfxHCz3hOGkCG/Ft+OqMFPJw5ssif4TfQ0U5nb8v0xKhExSlY7RyO5XkuZpdLSUV4wiMdK
2BCqblI+LPuX4dm2MnLdqeB59X0P2qRoFClD4D1deTQzDLfYXvwtDyeYJRi+Uk+19BpmDlDK99Ro
H4G0VGM2IENyqBlS3aOP5p9Ch7nfWvcKnLBA6okTsKWOJ0dIVfT8tDWejnRvfdZ3CHuA//Z72cNB
BQirgfq6c7pdGDi2p94z5lsbQDtQoRIsLDpyZdiB49h9yScgsjGoQb0cJd9/ulSMaN3EUYsKYHT6
L0OD3gjDH453oXyVKIgmm5tzt1ZckPZjwgI0tDoFU+BHVvrvAN1J3ru4DQl4DxNdH4jeulwyco7R
HD6Lp9sonzP2xXbvQJP8wPGVUBrcIfn72zlOcQJ1icUaa9GkLpOiGCrCr7SAvTwx/X0YLRJMTMs2
5Kz/O/m+yK/YTlthXtg+ii/5tLzGXpox8ItPifwrO2xehyQTOddYr2EJs0zjwcrFEpnQoCnkA98e
zm/ezmRVA0cdMMEdZ2R8r6VLrJj1CLDIVZ1KzgJ7QIhRN4SOHjt56lSHIuz5oHKnHxMCJhFh6xoo
vwEZPIjyq5S5xxJTjpSPWEtg+TJ4XqvsTaDzIHR3U9qJOvLTtTWGZVrg8SZVh5BJ5o3GsNrKHPZB
z+5CyD7jBsX5aKwjMkrFBkUR3vs8qQZv2zHOzbhvcyPxtIQObdfXdAvwc/9u44k++W3P98booOuK
1MXx50DSc/UVUgk5UwyAAvshm8e4EK69RqNloYl6CObfmx9hsV69Zi29Qtc6Pg7tjsScAae1yhCS
M3dtl3oL5J9eFh/utGgpr8yoSaPbt43QU5RMncp4rJHhMak/9fehwzhoxbk9FnBa5JG4Cg+ls5G7
AzeUzWM//wOHLz9ao/+ft7IU9+SRb+X/QyzxRRoqEXr0/D7txNL7MTQif8T0hafu78RVSN3Bf4X3
eUYzjCWhrzjNmLe+Zz+Eh3sFnxIjt/3v9EMAzrNwKlLAePEDXvWRg1BYlQbzuMcXutkVKH1xdsDY
CwGppBTD1B/UwzuLAG6XdgVTcRljeG/yD1JLJcOgdOrhQ+J2BhtEv/6Pht5FmZUavRN/eiqjPOTL
8JTkMthnglMgWhsmnMaaFssTlOBQtofkH9l1f/RoF6LT/SIUSE+1WfnBT8PJF/ULXso/73+ihywz
SAkmKFJVCCZeb5nFnNQT82dUOsMYtjndgquSRHS7oSShUR0V4lIjdYbnAm4oOCG0ErtbUqAIW+I8
qFg+mcKuGeNZKJoRRAnyVkvwkL33I8A1AEhQIBk/xc2HcatuE2X+WRHNZGhJTUASNZTc3r7bXZus
2sbM1L10e99Ihrtru4dXeKgqrV33jx4YicTff3Q7FYBRFc6rVpBDTLzOyCKYFLK+OR82jcftXCb+
H+y4Jwqo2glpu3vo+ogMRCt+q4VwESznWUm+YYfZSD7AncZSLXR+u2+VZf1F/w5PSoSkHlyDPD3i
zMzTozpuicygH5nZ16+MJY8ipzSGyC4lLCXPYnuGQNprjS2LkJzgt/5ymdvKRFPmQ/zFkodG0iBy
8GWERiaLwU4SwHXrIIAYAeQZpASRA7gQ613pnCeI28FPc0b1jOEA/yP3IBIB8N2Q8/Hb5lsUYF3L
ViSkgI7UWjQsBCD2zra6yIQoA4C4R47ebLKuwGLMmWoymffslt69SrGkIiOODbUrOw+m6ks7TMiM
GGa4Hll6QE3zpJ9slvt1HvZY0o3kdKgBSMzWZNn55C13M4JzNvJHaoTT55UX6oAF+oNQga0YcCFc
vLjT+x5g7kUroc5ZvZmHYIJfegOOkVuF3R73jseO1kuaVaXvzTQJj6rH7F6d14hD5sFIQdkEXs8K
rJhYabWoliBpuiXReha77EPc7eNQiv+bJvY31TWxTCtmpKHE9jTD7V5Rg+Y6I4SxpPiU/Z+xZAvg
eaCvdI0/qHhFanWoyrCToq2/Mdo+YTg+EZ36vbiezqPfP8uyMsMfYGEHN6/4dfzl/rvqYvu+rOgh
82HildB6lpNVw2E180M8meJyny4Kvhgd0zizPwwQfM16SadbHq/Be2VlmIjSsbNEwKoUsGSwTPl0
GYUdhMqTUS9iSrNhNK3TmRGaRQ3H9ph2V3EWt6to7zqLmxZf83Poc0cniN8BOPpycROZ3qga4Ya6
Qcwxu5RGUrbnCM4pMYmHjjvx7ropJjMLPo7mgtm6aHrTEVeOiPrPLJsKP1HxYv/fp72kxrdNuhKJ
2srt48rGo4r8IqrTYr+bAiVIsI5etqdfHaOoGS42zl+mvadpuLNNTEczl+0Vva2PRO1Y+OLND/pr
VCG2jwi+IUBIq7/ROgwRU1RC5YKjvxS525JM95RW/2OU5Jr4JUfakGlzPjpAZypm2J25bXe6XMhl
MqD4WGPB2EH5v2i/UKtM7FokettbbGaWyhGDIbVWy89NmvGybxMSRgpedfVW10HuIMF4Hnz/8hWY
Du+2RFkLbNabIqTCZIW4iqQbio8pstIwK27DBmkQBrU+1mZRKVEQ+m8VooVpwD4v4sB29iJfFv37
0hJgnXp4PXwkRjRJpNq65sAYzI/c4pgw8Vewaf+owjT4TuP1DmzqMttasAT0SqdlANajN/ld0JLM
pziv5TYHHvVs+dYkfMnE9TI1LL9bVrAhqUMJEZPnQafZueOSK4enV7jAdvlWYzsXhO7fbqLc82GN
EZHibxz5GBbW1RRNpaI7dmpjVFfLrt8MIW4YvBjj96E/aFVV8DOty0NmxqCU72M8JgClE5Z5r69x
S/s8rmCrB1PNmKopq/8q1Mc6Q/7fv65gSVg5BvkBOeUD39ZWZGYTfdC6hP65OrBfkEMGK1QHz3SE
2mreE9wVhALKNX5QbjIGqoPHQnAmqy9IP0sj4pGIkJRX+e3sUkcC/m9neYJz9HQYX86ksVL+TwtH
hx863KpbGxh0dhKZNQMWS3eyVLBwLhmQ15urP8PGVpLUYbqwx6nNhMg3IkIGxktWH5AfHDk00cwA
apLP1w9bkRcJ6E6vcMXgipogs4/d9kiagjWATYWtcrmh1Cu+Qj28MCQquQfsHumhlHTj+C0FKPt5
ZVHPEGKjYIm7tkFi7Pxkq6eLB+PV8kH8V9J1VqfpngipjApsBVM9V8Y1UHU2TdbVlVZwob1XfuKk
AKrsb2Ye+l1nbDL/rH0Q+Dkrelg6LTlD/A44hfEUg9aWMqWzPmdApzHDXV8yPxhTywnEB/qu1u+K
JTlQ6jNruvL5eIlGoCznoSs04apeMdG6DA7KQBdXdVG7ocQ1aAP90zRgLAQOD+tQ09uiJ2EmShBC
ePkEO9JBBS52iFTd3aIDaHbne2l7uZ+AW/KL4hmW10eKeOezTnocAlM0LrZJGNBDDC0J4yauuv4s
6vaQYicJ9qba1erQvSm+gBDNU3a17DA12LjhuArOsx/DXbCKWt6DgvgfM/CCqt3lyqWklR5tDXF7
hN3vQ1hxiCR4lmjjxv1mJcv+viWU02o5ZV9LqIM9gsHU4kiciRwuS7s/FYqxHXOlf3gcAWl65Ltm
nggOYfN48jXWmTIgF3pFV1ixmWKbNWPSG5UhYWq0Ce0po7Grzq0Z9LXEr+n6bwOISrG66LJNmkqu
qF03wjeonAXQOzv3Oc7XpDthAcK3JZ3sgRX8I+yhcFukC9o/K8GzSjZ/LhuufohGTe4ZBnwUgJrR
GbNgvA+iizj0JVrjvfks6MU5KMJ5rAjhiwja4Br07pdZOvTNoSF60n84p9uPTOtA1qQgOuN47nWU
43lyomA8NRjBLQ00j+ruMKrpHoN8Cet9pHdqsfe8EVEKxnoe7MVyIKyODa9iTGF5hYD3EnFDs7lO
N0GfPEgqiTqXwKvc1ntSmKskSetDvNOZRUMn5c7GbzCUM0RrVKUlVlKNExxYscPgIS54w3OrYpja
PXHoLkal89/RGIPep5vcsqqkzXj6nnBPIqUB0hxGgwR3kDanSNdAo4/duWVr9AmYsKr5NkLE2x7y
fXh7hfEQeMcGxzQov8R8O6AZBBLO2/xkL7wN6fG8kS3QJClFdUAAMBBx2YpBzQDEn/PHlwbanItj
FnclCZ8vsKgRJsgD/gzjd3nr15S4ugyGCIPuOorqXc0X1gY4xS4ZEgjPCdoOlZwateekCIaCCC71
x2+STiN4cQLJhYbdgwfRtuhGpkDbzK8RJH1DPihHOh/cIv6LzyH19rMQNpY85qnrW7lBu4OTTPHW
JWN/jOOPM9H4qXep6GLmHhSXYoYstQSml07I2rgnDt5z75pHsO97E/XYAbh4E24ZEde4xf4dOtm9
5+b0T+PIl/NUbXIz6zYimYGzl3D1Guo+p3qNV2shs5ReGT8OEdx+aL9hTlpazY5NO3OJXS5FJPJc
21ZuQTAtxVH0vtSrCudIqPgSP/1GTbRAANIrUkCykZ7sB+WJbMoyn2nLCadPHMgbOUnWhO61It/y
l1d5bRXaUN4AsAi5ToVRfA4eRGRbDw5/Kz5yIOS3vqx+J2npvYG6xcnZjU8mlwafU1PWjIqZ8LaQ
A6picd86YiZa5QTqRay5sWJMbaAlbejzy+AEsqM5HSMdL0Vjo13yKR7urJTX48kg1OiG4GbCaUJ4
7ysOnVGrjH0mOMQXRcIfts9mSgfK8G+zLf2zD0UcaDtPhaBoL1rzqy54hWLAMH4sYlMmgFWNIFS7
O+VHkM8e7n7IS5JvpniUhjgl7PTAMqGTYKTMqR93fpincLyVEoiRobdV80Y/HT7Zyc86KxYQVc3z
7lCesgd18he/AkIAQ1XTtWSa1g+Q4iXBy6eqREGpB1xcH3Nr2Pnd02ttIsz1JJ6woOwg9GIzvbr2
NPPfa2zB58TiWxJ21nh5Lcd2m2I/RZ0+HNZx14FUC4yrYA2ePNXk8guLji686063oMKo4D6fZ4RS
5cbLpO8AT69pOw4jm4POSlbtad/HDKh2Tg6VOu0ERalEyBUWXcZsoQrSmX9ujjuMhaFMkZ4kJ4e4
65a2mCOrHJhMqp1SW5HKN02Jv1g40vNBo3B9DDdDnzxYzXKlpXWZayrGPj6kTvkgeRzag40wMDSv
Edfee4cCUomS4xCt985tk19PMCVytTY/xm9oRl3ZR+1PyyGSTJzjaP+bnIbU+KPF15LTfIj7G6xx
mKNjjSeCe/0D1EiC8zwpUtRZmsFPAqIv5OMM6qmYkxjgifAEcKbvj0coWHOYVOrK35HNMYrWZ21k
4S9hMkv+e8GyG0hzVocMsEdmgW+ljJzHNjnGziegYGBG46BBi0Kj/sDTKYx5jH+sGv1VZksHYXtd
rvw1e8aaYZZRLIy54vBPgWG/bc6U+loIQxgwcWaQEt2Ktlkp03xoBOVqcVsx0g3uKny1z2M70TNF
ffjsAFseo2e5+6iQK0nQHWn14xO0Sj6GatNVV8YhBHC5Af4OWj55HXBIjYdifqt0gSIxgfJy0hft
71oz3n1fycPxb6rjirjDIab3V5vHFK6lpGbTgBNQJ8s7DtD3u+cbCgAjsXdtUbXx00BPf3tF5ju8
bEDZEuSE2ihpYEoUXFnGYPwmT4yHqrzWO4MOsRLSPkuWNolMQaZD0Q1vMSDfF+kF5y6Jq8QztCSV
seueVQYPvMJuCuiXtOHK2cSua68VneCK13Wuo4VFZ593+81Kv9SgJ8o/gPpSx7FL85s8BcY7LLN3
OlgPMNhrVf53fuBFRa+xObYi7QlhFbZiXKSN5iepLdWlyfNnuX0+QDQrn4ZLoTJhu9X6ZxwoJFBX
xWvkuR3OV8GZOSxlIfdNxQQDY1qKQGFf4epzbkWnlFsc3ohVb69vuMytrxQ7PLqolDifHDB9tnGo
6yFy/ExKpQM/dE0wOTUYm1z19G66fu6e4if+Kz37f+5Mfbotdo6CjEp8vtev044h881uXc4uxudx
LraNNJORos5GkAVIAblgJib1EpvL/WvTI83HsdcR7gTMtKRgp18luFd2A/PGzlZgCJ7RMxfE7LtW
hT1WUuMChqt8Yyf5jdRdZd0G79eBWTmDFaQJIoEVmz0t/ZPmbSZQEJy1sa2J5Ufe6FH77PFjZDCg
e4U12T1bX0h5HslXRf6AJsoMuwW9xOB/wZG8N3Db6FPotXV2DfzYXJgEgWcRR/+yp13U/aKvj3pL
Ei1iDo4IPcaN5klwlDIHvk+5JP265F4BqDaI9CdhEojbZeKMyaNyY1y67D+hfU23vc2OHfqXsqXy
DID+xRetZSFUmKx1K6YLmP0oPYIYLfRO3MAYGKL5hGPVQG4x4NUIikMfagznOYz3flU56+P+Zz93
00ejIxOv51ZunBdfwF//7X56F4XqvE5zz6VWjBK/IBZh3kTt77iL7HmCZSUsLmIyHuyZvTB7G1Rm
rMMzRYznW0TMBqlpWx86ZZiyILmuXoAwJqCQSiV9iPbEAmSB+A5TADbeBKQdEdwoM+pjymwVRxjb
KGZHzU/kkd90Fla/BzTAcuyWyasjGC+QVUwDGdV93czWnmYxR6osYoVrVI3pnhBF2uOOG0jsL3UI
dAB6z/WKLHGYxUQDalrQ3E9nuxI4EWDPA9b/JR5CwBwyAWjA/XRU+0m1jg2wG+FmG4NoB5lFRNX1
BDnlXlXt/e8lVLpUNRk/gnvnWKjMdF67d+BFoNs8KdglM3bAIRWimQCrXvhjTEvu8JqUMJ9aBnWr
6mDV2WjZzBx4D7id66vG+Xyltuou2W+mUWRxokaaTldyCr5yA6+uw07d0lP7DpXAaCzyCHIoluIj
LBLndtiGi0F7EkFORTWDjE6y2eROBszP2JTaIjqDPQB/y9Fv1aE0gArTsvJkxY3m64NH2z6XSz2c
GEvcRKRy6jElfuALclOR8WZmKH/ittGn9PDnwhJS0GbftZlyngVqt5uWwJ7bpxZ7CJvxuxhHl4XI
8bVcUUyd5BRxpAK3pzuFxdEKSXMIisMteeewkbWqRKG7hglN4hvl9iVeyV9ZKm/Zyf9v3gdud1Gy
biYtVQe5qKd4nfm1VWPK83GiJJonyyugkoHlTzOiLTuCr+Bg6jamISsQWZTx6HEGBrg/Rx0T8X9j
N8GKc6vPvyRP7YQXYWQCrNMkE1u9oJQQAoepf+h29fU7jc7v/oGQwUfmQPi1CXyxPq0hfMkuYlc8
rMadtR6hP6MYPWIevrw5xLhsqohu9uS+geDa44n4nWGW2vPWmNev8zl9gim0lup5wI68MN51+kaZ
8rOwmiW/DUegOb2mKamNPVMRAUORhh3JtOa47tIJImJNaILbffxPlf/5Soc4noVi9rBC5FB7I4ol
D2omc0QvzGhypvWzPox9XwxNMKl69xtmHjOQSN2jGvmTwH9cNog9us7fcOUQqq4IH3nF8KUUGQTK
+YKOIlhyDXYTg0p/pDBycdd01YbYP7ELaODAvUeUrKXdr7j/8ljZJN+0vdCMBzBsDQxDSKDu1oen
5+OFAvJr3zJK+L/bOXkDuH3gIRxt9hRiIctCq9Xs6LrpRNSnF+f9TwjkPVUzSdKHPsJybbNW4jdV
K3ViNsunOK6uhMFH2dNESppgM/s1cf+DhsqsiMNuRzpuaI+NRWR3l1+YsA8gRFewQNg7gwiGoZle
BgckPAE4jylj2m3wkV/FDXh5bO2NLC+AYSTdhCmnBbpyFMj9Aqw725p1mn6loCczY5//jrylcT9k
PGVCH8/qX8CytaKSVHQ+meyxZD9G7EF/ulQUk6rKXgra9cieIUQUwns59T6oMOmzGNOqCjGW4NPR
lrb37miTTycTuVE1hci8hH9PKw20tDWWaOCj0wlk+NqgtkjZwm4Nk8sRThAtDYHmkpDYTllE5sUe
sxTYH1FTIAp9jtS/jA6LDxB18IaHphiTH/EeAZsbXpGO1ACulan66HtEbgxhiDi3Cw82j9REvUYG
i8AFi26uPrxemlVMdePuU3XpTW6hBIK3nZZWZRI/eqeA+ZukMiVwuO7GPg3k+LTJj/WjqgipWGel
aCaMSuz5ueFyqJRj/Fo16ZXasPmgBxbiA8HMXIZUX/OfwMQ+xrPGgFRWyRfbBnmYrAFcWs0IxP2A
fHmAdxodOVFnD5e2F7bvflyVWTaDP8aFem8MXBitZVmXaPakCV0UZAKFfBy1XljjfTafoqNVJde6
rlatsYobk0hNpT02CfycAXNjAF52eKqrcAi8Sqk8zaJOO5zWTb6PSEdReEBtFPRC+TdYde8TqsgC
TGUvnrgetT/SH3tDp7v7aSXuRWPv6gaA7gCZLRaowwnL4muVCdlcnJ3I4yy8lRoenMhMxlJA/rKl
3/TPn+mxuFN/wh5E91ojXQja83AtlVkP+dXsBWUfH5jJoGm/zn1HcFTw2Mw51WWq8yIViIKIucdh
7+4/+q8mlpiNX6OFMp7YTZdG2GCW2Cx9+xsACuO7ZviqUixI+J/ChFdYBzkaRk3VvALkbz4M8184
FN0tPep56R+U39sZZLpg32kIjNvfLL6G8dBpN7FDI8BUm7HB2zw8KNU1xIGR4bcwcizbCFoOr6/w
LjIlJyHSVzCpVZLhIyrFW45iRPgWaYd+Xkx/JEhlXFzWgpwBIXZTaFHVxkCUdaEKBF9TZ8zcLr8t
7GbwwcV1YzaX6BTFnMmZBrP7OHOuHhlS5yu2C3nrMNtOi92yC3tI5DLRoVM7Jr8RmHbdgamEa9eB
UJWxrEYrvvLY+oQLrnCgaUSaxqrmidBJHxC9eA39EBBJM7okY1eI3RjtXfArzj0ryI5FrO5jfXni
/oTI2ThXgIgt5Lyb8jevcbjiYY1IFqEpnxET94qqOLJViueTITV0acxtpZkrUpCRRLNICbrA62rl
yU8l0oDT++GcCnFHpFRfURRLOfExaGNpPG0OSVuHju3awFj/FOHsrnHCR0ywBfyppSExcdJ7dyGo
VWFwty+/eTq2PFUUxjHzdt1KBQvQi3fg93eoItdA5hQOLQW4uD7oE6rbxXNTajsiIxVUENzR7dzE
n8TBDH1/QZZUIWYV8okrmS76yp/vFkC28UBPvGeOJApzwKScdTmEoaVFsw8ykvHF8R85dAaxU/qI
gIBs9kAX/rnNUn6QiTsTb/clbP5JIS/MN5x3vdeHEdccfylPof/hEkOeVMC12h8SpSj1K12U6IsQ
JZT9cE9/1FuiYS31GwWt9UBn/HZcWIVyu83LX/WgUD4fLBXQgFoGeAS9JCpp4VbsZ6S2DqjdDbg+
RtaQfS2SsgQ6Zw6kCTYZNNNwlZuioCOQwOrbmmH529YqJtDR1RbaTjLAeho8Y9/0b0O8bo1ttpNi
yyzaDeHi7dd7qrTSkbOtf7nqyN5WYAKWcbzOrv17AcaLsH1+qKqT0vW05D/sJO1Waj9iZtk9v2Sc
In6n96JxzR/39Rv+HOF6dDnEBzJveC+Yc/5X86d0RUdM4U9/D/FI8to2QSMbcOikzgIYzF5N5sWq
aNpRleiXD6oN35JctAGhdqcSZxHR/Mfc2E8svJYiGllwrHGcT/ZES2AT8Pc/1MJyrpDjds7etE1f
UtbUlQ10mYsFp7S9YujkD3Bc980E2gsRaamoFqMa46BkZ26Lu8sjRxLc/bxFZekRYBy2TY1AvKdU
miySDMPEL0jmdjQhvxf0rMKq1JN7veeaPROVGAr7GmyITW83p/oMM7cCSli2dVyhdTO3UYwQzX+4
M56GP8eeXFDFTeiGZjOw7+CXvHugCCePl9LlExF7ATPb4VVPCEcCMmlMeIKMtzQaMJCMLUzwuyif
7/T+BNeu7XVtG7iZ6gIHFS0PyfpBUfjd8IoSlAQNj3Glgko+euL600dVKgurHX7nieTXHiGiAs+w
uk8EDd5GItUKt8P8/g4z83ezUkKJbPhsAI8PrA/OZpAQpCtmgAQQhw+Wy725uW3vSDfjwgdPpm7G
PnVf8GJRT/rpcA9mZW/AtThIFBskupv5TFNKn2sq0GpSO16DDYJSkfzkE+Yyt6CK8qQgQDod9VMC
NjWxz+yRispCvz4ocHie8OSLxc+eUcvy5ehyq/e077p5ko5LwWLjzE0lIe1whi5ruH1+Ydu/0mSL
qY3l6USABH8/YUYLpI+/mQtYWMZ4Ukl3uI9dK+OrwItpx+DIJrn5fi2rJD6mPz7K8ylszt9sAqou
zN7GwQr7zqCmBQw6dpPtB+fk4xMVf9EQqtvZdRC1OT46dvENT+tXRDcz6frMluOyVqmouK5OXuS4
s1DAQ6WWQ6oZOxYigu7gLP0wuHuh2SdGBAys0w75WAM8nEtv3mopYy2vjT7GRZJu8fCvy6rCp8Go
C4jRTMO2capshzZ/wYBCTxkbR+ZCLRcFbSJBl56rcuQoqGms0PTodwh29m31QujAviXCznQ0nrMq
bvoZL1n5YqvlACz8g8ID73GrkIwBNoAB/4lE3MbWIiYpCQI8f84wEbEai03cN3M73n0P96FIVGQT
q3mkWfacimSnwOLiPexs2FWbglw9F9s5JXgl9ALpOE9/QY52XeKEuoCRLR+vEyyirJgVMJF5Uoe2
stc/6FCvGaycx5lq7Zf91ij/cZnjhdI4HLc/YJJ025tHmVqKNMbXzj/CydHT3IF7gNcG9E+l4JFN
LQxBIRJy77sFLvUseWV+z8qpF4A6ZEmPN3GsSEH0dNEnCO48UxgSSM55/YaRs8JGoezcL84x3HiG
9HMihPcoFutcDwywVUytZiBr6zRLoQpkclcckx5o/qtO4Uae4rMuUxPJxSwGnj3hR+j3GxPeh8SN
7Vd5jbXuRNn1tGLZe7ReMbhe7atd1Ux5S4uCr6FmkwbN5Yu+FvZgjoFb/S+S7GD8mQM1ZmO/snZ0
IQ9jV3ej/F/IDkn9OfLeijcVVNJO7Zrh5j4hFcKlvxEOzqMyt/EtA08kZG5pJaUxg5tYvNMe0/SS
ZD2v7Zc17eylpZv8b6FxUsN4BpeS1nCBqXAJ+YO6DWHCuZlWY4VeU9LWlRAx6ZAhvDgiiQ/4kU6a
nmdQKPp34sF38vKCU8egnPTlkYyEsXg/jm79luKeTg310g1HKCdVZeEYCsQIxk3zbOsmIMYQls3U
q80cxgj2wCKAVPEjRTjoyN9ZYy+wVCWuc6j6HiLlmct4c+UbuSVNfcEQ3NnY1QYN6rrnsFRVuF5o
dJfPZ3JN/1qkYo2+nEV6ycnnpkmbX1O78HpCDe2mvjOfBUdeubefKMYs15FsIl/rtUEi4XBL+ppT
5iUfAG+GyTD/XHhJ9pe+PhBPyeZGCabkZUlu7YiqN7OCPf82f9vvdytQkgZLjP4JlIdyrD/bd3lF
2/f0dRS4unF1fakGIefQOEwMGd+I+Mwb0y5tJKCMYRfkjJkqQJjTjDviKBOBuWe+pqutW4V5s9gI
ZLmCzT1s8+K1yumEeaT4Nudf1ulfpyN64c6aeuPwCHmFStpWkWek/Gzpo6l87ot4VfJfHCw3UWNh
U2hjlTchiROudmrh2RjMXvni9glZfUvf9qQ6qQspVv0ijvfto5pY44VMmF12OzU6RTkCxBz+yAD4
rQOydeJib1xh9QbsEslwzuOpJeGK3JlxDZ9bKIUeG5eHVX7Tl1a01z9fAbGdOIndh5niCHE4Jat3
8GGwYX33qbtWBIhfm+Z/kBPwKsOyAUvKD7wa/dyrxltZHIgbdZH9SQPZVYPo2Ith+Kbo1kkqDi5H
oh4F0HlvlnBf7LwLeCR9Lt7fskd9BmBXAI3BxGMgQwIKxSBJgIkvIYBkM2jux5Sx9dpbRO6Pcfs5
Mpd6Dn9lHbGsH5kLv7yrB9qwYCILFRVHccz3sVhztG5x8b6WGMe8CUTfcEqCPhaO8N3bBo18s1V7
s576kkPPlxv2O0MUJJ9rFgSIU/HpevlK9Y1EgQhuPUuT38SMcRzE6oxLIhsjqoxr0YqksMKTUA1X
HIEKXgZDIKpzcarrTk/pm1owBonxlZGZaKriktncxhjJpTZ47w9kJJIw3oxAEmHrmoOlGtQD6Wgd
9kd+FAbo4oTjOFDfSkIGi/THwtddPL+6Pn/aODBSDZ9Ib1xJZW3Vfhpxls44xbULpiq35xNU8Wq4
BRF9uCtTVHuJJv4aw5bqRmYHqSUrRMj0vCPRvb7onXkRz6CKNJwV4y5AkDeSKDt29ECsV+tj2Gb9
al0yoGMwYcGKrCitfc5pXLepKup+MaLuix6shZE4sKNjBjsApkZFl8CKhIg4rRWXm0O6UzYvH7j1
VurV4u4byljKOhyoHmLe4iuggr4aGTDVBXWKgE7jsy5E67JnD/rrGgOvO2rUohmQH5TbRsbvt2iB
vi2DB2NcyK3mpaUSEKqEGOHkEMAW3CXmw/jZWfn0qKR/TL5w1JE+CimvQhyxuqaRjENyCNrw7aP1
wlHPooQjdCgnwzF7R6k8z2bLic1X12820ZJCGV8az+o+rpqqZtDC/d3W0S/Qql7/isu53QOY1Ofx
UHEO0eYJZQDXNmHTiunLlpAqwEmKn/UQsdmP8CxVgil7RpXIIynEbaoDFSdpaShlrWDhB9jDxC5B
wMrXPkvNM5BvtMjS95OGswyS+0nzSVJGGFuUtU3fjiyE2YrdJZrm4gWPOpUlXuF+A2rOG+y5tKKM
0jn0fDHtvGlgyIakzEclkDcVx6M+NttO18bf6/bFoOsZBXWWzoewjas+I7IQkM271iWEJJDAm0Ve
Gw5xWDNII5GpxYrR0AXLNX9/GthBjb3BVq1CWse+4c7zVc59wxd0FF43Y/NzmHN189Ered/SuiQD
ZRgabzH0iRoCOG9Rgc5uy+MUzjXB/ERP8yhOwZxj4tnIqendvajyA0fBL8LdEu4VLPHVYQ+M/H+s
icChQotZEYd/6P4DHDGcQX320dK8pOPzRXAUh7N1U8+avELTwyopf3cjCeVQOft3s8MpoL4ivn8R
5hE+ATvDRoJQimEznQflMv7xbVrH4st55zWmtJTiLmc9TDmw5JIxNVHW6/Bdr17GfmXMm6ENuxnJ
iLE4HTGjkgcyhRxb8cPFUNw3VkjKtin780M/u4FqrEc5IJpp9Ub+5V3kWiDrs8j1y1saD5XnbQOo
vlKUgr50MeK2siah4q31lye/arbyzFePcCONMFsYLcfl5Lv1OaxQEXF8NWlzPKUvvGn6rgDKvTKU
UAgBybcqYQDjCP2rV1Qy0EZy9bNt2p/BKWgyjf1keRHr3BVPKDmMjx2bRPoqV/FFpRebR1kAoLek
ULL3cL5GUczrhs5crNZqGG3nd1ahnI/L2KGOrlVXP1VZlkG+YeEDIJdadSOxJqj5qrpL8VJhqZpX
udSkr8D+Ys7z8m/P8dmrlUSLVk2yJCKT9V9gXvzUkTeB6dEq5z+Z0It3fGf/FhbW1wt54nuYa9qh
INfhrTGpJf88V1ZbxsJ8s09Le8xs0YQb2pLpeMdYfZsvGwpLql8z72vYscWYavrqWBVOTuqk5AWK
M5QqdeuIPUitHxI5+D5BMOutnAECZj3/BCnqJFFpUj3nOHnXfZYK4K7aJ5Z59c4o3UwAkBD4AYQh
zDpeatw+VRxsmrhoTGYTCNS7L6dhkQcM98u6deYef6UXeDkgYYdxeSYRalC2/PCZS0cvTzBlV84T
BucQ9VJNOv2KZPtDjSnyVhng305BFtW04x1tN4tdytIZ3nx1AoF0ldv17EJw5kalRJarxkbOmJXl
xQIG3QSQwL0Ihf/3fqng2VX72wYys5U8Aj8WjDtT+KJgaZP1mxtxVlKSOmeztZrSNh+vEMDfNMaB
Pw6DHufXm27w/F0jgzRIf0WkkD/XqpDQbJiEJv9XBzTaPgFrI7zGtJ4w1dwSPKJa1nbYCMdn7e+2
LmWE0kLuTnUgvHQ0IdEsJrPvTmh7fZcPCQCcRXlcPwelVBMSsc78HQCnuclG9X5A5JefJxav2RzP
sCgWxuCp4O1T9y9zfRhjhAkoQ5EBfRe6dC/IK3TGFJpmV8Pc5U0cDAK7qmiHPsIwkgqzb9SQ8LxX
/XdilyakBvQsQhaEBOk3/OOhFnIr3oZSk+BTFzPTRxB3H2VdGgaoCRBju+iSn4IwZ3eGH0xd+7MC
DH2RXeCDFmtrYVSNfVTUyhAxiFWgLd1VnnwbUlPGN9eQFbGLm7KYZXv3Cc5d8TJ6E9Cfv51jBmns
0p916oz1Zn3ki8sexwsPMPb9UkqWmy2mNFch7fvrQtKvd7XjDnCWXRIo8c2PxanTJUEjhDQG3pSD
i0KAlISY+Tho+zYf4fIyiR2+69nPGJ6mWPpjUbNe3gwpQa9u1u1g8g/6dEp3eupt6cYwy86Vwoe3
n1mZUWh12Y1fEE0lCDn4ZFZ7QqcZAI15uVOzhsJKGmvp4qxqaioVWCf8wVKBsI8tYagcm9UcMwoj
23lo9a4t9NAJ2+Vsf9qUOPJdoquxOGQ6wrzX03V0cBSXZoRZdvFnqDLq6DwRg2hyPFYB+oqQRmHu
+0oUoqGMaONDbdd4weGRaOGLqlWl2rKn1tC+x/XcIvpFYhxnXfi1UzbSY7Zyeje3brVk8fmFeZ9p
BWV0cq/HIllxNR9NKMOVFEQl6YAJBijvIQYJT8C1olY8FaO0o8lWLG5AfYyKr9XBY/EScQG1tBTu
sFNLUM3Rk7n0sc6pAuqZeGFUjjr5OqLxErzZq76jYT8P59uQc0efgJPD3+61v0kC3OPhOR5yhjLz
1w8XDvcTMboIgJK5bfdZ2lZbCb2ep/hnfRfJ/mClZnGWl0tEeqImusvj+jb3U1C4u0oHkVhQO8GK
P+dP3zxYr9eV9MvdFDmPSKU0o6eQsHvra0aVpJqQPOCzwPoateaMfsE5tXRG9Z6OIYbyBQnOpyCi
lQL52i9lHkSVNzC9Esih8xO9/kichPGcSBVRSwrxcz2H5SmPGVEWORvdZGD1R5FXJhIdNYEEbYmc
BtmySyJ+ZsqnXf9SnRSFnQkZ9gntUWz1kV1QBOko3Q8xLc/ZoEtSgUbPu4LYGcxu9SCKK5LVZmf2
Qp9KipdIYyoW+L4aoFmhgGZXC5qDo6dxoTzYlVN0KegCNziOEPBnP9xFp05EZN21Rq8P7ZpeK2RJ
ZuK/mHr0J4YpvHVLtSNS+rqbLOMOOdWFHKZVFd+XKRvnOiKSct3gbbec4DYsrTz9MNV+2EnuzC7S
eLIMKFkP6fpE37PyDm8O3CULXgNYDRTRbQgs+3T9A1K/YS+dapAOu+cRNmnjnFGFqlYLnNsT371+
I0Lnt0J0v8YKpjiARF/GKnQpM6AyvFmg1f9pwNaaY25z4kMswdvd9tAHgwlobgMHSN/OUy4/jRLp
LzEgQnba2N/gDxz/hnkoIneSFmat4eS9pALklNLiRjlE1yZe6a7ygy53Uc1AQHo1hg8HYusuegzA
zJeuHMGPrTDJbKhLKubrxmF0JH5r/ca+XI8puuhO83oEi5wAtYFFJ6eLfGo1+RVo8Y7EaOALiw9A
ydOr/Z1igrC+HDpfhioEgLJJLeMwNk0NX5BPI96O6sHMiBi1/Pn9CqaFyhxmZ0JlNi6MGKRaaYu4
1ZnCzxA06LsI5cBaTjZ74ZqcALJqEyeSshVBy+AEmtwoka5aWJYRlsetCm2HDB/69Hf48k7WwlKA
kbSXGO6fnioAsNQ3aOeVuDY4stfMBgx6q1pUP7m+Xs7QrPhDzRR8H6DbQLaVZrVPqW5jHJLyAM+6
YPpDt4fqA5dj0EeEQfNioBDhEc79UotkvLBWozKgPOupon2avu2CgkrsqvRo1WUR3NQICfliHjAT
caX8RrHDAy0Gpuo9Z787s+nGqt4kNc7J20H2a8IT+tQB/6qKyyvPZtrKt4KRoruzddIaXRoEMMJ6
MB3giDf0lbjNsgTrKj+2s8ajdbR63gtfHIAVUSZWeh+sIauV7M+GZU2sfVzq/3uK+03egqe1TBhQ
rWko0Pk7QGB/mRGaLWqIU+ptBR+WaNUyvCmvnZpQxNrLG75aj76Nlehg5rnAE79zZ5H7xFnAPEsM
/qPUs4mA2hatAnsee9XWi947dnFB9zXFfI8vPJehoPHUfAjUDiijo+GFEHmAMjMZF/tlNbIxr6Wt
n6hzw99cZjnUDsTL7y+uhbvPiFgCGf+KIIKNTFZq6Ya+MHA8bKrIFX/3FNa2WBJxgcM9ptpuKGV0
4t/HZjR0ibopz1tDLn+jki0JL+EABJU0J+sT/jZ/ZOrp495AzFnqlyqLqeW20W5DmDxfiURpBWTi
ca9L7XN1cTdd2eoIsKIyNxsGPtaS8FgCMLvAdSRp4yaazkzr/Ly69ul47Kui1zdIMCNmDi5ybSTm
aP6xAKwT6dlSmJJUaKMn5uXvo0stLAllVgbYHUsAOARGDHHyHFQ+SCHRkrIgppYtAlH+3xfvU4nj
dSEhuJCRIMoJvzcrQ/I9EzdKOEzzaLfmnALJdcGXjKCeTZAsAlAzImOMWgO+EsynMKngN5CaOTyF
C2Cw/KmZSbO47TnJhw7t0Z63tmCYh4Jk5H0ipppx2sv1+fsTLa9RzoGUTpw04FKE7T8FI+kWCO3f
Qq+CoBfGE7QyLOF8hnsJi1mc/TqCZYJPrKLzCaiVrnhNFysrmnxujCDkoeW5dQYmSysZaB2KGEZS
tmAePPgAZpeCkv7azx/BP6b+VAa14pi9Dl4mf7QXneIQ3Ap+1z5FfVZET+k1wFSnjsFudeut7ZAp
Yr87KuCxleIiubzz/5OSfIGLWHWbLzs3M3p2l+jhiEwWnOCXEuI1H2qKdaYkmpNeCrkt+vS13kfZ
yBHo2Yke2Tn1sTF4L7gvRgSHlj/2JdfHWzCvA74VCGm2WksPvpVBKNE/pLFL3b3XVCVstHSVOuPe
EKwg6Y14kxvQJ5dJlj+przHzzqji8ZDAj68iKQXwQ85gPIET3XWnqrMzw/vvPhup4CTeHLfCWA1J
n041UumG2DfHq4FZeOAD6hT0BwH9eyyrbPbj+zvQu9uRr8+sLnJng+VHbs7PfELCWIT5EnCt6iiT
xzIfGntuXlY+5Vr2nVqmHvLYtThYb64zfd4ygjvghDurmccJbKznEeEfUV50aWTui3JRZHjzxvqw
loZJHWcXbQXKJSfHG0xN6Al5FE1FzcHavkYyPBRF5dM33GAgAqxHJ2TBIWuou8UM5Ge7IGuaXLwi
Za3G2FZ/8tFG0d/YWp+DCAeN1S9EWLNcwLXHoFoghHjTCgqwMeVecaipFe8BSd++TExdwPENO0ha
PoXLWu0b5HlMa8bzYJEcLLZ+0uzkcFe10Ey7+cPxteinDFRLojpgOryFGpGhYiGsNyzxl9LgKErj
Ot1wur/QKwzj0l10Zb/w3ojn+EjQMlXhIEiybdMfIBONV/1QZukutcv9rZ6JmjsoT32dXOO6XOyy
+QGJEXZwlZI8gUDH0ulCgBTc/q/QNqEg0vY9Xh8wfMjgTH3GXKInvPf6k/dfyvUwyEQF6PEyGDSI
zpUMm3CGI9r+gVrOk/bZ7yQb7g6Bv61Cs/GMbcgEviXg/fMw6FtqSs8TJKLRh6LL2cyEj3xkhbPT
sL7XneilInNVTYi/B1yUtIE5goL0W8FUjxP/uYbYrT1vPo2KYSQ1xSafTOb/N066vtR5Hwc/Nzz7
dSWA8vMoViq312lsBGeCBd3z0uq2Ob6M+4QNFJm5MWmQVS6DrT9kRG56hLFwnPJx9rP8GEPpC7d7
n3gb/r7jgEJQaAp1yX/McatbyRxUDLFoheg0UaRW8onGTxe2UhFttBttBJYNbcvd92o6FhnwrHDk
n/XtOpboMvbNRJsoJBnIy4lymAftxtB/Pew/QMXiixn18D1hHVZH1+s8n5kv2xSmRAm6wtZewin+
6yNjJoUG577mB1dpNRLadlnHbrrBTX2EkeE3wVQbLbmx9dcjWLbElbfyi55EhwD/sa8QUREi/v6w
yenfqnNwHdvDbGigbcZW5tLxE3ufA5wNkpJmtwDNaOiLPZmls7a4Az3zmEcVVCo76hvS+6mPHoHd
FisWtQLLA0AAVRHXjKeOpo9jRpubYgNZFwUhPNexQfzKwcO7deZRNRrEtubxq2JM4NTFYqx+5sPO
sDM/lpHbAHiJXur7KCvqFmqkFbis9j5SaIYf++aTGVw+EOCwF636r5a8MH/djs5Awy2rnGWHep2d
qe8svO7WPwm9zqVQcXix2jdaRJACJDGMwkXoCNUx3YTMO4oyYJ3X7bpNvQcv4T2Cv0svJyPSEPaq
B3OyM6A6vmHU15MfC1Wq6irN74c6diRhBlDFg8wK8J8f4MYN2R8tOaKDO7TW5kzU3EULbzcVJ8ug
lhVgUXfYrdHI1ZJ3PGxshgmb1vTOVg4AzjD+LAE3hEHRYHxd1FaVLBqMATuHKAFtygLOTUSkjbcY
xa5fYfxkwR9pEXdLSVtxHbg9Z6VvKetBBzITQoT8j79VIBITPXu5BRBbW69P+A0JTnr4J3D/Mrpw
xFljksPmXq5Xb1mrMX5rUBHuMu0CTCGZXKX8Fl4uu2KNMhy/LbxZBm6BZaRUM+NRck9ml8MJLgVB
Rq1g/zNNTwoThCp2lvmbTzkIsTf14E4ND1KVlZeM21V4lfMNaBTGOK/XRF8/Y6tnfRJw7h42h0nq
5RF2cNXkpKsvTJ7wuQ/2QBQxfOWeuP/7yz5e45v6zP/KZ7kEen6GBAFEkdafT+e06m9GxIXYDBx5
pwRLE3yIwSe9cpu8FviWISeZAmmZx9fVLOJovAFNasJj8z9qY5fhsXmmNUzenfOvzZqH7rxYxsAO
IRrnLSE7HiS6ahpbPxPSmkBDPOVycnCSpVjywJlxqM3Yym3diSt5ISCwSJ37fxqTBw8z9CZE5Y4r
5CtvOA/lzjSSVYFbam5QUiejUDJXV1vbBf6ppscSi7uhrTamNHc7n5zy8GKVz6TCWdea8sbwr0+L
WjF7t+ayakf8pvqp88ugXL/XBMxXH+k8aMltgyZaP2s9S4NKvAKqR2gkCT1Cuof1qsRTD15R5AVD
v20NoxFi2l4ovv+hk80miK63f9IlYr1DLFov10bWdxEeLT6mssCABf42xh3bS/7j3hpaT//cYcpG
WzJgcwTDcaWK7reDJ78rEwXWGlSE2wtnlHFkCnNy5nbyV4woY7x9MvBfB+EV5zgVCH6hwd1M5f08
oXlXoEfPmMaikWDS6+uK+TG1fIqheonlE4dSiQFHP+guUk6aSAYdxFhKP0ZSE2C8/KxWCfYfHJPC
n84/NIzxpZW3+u2WqEUGuRNjUc/Ae20Zm4nqPQrb87+J38nPDyvwpH2gE94pt4Mo1hdISzHFS8hH
4B++4OqJ12WRAATL2qvN3wAHGAwLVU+7FvpWkjDnmxa1aphQI4L1ICb0YY6cWolL+yW/9UoNGhxu
GX04QkL4ST7BRf6M7G4Labui+EHdVK9JhKzr/iwb9/tz41c81hE3QPNqCGHSZeOFf8fMJGMmpe9D
5TRAONrdS+JLoohSFqge8TZb8BDLdcxo3DP9HpyqH7Ls7hsZ4nz+hj2VuQXkOCgXGfFTNKhMOiCD
KYprGFb0EHbHJXq7tchGad8KnPTsQFAy3+QrYWpCPgJxwYbT3ms+kZoaPGILQtTaPL25Bu5FsVLj
MPaUZd6c05A5FXhPdy8HVBHROoeM0GI42JPLA/BlOQGA8Q5XmOTP9+Xq6G6xpkJJIJU71vgHiFgb
qLTWa5E2Ubr3yAq/tEU2oI8FYzbP3xI9nxBPDzEcdjiKMvV68v39p1VJtiohe6XdXUo9SLx+qacK
uRzi0mPv8Xw+4Yre0be/lw/+UWRuPwNI3ohtWWuifVFRatm0pwGiqfHYjYmNScbcGFekHnDxYCOM
QXodvGQJVdDYlBBh8MMejbLBlrewBuuiHHCWIe9ckEb0sjsSxLqcLKaANF5cID0TTnnX4rtav05+
0znFhyH9kNRlsw5WCL+R7sG9qt93ACrWtg860ole39fk4rVJdG0k6ik63dzb89rH68DVNqzJmj9K
IgT/VFRZrVsogDYdNw952hOJujyM4aLPqtWErM4f6dxLGbX0POa+60BiUlkQBoX/ZCSXAsJ0seua
ehMP+ezc4fUeJWqZ+u4WjWD345ZpoNZwlD1R85K4qu4NEBIyo/X6ipZQyoegJAJGa9Yv87tOHclq
AzKY9cEdws1XJao9OcD1hxIu9jtAdqmnNLGY97lNH81H0+4nuc4SO/ciy18OGkTwqI2hRD4BMX0q
FuikNNAY4WL9bftZmfxhWvTpcpKEuRCFJgEhtHyL8kOacOUZnufuFjL6GU68wXEF8Sbk8nlZxKZ1
0TXZqzk+A9d12oXp2QaI/PXBvxEAaLuLorD/0nE4gQCDb/uhqvJlUq52nWOGqxcc2W1l3TzosMzJ
64B61x2CBAm/9ARECGgn0sUX5eiwRVoEYym+vmaEQu6sMRkatRPCaOwwz4aWhGZj+TVdmoayHPhA
ygM60ieKUyu0234zpy03kDZ89SQszZsR+dkPVltzklOvl3AaneAeybtqpKBcw02Frb0uIfmjLcGD
MFHUIci4RFnngGV0MfhTpfCjmwNQs/dVx/ySwJj9QkZtRH25lTEZhepp6EhopjIHz29/yxXbDOsN
AKrc8z5+IgJPlEGEKOx20Py1tiQHDBIZYGEukEVthNPojzd0zXsyl5OdV1C/3NlKGZ/85KcrT163
OQJwFFHU0AL/bThajCKqe0nElnc8iLMV+quhhw7e9qScI6qYLxYrv5HnqrVBcHO7zdHfLjODB+cj
OpnAfzY8hvOWdW8M6TIBQMFBJhrQqFMmJ3MWjTFplhifouO89o0MpZpKyDuQ+7FHH0mfsAYZkwyu
ASkUpMoPHsNh9gz1Ltw54Z/vANSbhXq5uqsK9lVATdbRF3/FVktFUWjVHpIx56uAelsOjj0MmeAP
m+p9DWOisZ6WXAgdkyk4aXDVnZBaqJ8i7yrrGAxFRX27726Hm0KoEg/Xb9GnzYtjilkKex+w1jJ2
AfwQ6ModKcYlGmHZ2iI/bvkSs1zJYtXcHa+LErKIG0h/kfLGI+zUd1SznsstEmq+2tpikygBvyjy
RIaXOqzmxBaipA4adkhfYHzYRs36vE5s1pjHb/gG69s0bi3rqwhS4K2cUTi1w1uetZ7ohekrUzfP
9Yd5amFBPxlwsqLHhUiZlnLmEOXDsiWLgxPDobclSxWDprCYujlssjWaTX/gddJ+BeZbrw4+shDE
flg+p9Zl8szNtZxqu6/F8bqkUBvV7M+3aPUDE6u+f8NzqPZrhTrTC1mZQBD7YyaEs4CcG4cRNlYo
JskuRl9NTKym5WiWH+h3Bs9I1B2MFnhD/tUs+JKUJwEFXV/Ar2PyH8sc6Mn/CLW/2szsrfXFTsBe
7wdFYZK09grLBsXB0oZJD/mbE9Edx4+Z831TynG3VqCVG85pME3BeucI9/9bh++8PzmHeCk/C39c
UW1Gd338Wakz+Ua9/s9Ct+RwCU0vS1Q/U9QZ+Wb4v5VhKEWrT4z8eMJFXAEn5Wa4s3dSvPip1UOQ
YqrMFPxqBt1m9q8Wq5TnVPgzwKF7bx6lis/QPl1UAAWZk2z4EsYX7Sk1/55N+ILlq8u4yrQ3sCIw
GeyBQHcqXpncUCq4zLZp9f5RQJJ/lB8ZpMECtwPoz17EgaVod1zvF/zvrlhmZnshtYRZIi4dYGNB
PaT1TtuemAdNRbWMcaOIu+OqxXp0kDflAgDZTQKpkXKkECNl5D4ndK2FOkjdw11QsNNrVRIAcw+U
U19SnfyryI1+PI5E+kJsN3fZjkZWXyphrtS329eygDA4jKcmQSjMP2pc/Fph4tBE7capLurZs4nP
gpgdr4HYstr/pYt/yuEtUeargAboAYV7cTCq8Lw/+zhgA82dws37gewrEBSsCFzQLsNDbRm4D9DQ
RaPfuJ8tIwcpaTd6GH3CpMoDknGmghjtugeai9ulrFl/trEu9Eh5vmKIeCeU9T4MJQDt+qalAB6R
crrOTM6rrMU3EmVyPMQwr8h4K8tfafb5VLIoZiPIoxo1aQvpeilwLnkYyjWi0ML/xqljap6fTBo2
Od2VMfOEqAHlcil9srz4W5xXCqozFsAsDrk73XkAYoKGGNxVwyALSisk30OizISObN8usck6WbK7
uidr9cKlkTvP9UUCHJzBH/nqIM+S8uH2YOitSr/HANTIGSPVMeH41eQ2IUENJ0saaNU7KStEPeWX
gGsRQRyxlaxgSdPQyoDlcbeo5EGuj5s6FoHwc0f6teg3mY3XMyBz9de/opD/cEgKtpvHrgi6s6Ob
cdVv6g7KTmVv9vsKPzulyHm6s+Mh06vdLNY26U8ZqeHy+NOrdcfdHtrDbCRiYnE+c7rHduPoCEt1
g2cE/6AMy96cDgEtxK2FXJVqVgxGdIP5Agca3My3XaF+2wUtX3yhSlEap2VGQxEUgrGdn0v3KnDX
gvMPW/S/OPZyszQYWwj4Jn5Zj2uZmBC0EjiF2xMBYx2wsbLlIHpk85xTX2Dp3CmdSYfigEzSW9No
qQAhimii0xRmD4TQkv+NpuAmrcAgYxyhuHATGeSS6/1EZ2efUIpPtXq03KsorOZYa+ma49l5mwKn
SHtsoFqEAMbfD1MB7LOeNqG0mzJC9QeFhunyJ07CLCfmVRKb7UuMEQw6iHN1e9NyVQCaD/K3N8Rp
kSDchmGEqY8Erg2//XFWSUiI7oK3WzdIgG7HOVaCD8meniqpgAgfRLctIBhvOLuOO7hJvIEtFT9X
ee7J0rJt+2MTbTuFgbW+KRJhu2nKCxl2eMjPfi6INg6B3q8N+yd5vEL9+gnnQLtwKLEKN7ChYNEc
r6fcjeSYE+nvn+Zjut1+/DQ61pr1DN1cxTBvmsl3XEp0l34PFx+xCNfiTueIypjNPBNwLc3MxxJz
2C53vuzMhz3LT7pVqhgHIqGaJRMPr50BSPXexmCiGGCGKMAjYqSmrQMKhlVAqNv0G/jM2e8lKDMB
3AVkgOSNJ1Uc8VYAAyDPrtr+MzehMyUDKd+sIlcnKb01Xp9QabGHxLYLG17q79XGfLfGnTADcVpO
Mmx556It+R7ZCpORPL//ekbzmZxpiKhsO4RG73d1gaOzNQeAercKdPEB339z44HqXW231LYAYGrO
WZrfkfaJda89zJO86mn8JOLamnjwn9/AUhhNibOldEaG1AkXjPMTYajzqdlRg10Eyev7Lk57aq5/
OHywXNr8IlrNR7OndF4A5+YsPupQyg8lhOgopgAN67H3J1XeAcJqDCsHCiKvLRlmNGAkKHbxV1/v
fWigpnZ83IWjLH1oesQCWkYdD2ETq6dRDae9Le+lzPvHLExTZcFKt2PvjISiDAmeY5TTyV86iI7I
p0WRtSiOhlt+DPoWSigGR1Y6S6q3ra1i+sfUaNeyk/l+dByd1nblTaMiexOnY0IMJD+5FrDQt6+S
O66hFqxdoe+GdQAlKMtHKDLEljB1T9aIbCuhM2ywk1zurnGXBleWxXOmbxFwUFZbPk/80UQAjGAx
b7v1lykajVt2cYAAREmi97MZrwsacUyDiMXYfH82mz26hhbTZb5jzATlzPUFGFrI7HoZwqDo+sPh
9l+T3W3IxPW+Mwpj97PfY8qKwKQln4i3JbubtECsB0M3WSfp38qfKZ6r2osK6RtdkY1gtaWNLe6V
dtBVQRExlWEEOmJEU3nHj/B7a1E1JxnWDiIssYmopCFsF2xaePBkHVriim/tdhV5HILkFIEeI6Dv
HXqOp9HJkvowrXErVa+NhkYMKpICwDj6eJsHrQd09pQwtWvqUBwlW9Zubhng0n7Z7cBs35qjX8mj
7E8t68K6S6G8nXyGayyxHEjBC3WEZ/KSHFf1b1NmF9JiI2at+CJZgbv+Femz8WHy33b+MJRUJt+9
1OwItoQijTBQetqbNuuRGDuHEtWmqVd4JAZpgzAAs4n6pSNIOZ9J4Q1HqGRUpKzOXXA8CTIxtCXH
iSxVTxjP+MPdW1q4ltwWCv6G0AZRL87Q2xwrN+GGPwgFA9TVC3aTkUwUay0o3slULXtJMHOe82QV
UoJMSSvlM5oroE0xYsCsEaSRgh3ltZoWBGF10LRDadOUdLV2pT5YJDCOhBMDRYJBqlPlAuXPCgzZ
hYUF+4mL5bcFtGRx/BlGcMlday8I6MuitmGJf0ukM3nFn6qrXznFCeql1E3ySF0pfv/K0a7UCEqF
DJK4F9Cfn1S6w3NF3zgz6AwLkV+OYGb8F30aSZrfCtIBKl2Z/FzlvS04Yc9Zbgdjf39k+alfpQLo
SyGxwaNmEBRAg9GEOq+wgu+NQ305UcZmHc7upT2e3iqwauhMBxb2zXFOddf7LONPf7CKBcpLUP6h
/HE761j2w2AuoVR6Y92rWRZjUcuqWAl5SgjwUI80sM9eH/6dcDelajTlYumZfNn0PTioUP/83Qgk
X0cQR6uiX5/QAI9IEbbuIOols2tO51g0w1eJ5DwlvMTWrBhIhmH4I7uJFs6eXaPF/FI68MYWm8Fy
mscJ3l6FZ1NNG3oJIXUIatXmsOaBPOM3jh/31DnqHJsn8GBRnxmrNEj1Kh9t1EeMutn68Wn+sDY0
ZOjiN9I+ltnxo6LnseO8NDK88pnOqbd3KMSP6XqafMqq3YXQoQTmHxtjsGEimWWhuBOyIzmcC1Qq
JuYJYpl3J1vWCWIqqLtVh/uCd1d1YECg2ukfoZjHr5hD/i1pjGSw8V1UR7IIP9C1lExbaBJMVs2Y
K/ufECMP/PHCgp/7tBKLI61f8NcqwnJR5+FSBtBZokJYcOXYRCjLDlLy1p8BgmFFCylOTKyik+Jy
1eDj1ats6XqAh2AKc/eOkwkCbS+RiuJ7PWayq5PNxJxeH0drKeabSuIwLznEtSH2WQv0zXYt+iuY
AW+gQfZ1ZbZhNYvof2s4rXU58vMg/dPyvXcbntBRy+FroC6inG4DOSo4ZRwLnngnDVBrNmnn7k5c
Wy3m5nvXsIHgaC3tgmvQAQNcmahUwUVzwQ+/v1qBCmKO7Cc3Yg++KgtPGEUk8XD9gQEB9PDCsHlK
Eq0LY6iWtvpyE7f/tLFLs7Y6VJsC2OCB3wg1qkPjDclcsRlPG6hHBSreFCRSMOJbu/jv4CqCCOGD
iXTvKXIlLlOcmVNYnxBxEpQWktr922JmqxVBHVB21ayQcWtMZRgAllCh7I0uPU+GnjH/3VzqU/3D
jDrJbCjKwYwGETZiuwv3BOG/xJl3Kca7J2fsU5E1HlVPIu3Gs1U5dCfLaFykFfje5Rxnc/xXLpz5
BmIVSb2flLIWRHsUA/LyCSGFm1VRz/QQ/tueLAsXnvqH3idFa9+JOo2eF1q4FRdXAtcv4610xS/f
iIlGHx/h4aohhk7xxKRSzAQ/puDkHTSJi3sPpOMs4uWkKVkcPnw+T0kGPV9qpH11wltA5DrK9xr3
u0QBA5R9qJZYsggPo5g6Jw+V0OmcmBj4orLoN+c9OEFaXTt8zsRBnngHzKay+9pNqCMfd1dB6uSv
VpAkEq0e6n9Ki0rTr2O5gBkyunWjZmoElVgKKhhd266tNQ/H3/Fa4xfVd4K5w+u+yQLr4hXFeGPO
kPSQByMsGBJs4dNI9ifRaXCxHnrG9XSyIdV2AY76pA4OBz/o+Evn43yeu1OjU6kXWiaFPFehcy3g
QDTm0mcFFJNf6a5BEoZpDFYlxvbl7c0eIaGIGIflMASfB6n8KvwWkRMq5fiJo2AMxlRHEaop/sZT
Y43WR1LRyNAJt0sdBJJR1HIvOxmL4GW5ZN/wi3tNHH/0Phue5B5rpKtCztsl3yogXGmFqf13/Q9l
JeXwrOg6lgTROSPmmLFDWyg79YYv5doA40FzPLSKNI9emNkCQb779VsEFNG/pbOdSJTLGrFg0bAw
slX0L4SRAsFRz3yri/1e2hVlezRRVoIHtbcC3V6kB9pEl6C4lP+KzIb826up7Icx8QCNoi226DHt
Y69uNOGjIjR5gNlgeN2CWZ/tdEMBi0UZxBrho6kfkWQnH51elpRqPjikMpLjWvgVjuPWNTW6mrps
hP4ChOzgWe7uFUSk6LnVjiO3snjyR8lnBnEfeumdwTlNa8SQHGJhvmk85EJbkgjnNn+Ahj0grFRG
ak6X+Rp2WXifea2NEiw+f6EJF7cLRs5OnOmyWCoNDiHlO/6Us0WAEoLSGAnl39qQ+Ntl+ch5iIqM
FjSnuCZ33rauTI2/DRWIbPBD6XOYYEvaNSCk0ZpYnTZdRZqJ9FGoE2D5rNdNFqe3OI6F1K0BR/X9
0pqq0teHzd9yrcxiWEvyUYNYiN0UCfwPDNgYn6n4OJelFHTnOrPPAo75Ve7Xz06O8OAtsilTCsHp
GzELG8AflsXrpgaU05p41j67cKfJNVTuax6Kmv7zXofGeuxLoUMLITsw2dZOhTssvn7ZqBNCaEZy
Rt2tH8sx5sgI0gDMG1zW33WsIAO2FsGkQkO0DiM5eOCa6knhJbM+mavAIp/cst37RHSPiW8pem07
NZ4gMnfdVm348uzmF10Duur/UD/2io4NxxiCt7A1rc1aD5Ku+nsM0OaN0bj/qRS6FgTq/Dflt8w/
Bp7VmInqv6DKJYDtYzvypqVxM2aom53E6quP9nwe+zpYB2DJPJFf7lskRCIx6bX+N9WPshAAqzOj
mRxhubD2ADubKbV1gQjGoTj/j+va4LNZpbFr3lck8UX4OO85N0S0VOBWjmA8G5g4RiAJBlr5/tt+
3DPYKtJlhufSAmWgfYdjIlB4ayMPnz3f3sbS9AXGMkn6yPsmUMXJNu6NmWor6hUG9AKoGCJ9+0rE
9RlpmPzIKKEwCbbLjfw0yFEntzClHcZiFD9p9pwkosanTIEg+eFq6sY1iQoWkev2Oa5Z5meTk4lE
yXLegUTZSAA3zvvzum4k+kPNGyVBPid6Wx71ENcW3qYbgjWsvQpgzOnqBRa3vyHZvJ8NiWtN7dhQ
q7SU5YqAoIifW6yVT5falAVygF9yNUntX7yP87ZAHsUj7I9Ff5//VY4VFd2f7K8+U5z94PxquYAd
cOgpWLbSZVePhe//rvccQ1TCtmtlqiv1JZSLcC8Ynsy8DrqtcuZC/FZPPWE6z+l6SYcCAFzSGNt+
uZwYREV96vXgtLX36rgTx4/XkkEwogVYw55LcBRBr0j/nFPelTt78pSfF1qkrNs5NQYUs0Pbw0dm
cePf5onlQ0iMQ5BrvE1KXzBJTt0/iSer1PeqVlFiKUEAeIVtWNL6Sldd488ePCC4rIC3XAhRFHQ1
Kb271Oa9ahm/IosG495pZd2xBBJOVFqMwMj+BGWuXeRKbgQtNMHXdLleReNp1mpETARpM1UoSTWU
jIeQMsgFa+FZNl7fTbSCnVRMkUgRXO7H4c5yIsOCGEBhz39tIh5cSik8xDrS5vkG7FJMmu+dhWx9
qQkLr3qKIdL2QxFKaveQVKIdqibuO2GGx60cWvi9mZG6orVW2RwtEo1NpQh3aNVspFy+GqO/mYN+
NTAgdZiFxJCjGN6RCrdSuQ2zXP4/wOlOSOs60bDHpf5JgYYuM4pD84/+9u8tymcAK2w06vQFK+VF
FiI+N/xnpE0NEfyQouEqisRhhLmq+iQvbSOA7uLf7OhFLI7/vGhFSCo7e8ZILc7weNp2Bm+1fOOO
FZX6tk7Bm91jKUVBoYa4pTJDPkOm6BlKwHwM/4XsEJV+R3C/Cq+YeoY8HEq8p8LvUqaBj5dGFvas
IvOAcRjA9P8OXt+iRGosRJYrbCRDt3GlNDrds6MSF/Tm5/DcMZVJ08ZOmbcGw10Shk5hItf8krvg
DxDpOdHjZJA4TNHvO12Q8wdaw8fUyGCkmrnpCGlzKzZUS6l2DWfrVdNJy7rLVcDb7pQ6A0XXZzfD
WurXwY12BBtQQwPh78gQyMoVC0q2WR728MN07/d43M7g9o/jbGPAWn39JThK/sHG4cpVAVD6Hqbz
03ZF/sQkSN3vVSLywMyFNBE+sTRWOiYfSA/e/rs4GtwoWV4rRA9XJfAQ6VBTM/u/bvyEIsgfuEFx
q2g/4dhwPYb29fsCFxCn45nlL/ridUwNiT2nZGLkSzjLCOdrN4pe/7vX9aGuFK0qwXDfDsaOByV+
8IAS0Q8wjGv7bUPRo0POAME6VosVrS66DdVo7fG3GZnvNce7eSjGm7E44lyosvLFc4HRViXyJTyV
dovi1Fi7J1e2F1ixWeyT1E6eF8sq1eJB8oLRKY5FsTKiZR1LBqc1LNjphaBCJKbbShmp7Cl0Cu7F
YlByv0+KHR5kdr2JblAhTCi9O9945Pe1TNv0f9Ksg5bbbN6SYq7R67X0xHhH57pl5MFB97AOa7Mi
vteJs+TlNjCw4M8ECulXFrOvPgugENWM+zreLqHwInxxhh2J886Bcacc5kmAHJW4eap2j+08bdnn
ExlOO2Kb40y9S9o3PjtR1FPV+R+EQlKZ63a3TdO1Z3AN8VBcBt/sarZAF8mHeOSBP0G6W+Bfkdp/
q1nmAQ9lsb7y7h3xOHB9MwW6xO3TKOnEYSyMSyR2SKj1IBNCd0JAN/5/wu/23zYPW+ra/a4/f8j6
mRbVER4lKYe4/yIp26dLTtdBiB5DKAoCCNWsHK2G79WyA4/qc7RJpuDdBkKUTww2iHGHrYmU2FeE
zeUEY1/xliBgJsAqYfOqM5KpNKOqxu8OxDw+VBBuIi+QWrFZdv5Amvd9B8I3Oj/p/8YMBUG9c1Cj
Ng/7KpeUOxz0VttMzojCiBej+cdCj+eXWyJfI5VadZwK5nj6uIBBVBbdw+Hd2FLQoyO0SFt+Jn3+
st7x1LMB2H7f4UvuwmxYlxojZLYkRbP90MRwqZHA8cpzQATsJhskjKK758LrL2g3C+aLiiKaV/95
90gf+gknexTnJoGv8XBKdeXJN9R0aDf743m6v6Skpz0O4DfUIdI8+ViuESl+ir21qrZxU6rHxn1i
yeqdlREGe4O3AfcL/BvUFJSM6wgs2HHeYyKO9lS5uLragPhgD8V7jlG+J8ECZ49yAvF4kZI71THn
LsYhkatxAP4/dwYiV9pJRR4vT8DGcp484Xi/OZOF62yRtTZGveUI6B2yD/tluh/WnnR4XPYug1pz
r7PwKImiaEu1d+e9khEw7oAmYuUmR3H4UMR+CtWyeNFOjntKkxFoecUppZsLc4g7CTDcONdxfpdr
xiq6gnNsQR3PDSbwlkDFzgzdREMO7nOVKTyVpn4ABOnUJHqHkhjGgtPR11G+sVmsDA7gfEsSqBdT
uiS8V4f8jfLrYIBzww89xStHMMuT3RGJFoNEqv1NSzXzBqxgVd2CC0gmRKmVGNFZVNDnBAElbT3G
APQmTcz/iSL39xxBhocWVWyzQvcTa013iwkZZNp22rwSvwiR+foHDBWzlhx+rx+dEAsvuPoS2iVa
nUkna4arzZeL5HGwb+1KmOW4jJW91P7IBJBItBh6LvXqenL84SUktkmsgAEcgBEzd8hRNLSF7bT9
fYfJUVKRjcP6l4blcJKm/A/HdMYAlezHW6/FPEfaSYmIic7iRZaFX+7PN0NjEyzyfF66aZmgHfIU
ox8azJffqOKRRQOv62y5rA0pf2PblZcH36metLjO5lLgB3oGexlIefwdFGbVAq37AgYX6BteGUep
BwmbWjGMoxQrL/QEAxPz/ZuGuilOeDg9VXB2vQCUCqrzoR6luPSNfF7/8D+CgpkGGHNLEgU2IUPp
Z9r67oSQ5VfBkJ0Ps5hzHQi4wn/ubcaj2Q/D8aQzrYTU52d00dIUxtkJiBWgwJ56vv8cSUQGKih6
XCmtZCkOXOQ84RlZ9JqqK0RGdpNz45f/cQzQHDyXmoy8YZSGl7r98sJaT481jojES3FX7BcIm36r
3CII4i36Zp1vw7dwBJ6CjISjyx/ePvrKeFUBYZ9WWLwx2kq74EPEHXiqNVXLh0IWSS+nc4aRjDuS
jJh8QqfYcpD6FFoirZLvoAyDTdO8tXvquuKv6Vy3U1YgwkpcrRNFlPVx6qrb0iwO6FXZ5u6DKOdu
ECi3F5G8fbx7A/Gf7tj+/07jcrsdqToWyIzjKIJLW+gOZXp6nV0D+zD3M/WUlzAH1pVXCWyIT3sB
AK42gwyuO8rRKdTYMgHnjIkcWgf5MEOsOe0jj2lHFoHCWgzagV3gi45o/4K9BuQrib+dY0qSKK/A
4k6t1gOfV+xsi0HT4oyG+tCOX7eer1lp3nQw06dTv9dNSVViXkvb5u0GQvhHb2LijWNB6727d6MB
DcgTym0cm5a4Xzn2/KdNZTPcHUcc2rxK0PCAFWP6zT5DrcWi2bFioomGWBy4Z6mIS2yeXADL3l6U
hNVEA2QlBc/h/kC6+AIyBBK7gw8HzA1PFg0yPWBYadGmSvUpC3zw4L1p3BWqHxNzGyRr0n7laBXm
dVE700I9HZDWBcuu0KlIn5KARZeLwpd/W1HCiOBWpFcXEmQPg6KRWEUe4cuMoaJF1HGsEMkqV5OH
adYHv8e2c7ecYQ7V1BoFutwEL03K25AeN5mtmnJ1aKn6HOMV04OwwE6y8ClyUuHcKnYX3dPtrYg8
8P3ETGjWkjG3ap+KDfN9H1+FtQ+od06F7vIOKZwlXt79cCbPr1wgpxJc7umZ5/Eo8Vlv2lVqdZ7Y
4X6zrWxj4Wl4UKzILv2DmQQTCMBkoD/ZqBQAC04yu+buJcl83upqPleqfsB9aj/TkifPWo7xlees
y6WAszb+rM8MHKW2hZFqeq2sDh7XKqGLMD+V38A9bIsV/Pg0CZjQQxgh7Fc36Np3lijkakeuq0Wc
x4A252JlWsBGt87H/f2tdplCsBomc16Fe+vtwvykei1WPFnlF91sR+yUrZETGoZbJYDpsxpEztUy
3RSUMKMmtXgmjhAGnPcOMmEt16AM2b1/3c7sDXoIOhpmzmEJAoJ6F5YQWd9uj3+4m+IqiFAGw/Jf
CZ3wk5C2GcCPKjgMcu7bKnLqftv14IEjZmmHnbbHCYuduFlJHEyuRfo7TQsP/QTa1YNp0XUzd06l
U7WwBYHj2po+rhMkFPHaG/k6lcFeadiXMzhFFwicrCDZlg04EK+J3eTo1oWasGhr1ICSIiZaimEE
W/hcI9+C6ywBnO/LKa+I5dBNGgLQmhGPYnB5A1054+OW9CUGf5oyOjOK8bWM0NIX/HZwVjen1nZ6
xPPVCBii6nF0EDXMyi459s2ztXKbFCPPjP9AVFOySGcLFOspQUh7ra1mCR4XVFGnKGJVYFALHq66
JOQ9zWfOjIO81pXmWqByN1PPCIgu9DKHP5a0+Nr6sF61f1oIoacLasXuFRVeHaaHdDGjeMl9o70G
3xnNlR7iepK1Ias0pVBskwAaR5jhyBV0FWd2H1mX4kQTFfbdS+zOCEp1uwcKQm882PsFjXwcN7XG
gcdypLLcG6xyA4Fo2Au+HFgil1p/tgfOaM+9ef/x/pPHqbVwb8FTTBO3/HT5HcICLI2E2Yja5tBP
XzKyr8rjJmUCTUkWJwrwF9q6EpPxxBA05BVFQmSjcMdEGNo+u5OUJfBJo9LqCG37jg8tIVEoTfA8
ez/rMDoWFQY70m9YEbzENwucxCvaSc/2/ZRrmRMzRJEljGX/Uq0KM16G38y3L8EbIFfzVAcZOkkf
2mRncws10lW/6VF4QjX89Wv03yocJLymH7SR09xYH29t9V2i3lGsOsAdCs0FbPTvZGyugO2vFq8u
JT3DTX2yu0muiurOMy/7Wmzv0zSm/KnOKn0TWDvl9xlXx3eFAMzoD1jecuAnxbAkqk9D7ircIT8X
BSOC+cuDPsmTolopmByunf/PBUhWp+2b+Ld+eAR0Xz5AKThJuXiv/9MJ8N16sQuBPRPIrVheQZsG
p/cYAifDxDrEZZWFnrBaIsEATH4DF/s7LXEqbK75LN79l3d+BGsaUXKfbwEs9WQqcaSK7/hvo3R5
2KCBTh0dDm/QUNUFM3kFsU7JxCFazhY6QtGxl+rhxLz9GtPvtj+RlQ8qzseRVsrSzxhIIwHVXTfW
KP4t+otmcc+wWHIXgO0Hk8g283Pa3CTiVi4b8VC9nISA90iO1Q9vRydYLmMrUtevZ9n5B1wCus5f
ravrtGvUsLgRJDZQvv/kCOmZ2vYvMjw2zT8YOPCIW1RANn0EsedOknd5HmRMtFo+eCcEHwOYF0En
/KHZHcJC6jjco1VI85enta09iif4LwawQeV6am0m5gLQvXRWaiVpaVODnaZrjJDmew0c+wIdBaxy
/v7ndN6wGLQk3LPB8pSyLSNlJ5DIm3cAyHzx8MdSbZ7mXskMtvDizBAHUYAZh88apJWCxfyqLibV
PcvLg2edJuBTTumH2wYZthsoF4/lagjaVtjhcoKjGNcFvkKy5mP9IdCHWNtUCJs6x2Y8ime/36Vu
bmXFp2ZNDXi3emsNzQ3M1kPnopYaN44NjM9s6S4xeooVYvbdyTaKAUNrzdM5dskdjnmk/Bb/IiGB
qBupnoM10k1MMhQqLYX2k6AYUclCjVw6NOnTKW34V4seiitKeo0593Gm3j4D3nw/v0669FB88jof
SL1pLGwmkO3sKB3OYuUrOG6GxAILqaATDPOUJ8iulatnw+rQ/wzWcx4Bb6XxZhFyqUfzd9CrZUKq
o6pfRhOlW61BlsfQ6h/BzTU5wA9X45obXMA5U7VieWxChjuWnsQHzXRI4hzE2X0YES/Dz1rzmvJ5
++1TbcuMwdpL6cF11Lm12ztYuHlzCIrbJCksGYIrF46UKXxvBp103J8ySYW8Q9NeEXcFX8QaFvgz
YN8/aqBfNoQBG2LyiGoYvpbGZWlJSLQ8LJ+4e9fBDqCP+lleLNrc2RAykZjphHaAn9hXMnaeXA4M
gHTNXx623vDCr3+iwbM7IFWDusMZu3BfjCIi78c8zNkRn7DsAOnGVCfjAWOra2MUG65T5heMCkyQ
N5OW2KnhZvMXK26nY/itD4fUP5wJ2Nwyvip7w0E5A+t5l3o/TuQQ4cr1Z2Wj8YKaorwb4PULpw5N
u98c69dhvCEmNaOQjrsdI+4P0uzrXFbl/IKIFkzijTaBI1CHeVzrQ4Hg2W6B58fiPnQPlPiH+bWL
ZF7rOgK10nt0UXmjSLKlvZ/xKt3gdojD1YqDOw18gXNraEmwy0xHJjSWSEFHYjDS4VzZkbHSnKD/
CTxsooDusybejsaP9Jy95OLOry+0emLF6glr4F9UHoSAa8mYEZJ39le36/eqfH3lXzJzhnPsKHXC
M+e3Sa3n3glauWV8sBLDT0NxoMcnomwUn6VAFDzCFM38gNFQWislin24LA8mT5F0t7Efonl+t+Ie
i7I88JlTE7OZwmv4W8yfko74oFbjTnvZ8gJ+RRCVUZizbg6fHKuXDklVW0CC9vgiAWKZizSBKME4
yC3N1PaDG0eaVbte7+s8vy4/IrT6nnuec/+R7k4DzzawfqyaDy4dT7RlYT3FWitqUummqTd6PVHl
L0fWPYMtdxj3SoejC4QN7gLUb4ahXmlPmuMIAadZc0StzKOprtMQ8ybWFOyEAFJJjfNGOFlp49Va
VOBr59yMDHorRHX1LQQ+UzKIZCaGNTY229kx+kQ6Lk0ie8IJHkrEnEJBjMLfILSt24vfPxbjuB9g
KVrHcpH338Wpx9OV78WIpc0BX9+Gxadm9304LTb2jlDJ6xVk1We2TGiOj16AqyvuWUzXgffyty7Y
ca4u+CNiXDdVCT8OybB7x6vlzS2LKYTQURc6IBSzrStvlsG9c1TWd13sra1R+Z/E7rhRnR9+StLX
Qqttw2Cy6BDEws8UiHyLOQDbBxZqYZ9E67rk3LJxRMZojUjKQhyD5mUmm2iiKQeMaCcBL52cxlXa
kprCRTLuo843Fn35cMqoG/wshe4JoC9GI1zX9XIDBjXZluv221bnVdJlxpCJsGuV8Dq28dk4+3dp
9KoYuuGr1G4zKjj3jM0NYInKtvO9bZx+e6KRQ5m4zY/mBzfmFWuF/PjLpA9mDZzDwDHRu5h1/CGs
4P5Q3eAaA63P2Hk7ad3Jy88SRY7c47F81pE4GY6Qej8wii2gMTyDSv5z2fi7dXtH2Vs0oUxK4iJ7
iN8Dqe8RGUL8++DMzTv42uTwFPsUHkVRbgJhxMAkfjpTBpYYTsfZDAB8mVPsTQbnoyZu7QzIB6TM
ZkdBKWmnzYK7+0Jg3FFUml97YxD0KapyUBsK1dyJ9hl+MSu8g8TyOXB1KpSvd+qMucWFEH+vpbDb
D+cNcxi7UiuV9XXrMUt8xHnl53GCNgGu41w56Co0dVs99vEIZu6FC0QkMV+M4P0Zr88FFhZF447K
UYQcShd2XQ0Xq7TVwJ4YOK+b1g1Ui+Ixgyjt63i9MDb0WW50QvBCl206DVtZUPw/K0e83ZhVxthG
ZwlKOBZ9JC3XeAmYn/vdG910eMKrISGUYb6JXVurhIBvSF4v8Y3yBuQ1Rv0b4EtXkf/NmhYtcN8h
utxWKnTFmXRHlu5HulChD8sFV42A4LI2+LMOAd+pe7MAyYWXMcOU/shHODoxsewRyWAIbymy3KJo
9r709Q+NDAt9A1TW57bPHZcuHvzBz4sWvAa16wte20QgRy7jic9sig4yOcpMOu7q4A5rr3z3zesJ
TX2nqQHiE1Ghf7nLRrHMZXogOUwn7t8TSn2xF06euFMPrRmw05rbFpbDlMAGuwz+lkOLUbE8ujME
fVsj8fn6bZcEVix3I8gcf8m5zlUZT1/0IRWGTfaFk5OT+Lcds/LRcE6FnwtXfnrv2rgXqTVUhdIT
Btg+DkoR3WFjYB02uAZHNpVIn+LCnpxINrFX4P9O48brvDAHZ2FHPGZB5mkyJteckZJHzHnl5gPr
SCxKVKLEoj5dgN9zjaiIDoou1bU5tBg1sRaQ5X/4uciCE1m46dYaM9U2kQL/VZ6F3tcAQ33hnFif
iH33kun9s8LcCb3AfKuHQOjTG2JkOPUTR35cczTFDJuGF7YMEIoxGNOgpUPVeIUyqYL94PIg0Wd1
bF0c4ixMyUvl3J0dSjRUqGHgubzieUXdzpkP9Oc23G0z9gVbOjEPYcrxdww8OWpyMlgenJcTZgNq
Lr8Oq3Jy652fyWnyO7GGb9KzdkzAG1eAwrs3/UPaqsZaYaf9qRI1Hc0WQNSEgRwMMed/V3De1qDa
Jcjod6ITiLCefDJlnldvzFluJiJ3sa+c57HnwYMprmkYHKj5rHybCob1qxgMmASyxam+O2kLYKCy
lTKH/5flQh+zPHe5jhSaO2RfBsMFfpb/W5IB9B2/I/I4TBxzAbZcz6PD51bQ1de/iiBld/MdSbc6
0Iuyv7eZ7y1yq4pWez8HR9G7/sGx8ZXWfgRc28RmySldD9uspMKS1wNz7Y9ibbyJLSlE7f1iRexD
AULwpOsm7Q0Af0WLZyx03m0MEvAcMN8cuYihFK3qnY2G4CjaRQv2KayhRp0XF44/JPexJFzmclTc
Nn8QBD/R2AE4AN/pqmYlo8xDmzWBFTkhMrtc7Yb46XhKRyUoi6TxoM3EsbDHdtPPlMZd1tsEpj25
4d9DK80KB3fXxTezomTr40rTp5rqlNNiyArnaWmztE0fTMGw4LZzP3tktILR928KcWZw6DAFkl7t
igv16A6t9g4/fPnqh7Vuv9fxi2wJv1gEltxtGriwK400M+Xkql54B3095osjwlB0es4Fgtw2ze+D
zKb86xUOIpn8BgdeU1+rrzdMwDc1ZL005y3ramyFXcfUzHKqYIS2lNJexdhZVwDh8lbK4yxRK52z
qrFFyHxKKr1DBXbdS4KOIw+H/H1oq6gwQuxoj8gOwR2otkaOrbr0y6dYB4tjmtJTr80BiuplarIR
O45PQ7g4YW41vyln0G/QP7bmptpSASUPeCPMM76C2IP/f4f6WI6t1fMM/ZM4zrW7cuIf3n7cMVcl
VSeJm/SN8LQK9p1TIpNRvfTKZSspqIxH7MObBgiy6iN5m94VQJiCw5gXYE8I9mcVsKsdd7SIogGT
ccx90/9k0UUaqBHObNBo0IVF6H1fsZ1kYk4LhM07LL2Eg6/PJ4sAVcRUjIQJFUX1LOkx4/QHoouf
uBgjc2bNOXLUTRBtvuzBhJ9LgnjIcJFzdxvgByIHf7HLZ+WSNhfk2nLGzXXXiC/wAjIZ7jnC3Gfq
RzMcc1NnsKvgBcPqZA7HSbVxB9KJVi97mOU979XLpJYr79Hd1WAU3rFy9jUsSMg76YuLkT4J+iU+
r0iYmgh94GpyMC/NDBVuNkMFbcmSgIXOOXzicgsu3MXKLq7SXRYMX3yiggFPEu55bYCJMYXS4NDv
TeibzO/2jovclZT2Qz6toRLIg4gKSxY59cM24mRTAFCSExah3q4waA9g+FNJkvuYJHp/jqhAOdq8
GqHdWO1dRYqs1QG3VJudZwpKwW5PVONeXlPMzKJX2PfydUWFq5DPystUM0v/20BjHStXLpZF0C4a
SSBO/in1tRuzSEO2/M2oODTYJBW2gOi6A1RcMaPvaaRNwLN5JjXvoQ7kV84Ci22LbzK67Z5kQahT
qDGcBOu77eQA9YyEQKBEIYFoN8t51yzqo8d7lCA1S+3RbqkVt67A7CtiZf/diubqjqj6XqwZV+Bo
EeKZVgfy4B+WDrDyPs4g2n+WMBxfqZDadtH6Yx9bmWAh/uzDDNJmK4wKF4RMxJ569fl5EdBSzYTA
v/+NmAfonJU5Z4ZA7beCo2EBzbyitEJFAQ3bsr4qKHOVe0KHqDhmMIN6Iab9BuxGzenTI/Gfv1JG
umxl6KFayq4IpMFHd1WTOa2OZturoPKlF7IGGz0mMy/KgRw7FRDE1UhFbh4eT/f7Egf+HwIWUzty
a8pziwsusHF8oVSoeqQmVVdT6TH45beUCOSxTp4P0I+alhdTsyWu5sHD73bDYUEwlgLRr1r/QqlF
GTUP4smwVABlQMhyR6DO33CLh0kaBdh7VxnRBpLFcXzvr2Uluo0qNkY14lQxo63F9BXGIugnN648
qxYh6Fc9XZYdgTo7nAbtabrdmlKgeRkGdRe5dfx8SJKWs3FBBcbjNIlGSSxxY6gRzx/1TRE4oD9Z
zEDzSE0u6hOuYCQ7ijFuzJnq7GF8dN5ldN9hOjNY+I91N4oQ8uSSzknmyNKfBxNCC6CiQ2YArkw3
1ODVJuzYWT6xJnXHNweY17DIvDibE33ZybZLky2MI/ceJnup7bThrRvVMEFJQ88OvEZF5UQYXxXP
kgTY91S8Q5NJCMw2zOSG8H0fHTjUMSHY5pOvO+kMfAL9myFYEog1jWqRG47UTMcvEd5Z/bfJfjyd
mP6wpzfEmGOM2D0WLmKFvsOIGoTm8wV0GypAPjuX9Wxo/l49WQ3dkcHtcsk6QAZTLi3NQ22Z7P4R
KttwtsFj3or1w7A85ex2kQ0jUaxrmsvL9AEzdJf5TPUs4Xyv2THGxbtCj8Q4J6jNjECjaWt5l57o
bjmt0V6xOSFhLfAZSDJ1l+1swSMU+boQ7BHJuf7vbcbZB1upA9JN1lLAq+xsWwUjbpIBY77NsC1V
sK4dJ/jljXZyagEnKLpIpX6WeJ1fj25dl+RQsRZ+kUkZJ2oJxI6pLtWKszLnVhhzz8TY0O8yfZIZ
t5debasBEU4yFymCEPTjDNx2lzVZWZTr51H/2+Z21hKM1qCGwZh+KmEvmEXvY0e5y5CH1GrjRkGc
b1EA8vZokFBkR+MpRD7KoWMfnmzbRGvMgtM1ctLjwugE89wEr5v6+Ooyq9kVkwSp+nPucIAiDqjv
F1QozHqX3LsCn336htgEJZd4F5WpiAl8SeY7MOF5OukgFxcHTTuHHktWpUXfRFEHPuDTQJkVWDaw
oaejvC0X3FRXCm1UMUsaAZbDi7NforRF8upI3TrCYWa+V1oXU7qRTFmOxuClg9eoSAwZdx3fhY7A
/3WFLl0cOlm0otJ4xKhI7G22y2l8Wc39CGAkNzUBtOcFXt0Cb8uXXXOlmySJJD441vrTCs/9rq7t
voMbdT8KZsSUR0WWhNWpnx8SnODdX38yLxPlqC0p1cWnh06SBXDUD9uQy2XQGO0dep2dmXjM1kjW
hhMZCkjLBKL9+ehH8+dpI/yr5NXHaCmPV/ngbcqoQiFguJiqGAmXR01RpSKyArc8bLVeFJq76Tsv
flh7Gq1P8uxYMzVoprTver42IFKOMIDLDzus7h1iHAm6eF/L+Vg80dmsHg9XQErD5VwwZmUoWtrN
EDjQnNV9i1voZSbKbtaPsxIuAAA/BtFGtCHbMQ6dhsiyn06EW9MYrniDMwDmuXi5TLEd/Ff9OeUt
u3kIk7TwWrjoZT6/rMFjBZD0+vHjB9M/IrjgKorL+Ow/vtt8N8ru+VvwzCbt4Vs83G1OPMv8Gbny
RM6yypOM0BVCBqIQ+747bXg9OdYC9ruSPmhVUf2kYc4XjhaOHgi77k1K+rIhQwjVvHgquCVuTE3l
pe7Cw5tWNqsA5Xyi1vApPyMujUSLmF/z+TM2j4cmrJT/nCxJ8Foq+RJoYYIGKYZKiFPM08lHebNT
7b8U2wXpBP2tyAw9aGKhnLljgkQdsag4Q7fVacGn3NpfOYVYhp0rLSIkmNaMVxDPo5HIM0NG2ij+
6pEKeVjY8VNlJTzS2Z0PvXzl4usrg1Fidz6ryRILxbz3W1aI/1XLktb4v/+Q81Mv64JRxZ6qRo58
j1kKV9lBOB9ocxkQJD4whJkhLAhiRuh7ZyMPvW78rqUw4tx2j8fr1Fe51GQkGZ9bneMHf2Jnt5Tj
HwxARrv7ordzvdEiL1dLMKFwBjIZ/SOoUdqvpuvByg7VabZoWt1QV7Kv5jf1Br3SAYPlfLN9fly7
LLQrU6SoKTfq3vpQoiPUoD/B/7uUrZLvGBZ5AsLalocDjA52NAeYYB+mJkiujsyLoO1LkS5sErCk
6Bc5oqguBxvtURnsVqAcWWmqZmMmGH0Y5ZLTlYTCsGZbt8tbBcGAdjqQYbbyFHO3AB6pkniFKMGq
E7nqK15pTLbYMisOSbXpLi1ymqr0OnkQEurk5MNBZns8sXP5ZCa+Vehzz1Qjc371/kStIEdFtxvQ
oLhmINeaCTUIz43mVT6V3F9qMJFpxhctyJMO3Ng4QXuDWylfNPV6DD4ZREtjc7aeBi0apUrUzcTT
/+ghLixP2DXWQKOuUjGHz3Llhpt2OLWVx8hIJXHpAIkKnV2fPuxb3ja1Rk9ufhYPZXztk9imqHQw
cTWB/Az8iozT2s1nxccU/CroiDTkPYTYXqnS7TwMf485dHdxndHq1SsgyX3KRdpeUqydUNqQTeOp
IHFYn9YDnGz3Q+2AAw89pQaTIPKSaEgGemlogyD+uvuwXFc2jYE74HzUokebs/EgXTNaojQQNoBZ
iPyj1IpoyZOiAzmSNksM9oHM1kGwohIc2bCR/LJfBOQDYdschT+0QrIyrIZbIw94u9by457rwYgX
ED4kBvN7nCbT4cfEGojiS2jadFnDPL5AEcoatm+8ccw2u/iaVkYY6jgrr4LsCHeICpbqie3729Wk
5P6+gsPbjM7UIOV+hfWChM66jfQpBIRkyjwPRV79EInpjmlOfEumpYeQO3Y6PDjLI0PfmwGYHACW
lqiQOGXlGV5+5MGC8q7Hkk6HrP88qZhqeyg5kZ+7wsrukliL+v3tToa8+eN17f7UP5bmo24283Jm
kY4nkZc+k7dMf/H97oA5l+i4FrKZPUzCU4DiK6yDUHz6m3dIlxjhIgBXKhnWiwbiJ0ZusKS++tp7
Dbs47SdREjc4DAeFQaX4MFGRdF/x6R1tiui8I1Nap5H3s52ab2bCGz0uwSGPRQZzQljcz3jBSflC
S5nA3cHq+SxZkb9Yz8cvsQSehGCd9S2D2bFCYpe+zOM4Ma0oHcCnxmhJweDoWDwX//ilrU3Pax8i
YRWKknlmwuwOl40/x5MQ4Jo9hfSeumUcCfegDfFBPoSShKiSg6WxJSFjT5R5kSq1YitdKv0vyKw/
FTPNwUFBL17QWK85Lvv2pp976zCAZq14A76ZcLrVh4cAg6fJuTPc3tqTMYOoub5a2sXyjJJ1jaFR
ruwWR/HYa/emR17k7lFczj89TK7iVhSs2iPmEV1XZKWQNVjxiDnj8Uxw6YjfGRLrLQxabz5KgEU1
Q2mT7A5WI7ps8bq338p2FF4R+7hjx/6uRDksqB4trAvdv8IV8+ZlV16LwedERgwUqTNbUz0IB2h7
Ajc1J6iP6I/XlyKpDkhCyJgdxN3aselcit5ga0QaWqK/+tmqkmWQM6edHbUyZ8Lxn/TNrvrwA98n
dOOG65/1wjZ//BcHPrsr8JejVAF/gMknKim6CfIecoH/weVHDXVDzzOvYBl7aGh8UZtLzU0ORus8
c63ekCDTerCei/pSTrg8MUu8fXtizptMw8vszMTkOBp0F2Is9VWJ7c0cvXIrlryA5zjIqtGJSanS
rdKUa/JJfR54BIFBTfz3qqSQEiayDlG6j9jzrSMMPtaFrxT3UfvNYDy0OCNzAvdxwSB0WT8STAAa
RhyoLC/2fHPxFKpP2ChkhAUIjzhGbpym+kCZ5HKF6CLD6L5GGyrhsbTJA5UAKtQQBfe5bnspl9Pu
CxQ2g48J0vRymk3MViAHYgHhZ4zrPYQNeflp7VRE6UIhK0AxcoB69oEj13HHmgIYJ7b9dsVqX2rh
+QodN/G5IDG5L4LrKN55X+3V9karpfL3wFwxjTdDZ0jCgt3NWVwJfJDXwkVQiE16MGvEfwGm2ODc
0kwsvfArb2KFj2125iIF2fvRU8uLkDOs03D4XbNWGIqKLSTP0yeudkN4Vjro98dPgh7XuQ3Jebef
CkdvOnjElWDOIXZPH7rEaPrjJ41qe4MQvQ5inwPwb0Rb8AW6sQjZ+ePRrOaBNnl++CJd0fpTqDMU
ESqN+SBv0ZfvwfcTrqt2rn/OCl777pWDXS3dcNEOoBeexMRTPZAzkCem95pkpZru6KEDuhrYmovH
6Qe2d9492LW0j9RkQFJm/lbiRI26S3/9KJkJN7X6C/3NCtjWDEkz2JFs9FV4f5c0XpF4WfJQ+dYV
SXGaHPjRcUj/HGGGo3sXQmVyjs/lYiR1HT5Ivdm5dhWudk2pcUJzaWiJ3nMZ0fpiAhW+eiT2cV5B
taUyqa3QDdA9L4IcCff7gbCNivl4dicKJo5pKL1yqrUorLL5t+DfW7tjFL8m7TGMTCyxkSl57TTt
OKydr8o7yDPfDVTx6Wv5L1XKII8Fmfp1lYN1hVdtDbTYALexlnTEsW4QFzHs3BApudnhXvzB5mhK
aBWQ1YGtkRSfUads+Mk3DkXfo8bYQqLCAQHVr4ku3DBg1eapP/5jlJjpN1oalK0iTswBmPONdCKO
8mqVV4FlNh20xyq8pey6h5/8OHZhrZ4bceZG/wgGN/qoNhrdFRcMdo/Hkp7735RnMfMCxTYj4Bml
+ucoqa82IxZGZdfpyTPQYtxG9MGm02fs9+jwcRU9TOfI8CnRWXNhVNbesQcHrAPKJqWtY7NZJVOi
0Yo9tuSMYVIblapAhIthdDnsaEUoLOnb7eziPK14VFI/HlM3sMCKzb6fkMCKl/KOA9zwRVuaN0IS
yqZsV4uslKu69cKTFQIWP+3Dph4cZXVe6Uxv7OqAB9WYTRE1UJ2aMhZ61AbbqSknldCCXBZoGiAW
Ym0oMb09DQUIvrToLhQKBiws9xsJXsHKXAmyS1lV82SfrYKCOLy9KqqAhss2Pgvx9POz/GW/figO
J6NlvH0Ls3CLHx/rVqqEL5/dOYnFf5/v+D0REAENFz4fzDQG8eqsmShxgxdK4Riyr7S19vaT2vWa
/oC5NhqnAdAhAsR3oDNRdlpLrmTNQZrKQ8K1zcFdWB8Qv8+Xc9+wlBcrP2HlNeZdxJA50LQdyBTY
1AzX2yoMBNZrmCuHpuCeHSq9Zd/mVVo+63r7YRKoHDQxN8b6Y7EJT0fTNZzqOLjyXcBaRqlkcliP
QaRB0VvREM9WX43/3QpBov2bH/nCaT2Lf6ixoP4DLyIdZaHNPJEw8dfzJLjwmOE7UAbPe1SLkX+M
KD8qsmI78kL/y7lMe30ndwBUAvBpq/MyMGjpBUZSPTta6g4PMS6qLloVzU6aXNT8VubnBl50N2/T
5DCFJs3lYfYFRfqaXTD9GoXVeIHDgyRpEU+JOC1YWRNvEDd2kaTrovXSRm/V9xVvX2mhhQ2oC6GP
uJFYXhLu/w5IiUqIK6s4gUP171z558HFIBA40ABYD+yOyvFZdopaTcXI0HqYEKV6MvkRfH9v/5wc
TQeEg9fKS4EF15YY1/nMHPfrAyAlhirWg/0ujenhpLu7yx1PVd8fR+QrmCV74y1844McIdxrnXqd
SrDZAJZhi7d4X8UJL+LAeuVCwFUTo5ZTMNFd1BovNx8H0kEGSBXcli6RhHGu5To9pD5a+4eGxQRb
ZVevo6M2nTx3TZBkJoOg+i/uQiD3wNK8rJsasovRZArJ4WOekX98cBUpa1AWDV2GL77tAPzBrV6y
f5FS8femg2S2dd/Pv6t/p/KT0PD9WBmqwKs6MxAydbHLQicppe7drAS3upaUFSUKyott0NbJSFEQ
pm6fWwoFJ9TDF4tP7FB3EF+DR56h2WBOJ1BO6ZbWo17fbYnCQuMDA/pU3mR7/J9b+R+Z+1Vo0X8E
8wK5/KT0Dyntg47vvtcDPAk8VO2u3FsXvUFwqoYuuwTZH0Su7Xn18STTq0RnQP+JvrMVmbrroHyd
FkDuK+thHox9Rseg6fzyJcPdZDZBcxlObEEAu1Mw5MX5lszqMQDfmfWAqnlecvvXsnXS5R0E5zAH
4GbHrDwIa3pr7P2Tt27Ben9sTQTjftZxyLl4j5h3YNhKDQL7IiDs+ijCnH891vyrxLxTkOxIGAlh
pfZv74pLiKXKAHpqZ0hcOn813tnnxoJBVSq/aMQx9swaDhmOsojHVY9KKkcIWVpq7szmlt2qAn5o
klXtxvhxWcmG14KGCnc6UA0kWtsJA2+aMfRrO2Cm8Qjy4YsgJbK5GrEphB9O+RKqifdSsiS7pe7i
GEto7VNy9qOEa6i/jlcJQ6jO173NOE5bDDeL8PCqEr2pVlrnzDhuHCpWjqwixX0BcytTDBxS5G8z
LxQeY5hAk9WG6Rb1XD/wb/m2wDH6bK5vlOpQBkvyaDcdT4KdR7VmCs5AaWEZvGAgTunVwi8e+ax4
FjUzNjXCt6JV+i9QTczsWFtxictNN4L6H6ON05S+R4eNys9O9uNQ52p7RvQUsgRJFmqGbgFvaOki
mNQYdZZMbalFEX19yj0KyWy79B1ZE0HTY8Ki7BUihILyC2SDC6PgtHXNrOxVFAJZgzmwcdCzSKu1
O0tQQrrCxplUhMtHh/GRswYr7tRzuvx4pvg3Z7fVoj0tB166hb2WHMlWQCyZN6jUq6ai7d3RRtR4
Rlmf4E2iHb7gmd3ByUeCPGQLjGOv5CH7V9bRL9tnGnx0EqGw3iJRi2Gz9ggqDS81HrFLmJJwoD9S
ooqtm1HG4VjiOfwe8R/Slr9vvGlrfp3EwUUUGn1ueJ2UDc1eBCmzYjbrwCsuUyFPqTyO6q53QZ7i
BNOxrkxxn6R7bzaifeDfUKyWTZNM1sIroe1hXzh0xP3XeAqLttoFKwEnoCRgl2+VsTbJXma/s8JO
qhrtEcIViHL+2jqO0zrzeH59VHxnhyApu5GNamuxWJNmRPWBuxbI2sPb3SFhT5qW17sxhLSNt/8m
fIpntEPt0GcCk2V6ZyCs+oAUYt7d6PPbpDy8wWe7VsNTzG/Y/2REC6nFhoMXphwq9c+gr10SJ5WL
09AQfDGwGcNvo9UODmQoJst353yurxfvsUNvnI/I0LjlCX3RO+W8aMCxCKmyvg5Xbzu1l6zic+UM
N5CHZ5us1/CqX42fpyceYbKdPhmpqA8Y8gJVonxvYqOqZVhAAwXiVEB12XQh0HdgOUDQYLABjZFy
58dOxyPl8YieEjYGulj5fuRlkRTK0xNE7g26rMnCbXai3i38qKDu6zmqaT4axTRYnn238oKfoi2S
na3Pg7OSS8dOxHdzavSMj/s98mRHQeDN6JVc0C//Bm7fn6pwKfNXaBr2cowJ7/VaZFIQuA82T1/d
+f7ep1v2fxQjtMqPO0rYidrF/YQUK2jFW3nsWkva/Gpsbuw+YBpYjDmUkS/a9ne6z7rsqaws0dZj
lUTMH7JNd0TsmtL87Pauu3DR5kGh9nDv8sohSOtFk77haxTX2uA7Y+FmYuAqM/49HKUtQ4Aa2mE4
IZAic2TPZVkE1g2ftOr09go4Fb5yBMBftKTEQVUo67FUNcmZJfdVntUB+TkNyhFNIw/Nw53ZjzYu
iCDt+KD7mKQtMuvaKn3JtTzdiT6ZM/SIcjaP8D0TqiBQjZM7s9Hf43ysVslaMkvZTkUikkuX9oRT
0mG/gOYVYoPXWkcgVUeXax3Ecb17FLhhflVDDGRNhtfxAZbimOtsCAQ4m4L0S39ICnsYFzGUqr5V
tXUlPmN4B5jZtoP0ntjA2H64B16hP070nzvhMQiywzlc8NjHLIvRjPmRsUt6xdL8ina7zoGWwlOe
YHeqrok5Y9tLHlnaqdGuATRwJfiCu3oQSJYVDhmsuOxxUt4fnGPhySFYx17vhEB9KVxd7518H9pl
qQOCFhJhpdQ725k5tyqyUefsJ701uuZEeXwCAXtzQa97h4Qem0f5vYC1EFN6+JgLHdx40o0X8ClI
hNy1TZiyHEQZkT/kV40zKCgKLhSYI/wvVftOzLG1tBsXDgdPHofjJQvvhdFxEcKQGtHOeCrSbpsZ
m6MVGS9rJHyOK3vXid/TArDZuTTSQ4nRsPQ/nbfROn75+KVaDsYyIOeEMLljrrcgdMlva6PYd3sE
1ZGFLjBOoyp/Nm8Ru3tigIfwyYjSikvRkt8IN3PpW/oq4hlRadvvs2EVRWxPV1PIKtRSubS7CjvF
teLsseDJwEQ5HlLePYwWw0r0Gq6CMKPpM1/k2WJsve7A5+4c80XmmxDCEqRD1T0Rz4lg8oFLJJxM
BGENgYQh8u0Bx69ai0OqIfh8TtC4luhwBRIvkTjwkvVhubYOOtsV4LnMsWSq1zhZwuxgjWj7bzSy
PY4TwS77J0YfKPWGtzfzOOMJwuwH5HP+HWJcvqT6PRxmYS7yKefWzZLt9GSj9R7nZfctdY/lL6vb
NuCfqXQQ3ejKMufoYkOCbrF05zOib1Vc+4cKRkpajUHPzzPUbVmAY6yl1Q4baf1cfwlRKdfNum8S
5d38Aqhhc411pK/w+4eja92vpqF3Ngl519f4RMHXlL1aD3Ug21eUYwKpFm9iIRf5RU9MbdCLMBgh
bB2qKRPVT2mqubIJn8rWm8uPitmn/9rIaMSKz0V9N+2TjvT4o3vhIf63xsgz47wviky0JPpDG+4X
N0uy7JG3Z1/yOtW6OgJbKVjE8ojosGDS4Bn/ZwuYRSbq0SuH2tPq98ZMpJ7BY9kf8myZ2aM9akbs
L3pmKBjsV6CqgTmy7ixKyejBb13CtLXigOcFogg3vntONdcXKnKXQlpcP+d2ScTMuFnloIEibwP8
5PTih1U17Gv6RXpxU5KNkBogRGQvouucla3SXTv5z/A21HnQz52LCqZ+oDr/eO8GT7ezHCmjf69Y
j/0coJ6rMDuRxGTTwjfrsoWYG2MpiaEj9MnqlKnF9ZZSB9KSXio37F34bfYgxiHfPvzpGGnOcvXh
T/s9X//0M8TFUz5B8R9PLLDJc/DgAZZZigm2QnEE5FIyd9gSt4BqQ7uFcZeppgqj8hnDm8r7mtDl
oFxigbrUFlfat8Rj0G77rMdftSXoqBK1d91AHxO8g2KSxi3W9bQJ57FsoWLkMocmOm0kXM3qY/Q5
uUbH7JyVRKxXhkxDWBIBXave4libBE3sNXewF5Ve9wDw37G7Po9cHzHHw9AY8Dom+nJp7wLGq7AA
rt+n4kbuGhd+kbjHbiPvW9i/kxNtbJE8Faqw2Sxs7mlVDVqR10Zio2m8PYDlvXZu7YlcGrcc1/jQ
kfL5cNlFCXhNtJ87txY7EffMhyrxrJaOo04E/8sQtJVY8ERzXaOyWrNZlZFyYCsO5nzr8KtqpY6r
9qbFNukbsCSVstFFO7btPWLRb784J6cuJguBI78kEj2WHKhh98gwNdX7JzZxi9hWAmyg49oRnH1F
qTeRIQs8P9I29S1t/dHAG9ih/DudhZ3Di9O5esFBZ69olT+vDFo8iEXxhLOg2irE5AhT3Aidl6Wg
lDiLBrDb+/PXmXnaAfup7dkfWgDhRwzBpsy8X1yfwVMKt7glXvZRb/JxPCrnd/Xs3gU5DxC3cRcH
711kHxZcLGxuHj4/PXFTendlBrBLmUBLpMaJ1GdaAodXFm7z2xCNN+eeFpRBNdad0b1mC2QkZO4o
krpppN5AgXC+G5F3GxbCBhvH9IhsZC42OeYYogwn/4Kz9hInnrDA+zuk4tStOqz9kvptqTiusJqk
gCw/xjgUgY3+vvCq3ON7/MdKDKwgsJJ4tMo+eyXiVpLCpVnjE6Vh+f016BGrxbDndqqHBjEa/EDf
aRF8zFytw6Zmo7Iaakb7sD8gWIbYOCFknL75tdQTDD3O+zHaFAARw+HqE0RoZGUuIuqf+BjptTA6
ogu/ar9xODTVbv2yqhonh9N40UD+3pW1IvSx4VSoY/Muj/5Exu0d5WtcquYB85bUJOb2+NIQpjQS
i/IUG/6eFPFvKOQUCMjuxjAiVEu5ImK8tdCzWnv5FMLZU9YQkpEjjGnAj5Z++g3MNUFRKGI29sVm
9LQYjnwxhu+MIiwMcJgo1lPiDHbJdSVq8b//LGkpbQXAvbsyqqqHDrWNtzRIksl8yOJXnkBkNoBS
Oc/NzEypLmEKOY7VlhVm8vVxTYCcJqX2Jrp6iJ+D3vfIJYgUcQeMUxFNai1NXiAdCijKLo7bdV+L
2uRuWV8bXgr00cPMjthTs7w3KUQO24if2IyEP2csF3vScImK/1w+qAb3hxSYL46kuZTMN4VLWOrQ
7wjGHCBjlTABGFTDanV7aqOmqtiSQFr6g09uLhNKwMz1x8oSweDeby0VeFr8IRKLg6zFP+HGqovz
vcBs+67fcu+aCx6RuPtWjqzA1McNm+38MmHAXpXNzcAhNqvLSC1sCMDod4JkBRAUshvAIx+BbSf/
+cJ7KAf0ffPOMRt7/Q43bagirNxrXVQubPzuV154CtxwA0DzuvUIva5nf3OLCqHAs87ZjBHU2LDk
PXW+O9GrNMoDdm+EzN+PAyf1H8Mc+nhtDYcRbA4MjafJvgJFUTSbCybCJuHk/reMBkOZOuyW9TNP
CvzmHWjjC0DQIA6x3iIOo58nTeqiKJ35A80uJaesGHGclb+zlGuBAfMg0wdHIhricCnEmJvBi2zv
ES6o1ovJBbLDfjbUzsTCBqGktau3Sy9n0Qc8U5gdbOQtMWpfMQxhAhlKqC+rObRoRN7u1eX++USD
9BCSRSGyUnxM0SnyOQn+V5M9RoHZJP2a0M9E0zDkKZayMBQdZ7nYOlRAelx9HZrXV6oWrVrYdS5H
J5v1jFRPyp6ReVMmH8VwHpEHg0pwpBGeDceClpLk5xkhs24FBP0U9uQ0dUQUIug7iHZTvZXdklHM
/cRCEzvkeywPWSUMR4ijmax7PEkxGXJ/7Q4QLDhExutrdZ0aNYxbSJ96qPbz0PAo0I8npHRb3uSI
q9C4w6pa5Be2eSEf9XRs7utOXE6+8QyZwrz+Y3u1Ln6xgm4U1EBQ4hLSBPkNOh5ztamcRunhiOsM
rVL3NrXP354LaZkIvE0sh+0ki3DOSKFmCVwxc5OcvQt4bOmcKUWPCitWRr9Fk8KxkcJvxpLj8Be6
I7cb41lmFGF+zPOs3V3CdpZPRdjVhRM9D3xInmqiJe1A8348wca3edslZoW+I4Kp3sQb9F5iqTG0
M33XLfkSeh22XZtquKTwk1XjP0ZXJDYDcyBxMwnzBicNcOSlpmkb5EJctD1inwCa6zn8Hhss4UIR
oWzibvHQTEeD1DnAhxV7WT3ZHa2LLc72H8hFC8kftmZPKvYBm8QZBYoVrMHQZuua1PmLfWZkz+Vq
vqupCg9N3/ue5pNBI9X7vAPbucnNOLVVFnVnQFa/KCLA9D1pQpfbzNUlx6WKXJnJM+e7UEJ390f6
Wzc0SKxy/Z1dfv59JwKYIdCTv0EuszxWYD0wnslM9Vt+ZNlaEK5hTDXeOfDPlJ1g/6H5vF4k4TKP
+OSZTqGV8ykR5aIGeBtTA2c585TMcadYTohB0geITLEt5CZ3FfN6txsO6rD5+lZuyk8dTiV4bqTI
mm44Y8TI2XohD4gLzdBGbwBuL6q7bDBxVTVvmz4+ewGowFPT/7ZdwYcgrtek63Q27wp5CcLhH42g
792kX+aMFoql/QrhfB7UMZbimaKYHR3NG0Jz+zAwWlDqcuRBFwLVqg8FAgktoD9Y6riDPigSX/F2
9+9ibXzuOgIZnYAlKl7cJ1PC3uQitYtrb5e3t78hxdGWKSwUrW2JzsDxgmlgxwih8n5RCEBPKxsG
SkZHtb6t1VYYu0EkyVVC2P3hK/cmkLYeunNrDR0yRE2RsbTuwzncrYueoyq5AXMaVmhCgK13Boaw
/pU/WRQWn69TdzsKhheR+d/cjf8p5uD0Xt/cauxdzlhdP0vFdnly9Db0+PtK7TfOhzw0bEHgc82D
ekz2vbcRx5Or+Gp503ZVv7qmHWGS2T0+5lIM/J4Q7XW4dOVoYOm2CwZd67iKm0AywRaGfAX2sI1N
alQYkJ1mpG/KAL/4zmHe24iC2OFT85yLHa0CDZpIp2rX2kluWTzQmzygddvATIHplhWjTmHH3D1n
01pOgGlZdxH4iBe+c0v9jnNHBl1FAHxs/aqB6+DNIof7HyDgIbV6+a9f13l3KYr11rXYqgzawnWb
SvA7HQcLj/3SoYlcafU+cZgSldNpGN6Z7HnTaTwC64+qhM7+MQ+VCcjF2wCHluKxv7PxWwY4TrOs
AqwpZXy6xjegal2RgigtZozU1NCN3bydny5j4Yt6/ma1CgH/d1HW7OaNraJSDu/xDg8YtmAek4S+
2aFi6qu2CMUUBpYq+hg8OS1ZAJhhqGiZ/m+YByr+RKX3Zom1tfkmIxCow6AsikyMK2h8X1nX9AkJ
ZmtpJHYlM4gR5zx9pKmFv4qAzPVpMkqK4OXYJyEIlO7PuDMsfvsFf/uUil6mDg+TO3K/85OAfEHm
FuhGX76xEJElhvn7sFVf2YWPZLNkZhTxwSwnvo1bn9PgbpkT1eSSWHDHWe5luwFtOJu32FXoJjQW
qj7FL1q0EwAk1DTU45ff70UFfrgOioRuTaWnhWxvXtZ9td/fgbumi/V1+IqAvLpRjm2OrN38FzEe
SQRsmFQhlvavF7/Tbsd+YagAo3ibBZnG5q4gjH6AvAu00P2OK+wJ56KS8VCpQmGR0LIRJXOsBCgK
7zTrFWXgWN6AW1Deki5kxw1Cgvtu7LYQHQ19TJfsVg6eWdLY3TUVkMrlkXDLk1oG6ki3JzPJdxgJ
31XVk355jttEueEppBD8FXdIV0MFeABfmLIk7Tb5obgEAIKEgZwWUAYzYjKlvSjKlN1s65jyMH3a
XPYer2/v6++V69PnRYJkYKfmLPy7IqZuP6wAZrPUzaOZIj1Se6MdA68gxp/e1nM3DrkJ+JYt6NFE
RW7kmOBT1M7aOdOLvA4abHFJs0IBDbmhdcbmgZp8IQAMh0gOo3v2kC4sMya5p7cENagxytPNoFX3
k6CwpRyvdKxKPd1Yc53YRJ40QGY3MEJzyFjOUrRgUWjPTn1kU2p+AJpf9vNagmTgfeoouMpm99iv
pD2/PM4BQU0ngkpCmUJb6I9ffiusf8NgIS1wViIfMbc0VAk2ybba24gjlQhXoKzsPeMxvaMXUWh3
eD0lgrS5lsmmrNTeJqqgiflrB9pVIgTDqrWNTV31C7IaUrtaoo7uLe7s0GCO/HNn9EDajcMzfj8y
Xxf1TPV39m7QC+0XpefkNg+OJbt9/2okBUt+LBTbuBv+6VdmbEwd88Jf0BsJYIz5zaXkstuIW64U
0pCDpGk52aAathkFVydye4v7gdTJo0ftj78A7gYIeDMGE6AbNlcoZIqpkBQmIc31Mkpmk3eIXpMe
yvsXpk5mmZr8YrihILP7veuA7ceEwz3ZH/ScEIfiMTYHwSHE2l3jDlPmf/lzV14s4hukzjjarEYm
dge+6oZhTSxkv0MjOWQ72x8ayBIv4d3XQG5on3H0eI+MPrOBBwDd9rX9HYG9X9c3X9eOTAhyPdBo
KmS/61VjQDaI87oliwWX0vUQmEQqv2/MuVfb7yeUbEnX9STeM/PovW5DSw1BECA2jNxKBvjjgtWq
Fl5DPExAcO7ofo0ZUdNFy+1OK0w8Tx3CZIjIXUPdL1pYKJNCNN0IVxDGKF8PfZnP4Ptzrhi4FX6s
xSmG2E2Q+3POw+N7E7xjUbTIiZ4GFv6bcadfnRjMO1py+zf+cYjsF4nhHGhzfNPHW9inJnVt+i+G
fepkH3ySjKYLhb0Gw1CT2LTjI4cj68LAElpEeSCg5qmeLGlHn2QgE1kFmT3o//SE1SUIi5abYSsL
R/UW6OaaAkLLe97kKrKoEF6wa8bF5PHxV7oV6qbugbFYna9Lkvg548S00SlzGxMOnLB/i+lF5b1C
1agMTBg6wR13yOrn3Y/nCNHz+aGI5+NUPzKa7pP73IrTbS8xSi3zUrPZWYhZSdrbcSRfC9w5jS/g
8tnFnBnu9P08Vc634PS9qWhbICVYgPgIDzqHQysU4bw/reLc5EPnCpAVo/5Mx4xQM3yoGjJS9XR0
zKX1ysjLwQByJljlZqHa7Usp9WYSVIT1d2H78pvjr2CI91J6PG7eGe41qvGytjCn4PXwsvMzrwZq
hTKyVNUqgxI3gaWUoqmrU4XevBEEVN1Pc9tZjxNN0DUoOaFWVXxOupSS+xm0OydA0fAns6Axe3E+
V/0EHwUXfRWXnEz/YXkDYN5WzHFbq3XMljoJ8/9DsuxdDulmLhFaZz9gZOYQ+NCfx88hmXmz1+9f
AFAj6RSOcSIDh1gxy+BAHxm4sO/8oTBMxsE800zl2O+uzAtL4ZITfsdzdNS0H3MPkstzcpy7QzKQ
3+x8pXLNah0xXDBeAyeUScDs7/aDzXKVt/Imfa6BqknZEsJFvXFqwXEzgxnTECfmgvZ1OerCXOlh
lrl+6G7Xue5NV5f2oq/x8uAHjALRkp4JXM/7RQxBuwr+zKHXQFnLbWpkmc7/5V4PGxhmL/QkWcO9
Vh738BUtUEiqM3BWCFl5XqiYJ9MPNNMtAKKwApOgdrTncDhQbv3+V4+hVM3pnBGfwQc2Dy5W+lPz
WklkM7X5FPyLvsxNirmHEEOPQ4Vmjv7ntjS/bMgg2UR/798zsGfY++fBUz7f5IRv6SeybzPAUGQ9
AoQyNa0ljOfoLcAIYSdCDSeQTtXUM6ZOL7BodXYZV3Sgcp1Dk0D1KIPzKQIf3ZbQ6FQVYs5S0+zy
m5FbiOcwo/q1GwvuTOXsNjDtDfk17z1NdcNP7cj9I1kx8e5IRCzKooHuPNw++O2YPnZ4yi/xBvLD
NqDAbRzNeDMHKKj86jmSjjrvVndJug6CJFRH0Puww012UonQLRZvkazTEo7CR13NbS7jQPS8mlbJ
+3xbxOuJkne/oS8fjO0Cjwu/LAkLLOdibN6I/DdZf0wPYqiXTSumRg66BE/htvLVABZQOlGmaGWB
lRPmtphFpkLnjr2XpwgPNG2fhru0mQXzbeQuVBciV5u55Swdp9j9t6DuweYNS+U37SKf1QmUHK0g
5tg92kubISlJXDHt87I/AxU3r7F2qwZ+FgUklSiT/ICvUCs8gyzxIpTfP8aq+UJFBbFuyOaPt039
D3B0LeBizbT9+obgPwtSYlKAl+s9JoqWvM6P/O/f29B5qbRfmbqoaQcTcDKluSHAG1/CMFOOxoCH
LCpIMFoN+1uLxmiSYLXiPRo5N/Mi38rFFMKsq6k3/yTgKt0bV1dx/ibeK7u5/hlzWAwbAUhS6Mzz
b4f3b6uUsEO8hQeNVap5kbB73yS2r9Dnqy40tkHxouyK9/dy1RC32UsVPIbysMHd69qQEmeZwOHH
GSI0U80lw1g2qnkatzgvKJT4xfCSPEW1OSjvuz7DuxAP5mxlZw2rYSvO7BGh/A/wJqbIpbJYSujs
p2GdZ0B2ej7ZKu2VSV+KNEM+iyj4t7CK1B3uxq8iVHZ2L0XLjeOiJ5sOCey/RC5ISBPUA5fC+RnN
1kENtldWmcEifzONiQ4lsEWUCJ03DyNYzbz6cQijLXZfyc9HdfnmnAoDa15L005ZvZ9rd+GoZr5d
rI2AK6xNVttNZNbZ08uqkxGYBDTFWYVOvIXHN88QH2C0VcWer2/nYhhdxOyNPDRdVXidAL2stMuq
zFI8clLpcSCkZ5mHXTNeA+6rute19U6njV5JvkyKpkvXo0BoiWC5JqcHeqvf1MPKdnknB2tPC8kL
nMPyiea+JGv7ywriCny0GB6dRw+yze1pOwUI9CtR3QhSpOmf2Zgw1dzo2thmiw8FE9GSYC2izjNX
OaM9I1kIl8UBsV06ZsqNog5YlZ0upvGEpLeHBiqTHDgjC1hODhS+9sxKZhX4kaqIYgoTGc6fFeL2
SRoplRCl5ieduhaM8HK4n/QrqRFyNMc7LobDC7QqlHd7Kr+7JvHjm4YlRHF2k/1SIvfx08/2Gonx
HAYw4Mu74NhiFRT3im0QMybj9N073SsiCPL1OboYF52RSi/8RSnrpwamFhQhZsKrSjRklRPqFX15
VHTqW1wTxddaihmRTxQe3WnBZlqBMR4cghFf/cH+rdAF6/E7SqwrOibvJBs2J8LkOxrRsVPtVgR/
bmumDtvtm7pUIcaFZhtzSSyPKgR8wZQ1FlJ5Am7Sw0MRU2zN3O0M5ZRqy1DP3a8Zp7Um9shLF+XQ
G9xeIfYsicNMULEKKj3BeKsNt5EislvOpg959MV6HDTn5g21d3Sr8YA9L1ylFxd0YoXYqXNxe8DP
H/7sGNK1HWobiWbklzbAacXUC3Ht7y5HQLk+VwijgzpeUxLHkL+ty0QjOj7D225fNXSF+69wQXYn
SreqnAYoaw2MyFIdUaCGMpcH3t0YxSKTip4fKK/qKwxzQkaPBphH/JE1rQQUs+Z6IbSCoFe++inZ
DRZi+sMJgBcm7CXbr54eIgr9L5rNnpVuZFNkRw1yRjfokS/GALeHiHFtfgtwg5p9E2H2p0TtzPLr
ofF4e4y45tH2+W1ljPLP6FF0iTpmaB1ufPaAzmPK99lJdyMIMT1hq3UFGqaZGNyR64lkZST914Ke
TwywJryJ4WJBSfYurv1TbQF8mb4nmvMpRoPkUU+xMYmli2wXKddMdYacTeRh0W4wPhpGDQUb9xwb
fWVWOQv3/Knw/tYPnBgZgwOBLI1zHqUAPfHq1EMDDIJxhy8rfpayUtge+roANPm5wf4uhRAeKzRT
msEa+eLS0lsCK0uQAn0eYEmmQ7kAhyUoA9TT+XqKyB0g+mt9ykSOJTOHb1p+9PlsXhekNU64n+OO
bIalC/6uyFkRvlBGeoHt0xsJxgDhzH45sakYQTwSekzhcuMrA5SZN5j2vpQdu4Dl9Ei2f/wHMpCe
cwKBzfLsWuvbBLaAISWBns+Ae7Wz0vv152NKqRcLH2xawV3eUfhQw6zHOzya46ZAtrPrcPh/e9/v
v676ss4NNscoPfdui6YtfnFJJJ/HXGGQpXBMOCDnIO7lCPJiGsmoWNOzvhySPQIIG4cKzr+KSt7v
cdvzxFWahyq3q+C1OJ/pfK9VqdKosEUp0rU9MnfQ5BSo2iqO+zztqeQO/7qEwxjY8OSWGhkB6ksX
xCAMmZu1HPFlrPpzZ/n2GAfz92z6IlUrNGg5ftR4lWHmBDD5aWfflGaaW9vW+TKf5kp0R7I+Q+y8
OKbIskzlEf9tTmnKAQal5EBax0WYmXAG7o7vDlymXZA3TXTIBAupSmJxSYO1dzkegGp1kp5Y8pQS
4aUiDyT2T8OrzwNVu8MnrQXcDBPuDeI9sqCcGwA5ZG/Lq72smyc07XzK0SOa1up8Op3ZlipzqNes
vVq6NBKD/mo2TvIrAueSLUmol78rt09Os/+JvjI28u973F3BTi4YwgTBw1mmBt1OZ8+6EEGrXlTE
3UArMwmTB792c/CI3CP2sFqCpT5PX3o7srhxJBHL6Tr1vsXdkDMZy2jiTWsb+Jigv7Aa7P0T7srV
yqIBPyZvVZaQBVqIY4mmb2LotcHMWf4xj0u2H5wUVUMxNM3ytYSNp37zT+wHAT2lGAII8r22B4hc
TyOvr5+/xCUF+UYuTid3oS7HQgO9mGm8imErvDSGflcsVVVgTmDzeU2dI+4hWw08j1v1lVyx+/8v
Y6ZelaaxgmwRajnmD7UaNNQ7MP7zRVmFHfMTKCvmKpqTL4mCE82kokYELK5r8kyvRY65YC73S6PU
LVz2QLapYmkdu3kltsY92CNLkDVMp3e7pBtYF4RqK8NZeNA2DmPP6M7WdNS1v2DP7WvGrd4kf6zC
bMb6aVz03Nq1RnrHYWxPUdPy+ri7qId50mCL5ISzIwZletRgqKasKv9CII2iY3fCv/gW+HIZ2D69
I5Dx6t4In4KfdrZPJzBIkaKPDqaaFOsi0NBACLmneYw4mE+EQ4RteRn2F04CIluS2x3IVunG3VhX
N5QBvwIu4k2MuDmse0UA3Ibq0UJuq4t/G37QH3kbsMAKMJlOG6qSb10Y7PjYpFJ0Okk1kvfNgLlb
C7ozjTLwFMXHYcuSAf17Kt0wl/qH+MuhPd71s0Ot3OX2HtDFquK/EEXbe+Ywj40KtNDbjMuzM0a9
Yk6GuLZb9DNfxsnDi59K9Fhyo2IE3CFDggLrFFYOCcO6d/CtDjaq9Wfh7NDJaMk69rHCGjffQDp5
bKzvZbAEOHJ1KsHkL/QBUgbQk41NgPfxw+NQ7Va9n8c4mJV1N9Wi/UrlzEoWj2Mnmq7pskDuehJe
l463dGifvTigAu2aBvpbQ6TtuGDGrlW4IWRWMbn8+u7prAZTFzuIzFyiCp5VhHDy4o6YjPTbWLDS
J00JjuywSTE3LgqUXrhoebenOWmE03XNSWtYhITMlTe/8N9nf5rvobKp5XuUjUeJDDKEPsfuUaJs
FxDNFan+Xu4ofZ7CKvF75bUcoHml++t9SbUSgl88SqLYdA9xNP+Y7GfnunrjE3MdwTiYukzY18b7
GaIiU8z3fFPPdPMcN7ncWMvNeBhT2oPr7GigD2/+x5z+YTUCYCxQLM4rE9S1LK1fI9u/Jl3aHpfi
wBI3nd9BLnxtNRDzDvJW0Zb777ZpEgDDQf+M639nd8LelN7Od3+rq2n4R9u7DHK+nAu9eFe0i8xJ
sLNomn9raXj6JfWvYSOLaFtoejxI18xrUxsx8rvQTNV5HhlcXmiLl2UuT+8eT41Q4UjZTHnpYQrN
fph6J27C9zcgHmRgpuk7+9ysGq2vOv3IC3NBXxvHPg/1RUQAQT260Tzplm0D0/Uut15G84i7p82i
2pcH3lGT70gXCNpTD32+POeCXhmYMmymSC5vqsUzJ1aLwOGIOIQHhkayICkNM8VKHKQAz0nUyRjQ
7PrWi8RsaXPgIz4Zz4pP4Q7T5QcfwS6jVWx9tHZIWm8vswmdQiDwkP2zykWlZxuHEveJp83S5n/E
fK2/S0BAoHQg0wWTeb4WhICwaDCBeAyXRB/5Gh+uKsL4Oczv7o8tGm63kKrXHMuIm+3qW+YjAmJ4
cmHdAcFlNyiAdQ4e1gWvWMRcLn1KxO4HA/YPcHSUhkNeFJJTZ/XU0cJvYGT8wHPegz5y8q7bK7wT
Bu4JGLx2y5nivl0vM9CkKaWpQFTQIZrSYKKsqj+YI/fQxoAcuLeNa3hr0PUN2GfCTmG/881dczgQ
yNYH9kJio7iWf1eU9/pjGorILQkii9AID+BkGoXqHir46VdA9wTvZiZRoBcIhIHV9Y87+LO+qdTM
wLG5pnLZavXnPsrh+amCQk0qp9CijqUdgY4e0ajRbMi6VITrnFclfEUQFERoRG7d73rUf03x84bV
5XVslVoLmoURJXLbDR8GY33n8Yc56V4f8eX2Ah5JRNu+gLqGWgofkD0ZxEm6uTRD0vskkO27f5ed
lxZqfRgS1fVyVD9znKLMfCvbwFljsAfKwGDaYo73Ln9MIQE0dh0RhMEusu0JEhNK8KDV4U+C3dnQ
Slz6Cf1GaVCdXRkEM/NjT0bgWYyse7ukptAQyffiXe32eRuaYaGbe75y4o1ag0Xll0YHEXYpMK9S
S60DKHyZiAgKhdM92UvBZLU2K68V3R2K9kvmMUBx+6ZNNLFjcL05OffW/wTByH0KWVTej4/ZT1w8
dihgJdw23dVoKj1vbO95+n9SXPn6M/tkt0d+VRm6BsQoRZ5yHtGFwd70gDYFldeb5Q/qKTHu2PSX
4mJ150QTGTJCOGYblM1hcASVvzowEVdpeTKvNWsUACbv1JzxTlR7/+JLYNyXJlfNgYlo/EoaZAUi
+BN65W5ws4tJJKRjLX1YBWdaG1BL/OUmkT71QZq5cSIgTXfItzBFYZpxF6EgEjsqlQ3yUs0G4iq8
JMMz2fydk7f6syWMuUYqSDJq4y9i1+THyQeAkrd6Ac1UAHllm/h4UEEIYKhc299zgX1iLDeox/er
kxk4AvA3THuDG7ProlG+kAmg902Ca28kVqV9cloHMfu8NSA3Vf8fQrfY7EgF6oYxiNJWYIAkVHb4
sUhCqQ9ivJGJ5QPQSHE6pRMJ9q6Jt2mWi8bTOt83Et3cRzk+yJNbcnhf6vKNgDfKqdPcJeBeX62g
430eWFGgtV1aEiZLYZm65vjJxogT1qtHuNYpYwdR5oQYKVP4HNYY8T/QQ49A0A6YvVaTjrfw8Sae
s3hH74PWnz8F67UMvdsQDHSR61eR8Tp97pdzrN7xM7+VAb3JBnelRyOJpdwDJTK+13wqD8kdgOe0
1iffsGZo1IeepvEN8RLEUDDxosrgFvchCYfNZuO8wkpssuIBAkd9sRCyXU7MDv2B4iRTfHoABAar
7VlBtxBG9ZjsCQUW0PPzTIp3rrZt5PzrfYfEXfBal7ghiXsJzaZdRlS5hHCbOjZ8NymUHxWXa2lB
aA8gBfEIQf+MGqJwA223irtEy5e0sysqFNzGGGaT3urL4mcE+wzxj8foJWLG+LpV0YYC+6saCapf
eZCxO5cNKF3ePSbkLiDzacZQa8LSL16CCSoTC0LMalP7h+E8yrGi1gTXDpovpbJuZU2HBi5/GTmI
LvF448uC/UThY5SlqEZ0c5PyDY5Pt3r3sayXznpAYZtLPVINXUfGM9rGQSUr2k/n4lCI1g3wpeLM
MUXSCiR1++cTF5yv8BcK7SZG003YPGERnwMlxVoMF3GLLhCR4hrGVCsGtTLVbwN+SGf47+uMH6Q7
hkwaojGxUJESeFR6fMpvkoV781Kz1E7Kn7PaIl6CXtfpJrO/MimFabmTK1QEmtGaTLdDtvJuPs9D
DLoWgghVO3FKaTKunHziPFsg605ff4MLNnSbd5SPLAHiQ6Q31VXXM3ZzBC2MCSA48hFeR8wAq1eZ
yGUwsS8NRCN+FrcWM6TqwVtgTneJiSNFjSqByKgbf5wQT/3AOb44ll3wF0mNXNXpJBu997kNvCgo
uG4NqU55HcABfW3aBFE2Ni5p8u9iY20P+41ec1FIP6zzTPJUhWdpM9ebEmCcD9m4r/rlBvCNmEZp
kSGfMuDdgOOqB2S9L8L83qn/+u9TY9HVOjhuRjOrru4lf3atLgQgj3r6fcNJHoCYIWtxKPxel2G8
YzZOBWJzVcF+fwceZfkSSMOnGm4QdMyjJVO2SS2X06R3s/E9oHT+pJb3Q3/ZZXJtUIgpfj92HH7V
5/mSJSxZH95RtCV8XHvoH5P7DCk1bduhRYrmuNnXIbPk5Ue/c34q+iLh9AFR+A5F9oPc53cOmu4Y
LVJgEj8gKDFw+p5bToaFpQEczP55FBeiR/Ntt1tX5ht1EccnDk5nRIGxOB0FtPTB8RIt+HWAyzWZ
Q2R5ydFd7t6t4KgQZN0Xhq4pShRHs51pREyNa05NjqprIrSqhiRzjjGh7s5Euj2m1hCCD3Pzeq/S
Ym5ihV3UDrN+/IlCX3W4UMby5Fc//yPChoGd0+d4r5iEXckW5pXQagak6rowF8tXSeGXF8j9AipM
7bpqbNd6kTqXf0e3x464kU6zamCVObVMRHGbyhXy3DuW1K6AO1R+c2VdTKFbdlPSRyg6Ueb9AZvP
viN2uiQjI1L5JNRqi6LXDkBgOuJlUAjwZTKH1/KERzi4yE3jWEuC5QpeqIc+wDKHNb93YHogFOOY
s76WV4j7NVhMhR7onTb6mSxcISEYcjaM17UI7fp9mMRm1oBeFblX79oFu+CMbyRaw/Tl5hqj5o/p
IWVmc3FYknrD7DvbydLrjQOfnGrZYGowlEGwarClkncomY5DRcJKPqtPZyDC60WT6yzJB8tnx3vc
jAtCdCpiU5jZUnWcD6xp7h3YwKFT2phMdbyNc7YB0JInpB9FUirXFLubIEk+Z23tsukKae8yirpu
MwiqPlVCDgKX6E7TM7yg6muOzak+r90vxC377mYaoYm1pqTQxmf897BXqEgSgXTb4yNZ1oflrweT
4moWjgtehKmdn1fQSINADwMxBGic05+uTnHnLX741vbmqpaVfJs2LhDD54KrgmNnTZSAwF0NUmdH
cF4PLomHoG8HTgYEM6c2SCvedROs89FUKq06UZWLwt1jSEyHIpszppA6xckvXAiSn/JGSwL+V5wg
oZ2TvIbJE5pYK8Ikx+qWbYmw9OZ2LpoCYI8HwirFvxDoerr4CZVfxeKRhNv8Q4fTh/tAzB+fAJKW
03zvJDJD9dHgvwnxrbMW/T/LYkD+eVhJCmL9mv8aQrRb3+ibVkge0Br0HUr4tnd7b3JZKVD0kPUF
lTmnrbWthvaIJocpbrwElEExCzmqDzHt9GJIYW7Q7jXjkDmTEXhwr04PE1fUhbwVtaMgJ0CUWj6i
TG4TIck89kht9MpW/lX3l6WyeHU1pykegnNTEXhP6mReWe7VtWgBDqCmRLN3lLK1wDaBzAuNO3Wh
97cm96HWJFTanKKgA9lvfTJXvJDZ5rHT2XPBQWwHsSJuyy2xKwaxJc3bzas5cSPXVkdKeJCzaYCw
+zdiXcUPJJrJr24TUIwpD2nEsynTnl48HExJ+HuEhdmhntdct43ADTLJlPIfP/COQtIuqR/a8GbH
YLzlHML9sNrLNxTPUbEVKWWRwppsG2ZZSYx2GTl5m8F9lXFDAWqIbe3sd0lkvrlBr9NKTmqhOrS1
7Ig/WSOlDPNVvTaqFL76mjb0O+s61hjCvyhvXvmZ5qr+W5jqq9nYxb0XIcH68f/zSm62uFv4L9cr
2ignWJ1qo9nQpdnah3cSJ2zOMywoZ+xJnNZQVaE4Fdl+HH6drG0bTYceeUG9KF1dhVHA46/FzWgs
uNg9bKM4ohpchVb0+4BWrTNCwcdhEh5FrymTaIXb1S3zdQEadlmsqjvWAXgaftCgdSQS3l+P0tqV
E9kdv0U+gr8jy60i7MZ/Q8maqk9U4qifhQ8kidC6ctK0ws1bflvB2sPz+lY+mFVXH8MhDkk52EIJ
LZiXCmLO6eyiGpiZ5ZamTPJ9OIYty0hp+b7x9JCsVyz388LcF5Pqjh3p7lPbSesw+hBp12TBbfox
wduWEewnolKR+ttVdKTfQfe+50z29hLulBE6h2jkxzUIVQv5AMWXyCi+Vs7aO68Dc7ofqvgmgNwY
rVt2y5tLxegjLyJ+sGFG21FkGYMA+vGzG+0RR8lwl64w2t54MZrCm+NApVhHIHdkueW1zreJKa08
qbpNBcQ65kxYmG0ezemPc+umvfvzAAkvaiTdMbErlcjEzAMLYHOksVFWuzGQRmyEZ5A8ZBQKkvAm
RNxc/mamfbynd4R+rmN1HThK8ea5O1XKDHN3+zmmawdXxlA5ARz0/N2eZiMgsOXKzm48SVCPzZPh
kJrAyqi/ttkhU88d04EWaJomFrjuWDDltphHBhYHNIvEOrMMsHhOyhLjzk/c8RjOhvAyzgnlbiEl
3McyqlVHvOd54O59Wzmq1aq4elUMkYMQ4hm4DYuumufzV1et2EBJs10Naytzf6A3H/ERT0Hgu0/X
rG7zPm3+g3SewiXGB3T2+VlHRvIeCINmsXa6xKYZWhMRlGL4PXcmjz+3gnaglNtxxjhHjafgaWrx
X2hh0mYypMfSvSUEWU0jE5o2amrWhpXPNoVl0MKPPM2T5QQM7FLYJCkGP4jITPslDGdBU17Uif2O
lwT3KO4LRWVOoBYpeUUPJpbo2KgBUk0yFYgJpVtVepwK8RLVyHhrkJO/VEL5H0QkG1EY4LOH64C1
8JtDIaYt+zkexirpRu3xs9UXUATVbU0CUMFJEGpDMWg0OIlBgCjGpf+5L640vBSA96hpFXHV/ekr
6IS+6kgh4CBOXp7N1y4fRJD4pvV4/L9QSVjLjXxvikf5l4qHcpzdWrjsFHXDNmRRkYq5ravyZ0wM
javoWpkQHMRj97KiznSJVVwW8QrLdiW5cXVCxxv2kZz0zeXOLwtyifIegULTSM6AifEEzGXgNfaH
yqrQ8mSZjL64bgMCFHMGn4K6h/il+O3Mk1FIrAwslFTftS4GqRclCxGBoYpv24PUb8IxT0NxSSz6
IxvX4cMR52VJ4ikogsQdxYmGmZXqswtPBElRf3dl3SndEyGX6OFcx+8LEU6Fbr0cfTmcFjWggwcS
oEcY8+knaUAwxZo10LkWf2DY09D2hzXtPlbeN35O5Eolv7n8UlUDxujVXDSDxh10/soVo8Xvr7Xd
qOB8L+BT2GHMcYUmgjvzI0WmFI6T6gmPD3r/0KOCNwx+weJvsXNMvuIb7PiSJyyuzk14Xgriw6bz
tNDpYgyrLDjP/p2nLg9sSAzQZ+RRGbW0KcFM8BTReo7W6XZofzTCTp7/u1p2PadxLuBLUm6FdgiG
G39N/mKz1PZQUJX5seChTBbQoK2ZC3LmnmgTsgG01gTPy2AGifx4tv2AXCN2/XXYziOamCcmRXtj
0GpDh+VBVxNL9HnuxGvMakdY+v57B0FxBYcld8dg/+yUC4Qep8BCGcmL3XSCihN7MJUiHBCiUVU0
3Nhi2zcrVKM+Rr+mU+dZq5B7B0e2u4gdX6G25+WeVSRoc6kMc3+C2bB6NgXIR+VusK5mjLrSZH7G
bLhgxQml7e2gMGxHPgwC6RtE4un37adIUYUiFzoeSKDhEpy56+FzJnbN6UrkjI3DuMpk3LO1UhYh
ssnlt+hAK+be+Wi49u0sLZpAaZnKHcsegdfLHQCwglQ1x6lUk9d/WPJrRxrwWCCgG/ekMRjyay2Z
r8cHVDs5ncnO7XbFMAheDLjYyLJTko8W5aPOWDAaZ4aB6jcCvzbNdCfuZBbZ+d9JJMOS/Hah3pdw
5iKQ/4CQbLXcE47rwtRcorVap0PUoQAbLzBkticV3MPO0zC9zOHjFesG32bWSJnuotucS2xkCbdC
z1d3VolwwP88rQ2QQwjv9ys33Hug6OBzks+2RkML3wA6KEEyAZtD8OphP6ZncrbK8IBDBP7i73EP
EBpR5xaRPuz5UdAZm+ojMPliJTuSlVIFOGm3OU1Gr/TdJoA13XIVHpjjKXD3nEmlY6lozSurWaE/
hd049lbWB5lkvAAyYqIn7t8iCOKQHlaIgB6X0rns7PB+3Jl/3I4M8fH6o575sqwbnA8Np8MRi+Bh
8CCGopW0PYxkJe0+DN2fT5uj/ls0P4OpUCEv2K9u34gm2vMYxlqhID4WjbtmtVVzA7fiFT4jskM+
c2jJ+1WKOSHTpZmpzjTrgyQxzT3LlaUjgppZXhcLAJLV1+9Vzp1mjHMeWQZx4mP4JxfuPVmhxy5i
XriDyi6i8FJPr04VqKZnS2iUJWGlJkzffuC8Y7xtYysQ6o0fNKDCo2i+C2X/ROWhJgd5gXWCIUTF
bgdP0Yqa8UJABXzeSXALr0gl7W3fdWUjP2YCYfk41Vl8Fzfg4YNDVw7vujmIpSn83xIzI+Gs6ME8
ocS78DRdDj6TbGh/C95LsTJFJUmPVwKfHOg84Iu1u728m/+XBjVqOfT8kyscwC97sSD2uRilbs+a
c6eEENAF8S0rNGJdzpMvxBBtLSaGvCmXrEOSkas6aloOFq4qdsPugsy/zcITkKUdsDsBMuWpIPME
y5KSnyISgSyPG/wF4I/wfe8KV926ilntwd2W03sFz/G3jOpQlvic0FIVXBxBwZfzpfF+jI4hzR2X
Jq4igRgBJnzWyIB0MzmsvJwFkvN4J0GmZR+zkgY9+uI3KtjWSjIk0H2qnlVMBXbHe1ELSDwn3lDa
E7PFLQUrT4ooPHjJGf/LEJdlzZGn/9x1xVDezhRCvQr3iv4TqRX1gcxIsViuT3+Ot/wKgPUN4/TU
Xo4EAcPEv9uPzNgRPVZv7CTuwo52ldK2Pu7nYtKoWCuiFXHmE8EiPllaC5cOfNgkPtg7PxT13i1T
bwv/PJBoB9nhoEyTnxaOZKMeP9qDQ0Pr90BfIb79tfyVPyLRAWXLgNk3ljF/rcrO83b6Do2QSXEV
gkxAOsJpN4UlTx9HhuRW3bkzOdGP7U/Q8rABxlgPwtxhGf7LNFpq0w6jSiLKnvCaXssTnH9M/cUS
ehAXZ0Wcnj5XRO0JkOhLb8vK1fGNMKQ7wGGLmZdCOIc+JIChmS3kP3ml6is/mEiEmR+1a1N48yFH
vPs+61w5FmnuMnK/Z+P5MTdiAgOB0RxKlYccRcDmGdfM1V1R8ctiAleI6ghKt8UnmmeBMcXgImGo
9AuLM/cI5qeL0kBmD17I9WZPgXvujIKaV4RtqyRlsmIWKYMjTigsEdrF+ysftYBcdbZSgOzU2SlQ
5H4+p5pB1yUwAHlFAvCInAx0VOs/BPf7EMmiwV9I6h0f6PuEeiwXFFP+by/kT9DWsiEd7ay7n/pY
6nFFAhiC4/CoybrMYIR36RLYCpLzR3Uhd2yDyV7cCR1GBbhYu4z4ud8lgcAbKGQ7/rH9g4FGawsf
oODuIPfvE547MA+NoZ0cyyCQy9YZTWKXdu+Jy1HM7dOTSK6Q2EgrY77Eq6k5bEKGiPtkX5l+KsBU
ORU0EZiUWHqUTjeHCMvU7inBtkaoiMciG2EfS+LWHtn83/7g3QnMAAR/iYBZctlsG8A7zUKeFtPN
dKLqqKZtP3jCbw2E9O5Nbso32KYEhtTCxngBaxYY4d2GFrXD6r7bKckZ8BuiFxmmVk0vQDMOauJZ
MAdiePlEHCBxdoHduSrQWMOtfnY4RDYU4aMnw6sEc4liceUiYrvA5QnOKgstuIFde+W/rfdaFmO0
ptQt/7pPl9lwlRCUlHAl2ycCu6jO8N6Qe8+WnSMYQr3CAWn8kS4NqUcl7BB4dXRNWLJXS9R1olpp
fgLQW0qB870NE18EaaE2fdqDubaGxs1Hr6ubpXIqD02nUdfmc+ml4tY5e1/1zvSMRbfoPeCyCJaG
KDKZfqDKfn8s8r8NiVVK+zQcmtWRcN9RK9ax6KCk5Hy/a7WRdMnhzpiVVDNBvxmE/Yh3FGzoUx02
fghw8TUMHU9RrRYLLsI40RrimGwcmFLAFVp/3pnhkJbumkqOfTcnbqOz1aVzsN7P63BmjB8W0vQQ
br/oGfoTa/G+DFs92O+e8s+q9UNTiJSdwVc7GDCzZ0clj7Exp+WPTVJtbC6NQVfEB69KD+B+WgUj
sD9qPn2S3Y3QvE/CxyPmVWl71FfoiIKdSZcV8XY0qNP8prK/7/v4474PZHsxkEJkT8CkkT3aNB/e
GoX7TT9Ly/DdfHAIsZz0G9mGqLxZy2KCnA69ehF5O/rbcST9kgP6wWBpwMgpUB6Sx6LNZkFPaY9U
uk+9KP8F796MB/spoLUQhOTHqhS8idH3pgNCNugG84XFGZX8BYk5KSf0SU5bbnIJdtAg6NtMN+ZY
KqgPaZ131QAOzJkdrlHu9hYRBtK9Kr3mNMKsoZIR7dQuN3RvYjWL/DOjvoNuELLBrCpjoTeJHF3A
HQYSxDO3q0ErnD6kBg+Z4JWw263919dmmvg1U/U6vi7CjkNNVpl0ytfSMkOpP6PcGpb5/jM71tcs
qd2lCmCWTib4GpTHp3ZpYe0Uf6m4s41o0EwGMhluBAkl0GumpfdVq8aVBwX+nqAv8NJbXz9C+ifw
7rdEHL0oMiBKiH8cPXAzok4SUkrDTDYiDQ+/lAYnJlFAQvqflSnFqdVmTl+T5E73t5Gd9+C8PtAe
NfE62T1v7gAR2pANU/jFpjR7chBk9KsNbDC8GaEBKkRJIksj3z4THr2nQ2zguo4AXAaW2QCx9aGc
6gA/E1Ze/CVeRMRjiVcAS0VsJoIHsBMxo9ExKnhmK5+R+5f2MBQwp77cgvflY6aMc+EH/ktxzBtn
QvzT0VX3zqIf4MUH3woENPLqLxyFz43KMmP5VzpPJuaUvfzOsOOhDoV05kc2FGttfQ+9N3tcAUFp
NJeHKQQTPwBMTIqAdswxtFZ5J4z3wxH7GH5Rr41SgyECpCSFGbP+xkeU6wRLfsMUbBJ5w508ZfA0
KDToBdfZmSmcLT37cVzzsseBucI1ox8HBf1BiEYIC2N9wAGZdN/oAJY/S1Iuubkvkjmhdc3tG/KC
CMERAEDeSr8t/KoBHgyQGIbASq3faI1drxWbaip9zBun5zF+5RcVQNLX/9l1We6o31vgVJKv17Jx
Kt6IymKtUsB0NUu5rO2v6YWMurQ8LiJqNx/UvBht9IAlCLn1xChGNJgMXSGYG9GWo+JlypO0znKG
jjXaBJUmUiTkY/XfC0sgobj3UUl0VgChF9FR4RiaTdx2Q43xKocELuc2FZGd575MiSz0PbdOZ3Aw
eNM0vjQzeOBNtK114PiZcUW60jkhLZqajZ+/Qt8lSOPsmd1Qiu2fcXrE9DmmyVCsMRhn6MbCBJ5t
+zVMCJqbyK8PJ0M06Gkh07sip7n8ytm4u8j9SbykQmsTAxtEpJI7kxjLl8m5SPLzmU+o8rdtRiPz
PzBCIJCSHrlDWrnUpTeUp4XvBgx081VlNrx0nyH3hIepvkiOiWcxy4/N2Xv6Y6I2GUoLXnb86U9l
f8cbm6KewmMg8SOn57BiFq42oPuWhPT6jdUnTnSlmRrzc09L3xJHWrwhTuUWShIqFKoOziIsmk0/
Cz8abovQGY/tdD2VF8dojTSiDtfrr6xmL/2+JRtqvIEbpJHkizEB7j9e7hX3PXdwDjNlcb6yGcQU
RPTv5/Lw5M5immF+pGa84kQBLPYloP8Gp4LPk1uq+Tb4pBm9t+cdsp5GIKZT1Q3KSFrQdmOnenLJ
ydqJFZ6Fr/jkSGJSBqIM7DXz6UfA6WEDx/4KCYtYBCaGNBrhKHcwn/9g6cBd7jqvRzUC9e7K4rER
O78ko+cCndS3qAEXJ49jUF9iB4YcDE9w2Qz1rEfQ+xr3qEax9NddkLAyoiNNwtjoo/yKmdTTpkUB
kh5fQlSVwYhIVfo77e4+BD1OxGuJxS3BsH+o9N5dFL10HCRl9QtmTQtBEvfHIRpzna+jPo9SQZz1
tnw1je6QIYcyaS+XWNssN8tjOgkQ9WITR0Ykn4RAIq9TsX+TweTW9XlHMk2fwl9H0NwMjmilap1Q
bocm3J9XBD83W/U8hGE9SziQnzXVbbwpis/c6DCWwfXmuLDss6yfhcyBeg7K7iFoTTTZVSX9Leh9
YPBQVbJY8xc23Ywq80YbYVVohrQMemgOEG5KPTYbpzYz27GnFpJ3Z5ptCITkoXOwOrtVTvoUGdo9
XAxrbIQjYJgnc96Scs4ko0WxxoXdWm95C2Z4QBptQZ39Uo8pLsWtIS2Y3WcYheXyJjGOW1D4SBta
16ZDSTl/fgPf/e9/uYbbw199nOqXdPSr5fuvIL0DYhHH3evLjn8qoHVGXB2vmq6+8WN5VHRBhPsn
2hKG4JM7SAhqOToNErVhz7N1mQN0OZDKzP64DLoEe2SCSB09jB0KH0Tb+aRsHaRjRBaqeoM6TgL1
oJTGWugsEB9Ugb5nLHssZsFr0AiZ8+sCcryPvmCV+731pzEY9YSEuK4I09m5WWxaE5DinA3btKJk
FoqJioZ7REKvZyfj4QVv1qyoqpIOjDrvWlEcSP/Kdr4DQrGNd848s5bU+5Z55na9aw++Erg5Lu7h
N8tjtk+GviYAN2FK0HAnRVigf7Dw4VJn7TVDqtit3cWV57OZe6gD8aWx3fd8lG4ORurumoKNX80D
B1UGvTai0XZLXuB1G59szpZJBW3HPy8tkxvbOSCDvKJlFidmJzUOug6OjMgJmKWBoRfsUdR6jb0h
qB4oY/Vbrm4skN+kfLidlVrQzwFwcLp9C3LnWt8P+9IAe7vJvL8h2JpUEOvK0r4e/E9vhouwagg3
kBFU4yrJahs65DIIbhID7+dXWx1i3X0Rmx7hEn1MyiHd9LyCpsPxwrl8m+vJFsDKSff4QGbd04NU
FQme2LgoqIYNcj8y/lUoY3+Naz/I9QB7dlu+c+VmTkD3FewUVtuFwpB2Ua7/TedNSBbkUqvPO7HS
pZwTVwYC5v1fyojrLlaMzqKNCK8I0nCnISaThsYpew/ZGOVJdqKqObYt591Iv9Hz4P4mBkSbFIrj
nFSDMXKKXK5bSOqXMS6sy8aMA3UOm4GhEdjRq92Lk4KgbL20v0DjhQvW/A/ceSEs+ofm49+3WweQ
u9Xwnr+OiMXh7BVT+SHqhPuktCZw2u16q/hqGXA17TfYfO6XIB8hva7HgVvwVdtFSwoHxrBX9lHN
HUZFlTTr8m+q6OiP1pxzwGnDmv5owlTW0toNVc1RsYMaC5wyZZHfEJniFamJ+F5CyDnGwxn6tWTk
lj535kaEXwWlyBqiP+tM2NaY6u/nfPctVs6mZD3zmHnfC6FdWG3Nt0heHNzs0zEjPwJfXNs2IunQ
tAR7IEqEU+EPi+GdUOGA/YpA26h+Cm8o8kiwUqr6R0lnpLgUtn5VJaOXE+FVGcEtWMjnQDmpLTwP
lf1r46cdfISAS1DdW2XFPQEH/Is9VkqHZg5sm72zciMFlqiQ9ymMdxPuQj/LDdjjezGNz+Fw43n7
8kLjhqurgYulnyxsOpoB25ysvSwJv1e10jUZRvcjQXWOBjCOqQlLHd2cSV9k90UKvWEHhMotXsSI
3JhT2tmnA6MzA22UHhlehkIu6RP4RPm/Frh1lx+J6Z3utfebAJGnaMSmdKmmPRJudniXhx0jyST6
HoH6VOPYfREe/DDsk6CgCzV+GbDZMUTaemr5p2y6tXPYED7DBX3PBCYGOgsy505KpDS9SXKcgV5V
oxOCHlgo+wqzlf0SSWyu1d5TzmXYNh3NeZPTxAUirHP5xNPCeFUlQKS79yCJWqEnh1i9rYCxLxMZ
xCRhVjpj/FLenLxzr2t2sSGPRS5iu7DJ8FpkYbUF8IuqSv7a36aiUbb2P2Nm0r4w4Rs5lTOLpedH
XSZLohuviFFUFn/kMEhxYYeJY2qTLL/D/yyMIffvo1ouxlJZksasq2VdKq4/dfQRjfWJTHpQtyOj
Oqxpv266qCttruuWVZl/ezRGNsxfVnKVgbcFRXHaqHc1vXhUnq0IiGAxSDF47z1pOMhzwWMKSmga
CEbTuz28YCsXjn3Acke+LilgVNuBGlzPzAvCw8OiYnHxXf+YUdc9PA4nLrZJilQkvLKSNRiKtjhY
60jrMddWJx7R+hvoULqRTW+yaic5XIbsJLhO+iQVr30pFDcD789y65dLhvv4gVIKbItjl6nF3l3B
WiHZKm/JelEVZwCuKGnPiX1beT/81kQf93huftZukpOXupY1Iis2sX7ZrFgorMqq+qbyzLP/dUOq
pnmNkxvNuMrAx5KGTEYg/W3kgncbaevvDC+PwN/jcL0Wfp1J2f8/gOxh0eHk4AJPfDx/7yU9b+SN
w+h8T7nkdqEAjg05nI5VLGQ8SbTeRipH3Y+Yqp94mIUpJtysY5na+nAunnagtRNBWdMzwucLR5JU
NN7UbnLmYzA11AKVqvuX3t3EpJCoed53Oh0ZKyEqKqoPAWgpxnwB4odcAOQVtkOJQAtOwuwqD/an
ROvVTxdQv9thQV/uenoHjHcE26dpsgNFszu6naBV098upFYmfOrcZz6KKvv3mWaHKgKBccj2EUCb
P4QXp97YVI4vyd1djOmUPhhsIjjwvPhyJPStm23iw05QuQAbdnCy3a6YVN4HaCryXfiiCtq/2+/a
aVTkeZFP4pf+4eUtg764i7uqwfhOp67yKAwhGJSy58BGO78PiE4Yr8ZQJaRYix+OAd2o6ZzRQiwz
IsIFG15/sygHnJ2rJKP643wCKSl2HkrEVfwbpPelygLSoaCAS1tsqc3HfR4PfZLQpaBShdMpZHKL
U67rxfHDJLh6M9sZkWeEF0pK4L1xbWmwgrp9r1ujUdnpE6RxIab5xY9c87tBPpnXcAbx+owYZ93a
Sdovbhew6LeeXBbqskyZpykWZbkPaaRv3EscqYaYX/5hbz0TIDpnLZ943ktMygdMsB7Blc2PI8aL
vH0WGrL5pmPvdGbDgaD9lU32z5UYP6ExOChYOCdeIOmt4iJjrTue+KlhdAa/VCNwDVwmaIIdPdlF
/cWm2rsgJONjfPsLIjEwAatJd+AuGZsznBZqEmAIP+QPfkqzmE3wOYOlJ2+p867ApDXOTzkDANUP
7kEINJrdeY9JAljZ7iCaJ9OVnZbWZkIcNlCllf3hlwp/3j0/GB78WE6BqtUtSGgKtxW/ODiNUkni
ERvDA2tLzioyL4c3UHVCOMvulJOn6618njV6l600wsH6RJj3ZjZPiMLT/aZyCXBLUTyH5DbttcsY
7Ay67FaOauKF+z6ajUOwOKOE5JqNPrAjApJanVslNtqtRO6XOeff0+DBt6eTpNqzqL7UIsuSME4Z
RfNl5EswII7wBKx9/ltJfMzHBNu5KIvijKSNrgoV5x3PQne9H/jbdFtD3/23n+Y/n0ErnjRLhh4P
l2wMwwO8vATih1g8Jh3PdjLwcum02czYEfN39N0bqDFd9PhX9MPz1KpJBx89Ufoin0sDLN8usA/B
YjF1fzq1icu4GVL+KhZqOKqRJxErhSQijSGz6zo1goGeo3uwYLrkPaNyS6K5qstqK6MqWNjM3w3w
G/NgF8zhjS3X2ZJ9Q1tcd+4e0Qot9ZkwlHjI7OLGh7U/RQEsLDsc7H/hxljJYaTZqq5KS90IW9AJ
u3rPG7UQEkPiLrYuaxXeYIUHfKl/CNNpqgiAogmTHRzqpUEw3zha71vVEY2yW8vaC+y/C3bhYQof
3ugBVrdBSQdozS67sLcE624rELmOExKjfyARSHaWJEWOaZy2TYM/O6iP0VvDlahXbLjznPPvkpEZ
obdRVU7K0nB+5FHWpAch5bzEz3rD41aq15F1bu9mSawgl+IXHmSYBhYo0PL+5R6e0+lJeganssuZ
2HmhZAhXiC6tO/2TSrXdCwmFOQac9H1rzzc6KbXL0e6E57VYxHJTsZoXkYSODOMkD/XUuZfoCfSF
1lhUykgTyLfUSjr3Dq/eUZxCjhLw3vfA3nRAocyH6UUaIv1SIrfmHBZMQr0Ghz+ZheQyOFJLr7gt
eoZukYbUgBSEtPTEXFmn+WbyC/rzqlzNivADWAk17ygyi1buYbOp0sRpcKRb2ycEcmuWQ3ElvDGx
LrPbYpL1wbQld/941lPw8ygtmWIxtknlqSYa6rlghhfOGQwkV0vp4gIKaFACrb7I5YXP/oHAOhL6
/zsYX2MdRfZXId+6lcp1mqu3FXPa1syTBLh98u289DdeDZznJrzKMfpVB9WU6ObifmFRhNz5NxpW
tnoaUPiHk5MJe18JkcA3Ek9GVLI5Bi5paCWZAqbbKOwjSUy2Z4JupmnQiK2EuAwjH/TsptEuCRrS
tuXJTJ11z/++xkwI/AuIgd1RNdxacbcoGNEhdLile0L/sQ/iRP5scfLDK5FPIyfqm3SmbusfuI/+
Tyr6HZD94lB8ymaEmHgTvPR1sfW/l257D4hZIrT3A5Inzn4Hhz74PyTRZ10NTLD2PnsdMBo2wOF9
nV2avoL+CkSfFqFXtmC0pKcBDidQyecp/0tzWB72E6nlVwOjCzLig5ISqwNdeZ143aINXkfGlhtr
fXaTG+LC5KWWaCrc58RsLjEBc96hwD2LrAoMECLFe81t8QcFLIP9wOJ+48dll8C9GZiVUjxLuZ/j
vshQq4DrXxBefu/J+U6PC6oQnaz1/ZWCBUgEtij9XxOxkPO5Wry/ZuRrVPnuQJAWlErk/5AlSLYt
hqTvKz50MczR0LWkG6OEi3Vj97guK8cqEc9MdFDrFAdwCBwJ97wsO77aCptw++zNr02Du4NQtcT/
J2Xct5D6v+BcjCJi+A0Tn8K7/2antiQMexry+oUireSWIHXAYoqA9WjAelBYl1Qfq2Q9hPQng5Lx
pLLQNsDOwmCMwg94PcLahwL4NLACnV0Wc7VpcOJoA8wCV//S0+H9xgcYsn9ZclQwiElYp0txUoJb
V5ni/8cSVe4v9UUMyNU/+DxI/3UfFjWUEhv2KB/7gXepGahEcrI3DjF6nbIJdc7stit0gshY04DP
gAS0FE2jhLRHJln1fKYRndJfH1FdW0hwjOOZlV5vyx0OIFR70H8TDPK42iK13rn+UiLfuMJs1QXv
ve8ksPd7l5I50flZnljoO76WG4g8CAXDAbNVClvktURCNWSotI58niTWIV5VGYip67dNQdeEtEup
SoJf9zXiDYywOl4DYw5NqYKbcXbj8G/sTcshaU186n1lPBTAoiNtdU14H5k7OEFUQ0bU+E3+cWvr
oBsCG/irHYgxstkgrL8ouu3mqBlPTI/pZ25DE5Z8NayRkNk7PTlk2+U8xsK8gUv4bYwHvIPWfVwk
dni6y666RS6SsjIcf0aQB5Qgl97QYIV07+PQ8lFJwD70sUhF8w4pr0o4/4EiveHnIp0oIe1FImgc
Ku0nNUfyJqqE3XOyUvf7bZWy1Un4KmnxjH3llwPQTKBc33WN9a7nHdgfWdqcS6xuYTwb/nCCBHe1
hy/lVT1/TKF+3v/x4RTyMibGwDsq7ZRFxT3mhp0Sm+DQAX5WH7/bAx2k9Yc4IcbFAeqJIPif7l6F
t7xZX9g6h/MzboB7iDyT9a8FZyVyKH8G1OfWD6ngKAopkr6O7O3IVwCqd5oTZbCJDncy4ZRta+AX
TO7vmDtwz3jWlJ/EUMcmDAggiFAKs6d4bvYXQfO45BC3826On4OqxJMfoJ02pr2Z/IgrpCAU4M4C
nxeizm2HGiIdom/nLt7j6K3zsQLuiUBC12zpM2SiTD9AdY69RNHiXy02b3tYiMpQKcTByIdwfzRm
KmwybM3blKQLBTP8oFR2AMqvjHe7hpgFzcbnUJz6gCo6OwEo9lEYwjfUA8UbaVGJGAAT+wiZNgg6
EiZVYpwyfdpuN21JhTsuQ1HlDHgC6NROZeJAjix0oMo1gJqm2Ik71yWIdENesEGUxkzYAF1wsasJ
QhqweaJUmKJwLeQ78LKWcZdxNLx4+AICODzl7U8opVvwtxI0a+UNhJtpZQGUsKgh3FGTJx0r1RFi
x3Okfu6OkT48rdiJm19WmzSbdoPDflTOHeK+Qy3zcUDUCBb6M99FzesykL+hRmMHRS9Vwa8jzXNa
cY+1CVl3rcNIftVLMq1z6xqp0SC8Lz30u7UGhYs6xTqSyXRnSSVmKBtH8ZrK99lKKaxq9oVle//0
vO9CAckyoludeuG4Leqk1aPH9vW8ELn/1lSfevQ9N5zmvyf5S2qFOtvfmLuObSjzZ4sEVEEoVVNC
lOmMbqZVphWksA35y+bXmbFzAFyO7hKRc5r3PX0DkBxXOwWHSb6qLWkiM6H281pY78U4Pl5oecsN
PPi6kKFvcDWpZB05NJ4xMN/qxTWEqmGAcdpSRGylmbMgyPC30nZGosKD0qPqlB3/sxq7JrVDr+RS
8Yy/CO8pOd5yMOkSmXBfsG5RFSvW9oHreoS4CleOpYwp/TeWav+Cho3249VmecjLK7bhtOgmH+1s
C8jl15m51zLt+thM7s4y+SIgT2MjM4q0Dt1YAWc3JMiVhvgusN6CWMWHJKzRbXB+dnDu6qVYx/Um
e0pLROAK1+aG4u4RJhPq6fUrMf40uupwSaMsB3D9hLlmPU/ilx+/WmSnbctr3gsFqXA9WcW4Sl6i
KZHJKUkfPYQTnJwrzS+hUtVZkWLlqixmgeHNGV2SMhRsEdwvCJRn8pdZTnyW61FOpGl//zD9T6d3
uYk6epvhf/N0I6SlvlZDFX3UeinUWuuxNRpwFjvprp1UdLCxEf0KwVUiWCPMDp9GAc0+yQ5ufb4G
gyXg7hLOxX0mmLgz8Dlm6KGugDs3KW+IBBrXWJ/lU8sgfGjsjgwPxbBiYxWGmCk4x2rSzeuo23yY
f6zjG2b83azmjXdZI1SuQA5eBSdb98xddiIal7vTq2gkLbQhPQuoPMgTQ7O07ANRg3xjKJDe1+HL
Bi0vNK+1Qyryh5X4fg1VhglD6RIo6RWk7Ect5pChl3uaqA+T3YWZJxya3ynH/voJxdOgdm2oNDyh
mD98byVQXcc7b/cVqzpP+jlljgs1CWqwOo+iDLRmWjuVTY249ECffoYy087lRAEZGAp9F0KxDvH3
xsFC3Akj9XZzC9Y9wyL7kFlQQRpoBZ+h40dyZUa3gOj7dhxzw0PfdrJJyBFUgLq6aYro3J+E6oUm
uTzf0KzVD0exqv3SVwNjS9/EngRArca9R18tndY0TPnO5rcxIbwI4eqHyzpZk6XhBu/iilKZcKsN
LIBY1lftJdktDSQYt857a8yK0HRVZJiUFt+ronF6E79VW5n18cIu+jSaDbP2il+IHb8IjNOqpSN7
7rBTg6RgFMruXrzSHTeow3GsrrrxHcmiVuDqBkJ8kJrG1wpcXEGuRC52P4U+BvTwCggeq+inaxO2
gHsEWUydGzEY+JfPuO+0Y6bwJ9f/OfdK7qvQ6xy5nmWwVlwfW7qeO1fB4ZRaLEKuQ6HwUREdUiXs
rlBSFVxR5+x7nWrIBez7OcnME1HIYO4I33OoCT3WP5zIaVFo7KP+V0azmWlEBbKtM+0hjYB/DxId
5FjvDumeKO3SOh3b+YHgMUZWcCXsytQZOCFo2C3UyrlV/M/pz2YmKReiyQAq4pjg23r/psT2YvEL
j1O92Q9bUNr5oaif5WrCs2tJ8BRF5IrjXrSV9chkxmgkCnPR/XtJTAFJ8YUBL6gxJjiWELmFiHxA
EK9gfDCW1UQshPDkPX+NpRmz8uTGWRQEzJKRM6Rx6t7hg5n4+oZlTBngFmugZOg0DRuOS4mS13ie
IN3TH8QK0+PCYjPsQ6JTqR9pcSuTLa4UM+j526m5iDHDP1y2wNM1eNwJqpQyTXPlAZ0wEzHKSHA/
gb+D+Xj18GPZZKC//6Tapvs9IxtcmerLlpskStrgJPIua2cJQTqR9Y1/3ja8dnqqVLsuDPWjxbXX
mt6gZqnV8UJrTO2ILJMqBbtSsoIp/AJ5Q989CYzVh0o9j11+8lHs8aqYZ9roJYld0AY3nzefcYC0
UEOdP2ZNKqNEWfzP4JuWSWtfuGHwwULgpEleLxz0CwI1Op+BAKO5CkstvqfXYERidOwHwWydnF/+
zArGU5ScBDFYoeK2/t4NTXIGZDfskKvew85smoAdogqd2P61y708Nj1rxvi9LYIeQ9IgAJ6AnOYq
HWmisNs+Lq4qgg/3w7/pLpBBMbxCQU/vkTsr5+NdhY4syeitDoxWnjRjCPmimzcnYRrqLvAJEr0U
1D1prkcb028Fsfb/yTX+N3jlva5cZqNwJYbr94MsK6LfG8QMqsrSdIsvqA3ufr5IR2qgNoN65uFh
zJzSD7Q6Bf/MNqELfuLfP1P1csnb066MTEd7Heh9QMqctDTGL78+m0ifEc7RwLA9JKCkaZlv8vwL
kci1Tr0AW8VYGvhmzuPKhZ+wa4xXP60UPxRg0fKDFm3G9JOEYrP3UTYykOWaW/O9YuxnC3PqoU+O
NUFyM3/QpNxqU+I72o8wnx/jWvhYLbQK+l8dx3ePGMGUch4TzbkkfWy9PanUMYIdfvCTliuSbkOZ
ebzAMfrRJKNx+Y0HRB7MDz6IUdP3baXQeDr9wxWxSqkJuWue66EiE2JEYkh9QMoLVM0dMZmKwJXb
qi8t2qW8pIBYgqiI67BBr7Mhww1Bd9+xzfZ6aY/3FG/5Edf42N1m++IecJev37EqDH3dQ9GIxG7Y
YSuNTT68rXbIDVAGZZQoLC3B77uYbeNjitXqxrxvvfDDE6NAeLOPGq0vucLqx3uHdmK1QQIRiC7X
nhmRFDR0pWsFwK8WVwPkhx2BLbVobjmsJfs6nf9o1wj/StdBDGjmJb1+5nTRERCs12QP4V4eRVEg
pzyZhjHz32vkOm9eCPj7FmyC291OIMTV3AsszoLi79VPbMm9Zn3SesIK82ib51x8L0IKwrYwMy+Z
DwL2cecxGLgPBdLkZmQjViwKeJnWd2em4KkaD5Kj63nMuZAAqfNAXdg+YwCEtUDRD28hZNqT9OHL
Z1WJVhujAa1zAZP7oiz4brnLWz77YSp2HadYOfSK0XiLV5YlbD97B5GDsTGIhz4eRrHT6bFJbSjR
28RCbOt07UNRpwYZ9wE2h69zbZoi55q52cDjnbwyi12Izdcr4/ZzIFRbYkStKhj/MJC3IepiGuuV
A+hvlHc72juutxeUV90vmHRhv+gsdf57TRXHvUEAMImCVhKpfHHe/mYrO91pOJ2TTlAmn3TarxC6
dLqjX4qijCNXRd0aUZbP4qF0EVJv3Ielc5m3RGUM3NPPK5jhZeQOgl8ar0uiIGATIP9KN9YjvC/I
bQjA+tXKV/kAjR5KDtQ/31lUKcmylzWtDIMaxYkyjvCfKAxpx4lxH/yyjCgP8D8/IDbOSgEBw36k
oGRft20UM+cVcJiKHVsrfTRAJ3Jt55GuFPPbmIANk3J3SBn5zJ0QL5IQxnoRmVV148Exx5syHVo+
f9Viddz2cxRQ5Vv/RIgkyHlO00mcPHRr/C/cxhpfE9IpgNkD3lsktl3ANsn7NTP6AMTX0AHhmn+F
YYsa8/cEPddmxcq/tU/cb/VooOPyPMSmxx4Lvi6KL7PC/MRBlp+adfiTgswqKh1vkohldlfzl7Dg
fBomv99gTFMVcFYnjFSkYtShN1O+0A2qeHktuSPV3OYsuyxJWhJ41tUY1wQffk2snIZ9O1hfl/qu
/UJ+z1P1s8N2z3McSTzc3zIwAkho8tcxqCVITsyJxQ97ZbAokGSprG4OKsfm1QPrvBW1Tr1ItoDX
aaZJ9m0u2QAa/3b7mJ7pqCywbjcwhvPHMueB6sxNxhBzD/Mx3idncawyYma3PYAJEEcIvAmSi4O+
1VtiNBEhAYL/bEyAxYgcDbLrxSkej/jqW18F/WMrDYRyajkhLs1hWQgdrVgkV8fe9drv7y/z3Y7K
B5s9vuwiTs6gd0MKZnd22nN7/eoU5eMDic708M6QN6gLsJSuzS4Jf9GibHr2RSz6j9Wk94z9gUnx
OJGiF1M/MKIT3JyvW6/ZpVm5iV6zlGlgb5ef7ZK+SXYyvM5qUmWfKsheHgeexl3I9HAYWykNiqP7
N9nf4rfxio9mVhqCzHvUmG8YAPDtVs34+J7dQzzc1qCzqMhia8zWNatUKhj23z0v4EUIPZfsFYSn
gZOJ26fiJCLzg+3Ff4EGWl0BvlWaUk8FPb4ji1KAdn1y9nM7XQbuejb1uBUAhCNMnZsGTC00Fs7C
7toej2nG2zMnu2RQ59usIUiV0JgejkQ0zpiL1BeQoSd3cMKWZtHcB1rovZQ7CK1OQKiJPE+u9ALS
bJXr+hGLjXvaBS35G0BwwUPlJZI+TG0r2/ev6yycinGm/f6+NWzFpr6CxeOfAadg36NNXJzpDQ0N
3oWA6K3Yh8NEAOEg5rSjX8Y7zQm+o+uvu5Z6rmNLkoMNMLzR1RjUItYXT6YxsLRQ+6UFtx2PgV4t
voAVCo5YWvr2TYR1hq7MsShSZhDwxPHGKQjCsItULUZC7SY56NbQQKu5LaqAmMBlI1g8ZVsBacwP
ELVwzHdKqfeLLCeUAgQoSKxQdWwCBAF0Q0c0IAuQS9zaodBU+NoBeZuH5ujChXSQNx9NbEOPOt2T
abCW2/nFsrCkwqv4oiv428mFwLXrhqv97tiykVFlTfAR86OoJlkY1dmZf5vCIORTO0hR2lXVHisD
q16NUUBiIMZDFXWLvIGs4iqUXY2mRSQ1mVucS2xfZiOHm7Zl0wrkBuZrr6uzFFnQ/DLztEAoxY+V
S93RG/3mtvqBJPP1uiuGcZFIp+QmmcYKEyO3fXpaHf7fcMVAupX3JQcOMNq3Vdfg/pzlWNjHK9om
ZbGLFwwlscAx5wiHsgs7EnMpirY2s6ByAYXP9I/vLjEz96aJ5uedy9qaTxNw0HwbFZ86Df2oH5/m
anPNj11zxBWOovgUwtldUGJYfOzrgb34L7CvhOSNjYk0Ra2c7NJIz4y7D5L7EMlFuhxxUelHxRka
l/oJPalwTnVDUri3qObe+N6LjRkEn2Ja3zIrOnCMNVdTPap2RazXSJPiG7pWkJfAZ6c1TAdYt7TG
/10TU0aBpCOfxMQY37Yc9duaTwR0ZASngJYK5bO3Zj8VeqwKH7aJbG8IuHy01CdQwJdG+lARKhS8
RqEo7HAYTF8TTYZcAxhMxyZ39QeM7Ql2EgH8aUXU85YB+AtS/lTDTsyT0Gke94NMm27GDvDQXX4K
3OaIhaBNtbBA8tAkz3fdd+ZCYnqXCeirHsz4Ylvv6g7RWy8Z0Cb/LLViCzu0SprxnAM5o+5Xzun1
WBCS4h1i6JBeW7tU6U5U6svXbmpKtuD9AwlmVpTUus0KP6rAsc+uP5lVCj9m+M9MZIQ3H8e/J7Qb
uxvRm110FlzS10bq6X9PxRb//PnF50LkUSbHiUOsNlbzSU5rWkTdwI6ZpaPg2gUarDgMrLAyHCBL
fFp+Yi9tFgC6PzbKqwVSvF0dhAVwWB9GaP5NSAqRXwf+WAAOvG2GpafhQKtPGE3HifjoJpCF43aD
RLafzgiDt6yLBM4vQhIdraZgHchuIregWaCg3ceOoT7wTHAuEg4Kzbch0lssFNEzTQquOyS0gXLI
adhBjMg3dSi0dqYTQoRNPbasIHetU2lJBOq9Pw9YmHqsKdpvpUBD/Sg1objoBw7kztKJFerMmrHw
7on2YlVwSV5rOBqC1FqwA/EkxZyQxF6XDpp986MAsTMQhJWRvJQIbZwX01BCxa01X0OEuZ2FrsnM
w1gYESW93H0zw+GR95tgmpXWGP7yMmcEcjBYnkHcKgLL3Wcu231JpwwlbL/lQL5KQIHwu6EXJLAY
dHHusGn6+/FJFrNd6G+QzJIY5+f37xs+MpmISNxdpIcPQDHYrFTpnSDoQCmRzwaVLPMbe1/Ua3P3
ZK91LlnnXG6m3pi7FDkXorSVR3ldc1/cqsx43jLO7eqHPl9tcuYtScGRN+5Uw/IEAQoA5zbTj5UV
Fy7UTnQjh5aOi/N+seoLsZKdPUfeuQQXUNJvMznoVq89JvrmweiC7zsZYSuMqaohE8rf1QHkHvqE
/PPOlg8tCK1L3qo3x3vIoiU+tEzjXENSNC8RRHcMyHqeRcPhdBErmprbZ6pObNOHtfTXDygLSWEK
QWHHeC0xgqqZjOXVKyihB363VTJ9oRTdThHmli5hTI7D9ur4c1NWJ5dHLz6EIrSJ+2YVqED84MmN
N7/vWPRHfS+ZEtz+Mjc7T3gnT3Pkw7V1EfUUg3jeH/VGe2c5XNixdwC70vIdi7mt2OT3UJhvtQ+4
tfRdvyy3ZXif9adq0pEq1txpr8Fhko/R7IbkeM3OGY01mfvIqr1k27neCd9CD/pnrGSxEczwx0Fo
d6gswyzEJD1KZ/k6NOo8owpUs4uVmoM8i8Q8gP7NEtEWD6Wj/K5P1Ht9U2JGr4cmzhjJwbulodii
l5j5g6n45c5QMBVn92N4nxHw/5YrccnSuBYk0RrjGE0w4hx9p02aYY/gOYpf4UWG8NL5pF92YBz8
dHL7FvK+UW6q3zjBv7eluQzxSIMd168a64S6pWk1FRdfTkK2XWaXXuwfBX2sdVzLRsFrUBq0H40W
ntIcQVfszmfSP89gnOFiEg01xLnJ/hOG1wOsPDbEW+HZP7C2v5plaYeI9btuyL/su2X20dkZ/6Pf
vqUV3m6MBxOGzy4YMyYXgI5V4E2lENJ7yJ4aYpajAafTNlQFZVk8/oEGLslOiu2nGMKmtwi8ejZK
Lgc0k7LmJk2/FNhyTrbHbzBcjmdes39nMsEjGyvNipIkIBUQXldLPAM2DmiLSlYJYMI0DeM2zvvU
kRcu9toIi5DQwOjsMqQXKKY9bfFOxlg3N+KfzMJfj4dSxbiM7rM1pgRma5TTqmt9Y0erCYRhnjWE
UwiNc+G1v3L0Ch+t9seY+ESMrIbLYomqBMykR7Qz/L2HzvVwi1RjXGjlpen/5H9oO8jmC85sM0VI
UlCVcPeUPF0EfYJ1tecVCgiRTcJcoNr6/H+j/AwlARZLKe1Z0pvNaKDdHySaM3jTACAWUcqzG16/
qM28n4Oy2V0eE+M5Xu1H0DyVU4V4WqJp/hp8R2KrjM4YiafrWTKZ0GXVPgSRc+cCzQXKAaTRXXYr
Y60ScO9x9m6r8+RvyyIbHjf1asE4SgVi/IkjvoEOvSh/scsB6E4lyuPRtqqYjQAtHwvqwVTAzCh8
ZEMe4O7Yfwi/jH6VckHuESqgAWjcgK6XiTO/oQFspqBPxz32b9tZuoQpmmYqHjMt+a3r1kW1demm
XQtS9EDTT44zYffT4n9Oireqt/pJAeuucP+oglQJ1iZFf0Sr5pQUgewM666R30KW0RVl2dBKkh07
4vn5F3Jt6iv5XavYbhJjB/+oyO+kB7VYZnPA1j2L0hFmsFYo/R7y2sBomkxYonKqs98Cb7h04mqT
DWNps9eyj89+jlF77Q9IM6bxtKfGRqnrYc+qsLCuEpmA1Y0cZ/0HT9m7SVJeIWtrrfM69gy1lM+Q
ARbsB+WpIsQcegJzTLZ0AkKRMNXct4JgJp/6YWwnU1KqThnRLcIV0w8Jtx2CuM60qWawLkLHQQnG
Ryrze+AjMvhAb5BNKiUsq2OukmcDFcAzijKfM5jpmOaSsFuFc0cvvMm41t1w7E78DpuOkLcpjAWg
k0T0GpNrn+eHbmZl0RCLB5XzEvyFg11dIo76BGoJvJUcjs/d9DeOTIpKEus1LozHkozjcTWdIJLf
nV8doe3prcbkuQKEI4JsXI9V08ameqA8DsTo9VPcmcE+JjPfXbhnWDYNciJrSv1i8SSKAQs+GB8/
jvy7m8Lojz0ZWvTMK+Bt7x6NKa/Q2lgGt2R4O1yBPnyaztdBqsOJwdY7ET0RHsD+559q7u0o4wNQ
fgzQWtLD57KqHV7LqdWOXS/bdCSslMpQh7yZHmnJIqkMVZrZfo5yThzEUr09/ELSc8VIt2Ctjlt1
C1ZSMjgxv251IjZ/Dw3FzptMSeCWQgZfdp0WtEgBh+7C5iW14DElRTFTbZ/GRxrL44kps4ig0sp4
Sh6eJxC3Oj7mNGRn9vN6BboxXgDBHb4ABMPFBr0Ff/3ktmT56ViUUrPr5EmxGIYwBstaXcxMgPL9
UZYbjCM1ue0gIQXwEHWumKwNcgv/b5LnNQi8vJXRaH49fcZ0k3IXIXH9HJhqLoN/NKxInYbJrJGc
PGEQBtH1kSWXC93TV+YbXDod4nL544N/eg2deAOgND5R9MzrRRhuogg4EHyHswV0jlv1OIXqV9ya
CUJodo3bj+PpkneYEGiLR//kOO6wU2az8YYFbhEEf7LNdi1wthtZa3JR3W0xqdpLO9uwuyq+vMAz
wGJCrxAi9v2IFRcWKfWgH12seKWgkXcWSOO9Nj8EqxoRy/Ds28816+v4ybRK3UykQgbY1EJmxd7p
b2Ps3GYMSAkqbPL0IwgulXqlSxOciwwT53HHIt3gLu6G1wENLEFfT2b8zetrWfqjsy83e/WKjG0c
CcfD4K7IXKo+NYuwAEZ2WJhDI+OlQ4HdiY2EeauVzuhMRcNYhHPpyF3YP+qD0Hhr/BB/4zrCACvz
ycmn10v3VFg1SwymSd8luH+/q59+2Ik9JA7Ksle7nKaPXJLXJ1tnDKcRokianEprQ+Duhv9cLSXa
a/vt19vQkHL990gVRbXfxC3y7oEl4ksLDGqLtmCMZpAPxP3p/Sb1jkB+qCWud62B3MIcuYbqSiUd
MwZd2vpN/wrGRmQ/tpNG8brkMX2rj6hh9I71kbxeYe1JjN7Hs5vDrkN8L9StayMHuZ9w3rZcl2xT
5XuPjev0qV/3/jdrJBMwYsfndW+BtprJzmSVu9ZqpWtz66lAHpjrUvhzF9IkJpIPOYZoH3eILNWC
s+PijfjQdebPVKn7QuiRJkVfV55RFKmmqRP79Gt8dYz1zhh68nHEP4Jz7TKK962Z3tTJcYezHqWr
wDC9mo3wc1EaQ6OI1VnwzWDIqj0z8nF5En/sSuLTwMoaqHCnzsQvsyRJPwR4tKRGSRr2AfG0BMTA
WwXUZpDnwileoXIsDOSz7WShRxpjyAbhvShomM8LCYCZSkcAXpCUrE5UUzyfoUXh2sPDOBeIz4kq
jdmBZxqMT3v/m1CcSq/0xpnSIJ1IxMjftEgmRAAdk3nC/mHqrGvL+OCHjShfdQktc69KE1J5PvH0
nIZne29vluFmQoIZGp2n+HUe8rov2JHr/N2o6VxywBurxC+hKEsrBoR3Tp66bThf8Yz4mBTCjX7c
E09nxG7rjP3aW//lRu2bo/60xFgh/Scm6zG2Ag2lrGWhEqlVjSkdVxzfoCyBS1/Ra/XzmT6i5Ece
4BDZ9mJtgi1ffp4NOy9geXctBR5+DE1yA8pBg2EGT3BoWL5EhQtIqDj5bM24oPF9n3zUO2aaamSI
dXzgqZetmOFMXYsztTolcqq7dOVKyI9wVKoDTu3ZV3UE87UeudiuBItVgm/bIej0TYT8psXxZ2xp
ZNLErlVvICpFym872VY8KiLlykBN87CoFU+kMs4l/Ogkg1MTxiqVCBef11ex0dEyGORnNlqzcxaC
glEn8gkr2S42ZzIPiJtBbq4MjZVdCVnh1wvQLYAtTomQVy2ZpKdiW1KhTWiEz5Cf666pkIoVRPuR
R36HkG1BxlZ0k+Ahx05JU6dNOX7I3PqpQtovdSi7vvDcMK3xTnz8V81DWDCWmdRpai7A3ePCByxK
URXHUWvPqNIuLjdRAdTK9nRs3eRac9bor+wyP+GKM8vcibtkT2wHaX6gEiR2wHA7eVA2H9tQgRq6
JKorO82Sq4nRL+9wDGdPynBaTyH7tx0Gm1YBc8E71TFUNiPeXXNbC2tAhVZ5FjtLS1YvIBFA3ERV
mytV1FtrEVvLgkEnUuoyU4hOCHT5ESrW1tPZMIM1MJ6cNmZkSZj6NkwFFzirPpD3GyiJlOfIyjdu
UXu89RWBU+loAKXKdhb+p9e1sk0MdzNBqoSuXQnFl8EV0unkDNiZ3K1dnUZYWYNdzPKawohqIKq3
QcW7+EMaCQFIjyGPvsRdDoSWwgUrZSSQaj6JybtFKbgbZY7o602vuJRHWqrItNzb+3D7tnG2+/O/
MhkDFMJvW2HGOKNkClKxeALZ8OpH8oB6dffObyUKaVIjtHQyfDWgpdycIa/anKd/JCis2mqKRX2i
XtRmo0jxvAcIMpE2NiHZaO0/XVrBHnHJ8hZdiz4AMG2Gf2uLY9SxdSMR1FWKUNmwhQisRbSKbC6C
Ia9M+2vyyyio0jXA1VCki4GKytV+Fed5YcGTjV6plHiVkZcmkse+OEGwJ1rdwknhrznxkm8QJOqJ
k/xG6WFX4OPG7yUYbL+O4llgFq84GTu2mZ4Y5TYBG1oQcgvnq0C+n4Hm/yJsIWDuBpbx4aJw2sgW
MUuDFf3AQEafoERAnGRO4relxxOjhHf/UoBRQJjL2kMH7YSrVeyRgB6XxXASr8eE4uQaIaYyqIpq
KVAoN2hXKrtCW3r13MQ+DLl5Rk92aSH0r8AxpZL+dbJjun2TFlHiuaYQx0TAiLEb6zgGt53eA60s
MeoNBKu+brH+xOD6jz6UZ3U6gIpfuaMpOYsqJ8i5SYYpxqnavdAT/U3b9ABjvJZT1XK7V10fu3P7
0ItVkhvF/MFT5thjjhex8V8dybv9vUv+OTCBp1LzO8kutD5C4N1YHcSVCGkGi1+BI48gsXKOFI6k
hSbL6JCy5jnuy/Jx+GPTEr6ui8AJrgPJY7Yv+B2x3cd5gnpQmvK8Y73VQDHE/K7AEt1AypDUMlhn
kj1CAwS7WnlOpXGpL8H5a06yWoXe4iqz+yDvDNKRH1d1/Ss9xp34sqna6jL/JswxO87A4Q8eNKQc
TXzNF3X7+dIVSrUy6sFGqJ5KNsst0Tz1LprjJce4J3c9e4kBTHncjl/Nfin3gANl6jWamvK7GmGj
H05qDw2x/O30YDODQqjOf21u1h5K2s6xBjwP5u3NhKY7GVUMI6F8AQaKfGde87ToyUl22MbjPaDa
mVIIEiw1Zp20/Fne2+2DPFe5C1AlQJOAqXwuXjuVqLWxrFQgclyPh2PSpcUc3ZAa3Z2M3zsC0vzA
1ie8DgWxUtbr2mCkdX2iqtuFAf2TkLQ71+kP4ljE22IPJ55OtaefcqBKml4qctaj1AZfxXWjJhM7
xfO3te5rt9F7Pir0MdqPL2qTVht8O1NwEF1qHDIc0KcfFwiuJWO6hnFWfoTKnbcJdF2RUuXkRsfD
2Cjbq0PAHlJrXhp5YHWExEdqUc7JxexYrp60zO/FCP0XJDSuRKziZxgH1cBt7CotgUdDgNilEzYR
lyicsJlnhPBVdNpmUCfXdfouSa2OCpTF70H/pyINoFar9i76/WIbxzV/k8/rjD1o4Wsx8o5SaBOt
+JuUMztN47HuDTwFBDMhIExPkK+mSeGWM72a/ZRol51D4IjTKe+v/ejMxB8TvNq5jNE0uBmguOen
B6VK2Wz9QZ4vnhPUgpbwKNfCVLGv5BF8JfJoO1XA1RWuSJkc91wYNdtJfM7QockMuHLZJjaQ3Fks
jx5XgeT38smDGR1Djrtc0W8+ovcWL4VbXr9OVsqhl3yMHN7G+AptCEb+pcuMdhLuOrNnofrsHevF
CN44hT1jLAwbtXUkSAqgsC2Bg+CFeDrRTYlm1tkaaXKwb4ii7uIlJEOEz4gIZ4lL4DOgzUV+UWUS
vs5sguqr3utJqHlKmEbl3vL0NHBkKehDl3+kcXWVizXSUxmpbuY/bMuCfjrldJ28dPsFqJoVoWlu
i8wcC8nj3HytmVJl21kZT8ftpXEY2+Vp1jk5BbggRODllCKgBOOUJIzFLWoG2ocikc1ANeljYM79
FTj3rhc7nohSLDB45+6zOsKMwSsDFZSxxITr39XXGyXUL2BRxD56+gxQBywuYP7xYdh7sK4NJJ1M
7kN13mXYw4TyyC/CQ4rvAyScCKCJq72xhWNVlT+MMtNk7K5QNScNYVa+3k43/rtSm6u4SpD2vI+1
LUJjhXI3wfYEAKGw2XKvT+c9s61dwzKp40towiScPG63bPcckdw6vL4/0cJPSIKFuP6Pboby0z16
Gs5hWIqYozE31Mr9jEXf1gzhSFyoW95WFSZXlGAoHB+kzln1CWOHpJt0MeNa315qw486tMqus85f
f2hVzsxLDgMaMQbTF30qHgc6IBXblvD94qbTtwkMey2whnHjtfNcx5Kh7AlRi695bkbYYUsihHgW
ZVRrk4CY1tQyNJTMxSP7087SnzBQNRF9RNlLQOAnmFmVyRchXTPxZ2pyekiTplOuVOhhFOibSUfV
b1irMbNRFiVeJSg+w6kCGX+WuPApLhRyzT2VnQ/566kfuNPXGlaT+mMoEpgz9nJRjyfClcykh+v2
Fj1n395USlIVLUmwRM/KLMmu8zNOOEDyAylFLuPCbeGy8/gCvIrcIFm6XjohyKM2+o/0ECbwjVrB
qEsG8mKXesdeOf/5a6iufvtieerRjIbJsU+ajDnL2Z8Qaj9I5NxMhBX35ViVy0ifFc3GQ0u2DukD
UbBIa746/2Ge/ib1y4S38TJKnXUsY3v31tA6XV5tMaZIY2Dx5ZB7T9nC8mNnLfgRfUF7n12WBKvl
ajMs679J6IrQ/CLZ7bNh1x1QTPccN+v541xOP0Ib+MX0q/LpUGWx52h+2KhCkvgF1CyoqsiX8pPB
FcoS5tswcVCTh7UT9ZUJK6dpPhtdDfXpN+9AWkJAQCd1NNSfJ9KblyGS5vulagBBi3UY7/DTIEff
Ot29xOGiDmpHU+xXCg4zzJO0aZLQV4fyJb/eNRaAhDeplBOTkHHdNgSrqq2VhIEAp3l4F363LtUo
8KEqA37hdlQjMpFoG/KFeiWmhX2ifduTSrUXMdiMQGjUOAXZEr7a0/HP5MHAe1zlbBPyB+9zMKDz
togZdC0vQgIJ8CI7ClExNxgxLMv5yllE0C9uwbK77rR6TeloG5+u4UsaNLq9Q8uAMP0Sn7zi7vAy
qBi04MIQiZW+8zhegxFc0/voBNEI0uCcrhlcLnMX5rrry1DDd5Xc4a4UwYthxH62d6IOIV3Q5kRr
SAYdK2/gryYv0r63MldFSQXH3uzjbol/70CBUBS/UGuvKEPA4KtbehyyqmDH+To33Ue3PtJ8SGIC
SYYQa7nB4eUESSdHIFmrirmAO0wRTYclB3ixBvgPNSeDx7Z8cCS/PY2EPOruBeIpTaB12cjSmVhb
ClK1FwiLP/Gv8vdmUdPbJ3l3fkg1S6lDMScm5sXOgK9ARYNBn0lZj4PZAgCVEZ5mt3kn4qIs/4Fc
xvwnwgRwKNUKpZ4DOv8UJ/M9cKXD7S3wgmboPQ4ZJqy4qqFoiiIwWavop7Fzg4shFranKuY87154
eFEfWiFDQrduUb9mijjEHaMHyHljO1poQaJPBpui7iqOhyKDirSdytRLRx+qqg8DvXs/woAAW2/f
g7zIE4sxP9z93kba1f0ex8QqRKxd5yGCsn5UW3JXI9PBJWX62rFFxC0QfZO6w9YYc/x5MtXNanpF
Qe00/gFofonh+iUSF0nF3mMRsLK5TJilvQOP+Mg8ofFeiRIzocKznQCsBBNPiknFT/wjBdbIpVdg
x/iqIr4P6tA+xzhTgRXU8//rh+rzqemLbpg7IljzoP4h5KouR2nQFViJOBY4Tw2/xpoaY1Rhhis8
MVBgP8X3A+ChuEcB4/sHwa9AqLq58FfkWxD96TgvfvI/7tP/J8qd4uJWJTEg84FaG5SM04LfudzL
cApSYdLUluzT8Yhwy+Hpno+SYqkhMYSA2D6LgeNXDcQWSMdWO5Kqv87MUkgo7neyXLtpE/zB6V/p
oucF1h86qcM6bp+KmmD6nYAEyt3wH1PsZA4TRDmNhiz36I2H47tf2No0Aab4pA7ZowbDwWdsBRxT
tQwlnXcTNYx28j5eowr4RBnCoRGTB5+6iUYOjhw/TT3WOvgrAKWvPU/sbaFCQNGq6JAeMc/Neqlc
r6Rci98ujJOtd/Z8+GZ/CbPFp4pohDYm+/VRw9wCHz37gN8jQI2RTyFfI59dY4DgKBf+Fh8j1rdn
PbcbskHI1rXa0tt9dGOVGxONUwN+HZNktITityOIFOvEYACAYQawOMZJx1QKw27aP5YQlNHzicUS
ZbfI022BCcw1rrDubprMuy7SXMQXdNfyuO2IEL2zQg5rfPlcgwjRP00LWjattF2ZV9TW5VKwHzq2
kxDaNBnPKrMenVbuTZTZdO/1sZ4RQhpvUeymHE/73NR6g6k+UUWUcvG9t6iRTJBe0Me5SKmW4roC
u4Tzmv8y9E5Fduxu111LU+laLr+pW0tFEYU4JUjTtJXw50ZargdDVyujZTZG5r1AYZ4QAydtuc56
MxueHye0BelwkaGrsmpu1b3l3L4bsLfKMZaJwG2i+hkjLQvylk2+AKYIJPjYKCiuL4de4srzu3Ym
t3gBsbV5/xZTP+TxzXrOSlZO2416J2ziviEq49VIVQZMLyB4DCvdwGbcqCK/V/m7WkfO7e5pAFGw
VApzZBgGkNdKi4lV5PkVuHILLH1Fd6Ts2RCK39D6xI3D3J/0ljNB2l3+s18XfzlRfwySqIaVdtIw
aNjqshR3EqXd7SJAl0M1T116S4zzH+Lbr8/qsG1b0GpfvQjLzB5qwiRF4bDUSSQvmjFTdFHJ6OWm
Z4jYTKDCcYU1rWXhp69ZiYbsPltpqFa1MS2HZ8PTaEWHSyx3rwzqJCzEEWDVJFuuysrHp9SY0q9I
fCrWetoewrg8WxvE+adK9GH7nuVhAHjIjX7NYHj54DLJGqPGks18tp0jjisigNmkzNJ+KsrF/3YW
Q1cTfPdLX4xYcZB6RkHxkc5HqaDzAsS7uY5DAJmEyO0oa2hkCgNxU8R3s9LJD/p/nQ/BRjX0F78t
27FdnfXPcM4RdOhtVBd/AsZHHSv5HmKngcG7QRLjqks9TaTD10YKIEel33SlR5oBLFCv70gnK8/T
lQCQYJbvoEKRYUPjAlIm0pFi/5WOD6521JHjvCUa9ozhn4Vy7dMUySCeRnTbRqE+9XB8BfHoO9Ue
9wpMfrk/m5eS0BUNBJ5TOTIgxztthbGkVe3mlCCGDtrJVq50p3SdXwiPxbFT5NGfepyCUXodc8Pj
xFlnHB68QJyhce7dI3OYkVxA7lF9T2HGraC+1wwI8FlywrdRcWhbpfSQOwFepKY8uUL+1NVPjc1F
zfu7L26ADFWODc0qZQJVZWP82xfjOdDu3F0RdgoDcxHz6s9e4Yty+iXcpcwTD2npD3Y3ukOhllPb
oZP4F6LIIr1C/v+PqzL7HPNrMmx5QwRiuMi4mv+r0/57H4ANOYkvQCx5TYguTqgUEDuJi0hs4atK
x4Z4VM3Dd1AengkYqmmyxQU9RGJ10wIa+v7A6BzpNwSaUjLZNL34rrGRwXungDF/fvKQt4P6qEDl
TgADaBPG5FG2dCH33SXSjWsGsTFVTbQT8f7YuErFk5fqHhlkdjdPYHvOnrgmw7A1ujbj5H6NzpXH
K/3++8vDScqwo2v0OF+TlztenMPP0pxMqrqyB+9Lxt8uJV+LceLJkjk5o0g2t6w9qfvhJ4hkPXGd
rn5c9JGOqJkJyb4AikuchEaoMv/N/+p+gqLDtOvI5mh2uXzDZ5OXS1NXDxH+qgRltM9lZ5LRbh//
VayYW4ppjngpSJ8pXLiH0cCSLi9An5unLH69kqbC0VJAb/EwtR8DytszY6ZJmrbM2CybdTDJt5NP
nQj11AMzFYdg0skKg7/tSqIbjeR/53Nc7cQDXLoggRZMH7mI/TunRJARF/9Yth7jg58ipthRY+eS
pgxExagloYnl0WDNK4RaBew41If5m/zr6ZMGbZynzmYsztQjr/XyB3+fdwDmQ/NO9mwHEt5FmcEi
fGy5z8dJ+YcmWyKOfLqnXgPwzWyLlzganUKV3LSSXjNXRXyvdI5T51S+PK4Xx5ca34rVNGFEH+uV
T+e/T/HrSRDwqqk/WvVXGZ+5w25SCXcK8vmtuncy6VEw8VXy0wYJFAvuSh/M/z6kGFG38ZQeUnpu
IUNzz4+H7uefJmIcERb8CYcm37V0VunZqRjwzitKX+i6o69RpKvUHEYANEjty24Vo5bWjoinhBeP
uMB5gizq7VinpK6ot1md+bPmaqE9sPetS7UtoXYYrylB9Do2U813d/YsSV5Wyzz4huwOi1IbYho1
ZVGCLUGFnvePcCKwtffEHxVCTeGG0174fzbCComwpxPUsS9JLU5hPCCs5UqCFxUy4zfYAg7Xx618
r86PDKaO/GoXRG/50udQacQjJb30Jl9O6pQ5Y7xzASA9jc0kIu35feMI4ITYqSEwQMkoG+K+nyaq
EylY6yuj1SIHLTnEkUxwPhfQcWMx5n2Jn/CGCfEVG17ZuBAwi1OQNGg1rt28XvT1RIGsuDhGS8uM
yCMrGRo/rV1PUjFzfAkj8owzdUZCeCgap4UZc0YfQfJ1GR1+XWe8GbwUMEYhLGYhAXXYBhX/b5nd
nm97H/LL5m5of78wZWxW/LHJJYfh7NO9t6Bk4VrH+QcA4R9kObOJjMKMvJPPmtKpMmOKsp2cV9Dq
IM4NIs9Glp68YoufJX3TtwIWFY2s7+jYCfYgNrWRiX8jmx9pQ29uLxByqz/N+wysvUzcJolPNNTH
+E7H8Yk2ZIglQNIj+qFpTizaeI4pFm440a1gXNF95OWKFQpSR8qNFSjvg/JjfgkVm40X+LNaliHl
kyS2dKFRbp4ghLoUnRz75Pjf03XUuIFX3Wa7PBIffbqJangq5zCBQu/lXoVtHaEi4EQXyfDuM3IY
wKHv+Z/B3hXhJU8LkRY6kOxv9S3bhpEl1Z7OBmKXLJ4YeRDPBJUS3lzEwI/bURA66eljflXaq80S
USknr88WtsyqYef60JeVxt1ZZXjYuqz9Ttn/VfALh9b+2QxjY8gAwrEiWF36qpa197gb/2FbeqBB
SqenqRqxq2m9/xWuftvELnQrz2ZqDiEeFKdu+lTKOnsFSq+8K5xd07WJXeq1zAmL0l1zl+qdr5kr
545WjRwMCOR+/3MUlRrI3Q0ugG4rFsJrNbq85sI5rRK/+o2HYedsrG8YVfxmxaGsQYSAMrOYNtMa
94p0G/aPDY7MYquc7HYs76UqLqsC2nyFhij4se+8rsEBf9lirDYP92xHnWnR9GPgr7+dYbm+TpCb
vT+o1KjCnEibQrXmfrcFELmn7nSzi2sp36lRt8JVdviR6OUItsWLzZyeNsrPT6ZqegJpPc0xZZMF
fOUZvX17Vec9iz8mz2hKeNENvfgLr/gAYuFjg1cmvupMg3Es5YPgj8TooqHnN4EdxLU+eUwvDSk9
v21IkXGwTBQAZqaALn9s10S5okuwprWLfFSgntjWkbSeyKwMhjtj3NEQP1a/kBVj67v+pCmXIuNi
G9DVtxylKJQ3xyywPhnBRJdMgHDGTSNIKtymwq1PiP+OU5QD4M1Xt9F1nXb6FRQdkEbMmDxf4x4X
RczTyZ3AzmZ+tz3mCu/CD0dmeZ/tOT3uGjZntKWBDe7ZGlwQSKCulyRhcFVxeLeVoy4AZwe8hIBL
/yC1UN3sRc0pmD+d8P6Ns8UdNEY+jnWz92mZU99qSqMDD0wjRpfBsL+SOIEHnPCG9n+dijfojhoq
v0qfvV6ouxoXyblH2tV7TiHd/WD7f906ytCjjftx7ujP9edhFF/9BzcuTh878LOXxx4kqLm4bGZn
nbaaK5LH1ZqTa/biMG5z3srIFUtPCU3sqpGGDdFj7wD9F384Rms2r+Ctxw0b/+kT2Y20VGbZqp2R
CdVf7gT/3RwwsiTVlA0BtJSPmPp8DEo9WaI/+ZdBTZ2d1Q8Arktptiu2t28vEnJHJLzi4ID1YA6Y
fbQBQXr3siqj7nyU20SboqE2PPQvo8mMg2DEJP0qFsGTy49VVFXsr6zub61pFvciXHZxGTScAKt8
Er4Pbk1wHrTaUgTvFRa7tr5KYQAT54EDnTWX2Y7yAupekGGbkYQoojasBHrsfvMIuGpQoeNKnANW
7zWFjyE6ZaiS8NNmzbes+QG56RwD36zjNl0gYl48gehcgFwHqEEDlUdb2FDeC1B89STGkWzZ03nK
ZIqLQw4ZmsQLM8QlQPDuMzCjlfJj0Q2Prf37/ejBjx1aGOasiww4UVPGZnDBb8RIgFW/Bp7tsP3a
FkXLg2G1WQHxrMavZxM0QHMziU7wWmf0SDF9RDatcJxB4C1yk/u/nhopz74bnATfu0ut+17UAyCQ
4HjJQmHR6QJLzxjcV+aqqxP1fgBssRTCqaGquBN//9Mh2X5oDuo0Gkrky8UP1zLsyMb3amzWiLtu
KAZ5ww0VCu8L4jrRf0muCp5RVOSJNuGqyf7L9oGPY1eNcHNa44gPpBwV1Js1Y2+78MEpKpZjRqIB
E6U89bwoI1L4rVyE6IvRLEZKL+rSMzpTCaAfFgpbsFC99u9qNSy7Fdxva7BkvR//Ehom/c/oFzyD
Evr/9af6QXT/rlz+hD+ii4MLID4W0Rfl9Vn9A4sFbAd4USGiGCYlUKuRTDYs643pFx0IwjX5EBEc
OPkWGTpQ1TLwU337wRIxwzSn+JAyPnjzckKrg/Ukmt7iCKyl8qiinOv6OVLOUhy+brpm3gAJLKWH
ktozhkqZmowE/WbyiukSowtuWkAdRrNaF0O8lWpmBKVXvKhw8tfLCsivWAmEVNSUtR9KkIBQ3rt2
pWbwt0vQ+gJcJIy9h9lbR4osysR7KRxAG+AGa8XXg80CViM1mmwMCsFhQ49T6z/wCQ6he4kzxBBi
/7M9F4zAOsWHyUgpGgMq1jWDa00NTFfoxsBBRJcdghxGSOQMK3RJbFJpSMyNxuLXSZx84nqQX9kg
5AtfODiFNBo2jVD0m5oO8OriVdfl7O9fxkdX+xv5s/avBk/UUeaFv/rRnM07UH7/nk1kDVJUSviW
6ZpsxbuhG5hnFgqVTGA9KfVTMbsoTe8Y94pYprG4ubD0w5gmKP9uM0BiwnaWSRK/9xAy/xbwZcEu
25d3aBkOTZ6zx64uyvfqZoOv1xe92ksPhFbc/KKa4hJcAdWBViZfzNp4yMu7PQYZZ/OBdeSXiU6O
1OmIcXA14a+Xozhil9/BXzEkF2iTAAND1Tk3Q1dmdCvRat37g+ROu9iTq4bkLIbQnDzdQuuUbJnK
Dfw1CzY/KpXws8RiJM1Xn47pwxMy4yZHZ8sM4Iz01IoYhVonoDbbxcXprLmr2rREDTfVFL9d9L/o
KKgxZ9pkt04j5GkuWzZpFHaPHhlqHf85BqH0Bqg94vkVZHJevIscVEeR11loLCtJLCzNlCUevYDw
Tun0YIQ4b1fdrbji5U6X5Al6dcbaYakt8YRRjnQQGOGkrR9Zk/AcU7w0EoooJMzno6g8neWs8CUN
IVznvD0e1hkeSBiBV7ccxMBgL7RaAJjP3JcUXCicT/ATFUddhPFGals7HB7hst3KKIRSOhDXLkJH
qlRPHkBvuqBNjcru9UBFsakWIHurAos7iFonuT8j+DXryCfZMYujVT+jf8+TIMBNeq4Gig5WnpJD
G15bzHZBg5baeOYhXLfj2P8RLu72+zT5MB4u+9jT1AVQNtZc2gOvBZSzRwZGqze9+bPBDJ6lmznV
m3z8LS2lOKbxxm81Rs2qgZ372Ptgir5KVEvPcyRcF5BIxc0T69mNRz5qRkxzkV4+TWUMiGVTCuLb
ES6AlHvEwxQc31eiLQfV0PpeC9ZvIa2pIreEiqZ8Iz5WeTR+aSY66sVGSUZG2jemzGDskIvJ/zgT
Sd9tAmsbk4C684or2iqR7UGSUBMklL3F2f+N6jYd4kihr8/qO+mH5VgTLjp85C6UnQcoVmDeTqFO
itbDL+eiX7RM9tutGWaXNbartczyV/ICNSaNt7k0oJy6fm0VgNEEXnjno1CS8UQ26qFWFUIG+hWq
VYOuL9LOInSZJlpeWahVDh452aNRuqxsKGro0yGScCRndkgO1lbiXxtga4/lc78BQd1/glFQzVc1
BOL0q+EYV3jUdirF+UolgWtXrUdwbKY6iBlRRb79Yt9BtGMf+A7xb9BVQH2noVPW2AzJ9804tl5H
Ce19J9KFL2v9i2JwO2ZN34GUOan0BCGormPQAro9IWRl059l3sn1feYoFwjrysJLDCQ+g7qh0O34
IqFrb561Gg1i5ARVIh815f00yhMfo9cys22SdL4eOP1mnep1G1EerB/Rauq1GZqukcQBL5lKXGmy
0yfZBTr2ckmG9IvaRmHxP4lW+jsksFP/3dNVDVas3cXcDXCLMYfZJkYIV6J9XpPt8P8kGNGJ0mUA
QkPJkTvyNMVlfq//ZlmaykPmiKg1GsPMC/1OegIlYTkEK6EzBVoa0tlgkcDBsI8s+l1qve7KYdKa
TgsVN3/MR5urmtwfKtI35De3cGAV0U+yRnntPnMoMZZZVHBlt4LxUKR85bGK1if0e6QJNwUlufzU
pJUP6t6YWODKCxnCn77hzIzDO7rnoAfS9quhvmVsIk40TZ+fFiLK5OV1HU+buU0RSpt+T5wryM+D
JeQBuoPvKiKLo8vLTkkF1wMp5UEONWRYm7OwSAxcJ08PHg5XF0LK9BJraNQCQkcZkWhpk8r2Le6a
Zbswvr2MA+mEwA01epUgsjAewTKBWpV82mqeMrEKwuZhXHmV9Z5PdTxGOp5xXYcjSf35Ris9G0eu
x4DhkyzQuj2ovV8zgwXNhOa4KfwWRg5qthPK1vw1wZXBm0Wv+GASIMxqN7XXx49GrEoS7l1H/9j1
o7NpUtK9/e40Ic2QQLXL78FTIjs89mEnAD3Al9dMrWGOjRVcB88knFXdtcLnA2WFpQLJ06ohdKQ4
ukKCPqAIlk+QwO+JcpZnixEVbw4Cee87DjbJux7ByL1/7p5xVQHCoHkT7hHxQYEZHHLQmlqIbIyV
z7CzKHXW3hU/Yn6PJNo90FTB2NOaIjYDwQz11AwzA+pU7eD0LMRNTKnFsB42M7fPelxDMWQjtkGv
wLfiPw66mKnNuNf/hsEhguQPZPiclUVDtopR0gfxHqKTeTObSkaYkDLx9m6HuGcKfWA1qG1rnmdh
UFOUfZJWk1e/Rf4RDryrD7jOJqXhzy0qXTxgFcF8GMXq+Mm8i/U7svtcMeOtFTvEmpqYJ9o6M6Xw
wlVMdzOkGkK3lcONXuS2BgPFR1On8GTspiMrWrvp8wn9KXXx3wGWx3kFTzJt1vcdsqTGsRuYE73h
WcWm8EPswhcmc+XBS0YDI7bQqQd9NfO5wvyflAbMhbwoZSiajarv0liRhEqVF22rTBWrVD8Bsri4
TktZUYXbqKHR4tYDh9jVX1iEBxl+I/LKuzZ5M8LWBFAaIxuCj5kxe9FWvx4aNEPakord4rjDLChg
mKUVU2Au4Qk6oCBLHAd0TeK5s6KRv9Bo96DluF2ui6geTEBRwQsQk/bARFEBVrVqezCdQoUtRsfQ
MxseiG9P7EUsr+ZT3DQU/ZCBu/7dTLwhYDQnWv4xMRJ6dKkzPdnS6smanQzY/AiStm87EBM7MthC
ZkCSglXIHGVWlprvKLJ8Z0s80f4hCN6+Q4x+JVobGHg+d3P3TDRen6mDu8pynvsVUYvzlanH76wr
HHJ077LUTzNd9sQqTY0SAGYpeqFuzYf0kJKw3u3k9GOcT1vqvGZmfJrqTDucjXaYtl8Hv18blGpR
FlM5/gn1Zlj37XXp+fJvB+OkkayfRUvkyXRRPGmB3dfFaPbEd6DLTOyoTrMEHqbKT70Gbt3hoWBz
MVoyScXGa78Qjw4/J6imklrlY2p28heXV5d6H6D6g0VuVZesRRwJ/AEulw0SeJECSPpm2opxhkn5
YWI440v9+oZaGVqiKMDPbZqaZvXz1BhdtkjG4vd2wPIHZvwOHQHs2HXTew9F5wCJqcffLcSSBllX
tMYB53Px1DndCOYGu+iT20o8VprDn4Ctq4aOSesC99cXQC8zutFa0ms80469jJ5Lw2odTBBM++QF
sBHBGiqsriNvsyGo17hwcheCVAW077hsAuQffjhz+RAx6O6z4M4RrMHVe54pGE9LkSz1rfv4c7vV
KgxTo++PlQx1drdKNiqYAoVD7yyqN58wQ0oKXtNZ9mxuC6h9r0/zvWMZKq4XNNZYD86F20ZSe3O9
KH1Ei6ayctXBbr97aCfrM6jm5tAz80E0aDtmDEw4YCCpfZGzrCRHTADVEoD0MzXe9hBE9L5QchRd
cdHvRDo1LJCv87TB+txqBDN9CuMN8ix9PkXxGHkZhiO+qZvBtad81dLU3jzDCbMcF9xXasqTm2eH
qbDQKsoJhZEi0KhrDwxZl00tmJY3apc5+IoFxYvVRUXyIMssLNUpbEyFHKdIxV4267+LmgB5asQc
xkqXMl7cF1DnCmiY5Qu9Nyzyii6WVdPvJC4WM1gf6yeHsjBcxcqP+w7Nwd5D+1tV/NwJSyHDGkTP
hMBUb93XIZZS8rUtQty8P6xr+yt8XhmhQNjOPaCRmf7Igcz2xdE0oD4tDllhAxpQ+bZNP40rbHtW
17Cej/24CQ/dU+306d7gZ0Fze6iQ+5bSKTf6jDO8zASReo3VNZLR5DezcYVexOBS0xlkQx9BqH2f
/2k7UxGGEhoVfl24sm0c9KP2fKhHP0d/rcVJmbyKwDUa3kXDpOc8Q4rzEW2Gde07hOtw5MWPDT49
sXjmoZaxQFwT8DTwmyiLRA2Tw31byzCIOOmk2g9tGp/CtNnATseq5PThMHuUTn/yzIzwvJdqnkRr
zmwdcy4D6B+vJLQppAwQQtvx3OSFuuUsIEO121SaT9roqjBB6+3UzbjjfIXnsxa9FnAY4Z4QHHqR
B21HFqN8jj9mlCy76LOvSKJgwwvyK7Hc/cpS0MEB27Bv2wqZ+hVc311gHHg5ewJ32gCCSR9Iy4JZ
XJhBfZslkYTyR/bu22mQnB7E78NP4c5BSo5kQKJq9P1wRk7QAa8biiQpsi/eSKnzQlvlViXUJ//I
cQvwcYld1cSaq1POREeVb/Kamm+Fz721yoR9oTnfeDn++7CWuQS5WutJHX+7OKmHaHJvZEnbePfN
duuQHnH8hDNF8bDit81EA4sJQtwEc1Ttt/sr3g+yO1Li1j+/3WEkphi9aFj0yNVybQjHXYTENV/w
7ffMbZhDPbRkdetuXIDtu51RA1bh+z6DiGED3aXhguQMSXp1EuDtntZcjivQILScM0mzk7jFKxBi
7kwCg4Dd/2bqgJBUPb1xTUhCIUNTC/PgavU9K/SPPN1V8v9i2o1bjSd4Us7UE14R/aDDrZhkhSDz
ojKhjKgBrWRC6B0HlyRE2nxYKkALf/WXQuAlfMIyLWfacY4bElarBlJdnmnSAuIRX6IWsMwHNwGK
5kj5+tj1xC1KIQJJ7L9OHTVxx4H1ePvsq3M48yFG59gCBe3O6NsfRP/fl1uGUdsVmP44s6NaUAlx
k+CWcME6YIMS9RkR0s8EmukzySrAlUlfGPbt2EOmRN1a1nelOc5AFF74MjHFGy36ZzUfUvligSwj
2Zhw/UMXFpVgbm6TXiHS3Zg6mlsS2haJ7EZYZZ0UYSsBLQt3vOOdh5yOvYmYBcEMKjnWFmkMmKYh
jlZ2/Ootj0hyLVAz/8DYhogvJ/SHJ8XgQria+2DL+BFiffoqxn7nGsbYG6QIFJo0kQMxb3fNT0/9
KYB+ePvoiHhMjmss7Pe/7E1eRnxcjeoEbv0aNdMlFQ43R+aXExLgUdlyU8bvMTL+18dT0YhZn4ip
T4OGbNkRMsnW1zAvA1PHhoSgHaGCzRVaoE8+goQnILqP/7KSFaTqzWWuvKXHlLuhZr5Yqz6N5+EC
tJab/uM3Hm90H5TJa2WzVG/nfc5NlGIaod38kxvNvkBs3uZ70TLxip4PRbqf1yvQZTeS7fFWAK2W
IlTXAkxaUtYapjnm5NMSQ0A6EcpiQtOCJyvASXyNuHRBPoROgRgt3WUibnFujZWdDBaOQZP5aIS9
F5Zuaz4bWj977RK9IJNORkM/wjFqqF/0OMxo7SOkbg2gYNWJbtJ2xRFI3Mt/YN4qGfZUrxwYtdds
hJTimsFHviizZwtWpXGIFXQWIIjuv7Pl2esCl0/lY7ceaHTgiQNvl4iGI1VVyY0V19cLetQhKgFi
ImjKSFaMwqZ0TIH+y920p/9gqrAnIdDWP1ZJao1xRh3PJ+cZn3O5FM2AVmnXaAW7XxLr0FHZlvN4
AtBzy6FmRYG3m5/O9PiMAoLCUCFsBThRjNYieKSEjShGHZ/IuR5Doqvdv5xQhfUXfkv2ZD6tw1us
fmbSiVjld770ejEm2MscdQjXeuyb0loOfrqpgDJpyqxn7crql4dao8M5X+K8YQq56Pr3lrQtY1MW
zqItzzE7VCmwTSoasuxwrHZVgNZI4L54Ji53S6B9CjcfHLlwXTSdqRXbT8xWnO+u9oor3fBn9M7W
EAX9BoFqcrp1zISxiFxtaCEKTJMADXTld0raYkFv8H7e6Rq8HObqbBAbILwF0ecRmx+N5X8VJ8Ka
LVXnf88heLW/g3iSrwJdrZbUJrIxvrNcL9VOAcbyT5imJfpYaXSLp25kogNtfkKDxlID5wq2ePgS
rTwsx1Fvv9hVb0UxHIH/sLK2teWSNVfcnYeQIBvjAuWVkeY0yhgZa1oJgVySwycjMjHnE62AZJFe
aFosVE/t4Px5q+hNnAHbGplM2G99aR1RKI1NAhQvKeBOFJnN1cAjqm1WcNhM8MQ8ZFSjJbronrgC
tVbQdTx5cFNvF6q8Pw6FSCzqkyMau8j4994aeRQbi/LrQAZNK9RD61LqKpt4kF/PdYwJCRTAR4ED
bb7waVLCETnb0JRiX2NOOv6xbsiADuSsUHqyEcXngr3oezKfkJnZxeKjztY9v01Lr7spQgKc6ay+
mIuRFkmcrsBqykFZzu34V6NoE1jdpvT5TOufIzOnNTompYTTvy16sxAZPgKHlCnYlvHEpR0+Uylp
RzdBBrgaOMTghF2laW1aGSWvo8EeWeEcOxalD3ynCoqFL08i/j0A4KkLvWxaqBNtoqgxRrPhcOtH
OAzLWtWz4RZbMqfx6jswGKDIkhbpQK3X+wu8jF+7Z/P3TkCDBsEasVROsQ0C/lksmR5Q8EVGelaI
NJDIFigVVEf4HUfdd4tA80VBC1dvxCwIFAAq07RLWg/NjgrKV5MPbjRRTiz4ad5Nl4okl0aZnT6D
orkNv+TyVDX/fw74YSozVqohIMvTmolss1PU/r9T7EGitBI/n6rn50ngpafBK/XZ674l5+0P+ls/
GY3KC37p+fghDfqkh5ObOE9rBqb8Vm820QO9zpAUpV2kL7H9c65URbDiTgLU3z44a10Dm61EsdRa
J9IppQvCV720kZs5ERKyP2c2UIp20gyqNnAsO8k8MdfshUSKT2A5IpfXhql2ulCFSNQ7Wl/6M5if
GdmI9L1eSWcYFgOG10miTuWzFR1KoOizVeSQSn4pzKZnlNio2j0Uw9wU0kclcLNKmf/MQGayqQU5
4OZYkqHUzRY3S5LJWgON8sZ3DHPrfaCsQu2/ZncrE0dq1C4INbsUpK6bBOvgjR0Rfjx8H0L8mhxf
cWxn/V01Hij6pc6C1Mk/0vg1FqCSKkI2UrWKComeMG4Jouv1SOWQ2kd/AlYvw51easxCM8YrtLJM
wIDDMXYiKRkVmBRWGZdjnVxT5W6Ed6ykMpl31REYg7Mfrbnz/7RvFldxnQm5OAGelzH+YZn2W/x9
EbNcDjy6+NX0Uhdr3nscoTyAbQuYu06oVM//MLQ7eT6UkLDuG4+EKmWO+hMvyWoqc/Mh4WrZBbmm
4pWYLDjn9/uyORQgvMgKsTljix8/cn4ABHInlPRpbuvfdZoUQMcI7tuqE2fGP9wDMRFxC7f67AVr
UFGXSznrP1E73t/mV0ghPAzN5dttJ8/pKpfHgQltYTCXcQoYMqjJY3qoiD5mQYKc26Op6jMRQrlR
3gFnGo/D7ONoq9Q1AloF13l5qlw3O/N5bnfSZ1I/+XZKTmUy/1BOedTypuYJd0pl/n9MyVdcJa/7
30Zzpbt6RTRIInjFrXyAZAx4fyqYawB4rLGorJgEw9dzgqFx2md8CrFFP6eYqprOadHVX5qWlgau
1YgpEzUJPvXoSbMFGzUj8yse+fgu8Xr3JZEJHClVNOpBUPHwNKZ2CA9LYUeKTls+Zx71GEj2OWDV
3M0HrrKcy5EB0ockxU9su4NdaaziZK1wmUCgN8A4OS8/sClyr2/sfzri8gdG71bHYBkSXcyvwGg6
GS+eFso6YrMWYZj1MO0Y7dpoDFYx/O7zpcQHXYBU1KAcxOq9iiEMznDlibofyEXLZAQ1xquPUeL9
d1KeyKC1dP/VrutjrfvVq9mR2cYdlP4a+J8DL3wK00O9nEfucq7cfM9Aqx64q1mfBlyiutiyvGd0
NsQVB5IYGb+ThEk822m5qtWTcayUz0MgN5ujptKexEofaDX3SEuyGv82YKUMe8JXtT98xBqNTF0g
r+mgQrUDa9ddXY/6QFt/O5Msey6SR1qBZLjgcgKozVkq5W2Ry1M0RJ9NTozWjPC3Gav9a19Mwf0K
nVL46+SeEUViLfbhwOyqYMmF0MOT3olOz7kKgEUtiIuns77qGc2zVUsQP60Osrc7ePNdfgNjrv6J
P7c7N3+eFgkNxGOHg90wvQr9eTDNn636FYIpPKPmepywUwYzKLk4YvgGg/wIWaLKhRacW9AL4Ebu
trSLpdL+kWNUkCTaHd+Uvaz/pTUYo8w9V/WyY3wntIGb0b5lc3iUWjWMlYv9uU4D21mCI8x5Y3xt
nZcim52RC/qXlMbQydHOaLsmMaU3scBzSNFN3a5n6RC8nByjJAI+3RihPczqrJFNnOcE/B7LGz0M
0v/EXNvUXnc52EI4C11PJeUzoUZ80C+CG36GN/+i4dIqESYBchUTHXUp2tkBVpZeu5CuLt3jIYKe
IK7YUSEfNRMnZ5Kbvh3TfY8uragZjJy9uR1M0rB0wL0zJV8CS3L7Y5B2WdTpX8sS2cjQEgdVbuHP
IZgh/7g0yBaON9GyAOs8VoOI2DptA0HoGgupDxTSCMfx9xkcaN7OO1njjrEFg1qrKVH0DrE816xB
7FX0WfNtGACBIDptb7aRRLNQjCl72hmENvZg/V1vCYCBHxVVTl9vLHKMLxjjlWnSEiE/qUA+771a
0q3LZG9W1q4ldYJ9+AYLcTvTwH8c7/Dxli7yCgkVLxVhD6ohGXfeBFBwvB4hZQZWzmRImpKHjfBz
CriapqLUbjoKH6QBBzVyhd2/Wkocu4MDWM/ZyueCykkuuAlW2wm3MVxQrUoG/vEDeuhAejIqZrBM
MySy0aTqRTPZ8g7IENxPklc15KsVv6JIHpuYDY9maGA+PpQA3jgZlpOpLd25P7Pdub+Et7hZwdA/
/FU02xg29mgQ6U1wAmQf8Cuvmp/QzsUyxKdF3Q+4k+04LcWfBKMMwPR0OEct28jc2eMpIuUXPpfI
vMaJwSHflZpppfP9aYKGTeb1lvi3bWQLCYWZ6h4pEE8Qtl6kMZHvSyvfCRwlBXtZgbow+xvVYXMh
VLT+eHCjmL9BPtmryec7sK3EG18joSvYwCIBUI6CcEFHSATawhUyX4f1omjFD3IilEOJ0gAa5wKy
mJ4ZPe4zVTVqm8RlZ2QvE/RjoOXGV8cySuoMggdWK7a3hP0A8vSQzm4qXj1ks63XXAz5jGVhGMAJ
bqz3bqfTi/GBZUkK5+aNPA3r2F9JZcPcE4jGYO7wS2zDsWPKZLwh/9Ilq5F680k/jm6Jp3MfQJPu
b8yFgrnmFbd7AysmfyvflgA23CoYux/mKpuYzgQFKMevlHqZJFSIr9AdLP7FBUQzmcNghIbNDLth
LKu/u7HMFgXcSbZwojlu5LVQBL8iuQjI/Dd/sojUvn0nBZs/D/kNnlUg/fXqxmsnEVrDARVC2v+k
QFvCT1MqL9RZ2gRFQ7aOFsonUdZBrHlrAg8PbvEfRceFSUoTEKJrCzNV0T0nICaKiKiBuqC7hd7D
Cmmd1TZGXJm1+GLn5XmUST2NDMJyAt+JPPxPw6yD5/j/x9AFZNkzePYkHS1k91L4+T3fTC0pk8SH
n/pdMJm6Dca4PCfTW1Lv/aeeoVH/fkcwDPxiWe9MS+9qLJY25Lv/oF8FFw30j5K+rO3pzlJJgXLl
ydivoTgH/Ve6PiOj3PUxo66lli0Z0QeyXV2DKyHJ140IT1XZ+Mk+BtqKmUY5jGvUIFKau08FPXnv
70Yo0L2rg1pxZD7s0lblC+y+CQTSAFk31DEfv/u3EmK3/hyNpBvon4HV/Tgrd/kxyz2vcNAEI3Rr
6AT+AnGxwfKDVEPFgZn++0sEXfVlGeltnW+lN/s0pUTQI2FCNSHG0Bi/78+jlCcK7j9MYQTu3F5J
9YDxwOAP2C40irYi7r4F9LkZl7xzQMMZdXUkDXdUown6iQ46MP8+vD4v+MxjE4VMOcgXEGB2uXDN
pe83VD2Cu8LeggFuuEIXOUa+hGs4CHCp1kH1uhxLvkxz1cVCJVhgTyKHscsMBuil3Qr925kSRl2Z
Sd/zw1mMBUgAlb2zLHpy5uf1vHmQhT7UudKpzJEZvi8VO9lHzPkrWayAa0C47WkfyWOnhLoF522c
2nqhyWFmw+IsOqzcJGnu/iKwCEA4kWfVAVnKpMrbYKR4Bp91e4pFJBrWcOWV0qoQN76sET//bJyE
uMWhiYjXKCUL+1Icd51MHr7I7c9fvQTQkUucuSjeWNA/2gYc/fVLXmwfFXWOnD/z6N5N46l54rDp
utuZyMC/alkmlyagdfDtUpfXBa3quP9ZqdESusN5esuxn7MuzSfHBIGupg6zspNaO17Jk7dU54g8
4/YSCjcmqFs2Squ7Q2w8gcnUtFtLje1lf42xoIgZAJ4rqoVR5IqC3B/zahAHeNXxPqSxOjpeahM6
P5etPIYqifLrqadHCWUPLROmpTaHhoRqcaH1m/KdAaHLcGn92NBN4gKS8pEEvFkHxQJk97frhjxR
8xL39UwAQdoCqAOTDcIgW4OYknb7Xl7vEGSrjUAIfF24aOjNts4JF1a8iPE4loQfSR+8DWMg2zXb
j5kes+eri7Bbn7jxFh8SHjsbDo2LVY1CQilhGZpauqkIRUM5dE4gkqRDJhqIvIlDnwNm3wneYpHU
ZU4PI0qbXMQqoFCfNW4Oc0dRlm0oKNdxkPXWWesAzuKnwFboaVKvGp1c8Cmq1OnTobyS8rK1Tlqd
KaQSvHP22VkaTqjx3bYGDz5ZnFOXdA4GBWD4Ie7Xy/5SVOE3AklfoWal41UbIabONaojERDcYuLw
gCo7UoFAYezDXJ1wdVBrRq+gQBWc+3/qdcdtYtyIUGClvszsT0O6kDx/GebxCCxekuZu8y1bfVpI
xQ7EJJrjv7Q/PrZDmhksBBRmK1LpyeTFwJ7VSorXWHlNXTuR6AOiPBnOv+mudXuu/bedxQ9plQAi
PDAXVzcufuPfyKaygSBktP6EREu3ZkAWNRq36a113eR067Hbl/b1JsDL7up5vnemNfXzRisd0TD4
hshNHbno8RMd4fj4KwGue0Xn9OC6JYdAP+sAsIFLvqwPO0dUjNQW2luChvKHon6j73OWCLTs4IMb
W4YdXz6JKLqwdp5hdrdGwNOh/HTG3eHPbMHnE04MBmHSF2WxfD+SMAQhNEqSNjEiWvCcRtBGqMrB
MQGqL4TGLb1m20RorYPNchAb96jKnAaBcmmT1yTyOJPdA4f19/fVZHNUBrCqJXA99NwAcWwgfyq0
gmLRD5ALQIy8qBdl5ytmfgnpn/8tCsGMW0qMBzCQxRkJ7HeeKf0wX2sPX4CwNd02hF44P4WBdWze
t9B099TT0zf7wMZGOmwGAJ3UO9LINklmY+AmW+jUmzXvOnhnhnD10n1u3ktUaKYumi7EB1RSC7K7
L8YAKZheFHH14iY0xkyus3Wh7oyvQ1wAWI7BFkEm4Txss0Oq7rQ5V4tOeuMW54xJXT1hEJ5ohbRu
NeSYaQXi+7jCJhybeIPuvgQFf3SOWpYIFYJKUvWFYbWbizsAi89EdcbHytWNrwNfWLdcjl/5eRY2
IRRNsbLiV5aMj4iL+R6EPia/Y/D52mf7wHQCmQWvHSOrlBiXM0vNmaJ0nD6YPwyqDsh1O8OUVaYU
BsOQ6pP530osONoNPiW2yQ8+cmYDcMi+igg1mFfHBKKt9nYak2CBqzsx3W8LZ1cyZH6tfc37kJ7x
kXs21bVZF/aAOrjFw4EZUTLPr2ucjhxXXgvpqNw3p/NVicSJe4tVzkD2RyZSJzj0likOXbW3C2rr
NvCzGD+XmNrilc9qMGDC1qShmV8wVCI6Qu1NdPuigyqmek/vuOeOaOJocsj8B+v+QG9iNNLiUi7h
0of6hCMrWM3CID4WyM4Yw5hfT0OExobPqecBkamVsdODqTljPVqbOBYnhRdpmwgixIVgQfkRMtX2
qnc0eiQwvOBgaB7HJpU8wUIyoNZyImZczO3vqmEA1jULNA2WJMIJ9GWClKLrjFHYkhQJEKjefS48
Ykdxoj/NwT7aD5qMRbNnd21jpnXGglOeuBQ5Ppzy4a+Q3Z7oRL7N4rHINdUeKagPIqnWElrlNRm+
BczQSlC7bTygHrOpHxNCUC7zF9BOW4P7oCtNujq1i5zMO6+TU1KATnzxTFn+VUeE6iUu2OsU56n0
DhgGfpMGtue33EcDgPAs60OazcdFK4gs0yJrWVZ5EXUTE7elYeYoIRiXG6uDFTi8rV+HIs4iIoMY
5h7scCw9jQBEuBeMb9X5FXEZkaSYHwtCXRPg9YOHdS/5QpHXDRk2aknTjMx6U+ii/nBoXacCp9Se
BVX5U4f/M7w1359Ddze8/M/lI+FnPBfLPHgh1+Yygh2SmlR4sg6TYd/2Bc6I/Ph+nUYQRkwHWLu8
MP1auhk8lN+zZFZNetr/M9uTvQ18OqXCkvwJjJN6uT88BzajQccq/9sKPKsiZinkCu0J8nyyMSUl
4mVNceQD8UgS+5i26n+oYD/XsFUzc6g31tDWXfXwhuqd7IfiA6+M8yvR8YR3QD61kt44XscOQlhM
K4hY9+rpI82WnXKIzhTsSwNk1g3u0D7lBY62eTmtrsHNvkmSP2hDS704IQPq7YM+T2/gHyNU2w4Q
pf1mfHdWcMiID3BZY0dbcBv/wSXTVXZRioK7apM3fXPelxcUxxnS2DFJD/fpAE6rUg1stRI8rSIq
igtt6MZ+gpe2HjwpCDpKLLyZryq3zrN5MKJKwEIOd2heqaexEyYZc1OOgqrQlp+ipgQ1YV2jlrjZ
axGhIqvu+GgRhpsMfwh9NQGL8NYpQpf1lsdQ5nTwXU+An8k8HYzvP/phhddJxYgPBgK5cWu8TJSe
KMLZqhzfmrcqaRut/I35q+lock2Ggkaz5K2/CAdrj9APGk4KIwdcxGu0tQ1B+rd9mEn/F1RqCNqS
wxsDUIqhR9iwV9ji9rKlpmeEgBIVh66mgxfQ82gVKnJTz7AZ47ogPUHJGacAj95Pg2nMM8W1RAXP
0SCSZ2/aXJGBsVUId4kfOjYnTBmJAugvJJ0oep3p8fxwt2MBwHW+cu64Qy65DBD0f2peQDUEFCgs
bTXLuJT6Xdn+vVAaX8qmzUHiFAIV08FXGnqiT8Ct3dYxm/6MMTR5yWJ3bKi5WxVO41FFl7nZYvU3
v2w9l1CSP93iKUq3kcnELFzkH1VTDMaXLmmY/cUuIjfSyGQ7wQmzfXRYIpLjntQ5RxDI/Xuro3EX
xc0Nnk4Rh/UoN4YgiIzCYCE6k26VVm4b0oINGQiKErjvlPxf2KHUddSqy208ugetTn8GPXfBwjbQ
1UaQLxBgKGhPhtZMxrcG1HisGLGMLqnfAsk1ZFFR0Oq3X48ldt31WEPG9fAIud1MY190RmUJiUhi
2e5RnAKHqgssrrBcS7qlqaMFW7UKW0FupH4g/gcmCoTu2v583/QQaQTTGNJAo4X3FdYeowLNIxGo
x7M60ODKe4jiy/DF6dBytFGOwGtT8aLgkI2nkly+zZf5UMSCVkoJ++eue+yvp4cldatsQgjKtyRR
Va6a4t50hlg3KTgnNQHXdwr1eZyk18gxj45UKFNRI5VJJJXLbhKJK/RqIpDzbGjPDD+Uj/NceZA8
03+UN64ywoj/DwaOWplv+VDCGBqTh/yMNHBIBIoLxNBcnYW8BVsX9O9SGth6Mufttk98e2fvlpbu
p+NFGUD3zAIns+F5jp2C762ceSBOE7eHab6lU2+unOutVwLovBbM/qIsXJDWxx5tEhT5Bst0MW1H
UKyCreK8fY+kEu+NKEHj1U6XxgjovPRLYWGhk5v4AXnsTNLY8rlSwKlOGb2Nu+tuP2AsFzpkG/kv
NTzbxslh2M/VJp5MzmYkW5WYcSi1G4/HTdq0Dz+a4VDFOdTa7/ppy5rFhOcBOdGJ2A4RpWi9K0IC
08Zz781q/0QC9QPSdMZ2uWa8z+JtCe9Jn4cBR9Aia4CCN+vF34v1//LlJ0EkbfHmN1QJLTZ8I8mr
NS0dQvRixp7gDYEv8PEBsiNolt25SdxVUy1FhhICV7+TI7aT0YNxrRow2r1nzNPLEpFUzD9Dt+p/
0Y1umzbUCqzJhOuyUxWAq7JKp1S5vwXskNLgSBzFBdMS8ToljjI3x9tWIEwH8e9g4fUI9DiwmJ/5
wUVSA2VlY/sG5k+0xCV6SRRmk6zZs4UOLpthwpIs/Ue0ssbgQamEDpMWub6Xmjg44XVxI+WzptBg
UgLWP0jbkL1RpaizCCC1oLwDQyAJJGXw0DTzNwnDAB8LfQ7PsJwEhAPqMYPY0ixW5CF5yMCchqG3
36QOanKuodn/aO8W2F0+C5N7B2kht9IuFxhII6dgW5aS2ogm9s9dBUWVFcoMEST9606x0+aptRQi
7zOR9BEzQXb5JqehCzzRmlC+nRb+Ld6K3fKEOkHoeSMHp4hsNHiZd7a0Rx848k3USARqShJaDuc/
RLgfJV9O3yQ7MlQv+9XBrecUmOmj5Oogz+pNwjIZQjYmNZ0agjPm1uyL1v46ni7/tyj3mnZ30FgH
oSoqb7r4wiPymsWmU430etO01OIsNEd4okTtuOzIwr5zb9cVcwEkUhjTSm7/2qkq6uvnXwridemw
jdStm89Qgz9O8wZ/cUFWxty4L/vD7dzH0h8qzHRd7L994hgcQuLoO1B0vlxVTuHp3pj97HfsM5Qk
jNP1SL/B3pxifK0oB83FHFKwxiEhXVX2FieDIm5VMJ462uN7IupvEs59Mb56ATUGAG5roG0WptQ5
+MaAELXAofyFxzwjaqutEa5j5m40mecoUNRLk3FR5YEKdG0FCKuRLh3mwGPNMaHhBV/qBsQ2gbye
kDe7QGsh4jiHyHfc5pIfX04nB2KBeClIiu6B8WnlJdutaMdT2K8SYr1FHULyEjq1Ag+XdVqa6Wa7
XntQOt2e49eEjn7KdC5Qxadx/M7EaMi7JV8ZphRsXVL5dAd4fmSblOD+SJ3LEuvUJPdPEHqidDYo
l3Odrv07ojjVZ5Kx9Yq6FXto76AfEEUziKOUm/38kL4//sNh3oY7cKEBhFpK1rZtUNjCEX8AFyMb
YYDkaCeb6PoKP/fCO+Sdu6/8+3yDbNY6EJvQqcl/NufLcGoE/Kq93vSHIm+c6Dslcpy7oxWv01d4
fWl8C0KmSuQZwH3xIGgU/S0YMQkzmIzg69RToN3HwGu9m9CZtm06nlgpPb90Y41qdi85gosREGCQ
9/43VYJB8P4MT6ejvsKLmI23HP9UyYhdQ42/GqipM0SBb1KSTtvTjamblS2pKdOBF7lJI/u4jYWB
2pOXoKrENV6yxwi7vIgDeJPVhZ11zd7evyNFbzFNTztNLzFmH/8erJalxQhGJoQbpGZsSxe5KynK
WEtgSeQOAskJPIoM+n6O4DRB9qdy3zICZ4Yui0lH0UGU6vlwDGvGLwkWXW9Nxc1sB04rMRFL78Nn
FnhP1Lel4b5dhqQ9OPm1YIVvvLcVO5tuyxqnqCS89/cR/BlbsxoT4UPzW/jsogVREUJqVS21V/SR
o5eEbfE3RQx8roGfinecvt/1OIzPBrbBGV6Qni9vAAuWBukhKAb+bo1QJn8lET34nmZlh5qbwYDF
6RmyOPl8Ht19uxC4yx1Wn8ZOw+1OLBeJpC5byrk2reYulfTE/5ZLozKoXE/uPYkdnqwbSvltwGi2
wO4sLVh478LxqqTZFulwvNRx1IGiv4A6jcUeCmxn6COpgpAVUupCmqmyN9TZqvHWzKPn49Hj4iav
EFl0C7I4l2Cy5gqvZqrzLkavPH0hdr/okx5Cxe6vb+NMc6sBHyy9i8LzWQlg6VKxLE+HE45kIg95
Ota9X8bkVKAHg6UOibromrgivnY1/w2vQb8JCbqlJjXbm6upwp32UDxWxMZIRumiv3q0aW5LNnji
G8eRSRI1XhySpc8Gr3/+wvebNkeAs2e13qSPLLQBri7duLNSli6bi7851YstotLmIylVLD00F8qA
NC65wScv1pAxfLP0zaRnBZr7xeXhJjjsP705cPPkpDi4E/E+6ndpYpDMfFvdR2BbJwQ/fqra5JK5
klk5z+sZk2ngyjv2hCm+UJVocgIiKUJBdR9PwIKJlbLNTrsIzl41KXYHjZvKm/R4brmZJPG51CLj
uzWPoHWAnopglTBc57BLSl1r0ylKtPFsNJ+HPsnnm12CtBh39xh3abim2HfNsbM3mVdn1sxQD8d+
qwznYhsGIWzQhrcOgqt8NrvZeYWCWQw6iZMPtE3K5xMGI7cMZvDaaReO4dcYPWvdSpW0n6Ycdc/D
pKZcIt30ca1AAnPzQMXaJ36kVVTIXUI2xjf3BKm4WhZgfxtqTyOFNL4zFRz9WBlac4YIAnmWMYP+
X2EzdDbSchHGS3dFQIh6KsFdhGd1hLuviKpH3thF2FtTDcn7uyXvevsHIp+OeaFNzkFDreYdk920
aOio1k1FSuKkZ7CyT8/BLL2tHmYysiVasSm7kJL69k6QCiMfx2HhBH7HCIY4Gi0tV0WK1r0AqXJn
CpZQ6b7LaFU3Sbo85T4OJ7nsi6BLmh8wZXMqQ7Nlo+cFuqQf3dXA99xs8UGtnTaM/o++RkfUGtqA
yOVS3iw6s3V8wbC1WD3lOCtxsNZQT1swyJlq7Y1ZgqcSJbxsN73QqZLRTd8xrJfG8uE2hstGbHAx
7pdgz+xvAUHNmJgLlvdUacUbXp33U1YmZkr1x0pRz+emEWaxhVPTBCAfnOfh/ny9dUd8W68mfgg4
hNuEoz6WetfH8R4lYfP8LjBX/MQ8Ls1kRq39BysIcZj23C7hkVRjzu06SwocxOEZZGSPXFDYdaob
UG+Qx1xNHXygq+O29GyPY7kVQ7yT6XWDEjiXE1fDYPvqYigMM9D7FCXQ0hYy63VoRg4qOmsal2nk
9bLsg55YbdiP+xgyX+464hZLFSlJXeVrXvmRQ9g8p99Vky/aiBC1tP+ZMsdSHGFaEHYNy83YMO0k
scLoyWV5SHP8OYYdWRNN/Yce87IFqad+Jvu9uJmKWfMOQ8+SRWrUC5V77NfnClIHWAnymr6ROawC
UZgRQurfdjFye/8PHwB/eY9+o+n/a1lkpFmz15XfKLthjkirWXiD4XEwoTl85iynWy+TPqZCy7kz
kmzJNhFv1sdraZXP2+peQLVaKjBEY3Ttu7sXV6AvyRP1WMNHdlu3/QlVsAf7SNe2rO+J+ayE5tG2
AbV1xyTq++1vzf3m6oVE5YRaGsnVz7vhwvRcp4oLxTsLewaGUvxb//vMrasDN9A7EPm8GOiPzuF2
1KfDgNUgGyBLchqA3s16qeIbfQ8wAbGJafKtKCLgElnGy+q4r/Btl349/E225nBO4OhP4Lx2hzc+
Gv36/+0Yzh7aJ/RwB/eFkPtZ8Dtcy2lDpgUb44LnQMCqxVSCzsCjau4p8KX1fSlWJ0KFGSEek2I1
Ypn9OjuLj4EsD73U68msUvoomMRLYvrJjUd3RsNhSJsfLYNSvtse/FJTPxcDyZl1eCwGRWabk3eE
Xh/Sr7ZGI7K4D2VcV9FSAo5oEG+O3aBOjhaHQIYsM8W9+BTamGBQi9OLSn837IFWi1t6f7N9ZcPa
UHE6Xim2T4vb9FhLS4vCeDPVo2GlMlKcl10JpI/DD3sg6L24Fz5dq3TURSuVGzwR/KxXXBq5vfnv
Hon5cG3NxjONhxrxyplnCxYkChO8/ach6fPOsuqJ95ovraCWNf1w6wvN7iViMwofotiTogP8TMk1
/BLjjloX8nsdeAXO8tbThbW7nrPuP05OHxiyZ3vaTPFhpYa9JiemzK4WuYeKjhVg2HWkIZ6ZKpqt
z3cvzWwpFDpHpzq2tQD2+NdqcRskiPKodRlPVSC72IIZi6YVJIT4FKxh4X3YrV8KfcKsjHGN5647
7AC0IjUF8RI1b2laUk6gREvheiJm1B6YVSejYdfoo/TEpCXzI3R2Vsa1me3KWrFot0oPNShsyvho
UN2aNwL/+XMZcFH35O7KfD3D4ZRAN+JGuK+4O9ZwEyoaDBetcFDHKEg3gXSTFOhMfGjWA0TWQBMQ
mHnXmQHI0XKZy8zCQqW+GxuH10zfRYiBv64oU6B7uchJ13a409CuOjknxjCUX/qdqFDumdNKUsWf
TKDLhGtf/UdKeWU+1rOI7ipgOqXfd4gQyaCIZIAYUVSs80Qe4i+RqktGerDzCIItZ7D7TOXy38IJ
iquZQD9jQ785x/F7+XxoVohr2Q8zfn5EVLHegPpySWYbg22Tlz3p5zl4KG8THkGJjvkw5JnCAKdx
Yu682MTseJVHmLcQvdMu5rbEIIwQBR+GAuDxlStO1pTQBJ+OjgXFt/Y9fllHGJSWatUV463BrxQs
pPV4deZNmTfwUV8If0sDNoJxX+UdGaCF/3Ux9+yqhwhI8OmbqBRQNvbU8Me/OJSuu0AC7rXjbW/O
SJ+sA99VQJyNqEcAAU/C1f5sRUB+UvJKODTbVp7hsEtcEQ3VIo/wPnxu4VS+44jIfrKN5IuCnlsB
5zKmvv8Suo6LHagyE/nuH+MJjr81PAhnUeQT6BCs3Vhb9mti9H2j90gQQcx3GcMQLSAhwuWe6Rdv
EDjfi6t203DRtKoKnCshMIvXSr/xZ8J0tWs80f7JA+6r955oUUqkTa0KNth1HyJUjco9jdyvbbi7
iSbCIsIroj3q1VnsJdrwB9xKXyWMamvXmZ5CZrOwX/189r0EaJ16aMQqBp5DMFoYW4r4crEuU36S
ssF9Rxkbd3J0g/mW6sdoUNxq38b8CDAzNeOSjXETjZvDYuxl1q3DcflApvYMeuBAzWwNQHEr0edv
jbE9kMFotqoHtOquGq/h+FnzwPjFtdNPeZ7CkPmIa3xsbeOyo5NHgkch9XLHts0zwcaP7ZFcKzDi
xYpPsMr+VBIYcYIfu44p1LXp7yj5h4UfA2lvj7HkpTsne/hXtm3yabmysnWdvsTTAxmpsrUK+Bg6
JKDgsLCU1zKlBS9w/S4Q2TsJ4d5yWVzKDf3o4l8WQ7l70j4sT0CFweWe27+wpk6KHW/yGRXoG5KG
AfADQ43883R7EkGZvSX6Wkdj49VM3jocO8TFfggYgKAejosRe9yS2kwFo7iA5kKGaoqmo43mkaQc
9OJSkGwNNc+K1/bDBIZU9BNBIl9MBgjP0wgTFTKvbtWAtb4Je8ic4ePzjfBlDxNgR2yU84uHOKD1
8tMgJdyefgb9xmDmjChTTu4MjAAuH/J1lwFgVw+FTvt6PRtYoJ1MmAl0iP7HyI2TM6ae0/KKL3Q4
lJ9yTyb7KLB6pQv5GSmSYRsRpQINQlZheYVK1cICUtCD+RUSvgM3en8uKCtJc3aj52b1J7X1KwYf
2gnjKQEwBByRsxSweds5vOQwacnmft1BXmX2Pl95grFyAXW40msTVOdcW2VVpKjVcyV8c19jbVVQ
g6AjlEAwr97BevH58Qp60xmtrZ06eM656xcVLOcul8cKri+xrALKQSWrfHDHIzgvIRnfmoTlPh+y
MW0YC5E3UHMuAAf8mYZeNtg35hWwf8NL+C4dGjH7MhnhqQxeVOhQAU3t5GwQlHHisndctyIFDSzf
/+oi/RCw5xrL1RXpHjlM9ArfTseMdf6GceXZ3L1K+Ph+A+9Zw1xLc29PBQ1uZ2hY+wO9+ECZdwwt
D+sxJRUcXRbPxaIk0GNFzMOW3K0qj6QHkdJfi4zSNUIlnJ3JMKtLfCUE7sbGvqaWwcf4MSoo8l0G
mEwkRR2IJNGotA/8bWhMmw638NDinxuljPXhTxp78npLmwMU32ADYK5g3SWtMcmRduu9mQZlAas3
ZFSo8/xQ+clACkncwNKemUZgy+l7S7ZiNrHJ6+OzDLwxzCIBSdwehR7tXWzwpFyzP7jumSqvTHcG
fLzsygkQcBylqFj0tq2bt8ViKwmWAc6rmCwMnc+PydCjSO+psDKJyMPPAYd8Knw2bwQdK7wWWTZB
q60BcmByp8ldQGLBSAgn3apfIdaN/sx/MGH91xrqSiseOlqS1yM/v2h1lJBHIjPDrUhVO1z/ReFF
6no5+HyIl91p1sYuDFwM9XsqTqvOh3Q1+dJGeSiEo+g8GxoyOqD6SVLo7eOwOs6QgzhW6i+c92qH
0nDZesWq3eFANHenNvdyCm/E//+xnTWs2RKnraVqt4/W1Sv2h5pdx/A3vEQsKiKPDGDBBEkFiTiE
3Lk+A/V8QFmzGe2LAc4ifJdTh3PWrSSoh4l36m46/q5jf7CgXXCu+CpMfNJspzhsRLG7BtbrHtG3
mhLsmIGH38cT0gnvcAaV7muSXR5v6DhgHioyk5pjdSzmkqZbC04nOwUH/dq9dc1m0LU/NYkTEH/k
pCl/BRNeeKCIycANyrSs2lqukpVRyT4q5Sy/Rk3Oy5U9G92fGbYssvibGrSWV7vZ0gHUdPbzCYz3
FSWgMtiD7KG7IioJCIsWaWjIV7OtzeAY9jCRWAMM0mcF7kjt1hLrzSUEg0UgLSVvQ0D7Dxi+Ey4/
JBqlV/cOpq4m6Dvr9yLCgyIyRrUjZW1RqoL7041Ix1QvVvL89Z9my0cDaqu5tievbHNlZx8NJAxT
4e1Wypi4tk449Khw/BIsMGW+iHx/IkONF4VU1OJSVA7LLtjJLyvC16iCRVC6DWEaKwVCWMti2Jhp
QI3n63HF0Xrd40eLTkBQq66y7Hw/5+k+SsUp8iNMVTDnTSk4eXVAcL2T8pVk1nX2Yvtf7RQ1AXIM
rWp8w8lHI6yP8AoDer5WYhyEZlq3j7p/7HVYtYd2NX1Ze96YO/dvbzAaZATywRszjlpmVZkezZSR
SmhJS7zRgC4lAdtA47HwZZ7YLhh049odJEgumxfr//NK88kHwFZ8iAALx8sM6mY6cgwYxIfXJz6z
NavpRmkoVTWdPD8RQibRkTvr3FxG01lQIgheFT51mMLRWqCkDAfyMnrafi4uVWgPjT0V7x0NyZhI
m3G7CHUwfJT5c4pVPjezC4JHLf+KuBjzNEPnLNQQLPTYrw8D/yAkcPB8SDdzPC1tOYTWk6GIIiEC
ROSAeNv/GHv87KM7LL/PCF661H2lxF8+iMFd838heykUX8g4IJXIaWqwAGKVna4i4zXBeMUFk3NN
35R90DAUp0Xhk3ME4gHSyiueZQNjg39UYvwXoMchDt6NtVR6Mg4fBbCALCxwrQiRGGj8uyRZq5SP
j97w3KEj+TWtcWdqQOXH86R2BMM9uUuJFkwCLtb1boVnh/wCnEqUFXTE0smiUVDGKzPaKvcGuggG
1GZoo8x94LAJDI8pN/2FUn7iU5evseXcpZg5Y7BS4q1fKCG3ByYemkjEBgfWTtto8Be1HDcxhlv9
FhDzcBOp+9Pt4NoSjnG8r3QYKoXVyximI2G6E46/fCgFJgV109KwsdTGmDKbk95QQTUx4fWp8qu6
+k8rOD5IPwvFo7Zfs1SGwQzhWBI/q29DUwCp2xsOvWUBsTi3gdurXMiEx1Ie5fTCLax1JVVeV2PP
BPzjcRzC47mdAM+JZtel7OMz7KLhIe6v5Io2r+vv3Z49MjuCyO1bWZ7iOt10z4+0fJYZvGfP3cRB
HXCSDsstFSizARtZd8FzfEFDfeZqnotmROdFrSWXWKhsj/RlcYIiyTxSws5UrynMMk+S64nYIOGI
F4cYBswAVsy9z2OGzbnA5ywTzN9EuKtkyGfi9SeYbFUWiMLJDzGGHmTBen1OzeJpkahSDrPF9IWv
i0bMV4o/KS0kcQE6HVxBuDGO+v5/dWwJ/OZm6wvJILDDcHrol3xxrCIUaEdcGWk1AkSBn8rSCLaj
sIixwWpvo1PtVqN4SNsLrb50KSHiJNf+wH4KNAQjCX1KMdzX+H11eoCa7UDpdnknJZtSpYeR7TWp
Rz9/deS0BvoGSpzYqMUsL1CYjdKt5ggiNDFRc+d9eg1sFioPv/RwRy219pToKM9CtlZZSPrwQKoD
ejO0PA/O2OkOmqCS80kU5XJr/Lm3U+S7+r+pCer6Z1bJYHEbaVPmypwO+eHIav8kdaUxarENQcgG
NllEqxfAMMysxAfTV4Z6WHBPp3tKAifA5y+MRxURtqdITg9JlOzHjMQx+gM+5L66XYTRdZq3UAJM
l0hF9Cfx/NadCVbylwKyy8YVbvQoIn3nQqMMq958CNcNx71LSLByj71kXE6tOWbh1fnA6DEZYNF/
ArTrzmw2WiE0n7IXjggKgp5PoxO47N31jAIo1C/Rieds1qqYlNlDc6wwZqR7vVHNZzEbfMsVdpJ6
+DVMw/Fl31Y80Xs984RJOqY8uva7TxXzQ8XEXnqg9wlEnDeWDrY3oXQfZ+13MR9vayqnVrm3iP6v
PyDY+nhkMRqQbkWqLhbkeQZoUtUQYQCNaHNc05loPZGwUg5SqBbOHnmPPFPK5EMWKAmyKtNSgC2c
V2ewTHjvtf16QdXrL1QBndOPTU+K1uaEbrI2YRJISS8mbZkKvPG6VcwY2htLIR5Ag1kWamJroqQ8
oQePPgivJd2hU9r3YoMQpHGbzlcllTNarIZhgB61Mht4QPN4/xmpgIPdcJuNd9LsK5RHDfDkLTzJ
KkkYfg9iNVI2lsByX/DzLGxr9Qv/KdwROdGbq97Nqh0Z3xp63biiZCp1qmmyUy0+Mqzw8x+GrrdA
5oTj7vSwlj0vmIzpv28hngNs3RUT2gir0NKmcIjlUVNU5RW11roLqI6lspL7MfOkLlicnbNGGNpO
m8Cb0y7zjAZxK1UulxSVJaLp2ZOJNxwhrqGP0NXu3v7aVlxrtx6Ooy4v6AqMQT2oUq/yZ+JxTwdY
fApp0T5gquX+omGjQDSKLV909wnKbeU1vuah+plQIYASKxpMgAWgZBT9BqO61E+WZZg1AynoajgX
xWIZfF6JvZbuW7wDzU1umTk4UvQ8qtx44dhYnFWCQTdlZwFO/LMaNSQ4G++Bg3MbgD74Xc24254z
fmr95Bmzw1E+gi11EXtgQBZi2Bv5ieklpvEi2/XB88vwVDNBw92T9hgr+JkX5QvbcvJMpUcGzUnT
LcJmzSekmV5V6mj0F5QSIH63C2F5jgpQeZmtQBSJncq1pFbBBaun88lxNnoWHQ6wHz+E19gloJ3c
yvIhkUYxbz366P3AHg/3bmM2geg9W4aHiAKZBE14lgkRWtLOZTC689GvCPxZfLEpSRVB353Yb7Sy
NeH0XENxq0uVQK3I0wInhbnejtMOfEcUx+a/5DGBDSyjAbjmUahbeA55soG9f8AogXT4Tks+dDP8
bxk9lUN8uqRhZJJRKlno4neeCrS5FzmG0l7GjxYNPqyAN8KSD/eWjSajdTd7BgxCzHOMCaf3YNy1
QT3EZ9+FEFKOJufG/qLl2/vVZDRLciZB4ckxHBBn4qBFur+336kJa+4UF984iRiBcaRBTVmOCdMQ
bcUPZbf5XjkpFCsgCWac1qdv8ngbsyTzBnxMlF1qMcHhvisD0KQbYv+ttIVMQNRArG+4C+hcG4aa
ZDryi0Yw6INICwvLHlfoqBV063fXRmhgLAQqQtlIM345beMNbKJ2uiw1cHnH9SZiFzoaTh/aMhYo
eFZm00n4HD/SbBuVOdZUh+ULCoCCJJ1RUAJ07Fwxs0OvRA/wfmZbQUb9ZMo3yD8quG8hOXXn4GCz
uOUBbtW1nCAkxSmCFi4hlUUFF6NiQIHU0lP4FMQymH4O82QyS4Y3W2c+jZ5lP9w/QgkxQKbwNdQN
a+6kqn4iyGUGZnJn+uawwYZMh+4x7JzCQ22kKOgZfURQc6m5wu5aYDd8oEhTvL+KrFw1KnFEH3aa
2K1WAR3hZzPNys7cMoPRq/zXEOm6BhJ+B7slWo6y1yfH1cdjYUTz+jIzLRlHNmKty5YP9qgpOE3H
cWeiQ39Kjc3SNEGrhvSMzfF1//oCbTAD2Z/V1SIoLzTyKk2VDuyiO4OYUJv1NXbuz8Dew6/mSnpz
FYqES9FlrfcC68VhTuG1COukb06L7qnNQXgrLUhI296QvhKcLhCyeNTm2KMhf71nVfKbfLDyot6a
0drap+yBotGJ/U6Vp06feOIkzqhtZJ3vuLY2UH7fPa6as9VZIDkiGgyieAvzZpJ2wKsKISV4MJF2
Hp2yvTTR/J7Vw9K9hntoxGieF8dy2AeIU2Yi13E62YMLpWb/GPxlTm3ZpUkEtFMenKclg+xYjrGP
K9hnggZyLauTzEoBL3zLDKUeIVHPTvcXb3mXYknaW4fcOR7TRrFWyI0sObvYBqTAOI60GJlMOHAU
IrMhixZBnPC1DbYVz1bu061xtKAcc3vM7WXbjC4b86ioTMER0yrH6vscp7A1FPviXCaxqRS4ymp4
UvuNjaoHh1Qx7HyV5iHZEpOLdCCasM35A5CHBDm/f9nDwj+vc2qxcTQBdC+V7sfehLdIy6Gz+ST7
FS2egy0a/RYyT1OTMBkatfggdOCOtt8KmltYfZ1ySuFJDowt2m9zjDTSFgphjNX2p++onWaaaMAH
oCCyF4k4rdXdxWhvniYSqRn0/1VPHYjLMou9WoHa/qHmFX38fJFryEXZfLlDzqXpNmZtVU7/tX5z
s1tMgd9p6YGhdCvjMByoUYx2YqDja2drnYZAChpPXyVKZ0GA7yYmRA8gHUghHttXtnBEVH4OxzPP
XP/hZUh+2OIt+jWPyjbQJeHXfDBw8zvnSVI8pe2DkMSW85+IuadKuWPkV4QNVTs1wL/P9RnBUMEQ
S2WDBmwzK+PlJ/n96LSZ1K5KrzJP+NAViZJjHg/q36pnCxsuvlJLkOqZOE4iDc8JojNTEzKWLKmF
YOPEIpBJ2x0n9s5Gz5rfBAkIeUEIpgSbDUbWPzswbpXz/V5jE5auS3ixoUXvVPihTZpthHLq1bx+
y8kB5nz9zKIORzyHHK+z/YWm4Ro0g4GD+1fN20D+LN5ud0UUeB6P1JUKXdywGj3aHer9GQ0s/eDN
W8x6e1bgs2jNJCdTcSuYNzcbqS4pC8dVUKbmrJGkGoF6n3gcnGSTQwhosMK2mACFOPuqGiOgra8Z
jQOdzzBg7oGFxaKkkZHKGHZias1UFM5LmOaoE9o5kT1F0AC93Oml4j7w8TsqH8hoRgRZhZw77Smk
ePYdHtZ29RkZBrOMXHgwWKY02upBUhYTPb6QHS1dG1TVEfrMzJL+a8MqjGXyCHy/JGg549s0wNVo
ii6NJC9M9WFtN2OYIMAXFGb8mTQYr18YjJIgeLSGr5UAjAPRCGQXopvIB5wIroB59XQiKPwPxecq
9mhYp5SlIL7GPhYDxGaSXkfpxGPqEXnw/Bdi6RkwF3Px50oXKkJOgpT3DtkwEMVZxzIF1lSwlIZd
gCNHCK0E95v4Xk6lEeR0gRmpWCRKVodrWBSQIJ9HSXMi3tlRs//Y7DsFNWmYInNCpNBiITEg+K0i
ZtrK7qDlR/ZKvPKdrCCdNBlxZt20CRuzB82KzO6PI6ZEzic/f9sEYvRdvZ/f5fdd48SxRF7Ixw1z
woKw+jBf2hd7JhxTewzNP6x+cJVZyCIwWaBgyGpeHQTtOP1NrFMVHJo6WTxFIG7LzEDpPAFRZNC3
8J1GtWPwdrmX1ca9JWvccGPdvUTBk5HQgoCGLtCbpf673KbBPyEasYq61iXFwXi2+Cq+zfqV2r0d
2fFWUFk/bVKDPPcSJx7UDayP2Dmnvh+eRNuaoRtYPFa07NMzBSyozSlNpnLUgBuu6gOYn1OBf0Gg
ALT76hSdrAWGvHfVlrh+22Zs9+V7LD1xhH9+PldEC/j+m02LoR1z04ER+OrDBMPPmDYIbnLLlM7z
NLKLXjZDQUn/a6NiB7X0Ks8DmVYH6E3pL8pV8YFWYfVIOJlVhb7xQS16qLSNFhrXYOfmLJzgv+gg
1WJ4FzIqP43oK19cotKnoxk57JqdnF2SoM22xVBEN4c2lhHq0j2HAfJAcXQIFkuDIfXRdHVAKY5G
/2h9kVELJdm3FdukO+AD6bW39sRdRLjUbkRwbumKlZFF9grkNICV1II73kFiCgeCTWf7qy4lWjez
Gznx8Pgrq/ASPtXEXHiWF9wnCDtNM1/HipGVHPq0zWLyRFXozmLodqGFOIx7xZbbjUuU+ass8XNP
HFpZ5qvpqR++zwFBS5VSwoGO8Da8Vth1QhqcTYT//vMxti1cOA+A++/9fMz3W2hOA8b3Y3MqfSBz
sTtg/8MUt3MrsNZOts2YAYa/7XE5vw5K7g01Q6U+tB4j0QC5/1N8l9mtlrETJYeSVSb7Xmv036Jo
Xm4lhXysfPZc1mt/53je8EXAY9JYAn3wap8BkCppySnCQQg++DAUYpNgklF+1GQnoKZowcR/44Su
SK/A9yRUKMPKh1Nhd+jIHVhiPFsH9m4JlEp4oyaWtUcZyvFGBq6//wuB7UDizZCj5xRaxTffry7A
9KtrIoRn5tRMXmSm+JDUuj/UPLAqiVkAnJIDMw4l38xoaJkgcSqkhvRpMT5H8ARON1m8ym6VZ/oY
ZYzDeZxIEwhel9dYpK4R5tDTd8aaVy33TPdm0B7qO/oMF35enA080/7ljihs4gUFnFyyl3P7tV4z
2BEui2NWrk5uEieJTKsQjMQj2MOX1IDtwhtz9gscltNF0AlRuvWk6YpmIcKOYSiY3wzFfRKQIt4P
tOJdNk3PT1O6J+v5R2o9tHpL+W7YWr6gyN4cgj4l5aoftAA+ikLn9QV9yxvuzCcYgrpJxPvHE22x
ARV0MDt43+EdtjrUL8lgah23wjQKIVi6W4watp/vrpAoN04f5Mv0YwKikrfI0kOmzGGPdR5OmiGm
xAgQpsZZlio2Q1U4H6S4YykGFP26gqmfbmtO3mr1KJlyY4OvnJpNCaddsxRHR2kIJ2sWDLhgal7K
lBDGRfnzCObFE42ONA2dqsCJKa6FNobUW5O2MFZtM3aq1b6xy+aMsOUxXUYjq/O7UZY4XSHGkf8U
CcO4mxZiFF8buljXxhgYujXt0Zl46JyIz6Vk5yRVcAMSoqo6BcYn3ERNPOhNDlDi9CDA4c/6sBCM
Szmoo0asJYqDFG9NfOAr5eXQdJvT35IfrxmDDOSG0/ZWqqU3JKuybsNqa6Hs07tv2M9COnedKMMs
d6Z7S3ozvKcah4TR5ZtGny7onqwm/cL4FtqUPv5j9yrkuBtYHwRCc916k3YKtN4GNxC1TUSGhAAH
3v8XJYgpOM1JeAexVVmX8HVujKudsQrd9U6cI9BXEXjv30SU1Na8tRo0H41aXAs4u2RBh4AuytFe
IyPkxbqDAB7EfjH2jI/a8oiWXTnJvGGp5lO8DaNjeiMdIA33i3x3GgGpclOrtSpkvK3cXDkjvSfl
j7xo30OtctaUsdowB9GjPEthlkyzib7jmKxIWdmO1v9vhzeHVF3uPQNrfkWR+MixgkyH75834LQ/
dMl08hj5BpAp9eoy0YXul0fUZzbXM/raKdBHwCrNVYAggXUWbCoYqqoDswScqGitlbuU/PatWv0a
dYYVAS9cYXbIhmkGhXzNOseUQixUl/K+vr9AnF8us/5Ohg3h8+Fnhp2E9YxRAYTz5Ui6r9HqKC15
XkmRQWL/gs/f/jvI/WtM/Edv/Kpj0dmwu0DOy3QdrU9w07Ibn8F80xwL5CfjtSbVLKsYOQl4HB2S
YNtifw7BTpRt0k0s1IWGn29eFCM7afl6x3BNc3pR7X2iSwJ0MIY9xq33ZWnWIDg/vM91E52+CTjQ
3WwiZw3ERNwnzShryexyaLusTzmW6zY13ncckkyr5aoe02N5asS5YClVXBM51A2JmwGfUL3dJ/Ag
pVs/3T++KeSS4QIg5gYRe8NkpbteN7PK7sA6J3CmFV7y+n4ZLscih+XUu3cySzqqgZyHS31iY1sG
PBbGsQjplsAHIBCP/uDBXe3NEE3yEPSpEsz/BIwQUzadtTcz7DeAbOx1GKlOeBKbINc2/XaHndJo
lMeCChSSHqk5XVa4gfTYV0byRLvwNOUqrX1ZQiQl0BN3rnRALQib5DD0xC06OdR2UCPi1NbJu/eL
W2GJ/2lzXPLdUmUSkSU3TPZDFqaVXk8SGSyg2eb3cVnqUj4Uulo2h6tugdVHXv0LzOK/64TkKmU0
dy3yMXufzYmsYj+99Xflxx62eBq3OQtg1zwdBoS9PIFjuYYTy5e72M/toJvdrzUP0netd62G61Ip
wWKCPXeLInbwAsif3AZ4g1L46ioHseHx4Cs7QHduFGO38CnxPrClTrXuTWi7ZdATiAFVVVUrkeAY
iwMF4mFXi4z5z4iXBCr9is4pt80iP38ti17YL+/fwzeVB+4Lw28Qp9k7jFeD01t99eGT50geK/h5
p6/LnLyg2YNNRum4w8Aj7LDXNZ64HpI4zVedxZhTr0mzdAqzDYnXcVDsuxYITDOFcTwaFhQNDzYv
aXrrRgPU4EBpAzISjveoVrFx1SKTxrMSJYB+OUeFCfau1uqPtn/ypQKEJqi+H4tQI3vmCWSNO4zl
GnfCO4qRWkMVlY9OMMRIsN2+FizJAnhtdZ8ctetp4RhhFVePSskTETJ5UBvqXGFuTowJsda6HYj7
2kkWjLyfRPqjhCRvq5rbjAL05J78RADcGjZMRLLlttdQs+01poLBUKf4w/B6aQeXusbVfWfriTHo
F5PcF6gmEj6nWFfUQohvPdZbsnuAzpr0wkiz5D6RaGJ6W3fF4XqTmf1A0Rn1GE+dZH43PHotomnR
3RsKDIcRAHOIfZHyZwV1SbsIbX9UO5oajpQdNEoBdxM4AjhYX+4OjbJ/6Cgikei5uTAARyIDdwaH
i+vCyNtSpBjVC7ag9i/fj9j1BlaEbNw3FiEddq8n/ML6vss3Jeb4fIDADYqeKJlBvzaz4Ji700yC
jLjOcYG1AwuB+IGG3OdkPlowE34BgXzdC8S7pqPcbJLjcsAX6YsBbuV40oPkBjbgcrYW69s3xx+t
28eqUwJLx4JvMx6dTRBtBftq4ucAtrIhAcKDlUwg6PNy2eiZTgIWCOdFg1MmZEHGS34kDoq3pGhj
19pHCx0sNJOZfSdqP+FHmygjPGe/CB/LzuRsDTFd5Avn0rjznVAT/kwx+YQ0Sj2xurZiDzKpZVRR
g6jmVrUOitBSXfqpRDA5MnC8P/qkquXTuAtmcMA+DgrK3HMBbtDu3NjoA5ScADwPz3l4LIsyMzwH
mU/kpbxUQndq/SiT5rYC/iaY9VCrafPpzL+ksKzx7wYNxXnW56JT3iJ3RjTV1DI1nEveMfpmt+rn
ur7cY8qSJqDVxY+pOYFPe2uQPKkUUQZNGnltgMnvK+pJSM/7tAQNt9/KYR07bHCUc7/BIPABBbGw
O2BaqwkqEQUNMMiF4HKLiNxDtqhe5FR5FgyO1zLrzrRwoISYjEDxpfuWIrSlQsnka2GqODNgZsBF
ImL6Mnwb8FpQVjluFG9OXkPnIWXkfp4LTtTAaSsXslh+LrbwSlWRg1I4megDcqUdEb3Y/aCpaYmb
IVauHRixpo3xYorihWnCKDtyG5/VhoJifh4V4NfQFixNWZcVhL3MdQX9vQ8Z16gQLLBQz9BJFous
4f9mvjsPUUgeL7FyKUNz+pwkkaWQ3ohMhGRvrimM1P/tsNjxFlobMp2scJjvVZI6shkNxQby5PJv
WaYSOe6EXy+KTYN/ovn9v3m6k/36LNiKoiX9WX0UWFPNO8zc9SLA8oiWhFtXntjM91KQwcR+oDYF
o4NauGrBf25whhavgnHXlLpsg2J8VwyqVkl/Zn7tsf2upSSz3Te/ApTVnHhKcS/L8UozhcNFee2w
es0Xy/q1KIb6pfdXky53K9/BAy5N4G1y6hgymGp+aczwKi/rBSBpKpsB2438OT+qwvqozJa58t6+
PyyyhKgVgTXWha1J/ITORrA9/fNvVkQwwmE3g57P4FcItrBxB05bYzakG+Yt4eFfPgiKxsHZOO4Z
vQUm4Jqs5l04AqEokRBO6OYS0IDCJM2bYsEOUzvEAIay+ogOtu+YJT5xhIGT3MpsO9TPKwYsbvb2
gMOTqYlseuYGuvEUM7TsWUPs/yIRgrvybY1o5FtimascdT7xH0glVMTdxMXT1+h0VNP+r5KZVj/u
HK3KrlOmBHxd7UGiM2VpL5NG67Y5mIsVQf+gft4oiw/GFq/TtupZc6hIvBT7k+IFCytk1atdaQ2i
PXyQ8lkkpSg9xzlDWeR5nUdQAUNM/MBaGDImTJJIaYQP4LGIvaxE6y8KaIYqFeMX6AKH9+0MP7bL
YXU1jnOvnw3sSApbJignrBktNY1DQi3zmGarMIteTvPbn/5SK8t/O338h+zZBYE2GFIlImp6cQ+p
Zov3i8BXjK4JP3rZt30qF5W6kYRR6OsxcQIqNbWMrvG8zJTfPO0dMy6FIJZsJuQ/F/fxg3FSRhJ7
lgawUYOpixXdWuOg3j2UCBIk7OOBhjGxQ18YcUHlWFTub1T4LsAdiz5farPY4tedVva2OIdmRnVR
jzuN9MF8nl6nU7pNo+t+VFRUb4RE6Vu3/4uJPdX7pCu/zdiL1nDI8I1BBplpq67Rq3oF7hhfiDYt
oZlFZdVtaqPxzNXLg/6YWkmqRKKjvup9fTP3iiFJhdLS2rIZVL5EKEic+YjRwGzTj3TMjjNDyyHm
/2UUfNcuGLdWycKAvf/M74d/zlEHG3NH/Oz8y1/8ClcDTUDBkbGFHCAzyieUamUYH0j9mRmNuY0E
D9Lp3Qsdvb/RN3ghesGKjpbBmMk5z3e/+YhltMrUo6VSj7+fRv53J8oZSmw4raTxLZv5L1T/wF0u
Tz7uxFyK6bU4QfoAOp+6V/hfX4GNC1ICMjmdd3lDdKacg2bEOjBVsx6uFalkbNtiqMXUqJM0vwcL
ET4fT90EoJm+cdt/xTYR0O4yBQqwZmVOcF9pq3MpqUKUR9opVdhFJNrB0zUEa7pGTCwbH2kM/2A1
AMmKRu6ZSLLue9XnxFZux+J9NPWDwpFAdg0ZQjPrJtG6AvpVxLSNCZ5gJQeB0ytkf6VhBB0bFsFp
vJxwtbHDMJ7GcLIiMRdJzzoVKC9ctq4icnjgtkYyDbGcuLdygDQdyxoeurApKYfTYB/mHY4IaHT3
+Cvo/e/xwUnh8tokD+coz+8MCaTn8Ho0PyavsVc05T6vWP2Uv9UMS7jcwVC0crkMzKdpX5rk/c+w
Tp+2dU9gGUQNCZljqqcpmw2S7+U0lcGSvyS6QHVOvinrrgYIRrgtoVckfericAWgcoCB1G0bnayh
OleqTX9CVdq1qA3M7lMlMpPLMFRJWGhq6Oci/E8j9PjJHnWV/6i1acZttbULnOr0PSW8CdiKNFnb
/a7EWpCsnUntEjhXXZSNYLUuf4iib7P7IqNyCAPoLmJFx5mHnOLila2ICOMccrxiiP/iwp0ltqPU
E/WFMg005WLI5FbU0cU1OYxINXNOxn6LElTL4FnX8HLnNZM8ewupPYK01XxDjYMSABevpQiWbJ9x
YMxIl5ztoNdg8kI7VGWjXhBDLIUszpMQKhCL64TRaBatjyzGotT8YRRR62DV7JEJr/hN59WXyMaw
IyWguKH0xGpC0k7tqVW8zz2aP7N+T5CfIrYZPWcnMKNHwKN3T90LQ3ndC1oy565nIwYgSnwsITkF
3ZY+lEzWtgdas9+LnnAp3n183Wg/BM6ZWTosnZfIvWvXgYEQEhCKkhvjLqLzSTTAPFQPKze/Cy4i
371ByMeOznvlxzpv+lHkAOcsnefsPAw75s59ElNYbOibL5iiidxV+1ioDic53uIfb19Rg3xJXh9V
scyKvyiNnqg3rejrgt5SZYrkhb/OI9tB3k2YgG9WLx17SiBwIcX67UUlsk9k1wpwy9SQJ7rV5R5z
7QPpK+luMoszOkGkGfDq00dDadsmDulMiZFtYZhvCHO/xI8nWQAAYqSFJDedDpaU71sv8NGy/f6R
wu2WJ9WFaDZkDUQy7u1dHN6LPvIDmjYifGTCPr0J61RQs6HRWHE39OyKGFTLKEUrVNOc0dzfYEyV
tjlOGJgmhejRHBCI/AyEhP6eIbsXnmsgPuPsmKxzUxkn4rfYrTm81pEBqSquBKQMjr6YlRJ0YD3c
sWJKy3F0pJRupGAr1ZHEGnZx9NkIwIorHtltLBROkqBcN27KGN+lbVl0kFAb4s05ecNtjVZNPY3X
SBySw744OEZBF2K2LPI4WNxV0GVsj7NUss/W8Fji7zMl1XY02ZJdHFRLZUB04fSblW/6VyPPKeUb
VNobhtJffrawDkVmf/vZzzbYyrK/g1x0QKiIp+2kM6FFyePpQUVYjBsgK8WThNVr3Zv6GtLKU/+i
j0i16ex8bl05qEC3socf+sXTc7UKt42Et+VwBNksAy3PC7xEPNOiMHfhmlw4XkL0SoO9kNnYQqK0
lh3CeSYfpggHsvTEjrVjR1gd61vr+bQT4VLwjDVK5WR5JYHE6qC4b/65BxFVwCNQop2t2nAH5Ur8
gFntDNNinaIn/4ASllNbUTGW2op1CK1ma4Y2wJ6smvkPQcC+cVJeOMrvYGEAZZjXI4LhgS6AbUPe
3bB/6ktfV9yt84e26DpHx1yXuKzqiiwX0I+EteWNnW/uHk7zYxdIBWVsqtRj3aSFtSDm/ViCdO7n
PRpHroGFk+jiwPIzr9ftUrlI0CAz72JMcCil48mYV4hJV3E24c+1IBq71p80bT5pjo7r9d1OQlm/
De+Dnx85AlJh9AdrDw6Z8b1GKiH3tgGceOM/woSbXnc+J7KFO4CoOtJGoLoHuRafodXFnO4h6nPr
0YCt54tAjd1Q9TlWnDuzJIvzgyhB1yYH3YFXaJRKhu6sN5tE7fuqG1b3bo//QainFGZzSkojQFYB
uY/yFx90MPVyKUCZzqlvVxXbw/seLFMbr/NTPmQbT9NUNjkasRrctKnMZ6RBsgGFwa0jYWbb6d8L
f0VJ87u2IodR83DF0615XL4FA3r5OcTUGg6JnkNMCIJ49R2kjyNgfHfcPrfyz1z2fbbof2Ct56RP
7IQiqUcXAya2Z5Z+PyGbeKx63oJwHK7oXAelQ9bXVsPG/Lw+yFCfINIwLQ8rQuULSOVoVtV/F5U0
2/r1/8icWS1+ZBE+nU/6pEZ0KCVEXg4PwqIs2JPsM2lDbheNXOB9hMhS/KIXvSloLRfmCVuD3fp/
Q/OJHMhrgMhPOjXEHZdWL7p+M+OfDgxbgcvCQhcFzbi+bMDFQzKP7rJR4aPGpOB5S6VINU3xVJ3G
XIllWk+otFMnvni4UbeoeUGs/nabMGVfCGrnI+pj5xI6vNQVGCTT0vn+D5SxCTFjlrcNfMXt2nAR
jPf8Ri0Zxmk1x2u/459nbHlauMRAkA5u1hbuP4qZAOrPhfXN7yG5mOjspaN4UjDijjVQSeVSMTed
42r43XSHOlKQiz3g/8CY5PMEOi0k5iZZrEYtn9yM0Wj5V/gSzxLnE13M7MeBTCA/etzCb2fOnyU1
6/Z4twJip6rAINGzLJBHTiqdqPpG0v7yVih5CE5BzbhdbXs1o6N15cTlUshTkLV82JlF/I2fBdqA
wg0rKcD/0Y8WSsw00mTYiisjFIYNJya1o+ygGNKXaqkklP2iP+/CU19/rp1fsjC8oGsiat7z7zuH
7JNkYQFjEXQV2Dj5Sk0gwv2gPds27lt+mwGrTcQjTamvpQJjJY1S9xnKJ6YiZcI7vFUqGC3Y0H6N
8XrPX2FRSoUadeB4drCvn3MTAkx2d5nReSPSsMb2XTfRO/y5W7zwR2F1ayCUd3x3+fHxY5dTT2XC
Yx+23W6IZNP+OP6OUp5jMdqRSUxXVO7FTL8J+iEk3YnLafUs5ukCyY2HWzXVOCecRLPqI/wPFeob
GrJbJSgjb7FVyj6QmhvbW1CYEK5wEQCgRtZxNGUbCOyu+Mxsp7/cU19k5XhPqh2n4lu1/Dyy+fL2
3mwbFgTLm7DAdrWheA/yRkmRnExDN5vbBp3urjnTpJunZwirQjKhCJuUoOqqg8wtNpCCBdmPyAew
AwamJKzfmFyQCF/3fJc1fChZP4FjtA3kIo6bX5Y+oSW7uetjGcy4APQ34bpWlBq3xFcACMF6+nt7
40yuwSMJqcKctOPA/8vSCXuqPYkvJClJ9v1dwt33fMTg3bBTP5zMswaC3SQnTQFcB1H9aChJ4+QV
utUzBTyQli6nEF31a5TrfZufv0396H4IrJBbKN3IfzCeP2Qga2LjwklBdhfb6BaX9j5PdtgaHBpS
AUyed6lIwr3We9dhgZ4xZ+GgTMMksasi40vTlLW/mLzJC5/CRIR8wZA4DHIzzZTvhY+W4oTmpVDn
OlOLF0SzPTMnTZlHIVY/m00hu85RxFMdQfEEkdzSJ0rvxWV0e129rN3ailcXVqniRf4KLem/Ox5e
oyAc0kB1xcpQtic/FXwy8fzfLeZrVV0I60yANPMIQnv0o9XaMT/Q+COrwE8U2VTyfXddJkHSCNyQ
D4UdxbzyCKkabWWk0N4JPrKVsWRJHKYwyoQdnB5sDnpg0yk3TBuR6jB98s9zELhleJLfp5gwn9Cw
7cg4VyzNSlv6TizQvURt9AOy6Fmi0C0Vah7GSKRzBT9AsZabfCrqnacGdGeSwlUP/xyrQjifhvCE
iYr6Urj8m2BH7WoufDKy0nUyw/OAXpvUUzfXCFMa15lTUub820q8cTRu0vxzUqrAybK/lY6lwczg
jwIawH584jYp2bsSSpFn1THPZ1ASvLzF3xuznqY3z/glkyQq4Elx8yVqR7N0GdrqImDmq2PUJ7Ye
UGQ+TSLUFJ667k9MN42zxNfBTOKtevUwzi6jsikLWLo0CW3U0mNKoUG+iE+ON66ClYwYeqL264qW
lg2zEkgkUIv4mFJ5PyamgF1+hw1h3czzyyV4d0V2gTWeu6LIJiYMiLPP3EJn9DQPWF7/nnkrJtsY
je6wQJnmEuIdyHRHCQs97QIIuBYBNEis8Wh6wsqax449RwwmqIPufIMp+a+eK9TsBAWhmbNVpreP
0nwP1OujjQw5JbMZW5PuaUKK+kF63Qcm6L3gwGOcgV5njsnWeDgjNa6bbTgHipGFQChlIb+cs2ey
njRUewvpuiNKTMb3xS8+MVaUlbJwSbOa16MnXv7d/Cs7CrbC6KPYAc+HSvZthTJfQgxYyUgOyuD5
48InmpWRB0+cpuB804Z2I9kxI6bOnpe7ecOTVWbmcL86kTJ1Vo5bT/KwfNEo1AUGt1vxT0wuf9Ye
lxz7R6XagDZAeJfD6cFeB8jKUerV64zepEZ0WkEmZIfwKEt+h85smz+/EB79ZJpgW8G51l0zfND8
IJCxL03Lu7pUJxkThJ5EL49ZtvRxQWR9ODYaf3sVJ9YgDtqU8oda6pQFv1vSAzp6koFjTPopxm1Z
CxRZMtuYl1/YPdAbt/NoLgpmxoH3/xaLqMtNsGJO6BVhagESy8f5I3aZo/y+jH2xaPyXn4LK9hoj
plGmcUyZDQ4KXf2gZ717V/ykSDoFtwCBXuhA7oemnV7QdCKnMxjO22z1pxjHgX+7NvchdGax/w/i
Qx2Q2j+roqy51I2QXRdOq8O9SA9eD43VKkr2RuqFaUBmDL35x8lGG33hFSjeXKlitgABrX3Yuw7B
tKgp/OUuKNUCzj8BLFt5uPV3Zm+dyhEFNezDaa/kV4WRrRxXqeRyvItdc3wptsx8GD2Y7+3sd6b0
KviaS6zycW0Yqj701F4kV/1t68LcUjq7+z6uRPI7XPnnLvLG6brjxp8cT41+NC1Uyvv98EnX1+Ia
CsPejbG7K1qQhyJobQS2BGMnIHEJPC/ZvzBp54ckFlWQwGno4c6RRgaFc1W/6RrqLfahMy1EbKCc
T+NPiGLazdyGVx3tKtGLnS3N4IIpDxNjbF+UoD3C5QAjusO77S6Xiglocmy5c0ZcydgiDkkqkHIX
0N3Z0lN7+RofmSR2PD2nslfRgtXHL/5PFS/sobyakaqk+lKbdMpnC9MESwc7VAGUIpOumj5I/Bfp
63JxpCvDCrfwAulvOTPDWuzphMIM6R1hPiDJAeal24wnFHGHmb2Z2X0s7UC7DvdTDcPBsLgpWnRa
kneTZScqUFtPakVGz9Ch/k7Wgrn5AdCp9IlsbydcXwp2A7j2HVvEeoFkEYhfGH5qMrcLE7wEhGuc
GZzxxzmIDE9QOwnGYxEPCf+u1VlC38DPLg7dJCQABEWO97Mf5tYy1L12BtJBTtsmVYcjZ7B0JJRA
YZ+5orba8rInl0DkfmQeDymao3lRZNPMklBdiqpGPiArmBYPfL5yQavy+sATfWa7R2LmxMYDK8CP
QHkexUEa0B6Gh6ZNeM3sDRdCVJUnuXdU3CLqWq0ap46dTTOMdGhQi7jCnxAM2Hi8VnhhMqnLDUjk
lOjxiNaWqA5zwikg9HnDbOZB35/IeWEcsnDW5VoKqw44ifQHBTl7DWQLbcr82lEBF2xfddqOmBAJ
VaiUxb5nMvaWxTSu9vmLRlH1c7j/nS6QkXVwZrR3FFkn+Gg5ydBsdD93KrxT3LAuPNjQtDZh7dHW
y7JhpJbHJ81TpKh3afMO9GxSau9xh2x8SxuZ3ecdnwWvhtxZ9Tsb5O5CFEyFnjfCuAY1RM/3Jf20
camjT0KaOGIAZkDmay4bAxAd4Z4xDmnepyL2vyAOov5JlCd1c3SL3xlyagoT4fJAlEr0EWNBoeNz
z9t4oSfFzV4FVRbSVsnyMSwaZyZs27/S38dPp7feJlpYWjSndzNcb/3uZ64na2XO146bzApzDpWk
DvlryugAm/9c4Nt8Xc6ocT5BE5VBf5odCM/i5hCk3JkxH6V0CB3wSGb0uxFu2US+Jaqxk6vVTO9l
G9OddRoSKzBNeLg40RNraFcEhQVcZ3nQUUbvdg+vdEtZza0TaUWU7aZvg+M/Uy2VvN1PMkMaEMTC
7nBtwPutesd9pMDcGRbMAqneJVAMAeAobzsVbkjqvF8whPpfbBCmxecmFSDDc0rYNzkeFqS3xYb6
2tmViRRiPfssdUJGxMssNq6KzeRIlpuLjdP5yIxjywc+xS2qiPIMjqd7P+0NcrTl53N4VKurq/0n
o+d5aOPYDefiINn5GaPZmp0MboX7YkGlA9tyi77vA/5QVb8mUXLQY8eXdEXQ2t/GTqw8OMr5rkc7
mdcjqPPftkFF2VoCNPgGX1mNIqKSWAT7bsSjuLDofBOydhGuUZZ9qjP2yQkkSq3lykfBHPe2FQ3Y
NP/s5RrXlQtHdJBDkxYh0fFoRRvxD1rhNe2CTNvsBmjVWZiLVnVdwqpns2hrl6xsrKUyxkvP0fm3
nuMfdV7w6QQThcNrrtONPGx+ujqrXKHEDT8ZK/RbxxwyNOH78T8j+x3yezDqCeWVMWwqynEuyi2M
otaNkHdVjRgkguLc5Y4AI3oro9EH9wRLofVTwxwogymCY3qr10zI4mF7ezgsYVykOdi64Ue5sI4v
YQe+SlzdTmtS4EqDXbVpLC+vCAfDhBC49ACFYKMQgKNc7eQ9De7Lwf1ywdTqtl/ZOs6cbIWVt5JB
LrzIfWyDQ4baMxvFg8TTGDDNfp3s1a+ZG0K5j/mo5OXUSvzVd/b13xmiwolMvcex2CdKsJ9YxmyK
m5eSqpggkT0sotHJVWXNajupaVsMXE+e1tb3xFsrql3+gS90pozcDPzqLNTvejaFG1fFHy8GPNBM
FUzh8+ST1fUW/AjXsUiSOkK4a5k2pIMAIIILGC6ffEXKwExnwgO8UmR/RzCO5g5ZecScUKVHOJnU
X/CUC0EO8rYB8/ENpqPmUTYVczyns7iQNDKoMlT6jhVl3ecVUZhIotuAoW+r2urmDHG/1ynVBb2V
m/RteHehM4/KC2xuh35fFkUPN003xBnAbyPFfoXT8ZC/tEEXm5aU/fwjobcHyNOqsiKfjmHR2ipt
jio6i9KlhY+IImmfcbGnPPSrlCCGCp8Ab5V+F6gLGglg+q4EgIxxH1t3xBm7wjQ4eyAxp+NSQCwz
sAghD4BHt8EW+FNEj3nh02Fpp4Ei5d0M7mCO/wzDdykO6GEAoCc/bKdIW7c9zeDmvUhAmDpCx0W3
w4VvVWigHJ0Py2/WyikbHSDKvrDRKniJQ8GYxbO6HR7YQ1SJS62pGq/XQnpp1s6366MIn1un+KhR
HukavHwMTCjEi7k1XSjM84c17j9ga6PouIXQDiOQke0ug763Y/WbjOGMV09DnqS+WfN74d8wMgMQ
qlbcvg/zFLPEchU+eAbvxxfW6pzBqEGsjV0tcmmDAKhG6Lj+YZCapT921vc67eY0OR/zbTeJapPG
GECWS5x7Lb5Q3H/Zc2sIwSHwMUPJwxjMZOOFzZHMzJEP0TiNaQ32hRCGfz9RHEVqaPxX0q18AeWv
KDVc8TuVOm2qJlRulQ9TNmP2VCaDtiDOMkren3Fwy+YvII3Pr+D4loNjm1vlsW7Oo/7rXArkAJ9b
qlWylEYjbQDEjh1hN3Y1cW9yOzosvMgoDXz/dx0uVN4duB6Y7SVCuIxkESwyRjCD4SWo7LVw/T5g
waDOsLZrY+NCN5I1g3WzAO346yXoQF0T27OFk5bqZ9T+sGnnBpM+QjlCRN6GQfL4fg+3w8TCWAcH
xgSBlF4kY+Iu0CiCDqZpYAfE78KD4aZLp3copBZtqWWbbXKgYTWZxgCmg21SVuNMUV1e8gHiS9XL
WiKUe4x5ONciYz65I0jDDuG3mNN75i40r5XToMu45kZ95elGFwsx/MqiAeJMTbbFYHWPeuovnidg
5vvanLQzF5iglc+qUXuZ81mwPq+LhzC3DGVMXX5D/jYRpJ7vEPKSsikfA8FL7RurdhPicNbRTfEN
SLfcgY9oTFD7HfhMb1nSvq3eD7uegOOoXytgdLGbrwSNFi+7fnvg99BUPzWzD4ff4zu9+tSGq9dW
aDpcd4DUoTkV9pzASFjnjXZO19f+gAbNFJbYdBWTqTWR8p2uia4n0PkcbtGsG+5p8BMBADhs8eDd
ys8QaIx/zV+MHHssrk73CqmSK3bZMBXRUo3eynDMml8wTjVTHI9o+Mk4KgS95lVaC/pK/Cskxtf5
KLXBED1WxilnPJdAjz5C1S0usdsHdp38ekZ+hxz4IRFCeuTmxusBdr6ZBn2fxmr7SqALSb79LLuW
zyZRCVDqlVyHn57r/YRNBYeECp9hnb2PyCAmrk7aiOnWCIA4eKlUvnAILnQJvJpGBpp8Kh7+O6o2
ToQHXMQYVOoZSllVjrTBCfUN+49vQQH8rcCD2xKvt5P4ParWJYFJBDYmgrDNEWEYfHm8bonfLl7u
ECrexq/fyapI5QEOUSfp9xAc8w6Lp/xDEZyzmFQmbTAYlkQfPJMGnDDk9nBQPAtq/oQRcwo8YRyR
y1j2VvuOuBDjDfY8ptY06R1B3bi9n4gvkIC7i5EcAP8X6GnoSXzrD5huWqdbXx/aL38lgWF8j8Mm
ur/gbjqsrxkllT23nCM38vNn7cEedGbHpk9yN07wZyBvOVNJG1PKGD0HG+f7JMs0cYnenYsLMbhW
8tAlI7/6n/6EaL2wC9suG6G0bcjtuJxbVmEHnNQJlYcDbO3EDTUlo1O0oAMA6fnUv2j/ZPBa5u+v
E6T2hzgSKHbu/czfsCn+2WTrJH+X6jTeR/WTDXVlgcrz/rfScvDGv9CPH5ATgflXyIfjtYQPIGjE
1vKrdQ49Ne6BRLe4G1OTLTYx/Jnuav2rJz0wL3DH9erdHhLPpXbLmAvITDcL0nMVNSGvWUWqLOvH
+x3tbUEs3ODbCcgly7ZCB0x8SI9HkCjwC6z+6GSCibF48TTr59OVJ9MUwGeDF3zYD9a59GkAffp3
Rx8uHuPYXo8D73sAdms0uMRGelVdIgV5hvWMy0uDI9XKLKehHOY7m55AW35e7ng9qVy65vLswxvq
+PXNLyHg+V1BPXwsHDLlo4u3Q8oP7ZtH+FLLICb+VtgKiFcPG5tygifbgCkTeuVnZMMDGW3Z9z9I
Z0xDImDK2lwj/RvW4hiyNW9EhZv97BLh5/IdVxhiP9mUAFCK54x5/fO1A+2l62FEgnjEXbEiWMFb
sueyx+uoQqw81X0T7nq/bCPndhn+79zABMSQHEXkLE1uRADvqi/3HCh5U8rSKazBijmt1QkJI9bV
haWY5ybQP5CxnLrSWBdkE3VvQgms7+83ywWVBdhnNvo0eNDLoNVfHwWPe8BXFzIqJv3FV9/abcUN
olRYFxM6+PlfgiNDW9GIDF6mo0ZgVwGpZ5bAp6cwpxhkW9ZwdorpLy0z0tPl0/zLXIzbfginw3f/
+eq+OGMFnI8soVJR1n9Mj+CFAOrC47kZRClX56SnOWdPmHfuQEj9dFoGsONJ/HNHGc5z9i+3GZlP
X4RHFFsHQuxVtYpxWwYowUEz/rGKvo7nTxdRZIESqaLIVFUe7QI+p+w8mVlEZgIk5HGZENdwE8K1
CVfCdZ0su7qViEJ9JZobw2Q+jTN1Ay7fJFfEWe91UuJox9WiuK/3EtoTj3C2tV/MIdciCGZvlt+L
i77iylLe0x7cUlDa6OLRco6TvmJf4bXMD7OvjjSaRmlAPBefK7ncROuMOV/Ln/r05x0YU3HbiAEx
RbXZlj29B7WmRlG2hfqSmtUwxLPy6eQM2AOoFhQwlHrV61+SGX+D/ciEgJgJM8pezEqDqFNW+y86
HOdSN/syzKSBf5iLHe1djjLyUhox8zCTI0oixlbsEv9pHFDp/gQJLM0jGoqUz5/J1KnNzMm230F+
eVgoy9OvUZfAp8zJz4ZFWh2LRYIf+yulwNLc5wuIEe5fGx/eWcIa1f7Vjps3yJjspVchgay1SCSt
nrzOTLQG2aE0CNvepaVKx2fNy6vCo9gQaT/F0CN+MpNcOHquvvgF4jLl0Uk86uNwUqBzUQzxTZWq
Wdg8A/tPFhgpgIkGxDmbaJYW3IjXBc1/4SP/nTPFIqb34vkZpf5eaLbpFEvFE6vaQ8QY97HHPygn
C22M3+hYF7cwGip01Mf/0uDfsX9ZqV9xb23MxIRwMKODIA8me+wYlrOiOaitN8jiD/HwdhyGsksQ
fFlImfZKGLPBdr09F/dajJt6yb8eSQw5t8T+izAzvraUmNuRz5zNrCLqpGtOQuoPTz/hXRk57SR5
6CXDsBVNapQ8ocgktKc/Weu8m6wL6P8RM+++udegJCuI7owm2q2Cze2m4gFnMq5XJ+81VTo/5OXP
N3FDiKX6tXHAGTu7/Et3ufxpqQRZdclhFeOjQToJCzKdf5/tozQL0D1XypwDfZjR6R3XwpiTj5P9
c92c7iaIVJ/BPN1J2DGy/UIsb7twgEUPlHCRcVspsk8dwOIePScBna6rXJBHLsBIll/xlyKAQ0jf
sGC0MBkgxnyhvlnsyh1tVpuJG5SfK0IlEK39/MBIx1roLr6zTlbveWNsmhipQGNXmBGUz/55hsxH
jSZjtr1mbd0RqwYxSTo8QZUIy+BUyDbOn2PosfTIm1/zoMzj3M3CzJwr0WnhoYKwtU/J10f+E76s
VDHGKqdF/mJGn53BCkjL/x36/gOzja+LECW7kyDFbfeyZrgHInzbCOubGPrul/EDENTCaMTQPVRh
4Z23zIkx75KMCOhyZqwTI5IGApDyhJBQP45EhOhx4FpuFBUMVZRLTZW9fBMJFK8SXA9pT5717LlD
4frD1SsGe9Hb2EQLgDYLXIShCLp2yiL7NyP60I6Lc7bpJLH5PMw/SZqky59KrNaO3LCunOv5RBo5
JHg+J9ozOEcKYztTg3llC2ZUnD7RaUn7BNgkiBo2+aLtpeU0IzW/H8zFH7GohJm+Iv7gYz1MvfeQ
lm0MyaClQzCIWPdWGpbh+xIxZbOWDjICQLDcTK5hr906taBEJGrmS3Mg4sNaZLcS56MTMp/CDslG
Y0xnnZW6wBRBQa/3xTsD8dcGGTqobibDLZGOp5yBo/cGpsBmahln9yHZzmIgUyj+9g8/NdYW5HY8
NEv+QLLZsUAl24D7SbnwwOTnzib+F4hxUZbMhFy3JV1elesDDhJv4uAazVjhmTNqpQk0Naj7yhqu
fkveRhz4/9crXACHEGVDBkxadYMKsGFDnzm4XSeTazbUAbIC+VjtRG5EPR3tL5o4bv9sd9RHKL+/
F9NTFa8N6+t1DWHRFFvVANfabA29G3v8aLK2iHBxuuMIm9GhU4Mn3FZpP1Ubj1q/12DFvRhxkxGK
kgYu3pGHz4lxRXK8A9Bm2OJdKOJJwGHlO5bWdvhTGQrZQ2k7/Hj2S5jNSzytn0Fr0OQdJRxZFdIE
y15vqcI+VQMafa3AakwJM1gZJKBSyN+uW2MZhM8IWEiVYwYuhSnwQ+nncLN0P9tZQtW0R2A2vU79
TQXXzKzXOIrUcmvlu73D4sCuHihdFeLYHQ2qVlA1l5xSgAT2QuvHCdiHyTp8YH8KxudV6TkHvoEB
qN2zwdCSKTHWAVHENQwkTbrwFA9/yCETxEgZPHe9QPiiHY3Zj00sND8YdRJWXKND46lQh4bnJ6tr
IcqYpWHv8af37/KWeYhboBtOcMLehPgLSqs/S/3fyQfHYkVrY7NOzms9rgcpj+9xdPdkOtqdBI8o
obzZD39LXPmhwsFfAv4JL4e1dM+VoQpMTO98rZWWtQNx0lT7he1JS9nnaBeJST536atzH3oR0LHN
nfAr2ohkHEO87MF60LkQ8PXbx3Nqv5pyTnV+kx7Sje3m3I5cWfqhHYuUMSZ4jfcNZpXan/DKTP+Z
T+N8YTWpyhLWHvQGQIKZtTakKPRBmV0TAit5kDpy3QhzCnJHoW6Y9EFTPWRBqf8hU5/OODNZo1SJ
dn/dwATibtuvIm74A7oyvh1104/DHWS+a8RflVDhZy3/T6Cd/9IjynpUujmU7pe9sDQbPPOxWP7I
YQ6VaVf/W7Sx7SvT6sNxl2sLUgfOPifHuB7wrlNIjWb9BmsJVtTbcs6fvwyvfszVE5HLZzJinI3N
q0oyivCj+ABxSR9NRWiswy/1Ga50nZ5Yof84n2X3s2yzZWw13FzwkNyi1luW7LNYsiLf+ILExB6L
Mb6ChH6C2QQRC+WAGhdAh7enFSOldz5oLieCBdBVMkVYDsZ6FlFW5B4J+CJjAkKS1DARQwMTSIXj
7bkwf2OZfpScYaUI5PhnfwcoWQdhZbumG8Q1+Wzz6Y8QjwxtfLrkT4yXrHuSM+L2B3kC07rhjRs/
kQl6Iz2U6iJJUYN5D8R0EcgCtFRWCw+flklsXQuY9lv7bX3sUzLureXqJaO+JeO4ZuphhGNLtgBn
eCflc633whjvx46ZOwmX49MbnS5PFHORW3le5UwF/kTHwKbOp3WFFHbjoj3okdYZA4Uigc+jz+cT
qm3qgvOmiWZLPOTfoyus6EVFACZyK60gwhbjDTYZ2irDBLdBYUrTtcu82OmhfVG+Bo139wzUcSZS
RChQWASqJlLl5ddAIsBHyak8weknJ8FeFrtcT2YTcZoML/m3DJ9/ixxx3/4Jnh38uKF31Ic1BG8B
HBwK3l/xrJ7Oa8KarZrktoILUHnLrZTCc5BiYX5ISOMWZLTh83hskTqXpCTZY8aUuiStnARu/kju
SJkEU4gnENq9SIpEouYCT1NlHnWglQKZcDYvDPOZFBMEiKuT0SaIt9kJbSgJHsFyw0BxrHlSQF7Z
Gzq0kf8oG0Pm2r50uF3xgymOl+frg8CfuF2v5QBR42QsiD0J7rSMw5VqKyDci8vIRxNZtIcoQxxN
RRTBECVol5eDvncnkgzYgcsRL9DTU0LHeFkh5t5RdDtiZLiMmKZ6J5QP9xC5ZwS3jqFrH37PrZR3
hJximdlE+Dab00BfRTPoJEhqXwypyKeq7Ji8qs7LDAi+hhQM+exWqXI+pKpGGs0W2qcQe22M3pXH
H0fq0SSqEJ+KKB5o2UNncYjtzuzfh+36iHh4bC/i5Hgkyjt8/4wjPWZdg9gFUKwoSONKUOcg8r4O
SM48Mqqs94j2/+HLEbnrY69eq+Y/mSnYXROkoXSnBzSbGn2ax73IuSdptDVorxW7hF2dv3FRHNii
uLOeHmPlDrq6n+P+iiC2zvDVDxR6lwKp5FcpyNMYkD8yqpCpmdroQMD9iVaFcW6NU3X5wTLl+A4v
DkuuDtcASGhvbpQ5sLnrypEvGb1I/ECWIw/2d6B4wnfDlLc51OkD3m/xMBv+5ETkx/06LTCGU+1J
zPkf1BTir4a1KYXewcnZZ0Z/5HCEbNR1srLBZZpO5NABY9G8j5wPuSYuO3MKArYHuj2TkNhpQ/QV
P1AsSNG19ZXFZZYfdjf8ym4XRwQLEHuyHMKelZGQB37RgPZMRfgWX4GhGdimQxS+cqksMlXijjUp
D+PuJRm9s2fRcyghbO2d3iZXbvUdVMC7L2IoqNtxseOCwjXWWiplZOppuEC3GrUXEwOfdGPY6pJ2
VfySspt3hPbRk/PIIxPqHvyAtPgxjrOHROI0+Kq/SNMoQ7IbM7LV+Pucr0+L3VfBO2hLHAX3Arct
comKV5eei762djk7QzybD0873nBXTJ45SEGLpIDCehXN0iFBTA1iyUZXHktSIDESPzjlTdBrZiP4
tO8OimApHS03OBGbx5YpU0Cekkqcl2g+rMAAq1PkuxMVxlM2owo80lv6dabkrWK+iVIBaASQV2/o
ZXYZxMc88RS0JJLJ6AhsoLtROSBeF/YFdvWHU8NG1yNBbTe1nUJLSkCHXaKiheGx5r/+YGRXIkbT
9vET3YRJjdcN+DHsADUuHGO8dKEbYsKdb9IIrP7eUex/8CvzV6jJsIScChRcwPGa27yGPaWInLzx
zYRvpSzVFfeBNM8UEhJdAE+stp0sClqCSlPgyi/gTDgQZD1VWN7QsD2rtUu22cJfq2ObmPxaaEpR
r9faPHWCjAKieRYG8UZAx1yBMhcT0gzCcOa0EXxBqzrNS+2qfMzthcGl1U2IwOQV3x5j9iGHeTXw
dv1MxyYvgGGxex+m5Kes/EHbyS5dcYm7cFDhHu3pzq8WtsVjw39a6oH1pL8ddiU1jYbI2e1mUzuA
a3UW82+vq/4kD7KUI9/Qfax2dmlBBvi4CQHKFxLXxd9/h4ESS00gsdWY2Wlb93CL1fli4DY+ubr4
McizO/tADxbif14h6lG4kYbDxdJ8NydZCOoD+4CdHuy7KNABi4eel/GamuTOsty+0zOu1Nh6+ISR
36ezXo97FxcyH/b54ECgfeI53UpW/RmQd1xisl51uwpOsdkXsSy1uXT2JzsVQ88fXufoOt6qzGV+
NMLh3cekaEo8vpIkfOLtApJjkVb9Xz4qXPa5kbI0VVrFj1nGanIwfEfSj7hKVkXDUrt9VzimDexq
g2ylfWzil/pvjmLMOjmURh8BAVR5HoQLhEbGUXMqctOW6gxHxqT2GrkLqtxozeB1CWU/5QpZCZCC
IAstxY5J3B9KynBfj0RPZeBipnmEGbAfDJwdO+feAAFWenLxIBk+MR5J2G3OPGIqrvV7/I1uKEEv
UmlNNByKIidFAKsBGWa31O80z+HO+RHJpMv2EdOUlerjN/wwNETckbjnrkKKkH/3gjifpIBZugxU
r7NfO006gWmOPnsXbxbCS5i5ooJZpXi66ljgjTWJFzHlZbP/u58cga+Mzffqm1l0HUgxe8vm0j0I
DNTJJH/wQeo1rYikze0Zm/Hb6wGq/fx/DkQeBxoKifx/y+fLXFbYafK4Q+tarVQ9/QEopLjsbmya
NFhYA43J98LJos1vXRN/7kiuZEglUKLe6rk6jo9PbxM7ogRtNJGYX5/RE38s+yW+W1IZ2gMjT3/U
r1dDiJt5/b5D5kRgLYPS6yh/DHiyhV9dppsvxNACP0pBXE1P1S1B4TkfKK/nBl+5XR6y+9F+LaNk
TDy463IBvoq3FaVUs28G3Shw+dgQC7do8gZx8xtm/LKjH/eRF+RWvlQLTvz2fZidwYqivtN09who
OJxdgTAw3JOzXwr/Fv3quT0pI2LHyoWgHeZkgIeEONwfV37FQLgDLVfzpkwfQ72Y4yZbxe2lYG6z
6qS5iGBxrckdULkYX73nTphb7qcz1kL2h61QMFW9ay5yRIMD/6lBwPEzrIBVKZl2dGtEVGqjSfR1
B4H2LgW+ccfNBH3w+OxKRz1voKG0yvPhdFT+V+BUoc24jwTCP+42yUMvw/GKu2cXFXwYIKhC21QQ
ZgSsttVUfHmFR67fvdl8MEKJJmwPgefjH+QtOG3QxFmJAjjiwc2k9TCHnT21F3kQ/SD6bDyvXtm2
lD10EmaYWOINKeTiukXW5zmvmcBMIDB2QRa+kHmJoZ4QtsVTQxW98eqLujgDk4tSIcaiv0g4zE6Z
fQz8N2n9O/+AZSvJGinOqjr6uhUH0ia+ug5nY4O1sCIb4UI5tw/f4kKPQsevd4sIe7rhHZzzkDzS
f73Ww9pTBD+9I+5+3pLe/8vLXSQcpIEYsPDT8RYR/jWqfyBd9lBk9DPS3Qb+1tn0eGiGUji3ul8L
Bf2MqbOYGdhAxVyQJeGEZcoYqshuCJZ5T4P+YJfCh5QN8a2whjxbQZKLpyiofZgzyHWPSfhv9amv
sKZp0HDZf07r/IhEA4GOldnuEEUF6cLgPPfxad8NQ4Zx3aeVJQ2fWYKVxFPPr3gyX2OAWdU84Vbr
H+2V7iyomFW6+UXli8Uk2aLRpTKHhohAsmruZYISgRU7F+9NOEbtQaAuyOQBh8iILL53v0j//FGj
FBBVCv+7nzQTv0Lc8bEddf7SOnh4Nc/SNxmBoeJAPrpC3/2WBlNB3RMTkrvSwpflWZcL1AfwdWu+
VvM8IL11OvRviVdO+N1RqG+C7uK+WWeJ64KT5j0sa5bH1mecLPYQq59x3R8hlCxZrWXgRaSINmn2
/UXUaq/JXrgO404DC4MpdWXpxwGhoYtZhKQ/WVClYfF6cocYKIoM0XPq9TMz38EXczQPLnbPx+iJ
zEr0CnrMD1rTXS7HPId6mCj/LSPJq3JmYxh0pmof58Ri/hcVM7tk/aigFEdGFnaZLM9V5Kmj82sD
Ms7AtIQb7oudVdlcvAvxWOHgZXBio6V5hPBQ6QYdheyLxpw4PWiILrj2chJtRA9mzXWlG0f+/HaZ
eOnbEly27OpyBXgk5yjFuGcyJk3Hn+64Nhe0fr52G4yH5mLbvEB7YXPtMZrZ6Hh7xn+yQ31m1f1o
PMzlneUkliQiPe7SxBQH6jMBnSo80qxIzfluLleh1GD2/SHRXWDb6Vl2FsK/CJUlSgMD8eFU9Oyn
/MQoeiTdyDMps+Jn57QdZFv0iq2ZlJXsHcKv0e7rPZCIplJYWWrZ85qD6Z5T/YTqJrhb9jwSZwsH
1dcF/iLvxQURuOAMRRd2Aphscdt4niOmUxvH4avAnX2Id0BCr+E+r9UYI1JLmcbHv/n+zcFTJaWf
yc0t4DqM1DhZ4NLJt5hVXeeU1KQFT1Ov9CjYUIFctuhXBCuvCcdxarrRubCS67qkE+FYY5CeakN8
LJQywYLlcNgWFXh+BrcZ7uxk2xJYm2TQOb+QPTmCysU3Y9ss7aIcjMowRNjxef3TQL3FjfW+RMvG
6mwAXdRBzVTDfMB4OvCNIEWAxsdVbtc8fH/kLe2eFqkKCxV3ag1PHrNg7/tGzappPCW/yMP35d46
iGqUBDYkpotO/y3Y5cXEyUEdY6+YIMvRMiD9Eg8sesMwCOs+p1Vo5+12PG2djRRvO7yYjR83hqiJ
2LSlZomD6Td7VdZqeFwN+b0zqEEcbJxVVm09jUcJOQJEiemTdnTsz4CiZd4trzgArYs9fFYGx6Sa
WTC4auWcZTaZSlNusYD9ikZ155HZxW1Cak7Oh3Mdvh6EjztYip8UtDe2P1s2UHLR7IKPQXHipeWp
tbIyu7QQlsaLoYGD4YPokJPOLkweaia5RWeVDZYcwdVy/DXqJPMAKBftxJsCInkgrc1WdiTCyObv
Pt7bKV17XlT3aDAaPmknWyK0KtESZZsq6/cdvFEew0NdwtgkvguZR33coKKZ5mAwFekBMwYYYpSe
RfgtGHDCyu3KwkPOfgXEwilzh5XcO4p+kPn3QLX4QJBPOldQnZCPUFDOTMZW1XOyP3o4Xn+QdNha
QT9vCbcqSEBbaJEoR5v+lEnfgR8S8AzqxK+uewWcCmoih7tW+jo7F26waFPdHMjR8axLqVwQOlPF
sDsPc9u4wnPeYKIh5pHSeA9OLjk/VpAYWdo813MEzy/OJrb/EXttgcQbOUeTAPkr3+Sr++TPc6wo
5z0/u+Nzd3P7ghGy7Mj5YUw3S2wmDDYWk1DqsI/+NI4o5pBbmHgq3+t/T6PMwJMYyDXORm+I4Sz1
3fJ52/Ja2CJ+xpyfvQSdyDYOi6TgimJokIj/bgTxeIdswAEGt6SSIu+us+ooKheT4fbfggWLus2O
O2vll9DfMr5qbxEYSARgFrB0UqZmP4VhhS6o4iOonhCpJqznAWcogUSMFci3Dz7EqgEcT1uks/x+
E0Y4P2V4BbwjZdaEVkHWQ4P/fwEUkYKH24kuG+heg3AgcZkqjFHAXxPM7mf3DrOy7ZumV8VuExsY
1hlXtG2rDUB6F6z2O9VdRSlGeay0dlBrJKgFPjLXJ+gEKsuPlIbWSas0Q+t4QHkwf5Fg8MMJ3Hye
BY7ypm+/3mR9xbQrgSxK26dKuoHWz1BUd19ddVdoXaw6/i+AxpYu/ivHy4PXslidtsx+YgkflcVp
H9RtcBdp5+J7aQRpYbbJElIBrtIvChDVQwUgp6UNe6WTVapK7Kp8MX7zISrkxGxbVggLfxGlwGhm
ewZVjAz0ZfQk6xTG/UzXBIp/uIxuwgpe/rsQR69n5I4HHVK1dUHJ3QGBRxV0Srj9a0fNgqX0DUZs
4Q8Cbct6G+m2KqGjRvavffA3AQhfYSS/amOreics6HDKMOuGG1fngq2l/M70DNBSlYWQDRR9mCXy
i3MAySlaPsin3RJNEhNbMKqOXetZ5BzjXY655Fqw+YNlr87138tHKvzoG7cHLLL/VF7Qa5Ic9YL+
2C4qWpDEmX0HziEOhi951NA64YFcTUmrd20pr8ggTfhnSfsY2qUF15vQ6NE1W9SE2zjE4bxdJpU3
Cfc7Fw2SSxwvVupA5i/npLlHItlWo3UbYzaE3198ijNIfYAtkcPh7L21yWk95c2TySsosRKU69N9
1gytZy0rDMdIZQVS9hxxn3iR3942ihmKvLQhuywpOf1G3kBlY6umCFgOkWXOxDaKjGZVnSTCxBST
oEbz+etPi2jVH9hWdCZDQR29jH9g/uSBsNiYbxn9BaM7ZS5FzOqi4TiUnIokZcjZlNCtHMRCA86o
gEXWe9LRInI60amQaAWXFrD/EfFAh1fXAlT0VEazAzJ3BRCr5meP5lMM8fV2EsML2G3JkOAZPQcK
7y69ix7/likZhZfeOSnsyQvatZlQpB9961GmXd1oMZe6r6d4vpAl4wW6BcDUQQ7OGC0QXZrCl/2a
2kSwuI4lCKbIymD/LKVV/Txhdum71LFQbmr4Yuc1WV3OzqDVeQg1GjWKeaYGdacaKk3vCa6FRGjZ
owRBfguTQmKbOScgx7Z3hRcgtWnioN3lU8+kx0EVVzCaN9+HcWbDdFmUPm7cQKVcPRU6gt3R8Gbn
Pjs2rnmisOW5Hqgt3A2u0Amj1y9Kj4X22EHGA5llzGjVj3YnCVHc40I5AYWamj24n8nIglxa24H1
De5p/525BdaeHj7rWBawW+8S/ohtZmt2+e3lrl6tlP1GYCMerlpbpfNoyLaEgx7FOxIKI86+DaQF
RRLD3C6DYg92EXluaXgLfUA0gC/cq7/6BFPWbJIeJRH0QL06te+gFYRmoQwhjokcOlK7pashawrt
y5t1SPKPWQsv23SgoX75N77XRMcPEZkX+BaqIcdxB0NXti3skhYBLqvoZtn1h8HEsEYkzelpzOj9
etOfKzSeAJ9GldCSnApZ/pSSNGUlSMj6ezWIX3hZGdHo+tkbDVCGy11R4ra+/rskYnQsdlbk5441
GSA6HiJE5ROeRUDd6YZrMNnOLx3Ax54MxToCNM4D+IDt3TQrihJ/91Zu4bTRfwSE45k0G25NKVq8
RprABY3kf5Ikp+WIS+tMIP61Z8BS77UKuiQ+kvMmO39LW+fd0UN75E1GbZXCZFgY2SdaXcPNms7B
jPB86Qufcnglqo8l4ZZtntL3B6bOJIYjvw+3l+kg7/sWoEuDt5tfh0rWMWPGC4GK+OZklg/bQOoF
xJA/kHRb9vxor4TAOOnXA2GLvkieaRAqrYMGYgQM0YkaKrhSmW7F0EF2WFPWHVFKVczeXiLQDKbu
OxFCjgy8p1DGkwIVCOPFK71Maz2aW2sxublqH0uKPmZVkqh1P36gNjq34Y95mkiNQY9F6ltyPBem
1hdSG1hSczKkibY/IhiuTsfGBoJZIeCEGiQa71y8p5HDu5Q+dwUoURnyjv41S0iKfYwqtO45PrBm
L+2lA+n4krqcu7Uys4Zodbj0N3LlmW6yy+k1Dx+akJxuXkEVnW/+Lqjtwo3ZBRSzdzWUSqsCDsjL
YFHOakfpRGPPH8/ryBR/b8YuGXl0ZlLyJGPhKM5TD9KZADhkoDAV3sDLsFvz7+H8fe9m8oLeYKTH
KtgokAq8+Ff2Jf8RJqr5MV54bwwbwtmuGYgvh6P8VE5OzwmB/Fz+jANBAbsZT3AJLi0TUOJthFxJ
PlAun3NPbNH+A+9j6bl+2xS/xibTea1G8lzrvIaxh0V60/bcE3ORVqdrqiqXNTUq8stiAZx1hkn2
VekGrgzo0kZO8IQF0K26MZVclIyX3wT+IKyghh1oK3DSOUiW4Rb7YfB8yX+OYr4omLya4YW3RIT9
Cs3XKnT9lThi4PaKsFXdi06wz2KNnclqCsHSJgTVxdLePDaPtfrSOc80ciOr2g4vA3hc/JF4ETVA
HhgxIGuo6+SWOJU8F6G1jHfANDyw5douUOs7+OBIvb55vzeTc/F6h75quPLPt9yZHI6zAmZNKjV8
dEpWQI61+if4oaReXcJ/aLgCX9MiEUCF1ikqsK1t3cXtdocKUZq/cHR5LmoWB5JENEfE6RRBe4Dh
odmijlHX9JbsOQTZ5hb7BvzubeiN4NShJcZJflj8DF+rAC8t+5xWvfGc6P7T5Vkwh3PCw954MKJZ
ZyA3kgyn6xUKyojcZBx83vvBPq8g9wXQA/emC9eqEY5YHxaczwLVqJ15oMtLltVOcQs/XQd8ZIWm
2m/WO+QIuxhwu35HZR7YjBStltG/u9AEFCX9d3CImsnE/ObfkuI+tr5k5TkXtV0J2MnBpqh6SXGp
BEY+QFYKvVrxXNsFubWWXVP37BjxfAD30nnG7SY6+HIuDLdOnKlQo4+7RmFyT4XMverOnnhYeIXp
FlvdACZedOanktpaBBc0921VF/jJxwZ/wOPUfvqqY8z38jps3r/rtauxOB6gfWkUQkrO2x8jyBf4
4sxbOhuWEoVOVatDDCgxFs0kysMLjh9mIRU/GpkF+XSWSSxQ4nLy64X5ePYVgBQ/NcI0uFtQ2tze
89ddk4hsB8dRFKe8P+FQUHKBbAjTAgdr/v49Gxcbo6az6xuhq2b192/a3ixWX3lsT1zOCcajenpY
qvLOXtG03iFcb0KyrNINUgoBGQ0GGFWWzm4wSF7iCe2Hcf5wI4Lsf8uFlzz5Ys+cuTpz4dt0h0ZW
ytyAzWKKf2H3J9MD6Nlic6GM62Fo+KuG3wy5jeXv6NVlNNeNz1QAWF0rCNKfEEn4Zcfzuyn8EIVv
+snyiMXrtw3XCkwMPcvSber219pht44f+EolC/Wiwb770lEAl7a2DEHEvmjqzf11q7oEwjZE4Ob8
1mCB4E3UdNpe251+Ggi2T4DSHlEVhKVkIuuwjoZpjxG3KcuDeomUbn55BfiwtoGl8IvND0uzBkUu
TZnDXAC+Lgkyeqoa7qXAM85CXMx3NIfCGU3g4t+8cfesXUmabNA/LKVhLnBjeEmjmrc1Ls9MagzJ
eTNGMjbg93stdnrJMC676r71NEDmFpT2zgs1V9rROhLjCQKjg7uNAdU6iR/F2iH5IRl5Olu/WquV
u4J+727CduCmLYM91I3C1beWiqJFTqzGKkiPBpoWNRcOFL3EpkvRTGuxnS8Z0fMus57MMIlxGxqc
XX+xBf2cBFlLTVh55N1UBPvRYvDHk6sEqr8JkGdpEWsEeWo6O1u1z8ORtYWd6F4TsajaMiqOcUvM
h6JfVqOMyReSkgfiyuLV2KstW7WntXUoyI4q1IggEOFf4gBWle3fesOPT5YRf0K+Edklg4NED8mc
6PNP9XYIg42/DEh6aj/L3XUDiKM1b38/XdhoT9efuBt+T2rU2k/eeZuer0nzIbXyBvdKFUSJm2/G
FPYv1JXOHcvHslJmJoKiskpRc4aUvClAEFgxM7Ac+wQwpDILzc0NoJm0hJAZDyS4gvxZjdMj+86Z
NU8kVJ6V/ef6b0940XwffMWMgPd2rO7jbOrAB4WlttGMI5dpMdC35B5n8qwgq3HD1lZsRLO9AfQB
CN019bXyTfGQhgUVDcyZ12QGNmSHi8ntyJm6hTwnwHxGM6fp3kOWvIvEGfwm2yluFce8GgOshgcH
wnpFC0+dMX8uRzkPfLeP1AhsgPGwjqXfAoy9FT4T9Fr/7v5APg09R5F0zKPcPNYmi55BB6weiMJg
rEDQj3gndnaedQiXw449d9dKXt/DzWP/WLNFtOvxeYcd1YkiRgVqSRzDqkctBeHKkqEsd540uUQ3
YdN8eYn3wc1Fi3dyF6igkGukAxYkzpbVrrcjgD/w5ok/v6B+KrI6rnfX7HKcIzlesxOPTvOJxwA3
JKkMQ0H6TYo1blWms5s8+kTHPUj6z1Heu2HboCht9n+E7H0x7bcwd7dnxsANnfnw58T1Kt37I91q
6XIdD7XphRuGA+OjAZeFo6ohSHg/zcKIIWL6ZESBKmi0bsDQzPraja7CApV69zPQ40XzY+F6ahR7
Tp4FhJp8kbsdHaUCBnwBBDe047p7R282leL3JyWWewfPY7q7z89kww3IzE+USGgVr1gcgWjos4xV
E2MKq5fxS2k6YQ48yMB8a/QFd5HKS+pQ8hrSdAwy54gvUD3jlwMRQznJKuM+Vq2zz6EgyPHxOuBC
71uyQx9kA6VhTin2r/ftVzRqlqMZ1tMPxCi1zKL2OnIh4nnEf48sRf5Bwi55ai89CU9Fce+zQjFg
7kd5irYX/dkAY4MInAxmoypjlWbNnLIaZ4QlVanGb26JU5AFw+Eh8Wy4dtzc3mxT35X0RlJdxYQh
SBNsNSfZ0mVWTyjxia59w9OsDLIa4oB/MJIhBUgIJqBL3+NVNu6BrE6+rPKUM4jFu0a6J5odDzIS
GwzOK0jUErCXdA7NCce05RCNhvaCLD9afxvXMSXpaTxeuO8zBY3gjHdl0HZKPQW8GvPPIn54ahTW
BOQEgpBlNu2IRaU3zpGUDS3NWPECXkIRTqEzajaLeiIliYFv1tVi2gUC0zEhuqFuAMk65CB10m+v
Phr40Ll8WySO2HGpjdPAfAEFNc/DFCIJJj6EFW7go3i+ewcVgISt4NDfm8wpWzMBOngyG79hOH2J
DMti4GW0qkpgKQTiEDP2+MYsIWcLmA+e8qEZB/L7So4d1Pj4DxxTPsgjP58deBI7kfOwBY5dvYQ5
DsBqrViwlTaGlpwl+7ijjwcoOiNWELbrCyDmMCtWPAXssqN8NnRBefZUkuMvcgHcrvvkVbssRN3W
CqyXG6dhWk8rcrPSYgr5CzgPFs/QFB7HgOw2r4bDX8xkLHYGXIkAlIl9DatnPR+yd4e/lQpG10Tb
nmq5dJ1c8S/z4RB+YLiY1K6fbmA/VtOHTG2UvP1hfZBHsc1VKPm7nugaphEy1TSrxVQG0bz/DToU
kIAT0NT3O+oNpqPatAMXw2QOE8HjK53neZ8GcBfnD9zLRDq3HIDPZLqEfLBr1s6TlnXbslHVh/Z1
6msSOS+y2Ns7Bijc7pxubVheGLhiOQqkwvJusjm6NeTzv7OuKsQpY/pACbi2kvhI+XLUPJpnNp5p
z3ViTl8ZXekw5U6pj2gTvSxAusPmOimbyhfuIYuP4di0asLCEcAHkjcIuEk34w1caD5PwPwLQ4Nm
xyAbxOi5/9773gkh3fdbb13Mr86p0pdBL09ivqYd0SHW29jrg212lsqYKA0ExOINZgTXqoN8R3p9
Ozf5lkLG18dHBJ2WiMHTAcVeK/9gEHSt5WNo+KNycxmUWEaOlKD9heBx+zAOu144DjlcDV6hhFUo
otUThLmvKTVcXf5VpIjO2BpbSCX2uu3X20/KdV2h8ya5/dU8pvRDR648+TgFnBx1nh5GvwjSD489
xgY1xJ3UrfkK/KVk15/BwbclO2rP/dq0asgKipfTzL9aLQYY3Yr8kNXOF9ZEu/BGcLCmzV6yLdcB
U8JUkdCbppuqUndM3WNUmYBpatT2gsiNq3PDkFRFJN8TTxCCSVoIH5s7uw6Nl76eksi/xIfXanKN
5P0/1kUsEWbE4GvwJWBrrHSbX1Wepz9A6GU6rGH+09LqGB0u7DW+CLLscMVn5mV7R4D2TkmkYOx9
uDiMd+gFKK8opJ1qRsb7wYV8AkD9nnu8H+DCpU2987OaYolE5fFjr2riLUMABBYmutMyJ0Pu0jba
ckyGYgSW6GwzMDCfEM7Hz+bRkkCd2iPZZ4vEnmWDrqJVnHiYjkQ4C/fbFtbCuTM7Yey78zZwWuHK
+qh6CLPgEpYIhO5o+y42C7oiPg1/iBV4EkGz/8AlQK6eQoEXw4IBgdlKLLuSh5s66ixyWeLQwWsj
lOHJNPZSqAqYcSIQc7bI8EouRexipf1CjSOPgz3oOe+xYrLy9nfq26zfB9+iy9QUdxq3OD3v4KcV
qBfGLh5I8uxUC14NdpUT8+7POXy3JuC9Gw6ZRyl0SFroxeyXKowGw4/WZTu128IU9C1htA+3xQKR
9qxNQ4Z3b/AEEIGuV7kLiThtPzYqbYOeSX22zAeJheeGULPJ/00bB5/kiZiNNzeiGL+fi3WIFuar
T5CuoW5oyIl+wNW4h6Gckt1YtgZV+eTC77iwSayiWboZ9hhTER25DRe8qmOlvQIs5lasy+tlyNko
NlK03hIHy7gMltY4BmAdvXlOhXTWTkBVnPfLvNqBc5GtJfsS4yX4Zv1predBdnLno1rfnP5aj/Lv
Ms3kC0h6bvrsTX2dyTHfHdq6iYT8axnSmUpT8FCMGJqSPS/p0SnkAOqCx587XUPf8L/t6UnWaE49
k7f8CLSwmJEgbWmxCJQb+CJUmNN9pwlZzo6vJfdZdehCQFCK8yiogIk3903QkIoUOIHwuHTqIuiv
88BX7+V4kjyvxacJXWft3kPsXJe68M9BrbGRQAnNPXshZGs2Xz6sP9fz5ka7VW9gKHaM3R465sEv
G4Bhe+ZELCC6OIcQPAYtd6n3V0H6wtNKhEb0avoUA8rTqQ/R5U8VyhHe0XqD0Gkwglvq6nqN0Ufm
+XugVuDseXpYAfBaVwzHxUPA9yZEpciq6GdcfqaMRCA+rX3XhJnz2slNXmtGMrgKEN6yh2YT3u93
JM74/H7ODZsBmbNvlO5Iwr2lp5156maEPtoO+qUowaQkfQ0sC2kv0YA3Y2aYROC3NTPyMQVudU3c
Dnt54x5jy4JctbLLsaZNfZ9KoQ90wOWqF0KqKeJKhXvDcDXjKwqE44gGrbe+1xFRcCwdEr1TKAxe
d8Z6+Zj8MX6sYdlbj5nDHfa7gTwGhmsSEKBsMqK+ea7Bbc3+UJUwNJ07Kfy7OtCrRB4qpto1mxph
iQtmUsMjFZTOcff2Xc0q2kPS6joWi9YItuV0cy4ywotAwjsG8SND2YJCPQ6Mqc4lAHjsw50LcVPA
t10hz2qXpFfUEuUqQY9ZGGwbNoPu2oOQUDTzSHlXaMQYOyk2MpoL5R9YVV7N3wzhQXH1kILngnyt
s+yuKTYJXOLJAeYFR/nj+hYgCRvhMDlnPgl1lmvo99gUWhITbyNNsqEEdky04zfHBEebDGnLMa8h
RmlaQr6BHoGc2vAzzv7di7MQOanW9SKnKUIu81N5ofvJZGwzQftI4vA0K52vBoTDAvv9M7Rmsuab
UDnsN/4BsOFNCKCpPvZZ4IS0+8m0tSUcluFGVNlswNFmPS2nVBnn+YhYMXNX7VUaOSH7cWpWhJLy
gedJ71XebvvLgmiyhE7DdSB6Fksw+TQDbpxqM4+CSYqq2LCgN90m96op2R0jeec3YF4qPlnRENrm
5IT1kUq1EZGWEHg6sh/qc/B9VGET9jKvHkdEaI/3zzmP/ZbCwkcpMZj/AulLzRxkSbER+Vo9nvsK
t46Bj/MmvPT8rOMQBadcRz4SEHvnmGwLOrcQfAdGBxFQGmoDGmFeaGtKoxxEcUuevABbETJ5h2sr
lJpnLPXSk+b/YO53v8NsSUKkBhehE6VRqoOgYqW+KX2ZXhhWZWt1f4eSf4aZwJcXGVcW+PJ5y0so
Mhe0IrM7ddFD88fJ9WnP4aJ2lvxQNv1Uq4rvSl2Vs0Ku1ezKy+HbpMBBB41ZStuFh+pelJmuo9lP
G+aU0HhEn1F8KDrDt3kUSQkL0lKWCSm57/VLAcCzhPkrMTP3mQNnRsnxx7Ou4clV2pSPie+k29Cz
X/sYR1NFoLCOhhFLUt8qFyvLcpQ68g6aFW9JsSa6jIZP1J+juGdDDZpyhBqNKBB/8YRS3/eBeu/B
xk44dlmXc3OvGsQn4x92wXYsAC3A2LeL+Y5BwIjEBOLotf/vxrWqnyZ1/yPfyIfgGFnv8p0UUT2c
11hevWbtyktVt4hPDibnijCUU99krOpmubhEhr+fCXqyAaZkQQPDSIjEwF5Uj+QlytzkOniQybdr
2AXoRA26Nb+q58yo8DwXJTxqebuH0IY2bQYWzG4b8TGgre1SankZs9k/BvOQo7CwhD45/oQ4HOvC
/9zExIctodUW6kZR6bntKz6dXu1TvpZxNHVsFWOggzMYBmxqJQKTVcBB389CcjgpjFlC9+KDKHTq
95AG++iIWphRSB/DpY3GPMV6E+VzmzYlVrO4PBOrnQyDhCgoKCZezsv61V6ThIkEfflB/XZ+aEqj
kFhD6MYGaw5jKwOErY5upERKK1Gqdp5BBGjswQr6IJ8XZSiJjVbe1/FTaELM8UZJke/qYS02iovC
RC4+347xQw+qfFV/YgryIJ79weEvYQD1Op3EHgNVe2gTpgUr2EFN9pCeMlddOUjPBOXXQV209BmT
1sqa30FlBQbWz94jA2Dz1WpDGbRCWCd/CDYGaGcA0WEZMkhlCQiNbcELaQqlscHnZAk9B9EJqOHA
QLJwga7JjEf7zkrx3+UA9Cr5E2/bw2cIcFyag5RhSxkUjP35Dru8LAB3gERRs//Ywd7oIDO39Li7
MuV7pHwjMmPhXy1Udhzksxf5aMKZ2wJHATTr+Id8QuX3wg7dYlUFgcN7qCspe50AOcxKgW81/LJD
sXjb7YMOsWUQCDhviKpDJJL0vdOJbOi/+Y0aVU1gR9wqGjghX2Dy04k8xGFtweym/4MM7GwqqyJf
GYxbo/CHS8gWQWnPknhSnwtj8TTKyb5uzXq7se3yO4C3AubHf35YZ7RjcYlpeg7jR/ih5kmpNCFF
9s82bNCt3FAWCeDlynL2HCZgl20KHxkVmMEM0ZIp3QrBe+O1jV4V0dh+Sx8R9DNWUm2T4n1ErYg/
HD2zssrfp3x5C0ArddvRf8MfBJ7x+7plQYzOKAAppyRL67+1oE4WTXdwZPoMaZjSL3jJcxgEhjEG
ToH+uShcYWo+hnx0DhSAn26UkUwf7llqKst5VKQQtVF8cirPwlYcg4GPyLIYP+PFvqBrfHsZn08j
8d2Zl4tl/DXDm1wd8u1vlD+9aVB2+LNhzf8xQAQl00MzsywH0sO+CDQqnS+SRTWLsP6pjcr0mlpg
k+Rx9P/IRxtE+hyA7phbiMnj513ZiyBKoyNt7+VrshFyx+HUGWb7E4ytyXRC/fqKy7lQinaS6SB1
QfWrccZmL8Ye4+TlkUV4bN/xYXXkmuyU29A1Ciec5M/F+k4/QZEHL8SFqOIgmI8oh/pVBJuaZG2N
3ZLi6aaSZfyMK5v0ScAApTtD81cLUWNywHxeQ8LtBWU2X8qlHd3L7hY9qZYscA1d/6kFqnuKjnUW
5iqyrgmJgeTndTqcL/jPF5ZuSdymwFORZYSOMNaIpKC4niygAwsb89+4k2P7ql/TOZ1Wup6zkhf3
x+GQGcG9qsdJYmPneYnsSMFXeO8SRrr9atbOmEFS/MhnWnHBGiRxZ+IvjU07dXdd4ZgNDXRdDqSy
lZwOAQzfh+VKaiMAKoCsejonTU8nzH2P+aCOSN6JBPYuM1Pz+o8LNDSZ8kzIulvLxf31AN92anyF
z/GkTf9PO+ZNA/S+sTUV2RDub7xncmMzwQOiyX/7KItKSi5lagP1nFrppjjDTGMTMmxPjDBpDiUc
VprfcsUygGJSASSF3i14RwcFlQMy+A1YVPvn+hb07VHnE7zruGUVI6bcYwmih/uRM4sw5mzExNAK
I1NOquFVLdNjsHV06ZVtqIJNV0CCVsfJsWW+5CnxTtlGeQqaS2HCNdtnlpfUVUpWms8SDn0YzGol
2jzbuKaMCekehlvCvynLgyQS3Zb6YjhQqLxSE6z7lT5udw1gidY28Y2M4jZTvTJ77dD+vTd3ml/O
lVVJeynzNfCSASgHZ6lmMK5h40l90HvJJCozRV0SzZ6gE5ZpZheBzMIDJXd6sFhaa2+eoYormelM
o0x0ky1bbQ3Ax5DtWyoh16Aaacfl50t33QlhyCG90paOsXe1SvtnjGgYnhzMTEFzEoeGN6bgm7nq
XYU8/kNd90goCS7UraAMa5dB74dyXO5Dg4Ndq0fLwyzVehL0wk9MWfko7Bu5avWB9UTyg8NJll/x
cHWbw09LsB9bz6g+cfxPJuVJlguEQrqt8k5DBXOv4QZMdJLJvUlcY0duvdpw/w/L/K/ugyByiuQ0
Y6b5J5kKbEBYvJC3hfKOIYbXC8iFSxFtpKE2dlOrUwmaZYKaCPB+4iW+3HCuwgVsprAM8zecvIcC
9slQxdPdiX6Qm59oQOQPte3nfcuWJAW6xbnkWmEUZpND/gvk7zjU+8m/2Wj9pLiF3lxGx/yRbNhJ
9dl0Fj+0mhvpXSChF2pA9yQLl1CKxnO00LcijA7wqi78s0cA2nWaaHurB0WBdWS6/NapaPBO4nfR
SRJ+NZoffWjNFsDH7SwLd5jq9JhXsbJzVYUkRakXp5mfiphEjhwQTCjCg231f2+o54Y1OfdMu5zk
apUfszX/oslZ7YEWSuiLexXGpsCrjB+tsBTvQ1dJ6lm3O0/OJL7wqO3g+bM0v9HlAErxW+NyMQ2K
4ZMUg5wh+9rADzi12XSxhHOeeAQ9IGZmXg0yWsxx1QqT6K0FlESofO1HHvRjxF8J3J5yIWUyBlXH
a1chH/iyWcV9nkWwDJfb0twzc4cR3LcWBK7loi4tK4+xOSu3ke6Hop9TRUr+wezT5H+j2N5Um+wk
nYdTpgyNWKXLsAhEbL5iKN/uz8HRGDwfnYSdlHqDJpbg5vX4U3qBdcePpjUJ32tniavqJkuCgue4
CruorlE7sgA3kZq3NTZqUhjJjiilVPywKW+cHxteF/Ribm6WZZJ68BJU5MobggKCfdY432ihSHLc
jXeuqMFYiUnk9jsZMUoBOCDohDrQnLSgw2nrRjvt7yomIkWUwKxqeltoIfixDCKbiL5NsjBHfIm6
4N6RonFyOfCFidfcqlL0mCxFCUwjJne9fbX5iwz9PmCo1wKZqBG/X8S7MhEnkhXSFDnoKR1skiwM
SiaExxJCA7G2c/iUwuh/MAk2yuOG9NvvnNALaKu6dYdqYuw2Ks7KQp2TecTJyjIN4R77n2435twJ
1gASLJemj6rtVl12+U5/Hh9DsdjMkg4JmSJ+whzX5Inr00ZA0oDY9GNENFa3gDFnoCAq2p1E6JKx
WsI1CjdfnWGpSKXp9yjcss7ACIYB6cG2AQdFKJDsJ3ipNUPXklUZRYVBkgL2+nFW+4T1IkmvPh9I
TZtp1VZdeRbogVocPvfiOWEkEcOvzexlaC3DZ6Zj4H9NIlyg0WPadf/94AqMHTzanIJ1Kd0jO/Ed
jmvxkcBHhnMzXCiMJQChVAGYuXLYU5HdVClRlj0g1WD6OsPTirO8ulTPo4zCVDIYSmJkqJhuYdJl
7zOL0jnbxv1292Ve5mXDtG0Wl5XCxO/FJHSc2KXV9AEuUjOH2/fxoI2Ev9dnGwP2EiYue7EdFx30
76uakH0fdtUFz1ZrSEHWh3lP16MiNi64G80K3VmvUdsD1SuWVxRI8ePku4jWpT1VK60CTdUQ61sZ
xRb7izDxTV1mV+5CY46DoxjN26ewXbTL6pmJibYqnbLAj67sNLZ5bNcr2uEZ5uiurfILO9WWDZRS
jLU15OVrJDzdhkCXLHpoaBKFKtwHzX1wJt5+eQhVb4gh/vUxG3FOvJsOrXQWkz5FDY9mjSICeHK5
1tb0Ndd6vlo+oX2XLu6JYd6g7JmnTlHwfqrAe75Ts7NZoqohgO3eH43WCn83PeVCv3giuwgR2yKS
Opql47RK0eAwNZ8uylhjlDJ+aOnZE37p2hSgn3KFNuxYJrP+fQn9Ebck4RKWvMqPjVZL037JTIPH
PImfmUoflYiX4eHuma0p3sJhk1KNCUAZdiQJSS10hyi+XeqdbQ3mYFQf8Q+EgWG7iKcTtLTsdNbe
Rsj4z8jWS7CJNThsfiQjNRggw6l/eKc9Tyvt5kEPuaO8kS6wddHMLGHKwj0NCWyORN1mAWPKskEh
6PzN/rM839LVsnhuhv0omP1HoUYtm0IV+UFh3mjb5HDcCEN2D9MMe3wKCRxg0S/+t6YT/+VrPE7x
zxz9DLfzN13P8PWcIRoG1U1riX5Xqf2drZaxqF1lY4KQYLVcvDd0rCVHEdeLpxUtY+YTauaRUcXA
UnEMQ+FEEZpBjwKV5hcgl3nnz8suvMOWIcSzKJfGxNfqYpwr6lelLBXAMVPH6gQwpN+fe2inzosX
cZvULT9yIZdQDRBWQZp4ag8dhags2mk/vBJDO1WcRRuPM8lgwI3Hly9L6zkLs7SqP3ocFoKk94Ka
tSzvWLdKe2AsB8DzanirTXQunPx9TYBh/Gh2pWe/0ZcnxeUvop6AR8f5zhF1tAqaU89pp50jXA9w
o6kEhhu7oliIle40zYVFiWc+PE40rZXcokwRudbZ1lqaNDZgy/pEO8XvpVl15jVOFYf/oj7RYlip
C/RmhtPbTGtYt/0WGXtaX+Ex34yvSNVNZ3HPiMeTTOSd5ho6WILGDObHgXqi01iiYfVoWRWBnIQa
dMNyAlISPJnHv2zlqemnRbMi94ZsbhYBaTqSvp54WVgduLausIKUrj3irn3b1j4YnDSCPT5RINBX
gu9Hl8g4yHhjLysd9MFX5Z8XMjwA/DcnK5l4ZZRpmvg6bWaceUUwRO66rne99EGtu2LYnKSlRZHn
+ecBYVHh/3tOXUngTDa3Q5u9EweMkG3y0nyziGDonXzqNQZEabp4JE/BYF3PsU8RGE4HJhnaZ2Gy
RTmcGW8qmE4Fwn4n0+EWg5jQGq7IsbOLd1M3s/b5TXw5PY9FzPU63TqPfez6SdX5mwcWZmo8Hlot
VWVdDzzQeIo2/FsL/wf/M8ApVf+1TW/b6Tdrdna4NtINgtcSz5BwGGxvNqKM27GslspCMOOoDnmi
6FPtoWgvyiOfev8FYGAGPqa+sMFUlW/QAgLs4jWqE5HdZyIO/bNd79/cA8k0/pxBGhwLSWnBXLyP
SO/kmVtcVCQyoT7kCe7ZP8yMBLGGErrIdSkYG+EEmp8RfcIdzwK/Vf07gJO4KIVm1o0xiMX1SgV+
nTl6ZsBzCVmSQ0UfWvIHNmbVF6eFkrNHhp2R0IGdevTrzQyKT7QddU5iRZSV0QaJKqE/gJI0WsQz
ko6XMGeaCxy+wqX6hzh5B2x/a2Z+zgTl/E2Kf5GZa8hUpDfsfGhw8zy8er3Xe2tfz3ca9K89Y26N
AbklhtBIbRKGNNV83BoJmorUVLIrczKpwk+XKPYgM3r6F4dnPSs890vKn4uFk9o0+T2/DCACL8YG
Z7358pa6XbkoJ4dwg+HQRKKOuGVQydPjBiY/l7sRK8n+7VI4YrurE/B8Mr8jemyW+RzRen700z70
UOkZHYE7k7jmiPX5tQ2uihAHdC54jjmcJCLxA7xV7tmQV3dzz8z5jwLbv2p+Q3/FZMa8UMgO+nKd
ihTSbj1TGTgaoixEDSNEQC2HDFmUfKxwLisKz5ElcQ1beH67caw7zmb+uqPUyQoZs6U5YPuAvqn2
ETggkfmkLV9DgTaV2LVkZq99IsqZ58STM+JaLxFEy6q4Ozqf8+zS/wzz4LM0bGkKTqfV1DJAwn2J
U9XYXRAXo6vPJZDzE6ItoaQ1o7ONP91zgt7pswjCeKKM3nBbKvlMMoRgi/gEvEOFnh3RnWmKLY5g
JjqY0JLNZNC1t/pmOMsAsAJAtqwMwQ7dAdLDnLcIBiw29Ay9IW/q8CkOWEI4B6KHDuuPJvV5Jjr3
Ne+6r+f8wC1cdn+PiIV4MxQ2rJcYwAo797cJ1vVotm2qi4VAe7jh80QaIc7/UH5lFF5TlBKganLx
W4oz4jD1EaAflXVC8a84CbYbYyJOEtdY4f+cD+SI6bns1HJ+bASDz/1hFsrehV8f07twcyMpDJBY
/rg5sAFD5ca4/e+oKJzBZ2mio3iBqbeSeZYwUD0H/jhhE8YKlVquF41SXg94/zsPo8EEC/8v/zVT
5vXGlCHN4naCwfxVuPezPtGdxmri0DxRzNQCccO6aNFZWd8Tc4DvPcRR8Tgns9tctXaP1TAcXXoL
GByP3xvkiuW9DyDJTvaA1bG1XbuRWfDJu68L4et4ebtc7iUY2KnFFu9iLRETAXC+lVWirzrQaOTg
OePf1awBVcZ8vNVpKt0jvL4Yi/U+jT0DaTZszgkACeBJQwAVJwA1E5/Bw0m/OE4pBcqU0da3dO0U
+NnEee1ngLOqR5g7DAA7DyH5Diuwm8Hkq8qlrucUtc5WvGEdBP6Tw6LxutAIAYxU1lI9KOYy+oJt
r44f5eVk8h6kB4ORNDCNPod391GwccCGT9pogcz2ttYLE07SRWww64tlNIj0yEdJjgz7C43tdz5h
ubj2NytPYy0HIpaNXeXh4oRr3SRFSbTmc9VDAr+aDOqI/qYzOhG11lrHK3+HKjnlq3kopznwhM3Q
+r7/ZSPO40hftkIZYqq8Sa76nQbZW51NdOKCGtAUfSrg7WMrsUnMp6cV32ptkZh1Dj8LqbVAMqZ3
ZNcz2AvnItP1ENIokrlPJsaLE4fHB/4+Rbc5EjUATtXyVqbeb/QO0gpr6mQu0XdulkJ7keV7PzYS
wcQ9TJVwtvp/fgXCDYWXydiaK4tG8QqlaVYaBh+BwpX4Db2Q/IHjTendjvnsTwHuiA47rjhaPueE
rDVChlwluC74njcMKY7y4BZUfbzbHThY0qFH9oIYkE5gI48KgZM04rTOAiLf17Akc8KYYrszXOhA
Bl2PiC1AQbF0RdQ0nyNZKq2fN4I4cbUYH3vDl1OeZRNWY0eqefAB2SjQHR+fLrxEvQYVmzPQqz6v
ieqzd3uRXyr4cv3MygqYdmkS69ybb/aWsaeQaZq20rh97pWP4MX+n5R60M7WCzCCqdihqJVJwbvC
Ntxas4jG1pn8pdPuny3tJ/6uU0Ok0w0PL1Do+pp6Jx9jQ+L7SiQq57xVTYgr5VGByiMbLHXVM7F3
oY0zIeh5Irl6RGH3KMdQnHIKBaKohhasjXLe9Zoxl5clDHrbEzV3mmJh2mXV6qEXy1UcY1FTOqDM
t7iD/4effowsiMeMxoXElkYd6Y//tOLn1tW6Pg7S/LPdWMgOcRytlrnXrmX+g8DDMdh+ISAZadSw
jrXVH6okm42IpQUju4WWRbf29gn7DIcrAt7BMRbOqZeZw47ZREZ40kmSP/qhUZzpF74yEPSmKD81
YuT8f72z05X+E6DIRIQQ9ioe6tFzYL5vN8EoGX+oHYkee8YL32Fu/DFMnWYn8cY/V7tdKAM4YAiJ
gCr8nxviO6Mb5/XlXxvqxGbKmompElXObhNS/T1XFlSw7hNE+MgrqvNF+dqFXnXetUBaB8fYrwxx
rq4IBaKJxudTN4PxYTTchTmpTs2jl+dNCfKV2H/gwYG81YgSzVAwCqi0vK0QX/2YsYlMt3CuSM84
+oDupNremRMKRctR0Z+0/14n0AdIc8Z1f42AgmSdldsKukQhmbF5YvCWZ11zMJ/Wf2fTt+f+Gx+M
5Hn+lLyRJgMESlKUoa434GmdWxgdq7IBcXEASdf0NY0vkrGvqlRoZWEdvDxnOSh/2ZfwRH2MUnCE
hWvs4U9Q6/56VOGvwSFqFIUFciMbdWG8JqJil6Y4f79NzUD1WwpE6hCF36NIWJefg9VIz69dF4in
h43rx7y+7dlnpnIcNRaSsL032Sw5IX5Mf1ixlgzLDetZQLmYPhOQ1CfiA6BIFuX5edfpNVebzTEk
IHVvi3Wrwx/GDntwJGy1ZTDGTMqG271BJNFHq23JbUTZt592Jf2OVbyhycz58KRa3n6rkV1d0F8C
zk9YV/ueXEobV0Dy94PplIFlIJV+Wu03GiLUGpZAYtlgHnsUrUdqzuxy1R75ZlVKeusjVJC1u2wv
Jmi7pAT8u8z2F6kLZ6G5YEdxwkpxdbuI/cHdFCoYfPJeA4DlVxLv01O7juwGjBu+ewYtrds+ufeT
zwoafPWJZAGGkPw8aGZkMQVSItqfBHnKn7v5sqIr5oOL2pbqmD8e4RPSAxI52JPpUM3ZKSUgJ85l
PmbIo00t+6HI2wqBraj4sad9SyNhQ5gT65roVqBmDYEVjhVggAJ6grjK9RotfxSb5wz/+HH8Q4UI
0xpUDqqFakNZesByNHXLE8b+l1FwvA14dux3A8PSOOWJzI0IhBEFZTkb6nYDtdb5Az4rdVXI3vNb
T25TyJt4HLCOTtegMmNTXjMDoCCqsiyKzwPJPkibBDpoRjajNgKgZP2c9TBfndGJ2kh6LcR1vAie
a7kCu2UPW7C/MDA/9NX/msJIy/twZCD2rqwBLhYbG4aD80mJ+36IDMTwZBfpeSvRbZuYrVHcpZpk
wQU6T+o+HrdpiWw23+/dkw4oEqUD103srUeAtk1G+ZUFX9VsdQkzr13feA1sGYb6FsSHlPeCcFBT
fCj+f39kau24taqM22e+qZjLgdWm70z6Nh5bUln3O57ydkSiQObtuHoR9JHmZvWbVsGsohVHtElc
FNOaFy4N2zDTsm67qJ3kgNE/CV+PrO6F/eWb67M7jtYv9g6z+H9yWFdaUK/fiXCeqOx8HWpDH2Nb
Kp0taxVx/QPp6R5368z2D4P7kivtE1+QHm/Z7Qg/j8VkJNMNxW6igwKzQ0E042dkaj0H3T0yLiv+
awxIjbwv85sRRD/xgasAqV7Q+MofXhe7L5IPR38RpIZ0odblN85DwIWEmnRwxrn5tIYG/I86c67C
Yuy2V15WYMGgvuMSVMEMA2Pwux+T1vkZQAJMLXcd3MTXAY4tnvFkr18zfe3eYCOtMRf2m03IZcSa
K9zrdU1EnUqECmouglOLoHka2Ny2aPiIj4uGRO41ffo9Zk5T45v56Q/RDJ6n9CQr4Xls3rvAHnpW
VeXi1wPk0QXBIiW3bZAo+hv85OmjRFz/Q0FPLJx9h0VoX2olFlU8oUIaHIZkzulUacmEDnyTVzPl
eb04rNnsF61oXDLT2Bz7YlfSvYMxU43yPYxB+Uu1H8ZVlkzXdXm5BbkRZJxcFgQ1Zhl5n2ZqAoXe
z5TpzY4YAPUkvvg44DehlfSfsft+VafFHnnpavjqB8kKoZbDCj8jtuwnTXxLJpXzfkq0s0s+ntZ7
SaVlHnM/oMaZ7SCb/UmUYCoaaqmiKg9teh753k8etz3k+rE59r3KVfgSsMMcYbxI3c8pb7JELI9I
Ib6ki0fyaMAV4LyFe6u4+gxoLPnGpfBNCpt9JpXP7F75T2nXmf/Z1HpFeWU+kOMKaitkhP49mSPC
zhj7VpDPLZZday2I15zaOM6DkNzeVeDp9KN7TUlpszEP6yJeYLhPuCDqP4Hsp0nYz6oSifW59FTb
Ed4ei6iH2DRVU1zbotmV5fjVyiPQL0ngd/Qxmkw5oO1BBYNfbX8CkuuKhKMstZU137QvnJukFGWE
1UFvig82GAsAdaDZSBLPdUMyMq6xSPqslhEZami138aY6LcSQElj4MctVUxB4+FGNaiitWYwIDzb
UfVgKL93pL/66gWFTuK69VbQYUyPpS9g2IcASdboIb1als8zpsotUbar0npeOXfJCq3ni4ZHkml0
NzIP1Eny82xuBJbwQiV2PnGU6+/Ft0Bnww5FJCgpUk+2uHM+HPQpqbgElgBcADwRiGV78xuWL+3V
lscRA9oyJO3gXrStg4fkoq+g2zSrf1Dzjn+L/9ULKx5u7zpEJ/dCCt0pmzvyvW3N1sTYXWZuxBNr
NoXL3IVxbze9AeFJOlJLxRCSHYMyk/lKqe3q1ssWs9KK5Nn9tc/+gI03EfQ/DnIm2FIrz5LMryxJ
kLoppE36ykjD12m3dGTLDIHL6J5VAiAJwUa7PdJYQnlsM2XEe4z8TLBUaj3+sjMGH+IuPesox5FT
m2gJsCi9QlLHjh/YGUX9ce1ckVUQjXw+o9hb2p+bwpc8E/RTEbzx/Heq9IfkUi7aGE2g3cREojzK
AIyRc/wrp9GzlMNTvsq0Oisowu7D+cCHQPqyecnvLl6S4VWBIMJ6VZ8RxU+k0Yt3hcy597X2BclA
Px4Ru6hjNohlJ/05hWwz8BwvC/n548nkcHsKREYHUsYS8NAVCXzBjlsOakiQyPh3rL2nxtVm9Zdr
Eag2ILVYQAamDU94ZU5iH71dY5mZJDu6iiTHRIq0nneuU0B6V7IZ2EX7FCliqkFqZldcFd0C6ffC
L057+YAcq+U0lxZ5Gezsr3+20EIVSvwxPDwJdLMEtZKoUwNjuHpOruglOuWt8fp2oECgPiB+fi9q
rUaOas/QKwuDCQuNs8y9zpCYrqNEp4kdHUmFYpJ+mwq70aqFkWXP6QEfo8weWqeENjKDLmnj5bXk
mVgoga221xQPQMZRYi/jtHmWxIdfPaI7U0u/rLSoPEuFeUDnSJVzNrgZpywDAfLXsbhhmqnVXb3P
s9p8TMMdsYqlYN/Zb2x+Ys32r7zVAX6jcXEndWeXANWnaBYbDgja8QNvSFWygzwjqzJCGkTw1kHf
Fev7/tq3inz778EHzcLFm1xijp3XaTn1Sh1OdoJYHa/OMZJB9uV0wI8JdYLACbJnAWYaHxVrccSs
wDOpMxMYSVYTjxdpnkLbaCzb2rp6SLYqlTEUa0gvvRO4Mlbc9Qh8AYkM413iIF2+6CozfsxZz0m3
miXtM6N6iIv+v3c72Bxz0upt7xLjrkOYGUGwRoizWIlw9f94en1R9KHytPPsGolmxwXeQnDpYUaT
C+3rSZS/+SesiRDMjmd2BhHulT+jLWtJHDKMoozAXPB4lKqOosZSEciMLEG6mjJfRMLV+/zqUL3W
UB6fADejEqDyncXjDTnouHsMpcSDmUsNSftlYTjiQ1qOpLa64XOPfkGasg8XMW3yT30YlpHCnJEW
t9KwqpBPGShR8zppd0kDZaWhcnPf0HClEhoV9i99S+9JZj9VzU7CNmILJm/MNooNp0a/aC7SgysL
Ed4pVm5a/kVapK808fCZWhNqOdZLYBazD29ccFzyjGbR4QQ/BQHNBJDatFhyMSrwS5Hl3W/G9tjZ
UgXAK4cfbKCtcbTMWhOjvZTG8U3yGEvFLvz8zBqHWiI5O6Tg6ru51WkzOx8c0txA3LZIgRkBQOYR
oTw5juEApbm7w7V9jbSzqVbG3wo9udQOjgXD4KbQ9a04R2qQ9hizkfGvoSjtHtcDWaYp5eXB15wm
rJuW5nG8NCRN3yBf4ZrMSJ84W0hq0iFl6T3xK2nV6dzUyPKZNUDmkZ7XCvqrMGr7TAfN4Xz2t7oR
XZkqXT7xwtSuGh6eBhnqrtRej/mpTKhtHXqqYhA/3Ynv8Q6TM8CK2xWVElfPMaCHblagmeSFaTlG
HmVfs52I5SGC9Q+7sb8t9xsZxglL1h1Y8SzBmqJ+BZEth9fGbQrdzI2lJRfnbwnGoiJDQgcwen8k
zl1WVwlMVpCs7IwbMaOEHMxEfTlRLYLmYmr0rjK8wx8ldnNg7UTxdP9M/9omYl2FRuQa4XJlLEqs
EKQAPc1uAtXY0K1toV6bHJAWoli2Is7gxgHfxYnwGGnv/rC7GG3BVY6p4liUspSy0lqg+E5NC5Zh
9EU9RIWbqYopQ99aPEoJvxH28LNycWlCPXHUOgBLLSxvdwtu6SqIEtt4C4n19N+T1uoLHDJBDZD4
KEtSXAYuYPDUKiQwaRbgzLp3zLLmfj2DM32z6ufhpqDT44dKeXYhKru5hscDGPr9bRTfpno4Htn4
7n66dCjuovM7oqsalLuwfVhqn+59TrEqlZiC42vIdFvNZn5Gy5Up6WMuORSXHDzfEBKQEyXKftJy
ZvWNuOnLGg64ehMJm1JWj5B0A/LDp2gUNRzbhRD6y5n4rEOFyCM5GOxw8uGGqGa+SO5T90AJz5aU
Ou9xPKDfc8hDeIobgO+EZApQgxSBZ3iO+ow/MqMnn4w/rkVC7BEs9VWDs0b2ju5jWHKweBd1HpCH
rbXhrbS+RU8qAACKKh6V6NkVT97IHC9z2teXfI20UuSJ2rCZXJsjmT8ig9kCz0rwgjX2LayInu8I
61beKtORlRhqRPMwDZyX7Ok5LeC++YPjNwtQleia9DGw2E7plGZruIv2ziILY70nYIVXFYLAUeRI
wS9PHLEH2cHHdNjYgUM4DFpmfso3dcqVrZz33esm+fRP7AQtZNHZ/nO602SNCpdmXdT+aBIJMVfg
ZE2xlpf3pn328ZAEHmGXZNGdeMjwDafdDw2EDj9l2IF9MciDNINwk3QEtJfiL+IwgtC8NRPDzOoA
1Cjel6Lp0nu1K+mQQXcWc5vmpARJt1hH7nzeVuxQ48cQ04I9voOsWE+HvrPT1VXraQgT73XTUASl
Yl45T4tJdio5n4dp+dNRIZAwnmlEvcNM22ih/h42d9acrHgOka2yWpAsDD/05KPj0MLJr6bQMcEG
I7jTmpgoZ/pbYhEhk0Qvi3C2ajr0BU2lAI2TQuUbJpMTYgss+sTGc2jkQwSWJNxZpZ6XkC4jKhYq
gEoQhR06MP1hIr43Ix9EHrlRZDrelnkx8UxY5uU54E8Hj9nc+ulFFbRkSijmB7PSUFok/oDmdNSx
CPmYGkGqhuw5HKTa1Ah2Ug2Sg085+os+TVL/Qm3mdyRd4KL6axBKshLns/qOxYe/Q829HYdfHQGG
v7SagXam9yDjnFYw3ZJlNnDdy/Zvu7Rt9cJ6uJZ6JY+It/1q1VXZkGl12akOqrrnaLXXdhl2M71K
CF5+SY7+90FXbVCIgEVDK8cqE4vxnJQW82k/gOAViAwOjrHbDyrK6ZdE/yrfnH/tENQzd0Yj9JS5
RwyJL36KzqKybJOlDSh1EhYSJq8D8uypUw+niw9mp+UBwsFE78DWoaidZNjjoGmoRxGbGWegYF/9
cRqCvvOVuWIQR0jAETIUfJxIXr1Ko12kUOxW/HkNVyVrn95JQvQM3T7r+Vf8W8w0OWX1hDd28nmw
c1sMonrQ+A5h6dPshF0/EdLheY86s52qO/SMMzTvzXLqBvVwXk/p1ATy6Mdc0N2a0hGba1qhZeRg
VXndLAZe5L8YXoYeycnxvfK7yO8gngvyiZz44SPDIlpnRU0DLaYGgbvjBSZ+l4SQ9HiQltFypR2J
ovpp85xdZnr9hPNNJjfE/j0ouIklRD+01UAn4WdLnk/awibNr08lwdOHXCNtfYBVrcS3XhDB2e18
h1mnEgpupb1NqzUCchO5krYV3GNwjXCvjE9IO/A3f/g/PQdvqh1hdf4qESb+p48YSOk9Fez0UyPz
pMcLMJJMk8jRsvLAzY6CIqlmUfdDte30PVBMIEU6gmdeOQU+IOzAj4YegcbJYgg3mOhoQf8Biuei
oBqtZxSoyyfqoVpwVpphUDSA/XKyWefmLXqhjp+CFQucNkeg1uJyswT3XmLzA6wvO5yY/d/PW1Re
zx/0BFoivi+zM75WpY8PzEdGa6lX/BttZ3RrJqKcCAzm1A95AJ8uyvj40HTOt3Pu8Yk03yYAGL5j
ZUCYfw7wwwuyLufU2E6UQB10GZ4paIj/w+x/IOcJb7o25onmxsh5ZiiTs2gLm4uJuKgDPC3Vv85Y
VbIJCfnX5ybaBmrcQOzQv1qJg+h9v4+ZJC6dKNsD7PqhvU4C92sYNQq03soEtuy6asRqt2hsjTGm
RTEZad3Exsw7gpq1z5/cJZYyPgYrgezn2wxjbM+yXTQKtBwi3LIlTA+gUYZGq/7RE4m8oW1uXL+H
r9BMqbAIVIK0THr0zxyKIAuaVlTVMwe28nzwSuFb4XzrtCrFIws9EF5+vC4h/m31yLvwLaQ4RJN2
RupRZ3MzPFHV6xIzkSoDngQl/NFLPLJHJpveW3Ehuva02McVOkkxrCmjJkAO5m7MnlSNTgNO4g7k
Ai1bRKqMtLCQhHHEjUrM1Fihp+8nqzeyhiFHTvpDcVsi9JXtuXGtb/0c2IyMOxT1lspaim2zMtNR
FBuX5AK+tg5VrWNNTr9rQnuHPpHTgdPGf8WlaQCa/4MirACZPhlcxUmOpC83J2rRpW5OO9w6EfgB
wGf2lR9nLVGEY/h3Bf3oXwkoFcOIZm1FRicSnkxvYua2cLKvSP1JF+4vwR9xaKMKxuWBX8prIFhW
/esqWr/5d0eLjE1gheuHHCm2Pd0tYAajOhLqjN2cM2DbiWkGPzQP1fIdcJL4JPlfgQdjPbYEuzLE
0kOP1Qd/UIziFkeINUBthFXfzdj7NFiIpnIbF764OHC5Z0MDeZZe66tQXcAt4vn5P9brjK3A0y/t
reHbyIHVqp1fnamUSEjQR0K/Zuw69fkj7DEqTgdJInq8VOJErU/2R06awRcQ0iGRQU9X00llFLqF
mWvJ61sRv6SQ8+fft+gXzyI4TPhLUxOFzAQHyYSM5nVFB+kK9H6rQtSGh98MdNbgBRArwatGTnHj
6XuFg8H9iD0KyES94TxJwhu/gsDodXsjcbNvgbkJ1MB9YCdtgA3Tc2iAWwuNNx08M1tqMHoO945L
aR9zjNTRb4Nd1rcLVVDFtKXif+2HzRDkZZ2Y3oF59x0IO+dhkyDiglNI1kfCDumlO/ZXOwIbKOwE
I9Kw2JM18YsXD/qewaWUC6aLMtweCFK7v1hL9E0v+FW8QjX/t4Re3VLzmvYGBBy+MlgSDLo93Gj7
UNqs/wotSGaFiHGT9VlgZZXI9SbuVILowkIX3xhEK42g6RP9H7nqkKQquW/NM3jXwCv5mojToz9w
n0zgo+cab6lW2opDzamDti6QZRaT1fUAZ8KsNEix9HpP0xqge31A5VBXQUKTJhO1WfnQDMVUn4Sj
0clbNSATzimUhYOVHPHneDEZx6emtSYrjVo9aq3D+NHFIzTRXZWnekW8UrJuZ0wFWz4mYlFSUHgu
yTK3YmXzrUXpjFoQR1AA5ufU1wyCweeHiHTyte9KxdCYgpyxhQh2KqJ1RwNyqrYbQZ3AxMEbQKoP
aMRkyH4aPtK7jCQ2wArfeycI/FkUwP90+Z9yOlN2OAe4lIq/TDl2NmubianNui9WygKIvhZk/4xQ
c0Oq57f4++YINmKhnX1RX3LboCagH3vkv4YWv7oh3644n/YC2wnk6lMXCUMiNdTKU1L6lMr0bDqx
fv2atZb7G9gWOD0GDg4WLyAgULRDljLacu4T0O8j8Zj06G9VnAwCAUe27D2V5Wbtyz2kV7LDhErh
pmxajD6ndi91+Bp9pePbaytcyfMqXjtwjK26Zkm1v0/vJ7hp8de4O4tcfu2XQ8XK1kio8YKnx7ZV
bplr581gYQuddVzxAWiObYY02VuyKRc3u6ssKjQPBk1ojFrUVP+DTknzJS8+M8778uU5uOJxP9Ew
9192ck+KfxffudVE0HEP0aLk9J5d075276CwWkYUCwylWjeoSHuaptobhQCZb1zZ4G9PhPxN043n
7xlShBg8oyiFq+gCH3SYo9QbPyvz3+8lIU4EN9wD0lc67Nh9YILMBBTXbvrQFyA3dCXFRXuNIMmx
Hd1QfPqWLSw9MAuosHtL/aJdtISWDzguvKimLn6tWidKKAs147udY/dYwt5y4Oi0zsgm1gqE0hnh
4UNC6t9MCZ8N54r55E9aFrL2h7gYpjULzmL9XeA4osA7avMRkbY7f8Uw3FzoRYHSQZBugx3Wn37S
PNaMRqshKLQG8NWYnfbPnJ4s8uSxNN5I6F/ruP6FmhE41TrQ7si5zliVg2e7Lg+TH6Y5MH6+AP7l
dPAdGb4xxmkbUvK6PEfcrtAiPWLlzGgongfeLcyRmLuPoaEJllmdTHrxRNdJ5IFNRGF3Kb4kjDHe
5CP+FyAo1MDpqIZcynWwRUCZHDdWOa3Wwqcml0U3kfzjWw0jXxUf7enkYF8HpRKGd+GUj28Qjp+K
OT71W5+82Y70IRPg71rwZxiigPrkjKgpeyvpgeaVG23KHJMGZiBmUBLrF9aDTvaTzz1iX7NgCu+v
myyJyg78MIhQvgdO5/spu+vKQXvTiJREy1pnY+QRcKDwsaJ5wG6e+TO9ssTAVIm7YWqticrhX3Ey
jRsjiBXbOy61XeWD7yFnGhaWS3Z5EJwsrWP9bV4nwj8G2HRsPv8ux/ast5IVGThHwb4GVL6r6+90
eyokkJRHAh/o8ZtNp28KS3+t4qjYRwZF/+mTA5yxBRr7tu31QyI27tLzZsNtHH3PKzVHcUBUfK25
RD86gnTJZVErLaJozLtYFZ4DSp6to8yeLrA6hqnJHxL0NJzifqyRjH1nzUR7/OEL0zSzd1JFrXq5
MOUVlahWh+NeyOEyy5I87K2cnWe9+WRHJX93Qonn+ifJ1A/Ijni/6MxB3zB/nR4ezc5Y9OQdSvZ/
ybsStHFalDKGS5yDXBDvB8ny9Cz5dscyVfx3flS8JbCid5bI06aBKxYknoupOhAiQyn73W7S4avR
vwpQ3Z4w+uBRzNhUt/UM+QUH4bYOt+NwYl0TS+ity3UIhYB6hemxNixXlhTDLFL8ECchNdxzcdTl
rayBh+Tyitpp2lPynZcxECTNvOQD5G2F/PdoBiR01XuZKPWK6IUIBBKgHj2WyGoR+w/c785ipJ+G
bSjZE+X/2rmKPAxV/xkgn9yu7GXn7ydC7i/wkpRsrSCG7mV7y/inmPjGPz/0EsofNqzXjbLJm4Vq
7hQzMTOlORM1fAinoXlIFYckN50RM7ilB3HEgpefQLhMWTjWp4E27Q+z7j6hTWq4hZHjNsJSEuiz
MZydpaMeCeth107PX+IM6WMn39KfqhHAuTQbsPQnZRDIRlkpIdjnL/HjpOdFPbz2onUSfhKYrllD
pgpfjXdTrBtsrYNd9nCzs4PMIFkdTYjKgwKAq/A489KuvcoCOVK5/TPxCgXj9syQYGYuOqfw5rN7
JUCBAi7QeF+TxgrEbbGTv5scMdOzEfceyNmA2fhlbrkQ16mhZcwGEkBMG9inM1mtFtW6vbQ/MdFD
BfNwR8oa7723p/Ptjq+OTeT4QzsYGBGtyFdRz60iCbML32c/vuP/Sx8dUObbLWUYdruKYeQgCM6L
MfobxWdU4bt/nOfXbYnV7GP4OCmrpAFIZ9Xk968pSr2L7uIPUDfHUP+wwTDobiP0WHWPvwQhkoak
JPuJm9m+TG2l2MgTfrWKTMEb/rZ4a5o1y7a2pooQPMDFOkCcCkc5gIN2l+il2YzCoEVFRUU8CgGf
/ysVD5OMgnxXq/D9m9stOcYTkoB14yyiT4CvY4SW3qMKVe9Cm+d7hR5bmajZnFiMrzWQHTvOeagE
wruH9UyQJzbhJ9P7doM9lBWWfA+19sRI4m7nxF74quf6KxI9h0REVDvI+rh7LvwyWblBPFf9RyYY
4SwjsAc2prWSgkVaZml9HVfeys6UismriaIvXGY2EoYfSQHC1Siv5YArPd9Xn0ulbBLzItZNi2I2
5NKmbMlalA7Ga/qKT60YGj2QQfQ/ySfh4TOMVQrDO1ZUXAqXZBHgYKt0WT5q/1gR9bvr+HklsWF0
67KipqGMk/y9cZ2+AUPeudWYyHj5THL+8CwMv0E3vNsw0XY62jRPDGRJ/Bmg9iW5g8LbphvFQlIa
NU6l7GHN8Kvwk9Ja9DcrmiCUlobhHYuwt7cugmN3oDWo52SVUrRVkFgfg5c/LWXJwdtUKYLml73b
W4AE+2bGMWY5z7CYUOjTiGH4zIVoVGimz3oSdDB/eA2P3etXCoEsZmGQWUXg/NKEnie0DPOcaasN
473aVa4LxYu5j4+0pGq3aHeDCgN4jv4XFLYPd54WUyvna5wrXcqa4sDZrjoTiZF2I5WFv/X6ZdCF
2N/mEDxCI4wTP9KAiMxXBU1i0Z70zxMPuxoh0MRjdJkx+yTMG67vMSpo1nzKZVD+QFGC+01i+GaH
g8ikseJCboqOx3nuccTIqrcsjm76pAC5BPoWtCbPweKB2D3Ub/TU4r+GBza8NKKSY1TGsPTZMFjK
ahjv3PxP4HtIG9mSsls/sSkpDQDTQMwfd0eSWt+psFhcitwqSZY+WuFWhOuvPAvoH6MIBKJXZSGy
SQtg2tEeOcwdZNVPbfVH+vnB5mlQPPUsESD6zmrIItMy4B6s78Uz1kiPmnKU7SRDFgaFa3+CYq8I
SxuDWWVQFDZHzg4ulOWBNOssYpd5nGym5eUxyV3scalDGBOaDKg58vVbsrwrI7rj5n6KbGjmSp99
gz51XSdeo1L7ogu8NJktb5Dmh5P8sSmQlh9XOEtKddhvUMYjSv4VoACi8Tk4tjRavdaC8FAYAsKn
J+yOXYRze/DwtdzO9471yYXjUeUTxX8t0tDrs5AfE3glDIMi8fEQb860tQOff7NWaWhDPIy+nhzd
e+aR4HFldY+iIWi1avkYEm/aOOM64O/yNTyFN4KssDY0ayVHYIgeQfvy69J/MYwoDM0S+aw++THD
vkRKYvkrqsdXPSH2hfcN9571ZCUi8cOsX3Fa3WNtkerx+1c3bBkPtpCnZMDlLpjhHwZABjcipr+2
/L1v2xee1nyml+wZuPS12XhjyhsecktyisTqWpBP21ZwyZ4ySICTHZ/WQZom248u8elvvVQfsSnB
A1AhzrRMcz5tBAMQByZLTFt3cSB/LqQ1YhD3uxN1Fg4c3p6VWjjmqkuAjVjGH05deUZT//tYJfQf
OvC0trfF16iY+KwoGSvqWloqDEEDkWQOeeYARJLbNw0xcN3t55frnbPNYfCjmvyQodHpA3xyU3DX
reR4DMDP+0RPsUM0fWddpaiQ8yIWX33Gjb0106KpLZcazjMCd3bm7qc05wNorXEFKB4/k5vw3T5V
MyUJ5STJQ6P2TV93b7fgYojdASxJsVElX02wQyjWpsMBmo4923RG76kY2BJAchtrzkbWdHk8IuqN
HigY7ATEaWSYPqG5BM5EWbc1QBopep1kzBbpQ/0+IkU+8E+i21aDgabcuEFQSnbby5WdOEVOZy6S
4Us+BXXCPuKBHAz8EccJ2zYyZ+gIkukYQAb8ghr0DHfl3aqXvua19qlSd5wzlrsA0VFZAe1BJIwN
QzA386+yuA3oG0Z90TZZe9ma3LAjh26CfdEPkEtQ4/6Snv4uT6GiNzLLjRrLahXVWb1YNd2AlB+7
aB1VgKkYdKNXmI/jrwhUwCbWNggiIB2z0XN1h7llsP3P1QokOenJLGnTXx3O5D/TSW3ZYINcwKBG
epR40N+qLj9D4MTNLuleueLxj3ZlGiuKCpzi/WRscby9LrAp76GcnnFgLyOQd56WILE3lFy3K6gj
kjCk4pfUJB2IMbKrbH7Lm2+nZ0+GUuNEJIQDhi5gDjk1CdMgN+6OwgG1vcNa18bu+nRKr8eIcQA2
H4CK3VOju2j+2MoO9fA+4gm2dIRZpVDJZa1agVCaGGhg1t7YQeuSW82NvD8zE0qXgwpzjleP3O//
jt+MDlSxB8+Fn67CPbtzeNJVT6hiqMkW+8MFoqMngH7PPNhVNM5f3UjIb6hcN3jk03sS5ZAIl4kQ
W86OfLJJoLvxjAfEyaJtB4hnD23iPC0e3ju26F2CDYEzOtlvk9AbbIPb/wn4Vi4G1PDFLlqH2iZI
ab7g+9Y83iWGlC3wBm7Wd+aGW4lEU/Lfy9u1rZxPgQWkC0v6oNBJ3YVDEm2Mpe5c47SmBNrLlttX
DCEKOMjjaBJ1FazPkppyCxtmgLd5Z8hZmQIiNgLbE/ysVFfVV0bJQefLS6CvSc6rG89SzovVSWGg
tdnddipL8STNr8F+KFM6HzKf74iFhIwI+euXqtpwuQ5ig74KUM5z0dNEZlxZ/7LqOWsTNACJ41pf
DYhsnL4unr4vw83+SxdF1+MVRWlke9blePAOWD0Awiciptak0tFp/5oexsaOvp45ss5rNFWGuUYW
Nn7cvw1AGWW3y0ANWs5SkrF3JEbaJGX9+Xag27ribXyk2Ve0zbPtYD+IE0Q+1V+h/wiBsH6IOL3y
xPN5EGhtHujpetBUGDUMoZiY5FsASoC6H25A7Syz3hU9nfSRrsBwllIYj3CkB/KM2vt+DgjPfZ48
hVCADAM8K+Fa26udOYm4Y830+9MlGYJYeWrgnywiecr4vtrgbnxk55eRLkch6Wv7F8LkoU7Myp8M
i+CNkBMSBrmoNid01zF353wFnbpq2WYQhkoWn0jyS19lM/nup0CRwf660vJ7h0cnwUmkjZhhRAbk
P5pTGMcS1OrnEAyeha6s/Rw0+oHFfVtRd3ZQGQh4QI8XjHdTyMyjSKnYHbog1e/nsc9gSp4mIDAJ
1pGeNQsCjoaySUxSy7IaQVtJSwWkOgrHEWnIIsyrfth8t16BZIkgUMlPLDxyoA7ULpaUVIuGskCJ
uXoU/0a4cegiB7Hol1Toj6Xq7o4EcI06hZNCOP2BBUjZ/WrgFlPgZul0rsjzOKGupr4kVZru3H2f
5XOfo8mY4ecpHq30m1GRbBgjWHeaxZPtLWJhPyTWYqX9b7sZ28dDokym+wOf8xMgjB8psvT/SGU4
kfz2D/tWJncYtS3rm3jrcmJiej1UYi3vZ8/VL2FSkAbEraRR41mKAHb05J5ahtWxeQusyK+xXJ4Q
+t/AVYxMyk1dEODUSsTRdjphY2wXXEr8UUdpnhbo9P+OFxF0DpPqiapUTEwJDcY23IYChD9gFlbr
5U8kriZy2qwX3a6U9ZGsLJdZZQxxhEReK5SbyMqigMbkbZUwkS1X6+Mri3MyqWpYf3ENgsItGXqp
2ijjf0XQb6iHBCktOZuONTLG3bofobPUMSfYYw07tyr4up3O2q4TGj4X1/VZTRi5smKmRL9bfd+t
gvGraT71Agh7Qk06Al3rmmn7zAQ4SLrnRmlqQ+CIDLuUbFE5SVlIsMkj+N+x6rZ2VaE4JDLx0fyQ
oUCsoeRtFtwZA4jIt+B0cNLmxpEZuicXwSknIDBV0H52nphpuIRe756DIlj+Onrq5TDvMNpOG2XD
I3anoW9biB1JsP1EFrYlTTbOgLPElDzfY92gJmrbGnHY7QVUG2EldJKHCJzAPrTESMX94ixJg5OF
G3Dhbncc+igkIs7iJ6uATW9cQC/jOnhf9vA75JdO0ZRbknig5GL/OBRy3prNgWmU6P07cAWn6FqN
+GAGl8bgoqXJswd0ZnRyfwSM3vWQZji0Ax/N4RetRz9dH8fhA1t3+E/PA4kvI8/cBzpNkKjWvx7a
V3wL83OHqf9l+6wmKWqXA8WFtNzJc9kBwHQcKQB68kN42Bjt9FN4UE+diJsaOcRRnWDqhTyCcmtI
D+lLL2Asg7qiWq3dhW6RlpFyjHwbrroZtGITt5jCIzr0ZFeZyV7isXHMftAXB8Rzw+hYqVIl4HJG
rivNcuHmeRaJjJisbMVAzDrCaPel75flAXat1IyxhFR5pIO4jhql4j3zM+MntD6N9ecw0UsWcQOZ
v3QHYeRaSdR0k5MfT7ldwYzRgg2/AC5iCU/FNy/X07hE9fL83DwzYSvilYRPQ0m+5jYWuwA/G437
Rala6kIXMImlQqRX0WNqPB7zYP0SdGEACyGcTTjJWf4W15oWbdaxfwkMX6ia5/SBGgCzE3iA1Qba
PuGqboJ6WCVvHsZ2p28rcheAELNUMtNKfdGWvu/c3HB8+pj0ub8Z7jOTnd/m77KfdGojsBymuoyx
9cH1aQK/LkPXFbLF1RVpqh2VW1VVorgM+xMp6Ao7BHgA+U073y7DN/wQkEnQUPZquUNCG+2aw+P6
ZDEojR+0DyQWR5Cdqf/wZCNq+IN7OnczV9cl96Wzn57RIzjgEWAMZtR2OewaThPKKH1EnTeeFkwb
p1YWpbIYxeVzEd3NPga/KX2myXue+FYEniOnFZIt5V4pv0ClYhIKixo4Wf9jEFuIOqVSn2QTEG8K
q9jYfPW+EWLXmG2f19dkALDSKFXa1VXSSzZFx35+aUa9r3X5FPPa+QQkvJUgUM89aGpYGTXAQKj5
FLLriWzvYqtudOATeKqvGtXgVSEMEPlEkAQghNkCpVzSDkrmmMC6ikxz8PrI3aNOzZ367UCRVD/m
Lob7SSZEZQzvzL920z3t753SLEPEaDSRjvb8ihIEoMIXiG/X0/r0bWtnEbbL5B9evgpZ6Zdzyi37
Lor3d3BvXds8STizNJPPFLkrFgQ0C4M4VRE5EgFGCfctzB8yAEeR9NG7SFrxUxx9P7kE9BhqKZDT
X8nlTtJSEv9PMsZK+8+m4Nr9XK6vuQ0KgubUlwRsWf/nsnXLC1azL4iP3/3dt70z+Pq0HbcrK68R
vWO/ZkCbu90IYpFSknIegdFWu4CQ/s+VkqZmYxY4bqUVnD7GI03yxiECd7E/9J4XEc4AWmn4nBQJ
t7xLNyr6BDswqlB+TP/9Gt+PvbZ9MORlYcFbhbVtqtXCn7ppeL+qmi0ABH2plCxVJOghRkt4VGnL
THdzu/VzPCngsOQYcCZCP+7bHliMS4fMZSVE+cc+s5WN1iAEf43jLsi4cCUNeV9NuYZLZCxVSvaF
/YEgz9XSqbQM1mXxMu8aEfmQDMCuB7fMyiLuSD/CRreeElJeQ8oV/GZCuVd+00Xr4MO3OwctdSz5
VAmmq5D9IqYKuq/0iKMGf5EVoYl/WjlSVDMAm77jLoigAHVVUNsnLir9ST0Sho903iLABIloou7Z
qNefTEJlGoFRwMB8+2SEqKX91NE92Wf9BrhWhO9lOKmQ9KRAGZlq30TVA1iu83y+Ch+dFKxx3yt2
8xypnityjA4+B78UYD/begJsoQ6YAfCKekfHH0qM4hU7A3+d79Y3gyoWl6X+oBljzTaC8Ij0t/Cl
4aQ3+1vV1MJQOSeqUrMlJ2V7Yf7O5ewc+U0XAVsY/L3aa8INm+CljF0/TTBUL65O1JcoFe/HrijU
rauPSjao1mOs/SHd02KvlU6oeuTiAwx1RaUDTdPF+NxwP4lVYbdGyLNESpF1pSoYr467+BXcYzkg
wLQDRTEHOEnHegyj9L52Pn+YXr+WdpImJYktFh7BHlrNMVD3jB9ICknlbsXBgswJp/AzY/v5mSMB
oOVS+/iT2vUIAEsYrJGkIsvitEM3W461ZRpFCZtWffjuHCbJkFkmP37hv+pa6rJR3fEvkInyZclE
EUz/dFCMw7l00R57VVmTAV9tY191Z6Hr3WNdxsTD9cz+OOjaiyAk3TbO5T1KCPM1HGl0lNwANHZb
jLSW5Xg/ws8ZvtmK5zIQtCPjQbLOoEs9+vqxvRJxJ5qPsbwcHL0NjBK5X3X1fxlNlabkqtYZOYyo
oG/oJvKBsAAKTCOfRFS1lTRYRrgX816ZSQf7gaHbEdNLPcU51GPE2oXfAkaTtRMW05igMMx73j0K
r1U05tLvnDU64zRnG3CQOhmmjhPlpArEoAY6cy3zOwr1U1NSbPzbE+c/9m5oOkbk2LyOfCHFpm4f
78lSCCzjASM50lM3KJOeA2voGzlJea2MW5SW8NuPti1Z9ZFqoiYgQicMW4POF2M4PtUTuNjjD2d9
1N+MoWcrh76NOc5vi+eVcjJeydexlpyrk102NO0fVev6opn2CEK3J9pAFMCQGL54mR7tA1+5Kb7q
MXcwrtW9g/vEjfQoY7HyVi+F0duRbUgDt+XULYVO4dx9PlK/kBi8S0A95lPrA70EOMT1+/ROm1L7
6Bc0Gsr53xR52tcZKVzXMMcIAk8gNQZE4+CnSt7apIQOtBPYwGkZemPCaLyIuAKaxBZ9aAstYJg3
RNnJosAKThYWyvHVJnj8IJiBoTCHWfKUSNQQzFMEl5rsFhseGLeSyoM8i6lfa5WoGvSNOoxpC+Mc
PB+bPL92qx1FmRtwmKqYeLbEJeVthJfrnKILJn6Jp1oMF40Ng0DC18Ydi/ghKxaYRGWEqcj64+0a
5sO37i8+TuGT7jorL3ZQKtaOfgH6HdpkmTOIvhmxdAUoUU3vp5KHlIT2h0CCajfKz5sM/QJwH3Hg
RGKgI1gLVsNV6tsaKRL77U5eExb/7BGuAgWoTP48FxnHGKLrvn1Z+K3Q+lFO0weJPDKYB2cpRYcp
SqPnY0qzGrOkM3PM95k5c8dk4hZYndrrpk/AoWH6ejgx6UVyWC4KpY91G322WGw7Qt0XAk/h/G5v
ZBwa0u2m31Pxlfl5n9rCm7lMEONz53CUUN6EA3pJSVVqBZjrYgZaF9L7+2aQvR5cejRZk9C2v+No
8qg3Kh6mPvotyIZGiLMa+jhFXQcNUhCg3w6hA3MnG3eyI1MJ+ox8hYYw9DprCh9glAERivfpuKYl
63nFcFbalo3kiHf2sXBOywf3/TM0Y9CnqBZDIEuH9QjZoXxSuck2URCJ55X+MQyfLHIdWdfiapOR
iqrUPfCGqdLTfxbFg5jHrhpvF8zJKS6g/OGfM6+bE/LUU0fxu+yHVdwkvIktmdsY5yjwQHKibxPA
q4SNrOosgpBKOIwPN2tK+VohBb4n2CWGIFXvgL0Z41imClQ9/Z34f52hxUBkUSfYs/lUfu+Aq7Q4
KY6KeOsO6PCi1gLEIBmHgQgpXXrPI2PcbPQqTnU0Hc8rEZGduE8fqNp1NgJV07822p080rciFiFN
WF+MlAKTYd4lUBnf4TEsDb1cXYQWgAOQUYF9dkDtmVrTr9/RxSG+EIN7DDm+B4PZnZeZfNF0d9KD
2pxifYylgpJwIvg0bwsoA+lDcsO57D/SX3pYbBsvQPZJJCvczGPPH4PH83Q6G23adtz6ou2PLLdc
XEiABNGXRzGMr4vmunagYCSYN9irkHjn6DNNtzPYUQ6bapftDHJKgzIZZWFcWCPj3Da5U122Fb38
N7T2PUiklwK3NocPJ13zueCZExq5JRUqWHfcGnGRvrSuwZC8IKpexJcQEchJgnRlgsC1lMCGGn0I
yFCoal+cQM+kllXZJwvo5HeRsD+fIyLdU67rENZYISlYd3exsKRsQJQhA0yxMKlH6hQ7+RNd2wrm
l8hK5Nn43CaR5P/1JRP8F7Zj2gnQCzBIwFJsbDq8W+z9fwrWhzCy7JirKNB/JtWd9HYqvdvvVd0S
EqbAmajqGtB3XL/pQ9JCsAy8Oyk4Geju4+FcVX3wuPVewrauRfmb6cqODaQ2oR3ysBABEHSBmBB4
FaeXBTnwS2t1bAfzYn2+HFQRM6/n1bF3/H2TzvW1NQN2S/JUZB2M1ZyDS0iew9TTgFnCHEosQ6+y
bt3ZmtJeAxoUFffcqum0WT1oeWdMVNiwEo5fSyKVKmgvx6/H/A9kTK7sJVazi9cJnMXm9lhI54M9
ethCnh4rijpLlX53bfAYMI3EjkZd/tD3Rgsq0MMfnIj2Xg44up4YRDl9PfL2GKsBR9mkKr2EuP2/
yRhMDhx3wIH7pjq0T0Hds/npWzfO0k5H3L4tR/A/upobPxKlZ/ca+1hgx3mH8E2bgXBkiQWroRu/
JRekErbtSlclq+rjdVV4+cns1JkO+gCdOFOZlwWF8Eiz9Hn7RahbbHDDHwnmELGqbh0kRr3odSld
6UdTawVRRpKMXcAIS/EInEg6gyyOtRPsKKhaHZNfIc1yigU8hu7f5wwXTCvIhbj2EfhWLYjDRyn2
df02py1cNbBRLhWMSDzQ1VyuK3mrv1WrJZot4tSYqgsjsu3Km7awDJ8JoCqIyj0Z173iAwgJifbK
oatHvC+50rIQzVbSr6oCdck76n/eEmtVG8xGN/wtBvH2rDrQcA7UDr1Tb7CHbFbEWaXVaYFzXmgO
va6l4JhppFlLI+BYlhuyVts+bTkCzh4Omd2THm33zxBV3dvCgcBFz4cjy8XAv7URF1XeDEN03BBP
Up7i9jRKUZuBy9mH7HmaPSNA14UQLL1Oxv05RA91VLSalAPynLe/x58qsjMvSIWNuBr9NESyFTXy
zFVzAs6zyrW3eXPp//olZQ/2dMiCVnpE8+Lux7TNI9Fsu77f/dSvcHCJmY85R7dmO9jMNp1H20V7
W646QCxGIzlzXegN0yXoeIkYDlVZjda34lozH2ZaePXS7pIj1AMt0s1ruCUSaLpgmjeNa1XXauvI
puFyb7XLBSfNPy5UgyHL5eYyEh1YYoBUfKaZwwjq9ycuqNwx8yzoEShOD4SloZdYZJw/thE8biHv
Bd0IySrX4heNeP7wb+UyYJoy5whW48wd5SwL9UrqV9NFcCk5nmOWJ/GldJ9oevHVywNCXRweEp3T
QxrV90YFkvnc4sEipSrfd/4/mB9N5jKujB0qJxeALGewfWUT9OauTIXK2wriffnsXBH73aM3PC9v
pc8m/BqaRnF9WCOlKejocoTqdc4JbHZt/fRWAQIPOAzCnsd/UFAMofGDzN1BviC3OR2ZPrk5PD1E
nfAsrhKmfGem0TWkbbkkFI5nUxwYEQbmrFsxKy+vtSXQonnp6fhauAL16zuxYnxPpfIHTdf6varf
F6zEb4XGxvrFU2mRNSwuRsWi9gVX4MConeySR7lS5dX0g7EGriRc0u6t8MTqT8tPzDh8puO0NPfq
CqpiizrvUr9gNV+Mx/kh4YBbsf7rtvITNoo9wIgVvzmmbiMT1yNSN2lNzmx3X8ebT8VCkF8bDHwt
tiYS+3JEgtRDI4fIgRH88vlxGlPbf+QWxCXzFi7WLs/6gSlBZIFpGeW+1/tSIXQUnVrTZHxH0F9A
rKHpo8sxV/N0KWahqVJlJEjpO3nIh43tFndvas7aljuzfZbeaJsnD/OYdL+BvMCYWq7uusLKOoXz
aNwffz5VrTSnFloBkfaDPPmBiNXzyhtEoMhO0JIiI8wNJ6bxKVbnTHy/romIXqZUBXbP/5ix2XIO
BxHuwAHnsc7f3BNBsRu7fpckBrud/WHt/R8SbKEHxilse1XFkeSMYeG3X0jv2ztSH2wmcqa6uY35
Mqz9dWDZ9icTd8w939C92UpWLC55bB4nqO0G36soIwGQOAkPlDYZYs0Pkrbjh/kvs3lj+fl+yZyi
CQG88e5cXBW2GCUAhjYiNC3jfMK3fhSDOaBAg86/yS5HjhbF/yMM/B4s6Y1vQxXcdPKhnHSKMCX8
GtRUfwHC3adOJ5cMoPFo8Y5gs/gQypYft/t+6ZBytQh7jH2QflZxpOEIFY0YUo0A1nY118RnNGD8
5opr9IDp58E/EYH6tr7hkzofXIA6vhLrWoIp0H3H4R4OUnESt6LhGT3OVUSEAEpNdZFPe0bzn7bZ
QWwGyhrX1wg0xm5pakuNWFwoZikdqPUq1+eZWceINKSjyMNujxuhiC64olnG79yEpYxcHGEJV5/T
+UyvopY66bl8r6euBCZs0ZcuT/83WzTGw9A3LFUc/THcEB+ceoFQfYJJ3qZ34TZv0NgurxntNfhC
B/FO9gvclvL67r0Nu04CWFFTMSOs84AZ3Ek6AiEP3JXUpPWLIoeN5Md8vUbh8Q/SotB58io05SOs
2yk0b1kje2QvXXOoe2wleq4USgTR5TXWJqob62RpF9HPIgjN7rvJbcx+upYoMK1Wbp7UuOryjnxk
EwZl+t979twHtZqdiQyD3YF0YnBk7RrXcGBBVuZJDCkOespSh2TJTnWR5088pbD+x+9NXamim1XN
OExKjkTMDLh/trn+k+9xljM85fJ4fq4eqcMQJtSsBnUVVQ1No+SreUFuwvFBXDeOBwV3+KdGBs+I
sPnGFyQkB5AOMLbj73QhA3BE9JqjGwS6QYyJh2ZzYbbXXXrgY5xjUVoUfn2Dqw4Y+3P0BQtbrCkW
8+szB+l3dUiqYx+J5IqCXXIGfEUL2b+VDZsVyUbiGFmaiFXWzn8O32qKwVhkLSGDIA6i0MjcrbL9
fzJqtxal5Qqtew6wRTkOHAz2EKkIJCjfsYBqBZugrdBSCQ5oQmy9Tq+jVCq76xpzhiiXleqevgwk
788mpR0MlN3lKuWVIv9mmzmbfM2vvqy6fzxA9Y2X9iQ4kwVKTDk4WKP6zJPaLxQ7qFGq5Lb+LFXu
K3IDUO/C1TsaH8r9bDs3JwkTSBDZ97RjX5YvHSorp5LYXaWx+4Cl1+4mHA3+ejHhtNzGED+8xU5V
O3c0z8WseG+kmrPdz5Rs1eAt7ja/AFj/eBCpcenckQAJa9a1CZ3LPiwtJtCTiVdWSJ4l3x2oqNay
k2w9FFxLuy2F5nR+FDOleaVnQPFouA7xaT6kKofE9lAVKF7cOaA4VrqZEeT++hANJVF3IUpdTycf
SVmtG7NKSF1dOpI9j+zqDMRBKmXTXRybARXvzu3nvCQtHQl1qPWJVT6CglacM4TCkmcAoeUL25wG
Ib8dnShTF25WiMuB3OgBn7floDuscr6VjfgQAMTYsFsv6MVbXJCKqvVcXmukfQ9MKW6wkP1u04cc
9TzzilD8PX5ZKb5LK2VEgRz0z5iWCQ7FphApQ63poxruU1DaRzY0JTUJ4+JQxyQXMjk1EGiDHS4N
eGrp+l55BkAruZu/YKDyLFgPksqnkK+nKorqq7GB0D/4gRwIR9dHMz0DneeDPNwWpAc4NEbn9yET
ozEYmdvRlR3AOb3GhlK/Op3DqpU8dkJHDjULKKgFWvof+nipbWwzMLVrgyoQr5f+V/7boI5sU0fw
h7AhqmVYm/YX5sMwT+jB9NcElAZ9Co381sj86EwydODloWseVddSEkLocgnxlR0ebfsyXyy/lycj
cgUQu/Iq9pqrspBI7rhgGzqpFpUwg8SWrg7fG1u0kuudMy0AXDczKeaup72zrcOtDpkn5a8q542T
I9CelwEECL2RAy3Lr5IXF6dSueDNyTJPxl8zK8eq1rDR+43xNjHRKXJYUwHyuYE4hHVhga2nhNyu
/45FYUFWaxDGBjDzokxKswJjy4x1rUNMxo8Rv3wN912umn8KIdf/fPOlKtNAzaZslq+R6RPj8jBU
RfrarUB3rIZMq1KSjd9ZF2rZobo59vYtqLWjvJHarweRH8HoHYIFaSkv6nqzz71bl9z2TDrMbTF5
T2ZdDCkpO6K0gALnShw6L/0j6c0xhTZ43vypIMdYjUxWt7AsKisgzezFhnEupgXrmJzw1j/qoDzv
OiqXi/pOBgkY6fkHKbMq9FBvcrZcpf6hdbBcU+iiMe33M1u2Rd8Kxei4WPp5PhtYsQJK9mwm2b7T
mG+LcFpVWvUK8P/PPAnMHO0Fq+P5qcSpX/ELpzHC6VQMgsY2drlDjehUxunS5E6dsr2ZIFZyPsvP
RFBkqXLyGzv6t3NQ+shBn08xUI3hGotyvNgyef1NvBtPhbZMb7XqMbwZIRn1i8QLz1wd/az3PLIl
JrbRmF6dfW+mceeaGT+/C1AyoOam8G3ejq5geUMQHrWQSCzaO86iewwUmzOOfdtxA0ntHI5pSPbA
45G3O6mMxQnUr+3ZoVQe6X9kd8V28nonR2acyA47shgDkF0rZxDM7oM73IFaZQhJM31bytKQ+85w
ZJa+F8aYfiCdnfSOSVhAClBpyCIAXna1DxlFIiI87xqKiDnXAAaxhSPFNnIbDkfeL3+jn5m21iQR
iVIxbLq1dwIHPcwzzmqFeTTmaL6D4/pXCru9uhtLeYO9X2ZJN/HPc/cGOVT9q86/2hWcoka7Pabk
UBkU/1LS3uCwf3gtUmPXS+hCDJXLr8l9oXTqWeHfPIKqE2W5kY9l5CQJrDCMe4KbpNzjBEZL0WFH
pd2Tf9Wh7AP76vGjUavWeUYLezthwVse1UVbf4yCK372iTXt/a560qMeaaTRqZggWmpN+uryYN7p
QldfEn6jCGztSpOX+t+ONvzjBKGWGqqU6yX9i+zdc4Uq1v6RJD/H0rJ5AMupjtt6gMqLouTLF7jI
gfxaOmQWD8rufSTSA5aLNjdneLhEmGxVD1upfT46BIL05alaFHsw+muPG1zbxnn6czPYe1Gdpqm/
KQNGLqdii1SfX8I4fDdDZCHGK+QOVnM8zkhEpFDnORHqVPy+IDqP7fxA3RIF43P3MA74Vt9vrqA0
S5jlm67Tb4eAHR7xeQQNVx/CZV8PDeGe7vBpx4P9nP7g4kfByuOpyUoKWI4MDpHEy7ApUIOrSihM
+8FNh+Ic66G1rur4rBp3x8x1OjsEU0zYK+QvpkQ5wohpda3agniaVA/OrHu96CuglY1GXWYmGtpd
QqmHxgxyUyZsKg+1RUXs0LmHKvegcUy61L5uWadlnUFGfgOMrak8sLq1uYsaXH170EKQ3CLcPwOB
zDzwoABjGKcEd9dMxo659K3mko4QzPDM/6lAenPhVHG1lLpi/KHSUouKoYVH9PBzr77p+dfFIECT
ztnSuHkDmySN+6fryFpx3empmf1z26gU1FJIuR3Mwv4u11d0CZedhYsUeXfr1RLGxu/mr6wIi48Q
2zPsuhMrfq6xjCzdpGFDgcnibkDGNvNZasuW2TPyX7G2mB1Jbl/tnEZ+J49A4hv6kp/78eLHH2Nt
om1p0oe7tkyUPm90Q+lDrwTqIRz++A2c2tQ+nD7ofbuRYAMYDSiYDYACmtWEGFPq5/MemGdRL752
2TIapsmb6ZQckMflgUIr5kgYvpYFtpGp+K2tOhjvv1QUvWnoKVFTpLMPbCIsibUcUcwgRWyUba4L
yiW4zptfYqN8hOY0efEaArEuiz/Zsbr6ujGu0MRWLZ6zwtxDGur2vn13DrUfRgXmhUw9rO82daHs
AGkZ9ALB0bYimn2RygCFYkzREU8wUi9A2YxE//qih3iAib/tjDchRpIazjJ+eoN1fRL4W/8/FCx+
0+qX9eRfMUVLvGlqe/OjQ1/QiONlHgLbakfYzkqAY0Mo8BNsiOtWdi6sGNXr+WHDcRukpUuKKHxw
vhjto52ecq6mpqWPWJ3vTyQoXFsyIOBEHkVUh9aCkaK3T14Q8HYeOlLYgMINmk4MmElE2np4EeIn
UV0U/cb/mWMNDgQBnDudjyMGFlev3uzbnYGUbiVA49ILgz0NKdc2peA+hUIzSzqmU4kav5Q718Ag
dYk2FCinOcmuS59e7lbmXDBXqOIxSu3MlCCrpN50BZ1al5YKazVL970P1mRHjSzzXsW1GHE1CmY/
KrcFj4js4rcmsuSRlrCmgFA/koHp2oYEpRN8N3NEwsgNLx4KCCCsfEZppoy8D344BbheaODBh7i7
G4xp8CTwowdlv7HcvGoax2LAreAGVIyuFIaYKogZRNwrGbfA7PfiCJ0+59nJZzYuX9VVgJi5Pk1u
amRo0x1YSda/L5+2pmHNrXhXTxQSReElfFdZamgsywi/WOe4M4Z5tbk1XqfWAlOEPNixYB0LdyZf
owygMmptrp7CxeZCMgG038OwoG363VCDSc+fQy5q890ns9cBBFd0lsHUQ//Q9LSTyP8YkF+s4YMx
RmqoR5Ac+mbtIAAn2NhdV9pEN+JFRSSJDMjegndAaRnbyr90Nwj6JrDz4BuINBTd/dURUVqBZOp1
/KcaOKEtomTIYKix2yxeWvymXslestj3HgmPQLRImtuG9YBa4XLa/V6r4TSpyg+/Jf9WYwpS1Y2s
PoS22DTGLWIL0LT+z/6NHfHeWm5ZPqbnmjbhPfNX2jwf7AfB9HeqWnhzo9KoElBdReHyQ/PkQeIs
xJCFun/i8E0Tj+KMQU5+pMCDkla81RMx7P22hqBci6KbjIygC7B+EhXSDogzgOb1IYVJV6byaiBo
4qBeIimEyLxIBi+jH1ZfAxiGusP2AS/a8mqkiO+Pm3/lNzWf//lF1uUC+Pc9XR4h/E7zyOCdL/M9
73RpKOqiV2vB9Q8FbBFJc1wnz6z4LR7IiReyZhgcEYUVdEFHFXYlN5Fyvhiu++j9qqy2OhXDza5y
HPzL11Aj2cQ/Tq93/w9bz16m1C5Rz4ny95xu5rcUpE6Scc4qBaJ0/Z25fGimizNrqinJXbjCCVlZ
otO6vzQwgxMNmIeffDKUMiell76q6M1LocxPDnS8M4tZZ4o65wtxZEyAQztBodZOyLhu4P1oJjy9
T8fM22sLfS9l1eaG2tFWQHcw5jQLXp8mLzRMp3GS0x6fkOcOINp0etcpKFjuytjyP4ymQjk/24qF
FN3c0wcbxAGihM87wRmy3gR4/GVpyj2FDe8FyF2ulz8Ybi5Fj6JPovaToHMPD4jjivjZ8haUoFav
VU0w4URSKVD3DQOf1VkgzT8y8lLbD4Dr6vea+FqLv/iJ5Rij6moroPWpso8EH+2mPz10VWb/DnPF
klzygvX+KuC/bG0cf/1cBNCMyWE+3ExI4q+BnyjaCsd0lDihwZmmIxefz4NfkFR6z0fKb1yTE/vd
p5Ubv9mWKyzFDX8gaHwejs64rKRE25mzRaqsLPYWROVChMFzI6DWOtHih6i8fhS4vJPCtK9fhIia
XfNNAfl7JTKq7IAOvOxnW53hZa6ywO1WbB+ObtaWCZGEmt9lQJvxdLuofD1Vg0EdgoEZ/cPb7pNl
UavTqLP4M5PPxhQ0k60MGIf2Rwi4pY5Ki6AVCTrs/+0Q1QHZosfQxQADvFn348c/5NIWo5vuvAr0
qMukOkwJivgdhD+/sjvyb6SrroAFNegay/L+IRSSdTOxWYlXO1eacl3plXL2vdPcKh9l2GYmEUVJ
+EaX94Myk3K2qgYQjr7XZ7b5xsqDOmo4Y37YV3kykoOaKdZDvD6zcNUfmxORgpqDQhO8PNPCGgVM
eweNtVtrnC9+Vr/a3dcEY/5FNLDdDYaCfQF6SASC7LLuPqvgqhUFSHUpwn5IBQ9C9xbHcg6UyIL9
QZNGbxAgTCOW1sVtaEqBGdQUOq7XABNF1hCcFBlSJIAS3eJoWxQAf9l5NQwI25iG/c2F7gnTw/HQ
J8eXzhhhTH2v2NrwZlrO2qYQF/5bLYECxkDGQ6m42MDKWiYlheu2UtPlTE2aT96So5mHZONHaB92
0hM+pWg/TkzUw98OwORbQFS9gMzO6UlT7qscQ2uVh9et7xSu7jYsFkSn/iZo1CWdQMQIK76xv4Vp
s63/8/RBCLBNa/dI7f0/pEaEsr2sWuwqPxmZYWotNrwKnU/gU/CLec8nSw/88dyhQtR+Axk5/86Q
opun/SzbeCQKLynx67IjFxnoe8ufiVjnXKq20BLLJdTNctLH7Dq24fl0ZD3zlpdYiM7/RPGxMgQn
8ao+o2O9pK8Z1c1VftkgvPBFdV1Jm9KGLJNubPhnhr+aWwrLQK/QSYLhCrA6uNkhIp8B6OGMC1Vc
9IAUjMjAZQiahp0kxmBz0jMZDsGEzZrntes50p98z2YzOGBac7cP+C9878rxYbww9ySS4gUt4lBl
y4YzK7J11HmsbtLhtXSEvDY+h1sWlbIs1+Jb9G0QoDo6aaVAg8lqxf4FiJpfjPIgyueMUrMDuMKd
J/jxdjEbi6MqSjWa10rOtzFfYWh/f8oP+WE1gWq24kBOgbIUMAFAgjB5QCoGn+nPSqnFMYjI6ea0
SM9AfmhuqIxo4DzDCqiE0LUdUhK3kyOhP7VnrhTsiZ2ADcVyUhTHiWXU1dwouVjES2cKdZRhjllT
sM+yTju0uACNYjvZVbfBNXdrIlMlY1n3t/qHeelybaz0pd/X+V+vvKtG5vXq32atd4OwVHGttoZI
hIUS2qlfPAUO+pX7i/Dmr0HzPcQydmx0aaEf0cvkEx2fQtVYU6zwLbJittvcpoBN/CspCiwUtheG
5rLYrl0SbRpLDZa/5xZO76UCmsUXRSQ4slBndmC6dsd6pWmfabYLoNu92XCQH5J0uWDH9P7JnD+m
R5bE9HGfly2b4mB5NZmNCqo36gEZPS7b+kCJJO8OXgwBM//GAEgwM6uCwOiKeUSI5YlnhJdm1KTG
3YtwraV131W+A87y3SyNQe/ynYmsOH4cuZLdMCFWxjX/m0zhhvjxQozEf4W+a7LTrXkv1GL47iPH
HGxFglIyV1jhUgAVA84bmYC/GTcu3+AUTenDgxqltgD/T5xzTr25W+9QSygWRwZvLgRviGzE9J61
JuFKQheKZHugD1FiDeDJSQO9O4Dq1xBZ3edlwj6Jstrs5OD1i350mlUXvjw7SGWQqw+i8YzxRk/Z
vHfE2W7esZy/63ixEHBWDj32968TYSyfw6Dd6TJewYddKRMgx31jqYZZpJoLZNZ1pjgHxWnJAwpl
uCUwuuZr+R9DzLhukq/IZFRqnKu1FydU34xDXfKUPMy9fRibJ1qm5sqxTlJYwxSMo6Wb+W477+T8
ALMM8d4IxSyFhQhlYcgRaqAOnzYcCTY+EQ0zuDyp9uTpiE2N1Ubkd8d5qXgtFoHln9x+7GxmnuDm
NWRTLPWWv1CkMTjyFRWw5d0CEKc8VynDrrlJGYWVctaBNfxsz4HUKXNXX3oOAvi0zuMQzsWmPTsX
6WJVvvvyh2G3FIvu2i5VLsUGbJPn7uE+tEqColYm1f9/sk3bFlu+Wgjo0FHdVU3ct6j7uZSYvDMR
jK/bjQeaN5R8cltUvrMi0X3+9MEfD8fkpWxGttVK5bBVK7Fb5VgsVsR9Ub0ejponnYTWaktnnfKX
Aq+IiARoQuCx2nNwEUgupTU4JHN0DRYS97eXnfC2gVSkpS6YoQ7H5kILUV/iQCBsoWftGIqKgcHK
Ru42Fl5/q+CKY6SV0fPFfZUQyW+qOCk/1CU20WUIPbdyG58aG9yGR2LzSXZ0RL36fC6DohZPXSEy
AS7m9Ve04vjahKZbF5HKRyd5qTWALWBRkEQMOq2RJ/3jLONy5tB8Ro7F+QCvFbUTh/vV9GX+560w
usFLMYEp7mgR4Frtw3EzfX8qKZ0LafQd+7rSK5LGKyuqjDZOL4trntb0sXlJqUDR1Gt8sBKfnGaS
wbD5yEQkxCSooJfvEo6UeT0JHFVjFGoMYjWvopgIwu4oZ+ksM1HBaZUqb+Da8WbFsQPCnkimNZa3
1KR1nmnJIllanIIE+KQIHkBHU2Ws6AG2FMLSwg2lKsyOhMObhECSmm/KIxGGmnmGLYULNyxH1Zyc
jx9NMoaOer8kwIZl9j27Hf99J+Xqsw3jSGqEXJnsHwrYLZnlFGB2cz8sOBP8pQjMheQ5gF1yOoai
rN8zlF2KNcVD6AIYh8Kb3Wh9vl8d+QRhMhKTxr1doTf8S4L+W1uf+I9aaMXR2+cFQb8pZ6Hg7sQk
X8JY3whGw1HIEJBhjnZ3B1FcyCGYSJZpZB+4f+RGB4PqLyHsFHa3lUJZNwvsXFt/ihe14eEKekud
dPTYcRWsBGF5KGnXPADKFXHkRsA7gdiYDJb7RK+5nfle9yRN1imkln+JS4r4ZAUW0W4LXV6M0/Bs
a0saaFzs5ujivgrRRQo4nVzx6Z7O5ySrT87eSkAbTEXgappvahOc4l6gOVWjSQ1tRVa8N3uP6O8S
bRY77m2G95UAufueIgBqCPLF5a3EpXVMcgNWYKHINfwd9P2gwl7A8iLkD0dguIyiG55uqycjeK1F
4y15weVZGipttVnqibaIfZrbLoCi3NC41QDMYT4CEszdyyU9kETfXjKMyvymOVJtMdi20ZVQzr9D
JFkhGQxVUuh4pjg+ON5QjLoVgfslSau00407krJbAe4S9W3m/yw/TaCEGndUCtr4WkwFV+zy8egx
Ti1KFEzAWjK8Jy5B2dGm73Rdc9UlIqzGYb4XfqSyq0pAZmNWEbnMspduzOu0f17Wi46pVKMZ1wbF
YEk2Dc7bGF1QUp+4qsXiX6eFFpR6uDdZncsR3lAfe7mO9+xXcAhMMAw01uBe2ODEAzNevNri+vjU
LRa8yikKOCF4hWTnkbCVxMXwdRcIs4/YizwypmdQGsPyYNzWLMidseHddhlnSrapBKopKQCkDWIF
7ZinHrQj1kALAIpQKDmsPvGUdZPAM1OTmGetQflVGFoWqpCYB+LO1ve0MUc4wjIPvyq7xwvEaOtu
yxnt0GWrHJM0sBo8tZdJ4O0N8VfyBtAKoywMrr6SKx7m7oS6+dwJk1bAjXBmwIkW7mp2H4TTVzl2
hvA/X7H2Yj7EdErIYjJpgMtWrZa8YCfBfnWffBBJ/H0JN6RJz1GVF7OTUbOmqzTnsEuwx1H/b1Xn
0dQhvZZFyRQwH87JRlfkSCbj0Q1S66BqAjeth3ToyWjW6lPUZ0w+fVXeD2aJx8G1JSykke1e4/pH
sUNWfKXIMe2excAtKGWb1kMuar0xL94Xbos9mDwtzav5zVseE2JSMgglOAQkBuUx9t8pLVbhHW8M
lIB9FwNeXsAXRn9e7O2t2yVQuZS/kwrGveQ/ClssqDnQKskfLPZj4aB577EcveUtQO+eB6SzMcLl
bIP7i7qBXF0RwWnDw53s0j7Lx+u/B6+Hetc8246yuJigbcotKNQJ1D77omNSGMFnCwQpHo3jDGvk
CDuCCih7v405jv78IoyAm4g2cPRtYE6vO+VcPgnRMfsmhyK7Lu7gBEHr01Y4EX77EK4hAxhTDiti
msyGt+qnzQUspGcDczoWJ20Kak86OcgSuuvLfVJAqF+0CRZwd0xaEX05600u5S1fZZ//lIskDulA
fYUhyiXAMbVgCuZ3J7ECa49DSWHcoIzYxWWLoKJVZozDWia4OBehdMWRl2tthnUd3Tomjy+YPghh
r3finmjALFhHJ82WkRgYInnBoOsg7YJEKLlCSJyIk+CqPzqbEmujDhgJf/mlrUS8v5Ye+nm9i2t+
DZUScfqHhT5qge0ExqB0JLUNBT396k2RDdMpi4XjJPaaWXeUAfzphUUHGXjUKL2x8I0IiDtKBNnA
U4vbajZj0tJjivMmCttpq+5RFKXqLSgX2e1K8KedppM9fS++syiUcUb0eZbOMBOGF05w12J3NJuu
jVOub2MX+YHKWExJPG9smY+UeeC3rnXDRwffG67BCvnwieJYb/HF/R5mSkWkeIZ/kd71j2TdJWdi
VaePkjUQt/BmLwkD7Y9Y8feu2Ky+tg7WOQv/zOHerpyw6D52/y8t/YTfK+w5t3fP/P37BA3KmI9m
ELSE/OlDTDFNxERCvY7lEJDPJSMaHdeBeB+CKigX1wjE8PeF3EFiJp2Axuhidb+nQ7/CnRAv6RnX
5U+9Jp+Xa/L+ysTLio5mtWzqAMJQV2fc6gdscaHKYNgZMwYwoW538WkxhCfrQjZ2LuTrD7kkwpzp
y9S4aBEz6OyHE5idF5b/YUKJljIWW9VGtDXJNOvbcARiAGVMYg/ZOQZRjiJlMnQxGcabIzo+X43p
QraDbL+f2/aUb/qr963QWcImCqYFUNLFcd0oTFlGIuM+VjTF56Ai/bFx8IFG0oJkmiEVLUs+HZXn
CMzXVso44KUXd7azq/clHBT1I5KLz9ZVoZ3Drvz1aljXRKyVLaP4WrDmS+LmqEjQQDiAHUCtTWfw
ZUPrHyKiKHiP1XcYOWUqgraKKLx3ZlX9yQ/rA+dB+E1Q1/5HTT4Tylbic6/HBhids4ZJcpclmrVR
eHNEaM52YFiVggCMcLmkqsU1TzgX3beTor5iQi1894h4ARsZ8iPrCN5Noj8SOgSHiCo48KLAdPZT
Dai+XaMcIUCjip+YH6PlieKDaZ2Ic2sqMKeDJjvpqoryeLJuGSOhkJrbewGxTlakeKyE1FvpYRiC
YSOQZkn1Pey5ylyDl4D4v47KgwZO06rH6Aqr2tBZF/G+FCaNFdmubEgqPMV6M4J5NIBORrNhS5T8
F3qu+FpSOmiKuZLga3tb+uMGNV3Co90/B6z3tlOjiAsVR32qHCUggEpsRs5E+8y1nZ8oTm0YMdJ8
r7DWTShSj+nvUXn0HUSVkoOWcl0lnHoGCp6bea7+TvDksBqjNdVR2ZVvIlHub/lxyPgCJgC9GH7j
8md2PHZLzwvnqP8+UQIdN5cqPWiQsPq24fGLce7Cz+UpsFSXS1HELks4fEPm8zJiaZOT5XWr20f8
/eaZiKs0Cm1+6YOKe/WvJvYBKH0V7eVBSMCZwidLv+ybfcIHd6NoLnfQLer0WC0RqyCqR+umR57M
/OAptbeopW5bIGtK7W01PSgdveORd7sZk/s81DGUJMp3SqWo4cu6hZSAtyPAauLKoSR8hADFZm57
1TKrEvng1IWFBX+2Ed2hCWj6HbMfSbXkA/+qqpo1CZLNVAQCGBYdvln0iwH5J0cm9O8l5N4OQTzs
fPzKt2RjkVxQzfBbIgemO1Wvk9bVmsTEpRuA3Fzn8S4wvKBn8z3wJOEFqtI2PT6rQikJE4nfPePH
hV8kcH7N6fIwxfRen4W+0VRfOWaQuK8t4Req5IvVRYFinVqRbxjcm53n9QVJYcMRcQ8XdIhujkcB
FFpE0Mrq98tyXvxRY/7MbcOGPaJHoLy9UC2E0tLBJvXorPkX49lYtSQRQsTXBr1X0enweplJAiac
9/v3ySqlLsfb6NJJI3YMHUf8KPEV+nIe2rYHQ9h/TIllSslWwoqgPqzAADaC12i7S0UycvfgAdrT
Fryr8cDzOP/44q0JAAZAvTIl6WVv3dPyFYuOCjd7e+1HaD8eIzMCdA1eyfnwZA4mWc+PCKkyzJWe
GkhA9ff1eQuAaTlPBqEYsDF05f6omsIinfPpjPQAsgvqTpztG4L0V19yMFdZnZgY2e18+nbspWCe
7ROvGL2NxsWbNSokxHOCuVbr4DJldLCBrqoLZpIlNBf4aT254IQibXuHcVHonhMDWr4DIb2C7rv2
s9zfUxktIXF5SKbAJ7htoLfmB8VyhRXAcNqYpljP3N00oQkfu9HW1I8qN9L2fHQgSs7NCM7/fHli
4+0MWWP88mnNlWp84XjuBrihvB8KHQh22fD5i+eL9KRsbfNmfD06iSTKH4KREK0euyPslAqY8wz9
PlrJ9HLS9eFPtvh/P99kJcEHJCKf3TScOLYPBIyGt5aNBJOTY5LyIs8O1WnFg7k4S4uf36E5KRbb
dSfUzSUTPquBsxHZsqlQSzVKQf+SEvLnOYL3tqTJI7ECJkwUVndd9ENfRxnZHptWSjx7O7HQGXZz
TE6cn5LSnpFwxBAuLKExPzyPQL1Qs6JFGsPSbkBhEBnahfcZGOveQ2fBWa+8FWwNemRHSP1YBxVc
99zYtr1ERUtYG5xM5Gan+3815Mtmokbd9sI3dWtCTzJuFzGA4qxqBWikFK4j+IHzXFEp9ES6DoI5
mt00A+B98FtuGy3wf2pc+QXR2iSS/QDFVTp9jcAMw0p+5UiunWCrRBULMJTbt81WGhKydaaf51bF
jY3fdT4wpeR+UhaUZK9qy3tNE0ILQmYjq01ry13gq7Uv+KC413A7zt/BjDS7yiPsySZ7leX2ZdEF
YqupMtlduORncrEcesmGlieuQDKrurwqFyssHA6L8GSI+cEk1u0EPSqBpsgKSIjV4kLX3SK0r1WO
c+rT9TUaUqLp5ziy1MC9f/MwlYqtFmk5H7rS1d7BAwCnUi/tO5cEgpH7qyHBC/iK45rCcmcZVvNt
Lo4oNZI9vyBNT/dTDNa8yxjJ7f+fkYqtcGQbFK8XPy7Kbm33dfj/AiEE2eUUR7KsVxWWYs3aW8RB
K6bQKDVWTpUiNjvm1ekVvbs829kdG0SjTgrNDfYUh5BxzZMUpynbss1coIpXKqHa+qxP3HhF6e5S
37WyDBROLSEZ41VD46NvlfzmNW5kd95fvkGnYiMVHpjOe8x6Ax8UFCCkBpBgXFgn/B8UP0NEnlSI
rHpPXkMWiizoB8iwvey1ITHjFdUpZZuTIRlRwo5c3fNcs0Uo9v1r1fyy58oG4MbmDt9dZ9i1s072
azR4j0ZWa0QzI9fgk8plXUxO8escRX6n7SeVdBq2yg7apYd+GXg9WDfY2yd8JYD+TSzJN/BwWMb9
RZC6q3CGWRzF8ZdvNrzAuMWfQCk9jfs8D0YcpZr4jxCj1ymuahFzEvNgGSFpb5oKde66K0qR6VP4
RBUKhVFUE6YmUbknfq5brQljk3nJS4m9sUCSc33dxiKRKTM9o1fn8ntoaqoRXhXKAxFayV2cMbWx
91P0qlG9DKfw8MkH5b3EYDVGqSV7t3/j9PZORY/EfV5mJWp/mlllelSdKtfk6DHXF5ii/V0U6YJu
T44lKAcYvAd2fi4BeCycQ3yHW+XCkcY9fgr+28Dl49Ot1xTLQdiR3ZDUnlkJDd4tOmph3oJskwWu
ccnq4rHHu2UQYc/bbIOBpI8CjKKQrVijqRTWdCz6rDlmqBJr1KbXerco8MHeO9JGiBuJgHpfDuq5
NLI1TCiL2/qCPuRQMNeSo1PChyHKQECewFjcJ/8pcTpg4MAYhiTVVMv/5sqa4pys+J7csIVBOZfN
d1C8sCJKBw9IlbiJi17uiX5LR8c3WgVqRnqBf/H7pA52D1qbervFuBT+4DodsgXm2qV5Z0K29gbV
g7T5YGqvxzBWPwEZf/yIXnpn4h8zgrIvla+NMquhV7O0zLcuB4L0nwjRuJP2O74BGj0FJJIIQxjr
rF2agDE7BfRBuSd2h8DwKemqu6xFl6w4Y9z+e1BTUpGx9MswuT/lFQTRwwfl/oXpYdEaxQ2gh3pW
TtKwrsTRc1ysutILFvzKbO3I6IZJiQWyucvNSUMUWRwz6zEKcBX7Hve7xCn+0BpqK5IlWAa3kDmb
FEsN7FTT+Mfdv11SiQxm7EtBu4SprHVkXlKGxJjIVJQQ93/WXFEGmQtwOYa24hrDV9IfJqd/bFWZ
tyhR+Zn1QK8QzoqgIWDKrCX6Ft71lVoYXBvqLOoaxMvWjuQzfTdVg7OwSkDk2vBCr8dQubtELRvL
AQ9eShbwiFNHMgxhBTmEp6G6+Ggsr63gOuqh5FUq/2390sgLmkauDaMQ5kGJLTow/EdpryemswnR
KUevCWtjvjQ5Y7vwzss4l8am3fC6IBjV8NZi8MTuXd7RGJonFLfEhgmeoyL5daPGIpQs61HpQgau
cQiVG0X4Fwh9rru+gX2H8tm9M84XGdylqP34btAtzZ//rSup6O+jO/2QXOKIK9UdvFOFcZ51/EPs
fX0U33uCcA0wvEVu3Lmp7xWqRNyyIbH7LxVUxV3ENZt0cRbAL8rXW386aAI+hmeHLwnKJxSbDQdv
xPPkakrj95v8HwDejPHeEQ0tc9giS+pFdqlZpckku5Zh0/QUed7iT6UPoGkYLbG1RW8P0Adt79qa
FfrceSmZpDkv3iO8aYoQxxA4LSos0fjieVJWVssNOeZiT25ifFsI8nBv+dCSt+fAKOhteU/0mNS4
Gp+eZx28QMTPh2badXhIYttqXpuESG6kF4wgD9YmF1+LYiqavJyxrCSzP1gp5qg5H9XJWpTRYn5y
QF5qyPFAG4/OZHLrG7IFkK0mZ5gZ6r3ucKO0F08vLBVX1na5kIDkKQ1rtOVr9blYyxIIB7LYjv+z
uSsIdMFm3vkPB+TiULIbl94gNuZJaaBiofAQVIW5oFTJcUPXkcQGIHgNZDUrUR0ISYXgGSgyZVZf
iudMn3QYOpb9lKanBdCA5QqUw7Q7s0wnSyiXIs4tZg05kHr1l85CkLRsEqS2+pBS8XuW3Hu5iXhW
/7DxTBY3pqTXA/mNpB9hz6+wjPIHGj/lceOHJV312gmH0L6HJXL/yrq52choaeRf6539m228zfn+
uy9n7jDf1zh0ztt//H5dyw3UVv0GZCXxlQC3VZzJgWjblaoyzerBvpJBwAlS3jp6yWlznAju4GZE
vkKnrPVvrZZpW3ZwlQDHq1+tDHfJPhBT3ldgBToxbGIicjzPDgGljD8nX32Aa6GK75h473vyHhGD
8h/V74Ossq1ERaWQCphOoDS+dM/HcchgXfvhig8lOjDM2/IffOCR8cpk9bh4voR8mtpB+2pAy3sq
Up6rH2g8pWBnsuUr+QnIpqhpMlcVmxKOmeVnVcH/tmE1CEPTKhRszmVie+hgC+4zSrGrFehgaDBC
i8h61hhJJQpyOlYMBGvOCuEAyz+XROXdL2Iuj7wA/deAoIA/vrIAdFHw1LkU3VMrkU8vkKQBEov4
Lh9iSkezJVSIZmr+9mvxZCinp7ctmc8O5CqAW7Q2sa6KYuI22YdgNzRDwV5QrtmX4WuYNaZiOeAg
0S6coYAGGtt5dthwfgxVN0pbO7jeXIG1tqQs/luLtsmS3IH7rglcZsSJ1xkhk9mEE4EbT8GVduiv
Z9FTuzTSK7KG2FOz2+3Nb6KIylDaEsLUDevKwGiNeFTrEmGZrNwPaW3Bch0Ha9WaRdxA5uSa25CR
dFp0SwUQSYtVywo1lqbnHvfsbMTSPTX7g6JcWlS2m8oh5hV3Sf61hS6r2Xc7lf5SfE4cqVxXgljW
aiNfEk6sPvbcTf+MyVFkknVmg0y4AHcTWAjVn/0LLAM9lxoH2+UokEzVrNXCp/U2T0jYyIwJk8Q6
Sgb65HgBVVxqFmnhZCUoF6xPZMdsW2EuL6MWYGx0CwELcDII0l5guhYX9DtnbTZOCxagLTpRnUsw
KrPvo4gVVS86drs4dvN6sFwEwmoHovyS71S6Z4nzaz8LDlm7D30w0Ouhgpqbc5zb5z6reLGD4uQK
yCLC1h7UjOZR6SiscSPXse2Kex7SUZfEwlJ0JIl3oNUF85zqZW1bJzYi7KL7yuV99RhxzDrkfUBe
rlo7uZBuIsmBgdauY3QqkmrdMirKhS5QHtwNYE7c0GJoP7s3f0rKEcP9rokpLw1Atga+COOlcrOC
tnbuxi4Z6ygkMokLbIeFG4HkvltUjNzmzcic1NrMFqb9snWyShqW9NpGZpMectSawN25+7nby016
CG2al87glqWCNezwGazXj0y5eiYzlEpXzvSCQqIjqt0UVkOmccPJ+vNYfrD+21XXeeLL9rnIyrNE
C/5fNyt2PKbIAVkM+yLoRktByDbWf1KxBGjFeHJcLnZ3ulF4rdnxrj46xua4nLyfhhO+E1qihirH
WPAskrdmqPD9yewhY3VZyY8lsZGpAZXyELBWe76LJxYDNz608jsl0Zglg1U8FE3elv+5OCO1UchC
A4ZIkA2EcHkUh7BKociziEkDscLYuHAPxFKTFjy+lVPAaAJMTDOlL5fT7FDcFbTLoblh8n8XaARt
xq9NlvKSn/1ssY8yFzI61wlLLSPekAkgNQSIfZXK1FL2qwgDWhPZtY8dn1pYd5DzNbNx+s1aF+81
MV39u4V16u+JU2C78o63OkymqX0kNru6pqO/VgAOhdsoIO0U2JZywf6CrpNUy8hMc1SzcbykSI/w
ZHbHvKJnE0FNdjL/kUOamqYO0Vbnc3dbR59hyrgyAAgZg+glSsh9B8J6My/FVrTtd0pFGrCBF5Q8
qpJHfr2btKG+Oyx7BG9VC5I6wHFctxBfZdHNm563QsJp/SPhgX6NDc6OJiJHIrbvv+ppiRVF0oCO
GX3gr2JBRqyuGjbiAdeqjLhBHtRrmPz3q2wQihIms+cWnaljEaEw/S2diR7wJybfF47xwpY6CFcY
CJ0W+ecSHyqktFO0dGNy0gvBM9+q3NITF+6KW3uSZH0RUAJodN2Up25j6U19p2rLKUzNHWrPXi0j
GnEBA/55rzNRKavPE1cenKjrseVEEDQnDY6DrdpBkxox0rZImrZuAGkTDjcGCegx2huKW6UYhQqE
oktfIUopPzYDpxBUa5JDk3/XQJd7OoGOtuflHQu1EFRlyVcDXo2Cb04aXgqIhRO/w2E2R7zp8TZx
MaDgS/mwjA8ANM8D6c4xVMD/2Pd2XLCn//v0ShfcHA2+s2o8+NFMPEfxQmYVWEO303XJ2sxsPlTt
4RtFeewXoQKh4/90QN27n6j4xPYcfQkzDgWB9QdM/mgXUDF6bNoJRmmZoh42UQfhPLvcvw6zVm1h
9cR8aaXqHDMZrF7ENKM1cZ/xXGHbeXGUcfH80VJxCiW6LC0nOpPFRRQM5X+SGC344lohE4U0uTVZ
vzAkSPY5LNu9mct/cZD49y7FzBKKZ9ZV8dLFZrEMtdJ5Nkxdrere6+xkOAxoe/+LvYqYHJFmVZaL
kDQPn5gIfOP22Gr3evjC+8WsFGLHuMyhsvQ7yFQfgpcYvUH+ZwH5F4lxpcGvFn3MHh3CftL7gvwb
YFshs6XruT2ce78M5w6fEBVwK0gnWgFpJ2s+fb2bHwN9F7NzMdPL5cY8lIIw0QKkHCd3pT+D4liW
2hD9kuw2u1TfTg31VBYpzktmJNmnWO+IDHU3pNboBTqvtSEdwMUSY2Tt6PyBoUBbQWNqGQQhm6Vg
kTCPUfogF+OQyQotq46ymBa/kpj16Z/Mv4pXXCY4QQE1AyGlo2ksJ3d116HcAxVHbFqWJM21ajt1
mQwmL7E9n99t2vINGNMwMOOZaABFF+oK5DuKTvg2oeqHviRFW1yd75WQQZi8KihRVjc2Y+uZpN8K
pZG6HfR3b1NX6eRbBraCMOL5NtYCms98ufd6IBMvCvUtHtAW033suT9VvgAXzaFxlM+10vSrtq/x
XFZPWgoPUYgmo3wdsHYcrrAKQxRRYxyrB2rcfvfIHaYbwSPnZRsqhjHHx1znzg/K7LDkd+J4xCr+
IC+jN6ht8tW59VH3M7rCBC+IdGREG/9W/ERzQhTPHsBiMFc3wDuq4bBC9yl7XRygByE9JRNpzIpR
2ZVbpok59LtA1GGs33UcAaHhuh9doFqrn8g2TYUE9/l0/RW1gy3q2fr9Pm9x+kJlDEzxF/p/Z2I4
pop+pPHvxdi3PnD3sK89MnWM2smQ+rKsKPh4sDscc6l/yuilNAkGAcKEp5KTSmsH/ZhuTKVItXS9
h7pFKeDLiCTB2qLwZcTRc2m+6crf4TqW0HxvWg0iupjhnbU0oHn7snCQCwBvuIFmFStMEDaLN+xr
qioXW7YOQX8LY0SrSlzUOzOfNWyeC0iTM3Xl0cyd4EbK3xK/ay9mm0K0cANETSUxDBoR7BrTgOY2
15RLkdXFF+UJWI+j+72GXCHAJllp4Kh/542YI1K89eajWJrglUgaYnDL7U8aTprZfnJ0jMcO0Ejy
P4TZvkRzdkprJjnPXdQ21fxDrepzaWAWiJ/izU9hBgkUYlIh45ddFxUbkcufpuF/5F0UY/7Irqrs
6iuGlEOKrXOBgznPbnmv5MCzQJRtW5ZkTTbHYsTorKdp70dnAIPiXod3fwvZTQUF43widBRzpgoc
yaAuSdQp8Gv2VGWvgg2h+DYuLDuepqntdl6fp9DPZI/pYJ+E8q2zrOa4PoQNmH6oZVC+LIJZKeOl
Dz1q0rCiaxwP1eNmaUNb+r7DGsKm2zCrPcecNZ3fOUBRJzlMkbMdMM8VzzWUyHnU41mbDeq9j/2j
4OY8PjtlFvH2awyWUYqG+MkEuPtNCITzvFa/RMNZYXRRYX7v9TL6TENWz/iENIXJdmPCvYLSrbN7
H8Jb3KKK/ssqqJnmzEbW9KVVbUjO90LGjNY9ievSvaENZUN7rCEGcPEfFTnnpYXR7hKktUlM4FfT
MI5dMJVoZp7fd+eVRWlhe5HqXnjQz1E4MJbjfXhUEq9mqq0OCkDHV1+kwHOi3KH2rnPD/F/bwic3
A+Bh28s1rUvJ33PMo/JT11PZHg21Om1FyGYOCPe6lOdqs0T7B3n/mQ1VqehT8KdHpelonSrg7heM
1X8k/vv3EqcQ57tQFz9tqIjnQmWvO/svVL+9vKvZ8szgY6u8R/QgYvQQ4Ycm0GXtAj8pquD5juRm
9SH5dCHXycu8ojbhiRisWZW4SQaDBZhHUK+66Qdld/+NdQD9+5pQEM39RrPYwU4gj4cTq7oJyhx0
RM7e78uoCVUv/MdPC43nxs68LKw54/4fp21WE1INvBTNPdYvP/w4us4pqaH4RIpfsjLKFIhsfDul
oa5SXb7OZeJGEaM5VZnXgc7FH4Oiklh6CLCH2BvyEelIFjJL15A6jXfu1ixUQVME7sb0uLv2HoAC
KXcTqGJzmCYUvTHUt1uVEXv8GkojeyEZMBgJd5ROD6l24dubD2H3fGH5gWGFmtmrg6K3adPLaj3r
vIHQgG+yhVHsMLk69XQvRXKzF1DwN8XqZVN4hpHoj16aWfYopH5vJlkXOhh2ViFPIsZDlg2aYPoE
sImW2dJx0cltucrgI64BljBaBBdLARZ/zfdIROmihg7/xf6ECDGpuihn04rkNmjlhOEXRgWoW4S+
/Q/TiN0DOfHxFzGlxVh9MENzJJeUJv8ls2ROlRrIYXCQUzrMMScNDBza9iS7+rrtZRxsBM0YX8Yb
sBE2xGLs1UmJuQFH00Y2PHwP95zgbVZo35t/cZrRwSGiybeRpG46yYWIU4/DQhc7+uj6SfYOkkeS
ovoVHmhTRC+tZZoSafOdJjqdizceoNokNli/lCiK6gLoF3yiQoRXUj0oBEpFYSa5PhJ/ob8znZ5h
Sh0biG7jDNXNB4RLx5IA/YOeJHjJJlUPPC4Bn/2nzn0gGI1Wrlc0kI5uO3SxbyZfk2ztVjWk88r0
xCIOT9Al83RMITy6M6NESIdYoyWe1OrFIU9B8qMFcngcPhX/qq4B34KthbI+VUbtYh6Xx3FTuo5P
/l/afx8zQ972rOPOewWKeDM6wN1Wxu8nBmcIkf0EJqNSToPqvcC5B529mrYt0AwJCSJFWsS9nmpr
clpfNPDDtrnjfwAksyqDy0C8up7mdITOGj7vWPmMvaNSNUGODMqyiKfJLkv7SExudsVWV7mdKqLN
+SjHgKC1VIxIBtRjM8FHuUyMBa2Roy1zBqEvL6cDvPcOkwAxxBOIVw1erwHfM1EdRSR+ek72FLgt
T6srTDWDjnBMGAYW4Com38ed9AitV4bkXeR77o5SHuYV/z+rDTF9gpCRWChaW5rCe84Wfd0GTegS
sZvjCHNjYVdUhDT2esMb6ExeUKTaHFAlSTOwsAApaQT5DGbK5UXbN/gi2CfD/QuQ9zZroanlLvh/
hLBI/pKnHO41EG93Ds+fUz3nMG2MDFccNGI6ABxywaHHHkUe7My+7TnpyP3mcVvoTZTbpY58BGZJ
mrnuqI7xF5Nt4s6HBYu7wLUr9ovbmsi8Q8xcb5t2Vgs5SAyiPBDHJWroLcZQDfDS0QLwiePdzIyA
TVSAXfRM/RI05Ah7QYfBWuE4WeEPVeO8O8JZNFZQTldq3To62Gh/CdGalgYEvPsl9TxA6vC5sGnK
ANyFWxPB3Wyjmn6/cNJKFItwvW4pI8vZaeRgZEz1LSe1wr6lkVRu5P3F4nJvhuQ+bCENrA7VTilD
nRYyEuituLUKl84ECBTHklEX9l+gxDUfm4Va/Ob3Xrs9Qr+6g12/1C+A4OddO69phCGIUotRhomh
xmN0vPMQFRl6xiNuv8dSxelijrhZrsj8ZEj48b9J0Eg9qBSc+ONQFwB8Z5jzgbfRZwrzcoWy5eV6
JixRSKCmZ+EgT3dkGoC4lk4KPi82ePwOScP/1YHBXO3JZ5W0maETU1fBGiCHfN2NLtimQZmVP0A7
jvcveo4sKMlcxb95cw7CvHJBsXftMe6Tx/5r9tBCwCvk6Lzqr6kSMLZLQQPaRW+ch36mKG0eiKJD
h3sKRGTma84GUdBOIMK+jlNK/fSudhu/ppukwfa20my4lHue7L28MemrQUu6955l7mU7EXsJAs7g
juYCnwG728r3mi7miNEcXZku6CtKAuuZ/Q0/lrVlxG2tQ/bhqb7946e1Nwj4Icr2KS6JxL5oaQsu
NE/qIZ/Zw/FeAy/Ge06mq5ZTeG6Y7f1kEqFvrOQPZv11A86qGSb/wWdFQQrgqUiX1vINkzuRAIQf
HiTA/dlupZ2apQ8T5tnmdBcGy6pJHLLvHwMKmRSTf8Bd+7MGI+T74UDDt/v5Li4HIPElv2sf0NGG
3TsvBXFZUsgfm+Ugg5RB1LYC7kiz5JtoKoEGRJIykQ94jbLDWWcewqCxiOaYmkSMCtPUTtHNUcGB
Ihw0ng2V7DJzIZRDo1xAMsErfGX73005dl4AE0COX6cJhmJZJA73Ie51KVMLdx40xD3cSkriUJWi
a0Dhb6/S468vDabrMkTTfN3ZG/BA8mO3KYabfCvjt6iz/2bJOltTHaV+i21+wYUosjgbctN2NcR+
fQMyBk0jkM7qcddakJn3CBYSC32TvKCht1au6oy15FEz4VqNqOJABMqHMsgGuEAkr/5XP9maLowR
gQKbRM2gKOvO9B41D/6fRJiVnQzcxXR9GzNFKhEpLJhdFHmLrdYKTt+VSZdI+CAaZpOPSTMzM2eg
ZeyLI9GICQav1MyxzGI2eYn52E33w81/tSSQqoY4kelHTn/44sFJqEWO+G6h3v2a7HroZTqauq/A
Fq0Uc9XcyEuyTHnhFfRU30Jbj2Xe39LY/GYKnDeNjrGkaDYjZP0G9uOpE5JOtZPwRW5DA+G609gB
Vb3Dq5u4VOxvnMEQlZyaxQsVAsXjUCL84+/2Qr/xdzY020FJIac0LZlG8UN6X8Ov312dnWEyrDiM
DaXDuU0JO0Oa1u9qsvtocP6ccOlZuxiQLMEH5ZC5JfxjWvqTb7VT1++rtiAiGZllAt/S47wrVLTS
cldGSpZTi8JJYjWuB4rTGO4so9QU9UB9jaAIoSnbu9mJb5T6d+DH/iD1XvZZHf/JT4wfOqFt0q1Z
jttVi/WRu3Zvr+edU2IcOhheCLQkIoTOaMdyFbFBjfrGaMG79oKF/hV3weErrqrLZV9lDRrOW91C
EfL/KDS64qQMDgspCyRxXJq+1vqPmR8B9FefNETxD96WKgCvCCF34rItkCanteW0mYs1wlNnKtch
vw5JVEYp7bl2KDxLi841eJEGQndsav0/bkkwziv1w6hWVD9HWPsJLNBF55ovgzkUnt2QXFxTI6FD
izf7++QF5XszOstzDb+62kQs+ObTTL7PcZeNseBC7zwyLYsYovASPiikJVIhI2dkBRu3dXrKfR33
+9cLUwBDKREn+1CSYtPBVXGwzKt16+zSr0RoKzubefpNYMwy7xegAg+R/q9mXW1XmXnTzsiO00+m
jPNgqUItsE38MiQmYRSlLVdr0PGNW5MKiY2tDF7JDC5er+r0BKEhSJX25IWWDcLFeNN/M7ywBvS6
YUwRxQPEPE9y20cfzeuB0WW7v0m5ZU0HMm/lAd206M+sJGFPLGornesUMK/5+RszTN59FJ2OKjEy
lnetbWLz1Bo5s4sQUB+E9C9urvy+dagdwAT2rI9zUgcJAodGJ2AuCyzQosmzIsu5EaZsYWXGt84e
dKA5hJclq2wMrtZlTuBhE2dUZy8+3bbDqRiYwmnxFgbEOsm18TFqmCfIQzn7UhRvN8ig93SUtl6X
oc2saXAYFNjfCJS6t92whg/PZhNNiwbS7KZ9d/rfYP4VpvZUMOzJU6efs9QsY5l2tz+1IsUFzH4D
yMh8wylvhschYiH05Tr955yJGPVYXgp1meK/+xl/++TRZBoKzU3OucyNsquGRbzZDIZ0U7IfX43h
x6eC1uyq/MrZmbvZS7yWWcenBmBKCwmNJpJ7yQao0nRhTUKecXDazXmkew+ZbhoVY6d2g7FIPfXv
qycxyre1k82NSL8hlodgpLU5zX52nFQ8e83clbxPh+qnNv/3yAkmT9lAkHAsmme28JNH/7Lr6HpH
foLNKrjLgF5UPxD9w+sHd/yhfwUnvWKsOJkeet4pmCh8/fdHaF13imPf4SFEas6uei5B100t/L3q
WiJTDecwOlHMII+x8U836Iqx7XPpEasPeoyCaiTdeXrta4o07Gw3s08W5TCLkuSly3RfXB0gf0qz
PPdJiLGe2oZPvr37ZgA5xtdYIPVN+s8e7q/G5n/w6vjhEdjXfSYtvfTyrxFBSVH11wKiEWcZxeKP
psLYmNR9rPJmXHFx0ZJmKq5iHLh73Z7LX5N87d6oQ6Lds10p1rJwH6nu3rFQVe9k/HGzHWDHKjq3
PnpmZynxQJ596UUh0te92TxLpOk9ljGeE7voV5JKmVUKZqDxdgJIuJwicZcYBApj+LVA081B8nhc
v4hAEEdSpZh5ApCxinq8Qw49efbNoNSi5ZdePtFXU4jakAPovylnhyGAAHn0UxZFP+0USjoZlwtb
zo/N8I2UZ5EZw9MTMfetg+vHdfU5Fsl++ZYFurO6QYqDw+7u8oV3RnoJA2ow1dfSXfV4tISURaou
ysrB9FpG9iMaOKoq0vbBwRL7J98VIUBiHdlEegs+qRqqBAZq2b+F7EAdeWFfFoRFg4pLzucoEfYb
iKK8lCn7+/fl05p056fX5gOuJRf6fFn8mD1N6Tfvmvbgc6+56JT4NHCXsyyQ7pVUHwpA7hNiyAEo
A+ISOCPCSWazCAM6jwxow8OQicgBS2Y2Mk8jblXLZ1M1I2K8kyiiRTnxHDryDxJFQ02dGud/mb/k
EmKkoBuCVeinr4Y6F+baBQ/kjCJf5EO2XB6GjmDkGjKvPkAH2IKYWfcn6iRYN+DOyiRXnk6HRP+t
So+ptM9O9JnpskM/dSYBq7FoEpttnr0Hdbk17E4wejNstqiKdFtISTbfiYwxVBIe5gelOL21eYgC
IR+ZNmcoMlkFstXTKN2gAhiDxEk5yrbyXA6Iu5drsuErX+S5tUXtCeDwKOsORtF8u4iAURHQRayg
G2ix6Qu72DHnjG3kRbLCoWkEXtJW9Y5eCXmZ6dxK/sYSYi+y3dDAnOxd+0zISKQdjgFfqZFgA2Z6
remFfE0mZi9ooOCpZInFiyyWBYcLCJEl3M07MOqtVuCo1NUfbspazGLC3zHS93Ql1Ich8R3Pg+Gi
MuQE22lsQmdFio6gKiHCZ6sM9u2CbZu2hTNrw7iLdgQMnoKDOSwvfBRvj1tJH/OjQB+fnfgok6W3
4KyGYiC39OziGqFovoACj9M9Rokx/kEzZ6Y6CueynK4af4/zkUb+uTBiT6vFKxQESzpqGSAr2hT6
4/YscdXbSSpcilt2QzyuzYgvCnEVCKWQYkPBlU2EjMvzd7nqpX096LFL8et3t4ieePMqJaIUHE5K
XOwN3XLOXzNkytihxiWbJyECZmeSajHUBDdDAMrhXTmoTg3demHEDNnlSBfj76gLsTORuEGKbUAG
MaiERTmtUk3vAut6FtXVlQrar5yeGGTaaS4xDg9CSORkuPpHvNAJHe0aLMIE5UiASAvtQCaQzt0b
y/a2HKOMaKx2VmPT+rma6YMJQWC9mjb4oP51L7iORR6dF1zgvu2eI6daq+STfPAI9ODmU6ODq7aC
fRGylkTMC7WmWSxg9prCnmT9O+s19J9SREr+NT+FQOVGIv8oPrfXz7YUpr+xedcfDq/6SC0RrAe3
TjcZm2tOKpX93SI98mwNvdtLb2vwrFEgO35+CPV6+UqoWW0qLopHeY3asvJVGftWTeIgLd5sZNwj
OwISR4k40zOUO5e62Or7JR8Pv1Jz6muQa8bgqcX5qs2V2e1Okh5DBKo+PuzEkUT+w4HZCkIm6dlK
8/pbHsxGLZBjOpDQzk4HnW0n+XIT6qMhAKbOF/VEvBz30xt1omBOjPgpUsXdzNl+UIqzptBNw3Ib
VFc/QGYmIrBHsJC9JH05NiMhpfpeg9H1mtJZ3XTknl3rE5lQY62Hyib4Km3pZamWLtJ08lXbRrQN
wz8q0QUFPYbbjcOCJZwXvFHNYbreIv1NGAhXYsU+y0cC8AMFdIK/5tikuIyS0li65oPJBFKcNUlM
DOrxSP4B9bXkP9fEo/gHEl0yCNqKYMAOYccIb5ItWcwmgcV9tkipZy0at5COXMbWXJ7zYstQIxS4
45nF41BSn5VapKLyjlzHPLlVROgvfscL/yKnC28W7qI1b3/ZUZ8jSYi9TxYiU27Ke2C2U3Amr+1B
GutlsBlMPshxC91FNSn5KB5gEdB3qn9DIomULIccxVdsYvanYNHjjUTD4xK4JhinvCVspJ/gx5m+
zrcg0kFs+5DuW1ssoqQ70OHCr5NJ2aWq01CyyvYHqJUtqMUUc3xIe40t7Sxj8RLWMKEFbc1nLrTv
S/747ygXrHBwB4HqGSdh3+iaJuxSwJ5MAqUVbOytLG15PpqvZUsHoetBIudzAKg5t0oF4BM60/Ej
3NRw52EX3hyJkzjfmdewx7iLAnofn/0izX7V6wVMawifkPVUDyUzHKMldSgnWPCArxD4nrFH5myS
hWkeWHD2/Gpl8S0G4Evz6ogcTx/HjfdXA31cegQBUrZEuadmOj6MbyV49sz3X/toasVgWmQGAAmw
84unPcVwKeqc7Oh8GQH4eb0xA2ODOBx5TWd6fLeOQhWEKwawrrCqrDrjoGJooFM/UPGK025J3juL
UlmAUNhsItHIUWbK6Loxylyy4Haw3IqLGBqsy+s11+YDGiqdhudoUqQEjTHof6IKDRRjvqTChUNU
r53GmICA+JPkDKXYlVSvFkPwmUGYsZ0RRpQb0HDIeA591XHcx/7xrg9cby221Jfem0Yk0yIobfNK
d9XbwoC/2q4yr7T+xrdINZsv5ziWsNQsKoNGz4x23rOXeccdibb26ouxU1ZvmxDPfVr3AVa6X/Vu
qB5yeIZ8UJRetSF/g7rap6mCk56FvnGY7CxntWT7qUuHirtJEzDl5ns1R4TYcCj2QQsrGAYfw/tF
FSOn2Xs2bPBGETOZctDtsE3Dqa+40DJOmoyk70xCDGD7Yt76Xk1iXDJUQTjBlvvFmgbCZQOdmyMU
l1Buk7E8BlVy18OTAYEHduvS/pR4SXtUA0BRu8Qm5msvJrmRyb4e21axc3q0h/yfMIgYJQkw0Uto
NdPLCrZPnImza5tXV8jLYLjPZnYR/oWSnVDoadhhPrnzSYRnWVH5aZMtAaocPWx7cgVE+sgkf27D
pDjUgKxfKnzT/13vnd962qgTQwsWDixXFuRKanVVvQq/Q0BVffYplA7uWZtdqhaJzQZg2Ur+mCqo
vN3atXI86O8PROOKTvwduZybYcth2qgwLmrDUv/R9LUx/UV+qWS3ENE1oGfYg1mCnJ9rVf1eqbGM
jPyZpbO652Yg9zixJ+zUUuTufwihna3ag6+l3CntTIznp/wY6dRcgNBbJzdwpaEE5itykAf8eAwN
/pnsjK55gj9X8O3DRww4x/BZveCzyoJrZhSnPkVHGaZfWBkMioXF5SNS/UBHCzcJWS8p4EOMKSeK
qZSONk/FKbqui/ZFHDXpKZmweRjKqPXS6UcPopxItzBQ+VwxMiZZdc+tiUBmsYFDTxLEMnEuhaky
1YX4OUnD2YHsS/ltS3T7mFPbC3sOYt2kKjK5nA/FA03Fgw0psBXzE8rBVBSgQM4jfB/ns4GmTMe7
DEYIWWHhUszGbGf/jGsRZURWRdNmfi6ebFOPt2rNCF2mRrM7OdV6dsR+z/S0cmOLftQOTL8VvC3f
T7b4o0neY1Rw88hajH2jKajoauuEPOXdnTf9Mswho7RY7/l6k3r0hJ4IYjZOhtCK0Kb0Adcdrt/3
NhoCCeJGewXVkWfro/V+wFPAL1kOnoyoLB8IVYzn/I/4k+/18+Qr7M2m0UlvWt+OFG4Gd3AFjNZ5
KnJLuurRxGzM8Xs43P+qDS8vZMnk/4TcYFcvrgu3Mh1vsKslO16tDVMnA1h+vJYle+9NV64p5RZ0
kOxdi2fZMLvu9e8TQb72LVhdjNiDFtwId/KsKvHHzX4FHsJHzPwRDN8I8IJbLXdMM8lkdp8MUJPD
2BiDKFJigHT6dbU9CsQ2f3rGPkOWberwJyFM8E1l+GRutGX2+t5ViZbkHHJ2vKj8aB8xX5hUhkTg
8oHxoRF/2kDWQerR2MtJsiPZnp4+bKRDeGz8dHfB5jGaGVv8SAynkjg8/CZUob/X7t7BhQzciIN4
KR6fTvnTS0ibBSKnTuWrKr26cAZPh0tGg4b9wvdte7S8f4ZLniZhrT2EWT4JOwcWP8G0fZQlaHsv
rF5M8daRo3ULASPMt7aQ5yf3dcEHLzxPIiNUC1og14l5MLJrCUn+bdyKmiA8lDKYYFQouYzRJXTK
V8UCwgFtY1Djf48OCR4h06uEKCE9TQPLAXY5Vx0bJSjixBnoHNT2FxIMrC4KxnRFojZRkh0uE9OY
zlx1deO68gLeg/b9GIfbeGKNhlMbVSoMWETAz6ynMPTfCg2SFSubWxftzgAbFK5jpw9i8j9JhgMg
3Xln1NcD63MwUx0r9c3uInX40vkoZFrYOXrPeYUXdsT3Ir4N+Ttr6CsGN6rqFkcSqpb3mDxSYA38
IW9ycGtqBqbO6xLXDjZRRwkOpVbfPuk5J6ulcF5m+7qK/GaQQMyQmdN8UJqrazTE8pGS1jKdXI7j
YFTX//twSBmShbhg9pHDrP5u5KSnEwOdUQVzX7VzRZdtogdCRmprx/aOzHjkaqJraIkcfKscF/Hx
Cg9zyPAk4GvSqYZc6ACn0QfeDyVha+7HSTBc0CZ4KBNeAACm2NcQM0PLIrOYCGHYm3f9NdRC3UlS
wrN1V6Uz00UhBydwYx+I66Z7pgFrtNVvf84GkwcgI/r2IIm+RSpXGQMH4WJ7pBQuOgKkMhmcczSK
Jonr+500L93y38RDXA6dkt+vWHywHcjWz4Yg2GMQR0CFbcBpufs2FLVHmeC0XbjmdpthazdwSlOB
Lt57sNhR5wxHQaGIacsDlwjkxU8tajB76HM7O9pJaaYwhbN4LKDZw8OVYBuHOSpcsFgmqwI59PL2
7OcF5QJaRxqc5ErnYexygJ9YUIzwKgmuwP49ulgsMb9wpV6EuzTePUCXYcaE7EQ6RBdXpguTbqFs
hems0xWe3Qgj1RYWyt7jfViyymVC2bxcV7I8qgEyQ2CEr+lwYHd1QSF8MVbyUoPWKXMCCLY5usZz
GjHpKO7jU/E3xa6CN196DhYenKpD6192QyS6kNmkL8x5H6+fkfb1eZEg36YiszsoEQHxElFT5f2m
EHyJj3DjRjtpUPY4+jvkJ+noS6nMTLLZKtPBqSmBtX4QdhXVSILuzve+9MuWN8BdCkST4pPqFudY
Huy8ri7dBF/yovM3li0koEq0VR97T+siAVN3eLkUQ7QEl3DghW/+FW0/5KEFVsuQlCypcSlSx9R7
pGft2+29Le8yaWlqfH8mOLQWcxT3FDKXuiL8iw190X0rTgluEg/Xzim0BpERh2/97XbTu0Spvo0q
jaI+i2OWr7YQVw5H9jpVzkt+mqJ47v/UzxcZ00uSJjkrS8eIDqslhrFOdEg8u6nDW4Nwvef9urk2
e9yacacCBYLWRjz4pYeXMivPvP7OQ8jF2mgZyXjHsqWitAPgJluWrIprknLCGZnO6rSKl4icLoGJ
grEPhiIgKhYeBqif7bOqfDgo4y0d0ou83BGIV3t44w5siavTgXAfwZZLPLYllswi5IIAd3zqU7ES
f/BYaZL4kuuuN9X4xZS4Xh0hSKIh02EyXmzmhZAgb2Ys1/26GBcZPpSwNDz0Rh1svDMH9iRg/RQ6
PrK0rES6RmwlX4UdZVmCm2YoxwLBosgYIgT6EMSd7aC4sai+OmuXWknZbrw/BXntun9fImjsvqvg
fRDgyQxkTimPjvwRCP9SAVlwdAp1fvAOlbcbqSKdPCFEudtkCy5ZxRFmy0IM6RXKGqKbEcmcbvya
Hlvqbk2/4fuoEyDoyHoCZ7Gl9bAh7WuAtBAfyD+ZNj8KPRqQ6ElcvIaTfAAz5yAkqBGfiHUQjsab
VbQfpT6bsX9fBfqZAbPK+xRmjVtB9Uwc4gSewnxK41ki4WLgcoEh6hCEXNNLTafZ23mLfx0tEe37
ix3pN/nClHEiTFs2W23/3YYF61yKvhE9peeoV3z8F689Gp52Pl37thM5AlMBV6jUq9hkv9yeRWSF
k2+QFBksvHhAWdTHcc5iY3SsfJf5e85VTk+pTipNsZuEB7W6vfebypVDjW+eUXs9++4hJ+78fj3G
26GBPnVZO5mB+VP0BGRt1IqYccBTasdNdQ74TItD25cSh1HG1vyGB5qBoa9iiVG0Q4mVFXy/DdXR
1FV77NHCy+AG75WF9hjv0RZgRrd1amAekBthDyIFgp76sF5oj2TGsINEBW0oDjg0KS8sTUgFi0DY
nK0Vzy1XAcM+spDXNjzIAqo5NuJ0s20gaSePi+kuqnoqBK3k8IPbj0hwKYoZIaGNWPU1anqnDE1x
N8E5BQ8pabAaXQuZQHuGNzQLsGZTereE6N6OYJKv1/PENTaR2iVhOtoOuMYnZmtAZSbuBa6QVEu9
LbmB8oaiaZ+FxjQpxKTtpalJu0iD66rz5H9+QWthd3Ij0DB37RXImUu0XK/wDYUxRmwIqBSTXvlo
Cqwjkln7sG9CWeo77UyRO0oZond2jsWUe8it8dwAt5qeajtAEFG8VScdFKIRr3PVgztmGwi1A0oC
DpHoRH4+zYI/yDoIVXi7QOQpRdA8p4ZAjBPm5XnTy+g1CjaECBOykorhM3ia3VNgjb7XRCyGC+Io
aiBOEMcA60qAlz+H3d+vEVqa6BJ63LVk9YfblaHt+Q0g6zQU2V/7iPkPBUr05pbQGzRv56esFE7A
Q/OLPN1CYHI0cnubHUoBnXtrCccgTu6I67hT+4zuUCTyY3//j8gcfmfUKjt7IzQhTNgqkhDw1Q+Y
4IUwfC49Ehpd6/x/z9olIXYcCl+SWYLWgut62wkUg4jMwh3PLlGurSmXD3XOdfhWOVBG6qpFTNei
HXxWmyljOqKKBIU8RWi0vrTZb5dFCRXZ+vwrI22Z+IEDPNKGP+3G0WuovmNEZ5l6pJmAnCAFyF85
dOqm3WKl7yaRMGTt8PmYOxV/6nekTPqEJkK4rsBizTNBm/D5Skdx+L9Ea8dSQqFr6t42BmdrKVYI
93Xc6BCZupxcN3/NF3NLrP2dpPfWZbjaznCg3nfjKEgE5uMitO7kcmYu5KZPktuh8x7AHU0Xg8+3
m3hwrI0GRk5JSuqFx8ksnFXLN5zHsIB7GX3gb1PBdeZpxlVUIpTuq154+2x7X6mEBBnKB0W7FWKR
ZyoSu1zWNiXrxo02vLPU7IPIoaTMu/On5F2heDr9/zeEp2sAZv3uuCXU10shEtgzrNKwl4Qd8FuJ
qHU2S0PU4Gsj4z9WuwP+H07JADWy1+vJjkv+3SP9zvArJWFfbMKUzK4yQHsVnX9l8yz1+6xV7n7v
iWrtc70Vk43qcucJ4SXAPhwe0dgXJ5Fh2UnV9Wkh8w5WUXwy6VqEu42RBSK0VzyN6kPTFb/J8j+L
MT5VR9FWxE4EeWUWOFtUb+AOxRPMN91cISjvqtZUMitPIb1B2HhotgsMdnSUH9ZVkne2XfnQJd8Z
gnaasj7pU5Wt3Uie5L2DgOwO9UCBvbdrk3RR0jzXtXnYDY6sA+WGKE5dmjdsV3PBwL/fjgcxWlZ6
43GCQApWQtgdXoXUJsn5CQRfvlT4301Lus2hjikuTT8qfNNBxzOPeEguYym1BSmocS/m5/rmPZld
QpAnkCut7HT4rHBVQtnA7Q0fBONKp7iaZOtq1CIpZiwVN5UCwT2PjUysZ/qhZ/rLyrVtT1dsVb1i
qPZWGhZNd9l+FEZrVlQKMVykr2z8aqIWqwVnyPHlBEzcCVmyxWmQa6proeI7beMVFmlz5z8+lcpg
TIiceLVu8CmCrDagnJtDSp/JXJbZAfYz/n2UW67mDuz4ad6RJ+OsC6bME2ml1+TCE+jC6l8J72RF
M3iK+Qjhb/Vf07a/4WghFY+SYHwFpkNBqtyekpKG+IUHL7YEVbb4hjp5tCNC4k2dmcLJBjH4Urfw
F8Q16+1PVEfUFhfpwzNRvV5uTcP6DZpvvQ17VOWUCMMjbUMlzv303Rp9zdeKE3Nax78hsrwoezC7
yvl6SuMsTpQWLLyKsMow/LJ1v+rMJbZCmzryJeAmn+SJtZdYc/p9C/DqUfKevsw5Lbw7fxPpCU5/
p1oI1/uFF/EIgY6OVHqqIS0FucxwHSUZyL0iC3LQMVx10S9KKcPbODNg0rdfpANtQuVRPq+fL+F5
RKYKmZJY8yYvStJuLJEmbE6h95JDFcAfTE97oYNl2L3ovyDc8t5wpX7ISsMjHXRoAW9QajEsvUVG
l8SlvIPwL/lOjAFgBUVFtZDDGrcOIXbsrL2IzeUWbZZMi4bDWOYiJVaNMW1YiyxQZC0oXSwVzoGO
fEehQyzAdjzlSHKo3lTz6aDls8u0J/VgZI5iu6REzAJKtWuD4qwfQSU2MT1/25lnuSnoPtneOJXz
V4Cj7ysZlaLRbA0k5XlCjbwmkasbVPAY6Y7N0DNAehV6KywofT7Bnif/enHeUfzG5GAIlUQsNDA9
UX7vDlcvzG/VO+WtB3b9d6K2226MTzsnON14utL85gDFVQWFyq51AWi2/PjcMw/Gw4ylL0+JK+B1
eQ8qMgh6xbpVxJ5KT2vhG2NHQ80nFb2pQVkKhjEre2gVI+N0wi7Y9d4qRcIJkmcqdZh7AvrqYzJ4
wtI35/gVapIH34y4L6dGS2u6zwpbEZznN3gyTclrBsNQHrmpgRWCb55kTxgE+LM88k1aAZIVgUF7
g+6G58DVAOC3Rjdxu+ZhofsSLSQDw8Xj9qYXYqbk0op/7FWc95zsFrczpVTCKgStGbFj40cYPdxC
uUnZT3faH+DaMYoxUCMvkkSZZvZEbRD8O3S1j9w7WsP4ug0JxN/H4esaMNMsQl91Do4VncN9hIsR
m5IJa3xbrqpzxIbKqpou9QbtNJrC8fmsMAcfxUP+I1+2F9wyfYnmQKIhAMFEfNCgJujA4Yp6O9q0
QULbI/7tuNhOHxObKk0Z3A7ebfzjtCDPGYwfmxb83pegzNG31i9hnrLsxv2YB40mn38YqCNVZbl4
cTRdSiVzFH6H9pTs4GvM7s5nN6gZ+fCgd/nOUPlV7ZglwQfElAxsgjdtNCYLBKpE4D3iYQ7ULJbw
gNeXMkXDdJRoym+G8n0dI1CkI+OAPSQH5wjg2+CJC+sPbzByB1EP7nY5WWHbqwqaNVDghmpuF2Ac
M2v75yP9botff/K82XqK/Fwk1ae3f+7v4RzJTqoUaBa4fKgR1/xuDll3+ajARhOQNVr8uKS09Klz
XVj/VX2UBwZgq5kfgHULC4j9jcj7FGN+Zm0Zm/MLIhBkMv2Yq+lDlLyaUZDqJAfcpeRCBR3SjeHD
j966IqUdF8koIFRZOtW13qCmYfC/vknjkEr4BD/JrA5YGQJSJCkvs6SKG/fp/7WKYfaBGZNa5mh9
h8UoBYvwPYXqXyy8O4T+DuZsBxSX5Bp2b9aW8wNizH1pyR8OwAWzpi1zTChwXmoOHPSeJtygZlrI
FDlPSRO5k1UMFXVgY14wUFllh3Sw3SBXoWMXD9rtZc3g7N3FGxD+WdkWyIEF8WMlUjpDFubobXYh
lE72bfPA1PDEjsZtcfrXUfWmS6pWI90OMsfYRiY3nCCmVZs5+1Vbjs2Uxxpr0cZdBG7zgnVxhVlv
VxPM9n0Qt9d07oxx0NeW00mwzHgJt6FjA+MQ+OTqlTz0YxFDbqW1NhW4HOeZgLVDuj+sZp7sjoYb
TXUe7EJxzwIg94mlSGV6lrW8O7fc+l3+K3eF+ziYzkC7X1ATfahfm2S2xI/n4QTJnFjxIBXXFWzq
np8UiExxH3Q+iS3PNhadFp0Ed/2uDn310mvks+TKGgmIA5xaBk/yrFE6njCrZ12hAGxUsI1ypxCi
9eqMXIsAmHlybLFSWYEIaz3dOkSOSKNitl5C0XJdT5J+3swCxdlzOSHia0wBOcd261qpqyRNkqeG
JpN9CX2kpMv7ejEX0VgIGtubf3s2HyQ5/evrbB6pObYd+/js3x67F6HIc3OpBSoC0FaiXveoxjx1
qO2FT4hDeoe+2NiBTx/8Ir1Tj5oufVX2E/EujwHqXX5VyaWuNZMm48q5r6BvaZVUq+XCo5cQwLUq
0NqHPAYZE0/Jq9d8qjP9b8a+blARBzAEjvBdCVntGN31VD2KnNhxIKHX8q83UrAiYfOWnZSmQerw
38RpsqtodFKKbieqe/JIJVhweak7VSF/e/wBO3mre4+Lc+E1As0s6Gbz/FuDFLOWp3khX5IkxgkF
7mV3gVN2vhYOoxuNoR+KQiTSb/r4lItvx4e6O97pguE9iP/w13JfTrfhKbDibZma90Y136I8/0jW
m9GzviBeNgzpg7fWFP1ctctESgc8MXLJVfrZCAavE1d4I05GYWRGh9uLPC9+igqGQYo868h749L9
sx/XAAfu1EDUUIxrOcwEKpBsyUetBlIsLxLY8zpU2RIxLxzKs3+btr3NHjipfxR3E+gqsXSNsMTt
RYTW/xZGhY4F41DA4LB7RX6ZSiR3HRtCRukE6eN3z2EIXORSa0IkyFs3URfqsPAq/Twl24l8mU4A
5CL/GoDCiJbGJ4rg7iccdJeSyeURCIlDTXEg+O+YbUgf73TRRlG+2npOLhV6jl0iSCdXqGAkO9at
3QsG+KrPZ2q/mz+GuwS1a0t0mI1fzTLMk8xwvSnwQlrN+kg7Hly7F0FZyxBRYKDxNu11bASdupTQ
gYwdvzewnFX7sHOE0kqXrcztcVetHB0m1/50WqtPoBD1h5oCHjOHW2SVN+3ciHDhuq3C3SO4h3kd
1PM/XzcVx5pdAjeT6CqWtd/Y7Sk0tpwGNL1eE0wX2EQb7BLmldlSEWXNDEfJ5Kx15rncTulzdj2n
ccxyy1A76Egi1IZuSaMftRZ/DUVKCrJ9OmyBcWvyamNkZtAuEHc121cbA3XnG4pVu0vZC4UZj9QU
UlwFcNORLR/LAfvczAjPJHdH7b10WmZs001hpuq1FCRChb4d7hu5LG/TYOA1fX7NPcLLAxMW3w83
T1kw8Ox4ZyFkXDptDpSQ7TU3It02Ctp7sjKLvmBs7cY3MUQjhjjZeRWBgD5OKVqMYYU71t8zSFoV
kESSD8xlkldDoZebtAeVMf3p1AwqX2lw9VhbQBW/TthUhkPiwytGiEHOAkVlrpRnlai0Usj/Fltv
QrbDRBZOLG+me885egbfeGPCX60Dgj4MMUvJzORBKfNzLPyriVlcx1OAANrF/J11hMrGNhYUoleL
YfpyUJue6Se67vp/g+bXuNnhY0fsZmmUstTK7iACM0Q/0g9SCvRlphhM7gT2nuEV1oFjg5rg5tyn
n7hD452V+ATjK7iXnO6QRzUY4HjS/4ZiofQb7R3ZBWaO7oyYKaTGQZ7/7H4w7wLil4mAeyo7Rl9G
TeC9kQtV8WOisxF72REEDk4zvVNzS9Z28cC31KhzYJhBG2FzWjrWyEjHUjBxFC4C3n2cYA2JR8wY
3ppXFmSzT+yF4jcJmlxXzDsF53r6aVAydj9OADVDZPSwvbVBJVVuv/kGBpiyveum3hkjj1sbkzWm
h1lapJThrWSlexvnhN9vMkblUtnBUF/Cl3GKJLM1pObsLVFESqCzJuGhsO9PiJi803g+yCCEUTTB
mqrqcc6fiFHdiYQ8U1MmzMvhXqdIbDiUOEfCj76Q3CW7hQzSQ4uv/e1X229o4Ck3W8T3T+Ld3U6N
I0biOpjvehxI+vgKZTTJGxHXj7omFaIuOFecsi3tAmCKfnpGu8wohp4yjzpIbmsbTlWYQGojrPor
LdWsaRJ6zWezITyvIaiMKbzjEMeT1jkZ5HEj2CwwQncRzadfaBoa6FydpvLRLKtn3cc/gK4i+t0o
1Zrd5hUmPWlIRl1izn8b4Nkc6JCOq4L4LzYqNVKQ+fXfjiwg4ZxMNuRRGnpUbRakjPQrhmM2YLo/
PMM33RwEhWn7E0CIDb/cxfGFgatfLztfkl5b/Egao5+WSFsqNB3bcEcqcxP+AIsYyvYtBcVv3E+c
dWwR26Rr0Gh1Z30WPO4f7Fz5nCgphScBmb6jXBBQfrfVRhP0E7xCCTgbSFrscxnDAo8wjsAOBp2e
uxIE2Nf8IXj6z5TVPqPQel9A6Z2dmX6NRi7nktzml2b7NasxXgZGx0Ff9L7CrGZuA8xiYS9siF6m
bC759D27SRkPMbDUMtxbYeZtnXzh9QRZft1wP6IUu6y+uK2DvgcCLwzorep8I2ASxVRvVddczp5O
eyjf3zXaZIRBOe7SF6XDgh8AafcIZIRNwLmQfPgQnBcEhb/THh6k1rsxCpM40ntYCteCcEEOLpYm
MVW2zHPas7iZo03SGvF/JQqSutWLsMl5/X/SYD+knFiJjzB+o/byGdnxUF2aRfE+MhjB8Dnk5tsV
TJcHTYgspiAWAL7a29PxMr005mWfNdY0kfU4KJoGUsDBs8qoH3FwM+iNpMi0BUSt9QB8GbrLo5TE
vMrDwwoQrrQmqjyNxFjO8R/PhFDlxsHHVgy5lo4xmlWyncVgDATNFfkFIo+KIhUWn8so0CVcFuoI
fLtGs77LaumJn8XSs0Q1cCRKmq84D61RC33iQiru8+DwlFH4346UaU67DTJco2+B1TB4fjzuFZen
+9XlA5b5ygVg8P/aGO66eyGme1AjkyNueKMf0KFL+CH0bBWh5jxB+Gw6OLQ7ssMEoL9c+G+KJUlR
eE1B115R6qFO8kiGt46mU2ryFsY5fNvwUEhGPDSCW7GN+oqDQloR7EdKTuWrnKuenqsPokFSPs/m
eyCdY72E5uZEQUhJPWSUrX7+vsRtDVcoOFTsliCzS2Xbl4K2SRVaQEJd9ADmOFQ0Ml33k3Ubncez
uONrb8NXG1eAFhmXHK5UBFznrlm2sxsFUQIqE/tTonxiF22F647z6ZJ7t/MYg870o44Y3W7D0yk3
oiovxc1cgZ6I+vj/L9z7em6JCaOtubMXWC6P10C61Hp3NGqML382sk22KoTKZiVhe0qUFkjmUKln
XCJCkSK9XQZrBubstkyrsptPy1J9mv1rh1bTmpaC7Zzc3tPxgJPR02RhWtQ2ZsDXRuyI2J8UJZ4A
BwzXQGK4QnIOALzUTPwZdIQfiMx9RHSAW59bR8b7bj16un3C/QHi3zrHZAUnVcHDdKaJDN3mIGgE
rz8MRUx9cIxdfOeTO37JDEysXRe6mgaKaYZViMwPM9UQt1GbDWUDkT9l50ZC8KAtxivUIf+9mPBM
k6GiapADnQBIAW7KSnpjnijFAJZSHvaEd0IOMRK4qNHUCrHOHa0ZfO78TEX/nqITxZmQ78rOXvp5
Sr4IURb0+4fhyQ6ZX6N83VJ1ftOIjTy23DMMQhAFDTnmdw1K7CS5drnPW8Ti/z892NDBcEaMXW4h
wjCpt6SSim78886XT0iGZBGfhTuGwWpQvdDJbyHnAIX3CjERv02V6mmi7GL3GytMohaqM3BDfYBK
eXS/2nIP7BFbMIQz2A0bhy6vUvSEhItDHhzfo6/MqFctW3wN3I9dZ7mdzJGHIOxlaDV5VqOZ3xr4
xCb3IH40FnQgy96SufbpCaYKkKc0+yEm3GObejXG3jxQ8+GgCbdk2zB7JkTc2V36oB0zv6c1FrFR
bb4i2p6vuk+RQ/5xMHckwEKRQM4V3OmmDaNZDE+VXQ4LWI1NM7Y3fvrtZYovR5R5DI/oQO4tDPwp
/XRiakG7ekzCnw8OXWLDuUAsQlCL8ki2FTIEAp9d1DlAEzIISq7ycnYwMCVBAaAzUYyzodHCWRrQ
n0q9iNk28XOsAnjPr9PpeOX3K0CSpbTltgElep7nI1QZXqdfgjZ7B5V8yasIpswHp2xHqH42Cz9V
NAaVaM7uUw8gkabX+ZInEb9e1tpQBM5jetTfQaajsL1rig6mJn4Ifs1/mAw2hR1WPWTdsnnJtk7o
ibojFNzxhpMQKtPa0yIqODlLiUmmo6KG6H18B5wlh1Fp3wLLdJbbhuQePKQdQuWmMBBozXCHirOt
d7bPIt8l9aAYUnfcEkk17J7QSrpsuSeG2VtTWdPC4+bZoXS0hjAKl7Ay8IpdwD09SFVfiihDUHOg
uU84eDBkrF798ltTGGLMumaqjz98Aztk6yMao27YenT0iPvNyecwTOcHtgbPZmM9LKNpk+ml8bXi
cCHNwGKzvxbr+JZF0gJA6MLrmUDUW1s2BLkvDHROjQ1q2CEJ3S9tllMV1ON8gSGqwdM29p1ccPKh
HYJAHo7CFkWVh27ESiE0ovDeNm8akRrawPDFvGGhFJ8Bf66rQUo9yzwom0XxzKR0T9M2EuBhxdnI
FuUhHPIfls+WsqCQLTBoS6Ce5XvbTVBAUr0nOrYtB5+iaHtbiLqlz+9Kx8215It3DK0P6uEtSnPL
jWEI0sJp49NtzG+2a5Q9v+ncNVfCUueDk4Iw3Gpp9npn3JQZHNaE45PIR30mxQ6SZEwJ6YkG+qae
7c3lCjo4JDQpVao27ACeyMNja5qw44ou66IpGxa7q6wiyGLDGMf7VLtv74M/u566k8hwOG6wv0bT
xwYEGbnq4L8s7aYkJamxb1+j3fCabz0ZEz0V2SWBDneHCZVIx7BNYGtVEgPQAuf6Y9u2fy0nkjF8
aC2U1AmNkISSUJLA2IVdBpLDZbelYLnT8r/JDpnk3as0MUxvAORA+CFGBRqYCxWiel5QCYG/1zKu
a7aOs7KksOTy6mG+zErxWtAyxbln19r8EUHxC/2YrywNGfjBrw+khlSZIPqUexufZXVz7woTy6vQ
zs0LCK01YjyWC7gzvo9kEjb9pAdVEUR5KoHQRUkUTIdiwbLjqEBFnFn/bN9ZGhw7uucBynSYWoJE
YCH2dbdtO3WE4EpcMbT5538D3FY0O/brYpPQDGSxRUq4puHbZAJsdWCFslV0KwQ3NOYALfgeIAvZ
1GYJ8xEw/cQrio/qFFLiWE70C7JcohKYTQZ2gddECDod8ZcvoEi8vx0MeCWIFIBkoAdTfvieuVMC
eH/FgMnQFn30aADUWr5M1SFWXSyrLwfyUDdJ2/E35fe02LbwwaUKhsesFYBrCvCZEHaeDtRXysng
hoKf1QFjDKjas7k+cq8kVHPkJMtzD++BGZPTmsbD1e+67pSokmehMOMQaBEUXRVgFUiYpM4yFl2B
G3kJgUHP1xS8x+GGII2/zFlNn+zy80/ZvGGoVdv6FUOgUvqEL+QOMG+fkm/3DvADqsdJ6g/mX+Nm
JSfeL2GDgLuNyNFcLkyDUTMVcPTdFuXUMyDzNMNaFSrlAveajfbR4biRMArs16hrkCfJzb5tHWzM
2+hGSIJdSMFLPoa1l/Y5kJ64MLUt/KN1nv+0mHxTI7ZntGW4JhODxyRsvO+brrJvkqjkNw0+LHfT
oZytaU8BUEF3H86zxX+1OHPeVaiIsBApXh+yoLsZo/lghlmiCYuuDhg2CjDhfKfopionCqk/vs62
Q+VcfLksAiXSPcRCh2dN1541TBYMehhxBfte7pC5V88LKE5fyUH2CJWqYPa7JTr/dIFx1IiMoRKp
ZYGzyrRrRPBn4uLG8fORsq5Mov3qo2fsOqHnPFV5NewQV9vxFWd//imAMGGandHTcLHiWLcMSlNE
Pw1T7K7TAKNdXGwx9Tdjmm6qYwLhIs6ZBgOHnlH1imBl6pEIp6d0bcMkmqSk1GwRqQJ8H+pvU0xJ
eQIhWg2rom2tAbK0FUE791fJYj1hA0OZmgjWvfOSi6rTaXxUGUSgql1565NDT2eoICaEgnaWlFds
VA1fe7M5VsZRnJYu+j5InR8U1iBJqVhWPPkb2h14sqRiGfroe28BJXXt+3dAlA0YeW+k2nUU4B/E
Vk8N8oJI6gZi7mMREQSr7/uv10IZtO+5YlVy1aG+TdfinbjsBrNYxSkVhMo+q/o2T8c+Uj/NHnn/
WN98WKY9OMHWcU7dK6PBslS8i7yJJ1UmNqIROqRUygexzFxcdUSaNkPASrBGGj34l5fqBD6MhFd5
r6QjRojKyJZMkLmpJRnNE336wOJiQfpfs8XGUim9Qnqd39nOdQepkQPGdMmN3KeTF6/urIuVsNED
tUnH2MkdIO+INYARPtlzCGW+nkcSH9ghfEKT9VbxcubbOYrNRueFD8dXMDkxrKIf+F947G7gOY3B
dKmr9irZsqYrw0oPJczem30jbW6Zurvw4P+Bfcn2SjmDtzDzH8gxTjuHn6FOFPCiWSXgNB0lx1Cb
J7uswIru3qLK+IUFMgqNILzRLgiWWshTh2pAPP6IamIyh/d5zTYCrTwVVnio+9ASEYPCPUpDiVkN
d+pceNDvLRZy6cGlawdO8Zn8fktKxM8HOhNiTgfHAGKJ7/eYlRVcIY4OFQ8WddP0ptBIB/DewDO3
TM1t3B005quaDtzILrE6Kzf6JV/F3b0TwLGBCgMvsFuXf1fGlO6lZvelMI3ZxliiqdqyHssHsqfW
shPzuc/1cjLHnHhou4aBFguQwSgNGwHD1zyxKmbNPMPvQLyi2Xp467Vyjq2t+9tLj89GPWoOufg3
bZtJs8w9gQHuRbN7UTLdNaVkCqa3h6HU4Mobn5wXGLd9RU4QR5BKOQfT0q/Tf3cJc3CGDwtKAJaY
dxMva6iSiVr+KsxEx7UDgelZ74zjSwCf8YC+A0fYOzX1w5LAqjb07HWPdsIrPVVOX/v0nAyT5HAJ
A2cB3dOuKBqGP9EpeCz6hHF8O5gxFu0uoGRbNzjBugSChLLCuVcQ5Vdp5Ez5BAQZK2w2LVOOQIR1
8Uv/AYc+huhpaUh3J6unP5vn+P6nGw2Cx3evULrJRIjRBsR9+D2cC+IsqstZLSs6KM2y25ndfpMZ
5WEHf5OZUIwZ41HIoaFIGFIX2fp8uL+v6MPT9VDIu/df9pTyULWCz184Id4YaVdyrlt+KehWNvVm
3iEzF5cj1uookKqVWV8JNYGXcLJspvDBfi08NzThFOBiN63LHwuDTD1AgkD2/PsIG5Mr6ix4HPiD
GjETkVxjxX+DMrZ0lFw3rh807E+ipyXlwZUCVlf5IjH6JiaUBKKVvdBCueEgllafs+eIDMhYJ9J8
GFuF9jNjHcJMKJhd+vVuq/saWN8ajsv3Sh1scDPWH1WEea+WEiuWAPCVPp68eE22DzrJXdpc1UuC
a0kL2cqdyKnSeZtBz8RUvTPKFDNOYEisss+uY4XqkVz3ajseZESNSx/iEKgFI+tfMv1TydTvjdxi
P1Y63fPKoWtwuxl+lSXkCbNTWTYp+ESdH6NSeAYB9jbPns9sc8Olxo9cXCPyybxs5oHW/Pd5uT/o
Y7oENz5V+50G7RD0TkmwY6pbBqqAfhVkjrQqLMjFaBXZBFc6d6a/TzwR48sNw5BIAq9SiRyZf7Bi
YQh5GLZgWUZLwnG/504BKHsq8vBorgJFcFv4dFBdZ50CfRuadqxSqbKRxJdhqTSRVhtMpKecDLKN
gEcLP5vNVmXgwme55Y9w1KlE4NtL/JNfjUT/Dhdri27z3sCeCo3JAjOX+sBOqZQHNzGS7gnVYCZV
wR19PDb0feLZAEFABVxcKZTi8egkEERzZyp61WWsSxt55aFpJdqnTsO/B3IjFXLkaxlkC3BpyJZi
NEqUjFDNjTWZfquTsvB+KJ3B5Gf1IC2M+Ad1rEkrIWJNPI32Ek2tmREW1rlU0YfuEGuEXo36jVol
njLj7VHumAYyW/wCjYLXTe68+Eu8rA0aE51sbYlrLw9TvCazpeMCuX+5r9zWC9bhAiTOV6JFrKfl
FbVvpa27DecjOV3OcFH3cdCmx3N7NyFrUCZhjBGZbIOCYdQpU6KwzSVV+TCTqfNZprUgJR7ftns/
erKIATq5oarVx3XvswXhKwaN14xO50pHAqWXF0nzOcl1yH1oMJGrPO9FoeB4psFfZxJjQGBRDpZw
PeQJ/dCP3tYt8s3gEvifjK5J5rvLwxg1mO+mpD1w6TTlm6yLKgCz6EiVPLcHFKIBc+t6mLgxRL0X
ZZd1kZZ1n5Pjsa4bDtVbNE/vzSjDDf+mA+Ft4hGODRfK6qjMx0U40rE9Mc2xK9FfEi4VtDxRjSkW
SVI/9SjR7W4vRiFhN0zn9rdsomALoYibhxhC+fUBJBJzx1R3Xp+XKM7Gzvz9nedhe4OcT0pn4d/m
vD3mlsq9WuNvkEzfEcf2xCh04oyIfZUIni1KV6jZ4hrYLw+y3KRm7gm94xRiNKRHIoCkoP02cpiA
7XvWrwj0JU6EL+6+4nRsqOz9wMk1aETkZ+bYPfIrZ6u6HSp6ma+2E0CkDPJoh+DIAt87I6W4P7eG
uO69IY8bvrj9Il9pIxNkRfrOJS57LYIPw0Ae7VxVoin6ChsGGR+tvp9FRBsO4ghs7LSAwmLhP2tF
nHD6JMA1ehTrjRGu6igAidLktVUZwXgJbh6N62EDSjbfeG4SIYo89wENTFD5Q8UNQGjj0mTufkKV
RtF8Uyy4q0m6iy85jv4H1k5EVtJ17qzVHG7BA7fiMNTmvyec/6vOE36rFvtFRWB7whM0XmDJjFIB
jJOqxkOtpWKvzEih4/u8+WOg/x2eRsi4ooHaUluveMbniFsYg5wWbd8igE+yHErdAUWKzE26hrjg
83BrLBwvKP2/cK4hXwORYZJgis8on8IsY+ryPmFSZig2FN+NhREtWEq4PfD9Mdk/SYNeOpIfU2Vb
Bau4L3wChkQDzrtNx3oqmDytVq4CGZF6STixPTV6QQqtoim2akSaeWzAvjBQlwKWHmOBKDR4vk+x
X1ZlnFezWbXrxB2Dj7fywBSfHghATITCmY6Q08aO10EGVbzqz+qfLL7BI4gA/uHQTuRCDHvuumyS
cFBj8qEdf6tV6T+GTcUX+ZxinAGX28OLzsrxwqdtEs+BNqmBnpgLRxbecg0/jIzjgO6VJQ8KINzj
C5pjfqtiGtlSZF8zHz4QXXAyEKz9sRWRFc3Wna/IoQnrJDB6nB/eA/97QAa6NtaCRWWnbO5rorJ1
prIhefT+QyF0IK/hu9ud7dHj1bdtV638sVwBX5rP63qWdIaxYOpuZacdDv933dUOPWj5TuoTxXCd
5WCVpGWVEmcuLojbUJFUSO1IC9znZ1z+6uBtOaU46u+d0kUS/Lg+/IM4ed33NrxZrT5BKbHivGHN
82Lv6guXmvSiAsTnZl+ZtEejhIJnJzmcFyAJ5NajR7fMU9ii6+RFRRIFxskCqpFuoiSW4zUoiQkh
KWxLAAX+qCcMceCqrFQBqKTEGdDdD0JM+e07oFhDDJEKpHtn/QlDpOI8rSy7xug1w/AeFMzySlqG
nMx8TasXA56340fG1RiL0xKky5r0tj+pcsHe6KKSXo+upb22znl0yojrusH+HWoW13l0P/hvH3nF
C5AH3rfr4pa37lJrq2zx57m6RrB7SerHq2a9hR6wTfEZfwQh0FJKi5+PDCD/TB5NcBVkiilcxrwm
OfVeKy9Mc/f/4+RNRZr1IFSjeP9p/s8nODvKIXVNYOwBfTpSsdkQ5h/3niGQjFe8GUe78T+qsprx
uEc74WW6gVLLp3iItYZ1xoFs+W27DdveJ2ZxDOw7SpJMNYMl6FOKjpZVl+2ZDgOWPmbwosi4DSGJ
UCEbRbz5nzejTGdLEja/NapbAToIQThGQjquo/C5gkzkWj4dP5OBmePjTDw4VosfldefLCXqu3Fs
f0EDE0rFilxW/HPc3oB+UlBSLtHtVjIOrePi1sXi2tz2kZM8F1/MZvGYBeSneL2umyy5wExr2UI1
o609A+purxpu1JNb634znainUGJ1rmsytzM+F9QyJQ9xYiWQMbc4rt4xzKZ8/XIK3pdjms2wsa/0
PTzqbEprphgeTUyIug80JyoE2pWotsEZiXCk//jHibzMwLhbF2aPqvWYmsvGwIIAP7sHoyv4EDHE
jD6rSzm+s6Fm/iWyghF4OqXfV0xavyPH3bIUftXvf+LIQNaHxS/eZehOq8Z19sk+2Podulakf71y
3o8IGKrmUnCrzzb1nv2kVd5hIENtxm9AmxMqk4YtBTaOG5W34X3ZQiVnKbIMsIeyF/A45aPs6Q5O
sIz77Ha8Bti8Fwox3kXMN2njXE0flkt2p0MCH0ke/BPRDCPqMLgALEHSM3R2yb68i1D5y9MLBtKt
Kx8yq7gdpCkUqaJZeXtQm921UoXBlIHf7HfP9AJXMIhVsN73hpPr8LqAH/4fexpHixj6ZAlVfFbJ
4cArvJVze9jriLoY4eXCqWBRcK3wYEUn0s/PFUUBra0KGKX7nvvRrjYBWMrLAb/Y21EBkdxl3S9h
zU5h3ycmUgKc/3483y7/L9m7BjVIHjAWcmbVS/XmqSfXtV3J/MmyltMrhl1Jvzi4kIblXletg0Yj
sh1MM6Ii00xJIX6PTFSvJ/LL208eh6SaAXsxoa3EMi8i6IAntfzplPJWGGZmzFn0J7wlcBCmHg4D
hFoaegQIC7n1AmRICeeS7FGtESt73vD+jI+i1n+3ld+1VYpnx1CaNNlM+OQw1v7WfgpMxv2+rnpm
DT5x97C1yBlcpz4/2ffle+WIopogF3ci2uQlnI4j/rnaEf9dH8r5ay2hi1ENgf4oO/cQGIDUCktJ
0WuMJAQ8Eq6hNtV3uR2x18+jXtU4ODX4kV8DJzlHDeDQIr+7B7irZE/oC24doEPPb4dNuxqPv2Uz
DzcAVtdxUUpHD5Nf85NS4u5NJyL5VsHaS1JW9OUwxV/Suk5kEgAmnKnHniZOEL/aPigJtQVRjsC1
V4enrTa5SvjFA00uaUWK8g5JKx/cWebCwFAhfv2xuodCI+whWbGR5llYV9i0+TeruxJ0fycmrIG/
yLr/6ciGui/6gSjOPXx76xkW/cHhT+rHGV415XowSKvpEMmL6Kccd9CARjOhO48dZ6NZ4vWkFM5I
+qR8P7Dv1K25XVVqGSlN4+dasaFkoAXZrSeJwvmhuKBMkY4LEtOrZkoFKr3OJEkgdpG2B6e6uWH2
kK2NMWJlWCafeQfFQPPAYZzmGBu4YcJtkYrlmc5qJlrOtE/HjuG57/+YGpCp7BHTxQLcz1WixG5/
+OC2Fz8KWYlBWhItRyCM0t8i3My2IdbITrHXe+3JUcdb3y8TNYxuwMbF1+m9TjbmYjkDfxtj0oVU
449HtUe2x5nOgzAue06H/ulQJA8kZXOFowwg2qAw6SzQXHV4PxEiAjL/KPgE0g6Uc5JuCkdDsQYN
+utKxNECXMcEnah+Rp7YJ8i4w5C4ftQuMtE7dvyIggG3uVSSB2AOtFqy6bV2+WbZ030K+a3rx7C4
+R0iPGkMWQ8OC2W75ePeLczuCRp7eu+h+9pANnbWJFqgYWDjjMJc8Sps3FxCG+jWhuMlDEcGwc3e
WK98qXNzrVdhHmVAWsZ63khqjlTKMMcWUyzzOUb9WM1DW/q5UVEFqOpJrygee03vRO7bhtZ6OTea
Ukoe2jtPrY28osdF+dhL39FC1bFc9ax5J3QsbBgaRcpWg3/7TxH+ojNLwmUpbIpbm/vrKFKPQWCK
zP+vvRIGpa+6DSi9c5RhmDwtCZZZN9iLqG0CD5JVyQjf3HQpI0bExBSiMyXrE7RLaTWmkDrSoOom
j0aWZjBRzOtOA0e1r+XVcHqLs/lXLG/yTgSz4Giks34sx6WtQrjwWFEDD8RVjUMnar6wKQ9DzpO1
q3hbrshf/lDTSsDdlmcT1nnYye+OFk+z9/5uWNrwznQYAb69EvyhBMIcKwsB+rzvxNmdTiyrEdt0
vCxKKGUXQuNE8hah0XehaMhnlI3XrlC0ZN35MjXbEkmNmQtTsE8GlPy+/fxeEcT9gmU3ollg7LSQ
rlceIV7LYXF3d9Zbw7ztK6TE+vg48HYj+YB4fQa/9UWZN8UZfRfDibbBXgxF1/sEUcxcAY2qs4iL
ygAO5mwhiFsxqq4yDfPFldnH38TWh2vHrVRA1DjpF7kgbF1laAbH0PzXQpk5RR2s4kXE8k/cWklD
iGs06Ii945+DO4HY/bFkIAMiaiLl9fzWZIPyH760D8+X0tpT8c47jsOfwsQ9sCteS3KhEEwvw8Bl
e9ZNO4rAOtOTXOamsQNPG5sLtuCN0SwRMV3WSqCAqlVuKpRVD6Pb7+EI+mcVxn3s1k9PZ6ZekY8j
jvi1VUpStZXmKlSRfyKQT73OoW1ujxSqsqWqnUC9Uh27VPW9gIPkXNOwnN9YKF1nNlDHKnv8UeD0
KuPmYaoenMWuXrvqSjiSYdgRlomPt2UkSfeXOFXAyBCM0Y5oOuKBvq8iVoAUyNcNKAyiSIOo5Qul
SJWm68jb0JdxWSIVZsbHzNJXBmPYPuhNoUNyuCvaiauVA/ad/g3rquz96LMrWOnAhU4YaT/taaye
uRfCPoonCVa0/Ic2tN0WdM1pc7LjUru5PqYKAs93dJmOFN2XLUm0k4njR7MOumbjQ22N5xNPJ9At
bVIHmLH7Rr/lCkwjUVOekPRt5c1TcP0wczQEwCFkJ1gyEZBz/uDcTlBDJBlFfZF5NxTj+4I6G20r
p+4ETKoU4iAxwbIODeZeHyxEfJIKcuPtCVup8Ydt9LuIPhqsuQsDVVDuAqc2cnvPxd5mXZhgtisk
Z5FSTPIPJO7xq8udF5IjI1w/SSZIOLTqxkJtdYqjPk28DYzOIKwQnpPrbSC28cWztueELL2jR65C
36ugURczJJb1YQ7ttG7H8tOCL3NACTz83YNt21qOFx0ht89ir60Bq7EdQrruiAiCpwADJg26eoke
XUGVZBR6KEtDBOWkkFrtZdY6VfX9Nlw63gZHILqroTGbJUjUDLWI+/4TmEyboWVmph+Ip/BtO6lI
bGwAI2MIc/goSH1chQ87bKd0tx44BflRDJps2Yw7WlCuDfP8etXFf9PrmVrJ9t8c95WQV/6Ty9qE
6gcp+frdZ3fZRvfNu4IYFVqFlC9K31oUhvgnnnOa7RmY9mU46MnZxqQPcWoCieO0SKXLiEYF/7sV
pIWQt/dpgbkiER+aowWkBaNavK0GtgxDR1Rk+5PB5V+wjYIzVrXw6yW2kaNYuGeXA9aHBEdFH7gg
8eTiiAMSfzcQAQlr/wPzV5T+TFcdK+iejh1iWe0yA19QBIIW6ZG19HgAXgA9e84+nCWTdcQ/mpW2
juvowhcShrFN0VvPua6jITKzJq96SaCJ/6FvbWA3kRFLAF+bb2LrVTqyQqMFYW6Sf0lPKs1CM2cB
o2zk1WKaJ8D1C6fLDA3uTiMvDJVbpObRZbTVOXmarsV9O1TN5JHqhT8FmKcAUIt8j0vEYOoYqqWr
AowbkIVZnuNQTtNOT6w42SD/Nx8aZflQBcgTk4MQo89RL/D8hVH43f5xKCLH8J8wMaR52xBbGoh+
A72D5vZWOHNHxUD2H1fE1RqRiT8Wr0XmyGvZrzPHWsVn5ghK12Hx1Y5xRoKLZYWTmzUYel5H4I+K
jtwM8GJzietbX7A3Tw9Ps9pPfggORpo0DSNDWusvUNG1Rdn8hiPbL1GB95tV0qxPgnUe19I/t2ng
urUz4lmAvB/ck1yh1RvN4jJN/d7gvQK09Rq+5HCj98OSBhWPbKo/kgp2hjY6r6WhgF6eFEcnHE4V
7XVc0EGcvLlIOqzNmK110tjELlxwej4hGqKC3SGceS5/taIgmUbQz3XBw8/AOE5TvXzBbBA0o2ZP
v7eO0nQdkMZqA0lZmHIe9WllY86XT7WAiGmTHGciWKNZk07H0YKRcag/n/meSAMssFyt5aXDC9ZA
3gm8DyIRE7yXrwtX1goKDsC/oes3r/ELlVCdHcOIL1WErsCufMaKJOsqD9jXXCslUbt6n3oyOHnS
QaUtdS9g1xHqeq38/ohvfARb7dScpdm1+w0Rxk0HrAY6c4DnyoECqulTFZbE6HgPgB+Gkccc9z7+
toiKK15NlRXTgkF4aBcqIPCH4xEAXEu9R6cECiTng6Rq0d4fHaVRIQp4tZLxPLFjGeDWzsRWwwUs
PcCzb04eWpbep28ZAWnJrhJ7NMyYQil3hEDBi1KDeulWftdrUTeyGHeAA8JpAQ+liiDMfADYshZp
4cB+2MHXFNPvC40zlK0d7WJwdg0QRQMTwc6K6fq08jTeLKVbISzKDJ7Ck97CXNGianfaU0DQoTel
xPX51m7XmnL6bN+pcmkVumjYNAtiig5iK26JHPdzYIt9T53EchueKtnZkZALf2W0Bzai+mhGkRhH
5ACKZvr885cG/dMhobw88EYAHXoiDDa+sfL7BwALHuABgmqzXEeEQRDds3nlCYl1TwrAngmkv7ho
2Xs9HMF5rORx60Cj7WVCtdeCoiB5Cx+IfYbFn182dqqb1w6gU3YP8d2E4xhQ9SLbEgOSxbn4q4To
qduVtl92seBYZ5H/M9GGtdabRH5pSj0CA1wmgeiFQ8gREEzWMIhTfwwI9PTzZodkpcHNxR8Lmb/m
Lfj0y3b6Ev7JOBb5gVBUWS/8JM2Akb55x2p+x0jecJD1ZASpGUZ3Qdg4i0MQItSF5LxJTqaiyjWg
1Gyh7AzJaExCCUPkePRXl0JWD2XyRmBCHCC0e1QFnroqA0JnnpY4BevOpMETqdL6aZxy33OCAoYE
vhWcclcMOqwNLeSdP3mzZHKwYlrIxbe4SirsrMXoabDyc4As5CjusFF3M5QafcSYtlWjyMMmo95R
oJzXHzjiuAbdGtzvM1DpPkE5yRjsqpaBw95QGSzA5na6rMtrfMutLRbxEdhc53q14Q39MLzRmXqj
3JMiZYQD4lJumGFxHGi2HGi2/fykUq5L0fNi/6HBPQIAfFXKi4QxJZEHCETP48SLwdQ5HSa6JhCE
l1we7YCob0xa4etuC57lOJMww76TIeoLEK2BgwzjqWIeKLrThFhJluqJsuvCrrhjthTJrKRxqkkO
rvkKmUQ2sgAX4Nht2ib37IzK9ODYc/1fzor+T6QAO0uFC3Qdhk7Wl4F99rjChIgtw3W7FGwmOO3S
qBvoXsrGDCetOKrjU2d/7lWyTRcp7g4ligxEfFMT/WTFNJ/LjBm+mv33LqUBVTUyia/Wtjx9OSH8
05rQHYOefMAhVlya9RJmy13kHaCG3A0X+HL2parx4wo36r3rkEDNLE99Au5UqvMGaepjZnZ+wi4H
+TSHWnyt8qFq0bDhg+/Urr+2oHxlea8Y4ZAwwvLmCPbxE0wlvcYMTy07gxqjUtkPXQPZkkvgoKtC
jHogM13ozNYj/WoUoEbyJ8b+Ji/tgc78iyW8FnAHujZn7GPbOoa2Xjgd6KZYEjCQStyOGPra2zHh
s9Kt6Ps+0GYtscvBwQC6SgdRI4PAFayXZKbGK1JwILnxw3z3lgPVcNjMHwSa6NxlTrrf//G+8DRd
PvQU7M3o3rSljfWUN1icMJiZhcWeWlzjcFs5C0dT1udyaYAzv7BGqc9qa7WqVbqIg2cStt08tw70
ftSknXL6tbiDoaKC3IjmWH6DInUNPzFm38kxxKFLxzklzwFQrL8e3xHPEvJVijL9gdnKm0DHdDCS
YhejgoR1L3gBP4cbD8FF9jOa5FyLvEUX6NbEI+AY3il3N179rGAg8fzMkiCCNtwUBc4Tndl7R17z
2b7KMa8KDS8Dl+FA7jJO+PGyh88d+N5s3Cgr/lRbEBDVHkYrCeUXuVo+p/rt3eMb8nHqEsEpgsk7
lOJP3ahR5xz3TcmccyIzgNx1WWbMg9DRo5IvkzhWY5TvqwZtHFFUFOFbY3XWHM28THp4p83bJ+eC
Kp60wz+fk+FKh2CsKlCkggJxnLKuGB+CmwyobXogn9t9wcUHbc4DnDx1+VkQ5XZIOp6BW0MBQ/YB
sGGJsl1pcHNVn1psBszcqqp8dElqXPT+bEpvlofDl5/yEdxL7YYtUPZ1t4TxW5cYr1TA25BEYAPk
f0AFkDqD4OV/PV9Z3rJQqQexjrW4smnfUQ4HzMcdhILChVatX5cvDx9DwOZ9QGsR1SkF2nJrrggr
DHI1AA6RwgF+t0mEr+H58N6og/QuKECTO2BcshpJRLGEsI273PIUtnTzBhKj1R805D/vdFgx9eXB
nrr9hTvWnPeYyUiGAAyEbC4NlELJx48iZDBB8LQFmzdQxXrc7rWd69MKkIK81k1C3L9D+21ImY4a
0+fO7iCdbc6Jt4OLF29Ysvkx2vz4t9rgvuu5xQb0QeSBNUxarDRzUrOvqvwVL8OkCQdfebNe50S3
1BfctrovNYYIfcwzz1+VEkYMMWcdg6wZ3OI/02l78X9Pu9MI/50Byen5bYLCXpHJ9aEhwvU6t3fx
iGKA4M6cBmsiAs3aa2S/NvOmS+mIVABR6saeqkUBdWXb3AQOjdrEbsAZiG1DLHtY+zCJykVWw/Pe
L8lc94ZlgBXBnrQJzD8mtDHYAoI9wBYidoBbG2ynV4baLvtBcJH+V4Z9HiTed9OSHSwqtb3CO2GT
K3ep+43FwJDO2WGk6nZFOUGpIlX6it+4rz/ThAXRGob3x4+D6p2cF/dqu7WjeE02CRttpEJslVun
vMDEXjPGirmjJWm+7XRl0/wukS6sHn85tMi7EFY1AzgcKCXZeDnHvAq6Rm1YKyLDpgzsGbx65fej
alr97677oGD47wKCk5rxFbv4gB9sxW7FUZ2wN5HjW7BUB/Ff9oQhH22dhPKhfnB7i3qvyePNd00e
3GZIO7ebrPyywYqUeHWSBgUT1QTP/du0rd+sP6vYbV5eo1YspvNSFzXh9qdH7Qlf9VAkr4olVf4V
zLKJdjRBhg+aa9jy7iTCX/t/JMIenjMefqhalvqyu5hT7HO2enwIhA36ZYqFwNrw9ZxklbZ/BafJ
LJTUV2wJ+hS5UFKbNHrNAHWiw5YfUXK0XaxV9Wi0i2qzPHf9bkT3yed/XgR3GBU6XA0Yz0rEKYVn
a7zHbnCjEEJhO+2MonesVkIaizUQJN0JS2ZrDMZe6ZVcrm3ZfgxGI1TfJj9UaCOk225mDqrnpZcp
RyaQ6C3fGKymYcw1BZGXj+Jn9nI0eRIR8sfkhLPKQCB5FEoIXrK33zUbGbUcNsnU5dHyDQaUFQtD
N7X+0EsoyD7gRhZwR3w+kRyxzSHUJg3MOUaJy9pQtltyxknHjj5Db8654uI/BhniXRiMbTddTarY
GfpKOTo/E55F8BTKsFt2AGAciaMrP758XQJ8m6RWg2Ci18yZOz//uw6EKtKw/IdSDSM+8/sp63s2
ZTwzJqoGUozu4tdYXVhtIaZhq3ylzmYRoq16kSgOiiejLeAUmlpqZSfKHpfmcAIMMGOCRbm3jvAg
SI4bvfpobihiUXwxbB4LWDWfNTRhjWkyjX8LofLUCndsQJ8iUg45pq1u4wHaULidiMSAqzXl1Oet
9tQA2XHRU/8zF+OdB3o5UH+YEO2tejY2S4qzjT/oXB+Veo2E1otBMbvqpiWwflYeyazBqGVyXDgR
/+ewhmJBTosJ/N48FJlDX40j2kdZUdGlgGHiwVSCAOLP1k+0VpbcQtczrB186rdB+s62hDJVp/qX
NTIOM7rAMK/ugrfUkjJxeMQLOBwjdwVQoVNjhABvJ9Xn6Ngv0wTR8VvqeBCsIEGSk7lzTm2sxGma
PJCtBFGV2L/u5vDVVRcJ5Qwu1/tuvQIYfOABA15e78iI4AxkAEYiEUbWHqvYMsz/hkqq61iRkJOT
0xWZZL5r/EqF2HVE/Digh6QQ2eM7dFZE29JSGsvClNVHjtrha/xsq68c1T5OWw9uksHiesN0GIks
pkHgKcLjhpSXqCnYoqt5XI007dUoZqILOUUKWhjPAZVfeI2Rdr8pWusmzlfdw2WvgjIKcPtAACGD
tQz+ZXjx5JyJ2ldF03E74ol8t6QExb4nlGH5sP5uVdkd3QEEgCyb6Pw14zIlYqqCwHcApM6ZX/+h
GLSsowsqD4hSjpECk+0P1c86u4C104sTdxKmP3n7Tuu3Lr+DTlhGMpVhMnL3L9pqdyFh8iWHOXXP
SBDSDmjlK7OZ26ArT+Q70XYKRIbgtjyAmPbv7tJtpd5VHk9N0sa+M17VKFKe4wviThFDcx3GqYur
nvyGega3kOjbIvrWPqhOiIcFfYRwmSGv9hqPaP4NptXFZ7dqbn+FrHSOuJUSkx2Vhr/Sdv/0O3ox
/C/2kjanYxsglkEII8jfuZqY8ACoikFRto1U+MOGnOkY2mvkF7phfLsKsyrAYyK2gbwOmp4LWEZR
3Y91BhZeTVyDmz5HWmO2Xb9icPgmQB5UYvHg5XKKtzaS7CQlqhQTgTxA5ntc0k6xFqJAnkDdtwJL
ikbOZHUwUac19vI8MCrCO2Cuh/jC+gBiCDKE/sCR9RBSQe2Jq9n6bMhtjKg370n/Q+m0inMvFyck
5Nfuf8iWES6Oyy5jZ5YY/Rus3DA/Vec6qzEtHETSnszXdLdIvDZT2xPnPmdwMeDhojtCOWjZQIHf
K3LwGN4OQFDTYpwrSiGlKkIcnMsc+QzRSwV6HSldTziNbmIhkGz4DwSpxwOkYVX0C2LVxISp0zuO
My5cZMynOTAUPtSchwLbxmogkE3JVEuSoSajn8vWfUgeulOYsRUe6o0akNa8XF1xZ6HigTtPZqlM
LHc9b6lxifPydRWkDbf3xCHlJX6LsKlHfQmewOjial25B+Ks3d4mPjnpvPvAYG6oeYGkV1yNqjMR
dZS2MdSrRdf2YZrEl0/N4kCt1BUrJbHL5XIPe9OQPbQNFRFJyf0CaHMGkbjGjcv9v77sgLB05uj2
qsh48EUGluajPd1vDDZfTafRTueWvpN8lRjU4rA+Q2ijDnFPLcnrjo2EoupDAL1MA2nj1OZPIEFE
CaRNXlNBcPeWH6zvLTo5Mysj1htOcJka6rQ1Nx3xZhAl3qIOhYe0/hSfsI39XD2avNuUzsDkKjRk
2b9ODzKOZN9kgWhDKKr1CT4KRQ0dMUbgmDZO0QSh1c+CtADwwS4kd6jPUwPyjZA+AU4dBrquPnR6
SfyK8S9xBPydDKiJhodIX/9G6JNsVZUWF942f6xKgHD1OaM9OWOi2jE/WnevkHpvIrbOYVQQoaIp
IacCWMTGXgSbf04S5ccKVKqQYE2x0zNZOrOCTH2GHBoMWMaCYrBg3pegZWBKJjXA1B5ax4vUvQ4w
3lV1F5gtUCp/6zTBKpFGltoam/9vOU0IWETzrXv2pa0LVQu5isDrya5msN5qe+X6V1d+HZxybCrw
PhFIkfz3bj+r2Sv/0mCffT+FL+o8nxKgfVymVnu1vC73yy7WBKhibxUJ4zTXYOiQ1FpR4V/I65lr
vheB61e9AfKnFj6GXX2prNVP2/kjM2D4nznq5xY4PcO2v4IAokoojzy4OqfS2qkASEoV+xiESzgS
rKUNmBzgqUi/sn/NRjGH5xvHUGXI2+t86NIehRcovM/VseqOlVxTEm7kbmpLMQ4gbrPtlWGqDrf4
/QRfhKtl7iOCa/R3OmGM/ooNVSClC3sWOtDneh4qf+8TKaa63qmMQwCz502eOiAw3SzNASpnI3nG
VKvvDX0I5UaubUCLO67sMg/FR3QnZLptUv7wp/99nJQtpo0J+LHgBF1T5iF0TkAoUdXCyGq7OawW
xagU4dI45QCqwea3l/GtzIoNy2OqdDOXk+MAfLlaunQDQ0uGWfj8Het81g7JOq+xI9wpK/XWShOj
IbYycJqS3bpNSaG3nZGiXLVZYipNLKkCYhmCnN5T+9lEByxdA+RVDaqy1to0NBce+in+BRKXyD+8
yRtXed2qcS9TEZXtqT4RqsAiAsBSFhNmbeSRlQYhdfL8gncx6bxbOYkbaNMvJerV6PePtFb91R+G
jKSDa3ik6y4bsW/7mM4tmQPazZP38YDi+zjX2y6h4gx83BpE5t8hixR/A2lmB596+oJSwjJjeVvY
YlgrJR/PCh5m9dQX4jHLIsN+VMmYbThcOgZtZkSyQ18CgZEzuXLvtQFjQl2N4rj24KhX9HhAwcwo
4VPemp84BzzU/T+T2ArOQiKOBpkXneZWqlcAjCu/w7jAgyNP9IgLDI8A7WUM+Jgursm628GP/kLg
IABDxb4XK07s/LxzekvFektm3r64ECHmeToy8Mq/qaFwFBa8lbseKkhkS+OHHZh33pIvVImIKz/d
dDw2MXFE/5tXoPLv7sBgmQ0nrlIWOxEJQHnsrVC9kkrZduWWUyMcl4DCjxwI0kAkzxwIQ4ndsMyL
M/v5JQyln+iLQqWc/xLM9UezQ8Nl6HOXpTHyW937J4egqRtmQZ0SHX+xiR/FgTJoDRGevX6H9rbu
UJrawo/FPvWRFelJ5qsbeC5B5tGg64ozp8E89FbzAXHV0YHUrP3jP+ZliYM34qPwvx1n0Rva3TH0
Ch1mznmbfAiU6kPZ/8JMY64A89vv51ift9NGLiK9UgWTI+c1QMhI2/PbdkIj606w1c46DIyu4ycy
LgtNeq02nul2smnl5U8pmRZ+IK7Nrgdk5/8pSlmlYVA3Z4SIkUKTC90Tq2arDKFk62+NnT6s8bN3
3uED3J+knGa+iNWSwRIRSDo5S3psFS3TTLIXL46Vih32xeI7kOpeojmVsrCyVDSMsFLhk5loN26z
qqMuNihhLLBhxzMu1gdfckRXFHe5UaGIRe1BuazZuuNdP89jDPB2wI+JhAKeESW4b701bHeLpSss
IjDOk2fQ3uATmQDV4PhE0JIXh2TrhFHlRmcNrSMofHUXkE17wFLTJJITHPcBdSsZ1C/UxVj5SKZc
q9l5d1MIvjvi84/9URXCPAzhOahEKS64FuQWpI673foyszGTKtM9zG5vyksPwHdB8SKkHRNDOd+k
43HefDLtsOGBsqvto0u4JT6N77S2PJyxdM19aW7OomjwIZcefRt4Yvs20BXOnVe/aW/sO5Cm7w/W
JG6pNpUjCXuaVvGmfatDP/S9TE+Njy/GvrGi8MEJD9weUnaUEytfHV5jIseA9BRHpsaWG6IxxTu2
UKc9ZoaPLCQ+CftiTLT+QOUiaBnIeXzDKHhi2BmnjElnN2hvt64t/3o4xSEAPONTV85ZpzO7VMhl
sDHyrLgPpdSiaYUdEnUZ8UTBLsVU9p/ckP+HTDpnPYuHb1fFcE394/eWHoadtur+X2KkFa3NGiEE
pyjzuXbNOYtWiYOYOpsqDeGkp6PG3mtzmHfJSOTM7kQ6k0pEX9IMB77uE6U25fx63SabxtYOS0xP
ZVwrv71ClJ6SP71nj9QZUTPDOPV4rxlFzXc2bDzaLWbWWMXV1SWMfYRNvT0WaktNntTEoW3y1RM8
dN+Bqdqc4jm3Y7WxCLG+NmF0n5WpOmNyNFTYRJX46Lqrojdr5G42pP3jyn0eilieF9xbmYWvXZmD
TY60iqj0H9Q0wYsSbWnzn7RxweT4XBFW1j2LE6xrpRVdlL/0mu9n2EhAVItTtC4rPOOhvJzgcBiO
j5eMSkjegPOOnBxTpi0kvCqjFDi0hN0zUaaGLMEy8BQqXWnO9+mJG+SXjw++Ma4cvR1R7h6MFtnB
MU6R4IXoOo+kehvxvi2qSDkxuNskp/wqGzf33Q2+Pw/Y1PJZq/curhwtL9HC9YLveapDlfJlkF4X
mBf8RfT2XcRLsLgPWSeyPpgKTEI3C25s8RNbtz4wyRF1G7GRUpk29ZITlMSbCgZYBmb0DGl4UIRM
hM9cmF7lvVcWjXPDVlHEj+rIHkk0WDSQEUq04QDX619lFo/djek73H7ttafxBTksDGf6gDMIdWW0
q/xQTCCiWKwukzIA+x1EHYl72/3v9ezTNPqNeEbGxJURmHgz4j43hdrpQyzRl243GQGcWYpAujOT
4ffg3B9SZ+XpPQ5tmWql9zCQtEe4Sx9pxm5JNHWV7/hTpzZNuofNPlR+JdbBEj8z41gZqFs3NnYy
DoFjP+upKze4aJBYGgsarIU6L+W9dWT61KwHOruPp/efXMGxbLrDlOmf8Y9+c7rrNw3wxCCi3eaL
OEIqhM9z6El2MrryZyBUdjCqbg+L/EDNENmsYlYQfus5i2X//d68F/217j1xCEW3etwBOTSWeDGD
qbGt1LUjS37jbj2O0YahJclm6bJy9zYPn5RNqH2BxZa+d+EMiQjBcRlnQXyY1wyIY8BzIoi9EyB6
Q0Sp8bTCjAKz8QYC2fBkfd5AgoCl9tsoecc168lbnfkAID9JNIDQNNYGmg8mQXU+wvblDjWs5w0P
k47XkGtthzdnHMTfzTFFuXBkFHXDiSXvdWRkoX3GTPO3keOYsYrcr7lDkUlUXoOO6EfFjtyLpw/l
LIqb6CVr1QmeYjHfdCxb7BGYtSxQvUFl3UfikLoI/McLfPTGPUe3Wp32JUCG4T3FJEb+gzORgi3u
8q5ShtgBQ1kgHKdWe9XNPSnfbwNCqtegty0zTNHwLrKEqZk86qilfDwwMwkSGWWQu89BJygaU20B
qDHwjuZe8ToiUswTbGUQWFiAzwgU7SWRYSQLXCmBzhFBEiO5H7a1piBosBSJXEry121Dh0rmpmOV
S5qlIOB7iEDX/gfdRxqH5s8s1F9gr+PrST6xoNn2Je8CUPL7JJ7KIAl3GUOI6FJ4poSfl6WyUCih
yDtzHRmUPx0DEj1ORvBDh5ATJ4wC/f09oqc553R//fPkpvpdvlU7VrwNFsf/VbrXxZiGYdDBFe9I
jhec5/hQFCRg/jK36kl6tKq4nlS3u6w2chw7ugSS+NGqNuMtM0UJphfj3vDrW4z+LVkdPWD2lsI2
nWOry3KlCiQ3pCYLGdlCA8aNJDF+Q4Io9+Ve4VuH9moayqbFVff2Ez2AOnPB2zRCPlZEAkNwXtq1
WZoTbjLgOHCC6+FJ7BWAOg/do+wPB6Up+cV6O0fWxpR5ItniAQHLl0NmIJZL/fNUIFwyjBde8fdf
msn1sFnRXR8Q6XxM3vBI0avUCyRS6cnRNe2Ega3bGoR58mhNtwWTYrfnWgBXhpzPt3lpJaaJlB5X
7g91AJpScjGWAoh9mq/OeHyNnU+nRm513J808Lva+ndiTwHYDgcdNBMSIi6Inmad2Q7Rxe9H6qcQ
JLDhXOaCwXNUNV8xjJTptPOOmkFmivofS7tMlwhDiFrfCnWQZSuXA5IBgg3vdIMMt665RowTYdSp
RBwnA3gX/FVNF6qmp7k/y/vyxK+E3sLEUJkw0KsFR+0hdQODtBeZ05d4KmkARJ7YgQ4MELOCzMle
HmnaG29EvtJy3m7IptQgGB8393Fte6vRduQFTv7gaYZrRq7F96itCv8SUCx+NXXsLQayEt9M1S2c
PoAr2C7wqvEdXxfh67cyHVZMOFPjxFO7phzmPraX2S+l0+kSfFda5S+gE0gMuEc/tt560sm3YwqO
ILGQ5Hzzc8JSNIbn7R619aZcbxoVgy6ij3B5zGLCc3kBZoXDxtTNmoIp/F/hlrv4um87h3xPIO76
Z94iiVvQashamfGTbyLEGH+FJIbDJ27V2dPUiBPeYqBNNfDOF39g4VCW4nA/Vqf51kglDzTcmVcr
gD/GWJUBKlRKjA2fIDnaV6oiQc7UCXVSZa+N4DBqCxOh0zPPLbvqIeO8phzft4ow9XJrANaLl+kT
HzXhJVZreqersBvX/tudZA17LGhiKdKMGsL1d3bueQ0VnDYHvJJhJOoBq7nG5BV2seoRJ4fvuk55
P9/QJkjtlUoP4Li1NQa0ANKftTtVoaNbceTWR8GFzEfNnW8WS5FkyPEcMRK7xJMEdkd2ma9jaxAo
w3E37QsLCtzv1GnoMeOsOq0LRGS8sVYJEICWpetRXTGSv9lEuMYl1jXVGOT+JFLDbYXnSl2lqAYR
O8769ZGTbGIxiX0ZnoK3XnpevFbPyUZxV/G2jd8LBqTcxHIW7sCQtzSn/pmiQhHjooBBHflgzpCv
EXARttLh3zAn0xp1lfb6hVIwgi/h5ExvVbCjEsKRkoldl3EDnQSwXkjgix8DEPDh0SdID3YzZ/Av
AZe1xIB1sw0r+QIPjY5Pt5ceWmaduqTiCboLnkd6FGbf09bOaWxkfnj6apOJeX/zQG5SNMX9aD4T
iZiK4dVReKUzNdEauPia4eyqUWJa7sdUIdgdDX4paydJ7ApwU5BgU9iMZtBqHXx3DthXh7N2e6bt
yVTKfCgoUtXn3d5bow9WODLGJtqjaBKR19Y9foZ+zAf1cwuoGmzu6qVd4/VVBdhfTNiecnSg2jZK
6aWvGmqB2333AA0S5WKorJNZMiBut+AFnIaBGc3dgqypjW/3LBJA4lNq7a7jclP8zjA+VTyA96W2
WzxJ1GEgeqFpOaB+i6xgKltQ8DfWPeKTOleGB+e0O+SN4hQ+xjRnhDN3BQuSIvAYFVmGZG5pdO29
slspe7/AHj4O1NLfdWAWymaBtJu88gttD9ziTobUrfdNYEASOKIpPDVX/SwXV2WfjiZu/LKi5//T
UNZTIqE/ROgYWd4t6OINtLpB6VJ5yDIKqbPBOLrybT4pnmDZCqhXrOnnSCx2lqXTkuso//esfC7f
FAq7T2a1YRCWiRAKAtzM6X67aXLFoOs33F/zGUILDGAtu2qTpdBS9ceXDxSeIXDTGCG09SWbf3f4
vmQ2TgY/q11AGhbm3TWHC8t3yoQk/rce2g21hBW7FP78CbD8kklRM01XXEwEvJiS7tyP6oHkoiNN
RZFi+zOQ3Ekivx/0mlgJSJ6+BLYNM4HAzctYj0jGR4v4mt05V/+ihlQNqDCGaT39fYhN+xmeGNX+
hGvAuSvGz/key4ADqUFFhk4VeLGVt283zudAfK18KHXYx9iLdZc8uLFdQzcOQAJujjDw/92wImHS
4yec9tVvd1Dva27FdJCiTCtd/7JKVM1QobsqL57fMecjoq3aaiCdA0KTM8YIUJk/daJCaL0ewkj/
89vx4DAadgaM4nMH6pSuz7zEhCzOEeEI5fAHaTFzmRANlDSHsfjdZe6WZXN96M7dpni3W0Zj8Zof
ZFqHGLyfiW2cQBSVW4ZjBbVHEkTKQ/dt9uGlvDj5rtvPLovH+f9mGyEppxSqEZi0dN1nTiP/LP0d
9pPus2AuB/1IbgkUW22Grtj74Qab9cp/rPxQvOihPAstyxzzeRVTjavhP37X5Uw+OKTWuksYbJu3
+fiR5QGrbJpZnLx/8hci2BGG6xVZ5jt9kZ/5GS8+L50dsiPkKZXOGq/sBntP1EKyLkqIgFw0BJVy
Kf+GBl0Y1+4iEkzNckzP1a9tgrzLL7+AAStCKlEjslVk9kckNOKQYcvnVtlNcuPAoppyGw+HPUgZ
drnArQa6mmTjlfH4VyrTG0TBoJLrMxQZpJo6QWzaZNT1kR5TWd/Fs+O81FC74z5vIjrvU9XaiSh2
lkFY8wL3icYdTLYq9SMzPwnEZZGoNovT5tWPnXakL9mpu+FMl9AWShqCWcUeDeFi6HDR2hGXPaeJ
2Zs7dY+Kb8EnbJVMMfwxk3OXNh8YALvZE3HtFTOnmOfu93p7JsbN1Yw8wIhV4Fu2PFnmgmjpVB/I
rytQBlR4dhGZsuGthV4QBcW912WQ7OzsO/owO8XtfABpCzbRVq8R4du/TMPwO+9yRx10TFE3S+JM
HzJ68FKCnQRGZu4E5Ia5xm38fJeaPn+3SihOu7wno3lPNxIMvsbVScMPHd66JYDz/DnXevmR8PZM
iYG9UM0TI5s/frHbr4cNZP3vjb1lR8ji09QnyT45Z/PbkM+HQUGHQIRaLxqQC53CKxvGto4QWGFl
anPXRL7BZUInKY6Y1d0K2QYnIjPr3I097lcE8dlZIVSa+LcDHiOuiH0Yw/5LuVQ2B5klcI1m1+eR
xe55c3jKbe3qb1L4ddudCJD9sR0oKM0sDLQ36vyvRBA6YduTrpEnZwLkLd9BRHM+wxTUcFqICXTv
bX8jbLzvj1wZqSiAkmUWbmmZr3tOLrcrblfV5f1FG5VgmLGOjzvy7rLGluActZRfSwqPqstqI77l
ZivVyGpE6yllkfgQFGnIYvLn0n+MB4lIuAwOlPW6wfTrHZ1nSw4vARIOd/p9qvkspCl4B09rrN0d
+6mW2ZhnhdT+RndqpZvSNehG/ZhkGC3GDPgFB8oTQCmxgRfHDvNmA4hCUkDqJzU6X9QU0SOabXiy
8u4ZDuopj4WH1HnY0uZoUfcfNgKtjy8dxDvdy6SWcsUjxk0f1qVHArocJnxRnWb42DEAEuRNMXK1
bk8ZrqeHN2y5K0EKDYvq/96XOd8PgzmHZznWzgoV1GC7R7nonnpicTJ4F4z148U87OK9nXRabtxc
ZURUIPeOf7vMkAm4DCB6HaPBjPsU+rTDY/QPfML92uk0qA6dphY187bXr+WRDF/16kU8cnrW2FfK
hPmm/ZN6JhomNcamaKkY42j697XXG8tDruUpRDA6WCCBUHhB5YcCEov4MWCqleWJIHXb1NTA6+OW
sHMNVkzlPt7DAWUrMk3WClBnEYGBbOn/JgoOhU1uhdxHympcg6JcVy1Yw/XGY+zbRt3nyU02dTaW
H5Pa0i+ZNyNHXFEyL5/ahIAhZQXIehSjtTFduGQ74CkfEF/tPVCHas0ukIkiygj9s5iSvBjcgQav
84eQhbADQ1qTe/3Tsc4B2OKOgVOViPg2OXoWrhqKGhvdmX1TfXWJQjmT8fHOMCjg/ctCH876hsx6
AHrMJy2Etnab35rNZZFVDELWM4pckrzP4VwhbxiAINyaaRn4VbtCalLhQ46u7WcB5Db0wv6jJx5w
ttILwu24XQm+9u7QqJpX5bk88f9A33DzMqe41E1VN0H25saLK/HNbBygdaS1xbkXCI3Y8FYym9+D
0UVeTJhr1psX//SBS29Hq6VaWkmA2E3MVnf4K4IroWLISmKUjrsPereKxcJt4PZdm4ntu8eLsXkr
rYQF59xjjQZA3vOCLrZ6nNSpDEZQ06J4me3vIgjXHbMUD+RUKbry3Bf5y1CDWKxQZclGYPE9yW8O
dqB37fs3DDyJTjy+fMPNno/S8kLyeVkwjyMAHyWK9FlJaD5Q/IYKbmpb91mPlVZc78T5fWLMtxCJ
M8jrakGPoeJjGxcUfP5AEeHYf52n579oTG2ejhyTpSxHYF/Aw95k/dcbnRFVlY6ZNS+ATQLfaITY
LAlibUgiRyA0JavVKPimg3oqewFOVoaMRG3pBfYqh6b/FXJTM8RaoP1kSZrOBH6RwoMKXUXXSE78
kCTlD+yRCGuwI8a3x6Gr7FBXITx3z1Cvo5VNcg7O2zdTJXl54S4Hkebr787gppGEimVR29Q6Hwoi
2HVcOVZmlNuIMVFdJUl/2mUcyZR2St0NZYJp2M617oil09Qpuq4h+vqZAbloT/dVorAPxPPyA/ND
Dt7y9uSqZfmY4RKx64/9zSUhyTNjgNq9Q4o2FHRkYmRHV7HLH2KIp50N6IZ5j0sPBNZ5KdY24eiG
P5hzCJBsXf1iw6arZHC6mqQSw30PYsRXNsqCshn4Wj3Xku1yqZYVGprjqcHLs5Pm00xJ4o1eIGnN
m4xW+PxkiNIIdE5RzssjIzICRz1rQZAetuwM8jdqW6bVDiHF1DCX5Q3K7qcpwykApgw0wVZ9ePEM
LPlZPFWLNKHgLPk1URkmgFjDzoxuuNm/w9ukopQsUj6YloOuzjd0tHPaP5lp0i7j1tUG7uxjvJCF
JI8trX14MlkVUAgIv8ppIhyOS0xX+fSNmzyQqRm7EwY+WF17fuaL++ET19WM9RQhrFiepB5OCIIG
87pahy/e7PbFJcB8a3iQ76OiE9fPCgzwF3XXYgPBnjZDJlrF6OFEG/J2h+sNa6bl8r6/rQxnDw46
MY9SFCZC8I7KVI4U7cNxqjHdhPUJDrgoeUKMNeMywhEB974Vdrs39EhKy2enBVcu4RVTNfIRsmbS
fYgB0kf2OZLL+nNDX6iw7ZVkSWwq4E1geOaGfuIcb8XGwQaqpv6AyuHq9qVhbYTb2mEZgxwFScpP
pgJK09sXUv51gPSiHbV9EzrHRBne2zeVP1NXe4H6YRJjXXvnHAEgkWpxAN/EgaatZJlnqWI5363s
mFBmSnJkA/nlRWpFkLcODkQEoJ5edblGb5wMzwJy6PgETLROwLPENHKeJyd6G2v6b0lLBiRpFu7z
jzUj8VCdjjGdD9TncqpsV3V94d682PwJWin0TKS3Om2dXDCavOONFOrvLbnzLcE3CMJaNY96L+JF
hqdNH21VIdP6udqs2KOLUX4U5VIO/P350Lg1WVIh1bChAwEIk8CjhcfgGu25AKUMUf3E7EKRUuln
Lj0LalVdYKbrIvkBjHovYut5VpfPsQoSUTd1NajVni5t9iXU0SnyOOuswf7qE26BW1RnhlYQGZS4
siRpwtqGW1fxmf/31y65Lxa+/B5qYcLskv4omH1oyLl83I/qQNtkCyjQhwg9FX0JHOKEihwfXntM
8oUqDVcurLt4hi9TwWVCqtqtwdxXxZl++899TXxqpZpk0eschgnJPtCMosDB07XazrOpzOodJ9xn
Ve0xHmpYNXZsTcpVE0mrr40CSyglQ1hzjHjeoB+ZjpCLKtO3GkZdxekdJSRGUcC5nOVv7ZUSpBUU
kj1eOkAKIICpHp/umCBsw6lxgXwLB/k5h4PICxQ44i71FB/zuDrm63lIio1QIPCKQK51VGmWhTGC
FvZMimi7WPEm0Mv9hHoJwKNEv4hmeoj2r/Mn5kcPlcaRJglROw8DLB4P0n293Y8FUR+xBAqcni0K
XAzkMaRlhc8iRlTIMrMCWHxWMTGc6HytIFPjNqw3UUL2b+U++Ah3znI/aSRZnYBM+bsnXmGg5dWl
IuOd357PDGkVbilN0mH2ithidLtpKws50n8iajzNFMlFLDs+CAURP+Uen/khi25M3S0yJNT/GGjP
rPuT/2smlys/dwUR6n+J2RbZxOJM0LpFA3mBuDWLHjl6H4ym/F6mFZExj1wXmAsIiHu3dK7t4TuO
Bd4EmpG+jWyyFMSJbrJsgxFVIDs7lHZvsNl/x3N7/1XobU+uaaTa7P7LW6tF1ERPF1qXtJaJoEYn
i6z09wMNlQr343G4yTMI4kVOlMCn/BVZ0/SfPfi8p+SymKlbUkzkaSui1qBEwRwp6wYNwDj5c18P
DXyQFYPx64O4Y4n5ARCIQb7av6p3jnozdrtSUePIVqROh+OIaIjk0ZBxU+WvpPF6O0uDaDXDw8MP
bjNDQsPb6NHjOCvOHvThuEPTNs1AtAJzkHsrjeVBMWG20oB3ATyPTBoZZHTnw6kXDsvANVr9qx+h
u8PXy+sGRfXVUx+PpTIouorPLwTZBpYa+OJlsxRauEsixca3oVsPdiCUT76WrW1cvG148aC95yLN
KiVD3xGFc3Kme5MCA5skl+SuTJRhbb9QBXIu1v+p93OcIk+Uy8uXIQm89onj/Jdc9nK6aj/SxY9f
huteJfTtILmA4cmL9szh9vjRdptULAsFleIHvQFeFrnYv+HMcvcbFuDe+zaLb+mzl/+Rip5FGnFq
+wKbNs5wLm4Kpb06nhRw4YTD2jBAZLfp2R76i2MWfEk1grSx26whqwKUwYRYUBmQwdExgUj2qN2j
Ic0kigUdgUnmsWUPdqqW5E5V/RromjhtW/l8Ize/uNJXzt8NK/qlDoXkxA6cQAJ6xN6ZVFEV83PJ
JqyENAJLQs9T/GwVYbNn8F2+lMt728trr16++f69cZk4ON0h6hEHpDRHlc9fYWce+kqTNrCKidBw
icdQMuH3LohANwfUsmWwspRrTGPXQCkcbZ1U7XFk2EiOwhiiRJKz20TsWvQSMrqF7jfVPvYhSpnn
3ZktXm0hs6MEsjZeJmaPIAdLmh4Ainn2klsjTjx5jqZer4/uzoI/KTAd7kXY+hRtX14Wrz2Znhrs
Ci1Hy7URVfh0tKaAjmdPgF7vQNzAZTMmDzPwfJZa3ewmqXqZudrAO/oQexE6XtbY381WKkI5rcI8
vIuUwCrsGxYAzkGrq9QJIPbqPpgrJe2EdpEJJbSvZUmHIsDGQgWEb314KD6BkINWz90x7F1Z2/7Z
FGZMsnWvpGmrwfMGWCA8NwwA9rY+uGBATzkSXn3e2I6eZAoM4oQ8RdHzVpJ196uQQfo67bfYrIl3
EXEdFvv6uqBxq2rJ8gZU+llQXY/2VCEhqSFqYiJUxLUC8/3MjhfYln1balI/pMRQ6GeqxAa6WUWZ
clC7Krs7rtbknFdCN3iGCHvNFJBnj6i6cE8d0lOgprDl3JHdZW3hF8dkOTNehaStLfdL2mPyTKDc
n8STZJo68bkRRHh26WERUQxpJtum+2XLzUk14kVuUad9gakVS5Pa2RZEmPWZJoKE49ZkRHl0ByHo
B3q2vnS+uvOkch4IZ/YhdUkRDP8invy7Pnx9iLcpzgOdAbusEuPg2xhGdABhhUQv8uCto/qoYV3U
C3wFhnfZL038YkFhs2xEW8YzCThH4vGJBsQc0jCHsq9wjRAqSNYxMekglGTVy3Psw0t1rZxvvC+y
7nfWJFJwF2iPiRQIGm91V6MlUR3Hg5yrGg/c3WYyKZvfWP6jgDWOB0/tbi6j6Lu5rzIpFs7H2QH7
e3Zkon0k/nyo5jyydDhkBUworHF0/GkB6rfh75egauKmbRzsx47so8T8IkaFKfimZTrAzPiciEeF
7lVLjckPXIeK7dPeIehFXD8NiDDUaO1K8LtVroXKeUoiniDgB/AEhzD2+lQzquLSGdpjYAdI7Y4g
KyNBFdmzLBIFW8Jff30gMr1WNF4l0AB3PLtA+k2fEgGYg1qBqTxNc90kPLlFxiqlD3lBglZzDPH3
JujiYcnFnodzVPLwyF12KXJDaSlQ5r06hCXjgW7N5rLbctMy9dVSQlOdMr+tKzynEo0N2ck7mYAR
xr0Qgu40z9BKaFSshGaAXjei1JFCbX0+i2JDP9ucySuQH3YzzXqQi9BID51JV3qKoiF16hARRnfo
CPVT/VSGT2xCBQZDMffR+nQsAd3L0//aNufoXucfa//Plaz3859SkdJsdZty8xC+/5dKpeFyMpN8
mT9hdLBwjUL2ptXwOKSXxjh/x876VfIvFeXcjZMwHgp5ntlKzRsHCaPYRGKzbic25iIlQERhlF1y
QmQXah6DtcZKg/xyZixpsjHi48Um0I10I/TUVISV7hfT3mRK289pCN/HPnbrOnKRVzwmRKL9T5Fc
GzD2tAThYDcWV9fO+HitIgcvCoWVpV6I/9FdUkPaef5PpIv+KT7RyQbzKctixWAK1nA8c7al57GN
A0Jz14cbTF3ixBlgxwfgJihTh/y9xEVejP+1+L+91mQW1G2LGPv5w9km+C8tZkZXZiyabU7ZOZRt
+O5+NfVBV346VCUvKCKwifbexS1KE9zSwDJqqP9WER8Xt6Zuvl0IOGokwyXtPBIMYDd1ruvZjCV8
NphW1GL00dQHl1X0ozl1tq3QQVz+G0QrOAkA2hZuZs0nc+adiKky1UdcSMFSAIaCN83gb5T6Hfze
P0Rl0S/ZhHiL1xYmhv1qO1w0nyXaSzgDM4VdoQdlFZM5h/QAj0ETTP+sQFVTh3/3aXt5/W1pS1T5
BfvWs2+phpSXU92PqH0QSB0mKwjHV6SN/Iuv3nQTWeqi8rVJ5d7zrDy7/WsEnWc0Wr7KrDWiAOSw
rQWozANXp9H9tkK12ASbrSN7JqyiOxIGpfFASbLb8HaRugn9HrlxGvadSMFqQXre/OfV/mDzdWh6
IS7PZNx5QZrCukRgCDYfc/3lpNLF6ElzD0Z6DS4jEJjFFjARwpU0q+drtQXO9DEYyLkK8QMxIsoF
TKTwPS974ilREqXyAHXPfpz7eQ/50iRrms72s1e9oQk3yQ04Qw/sUA3ZEXxgwpVPGpUlLR5ueZ8F
JvQPf/q3kYy8vncZ6b8fV2/pzt4iNR3iaZ53sElEM52jSe9RQi0oJZ1ZX8/82NitK7nJphAvP6nz
tRYANlekP7xOCY6YGijMCQI/K2uHex8jABSggsJ+8myBj4gNFdO3w+3RpolNcmCeI78YI8xznTKd
ZzvnFcYcp0GMGf7K35H5sLmunUcIFdORX0F045kb0g6fRcLllG0zriFNTw2wydQgufrQRxfiQflv
mkBexz8JDbQKqvTYUvTS4y1bL8QV4pu3dmUZeAuKhsD9e2wOIr5spqRO+PVFhuTfqwU67RZZ5Yso
E+Dj/tDnACT61VFK8ap3GlzygQDTT7OxxD+fK9R6SuBMLH+fiqPfNDRM9btvq2Xat20r1sVGJmHX
UDcY/rbh9KxnjG5edD9gh4NUoNKWfGR3SVVH1zpEf3bNAfyar0g+MrPuSl5Hwg2Qzw0BiducLqw5
nWVspu1v1IHL5UEPzWEANNiONW06w9SXgNrftU+W/8TYle16qibyTemRWIeqmBFueFTZ7IL4uLBF
i5uV1TVcnyun5GAsvE2IpheA5nbgU8t/5h+sH+MrVCtNQaaXw2yHRoJV3dY9xofOt90a9U5mTxeI
MSRvqtLupJWC2QK3lHBJP8xwdR71JDSRGRVSN7sciCx6VM7P1iLaH2G5yVgYaI3sg1sxz5rWj3KD
9OBBDpIHdxOXTw4hrd99vFxOV+2G/eZo7tQQ3YjJWcDkdYk/ttA2huJMAKlfHqfpvp8WixQGDuTz
7JQDl7XKLJCu0xdCHcKsEQJRfwMCXBpC4V75HDeUs62yj2EwdidJuqo65Rh/LtppOSCqAXuA+vPS
tigHtctSyrmKF3wzCkUIIGtfPgzuFt5ko2NDB/aA17nM06Qc4Xqki2hJicJZ2rejlauWKT4JRlAf
FYAoG4wywMRZRDsgwM16vVzDgvwB4iMXRQL3rIVeeL1IgMTMGSF8BCRIxnlUhkFopmLmO3f1lFok
jqO9rRJUJvS+J4/ssq3Xr9m/TFSZ0DPw0JjZUD8bFCqG/qtuAMSa1IFEoiJfKv2xZcnGGizdaesi
YDpLJI+kxuMMK9NtGfOSdjJd/FCiaQ9S3ehxwX7qYY3mDZWxWwI8UDN7pEaX7+UJNzGbz8lXr0sD
8RZtamj+00YmdXo68FMojDhnUnmmDXVWY8iCIRGRHDMqUyZovQmCRWaBPPxnnKU2/7rmjOnlB2+9
IV5gOJBD8smllOIAxEe//Z+AxtVBgWfFmiXANSStVgdvAdFzaDTRrLM8zlywa+SXgJ51yMtwkFOo
xXdBaJDPmHib/N9X/SwipRT50TjppMnCfEEZ6s1tvvFn3yeE0edzbNTSY5rZhP4lsna+x/p14SDC
98rAjvidW2xBpNAjFoSz1ATAL9vG2u62p3wAy351aGm2MjhwRAdGzaCw4X/oSNqocdssdQCLwinu
kliEWLwo7AK5OsBBoC7oiaoPrRNEkKMQ4dAxrOPe4PEFAzy07o9zykzUWxkqnif1n/f7ER2z8LKK
v3RQMvZTAEYuYRMt55/LsrJhmh9vjVtUCCsHBsVe5x1K9i7I4KERLSXGEh7JX43Ntl7KPhw5QhoZ
cuj8+SfDCt62sjJF7WeRV0HrcMukP75HLI+kNmUSASNhXoSLrl2NpBvfu2K17ANkHoF3Axe3JKOC
xISVwVoqea/q/W7GAqJ1FqEQZ+RiprCBvsACvP0n0pkzq2MCjhFILadHwVH3gr6Hj87WNI/gh+e6
I5J8OzMSR7d8VAB040Ri5jguAR4y8xDpb0YqwWcUg76mTrg7FATHxZ+9yVl2TVj1lk+r6dTS0g8v
lwda9Ly3KQohfkQibIK35+S1/QGCCJKv8CRBYLDE/IsniVGsmdG8MxkaOviXbD+F3NJ+9S3TuIKV
dBi4G5rO22g1TFEPgbdzIuYiZvAagbjtzQJ5EJIEuvx4pKc0E96u+De83JG5UBmecOjgGETlT6ce
3GpHgDfQOiuutEFf3OeHxL/yXg5nmrwPBnYq/QGtbB9PqiCnPU9K1MfTGRPosOHpBCxqOOawbfMm
39ljy3fhIdoBHMT7vIHX+0WEWbzgzq1Pmy8CJ1TXZu3EeHCU2sjyx+e1PtUkzj8Z7HzRTS/TDTyf
K/rdr23j20PyTTMEVnp04A6WC725LRWq0n+KXmn5Wa3vt7dm2DWCbpEY4LLrr3z9E/Y5+Cv2KMV2
PHrg2GAjBHs/hSMM2UPz8KLydxWSkTFs71PVpFE6mtBVW/ioQqjWmbX1Sm8KMEzALycBvOOGK8ho
G6VbJ+27Rj+yvG36LIAUY5kuIHLZc3WdHdTGe6ImVhe+g18ns3wOLbM6FAY/fI3xtAlv2OdemJlm
YcbndKMsResnYe05SiRicxwDUinQnI1jhvwV8Cyj9xX420bSFDGGwRAruOjErttoWO30djtPb1Nj
VySnxNq5xLGbnN5tVFX1QRw11+OlW9Sdjdrdx7RHZ1Cm+wjz2woOMgc+UaDzf8hZD3gfRB3BHuZJ
0+uCJfPurZykxOOGetYenQGnD/lqsnU8ZgA16X8DufR3WF9ehbm1vjswZHSkLyt9k6hhOeAYBsWC
oR3cAa5Dn868GXh9lQ9b5IdySBN2fSpbfAmKyhV1nx1B2rDz99+GLW7Ps+AwA8ruKwyntuYZaTO5
N7uc/O4Os/8tOw0dcFz90SCWNWArMUCwNZnJTwWcmywVJ+yBaFxax+Q8JudaQ/wBVJV9YBdKgGK9
tkdo3eTboY8zelXlXf+s6UnHjLamf5fbVcmACtq2Pmb1qbx6wXFssyBr23G8gb1yaBusmsz5+0N5
P0UlQ4+nb62+ThFdhUtWHJ37ApDEksXUgpkDKhfGQwMHDn3Qo42dtD8uOtLcadmzXAUZMqvzKX+3
UevSApkj1QVd8WCUVgf91FscY0ZC3HF5UKc7ZAFrZqsNNy13eVn9mZvrvg6ojZx9sWakfoZIg+XY
XdqlEM1D60HGU+FIu01cZkpKBm30A4EBHnGt26fFcfbP7KHBU1NBiKFqEm3roExblpXdZsuBx6SO
v7Q9s7szo3OF2AYe00UzpvK7PzI4DF9Dod1HYPT/nyfTCaGTUNuwVdUG7p1OfKQJizubPG9RefDC
3+zeW6moZWp5D3RixU/pS1qP2HkLp7lpOfQCc5hShJxZ0DaPJYUTZ5nXt9PnPVgH9soPcOoxmnUS
/O2tjT1hbq4Sa++hOnpITVOMLQszTbLqOEbr0zhPEkQzvEK732D2I/iC5smGg0l1SYqdaqJBnjCy
XSamzuw/EyhLzbVpCYtt0KbwpDYMEt9z9r8eKm59HlcerWBGGMOdhcWD+Xtm9UfEnaVXnd5yq7j4
fMqL5hJbdgaSnexlnpdwm/9XPXp5Gz8xmhm4s1MeKPOHtZagBixolfzk2SUyNbF7d33JPv+ObNvF
cBvUp7/GEJCIZSks+/gkksDLBlsBsw7ZF+qX04dXuLwb3m5INevFOUMtxBdIUkdSWmWmGIQtM15v
vtQd+OSGFEvo3dyA/anKARVS/BUBJyRfgprgzdCj0TE+tNC83WglaFWJ9EEAiiriCzKZ93p7XCUb
VAaDvvogu8eIOTas5l2RExNeVpB2TIc1Tk5+oiT6wlJt4FZgI8keXYJYDIavsH8CP7DNnvsTGZB1
DLg5UchE6EPMsRpXXhs33DWlXfoXyYhyNnMdl3Agn/xBgBEQ6rerqxO4z3Kit2OhSuiASbw091yO
rBVOOXp2wPIR2EHsfFL1CGUVN1464LLjUCsST0V4fe5Sb15wTeihDsGGwu6dL4Ag+ZdmqRS4eFuc
QROogwWxs4ninMk0abGy2qym8ehP919ba90TINFJZRCozCSyCT6aUWCJZ2jlA9ep2ZfWNynjfr26
kxyVZlW5viyMJAvzPY9SESyXSCpeqUI8XZ1dJPbmUkGLgi7U2eaGLtar3IPWt5TTITEqwOhOVsbD
EBFVM1u1065ZtO+ZJXlVgO+ZkrTQGzlHhNI9WqbOV3x97g/YGBQKLTiEQoRNaGilD7gEjvKnAB9f
qb1ZRa+YdpF2CTYsNRySlx8Mypymouq8c5Pl7aAM1HJhanAInjwU29u+c+DxWrMn8jZpXY9fPNns
JR4g4eDBkf0HNPZmy4FdhxvX3sOnGNAzsxixRTCtgbM6HV7/mSRGi5CGSQjqER7tT+ihzIX4EQ1n
h69mUuYieYfAcUyl+gJwNxXIQNH4tT7Vwl7SQVWIKKViJ0G00AeW7wCT+6HDNDTe/riQgmw7ZQ+i
u1JnO6wjdVHvqYe2UoEuLwlyFNpOtN6B4aM3hsUUeXfK1+YWtQ74bMRH0jqQ2UaWaE78nxWO5XqW
ONyTpRWacqiKpI/Y8YYbBjERjVviZNPlDpA9j+q0X9VfmRLxsNLqlxh0Z6FOjgkoj2Oiht3wP1kG
U64V7Ylw8JRqDesLkbgS3nYQy2xFsrgsr3Nh6k4KI5pwEGa8kHNAKnUMGesLI1GzDCno/hw5Qnvw
EMjr5PMiR9vfQ7iyJJQIa/P4XfEhu44+jFr4JKpZ2kOVgHFT9XtdQkSxEYcr5jDbkG7CjGsiR15f
fI2e9syJ0KxxVGry0U6sxH19x7ICmmZGD7F263UE+ovTUohcvsVZbetrK7vpm3FYoMB0kS5+gl1n
4jTdROhQPlJs2ER4hzZCzaUdCJO1+T4V/NxodnTqLSvaL74GoN+qWtqpEmV7ZvWZkiG5EalLKNT/
cVL5klDmztH0/4tMoxfOjJg0KOB1zPbuL/I2ocLu5MDnbUTfYsoSN8uBJfInIVG50Atu3YRdt5qB
TmGEiawXa/oMb2D3hBXlLOaRRDfC7P5on7KaJVwPjAISOjwYVH/AB5Lg5vdZlsTN3GSiJA1++Kum
W56KINKgFtuawTioL3okW4B0f8SJrwFB2YF0HMtNij4SJ5UQ3ZAybCTsqjqKqnFl7ZOU28u9fxDW
nI4kmNM15AGnXuIQQAtzQ9cpS6AlHHkFzpw6AcRIvRgIPsEUHfvYs5/iaozfyVPD244QTCp8WSVZ
zPVfvO+E6Qujn7H4W/n28mOjnV2qNcErgaHzAixE0bnI0WoCVV0TeNmOyabErwQfeb/afL52N9nr
GBcRP4MoLL/8sWWs9ZfVbcS9+EU4uxDqwkJE5JsPOmA1Js22SWLbepXAL8UC+BZOpc03jWIPMdtQ
gwtm/25QLSBcNUb0W9jsM99LQFmP4w6LayYmFIwjz9Qm6vdVYofLj4ngkc7bE9eB/GOCTrXVMKNe
oubiCTre1pmCtZpSWZrx+eyLe+QgHjKlPEUki3p1CuLgefmXZnKo55wRasCLT8cjZkmvDMYiPZvC
zawiwdmodhaHrMxoTCnyvrUgJF20zuwkTTeEL+lqjyExznYGqm322VASL3oQ/C0hcfIDP+lroaRo
7aDMkboBFJFPdFbYN3uJzSti7woLECIJgATEXVLi/8TkMuVUW7Z71iajNUVB4GVS8JSoCW00uCNr
+FuLpXrzNQm107xrW4nuFC5+45m/XUPnQSjaE5W5rZycECLpT6IgzdT2u51ZSp4RWmJ+myN3ItS8
lB8H6epBlrdbilW5PPXFHLRvOsYHLI9QeTMMbJAAuIdKEfhoVuhRS5VxWEo/LcNiPCerxtZiCmNX
X6yB/vx2opkG+/1vu7jyi4D+yuQS5Z6AWGO3fQdrpZHxBaualtIbMc6x5R4btripPsLlS9OzEM3g
NfcaaZU2xJztjlNCdDFLC5pmzZQLD+3PbgvGwSDIkeS+FCYqPT6wxSjkeX11fdgTock0H6BBsv/Y
/ySOWr/fm6td28ZnEas35ybWzKPr3ij6iqrvDlOM7xUV2dj6wNW5rVBEN1dTB1FNg/GIx/zp6g0L
u9/EJZcbrFOYf82RM5sUevf4R4QCqaKucA8tKgij4q8r2SIjc/lcQYZUA5EjG9v9IoLqaIGO2ccf
xLmILdu5sJnL4eyqPcGjKbLrY/Qv05lXG5y8FEsbxBJj4loc7x641HhA0HS49LQbRnk/HfIkHo+L
QlLQJn3pyaGqLG9h6CBi4Ee4nF8oo2grSIMp3+hrqKDR48jalhxydsHYxYQfw/6EZ06VbI17rTM0
nx2slnd8Ir8OqFIIiPEK4Cin18yH/YIwri/6LE9O97n7HZj5JdP+gAHn/lIYkzqDPFEm9lGSshvQ
PHC63g2apbBvIoLwMY84/zNIYjfxkoOmYO1qtGh/s6/jeKZTTmuQY2xWoPv0k28GZnyudnNp6cbh
rzn9hTwDlXp5fiPWzUx5zR9SlvkgILc0tA8tNOlFCaq5mbVj4ut6pgMlq9Rz5CrxOizLAf23goH1
iVk8vSRpHEyQaqPRkPe3tLfLtAkM/rmqbRMkwQ8CQyFsGl3Z60ITDErfkorKIecob9BenWdhG/9C
XZnfgS61XQcPRd/HDNOSTeXsMAWHIGXTTk6c15T24dP/Py2shUAsgiOwOq879YDXdDSPkUrn7oYm
evMMcwE7PbAtIJUQmzFtrRg7NCLOvrQtQtIH6Ze2Y4uOYS4alkNblCGzrRWlRArFJ+eNivrt93xE
6so+EZ8ZEyF1+RmA2J+jYXEVQMyB29jyjJJSrdv+LO4s1zuu94OI1m5hO/YT4oozqdbPircYMoDZ
MMakG7+V9+r7JgVvoXshA2IMQrUkLU1Da1v/Ui6uS/OlWxwIYra0CW1QcpobLgwp2fRYUTdFQKGT
a2ol8vcSAem+pzB6qXA1T6XhUVVK+ZZDt5GtFsdUpbMfgYJlwsTTGEL+48vRiLNbQ0l1LjPGS1fX
pRJVD6DqipGmpvt80gO78CvdbrPVJizNFwWc2QLGTdyYRnAWYpFT7QFo0xVTxJ94QNIJPYzxbntP
qYNq+ITND24V8Qlped64+GJf7YjKwh2+Kx4KoPm/ZwiMDohGHfVuqSFqeVjQUEosmEefrOjNt2QG
iPN34WX7KCvW+1a/i8xr1DEr78XH9vyqsqIT0KwhEXXicUi/HL8Dz8ML+8InIIm5w/rMW8676wXe
mB3raJ0zDUoUgFs7YxX2R4HB+jOFcjTMt/B+pXPzXytjtkd9r2hbLwDPWMivXCGNN3fnhJDKgjW8
oQaFqeLk8cwbAhRejEGvSvo7zmR6CvK7wtZU/2W+qygt9s/ezYUBumWe5ZKdVE/mfJ4UpuGtwsQ7
K1Be5u6p0T9n5RnxMKKAEsqKOY1N6zLk5btfvWqCFrt0Hz8wy0xp9xn1DcCInz1MXfr0yB2YWpa0
NcZ+zAKMAv88M9tHA1PbHn9DGJJdJ5vETNUJg/YeSw5M43CsacyhB4snQHZOe9GPlYUoM28g7h0w
Eo4rpBlsFI0wOFktnaC5wESdHWIv8/I4AYThKXyY0VPI7RR6pKuEqLmoPEQSBSA1Penv+mtesf10
bnHub0ihpM+p/CBK9/slAZK3tDeKJcVHwCLl+Q59p871mMaa3UG9UFgFB48yLu54nTBzuHCm0oOw
dQCY2/xvr5KlFxGZFg7qkdmTP4kaMFo2o++PfnNPx43CepuiAhVpbUmsnE8ZQWbf6V1MZt5ac+bI
bTtKM/P6TIUTwk3IdmwrNVcgzdSpQOw1Y/zFTCYWTbItXDG9xY+e4pAg411HGGRILCYRh2ivgEbq
7p7gPWgg5Qh9LNc7fq88bDhSUn57Puvw2Tt1l6Rchxhc875iv1oXM72kb7vASKBsuJeyHxOsGsxN
8jyR5bq/0KTnBDL7s/Z+tc048txhvEfTf8EX3+o04dPSlNwcBms2VKriafPuuQRW/WR3n9e79rGV
rsgoUieOe2iVdkDGX3UF8x7/nTGmATu3fi/kD+y8ydF857n3a5QVnwAFKDTNNwzmX2RxW2lcfRsk
7dPVzYa/3rYHTaPxK2GUnr1v7kzzfWXhFqljvMGCgMjgb5gtBZ7ulFU++A1OPaUaSdqcHDzv6Trq
94uq3fabrAa+pFFHnfJ1PerjCe/51hIUJ23HYuloZXEz4ckJiEZzVf7+VAwSI/uPzWxD9q6do9CN
hXe7aURpuLlXJdv/z5Fm0OtSJRJDWB1RqQACB7TNE03ktW0YnZVLpLC4v8r4pyeC5yBWTkQQveso
nGUK2GnBOX6RVhcyPIMFI+vgzYof5c55i1laoFxo2sGbUm72X2i8bIgtyd2kU1IWRzsOeyoms14Z
IJtc7WJ24izeJFU/8dPMiziTVh94dAId8sa9IceXqK1KNuXza/Og98gLPbXxmDwyskYCfssuDkzD
REiaH/F6JQNk2hgNyImnz9DN/TG/u4TbnI5O2NcmxfLyLh31OmwWtp7Q3CuFiTdPyN07w2yWcDIU
5dzy45RhnP60hLiQUTydefkfnp2ZEC360TLDjAA+hgd6R4YP2qWBx/y0QRZXYDFNitt4l623QvZe
Ssttik9kgL3/pKOcYkdpsrgxFA39NlH6gTM4WDAU36eEDuFbOy9NKShuIbTe0UHFP6DWYUVn5bIz
H5xoHYDB+EA+Wwl/0G9/DIVE5Jb7HKaQ9qgSTUs/KCq+9iIAEPjozLjVEwO3c9E8Exzv2N7ujWZD
nutmv+mz2LQ0mHWhMzxLqUAxQcWyuSG5YpgSm9r47bE3XeBgg+SNtX5ymWLF5fha4/IOYzLjW29B
YsWJK0sOmwyEIHhERJeOAdaUl4CTE2etZtNX0pl7O3rDkvNUGEP3oKjMGFUcBf0wVL+N/n0XoYKg
DPOk4iTAty6X3Z4ZuFN7BB32VrR7R9KuRcRfA2mmZ6EGcnmpIrO9+cTaKG1TGnt3z8HKXEnhn6V6
c9j+XbaKEOFVnuiPBEKd2pXNrPGHELJN4jndHe5IMMUqTlZ23uXphogr+nCFF01rAhVB6mLo8i7c
CkKkbjtIozMjKda9r8uN9uTQx9ROFnVpLDGzkp03Aif1EHIZNosEyPntt/OKBFHiC5iYVJAVF7FD
fVTl4zTblPC5Bcku+fsup00o8QcZSq46OcZPoF2rdIranLw181t1D2Q7KXNF/AKwpWDsJVSFMmUe
/hpG/aYel0BHoVspuz85Sj/5VMtZoAOc7XP47bOlrKFH9qBqV83ISskot0BU8j6hd5MWz6dfK6zA
VMtCsTIhr4v3MOKg9yt0S0G221cd0CvgJpgEQCGrFd/9T9YymXT4QF/5wmcyxwMyqWBDYtEcdWfG
i5EFJRJrUM1k6idwEqWf2cZkv3NHfoSEItRPZ7KJuXX57BrS2zg4jbu98wyn7Zu+Ias7GuQ4nKKq
3d0Z8WYXW+GffL4cIRw0pVSIbsIAq3KHEMAnlJB9zY2MGqAjPX8S7umDoZMHeMemCKfFCQ7PHObE
kRXJQoISyGauoBkIj/cfiAxg2oPB/WLmvD3uDbyFHIlE8Th1UGrYClcIM+sabicBU+62ia/xBkYK
DaA9cNuaOGUnlcy+4epg+Pp5MM5igFaiO7NZc7QM3K2Ndjvxbx4qIsvK4s8DTZKtx0O2+EX4etRa
Jm+nJefEoHzwa22ClEMFFbRNA+t334TxvqoudoOB3UiVIco3T24GChN5dA553rMNp1Q46F0wKOSo
NlfNmHCZ+a63mIYEnVf83PZ2vbTy/eF9GvAglL/f0zSElfnY/e/OEkWfSiq2LFcSg7+AZvrYi79Z
dbfY/68K/dBwesBBr9/zGqGgNuz2FizCgSFmwFfxXmH5JSoCECsQS4RlrpMUzon+c8YSHQd0N6gJ
W4nDY/81BVXbUPX5QTVDoz/y8Y88neVycHWj8mg81t8E6RucVbKgYES56bubPPomE1v+tMwNQQJ/
GyBisUFDoqKqJMG3QGEAK39PRtmZVX9nxbinCYfeSMGBNgKTFPKLb0Br4YR/a9KDEM/ue8mgzBjX
S4qEySAgEWQfHZ53YYR8fixvgR44d3n1oTEWWb21UiSHkjFcNuflFj9lQpmKpPa+aModOLWNd76o
w/QENGJBEcEOWM+JHMo2X6AOqOZhODFn1C12VMu02uwy9SEtzZBqOQ5xUBHdLvq1vSX005s9zRYA
0x2BsF5+8CO2RdoOu5iaHj0S7HWyaGyW7w2mJKnqT2hQt/mBxZHGRFAxmODgdD9jj4Fs+x8kqKzL
RSs5s0cI825+MXbEJQ+fkJgyCc+g6kXkOUxy8HKu6ornWT06t8+9N/bE5uX9JKkHRcqkLYS+EV93
x0qbM184XUhmfd5mjwi2glzclYNg/hKdRsp1P0A07lYc+KU20Gy3qzy+tmZfkCiHNuCe2iXGXVO8
geaosBTwvfZwLe6X4GFkLAhy1UUcBHhmnwXD7+6x6HcDOFK7TYKO4HBwP/nfibQQnavZpmJ6rxiO
/9vvx6Waiojdvloq/LHYxbJKq8OyZeEKI0/vhGLMOYzV7M7awdwDygQo2qToBUXJdQQ2fistNixP
GfgkGApBIexpbA6HF5enxZJYTBQ6ZcvAEgHOOftY5g+17ebWSMmp0KXmBZMzd3kEh/D0N5Xoa4zg
u/CI56I6PLIz6zQEQySHx0h530uCfFX19DFGL1P703Dr68//Pmb+qzsQza4wiInHvylsb7Ltp+8/
wsxLnCp0IIdXQvnai70UahviIuUCbaLPVqjonuancOWcztTxP8ZvDeoMg3/XBbGCKb3V8sIF2YK+
Rc0lFDBtUF9MkgNjW/DWjsZmkkt2HQ3pGYdVyfqtjuH8kmzrXuZGEitPOWX6rTAqe7v4/3dE9xvm
Tyr/sfzmgSeazWi3r14/pxl9xYsZF0dkx12+PmrkqrG8vyUizqWUuZREv3ZIocesXYIfcf/yVIgA
bYXku6DoUcyquGoaJ+KQAX2Dg0BgYshZdiaprRBgqQUs1gbAZx/M61JpaJ8FcQwvkg0IaesGGXtk
F8XepOT8wvn4I5r/UgYWaH9VSfVXXQt9+XPkZnYs2srJ2sWIgmlTAoUJvKdnf0xzKLrYMndlDoBB
rsocxf+OdQWiuoT8Zt1NwfdJqIYcBdFLzLNlcCXVzsKbGSerWfO/w9sZM23p2XTeaQ8XQPMMHt4u
zXHNDU+inn3D756vQ37jiey49mkXg4f1dlOINOWOsyQOE53/P19bWPSKRTPUjxiBfbef2HcIrSMu
rJ79vy4YFMn+SI7v9A6bS4fxExWyBW5HeVQayP+rlekrd25z+Lf5xf4S/z86WMgJVPRdsqfYtUUd
CLzRGfpFjGKMQUeFNSWv25qcDEo3bNGxDdTnC5aczZQVIQ0+f01NejYEFaqo+bXK7OINauxq8Ung
+yoPW2HAVcl7UsYqfVKGxiDb5vMFslvnC+js/VF6WcQUhsKFs0TaiQhwfT3cuDrdYbN36VIOzLZi
NQYlnJfM6DV9LgWGHrwxQ8E9zFS7amsJ5SXNql+zjygGdPB5T5kG2A7fFbb5yJZH6Ja/rhl10HcJ
kYKpzaWhuWGKbV2Yw7TV/3gJyGs4h4Xj1yaNasH0GYnyApWJhsJN/21YLScuxmfcmA5nef0S3fUV
PvlWqyQTlumHTn2qacrhxRy3Jhlu30rIjAumk7DyF7t49QJVE80wNcILtcjaaohQYWJ6HwLhl/Nn
bxqu8ZvmynOY2MhapSMxKu1AQbdUkPcPBDEAuLiU0eYIqlA+s1w+ipiRamK97bC5cymiW7z4xJVj
l9M+ifoRvEkhrjtiGPbm9d19OTMeHeIRZ4YA6gRLt0XcpfWCoGtb6+diG9waMmVY0BE7NSauInG3
Iy9//+P1c3qOZi64fm4ZbhKZz4Cd1ndcZKm+ty6BzDTR1YBbqldfn7YwFsc2EWLYwJsxd9dcduUk
iKPpeOMPBCfbVnTPhhO8/CclshTp4NABkCNAShVkvOK/w6rsHya7DJPWbWIRAiH3ICCRIoxIHok2
OiujwAkez6V1EJUSx50+8Rdg1a7rPjYF66ncMVuHhbQ2FPsGb6RbJCa3yttnSygDa4yWreD5k6FJ
A+nAigYlWjf2qX9EbNh9OKH7B7gBk/2yuXXZFFDkDhZMbaqUncwdbEdcWJzl+7yFKk4hEFt5Cqts
KOGtOkxM0LJsBhtcgMhfiXR1i1+wR9w7CSAFzmPBQVYERstabvT3trtuqIET1y3qhB+iMQmtixtc
7RPFeH8jyNsyY9UitF7d5WjNiq7TNbcqIQhiSf8jXzHKxrQ0oqhsydH8Waquy3lR8zEVs+65gLug
bujSw3uEYN0SqDp2qgBHfSDW4vE+CiXxNI2XHEJZMX5poRHsYHRb59PFooD1qrOCJBG3a/C5zTtu
ibBRwcxpJzVgtcgxQPHldGurr2PvL+zgDv+oKz1a2QGxYQGqVTwsYqgIeGfL1Zw8hdEWYENET4s7
WdWgJzPfLT+to38oBcD2R3sNI02jvNerT0RXWiHCTo4LzIqwRhIYN6JKRA8oA6DZasf4JFDs4JnO
NqbufDydMBghP3Kl6wGCxW6pApBIh5xZOy+El4cTkwenmh/yytFimNW1p54HYbnGdQJpWmkBEbyF
FTbSnfDbjdKVVq8aKvmi+M//oAG5b2eyq10ZQ13uwMcBOpY5C+aMVhpPoEIDGo8sP71skQQZnzf4
QaH1zZWELxrD1zq4kLMWdQw2mco9sHu1Cz5JXSoMC5rynqGyVNb7Ripn53Xkuz+XEJpKWOs0n71e
CWgGpfAS/5W930ZTYCjQt2gvs3YSiibcmeuiIZS1I7uGyVkytF0jBWDSsme2Lm/cNDuA35miql/3
1Rw5Ng0tGY9/QgCQ0IXbNNmCD1FPphbX9FH9zmKgkUp33a6oU4KsHyz1MWR6544LoOf3dgRpQnOW
BuXhg+v55ENVfvF+o8BUbionHwXDYa1W2Lv9R7Ae3fWC90/6XbeezYlO4p4oc6876iKcHTxOhdTc
OSYJUnhzzfdWKAoFbbRw3+2Er/hrWSvqONeAka3V2Iz9qgx5hKMQN/eoPx/arQmhQtzvwYsNu2M6
+K9N/8OtTTYilakcBWvO82AwZQYVY0u/nzlNLfhyjmKXFYmJzY6tFsmV5lwg0qRvhHU27UrXsRYm
F/jmqFJEkkFLoLPEse0dS9yFp16TlTqmoB1CvG+qHtbT4CMkRFtId1VZHvjkmqtO8xDQi7TTIiL+
v/vXVmbsXytlQigQ0tMx9/WBFmdccZ5uGbkK954bm0fUP1IIdz2r1a2JyEqlqIELiAiZ0za7asUO
qkExxInQ68YUqDuGJ3tI3bP/dCzcrWnmAUKCzHAT+UXF3yWdTUCpSyxWlUKOfcTpyIXmdkOkkgjI
VlmCYME230G+luj5UQ6GIxD4jG67v9/Ofp3PvNtW14Ots/scMLwFN5nfWZxJeYRGl57yHsFMCMWU
MM5OYCGUribwR1WKVN4VdWVocMKwYu9TELzBf5uGLfHHMeqW1MhTir6/KE3RkkRm/I064Y1eY4F/
MshjdicvLIBDkQwOCkI602PHrxNZysUGRIS6dl5PxzOXl5uHfO+1iQh20viq9RaH8nJbmmYa+gc2
FeaurH1gEB5yHsOR1Z6vqLx+UtGRQhyqJH5jdbO20TZlQBG0gzl4ff2YrRV5jjH6EGvhOHPp0b8x
ZOMN5udG8mZEhf7c33kqYIIaGDCus+k3z/Kyg7TMtnOCl6jipN44wcCHfIZ44eSsl+hDDj/cUQWE
oS2bCQm/qA+zcPrvUwjP4zMVDWU5YfLyhppytijaN4FcMybSEaxNpHaVslNN5r2im0ccrazBJeBP
wTznGclYapzVQHEExo9qApW6YNq9H0OPCh2stB+tyj3wmdGZQY0RxUW+dpiM9iqt4llKopfOOSxb
sZSdpB62AYvLZFd381US+9bvOfI13TkmX8SapMEA0x4rndUKl3lG9KQ6bSDZtQqBLqqDM+O3SJLc
M0Aq7oLEB8X3D+pbI/2pbKNLa3fHIF8xDSrClPayZjc4rTTk2YStRsghoSXzuZVcQhD8dr/s69vG
0hzkX2Dmv2FsE1whaDOocDlveWMaByzerHmIHUoxERwuUxgZmBb7nC1Onh7nqmkN9fvO7Ul7LQJH
odBz6fXUB8hkaKZVQuoF5wcvYIAvUR9HkrsQID84L/XAj7NQsiqDtUf677UUJjCYdwUy9JM3hW/P
b498g9g2V57RUCHLXjeUM6iLKKC54ANNQaa0nr+yjUtLEINFZJ5E1lVA3eClGRKQCniM0YVpafBe
mLJ/Kz3eu3zDMr8rdmwJlTgq6jUS3236Umn344AOUPNjPNfTVGtxHTVDdQt9dNcSzpprB84jFsmt
d+cIs3ozlC1Ea4eGTomw11vLM1Q13zcxgYXyPUELsJqx1lA2SUFJvZ60KX9wpD2draCVYGC4ykOM
dr+EJ5ky0YRcKSDdu7lI2ikpk2i05JGy9YoDOwSGoLg8f02Ci6Yz5jvBLXo8WLqlOQgTjURoJCMS
zIpcbfxINJv0tP85gSplZwen76fI4MWnWz94KA7nockaRK2UAOhJ27Beb8qyui8tLkQWjzNqZ2fs
QoLHYV4RvpBLrosdq8YUPrhV4x72TgIHdSpi1yPOGNULT9imaBAAs4LQQdmAXsaZTcshXtAK6NUL
Ve5Aq5Kg8//CGelX4u0nhd72yKqAmMZZ3SwxvIBJP8lilBL1VG+BC6iBUhz8tzvpBtzeNYjWQESI
IncLlFMH16aK1gzlu0I/aT0XREGgS4rPYOstlkWnOaj+Tqz+nFgv4IteCI4N6vKbQQ9MuSTLg0Y5
Q93gxrIAgxFbzlE8lCd54HEbFhRsDVHD3Qgis3WIiF1nibdbGlpxPC9rb4F9DYLM8DK0iESatPRi
5fkS/g6PXKiauz6lUJxifsHOKRQo1CBTntFCGYsjqg7vwCq0wxTvMXrcspTMdWKmBoOXC4IJc0Ti
JJ5j63UotNg7WWvYBXtv3wd8AeBvJheUMcIAU0LJ8jyW4xmuEpWWagBDKoUPmBKvJDqIMGfJ4wET
TDp4JZUwdEL0MbNHiDEWFtt0tXk9gA+mVBnQpwTlP4iRVgpVgqLdPCEuNvDsQidLoRdTEqczjdFL
D1MiPardknHWbR+dk++fSVqHc/J7Z7vzyKMy84wWdDbKXe0ttN+o8TVhRXSEY8aQMq46bA4Aps6B
HyJMguKE0RnFxTcKFBdzkz1gPb3Cs5R7xB6AhAnb3TACFT643n4867whE7c6nNy3jcEKvwlSATQf
IFA97cl1//rGhHAn9JoQaHsiShdyiidio8oPmVZdErN9evNFCqJkSrSH78HxUW89Wg+pP/M8jJR6
eLuXbIN5um5Cjku1JwRIwtlEwZ1eziaL8jIvYnB7gqMlvnXrvTja0wiu8Nu5WDeZxNsltCwgBCzN
HbwcxDRa+JDHuHVkvE/HZ5szhc7+5yu7tAMBSLiUGDmZf+cxmhvaoLuPDqNDE+m8T6nziwgpMQsX
1jUCCKPhRNSBf9isxqQmrrxpgW9iokQaajISMe6UvAqBonn4qu52JTC9abSjhy/s6gqUGEcbblwk
Af4dAIm63JwpmW+3FAZ8yvnqOuIlkHyS6aYHb8rOT8woze4hJcTvJ73piZL5/jspZxZBlZRJu7mi
XxtXhRy1voGIv3uUOLIt151kwfkEFr/KNc2QJrumWDNrgFjTqUi9qo/ZRzJwsFEOHhMg8DKt2fIc
LiiWiJnl+hzzFhvoUpcy9jzRVCb8OwWZlys0/4ToytAVev7/z0oI9Es1Y9ZsfyUx1WYlSmOZnoMC
F3QVLlXwacbSAVrW/fLNM9GsUVvBHpbwRZUtNS4VmnVEt5DYyfAFEolnFiA1KsoSXlnnQ0JOzkeG
zNuqG9XlkgbbG1Brz9cxzke8Y+KrcU6IN01ZBDEjJL5Djd23WNrkni7yc93Iek7+7cD8oLxDVl9Y
TMzXIF9Fr2NN/NVv4Evd4EhJT6D58jAbCcSbgerc56ilxFBUN1cNLlA1F0ZafmJChPbNPM4zmJ+z
8Pr1W6AkMlH3Xc9F+IQlwh6DiaR4P0Yz0we5ew5pc7+PWyptBSDgm+SDThTVFuF52CMo5YKxLgwB
kRAnUDAxnEuXaBeCLLbGh7sNltEhNrd9mgtuBJjuGXNV09CEMRKc5YvVhc+tKgWP3yXXYQGr1gk2
GWh4nqDoVk6eDHlepJHXkb/zVBY8hkQtpe1XxKFTDejz0C0Ygjtx4ABQ7r2Alj5Flrcj7RYFzlLC
GRu8sCWqCmR5V2cF+aHaYFM0z2MoGlVPhimbsesNFrMMM0gld13KaFbpJuD+l/nW1k8GJvwV+8u+
OHI+kbuD3I0MUfGhFjuXodOxua0JA/6vIIjo2BhENPpOYEtsQv79DnngN+NZqNQeWQOha59Cz6U+
xhI7JjE5DnNeOBwVNBEHKVFkNzR9GqFY4diGDVIk2Sff2tNMJupuP5ooxacQtHJiaWaLgs0asoOn
4UdpVlWECZhRyG6uLXfuUHABRK9moV3W+8dnMH8ig50ESrls5EChUT2f+/ZmB39T7HKvPfU5x1Pp
WhSqDVwHHYdgWSGIUq+hhIC1+nQRQVnQcgSXtGj2AQdrsKZPs+MlkVMPHgRYQwGdM4FHvhXKLS93
uLpTRe4AeqgMmyw3RJLdca7HCrbN1J/vzZw26DgAHljX/yHBgcH+Foy32Z5HS+Td3Ky+gY4P6vXj
CkvTki9NDQyMQafeaQ9P9ajFc6jVisAuqkaTSg5ohx6re9GJ+pEpFbBa2m2xsBc+H34WjCxrycX/
v5AhvU2JVzdvji6HQPafBUauCA1MzYMgvcfWQhiyeXrjmYG5que6sS6ek7O1h9RyXvofVjMqJ/2c
XgBgnvsfyG77vsc3EvRKZmuOPtNDuHKjJYOp9z1DgX8em2cZ7kxVepvgEqbqsbZOUkB6iXvTi8Nl
t/BE9/Gp06lkGCct9MdZGIMVF4XLG8VcI8iaRfO7TEy5vow/iDAzrXmZC8krpDw/PhUDfdUt0EM7
lAB+Lj+P9biTR7kOgiUJDUYgunBB8GIxJkB7FS4cJGE5mvLA7sbZbU0V1OWOA+wlv2CPLbnhv+md
/f8xQBpWOMhdTknU4xrFyosoUhU1inxeaqU272SlsrNLFMK/gDYqDrF4DFoNe/CS5ECtwe+G2bc/
bI+cXfpDCoy/cmGR9KI5e/ocQL6QoTQXEWgSdDXVUbSGrZZVz1FTjwKje1w8ff0xbkUXju/O7Eoq
SQa/4LrrBdNFWvG9mDJA+0wOLDsWZq4vQdSwByu5b0NAKzvvbREMZO59ztvzPciARNf6/el87v+e
yFvTVCylucwjJhKcIsKTMPF+rRba0X1aQoSU/nCAcf6Z97rNH/kRryCufsymuQQBpgzp1/MQSUsh
T0RSNu5tkA+VkeN7YwByB0Jq0wvJcU/ZDuK6A9kSFCchW0G791XxYlFaUWqM5Rjv3Ops4hrUYpug
LvZdOBEQspj397NTr3pqv9JbY6O6nJV8f2dYKsQvNStsh4sHj30tFadE4KH2hBZ60j2P3QKEp4lK
TcfCeEZ8wkMvehZhaWPKc4bMocGcc1ugwA53W173h/OQygLFJK2jWPLyEgMBxPZPapq8Q4SzdFCp
ZfQ9lcM5v45VPQxfgduCse22W4YvTy3nhAbzf0BovG7IKi+OowY3wxrOJwlGBN3mjyyPawB6eYK7
noGmfRVlT4GJ79YKRJVmOMjEMwxjE/erXgaKMPxdEONkfuUEH5F80DchnJ/Ps7zqqGY3bJLRPjmT
yryGC3DLr2FCm3gh/M1mkDTSvf21zdMdZhM2vibJM7Y2rhGztvXnzQLQxbuJCfmCd7MSqdnvmEQP
BtlgIixkV5d6vB6pi4GrG0zfoLLDV5s5c5Xeiyh0N3RKkqlS7Mp67rkl3TOHbSWBzjkOKNeyoJjG
cjdodrKE/kXpEqclr5WtBmvTPVHwcdfem1YDmZ+75bWWZue48cP4AgiJzvduMg0yopE6WOK67R5J
mkXE6CvUkPuVU5mRiCy5ylqflm7ZzTr6EgTFnmTBBIfAybanP4wyMPaLiXYM4X/YPEJohMj2cri9
KZpXpPAqztGsSgzpnHVvuO7E3auGV4tL/5EFoNwpR/fJedCb9Q4PSyhRKZ59jqoi/4saOBIupNOp
fum9LgSqlgudrCWH0Awae/NyGz2anOmtU+t5sq5C8U7ZkSjzdNsh8jwkXBN4hLUCDjcvtaSGkZeT
Dt/9YosSplQLlEY7LSoKa1B/4ik1UCRIXuv2bmiWkpFfyRgavrOYIsWSPSCfTckC6zoiWdK7I9I7
j4KArjtRC6vnj0sEGz367EV8qI8cTmvadmUy8n0xX717928/UQTGNUxWK5L4zRnre2P13tUC46xR
rIrJO4DD5RNZ+OSg8q10hFUzq5lDU1tPQctYdVm1jT/ktIBpS9cAwNWagjg7YJuXPZop8vvmkTkV
q63vZbaQtZ1FYRG9Eowr+hDIEaKpufx5gvcc9QsQJIHl6ft4MfeffVRT9nRyUuAQk6HmbEwsMyqh
K+OBkmuzkL0+AV4TAV8krWC8Ws5IMRGSl03ZtQQ4akHKLJNhO2MsQoAMZO14LZEjDG8rGw/k0wRK
flQJptX0BjHAEw29vH1sLcua/AL9aEWSVUJsM1hZCjHtxuxA2PKU0VT+Hm3v53XIoDq7mR1uKdEi
B9LDsjdW7sLS4jiFcag/dapUWPuP12apUXb6iQ6DysyGf4Bla22jhw5hbLSd6jtYCrZX4JMd4tLV
NJBTqzWEa0NlNnUtBbWiSpC+9QmmtXelaPQIgAt4XSK4nr1sIyBFfUq3f9/lnr4Sp0o3qVYgxv76
lC5Fe5zjuIEZvSoKb1k4en3mtOrIXLh1OSdduUByLzV4Hgm/frLJDL0Gji1640J1wv8bGzKQEvw2
UXgOEj7CDpJFB3IHeqm82LWh9uqfYR+EQ+QnYoMHRqDGKdzmm+3lQcE03rxgxldlQpHdPxQLv3o1
prUOnsX2mjqeFA28obDL8SpmkQsQgQm0PDgwUHXWu+g/MWf7djp7CdVDIjjwFnyk9Okba1cSkYuL
Ra3BHz0s7th5JOfg3zAfdSkQsKkHfx275fqGW4rTP0d6M//S2AvwzNdHdR0gim1Vr8yA883DJ1zy
xazBkNZGrdju3JMWqquuPu9TkhqQrbvmSI2CIW1qc7VfZZalNHoMtt+A/r+i6bdPgfu3oY1jQdEw
QF9joFFftowva4KQUbAZPsdbTRLGt1HOEi/NE6FmCXBRK+sLW3VjoGnAgjnCjIn/EnFeASB5Kglt
uMI9EWEoIQ+e8BRzQyE811kxXkzMQRlvZsrQ4KYc6CA4+x1tLdya+KoE7vhsBvNiNeh+OI3wkw2Y
VS8o3Py+D+EKwRGnydXSqXTf7FgQHzQsI/8TRXID+BoFgbjtLxynqiSyYNZ0aqw5G4rtoCQpdIOT
2ECjJ6fdBmOemJ/eOSG4/MHYDZWWl5KbS5KRYpQoirqHS6knDtMpg5SNnhyu8WMDDqH/6EQ1zgU4
0pCAf6Gk62AzSi3k3V3iCtJ8PHt68s6sjIkyfFgzbdRvS7l4/IQb23lD2EcBYI6B+0LnG41rk24x
SOhjP8w421qDLKHx0Vj4FvAOCI8QygKS9tQpQzpGL0NQyLh1RULWtUHElYSkltRKmq2WQbcYS6im
5kGSyXGMRII4BsDQ9WDPhPZqKr8nmt7f0WhIy3DYlipCr24mWYheYCApD8ZiNejEr2B2U3gW/3JF
/anMGm3AHYArto2QmSXrDFtPBovYCsq1acUzZo77fxFGorC1Vcrnv92//SYaQb81INuQ79a/whyI
c2uUO/kGvm6ofAXruvX5ZayRQwQSGKqImk0xchPw3S8FTIXmhS0+qxGtFK70QMMmrrGJ9Ql/YVIf
NAeNBEy339FV3xXQhY4a5gUyDQ0B/PP+KwCFdtrf3YgfqIHfuCe25xijjKdziwOoTUEruFOJvYde
8wd6U83rjn+zhJdy8oNAfMOvRvEBiCOBoZScia8Ao6AZ2kMuEcn3GXd0ee8Bc6IF+lamGs1ROF+4
ZFzxPT0NuZml/VfWZZT9WrZYSRvAexpko7CqnYFxPQV5MRyXSttk65rvG8UOm/W06PDN8SVlO+S+
Tb2px4HsJHjEMwqrVP2Ag8B2lnYghXFTyXyTUd53Yjxx49i6S5KatLYKFUCeKiucYMh40xjeGe+m
g8VjDfNlKchpgk0H/sEOy9Tf+DZAcutpUKwCDYunacvfWovbf965UmsRsAS6o2p9/DQTiGA4J4gR
/5jm4CYQia14fOTfzNQ4Q7x+/WczeZKPZ+XvTbuq+dJszMMppH2nf8cedu+QqSkrpoPOuVg8DqWl
/Hvla5GY7Ygy7OmAcIse4ef6yiOVKFzQ5JHSZ8lYUX2K6rJWouudWE7yfEI7N5BI6/3Zn2YR8wVI
V/Inoy8ZOqKJDpR4+WEUa1NUbZhwv3naE4Am4OYGoAIcvgkdnAEuooRxIWRE66Ni9jmlFX51Gw3s
8mrqJdSQr5Ev+xO/nL63gOP+wFqk7NB/HsZJR/8XkS2PeHqpq4dt2ven4geOvUw9Z53AXGCmqCzz
Cwj888AlBCzN+A1Z9SivGWG0YAhGFaKlFyyCZ2mucldOZIAekQsoCBPd97sNGrQ6z0NCE2InA2KI
kGUOWVLJWHTq66lg1UVWSEcNuK5Sx3FzLsTmRUhOceT0C9YzgVe3XaHtW36JQgK5G34sEvQCYCj1
BuZwQxn6mkze99AfgM0DVl9w3fuMvCbGr9NXFjM9D6GokNX5yeXEiFZYvsIaQy3BlHWH4PAxzBlr
Sm0yZ7s7Zzx+03Vigr/6p0NKkoQrGanSbR3qiay6SuolJdZVmqOPZjKaV0lZ9Moxz3uqeGT7Ih02
TFUsgvVxHjWwyWBl2xiccRfkChRvCF4Id1sZW4mAi/KtNufZ3Jm4UZSluGcTQkNKsgeP2JalwdoH
MoJWb1tvkUYwWOIifntQ6Xq5uUrp/oy7M1RmtImgtTbLcQ26YU0R7iY94yvpvsxlcXvSIYNUP7zG
wJUgr+ZIx0sQT+1z5KB1nubNqBt0kO9ZrMDyLlSPvki3g3I8ypNfQHHjjjGIJGvze4wBHG/fvAfu
vhEEV7MnnJiLccQOYjAkhmw2weh+WTVGh4d8OQ3W4RJKEusA9ICOrxNiVmZkjBrMEkCxuAoLXjVq
K6FAL7ciN8G0J/vneZs9IyvTMGGBay2Osf+3V+1AKGpWueWo3ZdoA4Byoa/c1GqeCynIoxGUaa4w
elHgq9FGiOtvkj0Sp8Tri2EdoXuvXYoi1q6SaDaqiO8UhFUt4594x2rV2V+JLjIu3sgTs2R5vh0+
Cv+0LBlZNVm8tpXew3bdaZWXMDSDrggY6MF/v95aS4gdKvWdrXXrPDRLBNevP3NCQA6UwyQ6QgwY
/O6CACI1TTO/evFNOeDtwmzpy3E427TJsJ3Ys9ZbF3cpDuZ7FmqY/nwNixAaMcRAuhMVo4fF2Yvl
W2y2YHgWcCui5+bHZGd0KvyokgJcch216FuIjjMooous/RjAYDak+2Cgd3FJ5chhlpwYdP270QTs
V7O5rm878yhtUUl0L+VL6h7iUZrgNt4Wmrx2b9Zgw1mfk7xVBTw1Vh6nMea2O+turPKgElsbdSUr
4gmXeuteH2PhSw521yW+nnJg7QtZzI770o614pAapBIzOTcwbogFeNBeNzisB7ZQVr9L5mhdVlns
5BmpRwMwBKiA90t81qjoh00/21cUx5syLxk/XZguTsrM7O6jX/CobeMXO1EUviatWhWYJTCKdr1m
ObkBasoX9Yz6RoF5QMvp9usu1++CXs89DDuj0uHpeCaHwxKrkdDpzKogkR8ySydeU992n84iboBD
uWCNISUub4IzeMn7PBS3mF517IBNLf3kW4bhjBv0DPC0Mgwn3zMRnlxNU/vEJ/c02HdgLFbMFbGt
zVvljdI2+LRBKzJ2x6iXyV0bWS1pdafLhXWmunVMqvNnly1sFby8UO3t+doUVZTIwuf+GXfxzBHv
VwdjsRU0Zz4Gbim5VWULPLvc0nTaihzHOcqgpwU+YcXl8N8NWRagRy165bfnyR0bxxJ2/3xxnNpB
ZBccB39WR9Z4ek+wgqAmIrVsEb0Ueuo20fNYjx9y+/Xeeq0acPRLtcLnMBvnPjWZpcLu3MF9TsOh
Dresz66IwoOqJfkTjIbP9SDtGVDUbUrQ2qrs8BzGKvb6RFgAaXv38cBIohhz9MfqI9fKg7LQtT/9
L7bV+JmpArHhHtM5yJTW3BNIZw0/0pE/+YQf3G8fT+ZP4lYiUTdCyXHjRCEB+iLlkijLs/XJg1CK
azyuX+wubJr6OVbl/RpyDjYtnuhxBjKJeuvGIY2Y3mc7Ns/J8yy/D9vlIj5nA52Up6Pq5AErXWZ0
CvoSd+nDcSdrW75EVLX7LhfRtASQw+za+HKyW58bj8WC9R1tR2dGu7+4sEw7/pIaCCPfYY5pDDKn
Vf9lGLshIupA+0TNt17JG5CpauFskWZ5ngaVGuJuOtXjqU7VRV5aDzXT3cTJANCfpfNrCfjJGmuq
M4QUYe1fJGjP3MEyKWXzzfSm9FaHvaWh64NPde6UIU64AkguCuM9umJsWJvWm8Mb5YNuGD6Uzg3N
bVJwDtIQpaE0dPMEe890AwgL5WBnN0CgsV6uN7shvDNuEm7V8uOccfyqYWt9Lfmpa3QrdPj/RbD5
aTPlIZofyF7kbNH6rG9ZL6RKSfv03qLEQI8gOCPuP23030+Q3/RinQ5nikTexqfVequ9ehwCe/80
VKc83amY+1ZJtLk8NdLYMH5fdJqDo1Xrrbamy59AZ52VhGj1sV+Oaq0D5JA3M2mRamrkyQEuG1He
wBObI1Nq2mGXE0BDbgssY3T3C7aieCdJOPrCjy78w5E4/zPyUw39JTEiaAkqu/XMYP6UkgPrqN1q
nj9TUjCIMqrpcgu0IV2CyptXid/ElmvFjTMxwspILFyd4Tm6UZo3FxzEPVMzWOOm6YwwvwqFTc47
PG9cPEPc53e9hai4u8xF/SNAIf/63WmNv3rZw56vAyJAZkMGX3OJlsMXTH4rkwIUeCLZrX8zaR35
n6DZiZifvZG/zqGbxaUMUUCupElc8hZhMRtl0vKHrKa9mflGWq+WckDpm+2M61sBB2RSwOY7CWVb
zDkc+s1dpVLLPazf8dBTEtXBCvffAa6dTCU2j6wff1Bujh+m2iLOofaQH6BzhE7HuS6PW35fo7Z9
4bwKF+eHtcdp9EooQ4BQmR50r2FCSdSjS58CHmlFLpL/B6lYIvWcPBjG6hl38M8jpMq0EcuT7lpB
9CLisSJkjKmTrOwuRxFD8jebld0kkFCwwbY+J5M1i8KaPbZvcZHSHtIVrCf4tVusUz1gk/Q2QJTn
StxZ4/TBOVV/ieeineIq93XzblL9oOdTpqlQNUCmrxrpULHGAgVgY/hn1QrxMFb9VYzhUswKrI5m
gv70/oo1fWN3yoCrcoQhqcREn5vvBNZVweHAv/rYjsY4G2AeIp5FtfyqSRG4NAQ8VUJVNdpGjX75
HTISm8YMjiwehqC7NhYzYlxcZJB3RZ9QhmsaT3Xp7Uf54G8aFvg2Y8HvK7e38XuYDJTjV7vdADGS
ECaYSUI0Nl4a9CedKp3OcLVCM7Jxcl90EbY23Vl5axh6D2TPCfRI0+/aEw6tKdzp8QEhcim9IR8a
k24JVouCX7EwVJe+/3oJ633oDAKmgP1vZp1TlCPOqa99rzNp2hmNN6/nFrGbN4v8kTZobuA5a0hL
pqcYG9smq3hD+gLt1B9wNrfPkG5YeAongeXvYKMGVBrfRXl2RtMUVHJjbtj2kUu3PYm2tPukpVY+
d2MCEDA9Ms/c0FWG35nxig4AYirOQrmAvFVu+wQBW7jZG6uKmrqd66dmNR6uJF+/dqOAILKq36Im
2yIZ8+tCch0noSEPjH1+SRkDhtXAykowPQpJtchGQkh48s4dsqhHt08wamgnxE1qGCuclNkOQqCh
MVEwt3dpKSXw6wLQeeSsL8Yydh6k4HcMtjA0D/HpKyThQgwXWrJGyBsz/NAJ28o1Xqpp8doZBMdf
5yTHIRv0mwruKzdf0WhEeaZeZ+zxYp5aMeifh4QXPaJMqzRNS96Qz/7EdMFzJaj5rYZnv0POfUcR
r9i+ttLYAB0n2/ecUbg+wiXXYxQIbuhSFVg/iAbWy7YTJv+c7S8F5MYm2h5JJ9K9LGiB6CONmifm
HXz7D/5TU5sye8CZQr9EL5YqUObHHjsNqbad8576i6fU/88RW/O2ThYDOPwlNASCdDsdZne5R7gT
AzLoy3x7TReDFiV2VkUNe8ggUsHtDIvF0zAUEj+drz58awbNeVFgehgnD4TF4YqterLObekFkguP
0qihy/9CQfYm3HTa60zMwNGOmYH38GxL4snbZ5pvp5q7hQDVcP7chFw97TZkc4hF7fFBpHHcNyM/
njp4gk6KbxlNAuyEUZJqNgC1Pm5qSDtVhi0RS2jlTG62AZZStAbES34zQ5ZC3CYljOY3AM5lKyjM
i6/h0Tc0NtZrH1izZTnsz3Y9WQGdYohtP8gcjEV8CdIF7/h/AqewAOB59HVo/ZRnMi4kLR6KrugG
yddh3iprovH6f4v5rmKgOJmOUatS6pdaiJ4DmD/nZynRH0iEWCw83XXzCZ+OKI0099D6kVEsRoAX
GJerbEpBVe2nIIBclUmSiHmPejiaeUOYeN0elzuflwpwIBU/KRmKv8JLAqSt5L9BIj39RylMKnn8
WCL4tnWz2DTHR3Qo7P8tFlKNybCYuY7BGkBjGetqhwFl4wfQH7yXwXFz+NH0vbBNzfL8imTZlbDS
45CcwK7Q8SnfjuE7YQpxZ820+VtzWtFHXux4Bevxb0cKSD4DkTv57lbG6+REStiOY4O4Yjosdrt6
QiGEEem5tqd3H0hFfWkyUrJt0zCd3CweB1Gcw20JgIyEMzgYh2Fo5EKXqBMzBuLX2MkN7SwzzCHF
QPp0okbe5Svxqp056DU2avtnT5tBdNfA/GXSnVjCIPn/0iwBwJ+afnIk9HAgBuBbq+D8sy11ymks
7GiICp0XcfQdj+B90dj6wWQ56m1svGOrm7Cd+/WFAmX1emxq5gfwtoI+Qrk23nteIMI8hE+jCOHC
csh93lKsxKMqjRrcL8wGfa+XMAyDpNRX3UUrWygJT+izMYhiAYLqg8/2fHEgj8GgXn5efPApYUh7
rexGVF5C1bFtjAS407D+zQMZdHzd4lF+c25Qq7V+RTeQUcOYGhxLOdQ+p0vEcknsGfGt4WO8m5z2
m4GR27Zn/b9Mnb92FXlxxb11PFvbinJwryE3Sh+8mirDrwKxJtTGl706YWQSoVNuFw7AgNNpjdpf
zIKF2nJTkH1vJW0/h3r4TC9+uEkQbjz53XYL5a+whkL0wpBXvNT4Z2ay7WFckUAdxMT1avgzLBm+
eoZosNzHn9Y+nRtr5gszYgH9i3vXHt4kcD17BwbJfZLzvz/6u7ERLLuhXw1/JWI1DvHcfWIrdBCS
Bp4Urk38gclfby4SVaIK99YO1StOzMW3ZhqRuprlXd7QIqHFI8QOWGC5fdqE1yWEJkmoFU67xTNC
w9y9gzjvdb96kN0ROIATqNHWqEgkcOD1iDcoZcUMuZGFiodzsnNZx4BpDe8CDs/UZY0z9dumOhB1
GbRImu0NEoO3J5zExjUxgtg/Q86al1ggYXNjS6JBqDBmHTVT218Rsz1ee01VWwj2A4YQiINRfxBJ
AfM3CyeW3Hb/BCoG6gOxJDbctH/JkxhGcKCStSxmKSiOWQbe+bZrQ3LvP5e6GrrOSrl1HFf2kRkf
nNktYv5TZPrenU18Ni/hO/mzeTbGIHO/0xTtiATrHlk8wq6sLzpgSR2NQxUSvr/NF9Gl1cV5aYnq
qFdWTnePwspWYEMBR7T4KswAPFTkwQGkBJaOny7Bkz3sb3xyJm2OBtvMoElJ/17y9VhOD45BGasQ
vUDCPl5LAk4IJR97ZmxXOsKAqp3J7O45YZgsrc8TGx96tLZoLlvSJsQu7BrgyCA9gRNNh5PU8/Tf
G1d4X76Z0E8qmUvMN6TH463l0ldbmM4MXLiAELwzGqrqgxCQu8q4VKOHa2cD6BHj7YxziCLel7Yt
I7xlOD+p8ELhQc/JCa4gdpNqQslONiZJVp1gMGz9YI7V7StbZtlVHPZDYiOYFrIsREFcKSjGd3wE
BdBP/DA+MGiK2INsOR9Frwi0yS6w674wUsIYh4kXv4mj7XANUh1E6o50SRaZ9la/9pvS4G2X5itV
d9ebA4KnhbgBa3EMZMqVx4+JeEnoJI0LwMNLaDrHr1a4EAaVICT4pOV8BiDaSfYBY3hU3ZMnmlB8
ZN+S9Ix4fJrx0JBZlm8pTnjPquA+bJEWeHubiINKPnnKIJoidBEg8YuZIzjNElAagGN2db/0REI1
fBkf032ZD0ml7a0MnNbJwCbMcieQZweUB4vKVpUdsUxEsT4/X4AvA6OXLxD2LMxMA1R6JJx/Uu4h
Rb1JYaF/6cVroRyCU9kz6Z77mANZc3S5D3vNFIi+RnnFvDVW4aR6K9djrRwpsMLsFOURhVCrxiu+
L7MKr4in7y5Fx+sO+XMTVRqCzPWFojaX26NhpJAuilPjDGBD4vd1uha/O0pWY2nqTv9Wi58mKirb
nHSOam0UHA6TM/Yczh9+B/fdceqYScNvwoI+RBNc61nTOLQoirT0eQmvopDfr8L/XElwQETaxVsO
G8/EaBDeraV+pAi4LUONBwI2geF8IayyllTv32kByBt/49udIHTLYGG192I4akBRisbm4FVAIRwy
mhtSeiX/YZ87rv7dhBWMIgG2uvLOfOcIRP3mcDWnNBX0X7VA7shBpNfO1HZkeoNZjkzAwS9oXnYl
+r3V923qBptxpUJk4bRwtc2AiVdgNiVrKQbYpUvI1tXU9j0Kq6khA50yORE3OYSDfFqsGPpOjwwz
2yTGBC2pcK0KrNoeaORdLALlQE8TxGzyAX1c0VjZ0Rre1cNWPBuMeIfFKxm82KmPmHoBbCOqUsnX
rz7Mhp5edMuSo7QnMCLTMBVuU/3G9cU8k+ZeAKg8P5du5H+rcfkii7evJML5SQKfpQaMZN8vv/qO
sXakqrakvfCuUaeTvaD9LQeyJfPKmqyPq5TK/hfsLeCoZa3rYEiuyvhARwhSY4uxFr7h3A3Q9V5Q
SwcXaTPGhKZDi3tlABPjkktJYAnd31vWm+aQR75BEGVOVMmQnmRzsJGy9EgJfe4Fj+MJo7S0JL11
f7Y0dbejL2m+1lbQNmPJemIxyianSmU/+hGN9sFQYDfeXbufP0fy0PtbkvO5U/NaDYz8iP84b06D
RCkBiUGWD4oCnIW7DvK9urJ850ZnWmrOCavOiB4fkVZ1rsBW3qFpdD7m66iZvhYfJ2joKQoveUID
+NU8CfnRt6mNPM1DsDLiJ0wu3IR+A4jYaXwFNoBkml3ePoGDPJs0BKHYdOEtGkXGikUqieGXA609
etgiQLoURFkUJL+w5x3t525OlUou4VS4RByHejkofnRI5lpuN+H+ZjiiQDKo7q9+rwLcKVD7o55X
kUkbHhBy2R0dwNoTzVhZp8zA4tXaG++OaPzU//GTBB9Fev2Z+EBg5sUrEarAeStVAcb5C70j44SP
iqBFOhKh+Vt4fHncW4CpbmJBrNLrpn/nwopXV7p4g1b6qlRJc4OWiH342UBTO28OyKua6cgdf/AY
g+/agvwSPeFXQNVb35YjlY4WgwVEM5dEy94QaHsnXOVzDFMJWoLv0J+1CuzgCxdJ8m/8XVqFB69q
IV2zfXXpAcmMM1dOFRIr63bvyASbYC+yWIBi7jGYP6SaRujc3Aq39MywPK3pkArvtj+JkXyPovLC
o2Yu3uhmbUSlCxsNHe0bLN3EkVT9h9uT6whrQmfv2/NxTUxMCPFyUBzsp5RCsSu+gyplrq/JWmYV
jD16G2EnvG/CwrBpRJ3T2XXEBl7PmxB46Azh1H11M4o1IvklTRCyOIxbtZc3QxQcdTs/0uIFQH1C
ejDItoo+FV5HXo0gfYWoSbiKH1rgxll+Mu2lhW7rf49JIaR6RqaZTR0OgwAOnxy9DJnITV+jrC/N
itT5VmUDB55QFLyCXfv0x0TGLZJqpo+mznK/4+WfkuYHS7SJxCiimPFs0QL/N1jJYVscBh3LEdf3
/wFCzPJvSbDHTMCqHA0EEYLCEoCDb7NYuv90odYNpI3b7agn6uuULPSGcm1FeuNV2yodTbwzBfwv
4HniDW4y+AoHaVxGmJxo21MVtBrPXKpZiM8nHUTJ39ANAvBkINwrPd3jt8VFMndPP+xwLcjYSLA6
P5l0J/7sn3wO2cg9EIy714SfTHk+x8Rmf+l8XeCpOfI2iHdEwxmaIEdQLf70JYtslfr4+wNNslPT
wb+sJs7O1tECEruEyK9aT1mSclFFJl9xPgMSo9iMS3TNVffGhbuXzXMtO9+ZtViTMc89bzHZUwiy
Qw+Il8ypVer82Y/1VGrzkxGLJUEkprVX6cJoIO9yQrltw+lZSyNvhpIRnK6UsHiMX8fhbRmW05Al
eSf484O8OxiTk9tOmYPkPmssQgLVbweXE6h5L1wEaPCZv99RAWW18DIhE77iJI2EouPnEodoc16M
kcBCHeGakzDoXNgtOQxH2I3VMYhjnmnoWO6dMF406l2KQvBtn7w9W9CibbQlFrMTFAX3MThpPwMk
enoQJyxdhgDPZDrJ7LS5c6vTe8Li7eWR7v1P62usgHnrtw7sULjjN7feClLIaiukGohhLeVUdCWo
nXu9Dmt/rKxItL4Ip6RJGusGF31FaCO3zuCKBuluImdfoHT6G/GUNRUL/IVdihEzrYou7+nzE0jt
5rrCMzISjBHopGaPnpielRzItf4QVnV5HjHvLf7VsbLeNUBhXre9wwAGQqlSRatnA/VmCW9SRwE+
g+Zgu8mdf0sIkFhm5a1Vx//YnKw3UNbjM/aXsfndrwUuf3OHS5GUdNtbmZWfIN4D/mnZxalaM+e1
vUjfrVdU3PAuFG4MDTDUVHvuaVfUmqOa+JrS8RqWLy4AvR4DMz4HOnO+A8rymoSBvKIQQ0bMzxCk
m9DKspNb8S1UYj3o3YOvimdNjObMyBa0fDrBIaKE4JS7CLyncCH2Fcb4dY5GsA84vL8kvyHmWlJZ
M9FGQNpQ8KfWHIn1hGxQJBIpEBQfzJZKcl2ZugPIGmh1BPpSI4yYv9A0I/rXQRSvcj6wrFGwW1nk
tKlLGfGYbm1Gmt5iHohm6kyCdg6XDV/lZbZMKdO3+UstQYVBITNHjkpUJS3WVyGQ7Pw5T6Xnn7Wo
vakfrjjKkul+OtGNNJOH4O2ouxc9Ty9/1xNFGjRPmVKfefsmd0oblY7uS6ALy3dCTkEW5LZ5SdlB
sYPD4LsCNWtmGQGfa3Fg/L2d8/6uPVxklzQ0X7AYSrx5W/Zza9JHek6HhS3xlGSL01LZ12MlaqG6
PZh38vqoAt8JI83SulkBFbBYchSi4sVo5mp4fEyyuVzgq0X/2VK6g0QthctSBpr6HRmUbOl63axc
vWtxCqpPTxpwvV625ahJeXeN9d7XJO4RWBVf1BwI4ifIlew5jblm89zXukiYdCQBX9JbA+3F8Rwm
c2NywPgpOc0+220ly0JkSSH37409Dj1/V0JEj5hYaH+8GvZ7wjD6DkBlD93UY/viW1I4zEQsH1tu
vFoynIWYVEX3dhSoNQiQj2pQEnq6J1KWIvJzxgh8JJeGR+wcbvZGYwNYZptiwjehbczyCWVIzvcF
P+mBrgwlM8lpdKdtJ3/wphU57+AltLiD36KfpvDV1LyQt6kwOi7bZbVYzU+Af/LxaBfavVodGQFO
yYvRpTTFKwqv1seZ9neUBQGJoiCDPsEUsfVu6+tUru2rh4fnWbGhPn450USPSO4+xk0yGbN9h8gr
2YXPB7i+zonn0pe15GSUlIMezJqKrO5Km4oyqYclIzV1qoKvdoOLzcJhN6ZQA1c4EzzcY0hrK8BN
Fkbu5Ekb4gqyj6Jt3aBcPXdHdWXdJ8w4kI7hJjesLLdqV4Wi//3/1r45AbAt5x0kha/GiTn7sCQF
GUIqlQagFyOWrHLQ0xCPcrXGUZpXYYR7JjNMAV9Poxop9+v4Lsat3489InFtaQOIa5HTHZNOfeMd
7XcPbiT00TCejcn7u3puh7r5xWkEtaF0BQwHUECdGiNh6MeichQq3t+vzTUJlnR13vHLay6zbcbJ
rAYTUx6ipGqF+QEMVnDNt2Q9UsNFdb52v0jFADUVL5I0dYZRwSwoqp8fyfWPg7Ma4aHoX52v2M3q
GKCUYNKErvxoqOnA14xlQf1yyxcTLhR8IbKXx+eF6NRN2d5/PN/TjCCXvrc4C9k882UWP7fbw9Tw
IRTa++HhYPCFumZHOb5+6ZcseOQ+AxZn4C1u8PylD7ki5UBAWK08IO05njEFWPEXSYbUveefhMFM
hZk6ruqlBZBG6WFd53yWula3y+3X0gazZ7MEPdUgACzgTir08zMSJcJL9Oo9VowGMpaCVVe3oLHt
Rb7/5C6hHrS8Qaqwa9Rh/a8POJAS+BWiBOHR0mtxLg2FYNx0ZolU6qHChLWur6nilXc5/EFB9yHf
Kq+uRbD5YT1WJMopIGFv5sq2D2mnAXiReEL/toOw6+t3kh/3UNmjo8ZBusLj/IOVbfs0pvsNgKl+
F78d5lLwEKpRNtbQ5hy06hzijyq9OpFyzeLrniJ1vHQ3u0m8vv7UILEYz3H5R+GdCiJsagBowu4X
WPpSC6/SLfH9VtShDB/elrmgsKUIKxgeLv/zhVfzQBJ3y7jcRIOGUDG2P7Hg7vYbnKANzuDAQvRm
tUiWprAkzst+5dWpSnoLtk5QymOD4R9kJFTBeY8om//8jkxGStuYY0N7U8tp3VgpkPsXSq+m0ZBK
YktD4lyjS33WwnlsrqQWBnHFVXURS6SLLSqe4TPstZQIfpnojtlsjgqMsnIL/QWh/IcxOiphz7On
YpVgV3A97HAdzNou2ergHlw3E/1JuI1tVtJBGS1J+dP4Vs3f7J0FmOydi25/r+cSc5/FjGfnquhs
CMjIjTDFNg03UMMH/kXhySv4Tgcd/sTP1PloirOlcjm0B3wHpw6g/h6JFKLFaHu3Og3eHS7HO3fS
sH/zwij3JtR9HeoqehJs7suUsky7tOKBmbH5CymMigD6iF+c55ffOhskXZ3gl46jZ01gEUX5Z1lF
OBdqn6f4W3f7pvEDEt38B1J/ZXAQ6tnn1cofYMyNd+qw8XghHjjlyfXUq/E6aVJuVEdY3YVnlz8i
ucfZmGWxU3gclgbWCUlZVq/0yzgndYUjrbf7j9jl6deo1yVjjLvkb0EycSbTDHKiJjlIDbyMHO83
4M0ZhT7rZNlShs1fKsL5YMsqopMo4f/JKCGcKdyqC1gvA17NCbS70uAuTliNinyfNnA+gygRnImx
EkYVKDHZS9cHpKRRsPwXT4TwwAM5qkap4wdBOPNkERiskH/LVS7H7JFTTqoZFA0fjiz87GRnxZ5L
K2CUiQ1G3F/eHaN0KUeueUXZCnhzMTUP6jhgZ/t5BjPaKRhUy3Wf1zlsT5ZlQOwmh+1iAWqtetyF
oQx82KA2GXxFOCdzMkuaYsMuwHmqlUZe9iKJpzgBHercZDwho74cQiJ9TpqeoDVfze1uSyFApAh2
fTeF+rd689rGTlNkzwTZ5y1vcocLP3qJmPbBb6Z+xrXBUyaUD/kQLTCD7wrSQa7JNe6dFSjNusUj
TFfnD8LYq228DiZU3ldkchHbzgbGzUd/+/kemm81s7VGJDR8r4uHys+l0faqPfmtHoXPzy/n0fk5
j3h/4KRYh/iVEy+8+LooWfpnopAl0q1LglIeYigUdshACxSB9wtuu5nYBIOwzW1eTtVCHGGTBJ69
mW5Ml786OtUHTIWJ/uiSjp9JN/+O9ohnrey0Hm56lu7YcYBcX/UBU0hyhmb0ppcrlcbwIYTswxKn
OFvbX3xuijWcF7kHaf/xR7XwY3RwC1s4td7iolq8diIgSvuKHwwRkx9SECdhlk4BCR6FCl/9Tu8b
XaxDRYm+E8ua9X/Pv8TGaxj/6j3o4MhwD+VZ+6t5fER3Bwpzbp2XeemK/7Vagr9VhO4p4UszVR6i
MePAaao2SbotRIGr8ZgnskVn2l33hbQR8HO/hQX6GJW1bwuo4r0NCW+Ht0ll7euFffyQWrEz8bB1
/JFBZLXXfc+wEZYMEQdcVEtD6qEGzPQyXC9k1sKPGBYa52XKe9xjVUMMgcBuN4wYKscxPD96qNTL
NwmtQZrP1PwSmH7XicPVdmXvXCProkduAeTOhhwB/TycVdCIk6x5B7x0VXzrB0OBunYlhtq//UIY
QFM1LMl4UhN0BsOcs94lrcGb+pZXMvLpPe1r9HIvzmqisLs/dIYFjozYLEXpbOIXGYJ+193UtY0l
juhRBavA4ND8nDbO5tv39/JEz2Xe1frph8iZC+DbTqGTp/EYJjWZU5sNfwMbe6BaTKZNzozIyq5f
eFcFAk0rxp8nfrbGGrkjDfzpLpxd97/9zJaRQLT76mkSXHOGFc/JNbidx1SOvBdoXmsGcj31rpR7
asP5B8kWFMZVvGnENDB9yQ12M4NY0eQof3/pXSaGSZCz1sf8+244VUWCMyNkWtgAO7sPiAB8CLdl
ejw2hlhbWRc8paBGAsPUF4FZ++35+lzgu7A1iAgoMBWTzWc0f4CyQlaBedrKD/jaAIR+C7ltJE12
66Mx8tnyTIqM8NxNETBu4aZFrdH6uZYgA9jYMcaUj6KwEA8vlPTtk3DfdVOqgSyGQXkvymCZqMxb
ASqy/EZh8AD/5bE0dUm3tcoQ4pHaW5imh1vWnTaBjjbYRd1Rn0p326uckBxuJxn+yXrC07C9d/7p
hczvVNUywTiGC0ngAuiNl63pKTY5EWdVlKfpNnmsVrjNSoprm5npINY2ubs1m++xFlQtOpyejfKe
Xfl/qIgCNZj6Y4LtPQ13rRAhNLEOmjH0r4ifono8pYUVKXvSUU1aEtug0Crj380dCTrqeKFMWLjp
nMLB3/tufLE3jRxOK931GWce6DFJIft2+d7d5L76B8VUm6nt/zg8QDBUe1iQISzEFTxRdfajNfaC
nbk5mj0gGv/kQeLcXxd/Lo1flagO8bhrUzGMKR2t7hJtgLao6gaBdG7PbOLFGQadHJHro2bb4jrh
Z8vq32o9HKCaDqRW5I9sJRU9m7+dUXnhIFS9+ze5TgErIsmOBpHNPYegcCDWnrT1sq6EBRkCsC2w
xuHKBdIEZ3xz9ZW23yD7FPZPRWqV9ylKii4YB0dSjfvg/7WSvQlnGf/xqWY1ssuOhvPzpZpExuXU
ZUwlmw32NAIxEnzeJgdacKB1EtYuQIvnj+6QMC8DvG2VSPzDwZvGSb0YIUoiNVXiKUVgudqOD4Se
uUvvVd2+HcXnyVIuLn2mJgDn9J0cgdWSAu0Cg3uTQlhSLOhJ3bH3Ge/W7JaBFVoBGCSg/+OSteca
HeMXE74d+/NHd6pCDFlAqczUMzyyFVHi+EBQb5eRnESFmNoMq42C3nR5KZaTAGm/R1WTv/WHiCAq
Vj2uO5Zi7sI1pIppzUn96FTiiCBvs1hIIlxympHk96Ne5dD6+Kp/r6xk5+6ooUfLj0DqZ1Ho+Po/
PJWVuzZ4mZomz33GTuvzoC3g7twX3Guk8XU2j30sCVY696AqUocLPdfEEdUxO1s1rhw2cCKzD1pC
FPP4azMSiynYUlRtr8Wu2V+tTbl7y3Pq3FXTtRsCEY+UqZbTgzhhOFbi4HccNkgrxXXEKOtlRK2i
/KOkn9K4uBF3to5/qTHmbJxlEOFp2DD2MvGirB2ZdBmRntqo4C0s7dyZrvKIHqyHE3T98fuaYJxP
MOJhsgRyMQF3q/u50pBwn2WpZzIo8KTk/9uhnFDvCOO1pIt4nZeZvE2XyqYDZn4NyN9peKGT5Omv
UhcRGTs3Djom8DMZdulXPdN3pvsBIf0o7ELOv91ywZNv+/olozOQMtB1VyzGo1p2yPuNjGBxU9tC
XyRrurc8Gz/LugxuSEEw7X8lJu/u6TrhUNDSKUX9yX4cr1xCODCxADUcCh0uoGO1f83F3063Q0iK
xDDUj51wNcATMAclSJOLT4aNe3w3sfYfmjCdGKXTaQ4GhR+x6xb1IVSuBWtV0wYmLv3B7Xuw3hOQ
OrxPxs40DAneT+8ZttAnC/f6gGOmO5NS/xtzZMXPapMIXb3LpR7WOT5vsuN1Dwdg4sybaSlfmrxU
txrqjPEdO+NxQChHiY+RkG/soOXmjBZSqJ+G+5/wR6ZS6KwjU/cG4HQnvSaKhuyDsk3rz799NS/s
8Y4PsDOgIfL2CuPxPdRlAHNwsELgW9qZDi8owXh9ZZSU+W1g/QJbelKU4gN5NDDCEXjWkfzVawUV
BMfd/9nCBj/WDVPm2xj1o1WFeVkTus4gATnOGwu0aQEC/YrmhC3yYur1WUElV6f2EbAR3yhCJIzq
kGtuU5nSgHhLlUwS27ET9XYOLDwvj/r3K1efoACpLgiQPC5PghrUB5k5/Em/gKzuo4HWMVnviqsI
mJTDKaQSXY1ZwhQao6TPZhuoXvIPnhsIEb1FCSlgIijypLdtR/KUXTBfCsJxYxnO2FEUFcrhwwh1
o7lu3rtUhyMsHZmKgpPLIQCuAlDob/GTRpFe6icuKw98T1jPN6N63FP4GHlJPFIMbJbhrDGBYWII
NmUo8ygob7ongtPadk+kklTaIyiXkHCO9i2vtbwD0nM23IpDqcnZwJQZMgLEmlaF9WRCZsdxC1RD
hIDJ0rM9L7vn1dhUKCUIQrFw5jEkUD7irYv9reKP8mHOm1SA/9WhUhssux7LvwC1GvLjCyHIzejZ
3kDqCCSYNsT4HAI6WhI2zuP1jqB3yfoCYR8EuKLqiYxgsfj1A0nem62NIHcUJW1uMCnxqWTpCY2i
PrnhjRAbsJWicR7uAXu3TMhql1bMsqMWV9kt54/sqFf1MlGWMHmfg0LPf4UeHsNupaxY4avqPM23
22o8oGIASAEME9rcoaAGKO/Yh2eU7r5RiigG63gp5z+w0Y70zS0fUEIbDi+cWRQRsIdCwOWT4hlz
7PLkpOlbKeD81JEg8A0p+xg3syO7Wq8tToFxiGZDqM7p8OGx67xQ1MJe3+bQIuMsFiw/zvK2Ugjg
XpyTwsPPrU7gSVGCrpqhTNR8m6k6gmzBwvO2H1SE/6Av1J/gmLbLnAbAfo5vXmBRDHtsUvG93nib
5WXZg6D3rYQv5mNfy9DK/234t0q9X44lCfJfc5TlXLkpMf2dRe3QtZPBD428yq0J1fA2B4oqNfz2
oobenOJ8klPb4xJ74NQ02LCDkcurtLyde/xyfr8uU4btDLXrl5fjSfCVphrB2Y76y8p5j8dpri07
Bziw0qmpnvEdm1nUxG31u1dZckzgE3hDLFql12N1Gpgbe7+utRPUWAJBWPcniPPKMutwvcz7mXOh
5ZiN118GcBGZoBlZ4T9lSxBMol725sFkvrqISC72ti3SyjUXXe9/VgSdvhCks4QkHK9MCVOlkWhz
qYixNrW7MdU6GhGBZ/xBKiC8LsMc/CKjRTa+gKZApkTCE+bHRC7hWnsu8rL3o5NRY+//uUbcxGK8
1ihMzxPsG7NbyIDeLolDfN+DLrGX+xIUE+NO6yoIjLnRvlQsNHXfZyyWbuFQF8KmVaCgM/Juhypn
/ZPElbX8dg/OMPPM/cO7mkKsPNfRwEJuRTBrBiwqz2l3SqFZWjcNU9P7GmwOzqiiL1sVXtxxRFO5
S4zNbLo1TR2eOoM0NvO8sLr82pcZ50tFfqVYhQ3fqTs58IjjBWd5aN548GybHjYPMAbFysYAj4DF
1B83BQOdLIUQlx9s7Vk+8VQzCgDJVFeafvAhDWe0ZsXyuijgfZIlbzsZ1Rv2Oe3OjuBtHtmTk0oa
YFIwjNWMT49Q323iDs2ZO2DyDyBgnLKb4/ypj2uqm+LqY69wG/JpfQ7Yr2EOyfdBqLMer0NBZSqa
LrhHezAjNyn21AAgxreP82NmiB9jDXBzPPI6lIv+huksVPPipJ6qckv2ZzaakUJp+A/zN/YpE05T
ovMUmGiY7MJAqeoMPxBNl8CHhNvRYodU2c7SKooZvRZqb0monddJd22NSYlI80P6h9tqHlB4UcP3
JdNLxO7wuNDMo7y/NuMF7JuGK3Qpa7nLADMvvkMR8MtynpDJwx4Pi8nfmMeVtykkIvOcMj9T19Bn
TwKu83EJCOR7OY4Lkp7gLaBvwbQvkmsZxafXoGkeWyu7/0LwqUbRVVBaR7trp/FFkPvHkyq5sB/a
ZgndPbBmo/HSqk1e/4Rf+9FKXvE2n/ejGPtcbyoU5B1kPJa8GOny5ZGC+TZLTMpSbW8i43Gr7AGT
3yN6nrMhGfOIbKGsX4y3JCjVqqbBf9Sa83KZMQyF1DvrIk/I/wtt62BCHG/U0CoZbNmV8gujyjlg
eJ/HQtMzifm424dtI6D8LJa6a7w22jijaGPbH20tkBo+89b7FRGlTcO549jvI+6pktwUNkeWr7Er
tJILAvK39fBk26TjUj+/jG7goWRop54KeBQl87TJ0WJ/3vXm99AjxNB964vELS6eMLaCG4EEGLqJ
gcZCaY5Ib2jTF/ZkTmaMhN6MULdcTn6hxQSkM+w0u8zzysWvIlVw5/veLeNy5nQDeaD0kuYtDf+N
rOcBxsEdSve+1ARuuBCOBFJcnqVVCKxUSuA6yQ7e+d6xdmCk6723KSlkv3HKVAOZAe8n/JtMYalM
Fh4kqq0IzibodlVy5Q083zJlK2s/PVDezap9sU8HsgbyD7OMZgOvUf28E6L7Ej/FRnJIq3o/c8Ud
jfEXKA7HJtQ0vYMD62V1k3xPiWPYZwT/6I3t+ax6uFnxnqnwpe9eSl1ANBbybitqYAE8tKdSmFN2
UNwmApkUXCnUJ3JSyXQJjziMVK4Cguppq7iyki6rz2j2U7cgJe1SPdfI/2khXiL9qVNfniSxCweL
79xyIhERaQ/XfpKWEhbAaNF4MyG/jJ8gcFUW6Cuj/k/bNZWW//QMZYt3pgzPpjcR8eRcNyTwjAk9
QADZf3/Yt+bt5RvJMPgJ9a4Tdd0s/A14B3DTeOJ4BBc2C8ZfY8hR5ilRXodx5kJHSr1uKLKDa8NG
orW9o7fbmg7v311r0cWpI+1XE324gn+pC6NOEImJo6oTqWRjp3h51p93+laG9mg6sUos6+nczgv2
TJM+AEiEHtURm++MiloyeDZ5ajwGZJ5YRLM3IXXdV45YOvM03oK7udCOckm8sMstDpZTu0pRH6ho
JgnCJB+jB7j4gvqMW9pipI3KS4CiTq7ebTnqNX9aAOHlHd8VDb0qIBrrXHXEwt3CfClWHz+zdBXd
wlcoV8KkjfcmNrOdGqbQRr1k4Jq0i+O7OMjs6Qj8cWEBiuOq/rnfpb034mT7Sb05EF2yeK282tAF
9aqSuXOw1GtZKft9RUJFKYug7VpkCMLCPk3UNVB4g91ogIKsnLWvuETXzte3APJUM4IkTH+txSsh
7H95iBF3CquX0kQOKnNgT7tYK7UMpzKfJ8jZSlNMCuokzxNk0PtseOE9xevtXoZcJORFMA9VLCBR
VMEX9ZbQMSiX3yq1YjjyPbfRT69M2YE5wvpo6ns3xoveVIdiMl46uLrSPCFvo94jNq5SK0I6NTYB
pyOi0vZXI3OIA6wv6nilsBSdL/PlJoPUwqeJ5kPpH9XwSX7C7NNxIv62JHGqDUewHbcXJPpVEw5V
pw631pKyt2f24NqrtQTCAc0tyUXIH0HFE0AlRf6HxoL5Tfg22bZY/OOitl993cze5+P4d12uDCCx
e0rGSL8coQyWT9pBp19SErBbCHWHfMrqim4rVqWugRNR6xel27OzLIAtk7GY0RiBT9w8LVgwuGLB
gD6d04QlP6iChtTICOkfFUJgmDyLxI1il6c0ye4t6PxJbRtPi2n/5nGQtEtnKZUh+VPiFcYUiy+Y
V40Ilp4EsvXCDNM8ZAc7QKMXjueLDI5evLUmH9bxcq2LdkqMoAAm3jUxSYCFKWp3nI7+i1XLdRFw
zKcZnLghoo+2HFI72V6IOMJfVB0a2KTzjhdkPrv4UkfEk0NoFpGOmxv1pEsbEafivjqFiavvUT0w
UmrGlSBKs4VQ55EAZt75CBgXXEWc6HsFup5j4dtKCTxBWriLpYmMwWDpEG7KWeyy9PQ7eP6hyVfs
rnR2FKuEC0Y6Mstxqt6LvFP005O1JGPuroPut2KWSaLMEr4HF4OEHHOABTSeDShRqxYpWm+0TfYj
KUEmTZ3JBqcEPhdzxaMkoIdSM3mpFl9096lxj0h5gLX5ilh28NYq5rlZblY4F7nvynT/jFexXMjW
Fh1pyYQEfQos0fcW6yODYK33Btco31MCbRyHcoMfEC/R8jwVyOHBXc7kYDwup1WgDFGj42NeAI/w
kDS83DXXRX35LFmaerbfe9mghIptSsnHYvb2ISdcrV65/jUSP41pnARl8M28dVFy6AxF+0uGA0+9
1UY8IckXhhKapibVzP+VbIKeTKUOGVjkLpi0oTKbgta9HJsQR5M6nFYxKNqcl82nWuf1NJI22NNU
PYRMN1pcFhW1Et4REN3xjgNHaahkLL+/3lOJPqb+dO5V6if4+im0FZJDa98n5uFRWGjgS0k9aGEW
9Z+F7P9lwcqjLSXTcI4Bf93t6E8rT6GV/Pn1cEusPBBNZWbFQkFhnycXkiDhSdpP7VSiXEwJsBJ5
Irpxj73CczI1CNgzNJawZiCmHQ5pACfnn2AEglv0Qm2eAGo+h9FKLY26uLAlvXRB5WP3wxiX6JWk
f+rC5Dc5GON9XK9vUAUSkUooVmfS5kt85DoiKo90fuQYc0pPDTx9hqQ78hY7NADdhJ+ToX4M2ONm
jxa6d15HMFRpw28GX4xxNMu0hW7B1mQLxy/f/SFq07J7GVe22A57ZYSQUstKTcw8FrVkDy1y/UO6
vt61S5kx3aGk/8sBnvraCS71fx9DDl5H+rjIam+E9edEiuFDag/ZqLTf127vQ6X9Jo43YconJmod
UFR6J5Ca8LgrZZouIi5Xjyy1mvjqrL1jFczkkR9jM0G+/PcgUrDe46gTaef8nLiMDH/F1ugQ9W7h
YYSneiP0vMp+xfQ16eshg54QWyfKMmwBk1uK4tuYi2eyNhGV/C84tiKDRbHshlLwfqjqIaYV/hZ6
lKvLNjkrP0itTQ0/IkPtvZY27AyzzUpcRYo0KA+/R5bEdef+u6xvycnRj3wTSHEftlcjEa73Hruz
1RwIfG9rxjlsyFdpHsMSs1XQ8GnadCV0m/4j1UA+xHayd//KcxgMZY4gEmyHVS/HSms5RRX3/xlp
n1Q1g1mq7pb5vpwylGDc20CzdL1IicdDoaJXYsj/+kEvF9z3LYujicqVgYk/q5XznoRVKavrf/V3
CtIlpJsY3nCe4e5F3ifeVhkahEKnjWgcrRb3PBYTnyvp9iL19jcwQa25vlqPHWHfs39AYqyK8f9I
PEyczHQkIviB4y3Ah48G5+kYAhuBz2tHODTAIxSEn9qyeupB+dLNag9fswzrQ+cPYEDBSaKYTRxQ
S/gUyUXYFhBD87L+i9mqRUG+U/ez6HNHF5/Y5FDgEz+ACgDMPIIRJZn6copR2nOZzcT9o/iP1otg
hAimpS51QPRMMsiaHjMKSRrxt/fBv57vwZ9zcoeZzbvXOXR8kzj/+01XyjJ1F/+bL9V2IQjrTC/I
z8ddsXHQBQhXi5ADSd8fDGnfR71QJJ5kBwY+nhucuuxxjsRS5uUsfi8gZk7Tr4oD+HccftUU5uYP
MO3crpmL5dcllykyX2loSCc7vVg5rDxqkVRosIMmEgn0+3CePz70Ki9CYnqUQ0aK9OaHNd0WBttV
BtJuLLWDAH0fzLIpC6wcLKIcA6KO5UH64m/3xwsZy7s9LjWylV+CL+OpMsX75+UHFeOv53dB+KBH
JU5ZWavQf3eey4RJL562C5Tmn4qHHqbHdy+T4I9XPm3LFZN9whEfDZ5HQbt4mDYY2tnO2QAGflFc
zwuzBCHExmXO8egPC1Li7zy8Yao1OQnEA+g2zPvRU+echiyx2uf/Rms41982H2Mi26oH4RNTk4QX
FFTSej49vF9d5vwdteH1XQwmgi+Wr6uTza7Fw/ukQrZ7bdM610VU/u9VVaBZV4y+j69d2GVnhSX3
jvaGe2U90FKTWpw53UMlgJxve2MC1X7Pm2Y79fSZV4gYoLoyBeTMKcBHrWlukYimWZxY5hhJM6uG
fCAaViU3h+5rlkPUWAFN1BZNwHei2RcqFWTlECsDevkf2A+qNHzA79TvggSC5ZypHNoZTAfV9p0r
TWjO+nnumDv0I7GoAgkQVTpkZEvLuwRpVmAGQIJDJu5I57UwB5Xo/wKJUrVhqxignFKnovNIojD3
rFESmNbN8HaNTcuRT3slHFCpDR7YNkk2VXGkQcUpw2WdngXRfv0ZpMu9IJKkJLggy2ylBWddP59S
k727/0Yvc46I+D7SfD6pnG/3DrDp/yaHAUdn1PdAgCTqtrwtFYYPatzWYbrTV5VJRoC+kYxyPDSq
O6rtVKh+6rJkOB3/1i5XuES+4MXUo+zdRnOKzw5zjj/sjMNnTGaJey3mPOwmwUNHIpRVNDDC6Tsn
z2QI4OBRgK4e5zvABb9PJouGex2P6mUySRMRZzqd51p4i0JMpmZc3jpzyrnnpacKcd+8k7Yl6LsL
mwxi5EsNKS5x9E/Wns+qOpPZhI350XvxWmWQ9oteh2eRoIdgJnFy0CrXcUDI+n8UmYJzxuMNCXlu
H5dwAsfz3MldZKcTg2fXFtiviH+/Jb0tg0WbeCDr88fqwLJdoglYoZQNoV9CFwRTcWZcRk9qWLOS
/scf/GSOSR5xIymXemlhrGmkUuc1xvad8lA7Dz0iLmqWNSjJci4qYRSVosh4pe7slvyzUpb+QbJi
lJuUUckxoBOYnIb//dwj7Io+SobO0uCdCK19gs4CBudDGTcyXr9xI/BmvS95ZEgV0mqS2j6uPEmp
E7FT5VSdl4ESUarcHEISpBiHWFYebpmnr/vHOcUzDS/w9jNDOE2RYZWv5qGsuYIvW5acmA2/MbMY
mCP05LxOXkS71mdmbnL3dEAYbDw3GJocv2YXOpcCk4L5VwZl/oXX3IgFnWubBfWsxQ5tl8mGBZjh
LnACLvQmfivcwCAdc1NypuE5pdc4DduETLyGmlhoJIN4eYTrW2slq4Wtdp0NIR/ktpd9/M41st7o
rQSFUhWrllpVIBCPefLllrb4neZ8W2BiwikagwD8kI7ZN8pagvsLPllThakrkxICbtiNlq6wSNnX
LuYhi5oSuqYBdsHsboIs6ntHIbV3zY8vYNaD3/c4psWfTkppPktbKDCCoo804HCDvPYKvKsPsuKc
oIU6BIPG4/P2nsvQZiF74v/OYcE7Wqpdhv0XGdHg+DyzixVEumZdlAyNd1vlR0wZgQNjU6YMe4iH
0zU/dYH6b7675m0tE+mfUvAZVzepW0gbMULoTgEzRpyuQc3+FT1N6SCWOx700phbJhkiPx97PvOP
2rd766b4lfE+cC07Fi7Y78TKbHSMRyj9IJSL/7wwZZ7rrBqC/0tD94iA+SnV7aETAUMdLqblJ7I7
Uv0feqWA6LyVcg9+0y3ulghRV+b2hk4Yh0Ww5fwh1uKAORi+amXCzT++kMmI9NyYf/QhndFhxKWf
++JgFbLapwn9JCBhOZR9onU6OkHCncFOyNnEDJLloVV1wVlSkmOM5OhD+vQ8hRVBG1pXI3i5PWkA
Pyor40sqHS7z2uy1+0E8WE1JTmmSyroZ+1grEmjO/4iMmhlK8TNNL2sbove+QRjTSFeVwwME49m5
NUAMboVmeM5hWW1O9M0Ki1NK9lX/N1gTe5O/25U1x2icoMo1AJFjW5N2e1E/78qtyKdeKrpk4WUI
iHZevUNCQjSoo4941b3pufVE5ExNKgKE42gZEFaZsioEmhsB2FJPx2R7ZWPZSLUVdrVPtAPXIEXZ
r15FAY5MHzV+a1JA9CYZ5XPzF0kBQM0FanzbpgxfLhwRgWm7mDLjxzl4JvUxoTopowVknpoWDH9G
9hCRbhmzcjlHVhgVO2mtqnEd9/ZEV+rHNWC9Q0VMRSD+p2iJhKGzvRIJb7KFxX40cpMOq04+uC+z
/vaTyy0zKpP5oH0e3585/jI9JvLI5KokA5IP2mzdb/4v+w0+XWZsGDhoQNqQUM3OX8kN0/lpi2zO
3EPcVyo3j9TnjZrJ5sH2cieWbTSfdJYOQY6Qgir9f7yK0tLZQbpMW877Q/hmH60n1ssOXAdsqxYI
weB1ev+mLoZNIkodjGzG1DTMVbefUB1emNJmV1r7KEVMtjIqW0xKUgbjvRyivtBinj4y3AsbZ1T+
Udvz/CNfd/u4II71PAgBQgmG2UJNbufwUtuSEGOdKycqvoD5XQ7MIF0gwWR7ZxQQoceGqBAOf+fV
qMA3PDGZXfqMwAP679xc7U9iZArUtRuqWlvTb56goXCRf+JlR1oYpoUrThS6mpna7gmCKF176Rbk
oLiJe7GXPUOViWF61E01jHGP1wLxN1XQDWIA+P79PdL+dvEXz3L268x1onIrc7PhFTsXT72KD0Lw
QkAg7pL4c8+waHqwxzJOXLcZ0lCQBIXlBAkip/bvmSNvY1RL7KtRMWfaEBWyOKMx9UT4Oo5n6Pnk
+Fnl2uO6AwMMND126xmH+cyJnQX7hirRRV80PWDSqEjzLHqX/d6+BBnjkdswxdKC5TEJwd0oYJ2g
0Qw1jxxNiQaKKgaeOwNPkl70wBbYL4yGg24mtCq0x73C/21HO9xtNzzmbbUyPVuweMCdSKDaZn0c
q46M64vue62gHrQ++IcR4yiFcbDxNe7z77uZTEmJRjOBN6eBPQe2jOhIFGbhSYjub9HsCvKOxR5S
RxTxvsytvb8VSeguvFeejNwXg701dVdP7oJ8aInD2BqW3uPvrZPzQ6eD155/IyFKIW5IifhYz3yM
tM29fwawer7BH5I+RlMzJwJ+kx1FyqnSVog6YdA2qZOy3FkCK7S+n1Zb7S539vIvoz8WnXvtSFbL
2wpD7q1Ip6dwVPky7amQM7XM2oBq5XE7ysvatQc+HU6dETNA7a6tq9O6+jV3gz6WWG1rQ3aFP97k
UDuMYNQl02Fzi2ysiNlXJVw363DNKEAkhhTp6KjOSV4Q3Wt+Mc6nDGyTtsoyYc5ZzA6WoqFnQF9U
PSXERewtcHEqDmCh8Z6YlTFDG+/a83HckMPlBLvJJAVUDF5c2D/NEKyR1hmnQwEXdmaX/Ug8SDCr
Af/oaPCsiGYaKLolahpgDdqN5q8Jt6bhOPVz25VNrHUsnIJaaKgidfQ/uh83fThU0l7C5/5n9QFL
W1KocJTj8larI43DMQLHOLHXoLRPnvveEr9WReUJW8reEgN0b5VvGLJw5SaLddCNxN8KjCR/unTx
hZ6ISmqtnYN5iaAZgpmD6md2HbxMeXb1jrQcsVYnkai9lfWfW7IFi7FR9/YM8nyOImU3NrMA4zQ6
As8Ie5m+7e9DPOehbZO6fTIVD1BK89GPzr4o8gp1V7/jDlOyPQGs0nLSwRy9OqjVfppdX68upScz
CRbRFccfAt9j1CH3K5do/tIi5AtvQkItnPWKfNYIKcFpWd1xDSyvekMpUsf2YEwiU/pOdYGh0qdD
PROqzje/rgnwIPTNPHLk4SXDGMwEsz8/dtvi9AzMEHdAcjLLnAJnzsei9Jpg6aAUDEPs5YsFOe1i
l9EEijfFH+qGm4JsP5xN1kaRAtvCPxZuOOGQoicG7Jzz0/SSU+YT/reqmw7fhW3ff+B3yJitMsUA
C85GsWLEuoyaWDjTFID7aVqOK7tp6zk8dBSUcrSpM3H2ixSSuNdSWA9el/UM9YyHyO8JTdJujCtx
ARJueShHyZ5uv/oLFGofcUj/8n9C3yOWT//kLmHoAVhbT2NUHpArjOND4Rsy31mG4LbSHzUbfn0a
JiwJagLDMjjUNNtQRQ4HbyJj4QHl/BdjEunG4hseVAjfSqW8YOvS4uU9pEHNIa0wdmPtR4Oqhyy7
YSzO0Q6LRHUiQVyrQ8wcyimgzKcSmG1d9vX6337Oxa6cpIk2YEg2Qwk4nVa02/s81LHiQb9aagOH
1kBztE6xwtGAxm7bUSYg4AVCH/hgWlMErZo6tyG2DuogNtgAHXAgzNEBkFyKCfmPTNDzSBo9alj8
pxFlbJ9kHjVS4PTlP8wgvbGqZ18ti4okZ7aC4xB/v3Do1mqTO07gXiOa5a9KloBkT+N45ozxrTmv
ed6SUTrGZ3XgigjReSxBYYlBh4i7ofrTxhQLiRPAfXybkPYinXriVWeMUxPHIBLnBcbpkZDPIswh
uo60fO5gT2uZBbFeUEQM3c4LS8gG79U2ogzNtY8PcNm8zdGzx+TMM+wV+8LWJxBr/JTFRR8RaliA
OtUeZsQnor553tvnJrwdV4mhQy6rS0w0g0jwy/FmKSV7QtNneAflv37ZsAs2OLhNVwXjYGFgV3+8
5npa3Cl+BmdJknEES5Dp9q+1JNsb2muSdMTwCLIGrrNspsa/6MPfMPR2jfcZnYuA7MFVzgbHnKIe
SJzH2RUK/klKZWrffXG2qWrpixygvavBZKELhP/5R/RT4cqv9ICZZqOv5I6wQ0+GK2LZ5+kI9Gis
aVUVZRDFS7NrVuxNGKVLRGhMbSAzCGrj2C7aowcTWLl4Fz+RlutwujGhUiXgGSedzJFw7LMH8J3j
Wa7BMAiSvPQ+k0TdhGTSfFgCooVSWYDi5AhYqC5E9F9eoS1y/eZSd0baTId3D+6TCDrmmun16PQQ
wR15FJ+ohT/HdxsK2wd+zjkv1YkrlSfdJ0y/Jstu4CqfjcbPCpI2sCfBruJLdpDcj22qHcPF8oVK
lsEUDjB6NDbMilYfWEzAWni6WEZxj0c/rN+aWg6sK5BTzLggotlAeg3B4tED5IwnMg8xXvgU6nXX
tUyBEYhBATi5jMbprwRQIksZwbr4Ib9yeNPLpMKxh4GWwfzOQzhJiObk1NtIyhW7cMKY7m5KFvDA
4kNRPVORGv3KqrFre8YcmOjXLZjDlvImJXUYfmNfXH/yA6J1AHTM23ncCctkum6aQ1tTnznWdM7i
CbEM/K++ZUD7+CubgQjoxlClIN/lxp1VqRxdUeAJN/qgp/TvcUOsb9o0iscrLmRGoJn7pxCUvCVE
YfX4EE39bZg0Sqiq4SV+45yQ8Pao+3ULyFW31cLrULMCgzkZKXOooJG1TT0s7tASowB1sGEmqIqA
YoKGjLtomBBVmydHDEelgUmfHTk+w/jPLXTr4kdrx+sq5mZh+qYEz4Aie17MQlVv4P47Kmmdld1j
S6AJrgH0Sy2hWPARTiOGbUXlJ3v5xBoMVyQiiqNXDCcj3ImdYz/NQw4GUEKcbaSEGeH6enSZ10g9
JrI/O9FtalsnKvHGFjccF7Yb/msx9rom83xcEx1EuU6GtZsByBbqOqKM6mY1FEUdbSa3FD0iplmb
JPDqliawKyRkqIPiPo/fHnJyZm5VJAhW9RBx7HgEv4IfuHX5n6J1uClQPlYpsxasi+pjKW9kO7s5
ydgrd7/aghRdBcO0zP4CamH9CU1g7JQ9/+Mbo1kcfpa1l3Wka4yqbdYGvBURv+h0zonIyTYuW1hB
/MjKEZlB9o7gtO6en5K9t6H1ZPsL9dYi9Q3VsLWaDDPj1i9qxfQ+TiaCPLbAPQJm2osqrtlWjRTr
rV0IHpSEWDkzyTT9TUGxVvYKPgyqDYjBAQNSovVrLoEhFG3pNRHHdQw5muzvogtGPnFryXDle7uT
cUyQCQF3SXmA9yi3stTJnNmy8prl09fjivhMR/UBeqmuu1xgzI7Jd4N/qh3/xi7L1pH8fASzNDv3
5jvTHTWGiGg83gHfehNIygDov9FWerJ1Qn9WX+ieN02jdEpVX6ygvg4VXUoRuvGxTeqmbYecTDT5
3L0fKLtvHd8qRcRwx0EuKYyvlmPiJJ1HylYr8Hi59IS48T9noQfeojOTB3IKbGibRZ9fj5/6QMzM
giz+paOTnBuBI7iFkTI/poVfrSWjvRzDYAGJ1SxnRcxEN6VBUFtP88b/vrQ47wMNR0YeQGCTWKCE
ghhPh6CAjIvpOGiWB85cY/PdSUjIyHy3Xzeqlwny2QztMZ3pbwfaly0W+tb7d1uuNFcxVYoVKbAD
7re/r0at/fE4ON5NIk+BkQBFo7U9EGCUROsBAWSwjdd3g9FCyLkWzuiYW4x5zB9DIS7Qp8Dw4J/4
o0rKabzCE/8jN8qqlhJaULSWTKRmHgiICVC9XE+l/k96w+fEX/iZx720qZBNlTCHcqvKxAeinspH
F4NeB3PYy/llP9f7R5P99G90Jytyb+JESdH9dwVIjjUZuu7VtdmIsrmjdly5tEr4AxrKw1r5jZgy
FOcGLD8iXRSFrR1OXm7hlpqM9dwHH+TZgNZXJo/wQM7LpVi08NSK+q9JmdPmWlGhWtYDyN45Y4kt
banLmxZDrRACe8qxsuyJfk9iQbKclTVt24IVtnuwOpHda3YVoCUSNz/nUNASmKdYfRWLOq/kROit
geXASEdDX12gxxGlvFsfgLAUSFNkWl1OPCJhPOtOZKRqg5WB76QwDT3cesQq6YlWR0nmnDf9R8D0
/AwT/GZLPqQ1K+bfyMgtEQ54hBEpgQ570w3qsxPSeGuAJNH+n0ludKFPNEFI/gBOxCds+rMb2c+8
7aGYeZtRE0Bu3XaljjGy/fjA0r0GCMqb9PCaPJj9t9iF2O90/AFoDbveNruwxfrUiYSe5FaE3Amo
VtDGHZ1D1ezad7fYIr8zAAgd/4qzx1bUywv0QGZv3Y89OMvMyLJUpq4IBQqLRpib3JN/8petMp4V
IXahVX2iewDLR0+7fVMzgsWd+cMqbgmXjlH6axmK0myqdWfp9teswpKwyczn1OsZ1gIDHiuOLaRw
ZN5fRVeQ7OOMq47JhR5/obkcIzyrCcIBRQp3J23YiKG+3AIBf2uevVibV5P8gTqtsGh9IrOzSQIk
oZP9HPZnxd+80yWN/4q3z7v9ww8RZIL0/RxF5vFRZIDJTEeuRZXLElzFhkDo/+AVEJs6QT2DIc/m
03EwQ8hZixsqnyx/qmccPYaxGzXjr1fCtJ/tskdwcU3WYZ6QmL/F3VYDxIOyLd3skgvdnFkXCVVl
BWO+dKqff3ocXUGpzRbxn22UW1Er4Ssa4rKQlpX7mmvuiR+hyswxf4KTiKew98A+oBRTDr8tH87u
1+NFmwITKkcYWPnqFHT3cxFcbuhBF1FY05c6y01j3xqn5T9jbxROzafnkeqbOoawrLksh8pIkELO
tu5Aw5vNVx5j/26FRQo6iJ8WWX5vuIZrn/sivnJV2VhE4SgphqM1HcAjle97kOpJmLfH8IsO3PV5
jzm7nuDXk9/2YXWlJFdIccLwZLjxJkE9+vkPj2dYM0o2lZ3wVN7MqjR2MYOsdDvTJA3LP6F+8/RM
DLgGzFbeGynAiMTd88IPhh7QiC0rmLaInA+c57UFZtciFJkdx/nMlRiIK+2owMeQdrQfYJfV9sMe
uqyBoyFTpfHn9Sl8X/jjHnFNbaLokHD54kyXsogWc3UOk/FccyY+Xtmm5frp6fBooVjhAu4b4XkL
TpZ8sql+1c/Ab0Wr1yVamPZmLbun+wCrZc9gb33NQWV96AlewsFmz+gQb/UfziZSLz1xzIpSRGq8
Io1wOwCdcX4eNegbr0aFwDljxhZbfbdmc/bPhteQWU8Zq2TOnAtckegCMNyAqGEySzo+fhc4AZQI
oXr8wR9L0yey1E7ffFCBMSsAgdSUV9IxOm31/j3soSD+dbRUeX1nlDoNR9Sb6PWNKalfcKkxL5ct
E8/NYr08R61puyhqgElZCsf4efSkTuHN0IQMdAPqCBhUAd1UNKvwYxK84YGpz+fjIWnwhaN4k3x5
LIN9XWxt80Qn/eLZd+IfqVEk0LlnhLVsa+G/QVwMi4cYXPPqdBq5PXYaBGZfZNvNDozjPb/5imeA
/pyYo4uoroZ2mWQMyWBGgiedmSxeYpcCXVogtfPKCLTyrNMzPpP/K3FzgOggdT7ZZUmJ5mzbWrpQ
edqUU0FG/P8Na6I5FzB8pekWd32TNc6yz3Hk8K1tocuiZ07sNtrg+18EPh8VaLya8ICxejcGGts8
k7UoTvBezCgPaoczhNxhoZvjW/S0Zx6zSIh2NuftaDND/Pfiz5I5nVtskPAipTl8WsVl17xCcL+x
09vthS9aKxPNPvyT6sBA5J83vrmNwM0+XzxBTZtBY6E8Bvhn9dFtioEVqQ+TINcAD+F5qqCZdCsQ
9rWwCow7YXmNx94n2hbgt5l+37LKXUHngJhwBUWqVqFaNwahnB0Qnb4784pX18xw9mrbyNmxlg44
9VRyFOi4e38hPpSWrubQLvRrIjXD0NTrjwMB86YPXqXfRphRIbp1tCQqUKCARdbrIu+paURv5hUV
WaNk2RKGHgZp7xHNOhpX2EfYhjKRbnEzxUuFMh6gn/iogQ/2LZ7m04IYkwG8NVdDppWrWPJvNmzz
4AJgEyG9R3MUyTch0H1oX4B9I9GOJcw1ZpoXcEejRyA1c/h8+XIHwBAmv5Hd0vN2N0J8PHT68fAE
XtBnNRzFQxGBlL1tDW6HIGvvAVkuy2oA7SYA4p5iGzwNzAsxTYQB/nO9GXkeOvlko9W1bzhTX1Yr
wgpEJYj2+qHG62MTY5/rRYNOzhu0U792sw4J75xtLwFYe2b+9TwVFb+G1O8vrzTj8cjw+Tvk15Ty
2bLXRGIICRCoJuXVu6h5itLEceqj+TET/3z0/lC8PdAJynW9zQpgMQNhzIYTrCzIW9L2JVZMmXXy
8fasRjV1EDn7NI98WcLrRK2/oTWqqCWoGkdSW2OUQ+SzEThwlu8RAw7gw8dPadimV7UnjsUdvLWs
qOuLrAPLnDV/GVDrFqqtI5K9Or9Hfx2qa1ze7pa7ynE2RKLnPPwxX7ShWEPUUvsuIoGq9v5okw+D
1c8mcTdm/FhA7lT6knB8XUT+DhYJbUGs5QodqC3aMQOtgN9MW+1S65iFgwtmTUSk+EjN9lRHxmY1
Q09MZ50H7di9E4dVaBSrlxKPMoWyCaktjHY9NovhS/xjsH/y9yAfUT1E2G6YZ7jeFjjYgVYdFUpv
/jpMxE79ZOOASnE4JQOvMPbmv2J9fGUW2xdQ7nM08wwAUCOrvMDUKJsgeP6As8sbyrw/2z16DRgw
+ema9QNwdO42rtvPjbJyjfyP3QdCH+miJV0mOlM48czwbCO3d1V5MGTc00tCjJCaA2F6mkwG55QL
78ERjUn9au7WNDtZMeHzDfPw6y/hQE9Euz1E2nY5QqdHYYXLYPkv0S0EOxh9T8/X7qGSP0DLbxki
uYykgzUtbqLHMwq0Qj39CUob1Bn43ihqLpdMxVCS0is2mZXHyTiAivXMJbENFkMY949rp/6zpLmw
lBR5hElv+CRHoJPSwCDd2jwDzkTYAOwhN7Pr+G3SR3Md/iLZzROSCtTS37DKBpiNWB5t+lMW0Yvc
aBgv6qz7q682kLHf0KOwlIqiWbOwjmiWiIlE9j6EbDJFhbBoHN1d9sU1A9ZqpA87Z5QjTFGuc9K0
vKqi8qH2J59sDR78pJ4hZXCLJBxBisLXRTfPS76SgK4pv59WHH/0yShEmyCsB+5PSNNRyFF5D2sN
JM+JAZFtXYAHZ2blt2dczG/uJHXccDUSMf3AiUscHjFzcBvr1C7PKou72DqL+PAj+PUFDHLl1ouY
nNrBmnNCyphGaN0SEvdPS1v9g+LBToHAAlDjnK1fYYNR8eJUY0Jyq9bZZ6BVF/vuv821x88Er07K
18ZdrO0nfGYNTI/1KtyOFnI6D24ofugZGQAbRhzIGrLsZbS8C4bY1GZhpdjdNaMiHReNBdtwCVdr
A97JHmU1oSTVEdFZ7vT5Q50dCLrODEm/UEvLoTyfocT65LqSDj9UFv2ht3D5GyN7gs9T2REtqAHl
liXJakei3PpHFhnokf1QJzPzlzUM+YEUmBni6vEiByNP8XvppGRoUmLDAXWLPBLDQ6ZdIZFKptv/
Mk5VeAjfaphvL1bNSTJgsh/dr6tgw8nITU9VwJM9Kp2ieYpH5d6ilYYnwdhxJ7bTZv5Y9r0554t+
JdczN0HXGEnV8EAZbbc7wUi/4nVzu7Yj/geKiXP86UsFUeN+KfCsuTK9BoTTr+Jc6DnoL1gSasqi
BSt+YNkozvzBwEDezeTpVFQ+9Gb/kLHCxP2nggp3FSMcMqiXt/SYWF8JwjA4MCqoaDxFjVrcSipQ
Hd4U6fHlYaGh6oga+fsnZ2MRl4wxMF9QYDuMWa5nKpBbWPHBYEm0KY+RRzc7gcwnfDg/bYzT3Y6x
kC4BPoe83GUM0nDnk/j0FZ0taPQ1gVXF7ZU+yTEyRoOMe5kUJCMmgbuOMkSoz9IlA0G0tBMga/T3
AO/UAbbtwE2pAieGmfoxrrddqb/LTUyicDqJOlKsMzuKtO9r5m2a2A3Cg5i8dMJbIU99krlYNGVR
uQexkuhnUHImfnMPhY1IC7EG2KKclFsrLLSL8xe7C6kGi70vKCNoIq1JOCDqpkzl3cHK4up4SaNA
cGckVF4bszUi53u/zStf7K6KoIR9VEf6ZZrJbqZOcb2YpravUnXIQQyhrNdFHU7r25XgpFiljAJt
/Gj/MehRxDdUnFM3J/Igk4MIjSmaG1W3qXzcxukPHjBm0VWkJVPMlI4JsYRBbZ+Rg13REnajTWnP
Ne2tpDya4NtO5HpizinCab4evcuZ8sBFWfu8DP9OAH4E/f1B7AFgYOTvLZXPavZ5L5YKl21y9nJ3
gtWhPba2Y0JDHeLsbT6t8zAuXIYCLrOj2mAfRIvqhPgcQsV6+U2/Vq6e8NzC6J/BMa075JCNnrPl
FRKyXCwv3IwUazcowlJw6SovDjyHmMP718ATM1UI3uh9TtEuMeG4lKwugMMx9uox0i2fqby9hSxI
96gXHfXDZxRMpa6+tpsM5LRHD2qdHtZ1PovJEnVKXeSBiSom7cwTMlLYARO3zgjLk6vKCqU1dcoM
tUaknf1wB50EeZyVJsEcHLn7s2knm4QHOvBAXpCZ8gycdksubr+sm4AO5f1XBkMMR7HSIhs/UNJ3
nXEWLrDuRL2u7sS+2duUNDnpxHfkkYQN4BMfqSxaEopkF2Qr7bN0bDDiBDijCDXwNgU38irwpxKG
0fS1tN2elGkaF5NZOJvh2ebxK3pqTS9VaHgIIdoq1rc6Vg6Yl3/kp/mkl2cMV+pj3HUwtrmcvXoA
gl8D4PI4xNJRiWbjYpI5dwHNM4tHMiJ9RTmtMGxEPjcg9nwfgxEHKSVHghB/R1HxiTxTZsIdJUOG
eaTKlujwT3IiNJiGUCweiOvurvjIwI2ORzyezZTBl5g4/iHoLnbRBvvrvHeNsfsDRLkazKgxmbHB
1JN/+Rcj3sZQJmkGf9J9ZrCAqyOcB0PDcYbXKWnAxcrv6yllipPetKmQF6Y4WrfSYJuYUnl3JqWc
I5CbCMqQyj+RrQNAqf1ugjVHmSivRC3QaJmOiF8XxjLWBtowOZykCq0Q7zQ8+y6NDUcO5hgeA2ff
OxABFnhBfO8I7Tqxw+7h80AKAyojKIQVxQhe11xJbRcS3fPXBU7br4EzWV7FpyrpfUNFbEGMLtnB
6ihV+ROv9fUKSD6lD4V9UlwcoDcI7lfed53zy/mYldCIpoLUr5a6Ou4EDjxHvWYkA4mViTSCLqf3
AQrriHwcrz0RKUCeiUU/hHZtM9g02y9EiYVxGLXMRagxOuJkSF4v33UgXHZkrCa4PqPQd96R+caq
Xh63gAs4Al87s2Gdp9PfrMYwDk2K1ql4AVGOeBXU/pkGKfnVWVZ9So+5fW/sKAZO7e4nvOydYyCr
Uzr564dwZ6jdIM0VyO7hrsKnAa2Gl2Ra3ZJsBa/gmIRIhGapHE482A1PPmoHgp8Ni2U9zfKfcYpN
eYYAitgrZ4cl3//gGrEpqI7auRhLjP9KZBIDBYRUYKRjhia1vled0FmCDDHWJmo4fWmtYr5852z1
pw0UVuYHveL2el9pTX4fosikdEM8RQsiq6ADj4CkUUXMhASH+5GUQChON9cKz+4kAY2t0Pmg8NTy
IPWOb/UTKwhztvSpyf49R3l9g27ONT/q4pTV9xfmaNNx2raHv0vGBk/0zsFBVu8oBx52BeUuWr+c
c9ykgagvc9y+h3T75TgX1B/S2fh5zQWg5tGVrvkCvq7nlYAB/wPwqotAXTvaeBzJ0rtrmxA+ZrSn
j12x8g/HUfbfe4BhSfNjKsA1dviMx3ngYjtRxJtNW6c1+H+WvH0k1llVJM5Z5Prn4TFRCC2dzvlC
H67hJTF1pCigyj/NSA/WVCJVk7TIG/4gZG4NsTMhiwuE06EGihbRdpcK6qhZQ9ruAW5EKMdhSpjJ
y0fPAq7dhRtqQmTt16Y7l4DDYeCDShSopfo9hm9xUcH+AbOH+Ia6DQq6MnJNlC+a5Gz5wOqjiQmm
iIKR3KcvOtfp2o9e8AyZT68NqjkpubWilX+EWt9QIHr45AsCBo/k269s5d0EQHy1qO8RJhwrlYUF
sxb71/HpJ4f8zR46mrpq4xd2M0Y1jJ0Dtyjt0l/f1pmAJRuUi5sVwQe64hjV+QZDegk1gqqOfIpU
zl5O7wFi9xUuXrfLckhcnNVoWrBZOZSEfSSnPDdIciW1ytfO6KulhlwWwya3VbzvXzaB4nmUG7T+
BvahQue2l24D4v+cXBai0NVv5eHnWUckR3W00B5/V2LpzihQglYiAzPT/xOLcJHFkvb10DFTVeRT
NVGGEjj9GaUxua2oPx32zzrq01NnpQEOyWzn2m7nk4eWrSS9Uy69GB+1Ny+tYqZmXMZpgQqL50Uw
ZjpR8UWGjfYdnGaOCftfHHTOPs3Xq3g2tiwdrijngNY6bJB3bPKQYTrWtRDp17V3MbifS7y65ptT
384q9UFV2Uvb+R1hBWJJBJn/4kXT3kwq2a/C0FUtfKxiijX3NZe8aTB2l4xetM5L5fpQxvBBYQ8+
hnTmouuM+OVZxZRJX15HnBVTRLxCnB9xHMMFV1cA4gI/VpYMQrYzC6o2Ag1a4nYkDCNnwQiqB0Z0
bOHZ1r6dZfOuZqL6OeC8ab0Rltg/my+pjQsfbyeP7vtzjyS5Or9pug8osvBNhZF9X+20G6nGZJ+x
ailGPgzYvzgnNqVu6nRwKtw+4Zvt/uJOqvWK98aighziGQV6G8eReTOTR3XFk+W4t4yyrH4OQ0+Y
CChBlFaMTb3Ee2kUX2WZCm/wHZtXRCiAVTdOiIAecfLHC0ijYm35Cvbw9zks8+qiQGM8K+PU1XLI
E2+wB1nSkq9ljuWGSMVapmgauMoW1/k27cmBXQBLZafZANzZ+VFboL+woC/HWLYQxSPsRZRH5rhG
foqh+FBYF3O+enDJQcCL5qIhTUWqze6q2SfAz0XcQ2p2s0T2e+wHyTzRoSwruv0O3XGk2aOXEpDG
/LP8UEmSI9igsdU3TYU46im94fpXzH4g01DHOIjPep2m/eY8U7DVInGcV3BgMn1vjFu9HxJh0kWe
RypYTx3MOU7oess3/Zk0xdPzFPC1i5sAJS5wJBvmn2xxx3zeT7timydlqT1rq3yQ9bYiyX27Dm11
5hI3IqoaN9cvhL948EEXGcTRmd7wCGOTCZCESWnJBQwysyUEf86OrrmKYj4altaEHnEo6gde2skd
dsLT3KqIc9WXUyCqgDmeQGZ89sO/3NLhaAjds5d0S3vHoZYBybN6VmBWwXE+cNAgxd7/neIQtD0Q
Rqh1YGxFEoK6E1YTRJcWw43IIYi4m98ZrNezb3bv4k4pwTc5UBDjSBFtglgE29kkmsWPe18ltwA1
70xvfrFwyrST6kcbP6WHUu+fqD2poJiOD5u2vqGQxXEKJ9M47qCZSPSqfRa52M6Cg6IxRdIXcQ6L
KY/FwzOZo4K+Lqqujm4XAMm89SZvLZRqkUnfNGB7omeaMohDNtuz+2ZcbPqczb8cvlCR77bhILOo
+/qftGgnUCHVJAgaKRpA3USGJK4LyZlxmys73XGmnY4xA3OAC0/zJ2Snwnf10Luejp/2/OO6xFxo
8QwGqt0jxu+xA0NL3BdOJzzC6za0cDn+ND9pnGTaWlWM9kdvx5K4MBk5RcrmGp3FVz0NCaoMkPS/
LFIFj2hiWn35GWGeGh4h7cewGYldxhmZTDss/kFwUxCNjLOzTrK3pHZVtNdM/sLZ5I04zDOLIKQJ
HkwcqFzot4FGgNg3d87aYPZsOjCRJh0xAxYe5XhCPF/PkfmoU2ZU5WMEaoHSlhupvZ2VvnKfUdy2
q17NbFdggK5tP41s0rFqeZm41Gv6cQhRT2WW/BObkn1+oHHm63ikCPRcFM6/ulg/lclTk42jIujq
X2+hU7O+W2bfvQGbleGjGLPZSU3qy1049LU/KmAxssgi7BRSEywUIpM5NaFiiC+j/DFkIZ8aWrE+
LSaeeo61SjWOVYdtrTdmSRVl9I4qeifJt8vcbpo4mMKvoz78c9fz9lBg2rGBXM91GPzo6VwPiPSO
rLfvMPDOLpV0IHCWfZdNX4tjK9DfaNI4XLhOc3KhkPspOpQvDNL1zngG9V89LV4gH28YJoB1UFz+
MYfdKxZkKu4ZcC49bSEXKbPrzTIQOeMgV21+0nxQl7Z0wUcW9rI/eYnBQguP6XDvvr4fceYn11SR
f0Sb5LX670BxA3lfiWnIxaCCgdBLi94D/tJSuippFkEjYbASrlp8k6fwYYdI0n3gUqHR7rMmK+80
8f+rG6S3ZTkzbR08A+mmA4hCOQ+YM9BwSHFbTerfzgRMAJVzq1J8kikdKjbWD/z3HjA0AtZIEmTo
guzPPYV6ofJ8EKiwvdLOmt+oUUyEvyfq/I9M0UCmcjvnOmMJ7P1QRNrQNjPzpq4QMI1cjyL6+v6T
Q3Nnbhe4Cy2GA2anm2yc2tEJAZWf4Xgzb9fzi1DWEGW42hRVfPdSX3LR0YH8uQpuNrZkospCMS/q
iWv0JFusRO8W1YmO3jc0COBguupQolp/X50B2h8Rg+0e/THCVph5RLs9sFeDHzDOib2CoHuuW2a9
yfvvOxqjKz5EYa3TG5pWUFdnjP/OYUupdWvED0Nwe3scZYMOjvKTPNP0DjPScNXCfWfrLrE90IF0
dnijseD6flGrvGm1jE1Uvp0A/qfG37Kl5H5WRUKyaxlkE23HTQxJ+tXBUKwXWE2piqeEU6wGkL8J
2etOO59l76/+nOypXTRzgFCSIe3Sn5Y++6/wP3wvfRHepgPR8zaILhbkeSa5nrbw1JgdMvhq2OO6
4T6h0XGyOSJo9Nk9hG/IArFHyzIIuNJyWJF48UYMZDAI4OHGZMwpFG5lBZfLU8+eTGnWp/eCXU0D
0wo3C12M9a9WIpcFR1ZweWFnR8LfaPoHDFdBPNqXeDOSQtyib7q96her7/nqk0oKtusD0t7oP3c6
e39hakyqoFNGIa3yfTb6O3X7rNIDOlDeQN7CIhZi2Nkb0eUdvlSyE2/CVkfkoFTr4f1GQIQVWrnH
h0pmAjO5ixBK9DOgjYq96Q8VJ2sh7N9d6+Wavlq1El4CLmlHy1AgmzxD/nq0VcEUKfNvnV3FQuPX
1rEb8YMxs5ayt14YNoslKU2vpvPT2Xl3BAJdgAdNgMQ2UeCJbSgqL4T+UCO+Kr8ZHwnuA2MOL+Wr
Xw89KBrJJVsCwkXT3155R0Tfl2nIpeEdjiaAL7jl3wdCVy/pqH/lN8xWXspfm665IUpWRQgkHW1A
i47TQ4Or91d1+ztq9YJhmqXSPT1fl9w0LurwMfwMETAvHvB388LEF1vz3SOXMuyKWuUhqs3jcDOc
UJcXh6QaMvI2gTPeSjcjcZQEobPui/50Yo+YswBQ+/1Po8DtZ9+gx8RgJ8yQoVje/qNBb6yycL98
zjTvsXYVh3pfscigDpu8PnhMVjqBinuxk6YyEzhyyUddD3wKYgmXa3MUTLDlljA/QQxp2xNlI0KN
HmwoN6mZ6vMoNkIrS70aNUGszUKiIhgLe13q9U7g9XMx8ztCLIi+FD3ZZpmj1I9qMb8nlkRAkFvn
k+6QHi1yKDtpoj7HjK4Ie3PMZK00y4RxBIsKHWo4TD13hsw4VFEyHaK58KmjXIew01kFOLLumSey
alAjPlaRAMNJlY7F6wRlR6/pg8rALUoBpNVyx3MG67AZgimVedH9DNA5aSb8Y/mbJuHkAX45MKIP
5XZjlffSPCRrMdOP6bzKBcyHwRJBPjmmzxliHZ/Ymja1xAMwzQWfISFchKay4mRqzwzmiCc8OaSZ
USV1bfiocsYFG9ayjVuYc8xmBeMwhcnXE0D0JpZ1awPA6ytvl0UxpTd21BYw8FPzzEROGU8Cz3+5
WB5C1XfLr4xh1w9ny5SPR6YnMn6Aki3nhJGz0nkWfEdEQUXGbeD28Oet85xcClPBgxfKDc01LfsH
BhflncpLGswYf2rCTBXCEaQ/AHqyyl5fjsSqJFL5gLzDWNop7J+AFmmhgaq7c1I6e8Sy2cmIYmPw
m+0ykIKMSYlwZZ9OV4m545NHiKz8g1Xx7w35O965oYg11otXJb011SnHLBABJC3x5LLNZ+fnmdoC
tZnBiC4p0DGfneYSojhha0WYOZraJS1i1hzs9kBc3V9cW4EXYMVf55m7FMkcw8jDTpQlQ8405CAD
629pnnb8SvV2yQ05AuPaELeiZHFhG+ZTHwHOXeeI/F3sdwgPlTd/I9YZ11M6VvwvttofEaiaF8fH
eAILQ8NOXyIZPxY2S+9OPeckWoxEyoB0qnVdfs7e4wWD0YkxUhHaLIncyJEENe290F5+pJ3gxAs7
06xDIVPnD9fGTELkJqbpVn7WlYzeOQnwILqfSqkeYpp3vxvcgUT6k4dLP2bnM88kVrhK1DlfzJ2O
98C4NoDEi9BsXlC0DvevkPKeV4rBci1qF8647t4Oh/tlDO4y2v8m09+nLXC8H7czyoA6mpxZ+N1p
vG5l9/mlL3PrqDIdcdfLWHnsdHxhyDOOwW1/Mr2jnbtZS7J7JG45H5LuqcQrjN6JjIzDVEsausAc
5O/AdMmfrSz9oBSi1lVhJwwsy8zWvirkHgf1xXs0ZXvequ3WG9dioRrrw7RLUMNZ7ZrfeIakR6Cw
Oxu6PvN34ZO0aIkHthx5XH02stkiepS+33iIMq5h8rR6zDSHLIymDrb9sr9FHX7Hd1XVTc1FDd/Y
17O/xDhFx+EbwRqINPgRAy7f+Rg9FXcFX2AeA7nW/N6zWkbHi7Icci6MGpfzKqDvZppJysaIZAi2
cyvdspayCckJ0VkXpYjepRpXrmlhvSghPu/q5cStOvE4iDYJz35LympAdgLHKOVku2Vo32zYBZLg
bwB4eaXaluQKgNWFm1fUYtO8/QZct1hwdmZgkr769MdqZgKxY27rkP5hVBiR8UMnsKV1hhEBNk6F
jSoWXPNvP4sy67QxKb/LEsf1y2151mh9kjJLwIOgBzmZayozHeOzHoVMARGz7wrSK96OVkOFzJrx
xncZM7cPelaWV2ecpRSkKxkRjnoJEHY+LYBvEZH+PAWAvWAYRhi1E9ULpntTsvtXLRRM4vQJVEqI
fyxsGaThNRDYzzFIIjwtEcX9ABPWQdueSfE2p5rVR9fciXoDqFoyC+dqEhXfDmx6K5fnvF8ttBlw
MkKkEwdcXgsTrvn+dtiaUEaokyoUCdIysIClgULPpUi/bKMxsT+ZNPmmYqayssHQDrMcFOGCOJb1
jk9Xa7FdCJ+9lnd2fNY2QJnl0mkn1J71oIL9lpXfnQCgTE49gMrwwKsYrHP+YaaiGoQ2vbIBMUQU
3EJYcbvLQ0EpHI5iXT+Kat37iogK4h+fwNk2gIk6SKqQ5oT7SlB44inFrHVlkSRNbvKHgpVSpr4H
hAYpgav8uMTUbv/BWTbFinQXSKtDQ2giG3Xslgu3nMBrdafEach8EdiniXQShLLLtOyb3TLo/qzs
n0YO8s7Jv5tUIJjFz9NHgpK2iimL3GK6KLZFf1OPLJ8GxPlRkPiU1sPeRsbRIq4QzKuyqOOUnWhE
pSCRg7n6ynXDPy7rD/obhh772u5ya1KSAi8/z3oIWi8RjTkWA3CqXg+0X08vNlsn0JvxTCw/QP0n
Z+8K1sh+sxqxp4Aa8tqutLMP/9pWA8lstZk8aJ2Mn2XkkpCqjrfsEGbu40+YUCBCl2Zof1YF8psA
y065Fvb5qYsz3Oh5iK0nuNYrG+x49ABeK/0RF8qngcoozS0S/wky6uTv05YYZdLd8vAGcCtktbm/
POPgfpuJbeI3caA0b545jSXTVk1OXbRPM32w9QaOzDkXBRs+A37wlXzCwLpVqK/B2VVRNizL82+I
An0SF9X6bAhF0yo+sW+KKV75vkW/5IJF9REzZ6+hjEBB7QRcQviO+lP0IfctE1c6no2S3ZkgW/Cj
6PHFsErHi7GmEb1vnEWkm8DD01Elx6QnrXqgJqym29XJtvTa0s4EJ3t2PIQksVMtZhl8KHwP4GBX
wso8oJHskMRLFcH7ASrhB/kGbRTUnhKhaWs0mqcMkiUrIKw3IuFWd/cDkuuliT2s5lx7FITWG9WW
qgy+Dv2C8H+C6Ds/eBHeOWCOODkJVll+Pw59/V8O1k21yMpXMrWrHz+FGZaUwvWFeMAlsjAcQwyI
OBg/668ZiIUUQeTXr63zgxmIzKJV7K/2uhiCLfNETh1kd/EzHp2bcdgAZgh/gAwX9CgRSmhLU5iz
NOWpF551fR4ALRMAByARTW3rkHnKtWZSvNxBfcO/kvHD+cbsWczQxh0pGUiRtLHcJ+CMnvNEBg1e
mjWe4ePzijFJ98cFFAOqA/5F8hNcy5pcm4X1RRRgiKkaSm5GhWwglDbc7gaaTeZhiDSeSlVJYxLO
usxLXgLhV/ilNbOsQHIWV5Bj7H7DKuFjKGZrwvHdcudVCQx0P7CGIDWRDWR+40JIu8WSl0pw0thu
2PCu47f0cL9uZ3TR96gQzuq/4Occ+Q2lmiELId8+k7HtQe9MkRN6k4/v3wIDlWHfFviBolZaEBY1
dPnH1+C2KKI9XJZ6VEL2U2gbyb6xDV68/cfqqgTqh/uDZyur0x0RqQQqSHOnqtcQ6Fh87zZSZYfm
3NcdZReSt/W9DnU7IwRsO0wJZdjQ1VJBbc49BRvV6HuTVIxVyR03Bx6chsVj1+n45HmKC/MB5k8z
f9msnz+/751H8RKXkLcZjPNfUvCdy0/MQVRKyN9RrML2KrY+h/rld+psXLjqoPcBtln9pNFAHsU5
AZot8QETVnz0raSZ3tYITSR1pszyvly0M5nHSpldvsAyVsRC8Qdcvl2PwI8T7CGQvnIVdWUzAsz6
WM9bIakPaqahmtQrCTT2R0XS6hMMC7/g2ZFOwplcV1KJvRIubRn0aMt/NTDXGnHT5kIsnj5fUF7t
LO6lwfxVbrFRLStBs4yB885OQGM0EvfsAp/+5zWWnwgzu8BmxHlTON7S1YJD0zxu5tLa8NniUtXq
XHrJ5LeIDjAmOBq6aYXewJmnXHa00HFbSNMgl12R3oBUqH5+DeLcLN1y1uaHNB0m2S0C8ibsI/bx
BMMpnVinH0OI/JJxMIOpFsKWxwUfRS8krsbFP3d9zf7RciitTw8vQgXenO8fwwmAygrgAFCIZVGW
7yK8BltJkGQ9Ni9a0UnObVP5MHF4OyV49kOFV7JPHyPxiYA6GvbaOZnn809Nntgd9wNl76E0vicr
VkKf6821o/+HiYsMzYXMy83FoidL6/Cm6F5DyXCW2avs8m85b/DgHXc2YL/V1FaPFmghoIs5PaOH
oGrtpKXdSh7TtAm7CM1losJhJjHPSTViCAZjknCkE52wydZKgb9kvWKYFO0GVVgBqXmswbqcGR2B
bV35EYNRRDhjA1byUoj5rgkbJzMPxD8QRU4yAG/cfPiRO+OF0dYB2KN5D//JHvx/KdUZyTIP88E2
oArJ8PJgQSM9Hq4E/6EY9wTbwz8K3qmKgvhSeHumE6rfyTll9QqBLsglcmU6t+1PJvOFx5d5iMe6
nZQE9GeWhi1K8dKJO8cejXwrtez0GFZJYaxlDEiGLDEDT0HuNIRYSbUO2G63IXHTN+pwAQ9DHwzc
nhW8EIj/yaPIEexpjld9fkLf+y4J024n77WZ4B9js6g3p384Jtb4GrpyM/RySEwMxQjMfAEOWjaX
qJGUXFeyqyQUH0O8wPXTjwPG8vHa5APDeB5eRqlEN5YZ7iLNRdTxf8RW5wZCByR7Lm48VKArOdbH
2yI49LlIKiZdfqkjtdSG9Cm+gfMmCqpnzYDLRBTmjDP4KpBTXEhuPtlOX94uY/xKdtUpoGliekmN
6XIQAWGtpwCIFEX9juWxbh0F2049JFfyRTe9G9gvoFJgQdDr5Je3ZQh24UgQuLn57WGH+iFphGkn
c7LG7mUvTfugpMtkeD2ncso7yqDJG+tlDX4VMR1Ox+N1ILKgWt8tB+qtb2sIyPxHi1/e4wkiY9NJ
K+89gLKb9wuGInQqmqb16PqMjcyIe4CRmKGjHsPzQ8eDm2gCjoMptTeAeriUimauRq2a3d4J26Np
fUeyjydMlDStLhH7eazhSH4Q1Rjdd70usKCOV1vg2d84r7gsahMnS/Cjla/rkgeBYbjfA3Pj12UP
goJ7m5K+oYUdBL1u0dcOYHynLJjSmsBAM4LP2CPFY45QU9EHmaUx8d9jK57fhcNxUEatMgXcx/mP
tE2n0U2C2p9n5WL7yQ/3EZ1WdKxG0i7Jwb6xMBA7k3nGSkQX1jOzUWI3to6CrrPOX24LaSfAXKMZ
hlmbDiQ7kFgR7Lpl51yHESu5dUKeG++ROkSKZbk3dfeDiEUpWMwQlv9bI4CmPy6t7BxyRr5iCvLj
EBp9HD8LAW7luHUtOhqTmZC6KTZ8dVUsEZXkOXcA1EQe0HysJnaE34jBp5p2STIw7UDRCm04oU5w
/gurQIbg+tC3H0LL5VNQoYAvuLx3osMgxtLjglUNTww+Rj4gJt85HO8YJ9BdDwwSrgur1kCwuF4o
hLykNBNVOt22JKA8RY663wpygVoYXToW3sSKn9JZ2Fw78O37qfZUoc0A1Hu8khGealqV4xVpwrxe
8UsG/69G7+zwptnLQRKGJzYZ4qJlOonrjWQVgSTDTczPTGIZnEGcOn15PNnEyCx2H1xoStUjxB+E
dYL6+izJeUf/FyM4vdHKVbARM3AAcgSYJ/+GdkIv70cP34a+Ok+49kF4GuNzCBlS3etWZEMteyt9
tFaJsX0HDbLnU92CBo+qdrwQRL23Bo21hukV2AmidlLoCGn9fGuzli/bBPjNBqrF7ribGkTqerbI
URihJnRW8YkMh9hlD+8p9syyoQR4Gu4EMyFLvLlUyWeF9P93UHR7tYaSGAJMtBsqqUYrnSvMEL9P
ja76INUQ2r31aypiGDY/pOdnef0Bnq/uly6XFOHbrk1I+KCtA2Y/qDusVNrg+5M3NfntQ+yAdrPa
60Agmj1897Yku3qnEuOLPTgPs5OOuDZwnkq2903O7An5yrCuULpoZFpOFRDmOyZqf9KDAvi7TmSS
7MbR51ktCN3LfpNA6GeT/7jLhmsT7IxziBmw2LKYiNA3/6B60/J/yiOcE2FsA8ASby3k1ZGduhzf
q1y6poH3IJ8Q+/74mPlnior/mDUOzubedimMq3Pq/XDlmOC4W9uUCtcmp8FPfFuqWC1Aa6nYdEDT
Fl7TDaND6diMwmUTpDiRFbNj/+gfAnrMPmiY+arKm8hMF5XGy32cxmymNg3rKY3K/6Lz+rOwnmjM
Ie+euIy2huKcB/b2IKy4IOdF9FjUYgZYsiD3dl5V6UQZvfnjKcLJSgOg72Mt4bjjsEHXUCUxEXi+
8HkIcWOfHSncXIySKqz1ZLwvpMKTpeO62IgjpdVKkmXndK1OR5eW+yQdflYKcsf7/a/xYGCrv9ms
TFTr2D4/TlfPs+9qu1O94gjeJkIlISPYSbw0yYSYbf10uMw8ZXC23Z9843FB23GufM9KcNPIw52N
4IMazp3i8zZj10QG64LWl58WSrJTCaH/Hs+gNgKEuU31rE2B2OqeoJBUSqHPwzc2AaBPc6wPL+pa
sIvAtEIe6QcmGk91Gy/RKOR7+RSC2co4dNnaelAtqO4z8t9w96vvUY0nRfsQIRfmJGM0DKuJ5qAW
l0Up05Gb3nU/G/g81+UBkVAsSGq0hHvpMYdoGVP9KfSdRNl7Wmj28kvaoL96pW2UtJwj+mEStVCL
DyTQ02ofl5cdk6DCiyFb6mEfR56Yx/4YOeI4ikqIv4sYNTi74m4lcoHrf6fKD6CcNReSFbdIShkp
9wxhnJiCc3u2c8D+crae01G18h5Z5SK4ApgOtfC6C/201O9keOtyjXxjnbYZxdyhiFPm5Uyp/RO5
MmqkXt/f0ZzVi6K24oe5LiL6E8CN4IDMsoOmSF0Tjj9yL8G4E/Z3hPR8dV3rPram7YdxjFfC2B2B
96izmHiWHb+3QgLl49ATqYJoQ2y8qeUuAqSFt2iiQOE/qqWdUDDRDhoX6Kwvx8/bZsnfpYoK0E7i
CXA2/ML11KgzrDRn1BlXiNXtzFRAR2B+fVGPlXunof17EfgFVULMfjSg/NCpiaU2mQuqTGYb6Gdr
46xCoxUz+8/5DaIyLRMphPJt6yVKzehanHq3LZ1AYoo1sxa5fbYRp/qonRug0eGKobwX+4dP+0j1
72JVGnvvR7FYdzvzGNon/9ANcxHm3nF6wR86JDvnr45/jWlW43sI/8ZwHHlXZlUrnuhJyvDoxLmn
C6ozWlctfbwHkB/MM9LOi/CM87KZ7grHHGNsyKBA9kpXPQrPCDR/BKMYQiIy2hIYDdrvZuvskYH2
80iNbS/qvuobR7vUUwniCOX4g9ut/9WCgNyyVMvKmik7Y9/XKWuhBVlJyi877FJseQPMua6SxCZV
j1kQvD35+1RiIPEQgI3GW06ckm6sNQLlwcLUxbsl9VCr4UCmteTSnJSkwr52p81mw3qYy+E/SDxr
6hsYrCYXqxD6uY9uxt+dSFfecJKXIFXOveDY2vuC2jHg/KKbXXfQftoQVfL88unaNcnj+vQ7Mz4s
qnmS6ZGhl00ognHv4zduKlohKSdMiNACuyedPTI15PM99/9oSiXK98olxci/uefgmTwE8too4S1f
/Efh8bAdxdDl4F3HfDRmuoo2nfnjXDys0JOeH/YtR9UN9KgnnGn4NREXfN0fHPo0noM/QxRJdpGd
oWLnDVCKrnUbv27dT1lSBabnBA2lZ5O5hnD7ApyhseWbPGpkROREp2PtJALf8kRqAM4jn6wbMEUV
hPPj2MDEeJ4TqnW7UtSD0VzQbYfrs2+j4nNYd113IBc7/9vsLhSk3PLgkzAu/Yqik9oAOy4RRqyt
35cLZDEPy9p7ssylaCyYQVDxUdWixKO0LPzbTJTtp6zSppOFpqU8TsL4lvvlHiZHEyUC6vY9jqmR
LySDOHu5Y1HCjT8s8NI8oVNuyngi5WZodEALNdyJfttRv8hrIg4IfbBgswgzPPXVYN+u5iKE/XIZ
KRsiMoA0es4/c8Duh09qq9Idfe6HW5ulCJog3zPa6cef0raaokwPV+IlgBJl/7J0CYqog54/YhXf
VXZjsVG4JLLPlhwFF9GQHpUxZ81emnrTznrSiGVvNOVHvARf8S1ty8I8s4dZU/zWLWwJ6glVOJEm
ff0AI062dsiz6WoqhsfB7zKK6jjfxQMQ9h/44NpW7hgtpqPxJVZAi3hnzMah9cyFF0pmAzxPS63m
7fiYib6nfcMYO+0GIHTA7TNMSJP44jGrwCmhZpcK3X4sWCMYUh6/6BVCSBJWzyjemydbeR+aq22C
buC0yzcbprhp9qhHJPGGAcDF3URAIX58MYLOaoleQ/OCDX7X5vw1NIKienaR4U6gqCofTcTSjnrZ
e1GdxvCO/BdMDz042E50qj5btr4oohNvJLET8vfOHxCLtPYjgKNViiluc5iplDD0QWof3eCP3Mbc
LndOcBwIgotrfNgF1ccGWJQNBwY72ssp+fT3nUEqkA/WGI9uoC4YofwobhmrHx45FYJFGHcB0qo7
dF393twlhKBHzqnSaSFffaQKBjuzXJzqwuQkKhQ1STdvQqhY0y3QJky1SeZj0L6kdof5KRgVp/9b
cIozb+NvKXLt0O5ojrH9clLwIAoCTZTn7SeomVxIzdx64f3wmQ4Xdhu9bdKRFUS/8VGKNGLd0eP5
EheopOZNZIqbNpq0qIu4Io9wrR167MdcZOfDr5hZUta+z14Y7mNfYRiCUgp/HF+ZTFXd3LcXsV2T
IJDziBW/b403P8gQ/5bfMyhNLz+ybIsO82K3uUJee3tL1CDTsf/ztcGebhxeJGibNS93AioTHtCk
ihZADoU5i4IS74yVQMJlZVuX7lB05Xps2WwI5YUkKFCxpGi3GlnKi5aagFIPSrOaVyLAGNSnWGpd
ZV8kgAsLIb19hxGXWD/oCDnD/buCuLVMQQKgC4A+Pzi/kfela13YJtzlmNSndIPysXX7xeYCr8Mj
T+NziAxM6MJDQgmMiqlbxgV/frc9sVC6z6vqobsOnN9g69qubUrtUsle7IGgzp/xT0tI3EwF8zuB
3NsoUq4xvkVva46me14UZKh02ZufrEqwvjG/dJpoF/fmX1XQYwiHz7x9GQY4THCb4jUjO9TxBED8
gikPGcvT5jf945vhbrUJ6UdeOyWc18HpeSieRDz6kNp7eqAfVfpVhMPLKCN5xjrO2ZOCPoJmU//g
MCofx064gGJ/6FvlzPIE5gfZeyXshyjdXAfCnIuvGaMBcmdwfseDfDadY+OH5AsRu0KjsZtcA1zQ
gIiOkXBg40H/n21TAj29C9iDDO2oQDaLhgCMAUPeePEH1Scpgud59fvDx55QZMD/NMhU2H8WvAwU
mtJDNtvZFrIrBPc2yFDWTsEuiiQIfRQ+Ft8tVZZ2dKLunCkZXdMZe3BuwolTmIb77x9TYqZxQu2n
tPagzE7f3a+JL8s62RrwFj1O+1omPHs1Tcrncgpcx//frGugn4NXzsphmCjwaOBMG+jmXupnoJ0+
+DWwJ0/UR3ZXyvSj/WKeOZ58UNzbMQJTmumti0uausAfimDoTSrct3+NThMb0sEu7YqEZtNtupbD
gXarODJmsClcGsyXxaOGxzPRuIZpV25NFv5smNVwRfj+vnJHNd+X9qSxlPkAgKhSGqCamXO5C7fU
aYou8UhlJMbgfoMOCUcddWg5kt7PVcDojkuB+yySKWkIOTQu5dTs4ZjCwX+RAJJeGIzFtWONl9GL
KIU9n7lt9h2PNEI7yetgAhHjJio6+teOvGA3btV+jCzlW/TUNYMShyCuuIqp7TB+g2dPJ6IIOBgY
Db4xvvV25trv28qELAs1Ppwva5OUqmdoLjt7RpwliECS5oBqV+zBkSQpOyZx1kWOswComHTT4TJZ
MPXHjorkVl/e08cVkqN7KbZ93AsxAg+4WtgYdpvGN4OuKutUA4VW8XagxHHM9jbYpfKt5JIDONFL
X/c7NEoFTTCqAaM+crdfKpAsGTnKi09WSfmCuYKeJVbaj0JupA8HteAQfUHRgtb64cdshptND+p6
hW7SeMAQm+9XfQKbZBhrc8EYyG/Vp+V3P8l+ymhFTV4uDqklvzWJkIMSnB9Bqo8c4CQsLtRWTe8W
z7yOmZV0X1UOEQ8pSzog4ZnT2zhieHn9pms4GRb7gsA6urmJEVGgdIGnXSJxDX4dWVNR2Gxg1Rka
lwFrrALYPTHOqs500RIch3ZrkUE+BDFUcUUUoSbrpnWpYuWf6msVoXWRHh/q/G4yjJXdInxQVlDQ
Vz5kEB8mh3tUOrMdjkTB/hNe4N3AUR0Bnnrp1gxQ8CYJmblopp5NvD5RjZZbHCLJvu57MJ1m5Ge6
ZWpZ2whs0QX1vTAtKZSq3WGYcx1psfYGL6qlBtgF4nX4b+8BNAp5sGZcQQtVe4Dgm69tzhltjSlW
uXPkTKFJE9HjCZwBg4+T6nPLs4g2d1CTyBdr8ZkAn8Lx+6sOdxAu/hPtS8Z+L+KM9G5YWlK0BYd/
toVOSSCfkskzS+IRcn673bgv8E9ZngDICGvbs5iarubjBoYBg/DIF5SXF6UJLPFoKi/6eFATVDWt
SaVW+q8wQFumHnJ8fLnyne54z3ad8csOwYwTsFWORBrwruaedMGGZfLxLjpTsoFqzfHifbGtiHgj
oBe8IaIASFQMLrDDcGP0hHVhTGCUxlEPG5x399TdPNYlck+s020uw4X0rbA/yNCYtTme15660oIG
iNgytcdnnx0CQCvy5FZpssCmcLp0iA4EgiaDfSDv+hmjp6OEn74gxODecHPUYIQwTgTjNnLcgKt9
hGcdzmtiiNtWbCgOYHvBYkuYdzSWjoO4Tqr1degFp+J3lKfHFw5zM0KSaROi/yLVNs86YM4b7Npq
sG/Ws+81uuGYToGXpZNrzvzfHKJsJoNg/Kj2fBDpk2iPZVesXMwTDUPrPQD9ZSLor3OrpOmc2rZq
3nkhJAG1vexEqC7D5L/b4z98gAcjm8H6RpO9n/GbBrgCSJXZdbpZFLEqa4+Xcao/It7WbkA7K/X0
EgUWgxnk7DHQQ4VevtTBV4J+q35d6CITUbChIgmmX9crX1C4a+hojkCbj1TZUUPD+uyUQMFq/PR6
tT5Y3IP9x9aswPCsv1P8KacoxoCzu8D/d6Dm3m0VEVQYrKlF03fj7aUUBzy9shp0ay7Gs61Aq22A
noS6xKYJbxkr81fEXf3MpIgdqMy2HVy6Mbp6lboDnQQkv1FbXPEH+9et/IaDsjtTB0YxmT7OgY9Q
EC0YlAawVFZ5pxzg6ttseXRKHSpGmeEtYpCkt850Km+X7qc1DvJnrPHu/5fnfXsSrNnZmQBa1xhI
X6Cq7vUf5xx+5/2uZY7tuzJMchtC4l/btw/BqQJJ4sRz3NJnIr2/JopX6ZC0MCneCebuDQuFH42Z
e0S86ig/42BxixWfOZ+WNA0XcR7V4udLXJ1gAXg3GsLrvGuT43am1QrL2EjQOfJCt3/wK0E7Znsv
ya8SopnENHUZ9QZimQqOL/8BjvshDvNKEVDXwCLu8IOGjFNmNIWFk81q0/nHAlFIVCQO2x6vpna4
/VyOFtSuGAdPKmjSA0LyAQpsBn/r/e0U4pSkQio5Q+bBlIKdAWfa019+adEFd4KuRNmpUU8faPs8
6hhf6ioIAhA4opvWk0poyFXSBKieGDzQt6IMgGGJA0XTugs8/haYf8HwHrt0ceOQeVLo3ZiXrwIw
W9c4OFiAHfROgb2Eao51JutlA/z5rryIGuh5WYpNcXqtgyDbMyAR+m5UlxXjPk+ksxZxo7mxHI0E
fWBN8gFeL7tErZD4ha724zQ2GF400X/zy847e5jiOri+/sSAwderRdjqN+Zqq/bM+02d5cAnp8P8
w73cEx4Rd0L0Ho3QrRZqvGxCgMRtW4Hy6cXpmFiC5YTD+1cGxEPy+lhtDlgTvtz/uT0QMcxwTIln
WaGys+/OTgBqoQhGWHsOAs39BS74bpInaY7hMKGa0aRHsHleBRJmIetMN+rzQIyjnjuAz0eLcm1i
5Ro3xPvxIN6Ss6dzUCRZzRdaK0NOSRWkP9cBRuNBdlHRs0rocwfx+MmQBudDe6clH1CIxH/au67k
D8hJPCHTM0SzBD6dxwwrLDYBZkfcxOa7BUSV5rC5R+3MoG3v7+gyUx/kgEwfrmujpFymJ3Fs+CYZ
eXE7agnyptSSvPrItSR2mHWilpEpC0FuLKCGAWS7IJHSWJsLOqrju/mbULv99NnijtR6GUpOF4Wy
li7oTMmPG9TWxL+vOS1JZTVc77riT3lH4TKJXSvTKfQvnx1gKe74eGB9wlSGuITN75eefaGbw899
m/mwu7x+CHdpCmGiXN2Cv6ZKBY2oQu480/V8bTOWdslEHM9tEQdWyxSTJPjWXVzEGI1CkqmXhh4C
+KsYyP0dm0O4BGnS1yUA2TWEEuSI0NTD37bT2CXJL8165E8SLcEUUtfOo88Jq1+Asf3lk6yaHD5d
lIpWlbsXKugExy44tdf/N6p3CaeqoF8w8qpBUIrx70vmNtGKwcVM2vPMCKkQ5GNdgQAjnpy5kXEC
W3mX7bKDA+nJNXcUDS1Q7bTLAMq+aWUrLHKXuU3r2Skj/z2wqP0mseWIfUO0EpJQkgpPVCmIlGzO
5wTGKCaqJKDiU+ZgTNuNjLgpTbiG7q5Dv7THZEQ0UtPJE46M//IjxoU+k4q/t60heemu8Q3u5m2J
uI5IIv/oojZ37xPBURJQF5fWNHfbOnCWMOLVKrhwLQu+3kgqYvLyxeU+aRTgGDBRL/UiGC9DpndU
a/z3qcYB7fhDjNN44gyT3GqSl+G1vXba9feg2XFBcaLdDF8KarOX4uRhSWze+OLHZQ9h5Cve+YD1
fTrNMkmLreEn/uhLU6Dd7HmAeqLRj6avWs8ykpwazYuh8dzkZF1UYBgRb1sg7Hxq0ai1XYe2QfGv
dW4tvhv+r7ewDwZkBQRdcFK0Kcne8gVPuJt4nS9cpYW1HJKde+UU+7UW7YVrn3GkYKLXuBpYdgl6
jZVrWIaSMD+fC/3KZ11thgW1MQc8hk7KN+l6k2/e1zkJP59otAsEgyIDaTL5V1kbYWN61x0bWFD1
fEXX8Wia/YHQQ2xkZj6mvVSBhHO9aIF5fD4KYSYL8F6+HB5JdgMME/5vuGDuuRed/XCyONUItp3k
+Hd6aFvR9WvPRtSamvksI7Ji1HUDLB2OQ8WIdiNUUqKd7EwIUNuRA+1ZA8TDSAaSA1OYgbo4ZKcO
6+soE0CpBS62FLfTYK54+cORWOCWLSMxu5evpZdy00b/Op19MyvQOfg/4fgZcheHlef+fVhfQvKf
OLGmfBe3kwFdIKNw8nzAqlbe4eSzFAPwQn9lisv/cSOzfvORZ8KqiEQNYNbFW2ZykB4bp/JpPYoD
lT9JdyBq/RL4PdjoiB2KA2sCftQmYBV2pGvuUrxhUgV/IH19ivRTNznkP6+or+kS2aqJvrkU7EbT
K2zO6KoWlGQf0UYhb6b8pDykcdcHA3+KVaAPhpIFuRBUK5AQ5eqmcEBJdj7i0Clyr6mNeJPqoxK5
ERJe9oaGG75mgD8R0TJw3wsQ7bDE3OFka8/KdWXPoSoslpqLl3RbUQnLgJ4n+J0CMkJXvyNKE6Lz
HH3VseKFpho+UuqyVGS3eWso8UsabgwKpTqoqe1boXFLHkELD12dFehcmp7uXt5MRV+plDmstZQA
RNAGYibiuCXiCCF4Cp3JGgAKPaDsDUR5TYZX44v2QsFQSFMmf6YhJTigzOPOqrpdyW4KLK6VwH+Z
mUjhs/4t7t8SK3WZRL24dZXRDOTtsC5HngmBLYqZqrlg9BqMfq8AxobcETF1FjO+RwYePkyr//DV
PKWiO50GypFw+wWPxnPM7V6O3Pf5SnEuTVW+l5I3pFnDzpGfSnmfe6Kd7hC+bEk52wQOoOOhCUAj
oMAEnp+7nGiTyD9y6+hzhxSc+3KdQfRwJY5/PkAb56J6RC/zebkzpKQ0LW0GhxRGa1HHgLthKEqH
FMfBxHB0ZKK1HGAuRwlilwivuQaCj+n7DFYHgL1cw9VuGbPnOu2eCWwDnRL3r6aNpwhMPuF/HXpX
b4u8ZRKtYm2yvAUlhzcf6MIBI1TK6ikMPHpfq2A+afhGNMnPkmpIHC+N4l0bDYsn4b4hu+WpR5K2
RtBstf0d+PSeDVpLGLIe5TBCfAU0FBnjULzhC1ut8UYMmNEBvyWoJ1IfjG3P9e1vg5FsfCrqjWce
os/nhBKlYKsrSeHsy3/HVwW1/rxNkLZF4bhXBPZoS2Rm9Z4DZtRl0gzPiAL5ndzqS5Jv8EGITUvo
XHMu+j4zQ/tlFI7BCwghBE0dsxoelgNxnKe5r+ruLhGJ1yOq+4qqzLjIpjOrxu0l0AeEK8cv9EYU
3srMxGq/imw6BOHOzE1I/CqkejOg9fb8NGmxK37iOq7DMS/t+kL3UNPR6RfQCkTjS72/qvi0SxRy
uwyCqdat7b6UVSyNNra00L9Fe2gnBUjIjGOsHS0G8NugM3dI4ST/JUP8oDrZCOk898vAIpoWmXPA
vW2Pvy0RqtkkUBCr/GEA07lIypjAUtGpLHbwHZbyzVGlYPo129MCXgEm/NHT1ta+hhdw3Shj/unH
bK6SMQcCnYf6+1XKcIzfFKEdSyAdMlLlqA7tLIzY56dls2yAYWS1JKQDWap6skeQEY+Ws2Pk57bC
7D65/VHkW4fUkpwTQjYKeTSgMWORPnSLZiuiqMjq87oUQBf1FaIxh+i4BlXGFkhyKynUKVhoVlXy
T0lx5lm2bgCQw0TD0y8sAom+2btWc5Vv9tOA/5AYX2PRsD7CQcEsPZd0ta0fxN0pMAgoD4owm+XI
FMaS6azUkvbSI0hV6x0+wwp5a+VavA601ME5UFya5oTyAj7T4BlL9uaJEsiePcSBHJUv3MIf7OkJ
yjwgNuKT9Pj7eMXzy2rz6F7fHNdTYit4LKUBEm11mFrIbKxRBRGGF0CwmIUOPbH1z8H1ZykPCLUU
mgVwGKipp22kp0au5uxXDRwt4VbbSdpHF16Wi4Y8lHGADQxjG9M30JGVXRfBkk6WvpI3a11OK+xZ
fziAz6iyKg8M5u3BIDlZ43fL/Vxq5WI5ZPMBdTd8LYLAFpf6J18to6OkccqDOWwyofQG8vxBtp67
aSRwot3WWRDvVSSk0CcUPCxdi/s5ZCpx+G8hL/MkObBphDv+D3OrUO34EX0lZG2E+kL5tUi3N73S
jcjKC+ScMwduwCe9XvZvKuWNVtOczy2UchDh6yvn+kNqoMZGGwYaG1M5FaNwgbLUxZfsuvwQ9EKr
xMDpuyVMomkgbmamuhaTEWwPqYP464XOap7CxMFRRs3puM/wB1+L7Hjvv1JQGezWpp/WmDjBfVoZ
SxW9dL1IZWP5bqnjHGQm4k/rtIl2g95BNLy9DIxs6PyhwTeH8UVqc33bJAzbQyPM7rO5MChIpKYv
qCJRvb5qlVLGyRoXuje+rY924rAnRFyoZlVrckWQurDKMxg2s88EoWPt0SH+JSQwucuE1YJArfik
RB/icX0k6yxrrNRc7ODWdKNvHsb9cUAei18BQv+6X8835PRaqi5RS/2j7Cd2iAfpTOEmMxzcC9Q+
BSpLwGJdCelbXr6oMxV2KLheq1wB8gD/4DR7neJyQLZz8Ghtj9qFFS0MoCKNW9xIqFNFpqOEFEGm
2LPsDlNrb59rD5aUabCPlL5T9FI8lzIhsLPGgWuDRJ2Np+XjPOJbFmgyNBUoGV4z5guroByLDxRX
tOQpDN1zzq7qKqYLeVvo607SeG7vzglIjpAwX33MyQIaTaj613PRkHhRXKCgZ2zhLEjSahFtrYPs
iu9znvRNQzmf6pYpl4DZT0s3cJwkTAb5tS7bo+8BV/2gM2lCCdgfnIuoJrutHZhjN7A18j7IxCVC
IiGxnloRyCHsCBD22IUfVrn8bm7jw7+y4HcYgul66Y6zFJIVki9+z42tC/v7qrTn5mwhgSS0twX6
5vI2kS5pIK4i3xw8JEv/sKx86lNXOjKW8MSv1u/VcW8/HoyO6stpMYGnMfk2bc+64HXVr8BUnQCC
pG/ln+KhCMoidxn+uMzYVnnWmMz8R7Es6yPATlcR7v+ynP6yerEUVxZTUL4jSHp5/AtkMWpJy3P9
T222T6Yo6A7dWpWY5ZMkrnDlHExR6oI/WIBXE/ujSkiTMdBNX1wrzR01XCfHJ6TaCHKFA/RsqzRH
UjP6qFMX1zB+4D/FpRF8oDDwOZ0UXiDxh8ANj1ZEbguByjindKgvK9uyHZmiLlMXUueqNeYMkQ9m
O8GD7Du0RZmlU/fRsWZi7RW4XzYjbFWLXFsJm2MJft35TcicI7XXk/wSPbwqeM8GjGMpJflQJuSp
ycZyr4BYrjLkm6ZZ61XbfsKnlMzD3KQ7XlP97j575w+ueTyFTdhgtK+h0TEhWUzPOaPNAl6MkTPt
INKZC69lQrndJZQ6mN2xb1Zows8c0e/V8DXpLsuf/3RiML5+1OZR9+/+rG9iklJoGCj9tUSOpkyg
bh46zk3J1cQGlpzDqe/S2+coHmjRXPMqflD7Ypv3c2ktqXCn9K41dBB7+Wvo8CgYEPkVQjSnH+cA
ciW5I76otO6X7Z8/+HqsAq9I9YEFBUUfSaSkGkYcpA386JON7Shd91GcKw962YqaFu+Hthr8rd1S
zGBkloIAU2r8US6O8VYnAOJmj55yKEaYWZDgwCAKubUZg5su1jZBG4N6ynSYz/oSQlHNdZAlaipx
0yS4mHrIhlpuprlI/sogu0k0RvD+uLTJltWG9pboqffDQ2R+4f++VW0aREgK+kjLe7Frp1B35saZ
BIVo/0gpMHVKKH12wMDsGRY0M2k5Ier7k8R1ABumfOdSfPip9y1HITv1iRlymftijpclWVBiRGhN
zf1qGKleNbCyOSkXyhHeRUuAFD6/Zl/7CCSZTq7I6yN7FqIHB0fsT00JCdU5+DS/SPIq0NZ27mzQ
t+ThQOZfY5lm4/BknxEzsSdz7dHVA+2yky2CIVubqzlAbDS3IFcnR1EW4x13AwRzJTrFnNjA+S9m
ZpGBZI3+hhoLYLDubkVBfm0873TgZIMTL3rjgGRdKZ/8M9m+aGsZSqy+tiJbd23WhTlTUbK5UPGT
uG4mNUw2XM4nN/qb3wTKWb+F/B2H25VEDRj/FNAR0n7IDGoiPTGOWMyGSYFZSd9X40VfGqsF5MaX
umo6Lmf+SEjm8NKgr7Ssxf98VQP28OeU9J8zIcSFjLpMNQaKeDi0NWdarYn3a4GJX3PFhiSpwrpx
5CDXu97kXMw9EYfIJiNITbNGd2Jh4dU52nTf/WixiMDAc/TNnC0+LYGhs4yROfwp9SlFDT5riE0p
hRrAhE1ddhz7AEeg2G/cOh+IH9jQMqVTMks2lAtkjmcPiPSz/eYgqABc1QRlWAUU5eo8l4WcJYle
uvZwqy94OzmF4Ihh+zwBgLjiJyjLt652U2Wyk9C/Bf27iY4AAH1JkpiH7jG72c8ogYOh7RU3j8I8
+a3RWQ6sSK2PPw+8ZdGx+/d6NLYgIobTJnq1LVGamYjWQi/2MxBb3HAFUE+NQ5AC8+f7fuNEXtpT
L55d3mQewhKTdtyrSOxsfOoKyKXG9VOLxa7bsd1yLtzFI6BE0iKTmMBh0c896e6gMa8jmMy7p+sJ
Iilv9iE/3j2zfcGCWwthHXv2vMH8QCM6DRtxQGnEJuiq7Ng/CPFg2cLvgKBtAAOIJ2wFuSRJp/mm
H1fLD1CWLh1NSlEzwRGmzlsHCpMGSOZ607zWqKa8tRQ2WB4nfmfyzvDkKK2nx5ANQNUryHaB4bhC
3RjfSOsmxSiryaH/vZxtY221IVvLI5ZGIxYSZTQ43j0LrvbEldjJ7CXR8Bd+JQiv8Z2uhT8uWzdz
X9Cnc6+EEBV4ZDZsovId4MksPg11cpZlF+Qg1jdbvl9xOQZ9V8sDmQ9BDRTEgDlN1I9qeOkz9Hgf
iYHLgh1hSEAfTPeSou2RRnaLdHq8mPpYJKYqnsS/083HZ+D5RKxTf+mXabQZuPw8b7g3Su6sfflu
/nVQgzTc2DXwbshvfcHk4kTAoA+f5x0pZGXONjB1SHDUiUIqjjptTIhjNKoQcpYUr9/K0frsyb4S
FBxChJZyLuRilW6ynWnUZp7WPRA9Y5scA6haKDqnFRASYNYBAtuhEm5MmmmWP2FriPu+WrVx6xZz
jVaGcPCsS9Y1oLmVsU9uJGQq1pjQxwkjkk4FPe8WPxlcvnOtKEngeDAaL8dkMAy1F33hhcqf16jC
bGSqJpFKzloA6PhaY5vIQvFuGz89NJU7yW59etfv2pcq6gcrCxFbrdmEYrqcpKPZMkgB5spfb/i0
wv2ccuAAfFPmQvbonVvq3C0Y/2pzjSoPKyT98xlJTZrbUKi9RONmQBXwRIJnotkPP8XkVYD5hPJH
XucYaBeDA0VdD//HLjiSJyBbsQxSn3ZBFMFoLkckP0TkLF2MdeuO2DrtMmJRZJeAfTtBIg+SZYK0
UGyOhnYSPFOlW0KEWXbmTaqA3o7AEIv/TPNaNBwbxL7cPifVaN5w62v4hl7Dy20ipy2vu0m1F1In
tVwnaZfc8ler0g5q6GqNg+zt8SrOivRaNeKTWsHuTmfiu+3aEjMRCYwa2yTsIGEVd8tin6nZJfUM
HMbEfJpq0Oobin8W1D87JYVKoiDrpBunneE9PO7F+Pw6WXjMCaaJGinw1V4AyscDBq28dGGCBUnF
Ym+RYpcQ8LBlSLjihAB0ElyebcUrvTaMrxFsFGv5hm6tkzyqdoS8hSSZTC6PC7vI7sgj56OCkiTs
yDWHYr9yZx0vFXAJyvNNPnucqYEMK/x14lV3dE7emJXLwx/XmPqrYw7VZCv29kzZBsiAExePMxc7
ZkYnBwNbExybfsj77CdJIecEamuFrRV6WfFn67No0SPBny9ZoRUNMgv9ZttPmPtszFH8wG5ImWap
hlWI2z5EKenWXWYEpBjEb1PF27ml5DiLzu2bTJoafs8Eh/GGNvxU+iQ8FpKCWCuLMLxK9znpizY0
COsNMu91x7/okiwRyxHDErFY2tZpcN2VCi3FFtjZgj70xFBifRTziCn0wwdBRJm/T2vN2bhremJL
iYXtJRM/yIuSUkHHIrUY3t8BoVQ4BQshrODuG4rdBcMXtbz+JZ208iWuaoLKbZF3S3Kum/0p2hGz
+VZFDk2+m6C5CGqx//xc8eY3t3whZzpJYrliSqpp41aWzK/1d5dE9u1ETio69UcB7VKw4hE27dMk
jcrpkwW2XS2flzMJ+oBz6dPQpE61aQ80SLrC6SKh4VrcqbGjWEmnXOFdW3cY39T+bWxxW9pcoTzT
OLKYl0I8lnL0y+CFByI0kS00F07Z6Tr3Nyx31v4/NzH0fTDTXdfZW4bTeLmrdDxAAHh+TBtTJSs8
9yqs0YRCyNpBgNVYW/O5ssK/d/3ePTl4XE5+4hPSw9I1EbShojvsl2lUqjGjIddjcntHx5qq5xHp
YYhK1h4JoEJVP3crATgs92vcKiOkPeUuo7rGMpf0IEHvsbM59E4Kymn5RZoh+umq0NKXBaP+Xx00
xAJVkyAjfVpegMR5mqmgTttWaFHfYVsVUce8uLtQdjx0fctzuAXXeldBK1v7D7AAv2qnLG2coQoE
9m+s6Kml5w5S9xh38SJj1KvqDMeNau4bhvAv5ZNo4Z3AWFE0q8K3EzcfvljiK4yuZ+BkzvFqRZfY
xN1YkW/jog1V33OTNrrbVEl3HBEnhi+kWQFj5m2pvF91E/jKxBzWhD9VIZPQ8E1fo6lopacdPpKd
EFQohMr77Vbqu/Y6jY5SjuFwt0xYpqYioWua1vsNSomAOW5dPCVTzMEgQtkS00mxmyBUPkcsXCOR
08fyotieNGZara+kiY8xvgX1llLdbtqQWqUjYSbGOVw01awcMc7m5+ccg4OcZKk58iTO/ZU+o55F
/UFlD1+ctqpXzn0oaDkaMpa/StHbIIx7EFKw/huHu0ETTiB1Ya+Bz+rKPX1EImBcJADofa/d9396
zzp/+Iz81au+v4xNbUyFw2g+5PcBX3HYBOOqwMHsCet5Md04QP1Ma/MC66JG3KPadL4cgiYMRttG
4BQtaJ7/dPejwqfK7b3XnMF6Wh+C+ozbj8uDEGGYrZ666L59dm5KGe5fF971jiqD7pkGKg/4RSI2
MR/pyKWBDxibp6e1Xv78IzRLiRgRq3rJ33TeF7JjhYg73WKOZfAWKYGNp8PYmMwdkbR3oLIoeKNJ
u5OvZlBhQdwKNjRc1G1bfwrQF0ozDuz18sAhOaK9CiYbBiMwWVNqsw+z0HYTMzEMhiBdH8kXFrnk
EvzK8VoN1QfiN9nhwwQ0F0+tQ2a50/quJlS1dN1STnnslNntxO89JAYpmnFBH0NzUDBTE00dJsP3
DwT/hNP7J8pSnzWXo81eq0j3noPfpXFvMi0LKpyW/xzwkG+LsbMVqS30Aj/uIpV4TffzApjl9yJk
Thh9oZNyWLcflIV1RDVKCNyK4vK8tA1HaPUBa55W6twKDw5sH5XhUqiz+aC04kIy0eFfBlx9viot
YsPQ9GFvsnmdNrigCS4MnxyKCsIBLi+60EuEbvQrM2ZtfVm3LfRif0FRjSQplaBf03vQ3+gAi5cQ
Mn/gkRygJBpWm+ZY+DaI6OKFPsfYtI4VSZcqzc4irDMwgxB03kQyxFHSeSCT0Uu35uaprK0lmHiH
nAvSqDKC8v+NhUa01xh5k9zMjBRS4ImMcINblTk6gfXpYOyqwGuCbCNAl8OUnEJVQUthQANrSBau
NO/YZPTlqWIJMWVysAxStRpZnq2K36cBNLzNREsrxMFg5HwZb7hMeL/55g71E10O8OAuc8mVTUKD
bvn23o2ic/CvyL1rYFCcwIMkPqlYczZNQ7bQGrl1Gyaj3c/3nieAE2g5XtHWvN1t/grIL2pKRCNF
mTYg+hm/QydIcWDd3LQFtAZakB0kIU2/6vwB0raLVS9SsRUOKXdhPXLhe+/TN3pfJqABSb3s4o9w
TsNAgtBsKtmkWY78bT1pcVqX4qhso+qp0g+f85WN1gBWRqeeGP94HNA94S2SAJpLB/Fy+LTuKpQx
gFh4KZbWA7kRbH4j5VXnXq4qNtAtmkEdpIs4kADKSJ2MbCCkpr5ICRAv2pYpovbVP1gZ127AajqT
AG826xDr+Ms9DVb988e06LomcqTA5WfXCV02A2fMh4dqY/6uw62HxbqwdtzBhXYf26yOD+h0RjFh
Jh9btcW1pAUf1Q8hG0yvFUx35OyGgSHejgA5hTZ7QkZxattMhVSIsYky9WVFY3YQ7fgxFLncIc27
sVwBXotXFg2ipIuVgrXIDwHYEhBZnI2rKSc3rhu/cuxVopaKqtOU0C0p+jAue5U5Enym3fb6oIZC
kRo8zRDdrUztEtfg/zDybpmAiSf+FZCpF2jK1jDdnEWJxtW7s4tpjJ6XjqioIfPBqZBzfWN3SbeS
j+NlsKYzR/jmtw0Ht3AQ1bvHwjorFD/2uMwtIVWHQGWYk2Hk7A7b5qAgRvsRhFG2HNQi7xdKkeH1
zKoaX1J7by9jFtklFKX4w9ru9LrlBobDDvlo1/96Btcjt5pxGUqGATrmFO3xazuVTBhrQ2/gidge
+cIYphbJEkNYosUKRmzI2mm3WsaZbYO7EV4DjoCvr1h9Z6bC45XN424DFXn5WQd45oq9QDOO+Evp
9oe51HqcaCzQNevns4IBZOVDf/nrEPjgPrywhy6DDjEoc2EWzS2yFrwIMe0vanLosTUpmZ9lvaq1
npUlKxuqyoCF++zX+Hg+aEuvKTMD+ynJrmz1rrc9sSspCeq0q+b6ujIAPbw/MbN1wVDJJbrw8bLH
oCms9rHW5GOb2iFOjRRXBSO7SvRhJmbmzbi/0V2TWtr0RYTG4NGWYLqK/NE/YkXkbk4KBMmGKzRB
J8aBDRiIzid5UxOcIBcJv1wq/aSM4GkoD+FkgPsCfCUOnkmgkaglfz43nOkCR+O8ARCDifd51Khy
yYwQisUFTf2PHhgRshiI6e38ST0uiGN8Lyfmbwsv4BqBFZT1UqKZ1KtU2IT0C/CUYVmMI0ocheTB
PJgqjEeB4rNgKigw5GOJfuU0wFk4fizrJKpYXOSLm86Qa8uuJDOaiSm06WlmMbgQs9h98NVM25u0
xX+P6vByGTXeZS2saaBcLR6MLa+d8aZGUpBIqwwKJqWttJLfPnTlk2A5OWbFxwbaU8KOPznYfFYP
pT6hfnYc0EDrTK2Vsi8nCQDrleNt8nlcegXsmLjF9zr7wYdtTXME21yxD8SYuVg5YYDr1ScUdyaJ
+NUCs35+KLwZlyHmzxM6A5FjTgecW2OJPAIQL54CKvZvJqfWAKpNkXrMoSVyLWpy9aZtNcDETyGB
Gb3zNIlyQmFCURYLSDyAhgUF4rpaFLQur+us8BKllL7psW5czQGkNxZmxHsVewihyOD8caJbkkiX
aWSdBJk20k0dgyWPh0CvXOD1t6qx2kwa36bI5cCKRDLvDgWUtqzzNiy1yAZr4bghqioqIYc/dBcJ
uOafCUksFoiKNwyJsJK2D4uL/dyCMAysvZ3V0dMkjHplV8QHj7zGypUt1CYJtnWnuq38qpBHjrEA
WnKAyYfi/iBW5mAXY9upWFZetKG/610DpPVFoigyZUxyvkwCMKmC32qPGx2+sT1/xXqFb12CCPlv
dgY4dpQlobmPwmcppFRJcOFPKCw+qFiw4mkINS4pgL2A+t0rypZsdB7/569G7rEzdvWM7VGuGco5
4z9Rt/Ah44sHB4XdDraU7d15S5Kocbs8/lyGJ0XLoVj4N8dkcMpeTSsu9C8ixadZZ8AGX7k6vsPE
XD4vny1wYlk6OvnHLFFnPPRMWIdz2CLNF95Bt6H4ALcCZCr+JSf0r2Y4aqRx0F6KOM9W6tBYtcC5
grulAJoeH7vgwNXsP7XBGU0LNfnvPgk4tsKpNygVvHKvDaNqa2sTOWZl4IFg3wXR0HRXDFVLbHSl
cqGhJRz+UCs1zn1RDBIYMVglAAQslUvNJfzxmOo3UdlUdGhJuwQrvP7pdmKK+bCAuC0apPlqss0q
gHMcuQYTVlM5k6AhZyqRsG8e0Uv17If7aMZId/4PSToUVk0Tb7TdgQqlKFsSFYWjKfQBFghTCsqy
kNdrjoD78952vs3Wdw7HHIOi0YayldwbpC3Oco5kHH5qGU4BqgE7p7cH/z28guKDprFBjTIy4A7p
FcAuby/T4fE7f/MRFHiJFSHxNOSrkenrPThABrfLb7Y/z/p9g5DPjkFaobtwh4vElj9PLAHcx71y
g6An8ZQDYpS5voMMOlMo+Wub35TJFmG1xKLObGT4xtOD4GzVD8KI1EcQzMb9QzzzviH/ys/nHDiA
+l+B4sULnc9r0wHsviF9wgjf1XNU2USXhTVB/LvXnmB9UQHbfGm4j+S/DjtUlVirJxOsWTSIIHdY
2vWSrglTeUoQFdpAXXJ8NmxwNHvKwE6NCFJTaEsYTZ27zqlOVPpwRJWq/SaYPw9lPH+vR31bo2Wj
1POrlf0Tr14wwDHu8VjKHta1WgozIc0bqwAPachoi7xUCsIVZlO+GBfocCs5PVeu2b/KRptaW457
8XK/Kd5Hi+F6coQtK+Qqoe5tQf20QHo6zLSkzIjXyCdlHyjJyYln0H9XNQmxEGcxaufpFDuotDII
Gg3PmmJcmX4hBIIPbJj83v/xMPvwg/A/jYNVbm5mX5B1OkZ5UIX9kDQuYGYSFbtkFPwtDyc62uMa
9pDwKRPt21s66w9/tsBke+MP0HphmI2+ai6AKMqK8+cDpR6EurndxDmbO7/x+O+LbdyGWQNHk5JU
OVeFw5MvuPb5akyotxn/pEitlCequhR3TQb4FDB2Ic7sZ3GR9HKzwk+1lUNwwXNLFFTgxrLQ4MYE
iKB2jypMvVIcbNj7AW4qCbJqC5qpG45+ZbUYCR9LwzJ2p9Hmeoct49Fb1bNX5SsK8K9xiHywxIfD
0TtBpraqfx8t233Gl4NY9SYZdWPIzo6ukhTkvDK5XBxoPQCI5JNyng6fmTu9TUTth+lJC475PKTP
BZ8aUONAeaXDdrV33W/LFADAr8CnAyPLnGWI1OZbk460axb7+k7ESKUNJB3+XpFKdN5Zp9EJuzUF
qmWzpCgBnKEN3hJV5hEpF0joyr9wDI6oRKOoy2A+Da7W4yPTnWAPRCEzdM11K7aTrtegxjS3YUSc
b4nlCj5QdXxViri1/BD2maaQPwJEuAyisZX/E9OIO3Rnc2zO9gJvWARP3eqIstr9wwA3pz7NsnLD
zuFoDFnMWqQ+SFjOETR9f+22iP1hcEbPzxwKnOfM3XmdnWHewK6rlGlFDZh3dymCBVJ9sbc0o67m
a6ZvBbh9MrZ6Lp44rg26G1xLg/W4SKwFAaImEsN2Ph0clYWyXBm1C1FwX/lUhou+QKh+soZn/t4G
YT9Qc9W1WNIbrZ6JQOpXqM2tombpu5JfGQNMUchQLEZ2I6j6oCDMP+SHlES7cNnyfu8pAeOK2lHO
se6L4oLAzMSHGiN/4zwVNyI8NKzwczJCi9fbu2NXVvlC57qFC3A2hJG9qWKLw/vyDSfb1QSY9tV5
Jna+hH2C4/PJELm4+ksJUi4xxEoTX9KgWOKpvkLhrukQU+PBgYqlmbQUYYl/F09mfQ449sYlKVpL
o+O80O37pQjC0baqz6sgtmRUoMy3IoPJis4l6osx2vz4U0s4pSFkyzd5eKD+RZSIHIl9K/qLew7L
yp9z7xPZTVjpiLrz6We/Vx5TpnDTyB/OdsdXJkczNMprYmiGRP7fVTTDi1W0V6WyRJH5vg3cb8S/
AM+q6p4qZpmKPi5lf4USUkYltowsuf2hno8NvExmCRNRtIXm6JKECTSQjcNviD09soOORnySlAee
TTT1L4u6HW0EFF9AvksGQpUnpFu31uVRSlYARoioNyMI6JEwVPQ33IpIxS1TXIkKxIZceMVJ84Jf
adH4FTTbIzsNxmtScLfPrwXYYSqfTFEbeZRAvPCCSNm/d2q+6Dr40OqhYxnMcaMYfY7anQQT9lvL
YUGwIEYpdjM0P35+c/mQ57SEZtFI5AvYAhEPfMpznEQpZnlGuI06BB6hiSuek+F7fcC77vTURRuu
FKorJYjgIFkeSlAWOE7iTt1qLkm1fsAvMhHKOaRffAKGCAuwv0udQbDL8PJbCAm2Jpc73CUGrXuE
+JT63Sfcc7hEbYeMWdNIpSmlGtqA32YAwjAsD0+ffjrj8JZrb+qfLAWsQadJRLlnkJxvvQk+VyCC
L+PeSnsB+f5kjf6lqW43G6ztj9YZSXLt1u/BRXXqypFdxtXhFNypZEDFIoulsgPYNJ0ASo2Rart+
mujx+MpctFVwBm6vbn0fGsZDzGZDjTU2G5pLNoS30wKj4FN4VYHHJ7cMZKkHjdMa85yTDLhvLgsc
MCG3GFciMGvHB6UDVWqpzQAS8KDPysOX7G4XxCDtCjjjJ0a3EBm1OuXQlpHiVSadYtvJJFjqIoX3
YpVqe60CgnpB5tTwyJfIM6+5DFDLt29AiH+y0mO3kGgkuutWcbdXApIfgDYKpsprcuJV7BdRuj8v
6ZN6l4f3jn9txB179Z2lr/JplHYIGerWxAq4dIvCweU/YbKRPhOnO1Uus/2Y7y4NYxX/0mWmgbHJ
cCRLHWeLMs/bVYrQIn/rz4zSVNA0DHBTNBlWWvwqKo/Wmyrj6RZ0u8Pc9y+D+Bz/2qEMQZoAaTpy
g6wKAPtOoZqq3LMmljazKnJCVV212WgECWfaPBPQuMWcdmRIRm0m2ly703xZRjqbfMDVxPv9KdFz
AIZwDLxcLAtWHkqV131VU31BEyfg8RBbVaNkSEsDUPYtz2eTadX7qkTHcvyX7+hSiUaudViE6Iqg
vX7RROoC7QKYlfQ1r622ZhY67lu/MNSdQ7rhjiXrOq30PpUL19CzYNKSo+hXpKbUQl//FEhiAS7m
rC0LHL/fotvu0WapQcZ0yAgVODYDFHwxydGD4LBCzRQOvzGRjrj2HlT0voNa8qqfyB6Ga885dENx
fwIMo458FT5kyWgGbLstQ0m+C/qZNta1KCUVMHFKI7VLh+rzw9OP/hEJVpU00gwc2GPhP5afgkmz
mZLJ1WYbhO0nbJSf2NSrdmzp0hTEA50chJsIFQyC14VoeNgc4yhiphFJTbyp6kcl2f6hbH0Rzhla
K5LvKz22Ed5XGFmHpDpJjathfSmbtJtm1Pni6HxdZwZkInEmlIzmACnEBjbQkyMocMGFU2qkUbNE
/zGaY/vfiwsX1E+vdjYDhEHwbil4ilQ+iW0rQEWK9FN8BUt1lCSh0e5kpkI9+vXzXajcqmuYplvh
GLsUQmEyijJNN5F68KwAhViCSl4sZ19S2sLJtIzGdEAOUJysN8jxS/NZ0x91NLMcGROpfGk+1+66
Zw08yAUjPqXvREFWXySlSXmcbXLTDSgLnHEk7AtVn1PVbvz7ccbnu7e6QED7VZ/iVAHC63+eEtMx
Ac+kjWrgdqOdWQc9ut8AocWsPPgJyS+99K4FdriVWNJ8C2hi8wfelYHx1H/WT2XuacgYvmTg63l4
Kj8agPRqY+6VPq6cxv7jddBZR5WCxvLsVLf05ZmffS9LHAFiiPwIppWzT1m7rWn/3y1TnSZ7lFR7
+rKq2kFPpT6MvdPjTcEYzKJAM9OdrpSx56EpKGsBUtFLYvpDMzjUu8ESfmMYR2lqtvzhtTKPOH+K
GH2m3+orXpB9XFZfIY9EM2zdRf+2+FS+zJipXUDGTbLdVhHg4NnBJh+c+YmCUg7Oud/FCQkBfCWV
junc4/RKjSfL2cRc1AAPgeO3TZsvefPefE022/rQwHsPslpc1J0keWxEnSfg0zWKX1Bm0g957IrA
dRAU8XdDmg/+0w43pkerYQ37QCyArU4qyPp+gPy2tJAupg1rfAEHN+xyl9VA7TV2CPt8k8A6DKPk
ku4rlKgoYb/F4cS4l4Yw7bKLRSJD8nr/d+VKMinglT1yvK+K7qERUbMZGJDKjsws3TxpxBtoZ75Q
laOUzEqxOhFEPS90QoN4wKd2tda/f9yNqsKDahDO/7DFCtYBeWtT8ZfpTh7/OSzkUwdz2K2KY/62
phbFNLUSS6eUW41V3E1WvvOruo6LXyaWqGFIV7hamdwvRFmmy6jO7//3oYAjXd2HTS/J+kjNhN50
G20j9q5IJeeIDXH5jisWON+itjz0Sp6C21U/DEIb5BqS+vQIIUqaKw7rVgjWBqU2jQyjUIbFsY5p
nQeZpNvkeB6ECM1L7NVHzRcU9DFPvyZ9WieZnJC67aymha8DBxAQyl2l0IbQM7Ir0o8h1p/CUgT8
GuOj/ls0zUDxm7gwzM5tvOPpiFJFDatnKWHvEtvjEfh+NfTpKkSOGYb101y/6Nqd29IEtdipL7lC
y2u8atTwTa9K1WnIxR5kTvrlr12UNlK0bwIAAa8rwe1joR2vRWYrHV6NUHZFcyvX7lg5B9TTG2if
cjfE5NrWzyB6jMi5VTKoiMx1wFhhS9wiQwCtXNfy5UUR2wAkWV5QErZ5Df1IjcWg21uheCg8/DAp
il19i2V2ENFX2EfK9I8jBnTyEKih6iBH9YtS6nBtf+9lRnBhLE1Xk0PMmAzCc0U4k5qVX4dQWjAI
e1y9i9I99Kji+1q+TVW3DewMnwlrIK85Z7b98FYGnWQiwDLM7DuojNXHbi+/qnn9fOOD3Oj4ES6/
SsckhqIWuiLtvYbELUeCEE27//DmPhMZdZWcCTTXvhX+5AkZg95mJ8n4g07GgvUXz8rbqJA8Fou4
c5vvDCGnhE9mNSeaP0YDxXVPC0xwo7nTNcVdEP4OVCtx6qspBZMaIOfSiJFS70s7v6W1xssDFqja
PgbosSV8Nn0K6FsGs6mkgDAka7kNUK3wY0NVnGClpamT1buXybUPruAibakGG0ZFLUWziEHNSuXn
cXh1deFHmVF01AfePNtPBY7baXQDExAlmiCkBbTcOMZlcaqWUBRKt+ONQL/UKv/AA+o8/x0G1MxH
aNDkzx8+HPPk8T2Cf0hbGqkNxLnQwfNMb5AuYdGi1WSm3D3Mpk8pLBFqL4alT6Pw8k6U1KFSz8Wp
vN6m+X2D73A9V97V6XJN2zqeLcvPXzZMZF5Rlg1vVzv4aPQVkL6CO38/1v+4I92tnWHD7IlvKK46
IxJhUwzfAdZHcnuNyQVp2UjBnXXi6biJamne9wSYomO42bXTprj+skC81Gjxfl8eliZMql0XfqFw
U54q0oynTJvIr73UES+aYMdTM4AEeBcJ296HWxdfFir4dDAYwTaNBpDN2uYVy6I/R5s33cofyK5E
B+3OfMhQc9alOHCHu/LYTYO1KzNgzOTTDQRkV8YulzIPDbdzUflwHvN0Cn7nbUrMWqE1c+wcXLnM
Dw+GRuQA43lJR7fZCwp9JWG2vT4oPr0Wl+/OzpmouWxOQfpq6bKJSOm7nxS5eImMmGfPbjGnOo7d
YpeE95Kv1ROV+Tybx1NciFMcYYTUu8SawVMrFXfL+NWgKDia05xpPY13UG5GJtTLImmnAClpiN+s
Lr/ylBUWof+7rDcBwHlDzTZ52QcrOFRe8O2mnB3lz40SXXpvdvaiKfVr9JKWYddPD1sarUfA1cIq
1t8twGJ9tla7KLoKlCe/QVJpdZGVoB1tUr474sAn+rmK0OWt4LzYrq6FOCo0bAhdEpUY4KWpQETI
u6g9uSCw1jucifj5Q2vb8wzBgY5m6JvBvqjnf7kGIkDUtY25UsYZQbTpq1lnbuVA6PYsAPCvXPgs
uE7jNSVhJWlNtxXCMsePxqMQCjjo/JIHsrGtiLL+5YYxajjLrHs2dj5RV1eiye+EYc9nsLWts4Gm
8LSy4Hd0wpDHbc4kGr9G2b28mkGORQv9LTi7s9Xawz5a4vbnzjvhpKW5cn6gGBt86sEji/6lpfLJ
exBg7ib/h8x97RzGnv+T/uSlNywCuaXwkYvIIRaQ7k3GEWtokQMUOgdYTUAez1Nw1zHZsyCHFJxS
kArU3B3BKuPJ9XkGGHRccs+M7t7fBaofhtV/erwezv+wngmv62rfoVnddGKJKCZ0mSjVCldlQJR/
BlFndS2nCIxstCfoeMGXxkYo3pDSm21nIU2HoU8BfWnzG+nYRCKWxnmBrQ0BqjPXXVgesdaEWSs9
I4uzEL94k3NT2evf1mP195EF+8eBRX6x2RvXOmzXrav2h9FqP4+Vgo6trId+ZGufVwV6jqRAPqXV
//XE7+1IoFSGFxEUhax39B2gBsNWTGKFoKsplVDUBvTY5x0d+ih0+QEXu6Z9rlYeM4KbdK43Ajra
dwAunh8uudwZYSZaVNUpGSRJZgqTHIx/fnQAANdIRf5x5O9lUVmM4HVfsT0OL/NNjU2Suypl/qzw
w4GOtdBqr+BFEif3fr1mGosmavfWHdU6unC3ucqNOzvxQwR05+Hr25ys+/xIVH4gLsr3xUInmu6d
C5ZBqtiBSLCCsPsri1CccdZUXj9Dbq4M3zsEJdmqsIk1O9TMDFLg1wDiOCG59DjqeOxDkRMA8Qhy
pzZQ8YVkbudtohBdYq51r5qqmEFovZS032bc8NxjceBSqE4iG1gt6lI2P81xxGbJPYaTweaOUyDD
vlrYd3gdk5GZJ1AXJCNxU9dgqp+A3YS2JfDZTxg880uiCXoaD3Sdjwa2ZbTxSwzBht9R+ukl6o/3
hpfTDpJH9beadlyuHJtoJzgF1CTzw7Ui9wQgtgcbVRaLOQxRiPXnGfVFIADRj9GbdnLWKsSYX0hJ
FFjKUYfzrVw/sbESbhXHgS+tOrI5If2aHs1npBp4Q14cvQd8xGubTb9klU4gCgXH4IjJjyyr61zZ
26Y2d1hd/Cn8CEHMCnz0QkYrJwD97ZnBRsuEofjx60eOxVk8q77BH7I9TqKr9HE5OQoksYIq+SWO
YLv8nT7GTN3NwCHN7HoBw3BYePMX33eFibUA4qSVIKf6EcXaTQh2vqfHJYFU+uAGfewMS5vMk55W
caCTKUEyWqYQ0ndWilwVvjMexPpmJScaGK8+xzW9+67ixj1wYMnJjZJJoXEvcoSKWzaA0f414TVa
v1qMxqYe3syRD+cduwC8NUQpW02dDpcOCKeUNlEVToXXEKGsliIlvwi6LXCohm3G2RW/Lm2o8xV4
AwXvX/rX2INku95FoksgZ7vzGb4DqDV/x7xBbaP0fWjfFyJVRwUKRjd9FBv95pa+E54EfpJcY8Lj
nb1LXQBUZshkETHT9EHVCN2rdOnKa1D5xvrUc3Qtx+day7QBZFdZzwueT3HzDvc1fyLif3OpVS9l
/h0GOpKRUZftxGB6ZAZaPwij6K9SbwyA47OcyyAfBlS/HgkHhMxJ9sdLv0tKg5XbrBc+c54Jd7IV
mr2vA2tXqxIWchaE2d57QY5Dg1MJoGA2oIYF9V9VBb0RhQmjplMUrzK3tROUrDaimzozBi8jRRHh
/UeNKjAaDsuYCJcQr0pJ6BaWfLLOoYeNXyCUi/VlRWBSB05Ha+qbxfYTlUv7hyokRrwOhcIZ3jZ/
ITpq+USxbNjgfbP53fG3XTAPxdxgxd0R+QJ2Z0m0dbnrZxIYrqkGgmTNBYq2v2/kyaARhFRCJX6q
JTbV+KlN8HJBiC/TOOIES6iFUm83qsuIK2yQjldh+nLGLjUjVmowQunmi5uJi/TDt1xJp8hDHV0f
Hl408nLoPOE6xcS7bm7gspwPNcpeFZMLfC77p288BQJebZtBgkG+48i8XHdO0Wz5Ar5PuYtOM77b
Rw5cRaMzToRvBX4S5jvbUpBfWayDaD6n+mRMAFurpGnynVi/Ovxyf7h2n6PRfbhysb1YCmwq5bIo
ia4S06L+JpZ2QjMjv3jE2W4v0goA50efOCRTS0HQWd3Xw7XdVE02cY02BeHN++SATP+kgW3iG56r
7mB5/FRgwzRWQjZ+8X/f1rKEg1XZiV6eGrO7QQQQ58GBoh3qZfWvqUuLq6QCB5+ZefkIupAvZyLL
PoDOuqYa0ssPJgfSD8OMNk5OyczVd9L7XRP9tAj6TgoTutLS+Px2TdiDgr3bUQRy5aVsS6IRux7x
DCo0F2AKe2zbciYTMxBnp30NGOzKsxQEQu5FSQM433GYgeB5FPrvs2VguTOYGVJMz8vL/QEVlX99
xCa/CrPQ3oMOMqCKJ0RUpPSVq3oLGSdGDNOQSFFs1rvHjL7YJS/d8YOOVAfqSURn0yCxEV3BiXwU
0JK09YFrdZCzQoNPf8GkrYDbcODVtwHkm3CunIPVc3AepfJs0rxw1u6j+QotXX70/z2ix9eVwYiE
lo6U7Lkw42Kn+Uq1QWcw+3NAXjXA5cPq25/V014f3G/UNFpxjrPVzZc1Ki01hlqphoT6EZuLdB53
wMI/4tsqyc2lizW1lE2VU2LmGNkFTDXfYGhjTIjOYKbTmAC6GOtqKTTOrh5mWP68qJHvyRsWO/Yd
OKLmz/xegrhRMMmUXTI6slX/JdjC8ZMgLNPjcomaHz1STLFwoaiCIVU3oDC9miWdhgn/JTKDQdOl
RSPEko8TPIPHLeXERh+ulqM7bttZCnH9MqiLASflLaH22ylbiNsa1BmWCe9AV3ao8A4Qk3dParZf
qFRvZSj07GQx8u0IR64l0gRxAYNHy1o13h9/gioinpwKykAb9aDhzZTz4F2Yg3mSaeBOyyPI2SMc
1ohmDG4RUaVQppoCFRnR1a0vmnW+WWVoMsB9DkjHMXFqvjRESj/Szsd7Lov3lJ9xYdASNLo+plqJ
w/KLpx+D1f8U4n8WM7I89zcRS7OAeyvRQafllqjb1I14RWhau/GQAHNAbKXbiDm0SiOpDVubWLsb
L26v09jgPCQPlQjhKHwK27hwLJj0a5/WwOIDurbrYSleAQ8I3tJ73x8J5yo++6NAanfSV1oPz4Wn
R76JWCXQsOWVhg9G1dEHHQa45zlIyllpNa6A+A84iSyA6cHUgekkw7HX6PUcArmfNYBjx7dnAfDQ
exHBsVQPcP41k7ArOYrY4hmayBKVW4D6yK4bw8xCFl2o3Zja2OSlJEExyIN7CP7EG4tc0pOoOLFE
jM2zhXlZpBB/jW0lubfvodneBeCvn9aSxilmsKZlsAJOF8Pb/eNXGgsjPgYsR+EK8shBdqop6M22
Rs1POge4elXtVQpEqWbx7LXZYOTMbx9eDVz6TToRSGkE+APQvhZJno8XUs0DSg5i2CdBlqRL38d/
sYSlBZk6sfqG3ftipgTn7s1oAhjJCOsG3vS3sM+OqZXa4S/M+PZkvs+H+q2+qQoVc4+DSzaGGGpV
DOERQc8v/gh0MiJP/1oAjxdlQlU2hJzPNsaxTlYNjCOiwmM7GLPuMg3KOIomntm3LBzBJQecMsZ/
/W7TllJwtEz3JR2h5WutKZJFJCeZc7A6GVAPkzDIPVpNNPYV8Ka2VkqPSifBOT6OokU6qXgjQb7M
j4B4kMRMEswgSQ1FmdX+I31uZcLMcAJjVPVUE7Q8erzuEYZPa+30rU+GWsvz5s11ZNnmzoCjJx4s
Tw4LEpPXwWsxrBC9stavFoIOiuPsVFFLFCoKg2YHqA//5E97o5adSO3QtRSrx9awBubA/az6hyP7
aYnu9RB8OX9JDHMkOGtPGchwAjgtpqeM9r6X1BNbWjVikvll7tr1mDwQY4JAJTFunmO2aaWkaDwB
/kB33OFtrrcjz+7VDcim4UXkGHHbL9JQe64ovdQi7saM2uGxyqCPX/S38VxGlXif4O+qhVdM8oJE
r3bNF2gnE9MMePuMq0opLX1OW++fyaBcQNMgq+w6lD6NZCvD0oix6mSMAXfzANr4LrN0prw96Tdb
WfbHyFH6+KFmqQGhzeMFhQeAw6LcSe7QPjqgU+LtpwUzqMqAJSnPI2NAyTUAUQhYo5OU7Xxal9D3
fPvA42G0+O4p7thTrJibSqPiZad919+5JgtPllPeAK+60dcPZUgkO6fVDDmBxFYyO3uwCx0YB8nM
Xo+W1DuvECLZDtAB1BskST2TYKCh05xl2buQGMyxKvVyyBVui/I9O52Sp2FwQaeVACsIeyJauyn3
GmV/m8pAL5UY8Pz7cr0UxJ7K8h6AeCzCr5QWlXrRYyrCtTMBea228LHE1MfVZoGMN3MxR33Y9lYI
1DVnjOmzOJBt/Ih33ihQiXDw7ineZK7BU7OR21+YrwVGlVZD53fwMOOuFJjGSgzfwvuyogftB9Ig
RI0Lu5iDIzVj9enWHTRVajskAEdGRFMMFxi8ZweMGnYQD/zh5Feomb6MZjlNhpI+lzkHDbLKmjQp
DuopYGHlQ36e54nV1OWkuZSJLhbEknc2uf5T54uA77y00dmjMiuSF5rmxGIugHdEJqGISovYLuoN
SrbLDMy7UqAjrkvHUDZHNble+c9H/9qaHY86wq+g1PJgA7QnINV33Y+F+uADjKHkNCuslE1+n2dR
Jc43Ezoca8wgvetyHv+0U0lN43SNfVCqdbkpAwzs+ToVz9fACTs7wIAJdxMfKz+SInX6u5QDDswh
Gcsz7YAuTekZCIQ3GXqC4j+WtvmdKU8vQulTLJOn4gvFib1sFQhN5RDF3fevuniJ4sM8L7WrnbV4
tSTf311JWb5LRXW5B9lXkTWtvKVnlcIjFaWOuLhYl6i0v0e4GrAPH8UE9PMkBkZVQGjG9C1DOyDs
TxU4lqrttQkkFBSKtO039TsSyvLwjHqvBLafjp8NvT5l2KONi+Yfal6cZWmlk12tLA5dgYtc1qEw
G7Hs9IyXKFBBszvLiSwASOF1ybN9+7Ku4ETZxxTObY3+3/88golNYPZTREHmPBNwAE60sxEk2Sx4
+9Ufse3w3okMDlmjwJoAj38ayHWUFpw76yxhQD1lxLn1OHEq8gD/FVrphgzzDjJCDIIHsy8rdsMU
GVZUfryoKo/LvAO8JpiYSS2W3F6tEWJ6wZTgfm2mBDTXpKG6PiiF2jbV75mOAyhaWNBh7UEStPNL
RSOJQkOOK3D7oaBgsjyhcAVz0P2GyZipO3O+jrfUqFyMqz0uhW5hyiPR6R/j+EM0ZMoYorILj/zS
UchA9SlIlrS3Ng7YvBxiYP7KnAMtPmDziKdky3da8iEK+eeQ3RoFwn5T0ZfqAscVjGFvL5QwaNi2
15n6WrwMpEXr/2nvfFqCj1EOZ9nUAsNp3NAHctIR62/vMsKd/6QXkDqnJ1vUueifq5VADYtEbcQo
yqyXnjdAQvRJ0ZO1NFIjD1aO5W21nbY6It1rv2uctWgkvcseuB7IcKRArBE1H7Js6jbmUHyOMPGl
rOu0XL543CgMbIxh4iy4y7jd5rpLjE7rH12cSGRThQ7Vi4Z7s/JaFw3hyFye4M5NJyq+YCjSgg1a
74Gcuxe9uruBmzSqlh7e3y42lvvy85RISslPUW3eh02Ho/eXiswL8NQClMS03obt1jezW31TPUNc
+ldMhPe/o1fOu076IXYo8Pxd4KSbPYS3+q3qrdDB+0bpwCxwOynHDtr8pYvENMzo1o1bfzZTiyQf
y2PSlysG4egEubZ2Eqb4QzfNZgJEeEXYpRIkepCWdDguEdGYfyjNo9WMlFNE65sFO/+JTzlSTqf6
oPoybw+T5A6HMPiyqs2wWEWqDTuNvBG9KPwRTVALL+oyox7Igx8CAXfx1SAnfraKXXhZqa2pt46K
eU87pAnfoTs56Jh4cv4ye3qNVUFk1M7OU1rvIxamXOCFb4rYggbEnCbdjcXYYulQkP3m9wDXg4hQ
N857JbZbLtlIr7STD1fnajptMZBh6w2EBhWpPt+18dSDphUBduO46CRLfggE14eXk65HUTSJxZDJ
TOTRYG03Isguw3rQEt74gITnXbsGMjTDeBVqVVhwlEK1BW7SvzFQFNA23104ZSNJO0CZSxF4VKK4
JkG3w0g2Mta/ej8fX+7KZ8NB1j6Fbwj7fW45q6HIbuBW8ueBgaLSF//gJuz/qqm+3kEayjul6+1a
wdH4Qu5tsI4CLpRZc/fCD4VDTPoZZCR6ISpnrg4EZaDgh8woh9C057AezuTa3HarBvV63UBzbfiS
IAMSKPhv8Qd9AjHq3v9/+IzF03yssg4kBCSd00h2FqQGTHqdAGMe/A+sg7GWOthtBck/X6UPhm4f
VaFH4ItVAvZxhnFz9BIdlpVUX5gq62n75hwoBjdQrIzygg0HyZqz8mDg5eBH6lxGKdyA5iYpE+2r
YM1yf6OjwIAYrtOGjs7mEA75rDWVORmt+ZMJoqL8SfTrqo5/zjRokIaGFmclw7XywBIWNss4APyT
vX1fiQywlD4Mm7akPQE8COF1mBHqdxF9+7L+tMBjNgG6+HZPieGzxADVLzpcEwUrDWyRgaUN0rCV
iRNnrWt90NV4oI2pCxlOIJExoFBDToCzKvv5+PmFr94t/FKDtDFNeaQJzFOQsd/dip0b3+eMQLd8
ioO9+vBKDI2zh94n36btNVJJvFOeHjBCANCmku6jAhNHNt4Ci/P0rSLhXy9S5YQEATUIn4VyPNYQ
rS80bpgiVppSBI/f51w5Q0foqZmkVzJ3B78Bm1/0N3c06h2G6viV7Wf6ImV7iIC+lGZwNlR6rTBD
LBk9BvDSqeOIqL7QSgbXb7zaWFb8cVX3fuAMJ3sAV1EcfqhyZdsaJDJGGIPlgsOHCX2NiPHHauyX
ncQ4S6purXAubVq6cEy02hzLZD9wu6gOaF6hn3/Xh0faFFHt2Lg7iluy0JLCT+WABLPFYC0dC/q/
EAhdLbr0oByDJC3MLYlJLVKmDgJ7kfeSIbXamfek435VZQk8m7wOldeMOjmDo1jY6mfttviEWcrs
Jl/YvtgvAv8P+2zpxMG1/bvoltszTyu3uWwUfkmhSSDeMGWr8D5S92J5tChgm5uNNxd2oC3r8BDb
R3R9XrVxTSFIIanAUM0GKGIc4X/97i4jR+VNIqbCnHhvTi4Ua6/vNngLZWSFWKsqqrppdtf2wet/
TyNyQdTAKCvaLXC7WVVHMow2VpAl59W1jUw2Tjbgu5FO9TdfrqJN1MhwXVqByyo4aoS3d9iESmsZ
ZpUkKbCQQb/LREA+Vy+zjnt0iky5xaxdCoeFJH7XYTBGnI3CxlydNeYjmXv2+M9N8pDEbuFOGNjO
b0ooGhGyZujYoT55yqx1Qmn6+Tl2byB9lf5NcNSIA9xxHKjkRmBjaLvBo7ocCZGp2dptgSEgibpQ
jfN3fPr50feSqDK6AZBitvgJBkPxX1UjrO9dcjgmqYLlHrUW+9ycPDgyTKNvtTFqtN+dU53pRz9f
zU+Mu62zDZgbDV9vk3IcCkCWiF9tCxpF40xKo7w5cbN8bG2Nf8xN60DDGUsInvsD2USDli4ODK8G
qKUqHtv9Q+j3xfr59KDh6mC1l9j0Xlpevi3CgXc+gi0INIJwqQn51RSERvkluAt1aEsnLDugotLy
x2VeTSQipzMpzpxI/v6DrJdCHCZCB0AdtMZ/IopshhV2Ppqmp/6QMvn6p/Ur65yA++uz9VDQGva/
YLmLUf7ia1NoLbIbYXZ0vWku1IpgXI7ly9Tly9nuOjK5chqSll64Wiv66eDI2lh0j5uMKTUcvSvv
z+reIX/uiPMLQXlkMt5xqvD37Rtkm67NNWtDHvcG8wxMr1IsztoEuiWgCoIGZnojcqWZjcVtuch1
lSy7US0hdRJxGjijCkvzuyOj22QaU5JHbdK46XtGPt9OqWQIwV15X2iIVOOBIy/s520DPjwkATOV
stLjdRvJ34G7o5hPjb8DH8orAEobRTiUwzW6/UrhwUUjIFDRvQLaY4OcHhDwGKYgwmrvocAIdN7n
K0dyuk5mJ3mMwrZ3LHvcbPHHUK2QeRR0dedNsSa/+Wt+MXNR2uOwKOUohaQ4xlIZqRGYwr8gYB6M
AVqVyEGbpinyeWLw7/HJc0Pm6NY0doLltzOdgj9KVwoMFUU+TuPbg9RXdLE5MFPzfBRV7/MXLI2K
m6uNJgUYIMNUjHsdCz87QKhCxqWQCT0gEe0kz617bh2CT3hAi6nAAQz6iAlLg314wvVc7DojVfht
BEt+Mpyl5m/x1mI6R6R5T4FtDLI8wF1xjBXK5D5YoYJUYk/rCbe6QtFi1R+fovVP5SLnwjAovc7C
07x16ZRfkP1yziVlUS1AoaD0yNEXqsEJRr4KujWZe0Luc+02Ln5lNbJS1K3uu00GT00iBmxT5X2i
ZCsw8c5IC7KOLq9kBJEck0uPVA0CqCbBMlLTw8ksI4LR5+G7ikmhJWI4vd34yxonFkeuUNUGJqAm
iHwIr7jMVHWrAkC87sM+xVFiDFTYAWSsJSf7GP+Ns73VrqvkR/V1AwCJOJurHqS1L358oxWSRHit
90IXBhDcXAMfFfSXJLa6YLfz6YQEPRQlZ+ZQsqBmwjDizciCykkeUljdGj/An31oIktEqCafmfAp
LgQjJthDP6WPuAv1SuIyh2eV+CxvtjTWQUmSOWI8Civ1wCDS8aDJv9P/IShnGjb8e1LYQll2zxkL
qqrwqKnimQO57HlUbl/UVtGC8jXxCF40xufRqU4GxiWjGgDmBp46Btak+NH9DrH4XWq+hOOzuPo9
DHWyVmo1NGnsPe/xJS362kgdVzjOfxCF6CaYLVfjGMqFbnCFSYjEdM+CHudB/VkO2w5gyB77Vj7J
QmMJROusyyuqCX1XWKLpr+NaBwcOZRCiQPWQwc5jPU89Tk5Y1nwzUFhZRlI5k88bYOpo2BcazoxA
V9vyu7HGTyl9g+VeCp2H78iUTheACVgY+8qRZmJuGgQDuHe82e9ypLMTKL/fW5DfQaoqUWl029d8
r8vzNP0BGEqMo2huMEb/pN65d0bpzbHC9MzR7VJKYanyw2S0qPmPc0kp3BXVKn1WkPi+tJz1uBNL
EuSbfoF8mbk2nNQPxXGEzBFWRTG/XHWRpuGlQqlHxFFRr7FXSBf6uLNFMVZJ0TYJRfV5XeASVEt7
w84IYeyQx5BHDRHFnnPmRSukjVGvD9zAYPdGsX3uirH/G4Rh85dH+BVuQ/1H7ZpEBmaMy+LZjAfd
d5rYo9yBn3NP0IG81unTMbRBoZZrjnJcChRPkgTHNAt+UkRRLTgLoLf/hjLx2Nulbqo+lOcSwbU1
3VvM88U5H2lkyTV4jDlblHhjJw28UwO4cT2OXTzHrxX6CrDVwICRQtGVsYeEX8vVRtvRbhWokYX4
rgNFRpNaxthR24FSKQn2DB6LMJQ5uJbFHNci3Ck6ll0KgmPGe+81XztAz5/lDlfpTfLjT/d2dxEh
C89P8ZF/FtV7R5zhh09DYXXOopOAk4t7aD3K3urTVt5w8PpmZng1MI71/KELyhgZFVukLVbz0Ykn
xDFm3K7PpkvY1iBEHyyamjrkA7rCYtCAFzkOBUjrdRaZQUGEoKUVU0kmc0Y6ohWs03uecZrShC8W
I8Q8S73c1dqlOCggm4EAB/S07Z9Oo2xG5AT3LOO6dhTjGvQO2VY8skBDEu7AYnfbm0VIhIJWq2UW
IdmFky/gY73k1/ZfdARnGOtgrazpBASGrsMUyi5HQsabafMG4+he8zd6Z57CMm12XxZ3z77BA66+
aF84QkhGBqdOvGHQXYxIR5b2C5oheXVlMTmwvVwxCGaoyKI7RQlfH1fRVLTStin2XN+ApXl8mFec
B1kBivZrq1m6MxVRKWo+5aznq6FqJlZSj8litqao//XkKP48ruRN0YkX4fCGnbeYo23wgu20OQ/E
BbBLxZSSBlqEqXP0V3LHQjaoFVinsHZ09wU2d/n9b64xWClsPCO8B4nKU2qavQDNug0bMk/J2Eom
u2Db9aE4jJDGBuGOMmSileFIVbHiobESpqFDW2TeeY8/LMyjWaPjmjrdVL1JpSpawyWJID6KTF+Z
yYiASmUudGSBKI6aMvq7OoVUiEgodv3swkI3lyFs89X1tVBbhdoJbe8JquvRTWYhf3yJhbrmZq/U
sqKS/H3RC/mSbdH6XOstvORr1fXLAFrqJ2Md5fmBwlqp971whHTgXFiqAcAspLoLPLFZ0RKfosmY
Iqvp/0MD12U6Nz/f1XxCUKm8qOp5JgF4C0VKCXxuWbCxS/WY/dVzoW1V4h86mEChA5q+tCAEhJtW
CGaoFhPeciS0zz0LHPrpR36FVjDbngAN0l4QO+Qaklhg0P+kHboaUZlJLfxJpUSoWl7Kopozi+kq
5f4yrsJDMGeWqYl+uMBr/wqV4FX6Tc7ElJBrV/ynyYN9qqq1KxBTk6MRx8B2ZCDoHlSA5t0Tgi/X
XJtU4zZwKmBSQKbstbgv591nz26cUp+Y9yb+Vy2aCf8PRKpfb8rD2r8m9ar53YcOH438kErvu2Ja
HVuI6jC7PgUhpxduuE+5Ss1iws3qnzYoE2llus8O9dwq1BVl61ZEtiK40Jkq0fxRT/7Rh0YZhnQa
9TuOrkPaFRFBtdwJm+dh79/Yu7G1V9VJqUIrrwRw71tq53Xjb4ktvT6+n/912eRhFTL80kUDWgjY
mHy/Se2WwDN2xe0hb4zGBf1P3jDmUCwhuFCEzfJGvbsUEPzdf53PxtJwwOwd9c5z72+B17KlqwVa
IgSq55KMLj2Dn8HyQu+qqs/VqwJJDsJi2PdiaJChxc2tFF+gapF71ZvnDMnSw8qBmU9KqJK47jK+
CxA8zzk010Wm6trui3T4TATZlPmRmWgrMn6ZkBoQEHy3xfjhi3RFkRW2PIPfHRlq1nBZT20ZXLHd
SdOz87y1mn+rTWJcyyUnRBqZ6n20uwN6bzL37yp1AzMM7zJ7xKf16nxUlsKj4z/7gut9AxrA8vUg
wEIsFGNHTTOWXx6q/Z3ZBssnooB660jITcVBFSlzmhj3XsYu9pne+59sHvMA9wu+yj5E2AJwQP7Z
cxfj7RGIX7WQQc8Qp3pu2Eiuep6Hsmub0pN0qK/AdZMriB7Ig2RqjM2VovCLnhMha33R5t05BX4e
CNJ1B5qsIGDL54bjT/PDrrk0jwaAZAaRE6bZPnmeb9FFSrZT9bBsV/rtcg7Mjy1woMkVwWNvxtCL
PAOE/ELlNCf5S3mJGJEq2mtZbxlEIsweGp+t68AUoE1eGW4UFAMHt8Chj/Xka3x/RLlyc+SewpcX
ntg0Tn1K7CfVmTkfcG748fbnhcwNsQGDUntD127jid28X4n3VHw6gkgogCIXP+rD+p9RitIsCNrn
Tlc+ysL5nrXUXSD4mQdqTLVcKfXvO9Ypjw45rNPYMkmaOIc52i1zaB9giQI/koQ3Jn5ORIJ/x6rS
qEyy9vWC3pF+F4zQiHW+TvF9U9s4VZzWIv63yx3YRq/g35LFpsKKOZZjPmLukqPKwFSST2bIOqWv
NUzmWLeu2sOl+ZawR75XNTAzlEkVr6DrBom26Y/omxwJI+pHFxTbo0z+XER99yOxd4NoKs6WikAm
2qp5+ZY1avjmccpay5wDDTRgwELKVn8mQUs2yQaVwKY9iD9Ug6k9psPRqyOX+SC1dzntbfzUXn9c
R+cSHmHU3bhQ6AXH9zDWiqjdRm3uaH/nDL6T/KOuVZwcAO8rFXqXy/GxSrN3CWzKTk8dZ5XnekEm
vq2WvIoPSKX5IsQUBu2uLso0nb+6B9xEJMeBTFhuET/3ga9nxQsqmE6RdK9HCRK9m6ls2hxgqnI0
QePMS30UM3TVRU6oe6WMp+JYWE+IyQFLtmRRjGPj/2LmW7O2PO88QcKnfERvt7XP3wIlUMVm8tFb
x67pfJN8ybUSHB46lauij31C8WJRPosEC6HNaM1OT+eP/+DMAwICvWpI0RQ22K4erSqlmXOKE6qF
ZRwkDX7m511EA/QNGXgA38WfMdzxYezPoRDu+PBdap/md0wSRGhxw43EPVWM8AiEh02HOsJhx+9I
BISOCJaLUGxr78odOM47qmspriUdPmY6ag4SV3orz5/1AvISdUdCEHhgHFgE+6oUTGcAFDcsfzBO
OvAdh84+aPnMKqEtPtpZ53Wu8FsBhQT+3Z384u/aWeZSO8JIvRVjxJkMv7z8RVJgb5aSsUtGveA0
ySaSaC+G2P6sCzdivTATvYC8rcWB+g/wOyR2Ze+qsbWajtuix+vuQnv3qr7cXGynsImJgxXolKRb
PwyLRdm5ND6wTBRQCqxel0DexPRGiEu5DVplhIGpiZx8QTdlnnRe2XINBD+ygjxwU+vkWfxwKpL+
qIoMwvRJ5gG8QtCMojminGMJKJfo9D6rrclO9gahfE7ALnp5BMxGK3IrQSJv3Z1v7WA3EeYeiywq
+oxeycK/W3MMnAxP+3hgSptT9m+55U9ot4O54gNkGNbAni2qY45loJ404rQCKCnZRocEEoy00xtu
bg/kjV2BHZt4sVIpLeIwZuOcSm+zVJpLGqeXEoAmi0y20xAHj7cUFxDVCaGpKyB51q3baGfbsCS+
XENFQ/CGxwLwnLmrWESqLHr6nKOhdd0B4gr/LRXg3Ebt8Z3ZOWDg5xK30ENRskXHJa4ZYY/K+30K
bPI7x5I/TX3VxmtVsfvu7o3soCaESOEUIHOaLtRlsi7Yd/+Q7exs2RMQwPbbpBT5lu0dv5K7kGfm
C0hg5U3T/zijNMErbH/fUzx5MEqNVgof+m+lA283clwfwfirP0EAgDuPW3a/yuK1du1/V3k3OAEr
cZGWQ2vbzllW7D+uVOPfaX2iBwfICCoBQcsQKik1pksXuw1Cgco0T7qg7l0Wbc0PzRLZ9dw7cG2+
fN+IjvkAOPb4bbnb0Kgbu7CFGLPqeVf92LWQ0iqhC7xolaU9Xj/5wMPyFvpD8Ssc1rlYxyQZXR01
0S6XnjWOcOA/Ij/quXlieF0MEr0CQ51JyD2U893/004rlPRpsPJOmR6XFV1R6St8UH2lSvtL6UQa
ZytpkQBhEeV3N2JNCsDjuZVRIXtW8cPzB1IK4MQpyrJ6BbRwnac4ij0l2a57U4nmN4Qc4pnZPGFK
9EcwycuzCOYQFQjbI3xMoxT2fx+JqnQdAt2nVp4WWJNJiCuuln4QHGgWnrfzJf7aIG6WOZp7T6jP
ZKepR6Z731jPYlx34d9EKiyhhao+pCiDwLEeTzOBrVEia3pYtzTP1mCuN6BX5JnYZo6Q/491NSUQ
wdYbJsciZlz6N261E7AVjbMxHRsQTC0s9g30HRJiWVF2mP1jokKjes4p61UyP60XOWlwK9MNU+L9
ROlMYUQltC//n7CvrlhJoEcpKHYGdWb2ZhC6e44dGDFthxmZ2/5ZzV9MkXUPXSabRwSg3x1OSKir
bWmy2XE04jX88m70EoReT+aBTu1GfFyafP3JzeacNNDjoBn7lh3qNLHoctNfQMH8meXH4OvNc6DY
9meBOk8BiobU53rjWNt+Jca9qGFoaLbEy7Yy+2SA4RbzzanjY4NnWDf5BauG5iFhuuQHfHGDOfOF
rg8wnO2rPviySguFSpNeKfF0ZUKgMigc8KWn5I53icg5JS1XwrF1E1n+gfdF6ubNSwRtqwamlIxe
J6t3vXUY30F8pEqorv+iiUdSs/mh45JDhpHY1UE8UvuggDDyNOiaKe6rj9BdUhWX7u1ZhjNnfBSi
5rhYd4XWP10UbcMAMrHrz2PFYiQ0428AJGDL3zsHzydEbc3MqJ+cHJPcUiCVxyd0cu0FvBFPw3pi
MWXO5Cw5fv/VcbTb5KdlMz7OHutLVZ/ZYo78N2/UvZhfypY8HKvcZhjVtlb9bhrH94E2qMCJ4kWh
B2gYL1+XuBHgJgOzjTmSoojVL3+IZHDRo01Nd7xnWkTImZkPo2iLpsEaDeNjdgoNwBqW11/Vlw52
C0TRyA/F6WQ0JTOnk/1Y4JlIBodHISOUPCKBRmuCmYaJpW+70tdkZXTTpJXdPO14l1JEl0e8rXj9
p4aSg/7bxwOXV9B0XJGObrEJxQQgBkdcl0kZZJw/nPd1xtwIuvPFzlMbWCmeW59OsTR3yG2fumhY
y5afXI0sFWsyc9U7lmpoAGAgdlmcBPDm0w5bRlHZklY2EFQa9NrXbD3Goxsnnt+5Y6JfIgpfmEfS
S+trOqL5uK8ZnE7KZ0weTqD+m6/wHAYnSIGIVceB/vBTcZ9k8LLk/kQ4Pbn/ld4yhTnGF4/yMCXZ
pU40W+MKd3shWP/31z2p2QawyykrUQWDLR7RufdoKmrQ7kj7aWxBk7E4jq8bGUgMRw6y9xWU2KNt
v12LQV9GoWMGdhQTDDK/zqfFmt9ffzWHJhZCpiHiE1kuVYFG6AIPg0nBwtSbx2eK5hm2PDgwlkmR
i9Jbppm2JP4Ga8nKp06d0IXDq0yvpO4rFOxM8lDXlJovUQi+MkUu2uelV9qJfSr8AQHxnYilRBWZ
NbkN5BYTtn2DxMTHJX9IJ/u2SZDnnb0MP/GMgfbhpYcxPpt9GLAY3+eXsExnBJh8VK5EjyoBbUsA
pXkUJz9L0zAmnCBknZ0ZfmTsQPDW3cMOsAn5PcpuhpgK96xvkvItBoSi+FGR/sWSU7yKPNQY86cq
LxGPLwqstXqLateuf820YWJcQUBOf4/HjETRzkyOaYUZcnSZLZQot4N7u9btO9QpNKuoYOtdbAV8
lCyzy/JVJMFrLkTcxTws1WTfPYE3l5HgcldJbeJ66Dg/V7PbSLeArJRrWEGGvbSLG51ZtbB4HyDt
3Wgcmhgb45tpzxdn3LuV1VdX5n+y2tibYIUfLoWzXoPlPCMc8t2W4HTzI8C0lDYDlBRgK8wxzhXl
+VnDrYyCDFDPVjQwRLzlFD5OCiJHmUW1yObape/JWJ5p7dPpLEjibyzpTSnEfeTYMT5uwvHySFJs
EN3czszbBA+RKGnQs/C5FAKP2rpCbaiYpzAeBuzrfbb/vUI/6ymP9969C8DpNxj25j5jPXUCN6sd
cbw5fftkWuCpvLwVmsNTg8s7Yc6TSUee3BuyLEQNbNK7/IggxszONRruk6y62PLE7N6p3mR28dUQ
SOTPIFo3R0lsGwSBHxK6BWEoLtnf3VwYM8QKr0ok+SgdUdPDbxUMeJzsScWhyH+fx5uMNrULRTMI
0a3OSuK74ljc1Qn3skifJn06DgwfZvK81V5SH4Or8NapcKOwjATPF1zN+6dR92aD5TFliopNhnhT
NiRMGAVx2l0L49V1vp8pc9VC3kfBq5ykHtblIVkP/Q9xRKfKT+mJjuHVyyMri/7Ww9pj+0cmAWA2
dgjhckEmXReCCDZx83XqjcNrAXKgw68qMCXvGpV11dSP/we7TBJGj0elrB+R4BVuRf4On5UX1lCu
x+IVHu7v/RKjJvVTQ7VsLcfxxnZcMOY+/7hlPrYvb6FB1ckOiTE5QlU75fHPCRKOWgQDlk5pWlwd
Ms5fIStrFzFQTXbcRm24YwNx2daQH39ooUoMh/t/PA/IdudZZkNYj/1YnxRiE2fWgjQg2Mw+D8q5
UVUcEST8WZ4aBS+wKTCV20Q9ny2SyYBjMU7f01fNquFlL2AIKL8SWk67NgKs0eDjiPeAsHv5x9Bf
cU92s9kK5MD0LV68CiN9DsXr2pJaVsCjRygPpP/gmX5fqmGF34n9LE5RqHTw7Ld4hWroFIU7hrWw
4WsI84U3lIVqlh5VTePdlkTXF8fdbzJxTaxA5hFPhAWW2v5g7S88haGGnS0KE46Wrg0ne4q7jC2r
5Uovnm0CSbI1nQ7wF4ldGBaVpeLEUOSmm0+9YNaqa9Y7/jEo/BqGQ+0LrFvjnPRsrZPV57GGl2NC
bmGOPUuPam3+oCDyzNfSF8KMsLOpCyu3KLtcL/Od11j2KMP74FIfhxqMx718+Xr1bo/jo/KISfYj
Ca5fJmkF03YkQY4ao7s3BNI456+yoelG5IiDBbL03lvAGotzxBlh0fvVW9kQ7sFzmytZCTtWw8TU
HBpR8IqX+FkeNuWy8pG+z8Q/mU+ga2KM2ku2sCg9ye7CECF6aiw683nMojbPs+dx2eHnccZCEoqj
ZtEHF6dXrW+hQ62kAaf+Tz8aubwPG0eroR2oE1S/1nPNXKfUuC/PXAIuEekrpfXM5FKF7RiUXQo+
C5ya59qArQhQk3K3y3MFWX4ZcB1/dZKW6yKonyWmWX/TIcrK8bMfU9pEvs7lbjCN2ZZdzDZGLyhM
g8DWZas/HhUSJv7JOOaq5fa25dWXhA8O91AjqDbA4Y44jgZUwGLK0lalBNmBsatT2X9a72CTbKk2
sCL6NEuItW63Ow6n9ZXmQAIlqVMSH7g0UZMakRpuYE9+lVbZ0zTW0KgH7hJFLixF54utkeH6h9Ak
wlxWXgrmX4d9fO4coFGOZNPSUqf4ATlygCuz2+ekNuTpHCXHumpwRuEN3umVZh/Hrip34Ex6DV50
cdcKz6xAIy4ovUXcowwNibyvtGkMj9q78IDNgBxTRYB/AIDk9FtXI1deTd2i6EE363sXtuQV6838
to6FaW4oz5jtG94/S+yLXP/CrCpzURV5TamoHgAkCclhoQY6TDqYPEHYKZ+bA/hjUzTCj5nLq6WF
zJhLnXmtYFMb7n5dHemNsHo/8A7unMqymhXUjcYIm/48isjMkF5ydtiPROWGuN1U5up7kCH1LKSf
qMJ5Uq3+RnZGb7GNaweaOvsbGcqMCFum+IrK4buufFvm1kKx9ykLgHwEAmV1JTa/QPiGMtd8fssi
z5Q0SbetxgerS5akdTp1Y6gbUXM0I0HK1nCuxXs65jcyeV1bRANN0u1sUf3rgsFXGuWqGp2ff1Zh
or0G943QZAgCj+J4sCa44Lf3+EQgbTAjt42yETO3xmyeRcctTygnw8Y/WcfA3R3tAyeCCIZhHcPp
bPEC/fJTvGt30qhWi+IFNr1AN33EqFRZkwthzCSlyQyVWd08iilHTFv8cQmieBhp13SOsF0Pz5hy
SRnc5Q+J9pOm7bibmVbJ1dsIo85J3TzuNLsl0VrYOOjtnlSdRJfHnvo26zxXl8pFYBF4jn0S3/la
gEYR8uKOfIW7DBerIQAZK46NxsoqQMXk9BPDw3d3geXJtogNUZSO6+pQXLf6OkHpfsAafMXDBMOX
r402fLhh3z8eibiKIP+y9HrBfXB6TMeFScQn4eNwhUIA0BjCbbzCwbZmizjwUTjUMxRGz7vrF+lF
uIoIN7jEv1sd03fY3jrscEb2wfQdwswgAUjTa+XPPl85piTWkB7UE4Xs+tEPvR3FF2IzOIATKUSd
u0q5MBVYEBFttEPzIDdaOsZegq5n5Tdlh2QPanT7bNvgQ4jprgwDwo5dIiy9DcldzYm8vFVibx4G
N51UAiy6jkHj3tIfxkeVtIRdqAY0J8p+dgQ68f/GQYOynP3FNZ+SjDsT+yErP3qog+O+b+At35Kr
bIu50nvT0J+JQKgIh2eRQE0QtgVeWo2LIs3lyCpFR75YpuAEdEmk+koyx3nVL/mxexChEtfD8r1A
ReMFkVAUtJO1bitgfqLJvCZXAOloEs2hHGqlLQyRh+TsVGznh1YF3K6x5emSo9n3aBU4Rg2IHGZH
2cPbQyMzgE5L3XBJK1sS/ao5AJGrcZ616pnFqiYZDMwWdFjiyOCa9uEIXLtSePxIC3CjzOaWff54
TpEnHKZxHbm+MUDxdoNvzhnAp6KXHPkx7Z2nWU7d5dpNTO6+jIxJslrbjody7PzFXvKGKrq+wjPG
WSK/TzdJY7wcfsFgqhsfXE2QHF3gu9JgAvuR0oOlVBkZQGVZ2esM9gnV4gAzgSuTJMwtq2g4Wgxb
+5wFN6hug74vSuWDWcP4EJr7xLXRPXUvMqUf2CShE7BsGwWog3pyXv6ef1dsgp5Pd/IDtUkTQK7p
pHMATbn//c6cWFwRU2uT/iPRVoakLIcAZeTW2jLaC/uEf7AfduXs2IMqFWKY4KirNcJEgyiW6FyY
+yuyavaZaioSDJcrG/VBB5cr7YgR2tnvdBZIyk2SiEk4IZQK0ElYskpoQb0dJbqzjnFwXh0XHwEs
3Nv0rp4nooUFT2m0L2YNbdArgnU1SaW52ZjEpizFXVtH+y1y4eFMQ7PbSb3fdgygOPTLK5XTty/P
/PLPQrwK7BD3Ap7liGUOlwn1cWTFaVSeEhZfBpQ1E5PkRzje315WZA+FArWX013sWXagm/397mmH
baBFDQ1xBLdmQ3XMq8/NXcaBtRYYm+gGeyQwa94KCgmi/K8rgFHO+n//jjj8M9MjQKkaxobVuVCH
45VWjg2+LY6piEwQJziPg/7mwWrDXdMgyXlNOUGfQocbWee6L33jHTWOHrYGN0DCLb3o0emxbSsx
1VPzHXmYU5QQXkpzTGLAmVtukHiRLatfs6cWP1doEcKY63nACWYihrmIrhBNNovKo7AOEdEhssgC
zB82BXD55r8o+AxCrrJdIbzxoOMh6e/S6n9To91w5FQkFJ6+akYJEMv0RcS9CYvZBHYQvVYEJnk3
zycgGQTdO1C/1myc1fpCpD5zrfSS6pDh0+270NcG9P1XxfYy30cVVzAXVp14tMArlzh8oYTwXjv1
Jb7G3iYHS28nEL40ULCpnXP4+w1AgyA9hH4jHEsHeY/zsfu9spKlMREks4Ahcn9Jfp9uVJflxrUy
Kgy0fagkwJw5NlZyLD58ehsAfnNErOyfU49scdNDC7uI3XXQavi+fdVlIYKZXHYGc8QR2HILUBEs
enbl0hcgMBd2dtpjUsjN/t489MMHILcsmJ6MWJPi/CgtO0F4FnY5uG/OwlG7+08NcXRKg8kVTzcF
OWwkJhNcXMMgkaLJ3TvwHF7X6ud6yjZ5YuobzGox9o5XkbLFt5qIt+HMMKQCwDs5HbP6erOdg4FJ
l23pIuOImHNLVYzctrqHJSEFGP7ZvltiBcCQxPWNryplweKO3Wmf/jTH4c6AOA712+AEw6PY3kUx
0ONvqreS/bEgxCJUaZkHlYTtr5X90iUVNzsyWJiGNj7rT0mZjwOhlsjGdb+4HFvg206AyLGE5c1n
2q5SpDDdQ5mX7uJfNbQ6V6h1g6DoEkSuRqhHS0kTFsQMHLqIMJLs71x21MGItq371gYGSGZhrqcU
hfz/2lyGOKqS7sOpsWhAtOYcubW+WjZfs9fhmcr2sZtLqFJHQcb6EuR3PBasVGZucWdLbaRgeXR+
JOK3OP85odFtpUu6KrZn87anoGOxb3zLnC9SHwHRxVJ0rK1kZ9qO8gW3/TY/M8Gt7H3Bnk+hPdjP
hlMdnOVSpGVdCqqQCdElstYUqdkPaoYE5o4+4Ac7cZ6E197GeaoVrlkDPIle2P9XSAJ4IuLInHPu
EETZd2BN8O4i4eCsnUy4CObVENSMOeqU0SyS+zh9ANcI1lZ+QmYVghxp++IM+zK4m81cNZS283F8
h0ci9E8XSNboDrf978hKQND4mnBqcB+jcDg+4YjJoZwM583Xtw+gnf3LI5sHszFBwUTEpvbZr/EW
1GTSCnAq6ZpUFWJcVRMbLh6DN9Af/QXJs+kL72fqSc9xdrIu8UvEanUwD61VcMxI7BSTPw6g4Ssc
z42ss0MfpCK4gsylGZUKl8qSVvjT5D9HF6cQ2gdo6Nyn0/uY6zvrV0ZEv0F9KmQPqdPTYjLXtAi5
MzJSB+5FqDW+DAaBAs4yhEC+w8sZBy7swrMCjXolS9wwJOLP5WYsy2qXjQTkQE4nAqxhGWLJxZsb
16xF3Gj+qSUMdDJ12hnYwBds1IlpgSK0Eud53ojBQ0P9D5NlMwdsmd1VKo7hyGZxzkDsDH9Qr6Rm
7ud2GFajBL+cdDcYSA72yVDoSZx2FQ5RQe+hZ3caqHwwyDXqZgnYP1eBx8ABeCfuFpwIx1rw2G7Q
j1TWUJRTJH2D+AiLZ02NNz+SWC1dy6Vj8qG9s6rJeSQKWo/ESbkh2M8jICuNZVZvLmdq3O4Prh2A
FKwlSOwOONP3JsvN2iIeccaoGHdVWl4EJun8xofGpsmGqgE0BnTH1a5RNdzC945QnAeufLFMvEDj
9K4fsbWd16SLiUtQQHr5GRliBs3OigLbEpIH2RoWYQq/X7hQxxeYQs/OcbTAKIuoCzrk8/lpB6CQ
kDPyNskpa3TgrlIP6Uyn/tvUsgFGB08a0g33zCYeeXSjzpo7Hcw4J/B/AlXEdZ2Hb146avTOAlM1
YDW/ll0G3amNqyeoA8smy9YMQNPo6Ve2G/60ejRKxT3NiRllPv/nq1hNIaO0hx4S4o37wZy1jk/H
sJQ+97Xi1TLPmxU28b2Eivb7g9+ls/BfMsWTxvggivYWzxjArSjHEFh2/0wsU9SctBGmlSDmT6BZ
NoYmnZR3aGm4w7CwZDaXUOYI2LInIkETt00D8hggU6T+WmmDHy4bHXv9my5yT+KALZelEE8bNai5
iYJ6RqMaenaBq/QpsdNBywXH4jaJViqNO3Uj3F3n0/dMxLmqoCcVz7hu9jt03JPEuFqdcZhgEoGX
FKaKqJzRKtt4meKg2Qxldw+DGg5c6GhtsgxqWWQApBlhHfEkb68d1Nu/iXNJznQ5CUmr3GvIdFML
FZENt7KT8ZF13JYkiJ0L3nBYdUSy/+/pLS5LYy2xpgwT9qXaThgi/PLMviUjObF0q2YWhhhv+8mv
3jQ4trkKo75PTRRh11dAPGWALXkNNHgD350WZnwF6qo/t5RbR59TglFm1djggVS6s3hskFmsPVmg
UFlVgQCRkLdihSIiT+Rlo1aJhUhH4SKHZ4snsXbl7fSM2wOZdoVxa9+v9UUmAksaqOnl829S6GF7
Q0SVVB2TF8/TPmeXnWZb8k7vBFsMRzb3nkViD1iTy2SWeWp2XB19rMIO2NTNVdAmg1X3w6zRHIge
6yjmm4jM5CozAvm3Depu5cukNlcbCbENoV5O7vmYnwrWuxvLe7sKTTKOSL/9qR6YRgdIfhML7cZb
QRsKTz/Ly2bql370O0RgiZX5JaeTz8kmdcg3sq+nUAacaotMMk2c/ly2zUKRvhZh9YIvBv0uw+0e
GP8njSdvszONA5dgYlIEFFzVznt7K9kg05pEFeCg1yjBLwj79v0EV7UK7sadVUjsJ4ExFYwqNOJ3
jA7hq9INy73xoJVDme+22GrOAJZfHqWpsnZYHJ21TmFmo6ksebowOzZVMnPYINtP5PJIzPuf355e
vHhUJ9G9jmZ0f72WbVDkgth3UFYnOesbLbhyHi3LNSGVjgmcpF+XDy7/qyIfNSYWeWAuKh5JvLty
0kHRnIHwZZcrIveG6kHSk9jyuV/cAVlPihzQWl73p28Eq1zH37AbxcYorLI6F3qIQ6hdhNijKel4
7VP4AhDOmHzUH13rXlqUmlqyOwrONBi5AYjnf5N23pi8QH/i+1oJBuWl5dhuUDtLwqrQ4n7Tl0vL
9/7ky8+AP4Y2wIVDh/X35CpyDmjiKCXKbnoWNO3Ul53k1XQfPfsgALejo5NSqktJlIRG5slkKDIs
rZRFbZ1Fs9eUsMJNQX5ivSi+LoqxF7hWEKQGW4rdIEPBbkd97No+guGwIc65zZBaecCtZQLBRW3p
P2GTyCrK4mbsp7tQkuDiaYP0WZ5dw5wpvwkkWp0bWDcmMquh3zA2TDl8knqc2bDmig8qpQXRCCE9
VDwD3vTP0zJtR+Vdrd9sxOKm3RvR09BKT0VU2XCnwL+vvHz4NVPeuTVa9qNaoQTEfx+di3bp4LKO
HqaM8O3OHdvG82BHX0gcL+FDUlcCh9FMGPa9BeuwnEMvmNp4XVKBSY6rZw+WaG/Z0Gae5VcUtdSe
YSJ79IMIGkvyX6K60Hh1OjtZUyhQDN/1pUXncNME+AdqTXYng0KT8O5+utWQhP3N12eAJc3dyUKm
GVMJJ5jJuimCB8TzklcCUpBRpKuRNs3FmcjLmfT4jq17VfS1ybz2Q8MDX0IncZen81Cf00KxI2zK
FKUbs9G2LgaDLSxr67nDiN01gQgk7gyu9af6dlB9fQB7MYYmJR14lCUPAaqSGPC31srS7aHwEuCn
8n81n/5BH/bvPpWjOdXq8XiKfJunid+ng1CuBBEnhKCg8Lv1ALInzy0yul0D37JOtIeUGB9Pa1So
FhGFnsJajQkBYlP8FL+EZXi9ZIfzgwP66tKExCgzlRudHp5nVhuRtZoZg1p7V0AbloII3ngy9IDH
YTTFxGh6j8b0H0hPdKAWQAeuMl64qd0eryPlP3QeARk9FKp+fjtem0hKP0QzJSPj5T2RKqgd6AiA
7kHYBjaqfDXZi77Ni66TBT80jYHPjVKV/ZK0Z70SljFu8TfBrRgkcgFi6kqy+aWL6qLKMyZouWZ1
jSWkZEXN+SKTv98/zUR06Yj6zIJeex4zAmLdhbxgrixVWzj4nmKitczhudOsBCogwOW8UeTvlqI3
fdj/0csJHsK23uahk6F2NiNYP4rTbKpkWFmn7H57Q6IyMfMQmwHxyPLZgSCbQGLjFLR3fvOvghqT
qSqeNs1cwd/6zpKFyqA67cv5fPBUmK7S/eHyOzBS8sMHz9knlp1LNw+siNp+HGTiWwAVmV8BC93t
FGOSPNcHk2PqjcRplNuBwbjki+sZzjWTUjTjuF0f5VVT9JDGbIv3J83H8dz5wkU/z6b4gbAm1LRG
Q9OP7hLrVErGfYaOE3uuRaPHyzrmNRZs8hG0wMUbyTtDZHONcYAz6A4zy5g+kx/0zqny/UUnP23X
E1Rlf5RxTukW+F1iqSUnTMJULvTYuTZ15RsKERqOKWmpwEts/iGEWTIundQ/TWSfE6DXqfcAij58
FANq4GEMdo31nAR4Onp/JTTuByKb7sBFDV1T3Jjr+qkFdKg/4jOEc0+0cJX+WyNYOQySDkGwuant
Rin7DP6J7dBroE3NQ+kAkUB0rFeqptwYtMeaCN/aIU3ZIwRk6PIcpO9JRzC4GiqQXg5nmLlrhxK4
bYkMoPSUYJ5wXfQ30/0bjqp7zhQ9NfqBpxUpg8cJLfaflnJyvnBM1HwEA+WxicAXtICv1FEdZ5jg
1sAcCYOf7mnxvo1LW63An6fcvxzxd11SIPwmE4MENkwv7qAhdos1OtwQNCsnZeoXz5zTiuSEVmQg
882UDxjTqTv5lrrGZvCr0+8UjLgM1zgt8/yxUYaslvynDL7/7KjWdQRpSQV9t9YAm/8GqphJLE07
OVpj0trNtww9Sg4VbJiMlNQO/X9f1TPxrciHFx/G/fL+Wl2VbimTkVya0JKuGHNCKqk2tlmMepPf
5nw20eZhZTYEwVOPeB2HtDPy0m/io+C4oFdiNkeVUDfviSz3qUnVTNc7H/IGB+zs4DMUIQD1Kd94
QcILXTvscWZNaM5DNXnORrDwPENTO3wJglTSduj2SidO11bqJuqIoak5qd2fCvAQc2cUIf8VcSTf
Fe3x0dXIkGR0ZJL1W6c95Xz5CUAfuovSdFUtTZ95sQPTp8XC4Wb4djzZug5vtNGjgMZI8/R6YTvd
IwI4DtvR4uvdHReNQi5w3EV72pf6uH40RUOgDdeWtwjqOHs4zmv01RSmima2LwkKQ6MVHWH2BP/O
Ty95Bidzj0xfzz77KJr3M7RFySICRb55G9vGZtZd0m0X4xrE0MLXqc4iDafvPDabrdARs1gwBIFe
GuxGLzQ5b2IccDiTIEfl7E59E4/uC4PxZaljDc8CkzUbXkdLQc2cvKt7ylv3aD1q65ys4Evgyn30
o5Vwcy45VR8BLjvDNm3BfMEwoR0Fb0K0//n0awJ9eURUfjhndlT0qmoW2X3wUIhmMg3z39qi4LtB
YIbiTBk6T8U1StT1oJ+UqFTSuJQB35mvDKF3uRIzZcX5TC4ryqhFkEEtYb1CodVIopftY8UDpRnl
PA6SRtSAA/Z4+lQgDfXH519Nx8OOsuuyI3y1r/1PxAGUdZAVmOL/3xCxQyLeEzXdf1pS50PN+qkN
59c5sLmzYestb01PcMDzIj2p8Jx9plIb/azbTQbQt3yU3sZQucv8vCJs2NGxpeTmhrhIohwsxsAz
3qtX4B2Ad9Ztec52ZkQqGLghEOlz4Nzo5fiMjFciMMwXYpIBckgHtl7/m0D7cAXDFvMeTB9tZ6Z8
VysahbI031OJ/FBE2Sq4jw9qtxdg3qaU96CRxSqOZLqUiWe4XSWo6+l/3WC30IBwwd9DoOba9kMr
m6TZx669FZuiM2AvTilH7dPqPpbbj7gx5b/Fy2saepEHRm+Hnc3RFOwmVHvCRyY9rcrfLjJ3BPRa
6DDbTUgbPwnJr23zyScVVFs0PLLvC9QWm+wLqchJZlzLeVOzQSGPaXj4vlUM0r8M3jBF6IzcIfj0
piNb7vswGzjikeKvhXwpy/HSmKIRszWsX0+jUQt6JymhnUsRrcNo7TjQDefXuFfHWabsx7hhRNYo
ow31NfDAn0i6p/DWLgtks7+x3xx9zgS+YM3xjN8VAc/Zxr9jWW9a6DX0sct83ALBDhX9c8floXZf
1d5toLjiStuJtl/2ZQKogdD/UlNuGth8g7o5IhlyO43J2eQahJ6XdSoSXk66608wdQ7U1sM0XmhZ
xR82m3WR9NKzw9RvLaVfkq/HDbciucaf1/g60sqMVOTnFzMJSrW6XlZIATuR0LQxncKa3CGIfLOj
NhPxzawOHmdqpFYP1iADz9ianExraD1Uvrs2vrpqeXkNbHu0YGS3IYo8qB6uDaQf1lJFXgj4ViPB
tR8s+5HAjEJfldQKsYq+57Tr3ts3Iaj78wsFpSaz/iloH9fQHIzlPDEwE1uboiHADPpGnHFTfio0
6okMIKPnX51I1XwGe06sD7fFwCA1M5SAIpXV+unmcyxKnkBRltnwnpsnoGcq299FaMRNJ9FMs74B
LMImgDSS1m/fevdNvhutxUTKSRh/iRykHxRpBiqv+Xw2TLEJmBC/Mz7ugV6OBnFijIHB6+Il+vxx
kB/gMMy58tKkVRHQDq8I/VLvtpSXtn5pvKXdijv7fLTUtCjOjjwdZNoii0vgPZ9RmzF1ygnpVdmZ
gyczcTS+qKkDhKJg7QkdI/t4koN6WVc6y4MVpcoNoaVkwE9j6lpvp+6EHxMGfSKAicaBBn2dE6dl
rf0JZlIQa/R8REl2Gb7f/KHElxZaL8VvAE4V/LMmtUF06xZnHKx8icz7b6ObFhrqFBT4y5faptWf
6ilUZfjb5kg2a/OsLpdWnM349LimKU2CQcjkXhNJQO3e2nyh39JXTyoMF01H2+sm6UIvwGjOUo2o
qugMdYPWs1aUaUneAQtwHLGSoDvS+k9VewwBtxp/L14Bwgy3exTwQIqXCCNfZ5FFQzp5EaBaBvsT
BRgvbtv5zFIHLIRVCLsscILo4qu/hbLcwS+Q+6m6IN7HYJnzn7ezgLaysOlOVC03bKT8td8AP4E1
UaSCdUNF4bN6lcYiYy1BL3/+8Zl3dELnnZ6NXmCi/Yre8ebgzaEuGZQZWe5VE3XOq0GQsFPE2B9S
ZNesaAq4NofAZSvXn1KTF4svYsydG5FEbSNHm61S3CKQ3CyOm1gRXO2hhqUgN9bRt0q4PXQ2qI14
jGUpbGJrnN9qqARqPKa9HsRp+W/ATOrGljNIsdwASqZCBg9DL2v1o4RsUFInghVItzylO0utpFPs
cciPFG4F36w70jBQByASTo3dydRerA+aKTOhWimJ68q8hNBxDEag4b8IHeS/q5Wv41skjQG1TSrc
eUi7ZabgRksh8pq8823A+sjEIg2H9Qk+My7bUnA/erq3rtDLOyCcoMR3ExbBRjNY1XzU+K7x3TWl
HrhMKFaN0ULfzhmCrJeZRHogfm1v+nTqslq5WHwdQRIv1z0fCeAgd1jc7zBSf562LJZSJVjJ4tqR
GKDvV3detU40Ef3xjPDjU7enZEYdLA52mVc0uULX2BnIKRmA6gxu2NMQflYZARs0PBG1rRzzlp23
CjUxDHRHxxLalw6ZOuG5mXlenmXMrg2xTAAybKTEFDTo/P7rVDwkoSQ5FbJH8DWdcykilsfvPzen
SNpIThY021CHYQSdRpSpi5vnzmNc//IkeNU4reT9HJM9q8QNq/wPszclGU6hpz6GIz+z1ff7FjCv
FKAS7bNDG4qCK/4ykBDegvKeL1Thsc7arJxW+51mNDQeyMqdE5+wWBvqxLz/iRSIhzZ5A+6J7JBl
Cc13MZzUTvLJ4d3TGoN+EiCyIFKX84bLIzNvOMLLVOq65GPc6eEA/Xt0RSGlnMhfd23ueMSRLwNt
3kUzH8m0A9LZoq04IAquNWSLm0iOxLNTPuIg/HUdpSdKAenSYIepM9dehr4VgYQfvmohjxkRSlUN
JNR1bdMKD6q8ZjCiqTppN6U4QJeKwTtyWBcZCrhPOD4bBIDLFCMMoop0LTh2GruGMDmHFFmJXJCd
fVHdqx0rG7mtb1hXBscfsTYkq0YLTkbc3mprd00M+IO3T7cZ42nUbGtmPffLk2/iXc25nY6A9uYy
U2bM8a3WazB1Sytzc681IczDr/vGBK5jHIzq5FLEU+p4+y47ZFRFGuHaQG3nYnIGC7hAkYu+TpSG
eci7IoMnOF1nwCVWVmRgbv3y45JYTlKMFQBj7+H8ehfOVizxKoAY2KGe94zl34gGb+HFKB4QMC1K
9ugO0wLwFRZ8268T8bQ87Y67FwHc1xCKEjr7IlYtPuDxwGS4p7r/sLFA11Tte7NRA9v+yu20Sd08
PbZyMWQ5F3/TgSYq+Fs+5yA43VB/+qYNLS3TSrSxmxYsyV7Yq1rR8SAtNn55D+wBfqIbaRpCSCSI
AN78Us9HgQH1OEiqc1cyWLY8DA+juJyfaRmViPLSvJjx++T/UyoYRvWudlkuxKEBieit6w9/H78x
ZyyeYG2i+SaXGlrbxbzgVsMtRm68SpSsc/4Sm410aD4NrunwJ5u8L/Vs6JSsN8zzRjyw577526P5
w64GJ+zvniWETDQh+OwkYGTl0NXiKHdN3f1EFtmsmZgcM/CSl9bLiIMBuB165+/SmhgM47RD5Kga
puSHYOUat3sO2/tAvOH9eTweEhZjj8F0ZnkA18RaP3v5zp3SjNxqWC2m/CTruUnlCA+IO0M4bfpX
ziHW92TGg8xMZXiITUdwCIHPPQiXL6v/Ja3XCNt5LpXpbIzYqG0ct49ssHyIJE+tVzNrPvjLwRYs
qqtnixmCt8UTLR9h89gdFUQx53CFhRa7FNWvY4ZPuwI4u5YVtOUky8+vnPPdQZg/VfQfzVqpzSaq
A0vw+ioF7nXKhn6KOLHnqTjXoYmR1w3O1LAiMwGFHywonPyPk4I91acJ7RRlexYdLn1qRDQ0mDTS
ecaWXU6XK8Kj6VyGXIBH0Ft54k0iOzZ5HuFyDPHZ44cwI0EEKBICmQuSD/CuHCAaIno+q3FgkKuO
dWjpTB6seFwWWFC9zR+D7uhfBCVIOVXNe8Wt9QLmVr/pBnWZVOsOrnHdbf+FuqCz7qwnlqaADYus
Q5Hbr4i0/ySu+UZzX2ZIwnk0Ivj72uspVypHNW88jrgEQHxKCGMm3q0oxh9aAkv08I/tFX8qCakI
rlZJY9gf6O64lns2BquqZsZFNjhT4ubeVrnlew8txrQxoV1Bwyy4dr0RuV3nhtwH8Y/vJ9spAcRX
6tGSeqxqSMEQVOuU/3H2IR/AQNv/4BxS7jA8uwwCpRBawgR0TAxYHFlPEnv1ni4iPV03nNkYPe5V
1RsvF8dO/vdvLkACDoLxtF5RVYUGmgF01IAukupFMYyfSefo0Y4M9LgMDXmVcr4qA70To6FyyFlu
B6S79rRya3abCoWvWcULnIGcX22vatN9b5kRlQZNkdcQMqwK+gP0SEQ15ebuIr58R9G/25deTgjX
ICcnQrYo+7Xb8ftUBgAEowKBMIIHFecma9oY3TvA4/Rk/Z5bjE+H1Dipv4RVr8O3MKJM/e8AX6d1
JUhi5jCtVZ9TpH//cCe2SNjJH03/QBhj4bZATuwbexmbKxJfeLNHFUP9f2eVssn+Xu/1s4Aqo1kQ
31GkxqcmrsFC7CgsfW125JGV9/ln1h5xKgAJOzzOqNqBVLsXkQyKMqh+dO7mIY70JltVlhESvN6J
kZcuKBD6AHGGJB8CHZ6f41tzQqqZ3NB/a3hKwICH5bqZKZPxH0HBLpqMbtcmIWgVM8gqewl/IEau
O58jJXfcKeYEeLtXQLHKXMGh2be9CMzyf1Ohuvq1qqQjXqmx8xI/SViuhxLBrEAfvUn/MYlzUjA4
MLUet3I3jGKgpD+6hNb+akZh+IbH3Ut+xK4M6fjLQEXAxczRd4eQ+l2v2TqDH4Hotc+xyQaeyOQZ
xA4Xog5z00G9pbIY8um/CIz9inlE+oAsdPIn7lOiMUki7KAWrhpwtmiV+OLPyo7d3yyXJko8bG+D
o5B4c9U05X6sOAR1GXLJuM8n9s8V0fA2VQTozCc7Qx7RLq5zKVyb4YyY4qAa+rceIvLPHD8Co6l6
SFhw0zRo1SfJTLR6THa5lXLH0hPnXRubfJmLPdm7CbsQdSzSAC/WaQrGOfXK0YLm+MG4KjFvtenr
unx1rbti+wSdKN5ns12k/ZSyHjrJEHDpLtVoaPSSCXp5FeinRUpikW5eKz2yQ+J2Fk2GG3oqsvmv
8Q+uERD7sT1P34HsZoXu9I8NfaYyYDS9VPW/cdw2K8S6O3aS3fok4GWXCLdOzkpfwMo0bR84dKzc
Li2Kc66a6W0ixv/ggVk2w0M+gMLlbD/iJNpQJJ36wzKnQPMAbXDuH5QsM1ryqqF8Qw0SX4RVEqMc
CFrECw/hHkX11/p4i9EEh81VcRKoRJSFfAXTt2Qx53+K5DMj30WvYk4Jk9SBSaee9lqm7dxQHuhA
aP3CqGkOHDucs20zV4CtAXYxfl0ktdGCAWnXmFoUiVIEQ0oHc4lYDu38RH8r5m0IiPHHH4tvyCQ0
fgxyFjFBKvxunShZZjF/LISGYtoymS2UgiY1X2KA9iWfyq5q1R6hTq+YACAEOBr//091MzkIK8c3
FfWqaelKA7Yr+Xj8BV7aGedpnrGrUaneiL+Y397ebPlzM7e6Yytu+qQLBFtR1y19EqphGtHwZy/h
Db1w+LkSRtTAU+IVElucFEpBefxf+eFdG0sjZOF5mdYXsmyqumT0aygeUKLXQshbfng/YwbyZcoV
KYAkeyPCL8IJLjHmDzW6ecqG9M4S87WyieGzmraGw/2hN2KAp7998MDzTCSdf1R0QCbb858wfL9K
+b7MfBY2HyFnTNG+lP/mU7Exm4wXDihOV9U9MY8UQDekp7EAoFwa8lIQ4ZyzEK56bGeRizoZMe0W
xHoSSRZKXpUp5MMPyzPFEBpl0k1I8MZoJ4QQRZvAlnfE/pgMRb/DFYQwZCGTxm27qejc18B5N/CS
MYnXu/PytWZvWSqtDeODcR48EgwlxINB6BYKLe8mfd8GLn8MOuUpNheefFqTfd3DTQdRCvaeLckc
QWZzAKyRw30+4jl/klIOyyhr5TvbfOO17HGjTeSwKcQAZLTCD5XMHh+f/Q0q8U2SR+HGmnR9tMra
Y/VNaB1Xqos6qatB3BUCIrDV2N4OijCxZCzcK2p4JJuJ1hQmqV0oyVnMq7+VikgSDxmrAND8t2FE
2z3kgfuQPZqRTbn9TfkJOtSX8mOIxspfHgwMJyLiszyCFs/tUUA+KOhbPao8o0hkmmlQYUDR9nOD
vHHFHWXoeYxnfeEfDZTomMY1kHYTe9xUWZcN30QXV+7SB5DKr3rmNl0lqjLImbXhIpLV+SVyIBeK
OvbNh+r7MtLoz8GvoQn6Du7qHIm2oHnt29xi7cYm+DEdixVwF9WcBoCQdCDGFaxDQclZ3vvnya73
H1vAsE/UZDEdtEJnrBFM5ckL9coley/CNSlRImhWyLDs0bglrSeLW4E+lbPDC8HVux8YQ3ybmOPC
vj9PeOcHnHBpCHkGrK0nPvdPhkoKuUl76wbOluoYFJU/RW7ZpN0Sxj9ZFPq/fAxgNxm9x4kvYItD
ljpwebWL8y2P9vhkDYlPECoiJO134XyCtU9knvZHw2uxv83pfNE33l/2bEF9H8y8EguL+oeVi2IL
K/jyONxi9bi+Rww9W5wHXQqunDbap2/lEP9u88HzsdaF6bzDf5Q78ZUkSamg94NItP3xOKFRgjcN
CDaBxMGuLoufv7pZ7pZzh6MdSBtGHH2s3GgocnDYfj856UWadNxfX6mvcI7Yu1CyfC7boR+z8h2o
+N8OGlMArkt+57v7PwKRkHYXSp6+ao9Q6fbuUww12gwDgVDEHz9sWL4JONAQ6zETJmVb8gW0hzsU
GdmELNvuWWmXKabBuziIb22EgLWXMeaMiKh84+YxgSBGHeELVnirbCXFgnzBKQgAzXHYWeF2eB0I
o8cziDTlYTyhmv5k4xvGBgC2XJb3AUOHOGWCTCEF+Kp790IMcqFDhQWXJGphpxxH7ww7aXfoi9DR
ToVLyfl9ug6nAdXr9bH0rCJryHXTdM89nPqQaPN0DqViH9sCs2WguwpV3Gfckm/oXzlHX3zHco3X
fNSLL0jCrb5AQZTGW1YlCFSmKVBOUSDqG9C/G5Ej4jZJoUhnP9v+h8QW3dD2Wsd5FfAwnL4vNonL
bjyKiyOJlpfGC1vXzNvn513n0I4VMCqG7saSZqEeIYmeMIAjFXuu7/O/zf71BZf5lqsPJRxl/YkX
VeCokaw2gOVIg3zmSn5qQTEMsbZDZPHk8ZmKBgL8NTazSLaA053Lm9/SPMwx3jy4cf5pW0YGM+nC
YMmIe6ppJH/tHk7zIqgPAV8N8qDwnq0Z3DbKMxyt1c/a0xHKh4g659napCJ2ZJarlgSS5dhOP5OE
a0tilfDE0QXGCaoIIqB2m3UHnhUltoSXXK0BcqywuIVSaKT9ojk2KLhz68rfF/prl+Zb8rTSl2JI
+BBOSs+IBkEs83Yxs0fksr1mmAS3064+ZoJOFEDfIyPPeyycr24Df+HXneOpbHSgfzf0+92FPAVn
H46h+QKCc1zESLOS9w39c1z2GBypFki1o4jNnzekfpJ75VlSOEcftym3mWhKI4bE9lHTqsaS0uUO
TAsBl0drBsCi2oC7GAm9/sW6NRvMdYDyK65X3l21zmz6zX53daFX5gfQnjGRk1QIvIrZ8pogPnkA
hDIiIgmc57JplfQXxRw3Ts3dJmX8OdUBN9LBGS5kbrcFjJZpCdu8G6BuLnBUo7zSREg0lnGnoLmF
dsvf2XLQnJZ6FLxCDBW3Nr6yF3r2mVnoZazAnGUkkVdHTqmNIBC+qwq+j6NAZhNl41HJN/dgrWYL
RJwtPBAg1wCVvo/+iaTHvE+jc3QULghP7UXaRYFGpwXOvNJy8+tZSYQfy1SHvKTR3xcIrOVvWgoc
MOPwkvrHk1lfel7jsVCLlmUvhHA32od+a0mWJA1lWMfFHIlb9LE9XuOk51GnrdARqB/az5X1tzMM
w8bj6zqcop9ASbMNvmriAGnRWER5rdGKo9+HJJUUh/4Vjan2bQFl8StEjAvv2C7A9pS3qobmlETE
lsMKY3tAmnuxPbVIeRIA09w1fExmSXplaYc4OqKsiV8VcEL8pTPoUi6m3bkfNguSmBS67VDxcaBP
swJwE5TV234bNGDUL2AoBu7XKTi2MiIe5a9MUyQPV/f5mj5SWCp7CxNve+LLa6Rp8yAcqU+tF0JK
ExMCmqoGUWqYy5Cm0ILstCw0a8Gyk2rkX0MsVxNEKcP+2PunLOZoHxWLnr8IcphoYw4lBWzsXl9R
txNFPrYjPk19IA6NhG9IpNBZ+DrE7oHHh8mhnWWTHkBjJvU3AKqZiJR6EpBNUOdiRZftfZUI1ygZ
P6GPlmU3EFEzv2W4P97OMoncZoD6F7GwizvbzlYDMggjnk11V4d31vp10tieb1sjckvXy6Q6A9vo
FEg1Sz/eOvDP878izoUbFSwx3jy/e6TabOurCY9noaaoPK6sp+dkYOZhyAJ29kgQsKV1FzMjVvjH
hN9mp2e6r+7cyODeIjqykOKr52jA1bezRHxZouNRZ0dZlcjje+FaA1AJRI+j5I1k+/GCz0+icViW
HPMUsXLjbu+i8hA4eHLrNpFeA/66hutqUllbxhEPAyQZRczmQtDoejCsFxDj+pu3nYxVdwMpH+Ov
DzZNtz7RqywpL0PvCMPdRpTXaPsKkOHNTsFnoNFssN2namF1in+7UlVjDs8xbRomxCKpFzF+xoWq
RjlsI9yBmMZlULKMHUHkm0jdo4m8hUn+9Tpf+5q2Q9s9acK+BlhgqlL3b99l08pZtiiyepEVlYub
6bJgtdm4GKW743UvtWuKLv32dzpAiPQm3xOG4ye5Rqt8NrLJRyqGZxxFdFAikIIj+jtdOKGVZq2x
sqiRQBQLxRSxeunmzGpbFJBzSi/7REz5n1P2mRavumDSF6MWx8GX4jEmeAGTU4dPWV9lPxku00ON
L79qGHeMGpkkSYgnDcHyTOq/HVV08rZR45RI0jeYTQIX90v9eBK2P9q+B3ssGXAoCXsGNVQc4yNs
Wxb6Jm5HbJ3mGhzd73atkFx6oILb4id4/XJvQtlTU/+Sgo82jtU9yWhnUZFlpgzpVVRQqcY33J1G
BnSWDz7ce44WLSydGiDwPMGXkOisBnqGxcb4dY3soUXAWDAsc+feQw/pBNNByju/QCgKTomz6KJy
NRlBMOTCJMax+gku75MvXvwNi7SC0pg18sdoQjfcrPUSwCxKiWEs3QJ7n7dVdyXEnViRzu+TsQyH
s77uaLMtywRkq+mt6s7/Rh4dacXEdkOLtkhMJGRnNLcrn9Eth4uOvikq7Ap573J22IN6W6sKNf1m
hXOwYVb8f3OoX5jDT83lnlsVmHtJjFdy5LvnFjFwNAqN68pNLqUi65U4yw9BNURu6+nqedMQThwM
b28U3KMpJZ8T0Bxdtezhvh/IECZ6Q5C90sUI1owV4JpmZDv20ZUGgVpYn3fCIqnTvqAkWH7QPRkC
G1miexMfOQA9NVrO7p8oAHUIZfmHpur8kr0E00r6B5m9lWBVjM4UFZL/oRmuQ7mWr6HUFbkQL2eE
ZqO3Cw4OvHzIB/0iX24LfMIynRTCZlT50SneFetkKTkxrACd6vlnfW0SKMAXfx08r35FtIqU8W3Q
HZ/wLgji7yE5E4t/jb5z/sqOnS8SrPPMM0AkwcVpoy4oYtp/5wql6tIITSli8B1qRJ9g0WM/kt6M
KcB6/3FA/zY2NXFjhHJyODJAW+ZU6c07BdyPwK8ZGytxa2Il9m0Evyr5r1igiQrOzREiCQKBen/U
Fg9RkLwzJXXUv4ujCZe3Ar+WJzdYfe6CBC8X1Ck707cWFzSF5cqJV0vFbSWvXjigELwNLtmbgqfZ
9OKwuvKv45o+xwqkVPQTU7iWqX+fGYMU+NTQrfCvXjz02ur8AwmDoXXLksLu13uan87uD5ylQQN9
ERDllLbeCbTr7MvrGwA4if8c94m180IQTWWsiu+uetu2Mnc+7gu09b7N4rjJiBnssW/eq8IktPzY
4xxGLi5q1y868cf5uqqMaCELWdyztDrmqKndnYuf+xO4tBXq2wr3+/w+CydJYuXa6lHIvdPA+bQn
w4lNq0f0rKJnavsNFWJi1mTCiIncvOj6yB7XdqtLnwtQoxegZMVRQpgSEKFZOlJBAwDB0JCsRgFS
8hGFdLV3qkAUw9tMZpyTVm+OajHOEwqf89fuIEoyliqkaI4Dff2dbKZdT2OalsF5mmL9ef+sycWU
en8deOTH0wdDF+DT+EeET2QwYs6OJwfzsfbSRM/0umVLZs9FNGEes2Zmif7n2MvyTsbWwkFwcbfC
lamvge52TS8yWjUSpIaAjJfYNbJ7xcPC7vKt20yUaC/FgaFd1PVbBsJNk+EsH+5+hUSCVUjf3+Rr
ESO91vY75aISyyy5QnJJesed2c1LxzvF43563z+tGWCtSoRS6Uc2MWrxyz8KDQPke7on1glfrCXR
FyjN9NKIxIEleoZ00i7HffGsr0WTTh8jTpX04G+tSIvl3ounIc2kAseol+p7lgvtDVkMjUFKmZTt
3U7jmFR5U77SLzmkeGDlgKfDifAw3WuoXObnKS6VoMxiLxnhguxBZqBb5a5L0eZ17qebdV1k0/aY
duttPbWtGziqnWE8sgsgglNT/EZ6wDTofXDjNdik2XQgjXudiSb+xlfhMQzxzmUyrbp+BqhrxH0y
oIiTtarrX8NmmsyMv6amriAB1YHsjeU2sBqZifzQPNA5cvPzIw4nJ+3accwAwB1IQgYW7eX4NuYc
m0905HuQgzbz5w+PQDdhPZnaNyzbtUGA1C4arFuC1tLi2BXAUhUK/QiNuTk8vM3xFOm4H4NdiUMI
XJGGKiFqNxj33SU/5HWvC+cZkPhdUWtiGMFch3vmYrQhVIoxZF2c91vzDzm84rtvv3xYu6DfWOcw
tySPl2+kjZT+hPfHWHlK7DYr6cR8UaF7Iy0+FYS6dZIDZ6/5AIYWmPqW/uDW6ingmXKA/DaPnDd2
q5k002CFHnoHssXWiYdVDrwjRveieQgrOxUSAgC2Usp+1gRG3QdtCIHuvDxd/z9mDf55m6bbIFdu
b5oBamzq6TsReLZUrdFo1y7Fqw48pM92QW4wDbGPgokLs8olHqRs/1JZm6nSMKRUcgVl7tSesHc/
rywNn/+f7k7d0fritHNwmOz04E30sxBEMD2U42310SgjzA2zWUrC+DCPsApLoHefzzE1BT0wDTSA
tiAtTv1qMov9TKY7XSI4/CdQUeibx/XpQofbC28FQDIfAQpBUASeBZ6pz60E59VR6WicRFZXpl9s
Dp1E7RgSNAUbn7HOO+4hv6TlrYSNZJ85NnS3+alHi1gXFRRhpp0iNGeNVQU4KMZ53xiL+7NWAyBD
hh3XuLw9QIAy6cbZt0bYd7Q/+OjWarafhLR6FZDN3Iw3m8/tRSfQSuEucZZR124phtYRJ6ytM7LM
ccAI7qrQIA5l5/ckriGtqL3mTZdUln7XDJpEJ+LoT8es+WMKFbE+c3LXpiV6EWsr4B6F24jW7KPN
2b8hJR6OaGZZ2c7uQq/3GcOgSTb+F/v8bEJcYbob9TO9kKABLyh0qBshQxI1jPRB6wIwQ1Yvm64a
8UxV2I/MFZhO6+rbMt4fjl4mr+A8tt1pKA8tvozXqwdop8D2sGsoL6dYqLLjbYTeUbotYat/DegP
BUsLPeAegozUWOXAZa3dddjSAIIpNLiKD7jRej0HA7RoFPkL8WFAVyH+seWnSVC+Z0OAqfy3GzEx
IUil7vlfmHCfdnPU+pz+fqV/35v9t69XdQgByAq5mzztIHlvWxwfP+KtVetPSq8btJ25RKLyE9ae
RX9+0ydpOLMWQoG16g9KcsS6m35D9R22pxU8vpz7n1gtcF3LLnn+dTbHXUOqsWWALZhGxRoQmoAh
u56I1xgH7Nlotw4k7BjTc/uvoKeepegRRCPcOnAxHLmCFxRSEFdFRI7BrG1YcfGe47GQoUSXaoxA
kfF7QwLJF2YYpwew7dvU6vJXEX604B5Xjqv7rs1wlF0rbQSKx/6Q/QtRrORhI1KkRhRu2jOtAMSq
ZYa8/RBROd9a18z2lmTW6DrI82kUR7BDxNqak/sxwydoQWD+6X7BGRuYl5+37wcm1cc5n7MdaAZy
GRi58TQ13H965SQwBzRMHiPjsTmRufzFqVZlNIi35IXTgpeuqNGeFiMh46iP/WFDEbhqYaBvDRsJ
WLBxr69ENrVc+EgMCOkE1OxMbG4hVv3N23OKzP880LJq5hhwYi1/rRCHwmjnV9AulBf5QZZEa5GS
cYymXpbL5JuV1MBAy7CTDep31LPc9caGT6L9B0uA7vxayGYDSv5wULc+dFcyxQn1Xf7Fll5k16b3
se8VnhJ6wqi89WCZdQA4IW1pRg6fQcc+5JGeTt+aTrt95yUVQ96wjfanuMKfizkHfN9ZbDmTWHFH
EOZHq3gSm5WbXBKcri45/XUWn0tdFd98Gea7BOXBrxs8AvAktjaqRBFfSMOqiqOf8+tgQUH5agDm
l4kBIFnZCaE7MxfL68zea/fNUquPpWstYgNllruAezhq6ilGcgV+g41HWwyiTjblvqbDphZUj9Ei
0sLVFViJJGgylweWH97etAVydjUZdOajAPwL8zlX7sp7YQ19IwrJtDpfyasp1yoYcK1DJU2dU8C5
wbD48mvzcFwIy1Ys1LP4+U1EXaax/B7EiWwiHcpBe5RSf2mG/hvBnD9hPsWm06lzagRgzhVhhKsW
/OdJF0vzMh7YFs3v4rb0PEIe7K7Jh6DbMxQB/42dPfPcKzQ2ipgJrd4dfBIznVH1A6OTYOYALD+W
9ciO+bVeKb00oTLofHSYKR8uMBixFs5JZZ8I+8XgVjlmm4Imc3VFXOV6ZqunJBV5vv5AKpIg6AzU
7WET/WFaNa4OEHR6Znaf/lQxkIJO78qX6hfRiOKW2hAbpQhSh/i2E3lC9sFL4uCQ6cGWOHwNmO57
BtlCFAPJaYlPtxuUuRWSq2Oy3ez72NmsBzVfoqmvhhwDuoWffaKKWjT/YJSxWGzSj5sIbpvA8LvH
Dsi5rZ0I6MunAGlxMERkqRpUMs7DvocfyrRShnXzM9JahUT443KzilOlSXfNr0bSW8kyXykoCnvu
Ld+vuuau4n8nlnxIozG1/SgW3xyRpotWVNXcGgj0Zp8ztguEGslen0oNTYu7o3Wm8b2P0GiKi1XL
ntqEvOntz7tiQNkxt68BNerlJkr7pEDYlsey5G4QJ/5BOGD82pcc2A9Ql0nudswISgk/nSEXcHN8
4Vhcw7ph5kjAmImzummy4HxKb2D/LQIw7X4jQ0S56CYdIUeqy+ejNlPtCdkB2uYfqwWcr4i1BnKW
otPLgfud28qRne+c6aCJTKKulk0UTwyGVYSGUGUJZteSvS2KKCaSo7BnUycMG2v32ELTJyFtnR/x
ElThgNp5Cs7nwiiagM9mloB+Riw1v5wlTeBEG84k/fzK0g3KmClRn2rcpjIU8j+tiCCpodVIsHSX
wR8L+3p4738T6qobN8ryMInQpxxFcjBd7rUmGVdLgpTe5+F+i66qlB5+XfoiLW+RnbHIpnVOKM2Z
hMprA/Bqe9b6GHaYrd7Dia29ZdRWJgyKre9VezRjM5vfVqyaHy+IUfmLvZg/t6fKag4uYgkAOJ82
IVHgPDqbmmEYE/m1TZM9PWTXzRryI0Qpw2OuXSptODPQd0jGrVJRmfqz4yqN5WPvvUdI8t0vYkBv
Ldl7Cty0sFqoTvOWuBKHciktTW+ZOYPZVQqosRbRPOKNECqvjR7RLjipo3LHCZjB0Aj8JdV23oMf
PXmf0CNt1nljMhXoWS0TUKOIyMZM1lqb04t21GZP9YfQzyfguOqfdbJsmU2xFCX0brUMN7wkIC/T
49JX5a2FpFslg+RBgxVvU5M3Hh/Wu99K+mmq3RtLsOEWe+4pwPDAS8tIhfOgn0JRySPfibc5exlZ
5OnBer9z81IjTyL37doy54mXj+wxfWO8ALJeWEptuSi6bVq+WnglYvJ320E+ucLh7ihaFQndBbIH
WeS/5bhC4XPVVQF6cBCpn90plPYssvkG6ZWa3mUTBSH30916AKsDcPwk1TObxIEJ5trHWGSZpBr/
R49bvMrpmroYCWjCztXWeOg+VfH2d4TsYcFPwXQ2tbHO7hb57+SQxymtOfU6cktaULM4CDzR5mkD
OwPWgK6zQlz+7/D0eSyhk+zWOvwSKAD4hm/1A2LkrPv1B7Ks6PpXGMkUR43gIqOZ9iYMoXDmiW33
YstWRxcDM+IKPvdLYFZqKFrNpkNsQHHj69rVSOFcDCvaEx5dfqHSCWTgD17DT4z80D5huQnzdMZD
mmQKIsThPwfE+WpBsZ5W8pC+5GXTH09FixrOvNyVtt37O8dcIaiy1HZTYTK/gCS0pvVIO+J814H8
Jx6Z0fY82bReQ6d+fF6RGc3PwS1k63tN5SKDVYbnKdka/Y7urlaaLFgIUznoJAB92UJ+mnVsaImH
a2PdSTu+fWyEtiexhhG2M+x4hmfPyGJ1Wpto2aK5Qd49SWFlNC5Buusm9G58n3VAqISTicataU4I
OzQgAr1SXS96GKpFzoZN1PLw2/vspPuFJUnqwdQoKlUhodj/VAm95fdezpD6Fd2bwOY8GiztBdh1
/JaJ5wRsFl9L9eKxT8zVPqovzOx2IJ6lC0FGqHWt5+gCDdixcazmcyuCpyTYYeA2dzktaJkTdpA6
4+V+AhtLeUYsQhw4agHZotf+KmJvhpy4lekf4nCxtXYep+UwOkVc6p8YvP///heFOJMnVXkDK4sh
SxLGBAANaiGgwcZAxPOkjQeyYtrBCIIbPbDRh5MeOKsCowzmIKcK/Hho6oBEiqKULKjrWtPinXA3
ldi1BEAih3e+QKoJ6XbOyWIPqr5iqW4ya1wj938izcIXrmez8DEk3VO+I9z9qK0lZ0i3t28Fbwlp
E6v8eUrIje0kl/288VutdwNgNrY0XtMZgN7cLVN1jeEy9Us3CY1yHR7OGg9q6iGroQ0zjnkp9x/q
G9gC+K4lEB6miME1NF070GAg2RUHSL+Dpxcf1OwVmDqk7sZkJ1aPQKHDMhfDYhd3QYv2AKUwAxkL
JkAjnu0LWfRqiHKqaHLckMZdYDyupKmg5sXqvnOfTwdvPXYE1LQHE3WOILFNfBPBMepMhJh6f7hc
SK6YsW5ZCbGcKhyNYJ0MbQG9h7x5bcodzrLmeQRyr5MBurAyw0bghuoUztUOottepKTWbwPiJYvs
lKBGm2O3Z2WvOjbt6ajueyNbhS3bXNVL6kRLexCcI1h8fOR3rpL+7YBT6kihorZm6bKeJh03kcHZ
/rk0gSqp5LW6T0Aqqcu6sDgGWJSE6JAqb6Dm+59u4w37XcAX0t9uUl3BPX2c9KOOb+edVtuxeT1x
9NiHlmBcQV7LDua+wCGIVU+TJDj8ZRB22Cq32lI9UDvgkOcYUePcg13f9IrHHhpT3jggwIRa4pjP
5l9zwcBlDqkuWb10FeGNATkygN7Z/vr+fqavBB4A2uoEoqyzsePLIpLeoB2bmGcNm0LWyi6CaK06
g+yiqfWGMdAmEfsy/3DHSHKXtyDNYge6yn0qBJmYYWWyx7hU3Igd8mVMcrsx3xpi6X8lk9JIdmNu
CGPJMh5J8Q6QTWvf4MwR/3Ee8UPDKSppfhKhqGi3qrzFGycrNOTwluFe6NUozuXXd3xlZGx6OvVa
GpVVr1JONpdipbOySI8MZ14Qf8f33ZdcA8zfRhCvPVFRKVzOQqodzpLKRW3UltsO7byCfzS14+JI
AQrl/1ass2lVShzHhV0JXvQ3m/WxNxQdQB+RtbpeaWJMKc6ZGZCTQvhlZ2NqbXQ0+6TM+n0FMXUF
sfnD/I4a+FGfAC7xiMZXI6f5yiZx11mQjhBlpFZkPXPM8DVwwsbbeZCZuhKTVCxWIvizG6RopLHT
tF1qUV4mju+yQEBQLjNY218zoJNzw19sNWDgySBVR0oe4bPAR4RQ12d/5l/KtFwjkyK2IiZbzBxS
qsmu4IefaDFbh4gCT1gJ0q+GfRNrwsoB73VVnxvDfX4sFxzsA6fGPddbSqNnMEIQhZyOFZsAohlC
lasdJmEEg0jGKCDqDwzWSDse3QkSMorFSotctf2tUjiBEkbNb4SHSb9oPCxzVzO6Uma0KZRrJ0DR
sdgPqYK9CQko5/RtL002Fe/0a4k6wzSTRTDXsm0dHophwAKZjdPutpSQaTTk+LhgVmAC+iVwq3vu
R7VhqVp4yXsOXqnyrVfzn9Qoht/qHPAVl+hrz14N6YI/gqkXgCxXWUubwSsDNa7eDML5bs6i4JwQ
cjjOW4Z/mur30jIrWC0yutsxpKGRW2WPpRqVuB5LVavH9nasY/m0MtYnn0NGrDt5FVH5WRkSiLST
HqfSZjMTGVQ22NtuvuXGpT3S/G/N8/VJcjkypH5FbH8f2bfismuTNsns3PxpjSLMk3oQc1EfetNW
TEPo2e4NY79ZBb3DhDnxOd8Gnvh2mQdXLMeww+PSXpGaRD/5R0+oEzvZxRN9zzkERWLG2UJvbMSs
YYKDNrP2C2pUQ15xfOYr13j2o9sy/Q78qLv2BogwqL0sPXftwEqarryN7k5Pk/5gzkcNwRO/5nKt
2NkxIOAgmQHaJtjZJ3BlFI9A6zn1+Oymlwrp3A53Q7iScQB8ODAV5UGXgX93d3nKi44m0xSPmZ4I
3lKK63pYrnuRkyMgpjpMjOHK8c/LRULWsGGk30H3UJew413MJkI9xhsrZWvyUUTSJ4eM6ZIJ6ub/
SAYJ6bZoz3SLB+IY70rY3ZGPneJKZZLUX5B9SK6zIEdpVAdJjEfGI1HchBXKIszKDs8u9XYEHypO
gPB2HxEPhF+kdNSlOavON0GRGF5hZFwGy8Zlw9SyHuklCHtRspNTsrE4rHZCr2KoYzothO5d5rG/
vCFsFFE9nlz0dIAJXUlwVEr2HEP70CX0ONW9qwjgTwOPXXzocyWxTEcrxjbNekNCdDnbJdmRYDNF
9ZquFxvRmt1A+IqOxR9piuFY96N11fh/+T86mbTFy/iqMP4vb2RwPWqn0EMuZBn1m1tn5TC6Bdfi
bvNSB/+6qRzA9TM9czYsAopnKrDIqq9Cqp11TmiuDI6iqCEc7ROKtzxHzWUhDxyi7360AEZotNYE
h5bB0zjw4c3XTZO8M5FBSL1VXi13D5y3fwYyGuAGI7x8gOiDrAYQMftcYS+94GwDz7977oNT7ccp
VpBvUFQf/2357uRonS6ZUVQkpfyEurDtWuKDlIt3XqCQQhZIFmjhqQ7i8tB7sNIWPNaJgmMSlrtx
BYGiKhvuqd61Z2YW/+tnSxLAsIyVmCw7g8nI7qfaXIP29mF0CdFqMBiqpfADpSUJ/YpxcgRAYaVA
8Pb5HgZaSbnt0+c1NKhwW/xH73co5s65P9jM5o2BYJW9fi15a0tUMYaRim24W5DA4hRr5tY+I87j
Pn6FZhmoMoraUnQhMpEj+L7hl+CnqOFWHRk5fu0E2z90eCKZPwslKXjX3yhhTzHLM3e/bMcVc5xa
Ghl//KD6/NE+LLNWaKAzhaKWCt6uVVTXVTYjcKacpGPxGc5WxoJVrR+jssK3G39hI7KFnTzUYdlo
Rs48fSEf47IrgeqUMWDM3g500cbG2XjJarlyR9lUoDh/4RLyMXj015jAPDVStIWEYwy+XDFffmuB
OgP+117UPHGcJs2CU5VWPxFfPn/qGtYcmD/lync/Dti7nDymQpD9f7vr8ETwQfv7Y8VNQgQvzbHd
3e2lHDfaG+cU9kXOZZ68Dj7KI3pViz+j9l54QR/nmjbp/t5J2KbhcICmwWKRrT4vrC0lY9U1qIem
nToH7cId/al8fyJvuPCC5W9Z4gbKiRwECOYttY1lhmenME9An8txjZORsvZKx67s47r5ztRyyfl1
6WFGTaIZ5YW0bJlAshlUz5KaCv5NFx8mFJyFYUG9uL2C9U/JcuobGRF51zbcya1wgpzJKLLHdJ3D
wYGbxAejcItOccp6GdpnE6EJHAoOmjmUYou0QTQEoYZCLuHNq51cEBwoWu+9n3IQrWJWGJlGu317
DENOvBwmEQaSixkkT6wq7Xt9ck3glD846ykFiWPJUmmTX5cjC7EPT44ENm8CmiME/P8odR7z8cdj
hQn9bFih3HgYQ7ZfG2WTjvRouPPMsVcj5phtiWoprUyqXXOfGPR87JmcIwmMrlPis8HEq1VTfQ76
YqV3oATmOfnRRcSfYEHteRXY9N1IbMn2liVJx8L/kX+6GR3Dqac4nJW0xUeKVgECuJ8WoHI8MoFs
NTWqMMMuZ+yNW+F+YsTb5D8ij6V9qXXwBdBvEN1Lm78IJm7iCJk236EuKovuZsw8kQ44TcAxYKvv
ytB3acGAiWHad+gPb9ToQBIywdfkOtcUx3f2rT81h16lXMx5xcuFOkt2hwBvJ3Gzjd3yZGyAtSHy
NbagCbCphmBzTobg4K0cGjItWBkv7gGL9xGPjYPrXin9vgjusBj4TgXVHh0m2p8PNp9gtuXumKZF
iozcqiE4jWX2SHLUYHbFYsLKCpze/3j+vvvYPhzyayfRfCLUCNlB53SajVgU1jU3yZIel2Ms31yM
yXOLcnpyZdHVc9BmCtjqv3m0wThjVKtnGIb80gzj47+9OUyIaP1nYBp/De4hAOMrtJoEOF02U19h
I03yP6Uj8qfavHkA2C0U+HrDrRfK88v1XmjEiCeq9hL7NbI4v5AjyNW5YoX7f1EEteyf+H2LGj3o
lgPgsu0oDytL0vkeV41+dwWqnCh4+0J+/bdR1E19Cz6JNYJjoyRjPI+YdnmzITAtyl1uZ5750xuq
m4gZaM5evnXp+1vIaO/g88LN5n3hWdiJmZirOgOvJ0f8jx4By3Ta4IpMKPzrt4uCrl42ljJ1fsOT
rZwab/dB9UZxUUH6th5DxHYQ6qTb6zwOP4zi+wH6gIHy4YfiLZrNUMcewpiNZ5tRzFyEFnqMeQ8N
k2RCssjvdPgJ07A9HHCoED45t8FzIMhi03uNCgQMJSg9c26KmrLcUrgkNXFqUDGv33eqGnCZlhtB
uq+aABnI7bn+yqm6RJqCZVK8uDvsy7+aneDI2zELDGSq4jKNx4IhcgPn+vcsPU5I3WO89pfdRoad
TcF12CH99jRS3Qj7r+dmMmh4h7JPeyZq+to5pOVNquYl6azjaDls6/eBDK0xC0KRT6t9yGlYiywl
PDGb5sP2fxmaUCkVP8GwmaFiGiiu7gx1Ofe1CwmFMv12se0S1ig6+gLLfgclrHJ9lltlShnL6oo8
ukxPme16GbTYSaejuutR48Jr6uNBmzbTpjWwSAnCwj2hm9nEubWsj/g8FMfPUbq9YCAD7ys6grRR
zQz5kqDWlJ8y9BaVj2K59cdBKMvFz3IQgN7rjIs7Hcqb3iOyNof7nl9ANAVVxwHccXjKS0GT/mbw
YS23eOHNVyyaqKaHOgYm/AlOBHed62jgTEJQ5InIIReXvtsnsHjIGjmM4jhkeLcwpiCL+YW08XNc
xuOy7iTaLP3asZKDD6KQUMQVuNbuyl6M906S9Y1GX3sJwG/72UV0/VGoNmBJJU2Uirs/SuDZEood
+w/r9SXDsPov9qoGInsIpTXdwuNCAdSSBq0mPl1o1kLBh1gAVUpk7TUmipAc2h1dmvA5K7ilkoMA
TH8NoTjGOaEzA3KzGjo2DqjCwtqMC4Hq738hObtgTpuMS/v1qSejUH6SwrzSpJd4LmEe+K70uPJB
RMUSUolDDx8msyo5G7yjjMOXyYlWpEIK7syz/WUlCiwVpfedj4enJaVGoj4XYJwm2sbKxUXbxYnW
XKw4VvN6veeMFbTE90T7IJXxVGc7c8rHciIQAucwyXnSA0pbMmho2y8SW551u6MaVHottS20TBT1
7btDUqTOvvc0H1iU83oguB+XEBhhDFrHtIntkeE7dE+w8mWnY1QNPOLzO633ck2E8XYaES40E9oT
DUUHlZPmNCFBEeyKIMbptCHmK1C5rqpJDQGCahePL8DtzwMbY78yDE1z7uuXz5tA5sgBD6cDO7nY
tXis2yPZhE7MIq29sM7Zn63B1rmleJdE90JuLy2VfHI+EWk3786f391P5XRAbKMWbPpg9snKMofO
HSA68XfCdd+aeHVDjs3+aKyQj6EJhvqZnkASLPxaAx0p09D2I4y1gzbWIURS92v48Vidt6G/rzIo
BAbj/okcwOdtFmH0sk0jOJNEgmj5hHrg94CJjID+dzqm/I+nQFwKbcLt5+Di35Zx27APRTGSYx5f
WJOVkZxhxpgsYQENJ3NTaqnfRyGitQUPsbY/fNhYHMeoBFNCqQa0qd6MpGV2Kf35xs+kb6gvWqNh
6uxfL4vdy2PR6fqbUBLscwqW2NswjP8vRO3+gkwuq9Ty9krI5r8JxOX2r/PXHwo4K3Lke+bx90dV
Q6ifEIuuNsR024D8eHBpGigPHYv0T3URqQgIjgkw0B0ILZb4zSzjJYkszbx+dEDaXOb3YzLpRrHH
b9FTUAsDdoS5azvmhr5ZqCEAtOlN7pgfaw4BMXvf/DG56OFbFLLP+ywv4PZFZgv8Cl4rhcqkUqbo
5vkcOt6rtOQdm9AntYF7McC92iqwpEfsiFMgdYOdn4/FCUZeH0hzBPGxbU1cgOkX9x0ZkuVA/ibQ
JU1uUo9PBAh9uPk8+rMhLlGfBWSo3C1Q3dZpyWC2FRUT1GOtdVIFMhhsMuhXvj8Mo3r8BHN/9UlN
6dU03pKazVQOX1z4cYrkQoxZFnrLSyENiBoNYa8d2OylRZJcDPlma/qsQlfMGNkOAPaClhGvBwA9
wvf9gsjj7aHnr+cO3ea58oniVSqJtDz2f+DRtdsulvn5ik/VE3qTAOUi9o+/G8z6cTczOAN8VNRE
Oz4p2ZUYOlwaq5tCpwOhyai4l2WY78e/QrTlrrhxynX9+S120zaWRYn9fBpJv5G1ZoCVYBnj+ItX
jGqmSFFEiCA1sLvTT3UJL1VsSinNgDMNMHXWgi1F2SDt7a2oblwM/hwy0D/j+OQ5XuXIDvnlUdrg
wn5wY9cyBzlQ8ymSWXLOqqQqbtjeoCJTLIfM2MNAQfoF42Ltmsij5QKsiCYe867xQhkKKiYcBVig
LoHGp0GNozYqP5+awgv841+Th6O/hOfN22drJey2AZREVHzC+VhKwQij6eMF9OH/rd9y4U7SeF1E
iYZYDyII8j4L+f6EpjcnGR7mYCf86WZkJv1SxlYGD2ASPZFxT3Clu34Snzu2XZLIG0nhW9rpIXyI
F6eBuElpXvSLgkweSQZD49Ee9Eg7bZgFKiXvcxjcYFIDLtt5jH9+98tcSy+B8X/cXR/rt8xjg94d
tfkLXOTlaBlL2n1VHkrtCGjriCvBofUj+Y9H9iDk5vIiryYmi47qt7b4qFfHqKktD4lHee60x3iv
2NtkQ2djSBHJGvHGl0CD+nklb7sNQlIfexPr4/BXqQAYTfj3vCHasZ8jvMTuTINo+r5N+HlyB+dO
56/BkW3ihxw9uo4FHW82seGdfL2XMCFUOpO5XX7KQ06GhuaFQbc+5Uz/nxjzgmmIX9n61qYSQDkZ
ouowrqxlIIIMDvCN0f4FdijPU4ro15Hk/1vhV1BoRQIoWet5a+7pmZz6tPcgDIX2hUR0L3GJbnST
c+Mt9spPSoGqHL6ZjrbQmC+gJLUzTG9FemFXof34EndO1Iye942Hz/QTZ15OE2+gkwt6iB6yMWje
5tgoYC2WVGe7k2zy3UV3rT1tuXsLNMi083DUOKzxCeGSyk56ND74U82KEpO7nAg6Xw2au1hVuFry
kf0CisJq7xRlMb/ka0QXuFw6gVjL4M7P/u+5y88hujt3pAuKUMLpfUmY1898TSL/hsK1A9SUz4TK
WB/7EIisQRuCiw+A6kh9WgE2SVWQU9Mz8S8O5pG6VXMELJntv5xvEbVDQD1eFKIKLwjSDxD5rjKi
rYh9SyNJ+80HHmuGef5KHPwiSEzrNTmRNF1IPMd2VppTxAeyGTUvkh38feUbfsZuJLGwDjMskltI
Svq446cYO3WN0Sv2B0QSNhWuXLBTG0Gq4QhTfc1zUAwhuG24/ik2kfKcbRRQ3uYvIk3KciGHAxhn
+nao5h99foLv79uj3/HuQvrUz6W7iCbCUTtUj/rQGhOG+AH3sWpIlxNdrZrWE8uVAJaTruWxGqmy
O941lb8q0nJSwdEKRTcn6ymWdUIaTMvizLjp7a9VgqEqEX6KQyqAOA29L4G0CQnN7dHKiYe2m8JY
2fhIAu/OGq+nfFRYBiuiJT4h7JJ60utsplfM6NFo2R58Nlnn7VJBFMe58bdaQAMce2e/jXgfJ21C
h+F4KqpaXY6k9RdcoFiN4ZrH5LpaQkKSR5QvAEMrb44wMxVb7/bXl4BvfiGGK3T1ndL94imVh1P0
t2g5rVuoMp/RSDv7irD2HbdGwLiQ5vp7OnnymBlGGiJnn34FVzANZsb6mlg2Zr20oGEpaB+sD++y
czGFpeckWFCRtAg6ODVKINNowW1pTnOun4XEJ5f3GRG/tiONZdkUGkgdH902JjrQbmNiWur2g2xM
4tNxOQBJ/b10k9wVcpy6n4h8C0JMRdbChLV7szEclynupVPJp5atsIK1VHqT3nCRjDR15QCFPioP
Ntd2z/FAkP4+GF4hY8HPcQmR5RmPdwWkAbFiOf2+RaG5JE2IrmpJNLCWsDNk5Nm3xvjI0fRHlQqL
XMrfawRsPbZUVpGVjh2BXyam7IPIS6MI0NFotWrSfkVv344twbVUsEexGt+p8hPu32xArIqW73u/
1Be18rq5jgW/Xx8d8A+1YbpnF3GDQeUPitZR8wPiy4DXwOqUOOZr5RWyAiaOJOjXTv3DoMnvQc5x
0wFebUhVAzdxb5W4LjMB7EhRgulQNyAq2gr8y/qBbz2Cf+NOrYaFRpdzlHrVlhQJDbrZgqngF1NS
mC/p1KGJ26heBDDOg4TWQIfXtDkCYrfpDNRhoorlFaNrxi7hfpkyY9Xe8+k3VXgcJuUtB9Y/mAzD
9FyuXsDznVIFN1csZ0nTMXXok7km6/kdFqc7T1Rai+YfvUDcfGvrUkqepbNAiucEN5EPoAfLTOma
MM/gI/o5tlwq8JAU4m49tST018LoRbHDwWMkk1cCowovDfjq9SM4ebrgEkk8dRn0MSq+qT0U3GL1
x1cACyW8RKWcDXapOPPMU2R2+UBau0qQtRBNqlJy4eCphAruLiMNlRbOF0gsr/N1sJRVphl6ri3q
9oEU8RevA+UZHA8kLiiv3Gn+AwzVJXeXfkg2CAx2IoYZGzQMygycB5UCjcYl8GhvAO6trbZh9DVZ
fBfZMYKIdn30pfUkdwoywO+k879VjGsQwuVjNBoNuMcMqRAR7/I/xeEY2GHb8cSaDEbYDdcGkHp5
7YAr4JrreOZo/qTKdqNmfksD37G0HYJbIiIHwkcBbEmwD5itPl5AsUaW+ZIFbttlUAoMM7mW48s0
ukbbzxcknb37G9YhSKtp3+UYmRtNBb5Uaxixk+EV8Wj3ebEwKwdXcCHaK+5QtNG9KStwoEGFdzyU
VmKTDrgyenhFNPOVRZY4HKGJXDD/Y/ngo7egbQPNn7apTjXkepYrd8yeQlGiHmTiGNNgh7mhsVt6
s33/DCNEWE0EZNUly4gdHP//2ajVt7KWBftlUDXeypG+b/yJCdHwvDyq3sb971po0uwo5o24UOqZ
vUuVZo1qXbttmIdDpLHyrFFSN3dH2z48iQfCR0HZukMWrl+dAXLZbYN2BXkWJMzbHECA3Tilc28T
CIAyqBuW35zOcuoScX10aDHO88mykRnDPhHTlrUf7AxdGf8Y7jW8XmhbCKJ4mbqbnGOMbHfcr9p6
TPc/nEZyA8WBLPh5w1AuhaYGymFhL3nZkpxhV7Hf9wP4ZQNaJYFbboj/9nG0Jr/HloLWrQ2Xc+rS
VuJvqJePk+v3VHNV7axr+z2FbqsW0DN3Am/AoBxfH3pOgy4gVIbAu4Ezb2MClMxZp46+71sG/AmY
rrmRv/O10THWjW8IMrmrzeELBOFaytMv6h14jsU9FRLAN+RaxFHkoQUSy5MMDt0+Kx3xBmDVRo9U
MrpZsysKDlO1na/+N7ZtZ827tAXat5onPnRAfns3TdjMIEP8GLAGxV/q2CaBL+EMTqGQ87hDEqIT
OISIIOeyfMnFw56MPFknUZauUj2hQsOQyiBOiYPpUzMJv7TmMbuKBC+gMjr/Dq4JI6+dHntKWwke
//OWJZn44Ce/OVfWn45DiqmMd0bKYyq/Kxb+aQfsbtaRxM1m9IUAO1vF6Yf9Sq0em8pU33dEERbX
pPMXY5PximKYtPVxWFkUaU1pAJKqCd1lLVXOhIv7A9WnYICD9ccm42t46GYxe0DM5pxRk93lQO4X
vW0MPpCSIGRDXLPvexsYczreX3wvzIfShSRukieAK2nY+4ygFP+oRbvlxvA/T3ukHxDlYN7+fuy1
5vSOPrTomaWkkICVK6mqWTZqSoi6QVXcDxcPyYNPR2KLf4Wq5AVoWzIPVi1v0n2uWSqk6HcJ+hK3
/047dsvT7EQQwQXRP7+INZ1j52ozAd8WkTheXHRGmbCPAuY29fwi2KdiMtQG1VcZMKmZf13Ns8kQ
wAMyN0hIdz0FDS/rwPYmfU2+tLiX1COp70WSzTpxUsOC5X0XfZYNwDbaJdehbJE9TJjCMfsLe83r
+5iKF4cqDa1vpAp72N7C2+dj/lBkp40WSU0sbMCmyunh0Trm3sG+GBkdU2afL0mNK8/96vyOHIih
Ryu1UUbEcqR6Z4H7ns6P+YsaXEFYnrSYjvVA+7mA7Dy89ERFTLXIN8TelQWtK4lhOoP/Mdt1brD8
SBO6q1PvoDS1SHk8G7fkuBjr3Vw3AnqHFdyYKWFzi5zCoNz/qV5YqX4bYGK2Ad1X/+cyfwzqJLVi
kyPWaV04TIJYezvxGFc1Lq/Ue5ObTde3cbBbci1ZnTf6SHYP/HF2J/tk5CEYUvHaC8hwCXfNPa0b
4j45YPTD+lUEqma1Q9JH3hQ7/5wsG6nygvpsJpcBYytscjwGd3LXpW3Dqj4aw33yg14Lee24Vt15
Q+UGF1PGavV5CDC2tf/7UFFI43lRk0prnfkdE6TWamm+4jHYD4d3Zz+tO9I/2j7gZuBLUmFhcT/R
5oRrIOjdHbRo5wrWXWUG31U8elObSDXVBp0Rk4Xk8Kw6Yuwm8yldwnmVKm3uK41JrzLUBZCzUCHR
bCfj1V08JrRGEIwo0uvD6u9xgJzpcGlg2PkuKv3nF9e56zelK+1BINuljlIFK/bKiWoipghyn2a2
CuuGrKT4E8c0wR6fRSoaQNO03dkfHo4/IdVZyYI9E8aZbvO2aEQYVaoVe6QL3+4hoO5rpj0RuK/m
Iqw5ywFOqMjNm80uZWx5xwsqJDmsmHCMuUcWQySx+7SESHy10zmBMJ5vX2uexCDzSzdro6MTGxZR
8w94T2cM1BNPA2paDFJVCj3nl+ikqyBFkuL5xoG8uqhH/lKBRr4OUwTxKRSOUIu6bcMPS487UbYJ
jM8+zvYtIfYdxM2vVCzkqNAk5Ml4EYpbWwcf49i1T/ykQADnMWRR5YOGdXjMYSe57lod6ETWu1B8
3Epg5kujnQFS5UY1R7u4SlLNcNap/FTeZoJseGt/U8s9/KiTRHldT4D43m3KRqes+jXijd5qFLYd
F8VvUohmI9XN9xrXGUJcv7ob4tnQrP6KwGJTkkbUH2UxVlqG2oQ39pbfXsbPWBfC3NDs1i5dHxZD
D5BiJe9rbjvCNUfKJUzcUTLcvYvmG0h00DmTQyPmiadDhepv2zIfmO0/M4THTWqGm837KIJ79uTX
2DIdRTSF32hcisxODKbhcYEXGu4JpsnlgK3moQwbekqEi9UuwV20qwKde1Gdnc6W8ZW+AGg5Dgb9
K8B2oKKW5rVtL8d4NQWgcxsC1v2G8swbpnbzIm0CTEwt+Hc2IuLJKTXSmlAaEzTmNp22Kqnnstky
tClIxembiMfIP6cbioTxVDxqCl3rAb5S8m5X9uIizoEJubLidc/tJoCj7gJmTO91SiTKivbc81yX
gIOWjAUODyOsmmzW6JeFIn7JQgSfgIt6WyJzyl/o69yE/oxZdqZ0E9WwlRqvdoEFt21HZdrbHYLr
sd23vHfCC1lAap8v/Br8b7dEs+rd2IJYXyI4l3bhSSkhpPVuqPvXnikjd+iGchWeEW4ORMu3cB3+
D7nl++6QqGPstwBm5dZnXoq0fmU4ElUUiZeQnwnud+fa+34Q3ZW+hVZ6cWifHcaEgQv2NJureQpr
gU0r355oGO8LCMZEVv+tzay6lWBLffE8wZAwqSjtb/M6F33RLSOZTFXnykC/k33ThJmjxrqMybNJ
JBXnoewckItngEdiq4YlMBMCcPxv1/biT/W7BCScgjpban+iUE0YjY7+5PNRr29SFAP5TiEyc0PS
TDrbrJx1co4SG2SX6BMo31izWL9sL+dbRcPR0Jbjo9Ad2wFxzKuJ7QHWG81xNrF1acFxPudwqqKw
TmIZEYqah5xK/kiRKp1vDUNuXJjI/pMQteOgwzts+8CXQpLKdw55mmMc8T5DsPJ+c6SxR8PFycGC
l8a2TWO1n894RNkaZZnqasZFgp9+5GVcjrSyVzLc10xYh/Gs0oL+vplWSsJqWHi1DRkszuLhzrX+
vDkfPJtbydTVuM4wXtLs4EbMiODCKF6bXASkcYwAZLwgjuuAfpG/LTZPd7nhuZommzC7NPBq+y+h
cLpjdTkDLREswnzk2rYm/txv4j9EjzkRF8JnSOyKTa3RV6qw3R/lOMmwwCybAknN3A1equE/T3Eh
6Z3RSAevxaQoGgrjjYGIFQ74G7ft7GplUd8SizoQZHE1gan++BZOaoWrLbAnOErN79RVD7LZuMdH
XNDFCiMqvwAmyEMJn3inX9jTm3xYSTApiTl7ncBL0Qq/qim3G2Tis7AWB8f+27RbuBHYvSxfU2eA
yByRLh9HXzHhsmHyGRO2dXrafCrlX34jRuBIqvnaDgFQGmjn/FjYvgVxU1q5EismQSUnDvp7tiXK
LLW+PidbObIJozgYZzkzre2LoWZhbPCl9OMK51ZKqJJsFvlLHQFFuliBJmmxTc8h4rl5/B8wXYZa
y5Yo5NwwcKTOqb6N5GpDLe3RCvDDabnyi9DOA8EAL1CERRR14UBOn9ges7fIYe+6D2s/aDfERRey
WNPRaa+2t3Td6KB4GEGwwcrVjdC8bcocLoMBu73JMHhzhYXHP+KbH2Fx+3SyZ7ujLuzk6L51P08U
xcvGKH7vm0Di1ji3hnFKMin5aftRuvmxXijfJeS6ByKMlALPbFNKdrEtnco7IQX7RyM2jVuPYmjm
ZXLHfS1u6MPRYD0J9kPf96cz0wVoXbwV4Uxt4SXOZE0SLyYI0gQVVev9BZO6r5j/+i4z1cVpdwVb
awBvlvi4fHKhXv3b+CRi/Vt373HafueS+2f06/kldbHP8DlHQaRKG7BbEb48j+PiwJbBHJn5fM7L
4zdvWGkiA5DW1yOBhnfLmCFTiyi10wlJwKik4EIuQg4IWti13WmO9axoBGiu6vnAyrlNuDDcJo7/
UrC2W1C+WE7bHfayTlBDv0UvQpll/8vCYPrqDabsVSzaEtaM3EScFwUahj1rmbiPkPoOU2j/QdWC
rct2K6TmKarSBl812SdyQAZtvSi6NMOolSRK+KHl8IN6umoti/btZaMo7duwYKwUrj6YMppcGAtn
kzKhRELH3PW9GZWvAoZAniXM1eOlu1P4WJLCUKqlOyHcDZDv8A1iZvBA6iurpOJ2WjtjfaRy5ASI
+gFMqDNv+ttFHrv4YUPNkBsOyRXLr05N1C1hDFWj8wKgk0z9A9rOktvmCjw/wb2KR6uuNHermKFJ
6ngwoSIBCnbllelr5wlQwztKe5n+H1/sqXu2PA+9L599nf9RHCvLzrBORth/LC0Pq+78tc8L6DTD
AqBv2Qx0ihbDHzarQJ7rZ4zSSfQLHxxGUxZ8FRMLMapSb2Wwgb+aLFGCs46DOfU6fu5NRWRtzS7f
wxI1qy7XhXwMZailu9JMdh8d6fVSy7KCEzkHf1BEsLwE9RU65PCS0H3Hxlz9Rar0c8Q5QS2K1Nno
pfBC64jppjjr2XKLEP9L7fWYBK/gp2o7tdUum9S2XFFymEQIQyZxCkErx5GBmm8wWEl43nZd4Kkc
+B0JSj2kfkJL1BtnsSM84AIoGhwuCNxUnyWynK0fYGtIEYn6/63fLe8lvJ07nGlKNN48FOcQfQA6
C+ZY5jog9jhp5bWKFcEj8CThUmg/nj7/w2X74KcOpgK53G52RQPDQQUmwj13cQkvAu42UBthjvjn
ySXKDwUM/Zg7/TnK/RDjOA8kcQdIta2E0wGK57BERqjKL49mCQD1Ce/QjxsZxaAJKa8RAQPwwmhf
wj25rbJWKOgCQgGoUE00UL0ibbQpV3b8TMRfjb7gO8DqZaXasvbtawXZ3RfZgL0Dszf/oXlQtvuZ
Gq507LIQNPhY1hxjd/4OBqhxcHQ1y6RCqhBfO5r4K4Vk+9RwaeAsaBI3f1/QIv6qjaRp3+/S0Mhd
uN5lUw/8QiSJwLTOf2osTh67Y1WJ8V8B+92s3CeH6I8jKes8hPoFQAMgJP8aaPIvq6gakq5y64S6
8MjLIgdQlDGotezld5fcY1JzrIyNRUakyk5cMaESUcAmIh6xAy26eb3g0zhU6d8Zb1YO7cmyhln5
hm4u7Iuvw7QWDhCHtHQwV3E89WiHrZnFfPGpjokawBqzUfotaF7tv5YcqhRaA8bweLWVRHAjddgv
eBteg9x8hEqjD6r/bM0AyUJB4qFIT0DvwAiwdokzfATbbsCvWyWQ1a3uUSyQTkrPydKFI3b03JB+
L7mSsKimWJsZGEPU+Tip46C7A/WPw/hU99T8BB9WFp6bd7weX+lPwYQQMAtEd8Xwk4ZfUyPnLZNu
OQBjILacqB+YDUP4r0CC3cNYz5Q4xH5k6TGHfY+bU5y+3HgFV31WeXaff0UUo+nmaGnDfyUMh/lQ
xprzhy9PZub+7wbBPzYh1WgbDgf57UwCViU/C3EuQdrAeUomhq4+2KbAg/yzwQHjB76fhXaIwBsf
kINB+ZjMPpzcJShD34gOnfDZiKoU3hNlKB975Q56pDfPGDiF7zBmZd3fhWpPTQaVtESrwjUvMisu
N3sNNoyMtZgCqE55B9TWVEtViN1Mr2OWzGz4itbOjSTBpCzLAk+SDc3aic6i+dH0h35ZbOJvCKqf
qGsDXjs0kgfve+jt9P+s5Ggk+RjaG6IbDYVm5Wx51jBZ1X80xDcLWkZUyfONYkcX5jTXWtWDh9C0
zd1B4He7qpug36bkFI/MUtwVc/68zAascSJ0oDaP1VDLjkuUM0vZQWrpcvONDOloEFfVMHbWsWTe
lF5oms5ens5XRhqmEmgbUdx1/4y+vw3PN8sQWUOSFLzYwhGNHYRX+QgsN/4mAAPzeuTrNjkms/8L
TNs4VUiziUAOdicchQP11skamsm8kz4bgHNAV1fDeFF9B359N+1Os76lRwYgNuJB//smOqqv8BD/
SQihtAH3kNBycOlsGfnmyF6FXKOl59wgdv0XrAehidZ4IaHHuO9GObfa6+1EnX22vvcJn29M1mwH
VDrgIy2c+++0oqNrRQUG4q+40bym0bU0/0EIUXQpP/UyW6Z0rhjGk5ztnuz2XMYig6X8yEZTf9wP
bS5ljw6EkMza7GG/2OfHt5jK5HHp8ZpFAEjMlZ3+VuU3T4XrQfNXVTtw5G7YGRV9p29fTugV7MJe
qV7x6js/scTHvLsrv/8INwpbSzJp1F1Spre0NVRk1PiR8F68D4G5dLoyrmeDqGc7R1q+QFABPUmU
dfJKPWxQ9q+FNFQwWrUIovIBqr15eeIeHL01YiRqmFWCooaaPcM8oEJvDyUrTGf+m3/jbMB6fWFE
trCGF/5mhA48zbmG4GJHixiPMzFc3fGAKZyadc71vGnecvdtOubohoMxkXiCKUCOGCst/RtE3hhU
5fyO89FXkGBFwERPGYPaUz2GHoxohUZ6m8JkfIlHm91iCwAsjkzu/ADa0AAGjkLp+A4WR9fpRQtk
4g8p3m0s+rbJXEdWAbEPvL1MsLD3YP4G8zbL/srJTfrQwP7mvS0eT8jDpca0VWN4EA9Ph8yQ4JsF
/SZg3JpoWi3CHYqRXqRP3/LFKcnypqKLLpOug2iaipPL3adpgOFIiCMl+dISMLNdescdSWqEhiCX
KESErcvAptckUBvwCejp6UllMV6/sEqN8XaOMsx7U3UfXnPSFPjWaTWlaCkqyRukaGZOZ02KLitT
6Zs4or/1Yljm2bL3y1ttwSA0ULS/oJb2ffdU2pEa0a+VVJv+OWRxN589TvRzEOgXKqKWTyqat0IV
axOpfEGd327/KQESiREHe7j7zgBdfOcPCy4x2xT1Kzpt65zsHURjEILe/J3FVHyERwcqQ22b9fwp
eSMZAM3kyRZR+bwszsc1mbFIQTIwf2PWcp31pO72FXJwjD5P0oq7zcn5jrwDiZA0O4cfHGbuFUJH
bejXKzjdcShhu5NOldZGZp03XMaH+Hw1j1aIsvbBn0h5cyEwqp3bmt7VdNtDhbXU53tskinUWElQ
/7OcFez0PR+xnV/D/D1zbcb+ES/0Hgx3R5Eov1fGwIMu/8I3Y9UXWBdUShAU876+drJbdSV9KkEp
sXM0VjL2qEPGe+A3pMh71qGZaAHcGMNBlLFysqisjB13n/U5HdIkZoHd66nbSyOWEpiNgwrFD5vI
/udUjtPP/Q3FRRCiDFgWgno16MbMqi8cnGb90rgAyqTD5aNi3T6HKvVOf/YaKCPnjLGihaOT/sdj
IO+QSkcog4dif5xWh3ZMLD+vF3YBrG/r+n2J/gMQQ8pP2G5c8Sn78RHk4E1VzdCN0ff0v89TgV8f
fQnh9lJix63DoK28gSkaqxY85ow/uYclPhLhpwH7NkucqXvbxmU5p9nGKRCm+3OYH3otDViHp3HF
SIFdPgdMP8SIRAZN/5aBUSWYrRg+mp/8qcI57sb+0WQk6I5RNuG2xq/Vi5QkAbhNVTeRO8Fd9mao
jqT7d0dQkaE8r6Qh2i4pTXERNbBUmenpICrjaXKRsSqJpjNea3f3HiRHAi7W0ggqKY1VPzcfKN0E
LOk7NUSX4qzmniM7LrqhH/7qTb6VdIj0zn6VNJT9qydysArDGoPFfWO1ZPNy69WpSAp6KKU9xFwU
Mn6HY0Jk9Aq+2KbP6s/stJOw1DU1Y+yOvpvGxMOYdXMbhgvCyMBaws9fOtYsKG22B2/Mb7ikkWg3
qAwgpXJ9bkIU7ggRX83QT1zmQ00orSmJ4bm/vCcg16G3ZudiTvRJXgw5LywTbOWbU+FsdPQkh+kE
90VcEZyd3qLOhAvUqrvZQuQ1khCqycnw4ZWbdmmXmDqH4OBt3joCdcuacnf2tOvRKjIcPRrPUhFZ
mc0Mj/pxvgH5blZmpCs7t6OIlIjxx/W0hZL1G19WGc6xJtBWjA3QCCFGS/r42GAdfShIvCgFGvf+
cK0C5KLzgdw46fcXBdmIaiyW/KEzFiDHvs5L1K9QPVnZGf/ntyqyFvOAF/iU0YMucLa5mJL5xCtx
hh+TNPX06xNLgtpSPLrQU0G2ab+DZz/3k5YJ0Y+SNc6ANOWTT9DpsHSuP6PIlmiJS3FIfO0SaI9o
tu50cHYcr5Dw39M7L1WwZ0ezyucibkbdayj77KfD0iQenKGFia5EOg+f3p4S0rL0g3a1eYdWYdjP
3OZh5wS6wI/jn3TgXWeJp4v9JQRtVj0Crg21qHG+c+H83BPbkW/9m3kNvg/Ewdf13K2gZqW+lAqv
PB5Y/x3OoNMHxmL+Txfxd9JepvSk6XMw6VSQ2wLrJHfPWslnVCsViVO5cT1ZZnLwyl345CrYqYnO
SbEc4NVxN/5StiBcOl4nKchU9liQW8NrNcC7ld5hGl5F+Tb+FNRzzJJmKboBXDaMeRqNH3IYMi0H
CNElRR6N8wEkq9NfrgNewD7WOc7tm2R0KZ4hwF8X3gW7Zi/XCmlyb6fKwykhN7itEQwxlbGSnwxf
wNriQB7tmKqwnJznaEOrrzSIk5R94nlQMO1PW+e+NkgarZWpRmXK8j3i2PWQSHNbCY4uW9NELaaq
hGHUg65AFExwOTCp3EmLSTpCkettbCHLVEYETMw0cbrDUHebSAz70rOlHwLEwth5+Y5dbkrDBKgO
XUddRX+ugfwjnbMk7LiSXuJefxmJqjBUdSCOpc6qAMk7WlfDLgjtI0BayFQ/JlTCElMsq/xYIfzd
14UHqBddIWZ4kUr7S4RR9Rt+HRKXjMrA9M9slAmBj9Dwc9OfcCRBi268lK+yH7VMvHElGMRwvB3u
c70qQ0N6pL+idJTKXyof5ronBwAj4LtbRFhB6O7bRTwfwSChAlmjWmRXyhyH145OrLzKcsc7woKC
mKVVdXy2Cf+/4kHkEUay4NSlkS4L1W8fHd6Pbavd6DmmPZ3WKWjyQF4W1TwMOvV5Y9lnbqZqREXz
+KU6JmNEEhdJlPIjSgHlQJCXsHA3TzQCAF+X3e3WrDs4ESn6zwmqPiT1MaJWty9oIv52LaIoxcst
V2ISajzZS19I6Pn+hoZgGwvuEicxv9XM06RK2N89dnE/ucIychZR+6RektlC3m9tIEQkVEfQgyUB
TZWZ5FNSHZQU0fZGDLEm1k5P3MmY4uBMRBtmTrb+jEKAmwtAr3EZlGaWh4NjpHTpOIgJNgajD0EO
kUw08SofnMyoDDxIjiwisRbdta7wOo8CDdkTzd4zmhoQ2AOuyU0oV7wCBZZnhnrojf6zDkg3MFaK
9dzr45JUpkW2097W7Rdczhe5ZifJTS8pGRdJy7r82c7AsMQOmFJqhIAIY0qXbrau9dlQIERutPsO
ILDJfo/6uEgV+A3m8g6cyUVi8MwdTk1swi8W1dr0iODsyyUyveWNbCuDokOpq8YZDURiPPNMHOuC
y58vKGQ3YZK9sJPlEFu3NHhV1w2+uhmqu49NOiJAgOzPQ7pNfGklZiZZyZXOvB9M5LQ/3x/9laur
Zs78iqfH9u/GXTFQLaYL1EBts2h+0Ufaqu3Z0QUU3eT4f31lSKLmQNb69qNUALZLQa1re/E7M+om
Sh9y/oDz2XbsrB83VUJi26TbwS09DsoMcWYmuAZdmdREQTmlgWZgWNQrXdNqgeNvu+e1Uq/Joj/C
pW0cBobHCYeHnxtLqoBb2xYGiHai0vOiokTF6coOftO7Qrb4nEtXTAqu6ssEfZfkwUJe08pYTVXe
6aT3CQe7jzGqbqimTN3odjKEEx1RBnOUPo628sEkl8407yWF0tRKBjZSTlO9lGbPNzKTsssVVWKN
wtSrHEARt5dJYZpZ2Hsg+3K/FCiWcvqkr8hA01V7m7mu8tUY2v80Eff5tur6mLjy697YzKcj7Gh9
IUjzOllWJFkhFfJMx8iyJK3rwGBh2y0YX77bgkVJzm7p36KFg0tf11jBU2A+9Jpzt6NMv+Axx96E
uLNds2jVIVqbm03+LVSMD94PDB8YaHjP5sPneXTSk18QOUshgOV0fLcQqopJ9D5K5/3ZJO7tT6xi
gpxpnnT/5/a2jargN0Hcjufryg+0bey2tjxD/rPB3XYrQo9xzxFzT2bHSjO3ZGoqSQOhmYUXSFa2
qdDvgN7+QuiIIt6Eoki5QKZZXdDS+LmvRyK1o1EvJIfcN9F1wy91t8Rvl7yX2Dunq3zaJYf+8cMj
ql31BVvePP5yjTdlBeD4yix4q0c4H9IfV6sVHhByv66ocN0jSLaOfBwCp3xilCIix+YbdRugUlbI
Z2MUfldg5HwK02aLvlKFEOxsTZPANQhjccm6oOt9+6Uv5xYi1/SjKV0gm0Fx7shChSsaDeX2FYLu
fS8vXNhIQ3JlxvqLq95Kelke64g+gRHO5AWN1uYGAaJMIdmb06cHLFHxvVBokuZoFxaL/L60jCgK
0jHtl57QZeqB2NXU1WVNBg4GEaVVhAQeCYJsrT2Vtye0VPSO4aZiwrTpDM7gKL2oaBnS4det8ib+
DO8uCeHLG21oVLufU9bHFaHr583fJfQva/pXs7E88nt3mZukUN6V8pveYZycKZVPx0kEFFB2By8Z
ltozSBEWtlVKU6PPicxFuuCtMtbHwNG5B3aWFnihp76/vTFz9379FAJBJy+UTrkVwWNNva+hyK3B
eqcwA09njgX6FA8L8mob0oIoJrFPffhuBgKVlTfciicErfoaOgZTZYdBfCSF7UkF5fyK0dK7vWF/
uPDP3FvvGAHDf3+aeJFl1NzXxRGpzgVuAaWYbLXkLAgXI4rHbAEk1uHEkt8jSHbQiuEPmzwPnZeI
jmUYpu9iwtDAzYVsupuqe0i7segygi63iYBm9N5hrGrs5Lek0c5nsCks9piGCC4MkR36A2CUKAeb
fpVd1j3pBiSupXNm0kYf3R2QZN+9YaHSAVaWoZa4h6N1JYmknmgXGRHkk0rByByRknFlncSIpKx/
hT/jU6VSmtBuWgo3t6OjoIxHkU+uCiS4iRBik0C/ISYb1wlB64JEMxUTQFCAJBMmfjE7Ll3po96C
mQDxnhG3aVk9qRYSNuPPDlDK569kU1sRfsX0Gw7OAX74bhNoj0mopu398oSqYVIlgr75CsoFq9Du
SS6tLWUh9mfg02y5fyMfsHPXjapcmvGCOKSehdcZQzKGzsez1J11VjlFn1puAsr2LudJwMuC4mOy
bvyb5wSuCvO360bIpRe4mAjhbGpC6swDUwvAefR0NTIuoTnLgzy8BHkIIq76Xvn5v69oJOca3Yap
bGTqOFLeFZ7thRv73m8oofYXDJX7NUMpbB2R46SWGYaMxWFpvb6btz6q5QZ7FP+94ii+iF2X5Tj2
dadLHuk7bu4lTOor3HG4EdlHnCmwjx+1wsnQxpr/gSDw6Hly7aEOT8VjQRfSGmK3N9WZxRWHknGU
10yQF9CUi/eJka0O74/WdQM2M2CRjS44GojnpGmtXXOPSr3k1yy/JNcpovs1FtJs5B8n3TfMbbeO
isrpNjlYjYCWCB75b6tROm+aCPNJ03ucINzLCDe4AjlgcypYzLUnRpv2xlMEE+mAJdSxxUCc55LN
v9jUzM6AP9cXWYdVC85OfoiBvzqNI0EXulUhYH7YRrjLGhg7xnZnyGDujOeHA1oLgceQufX7rCgp
U/+7z6z1D18tJB/mVWj53PoIJOZxh28cN/UZQeMDMT97C642WH5UTFRzxmmud7r242JCvUjOOEUF
MdHzUtKuqewiBsMIT1N4k07kuvQGirpUOtOI0NF6/vyMinDl0CeNRAnJZxFfl4h84w40PkowEZyL
urDVxED7UpoFUJQxDJ8/qw4/abDuIFiiHV60pGQxejV9vMDFFScbZ/Bq/sQGCqF5dIIY4y4xCVZH
iiw0CFx5djCslFf9b5zVjktdqlPioRYQDUN31xYimLU8Z367ha1WMeutowlL/47lznslsTUBikBp
Ede05WiEp8VagmdvpR3s1kE2hUlmIczLBj9e5LZXIHahcfSHOd5kMD6soM4anaZgGcrMxyENvNcE
kBYGd/iprIm8RkenckA1RnEILyRtQdFTZG7QC9IDQijrbLpzG10Aiq/IGcVqjBxrbEucV5iQ9Nxg
CwTZQckVN3TAjzuM/ATKzEGdrGpXiVtkHZti3NUu4F/TKQ+9f9v5w80dPxN2hNsKbJBXYC5M4Bg5
AuwsblM7pBj5ciDYoN9OSsY3qH7EI5AiPzWG74nycHMFo7Yojwof9RtoIkLGGGZmn9DXKjkH8IIh
3lltwVI9qdlVRD06JLP/SMhzdrQ2yvu4gcZWFrYxuWRqS4dFY9Cxdr5jEnZNTAMqwFJith0uS7hN
zOhHSyE3WIxPwGoWTd+STum2ea5LufbfYYvwoWmUOys/bwMYhN4Qk+eBkHvuMMT3BlEs5ikJwu7y
OHU1SblqSfVMJ6uv+3wjUehvFYM5eMc58jUKO2lb0Pg4OYGP17FnTAJuNac6p1iLMSGcVRpKWUUa
mE2vZhZDVhWwxk/wss0srjk/SSmBEyihF0bjvuF92xApF0jP0nLPPo1ogiUKeNpsRdHFP31ZNMTr
ZEYBkjtdkLEfG44CPYeiKV9EmrvTSq4Mo0b6dxZVW2/M8f3oJN84QzSFg03OGD2HH8IDGoazDWHG
5FU6gn+1zQjaDqPasIvSy4ltx/ep33X1uU3FJUmwCK1WqrkH/yXOYquLPS4SOInrUxRSIGPfzm7S
Yx2y8SxLkPyLhiGgXO6E29d2SWkEAgLjumwROWcw0yhm40Mf9Kb8AAC1uOln2WWy46YJTfJZ5PnX
8NtYytcxpS9B/CXNH9nOKxZrXXik/y82cEVTm0k19IWHOP+nSFESDFaYydPVoVdCeV+xN7Z5nGxv
V7Q3MHXSUu+kf8aOGW9se1fSzzf2CMOPYG2HIh9eFBB0uaRYIfLG8YCnAyYSLhGLTuZTCZbxJUvE
V974ME3h8L9RAhtym8BlzaZDcf35ydmS11CWnv7AGbl5tsTitMhLTLrISajy9/6ahHmPr7ru4xEN
5lOoOZhW9Cwg1rE5HYHTi7RlYrYWNoUDP5k+1uyyHgJjg6EDxB5tUIZYB50n7xnbdlyhmPPd0/SK
AV9QvV60N9vxeH44NWCyP0dFrpdAyrUj3aCLIiMQ9EXlnMeCfhmY9oB7z0sw1QzsoDO7W3cDkTa9
l3dugRCZ4eKd2wIaarlsSErLw5YQWf4vH+VEGTlfpfFI2WBnR5LoIOe2RrnEHK97swQXXMKeIMq+
SbD4ZHsS7CN/ctjQI2Er4N3Z1m7huEGktIygv8A/4e8brtH3+useYSJibgCJruJ5btQfVnP3lHkG
eWV/MI1B/IkYcje3zsEtweApRmPzgewgOnmErYqntYJOPnLQdBiSSuNXw9Pp27Tk0HtbxfDIMbn6
4962qrsXz+xGdvG1L0Huir5RwyiisGzJ3JJ+Ftf+swgEy9dv5DZL+10PErYTZq3yPW7xv0pMBhzI
iSghTMaRpr6ssDIsIOom7DgF/NY294uUu35MLglSCbr1eeqo89zeeXxeBoTH65NDfw0Zw0/esU3t
hkS4DnC/QKQVSx3kUDA4RzsvZKcLF7u/neuPtn7XySiFP0dAmt6In1fCDSsdL7apHCuo8McZFUHE
k/1Rx47/8PlyCL8LsmHXOGg8Rr13itlWs78Bf4GKjLlIh9ZXceeVipDAd8A/IWWLp4+fM/A4cTuE
R9pcfkBSAHVqVUmsTbQBM86L+p0MrPbLGqoucAveTwi8KY48+rSvOeFU22srpcTOwgKyRvcpkxGW
2DRx51KUEh2Z70gmS6kv7kkFWrgrGK2Duc89/an7mKYty85q5gNSOd1y7gcJO1DPGOv8D2CYcyee
4qpVRs+v0nHip8Y90KrITBg0z7+3/btpkU4w0JFU+CA5UkQEEHObu0tjPc/7x/GN25uhNfgpQLoS
EJ02CB4CAtJ4CeLFIQluJryfG+4trtYJHo8IBrUcb6LoNSbKnIrBg1w+wUKzt3M9Q8KHIau2W7rG
dnuA/RqP1iBLuAjcBRbo5rs7No0xq212iG3M+5p4bVuvxldDyHPxDO2PiRhbuVtyLuTHJbr3TwiC
XVWywjmV1XGOZudw/JFudBxFrzHckAN6k3P4rrK9Bl9kGWkAqfCgrCIzDN31sdhaE/gW6XMVX34t
6nOAf7RLeNI/4W/Y9d3vZdg1YC15IIgqN88xFP2opnSi9McBxA8MXJ/SN70qUqLt4QR7bAemJOAq
+mLQ4MqfKkpmch6AZOniewUm2QZYxkCTTR5NEeZCdjnSIV6nunLPsWnkS/5etJuvBYkzeLGzD3Xx
gkbvSItsmeipA85IwM78xnOoAhYBYR/dLagjNJvfbSA/ZsTdNOYRpSXVXL8cfAYJ5Q+pZZIJL4Ce
C7jDY+3WneS5RGiXts72pcdlWZWwEiuQWxcLS33ntvfkliI9J13OtCO2U5Q7qBZtwSPdkWB2g5e1
d/iUmNcDrLswlyvAps8h/eIlLOmp16FhJwLPD3Oa6bqZ3IWqFsfzt39frp1T2uZYNqIuVKYovEMh
uhx+7frfz05NkAig6rWP4POTyVBEcay9cIzSzdMnEwVo++1ojihaFT1y9VpbqBGu320bNqxFwOX+
0FOC9TEGkuoxXzGQJftKP9PFOzxva0gjP9bYslNqAAX7kYedWbU/F9wLQmRXW/Cb6MVVKJyEMTgz
dtlORuQ08tbatu78cvLzU2k9txdrtYDCoECVxpbu+hg2J7KMF0KN25vKcL6R0KtoHiGxGKLc/Wvf
t63AucE/ieeNnOGrI0AffxgYkHsHJHiYWiEMBcc+veGo98MW/tBumW88hU3mjWreCc39sO4So3ER
pXtXMZWaxVZK1e4HTaUzsDwFzJMCghAbwA0M3PdPbderJw9EzZHBlnyBwrIypWfkcGlMiQ1et71d
tSUlPyYmY+80I5CA9mKotri3NjEpWjmnuyw194xsE9NywSjeLklR0eFG90Zzdo61Y1JVvm55RvYV
Nbe4UX3rvzHZK+atJJ2XNAINAuAem37al2kvTPnRWuYUouFJuHY2uTW1WOaDF6oylIEQdxwI9DeZ
Np5AGEL6DAYEcZMYQpA6QA63OBzXGRYn6CLRVNFueErLHxVFYYcqC5ikE7shga2ps5LJx1vIObtD
y9Yaf17KbwPCI0jHbypLtA1jQIr5RCvgreTzp8UUsWehv74GZIlmndPQDecHInb9YKm3GzSQH4my
QfDAUWplMUM/Ax8iKJ+IJ5BCewsdNvJllOiFTg9vpzUoXcsnoAlykXQVC7XOwKJMQuznSi5bCAOo
IZbOXgjr21RcwZDScQyBBmlR/dvG8LHtw0Kx7mJqPNNKh6yVmsHqYksHFPd6eKyO+JOUKfSn4HRH
+DUV8k0qWNvyINii0Z2gS9/gkhxv8mtKi2emsgsImLWY/a1OZ/t4uKWhiqUrh9WoSy/7U1W0lmQZ
9zoUGkaCSp705MiZohuag71pV7A+WJc5srj7HNHMJPErd/IsqU5uDE03rO6i5ywdJu4yNj3gK/SY
qeGnlK2fsUBl7y55RCfG2m8N0uWzUic43FI6QfpXkTeGMctJggbrGwOFtQdZ0fTk4gLC2rd2mqRf
N47GD2e38g/WzEhfEProIs8L1WE/rlbEyXlP08mZhlB4+cPwhjGhdTzh0qZ4tHfJPrQKlOyOtPzl
bY2pUlDnEYuvNiX/LU5wUpM0b5LLR6Tet1VZRZof2tpw6XB4hOCmwqOZD4TcrUhA1YQ6RAqLj0uI
6xyVxnHJIpLv1iYUDTLhJTQKBQzunGYZMHX5g7u8HmgYvb4SDhj3Hf7RLrcbXLe75PMqpa4jMBN/
fhV7F1RkpHzm1M5JlIa0fH6td+hHzpSfpTHvgI0WavnVP0Qkw7/NHFqnSOWMCVVo757mVxRDLSN4
0v401IqdpF9ZbP3Fhs8ZGdsicxGZSIZefatEtfTljKDOFpalq+toEoHJDlBo4lqZ9F23aE4UzF2x
vlmmXNq3AD0Tz0sCFWtZmsbAgEOeK7C/4IL2oTi9dHuPZ70XCCwq+y13hsuQFTVqRgfGJ8xW8c0T
4OuBbOM2wxtWsfHUvereFyNg3pPb9zkMSCXf8NzwAOKpqIKgGcgXuR66xjJ1Me33k5ySh/ltDOx0
yCWVtODtH+tOzde6ZfIXmOmyq5tqqP8NsfzfEy2ROfpg0LOzrodaxvl8Jp1XJGyu2Bor9Wl1MBL7
ooeTZuep4C0a9j9EIHy/a9OzPVrcrQTZMbokKe6E8mK0Rh1e+mYviOVp16G+5ANAQ1RSV7CmGPWZ
tT5uvGkG0SyB2FYmIK5t5Bj67D4iV4gI6Gu8piDBK90S2S08a5KNTbJ9YJRK2F94Q65DRy79iprt
/tgXF5cIIU3gBZ/DnNU4AkLvd4/Xd19TaKET1GsPwy7/B7Iw74QJcwcUvfmPHAwHfvbIGl6yVsxX
NVKPn6p0csnkpCPm+jf9Z5Ozv6ZQqsqxjwWIZX9+yqFObl+30GQ3Uod1hIPkHxaN6o43rp7PpVCh
6SWgCzcklCaWJjLU/HUm8E321BZ/1/NNR0VnBkf26QMH4a9Lnp1hICCmdsojDvXn+ti5c6He8pgF
qz3NIRiEsF1hGrWjsAob8ZrwAdzrN+/hqgTRiFGttQ9gEFeAMJAS8lMQLvaxP6mgxJQ00sXpCTbZ
gBhXKEr99qhRIB16isoVzHRqW/EROLbMy+eX0znmz+yUCMLEaLO1aGJRAqH70ttz048HHZl4m4VV
IetC/XhTdrC3VQgJ6+12J6mp5JZ/AjwVPJbB3vgtt3EQMF9iE117fC7dFeRwUxmzLjh1xbUcj6hC
quoU3Dx4hUcMjHozTEdW0FkDPIO8pLoMS4f68m2I8adgnF30HBBEDA1ETbtHiDDdgcxCNuhRG8pt
r3neIc5gA7PzQLM2hAldSJbVrnrYCmk35HRIvfXCEXrco4svijmF8rVtdrr4Ci7UPHJnlCisU/F3
dBFO4ZLwZs6NZXGTNc3pRf29j9876e8U259txyWgueSB4pSI85wcuT/KvK8TAuDm2JrtMW28g4pe
PYWlW/569zS/osY9pu6lKbq16j6F6xAlk4IBw98boSZFjMyHhccW7ScRPuE2HamhOR2iQMZnUlaw
FYQnkFKeGcJ/D38gOjK4k6Jf1/sR8cOxgnsdwVd8LYI1SJf/UFj+SNoMWWSaN2IiCmHhyUnPq0dj
Qz4L+bFwS2RrrArL7b1DfRq217rSUY/r6S+lP1GuD6iPQkydYxC0A7QUHoGjXlW/XlkIGynTCp/s
Bym2l6lxcvvKLAlhg/4tUWBpbr2rCzsAJq88d0jfBOq+EVowUtMKwZkZF689p36dDpNF00UG1tVf
P7rvGxc8vFweYS9KeTovIJwcjXA3KnWn/iQ8yGfuMmgkfc8AIyA7HWNvABbR5ZBxeJmrMbZ6UHPb
Qqg8bTZADPA65kafypTuZxWDJ8k5z3caboSj76WhK3l5rE5MZZj3jjW2HU0jI8cnHDaoJ8121+ol
P1hEICzFZh2JAeR0zsnLHPxJS4oOsnWIWDsAcSFjPZI53ZAxi2apwIvd8jnvR4D7H8oykwhQ9ZYk
mKpCuZq0GqHZumbZ/UBRaJdrSTPOydrT5G5B0ei7BN8h5dKL8zo4P/yfwaH2H7r8cN1pz5LwNdhD
zvlMMtZSKBqavWEiMvAKT0fV62riVdeg4bmPaGfGv0n1ZxI8Q5jyYeoAbhm/2xUup5XYTsEqi8hj
5GTerpxuz9EzplUdTtexRjZNuX1azx8PO8KR7TVDbCAIRhHmycxwq/9A6hW2+Y0ye+n092qftYWY
zo1Oe2bKhv0SkBJgzjbmVFiTP2dizT+Er8IPiHD7rIyIx9bmhwS106TLLX5rIwsUaKtfALm+M1jV
aUxrhau3SPnHMXdhBM1L4hgs5rTW0KWFIXS7a6dtWDNitYS7nOX7dF29gBUFgMiqMBmg2vq5kKWV
AKZ337jeoBBZDyLV1BDtKbj48byeibxYyQgEQ/9rdgKIu1pY881eq+EjwamDCH9m333WZc5j6v9Y
STbzvKWXwTsgeQxLqqjBay4eJN5HY7Mti8ev7Xw6v2umjNqzOapu62xaDB/7mcCTdMgbHa3jABt5
vLzGRM/dMbQjRxBXYPJaSl9pERQ2EpyO4BC3Y2tbGmVuHPu3Q98XlyO6P/N791bze5KC6N2WtF4k
Xps1bBg4dfyXHGeLBHAdeZCKvEOxlszvE6Xq9H6IukmmxfN6kgTFfxb8gWUal40usPN0amNJjNP4
gx38PPkqcEQoYp3V6SqabafmP0M1wjg/SKhZwrHHXXXnYsbuzn1lycrHSmMLaZMqt9kYrWnYNTJL
7WELhoOTQznjOt42MnX6ksu+SpYhvPq7eGVXi2O4AfqDG9KvgIFAi3P1HOLRpqDAWs3GsuHjJAY6
goclf4vsK5CKD1UvSGB5DaTU3CTtTgupKm3yThxC3s9A8ID+LmhgbxGPh7htKP2y6jdYIsRrezOb
HYwyowerEr0JLyHVysu+HJqFQAnNZHsyUqSJTtIIaxIFZ9R2rWdzfZrb1Ea/7Z8KYD9QCeRW6fUh
nB0C7APxlTGFsnKn7RajAZcVJ9uIlEAo29mewgvyBoNuijodb05hcba1lRG8RyqYziLvB+OuAA9G
Nd60Z7ocEKrzUD91p1hjGoqMukLHdTK1r88u+BZgkTEHdWDTcdF8A/6m+zWjXAYc0SnHUKiwG4Fc
pD7eAUXbWEW5JTHH5PpulLkZYBdTEHvcuYkp/Kd7n3xBBmcNm3V9b53hISl/2tnRu1twsuh/bC2U
aaxg1LSL1cCqxYkYHSMwZUyHWBOolaPsMVJ3K/PhgsMwqnGE7zSloToopkMF7S55OueguXShVQb0
NQfOhBlDtbzpmBzvGWHj/Tu5mgceCIu/QmPn523fnX9uLcBX4B1uP7Dr0MLJY/FsmNHRt7QAI3AV
i6xjm3Gz9ZllRyAyUCwPfIhmQ/TYk8/NN96eNsFZUQRH4Sme6vv30ranbs/4coP1CgfsgcVOAKfy
OOL7028BAtdgg3FYGC1UdCrg0GDXiwezQn9ofkVwWVDn/p5h9JbcFfTathFBALd4RlybwvVAVnWd
IFyajwrA7ftsLvUQ8g7cFw0ibcngOiz55TgZORaitbPiPUoRRKg0Oqs4v7RzB4/J6qAYm7VvR8CA
ERJbFrw8RPd+g5138ebV5ljSqxgZ0+X3JKdVDdZfX3r5VOZuNkYFO3Dvcv5/BfMFA+wk3jPFQMEX
ZDlUE27tCVcOd0gx8suxDtPEGoNHlROVWMskcQ1eLtq4cKTuvPiNdU1UUisciHQ8It7iaDZnjMfg
VyQobaHIAwMprwMMfWWVFszTwOycasxZ5V+ZrUzGBuPYQkalQ2BfliMBGIRb5J+nFZPe4js5Q3mX
Q2MQGb3gCIJJrdYPK/7AmDI3SF3DB34rvBudgAZMAmbG6KuMcHs/fYm0R0ka7gh7F2xAdLgpd8TS
Tb8K6ELy/Smr5dBVVWc8NrZhs04/V/S4jCxZnebE8rPsGnw8ocTmVheSxmFd+vX6ou2PiBvJQZx3
jg5pVXBGbkZVVeeTaJQuSQZDMAgT4KjYxYWjHsQm9ae4yhTHrKR47jb2ULLMOV1Xb951BYoVRcOG
Wdk1rgsyFAWQGaJh6CARDzcD0omWmMFSyBXChQLkxgHtYKlZgWW1hOE61p+JA038O88tYr0rx++5
82FWc7f7P09JYUeG5hzW8lTrz11qnXkymi38HH3VhTqFc0NAPeV7t5TVszvBuypfkV2CUzYYTqDW
x0d9A7OwTsBmNOi8vmyUO71Meziw8pgKre7SfQGudNK9PLVWMwHzpPOweMUnymUwyUoRyM24kj2u
nHqj5cyIuQf2P5Jvwk09XH94cQ9MJjL37BWWkRAX3Hi2JBYZVJOmlU4mv2q6Xd0ceAcgBmEh50Bw
TB4S7n9xul+duV7bTf+eEQmhb1VvhOUsWUbwp2mYHSO+3ZMyPK4J0cdcUgeSPzhRpEoKd5uPzSaA
4/T8enbV9kica+4cozF+BwIWh04mrY3RiQwvNZNqKWnXpDkgNDCqtaX8Qx/BA6KpIlYJPTpf74tX
THiZMxvH0edAa4cT0szKi/gDnBeilUsgQHowRmZY7EL9a1PdaW5y1gNvQjrK8xf872+zkTgGFyrr
s7xQz2v6iy6lp7YGyZdTKhBqHLlS1sQV5pN6xPl+s9IG2lV9gE95Sr+n0O7VH4IeaLHUvXWC5EHJ
SISlanvd9bEs5/w4gx8d7jSiOI2bw8PhpnuYiCb/Psc6c759NbSib17lPxbwfbBNPhYn0gV8Z16u
QXcr2/bPgCwj/xg3cioqzqPE+OoWvBMJaRijMmDwbEf5njcRzUSlj4/d8PalrOYTwKJkxtkUvD/M
6g/yHM9UdFAN5VV+FCQtPLpkmYMQwaTQ37nN9c41AzdEGQ+pKjGO/4ioUg12fGqzFvFx7NRsItxG
z8exii3rpPnCGvfqFlsjOPvfK8kKHydUwE7yzZ9WXyN9EYtMBRiWVnyZvPA1WAypoRIoqQ2UvQaA
/1Rw+hsf6r8tW6WejAjHovtLnhB8DecVFoRVIjjqtiPvCCFyhyBd54r9bBg/96E1HNom7usslgZ9
R80JQozFwiP5hJOEX5LNSp15ZwtxmSFygyiifbl3LyrWfZVjBRcV3C5gQIseivfGjyIUOONVpr5o
Fg4Il1nroZZqG3m94LAH5VCptbhvSegFpKoxHPmMKDXDgdxv32PXlRKX+cMxyYiQkO1E1xBOg1pr
ie0B64DfhVABPcjhaisBtzid7UCJVCCsVgBjGebSpSPUs/xj6PgLi7r18Vv0KvkGH2cyr7sUY0qc
ceGdrvBSvajih2bkzQ23nAugECv8SQYY/FKyoLzrUJw0cDFUZJPWqQL5arYa7CLfMqxFcBoASK12
78i+m87cxvpi7Xu2O4rJfSrzu3msqE0eEyzE5ZZwxQZIAnztOv9eQCi3ccNKEZIB0GoriJQuvZXV
wcZwtcVmJwP//jiOCXmQjJendzXPs3sgm6VFgrnyAQ6eBcCErjx/L0e0N14VCaUQexXSpmHxKHy1
uJi/zEC5gka8et+Ig2wZIHqQcokOQf2OZi0iKF/f/2XX+wtmn/glSt6A/RfhYObtSDdaIZQ0udTT
JACwqC1qwXpP09nofvkMTXb+N9zdDtbHXBJfRsBJRyJfF0HXnuWo6RMoZgvDQWrGK3SZ1mRgvx4I
5UG6X/LD0pcCk+Z08lduwiQerEZgBlxSvzC05JsKQsh09jfKGChFr+9ikstiauZvZ7h8ZhOSDaJG
HU7I5f3WgtRiJ76XZp3sV8J6nNy8TUNIIpBvcLYnYuAa8wGP97Opwxrf2lDaJlzSuHEl+a04kW6e
AX6dCPbTcU9mzG0CVhRNqDQXg0KgckZb7XQN8fE9wqlWWD2p3M4b+0KBNE1xkue/VNIqYwKKhOq1
pa32ZT2U5UQbaC5yS7oi7v3Nl+3SUiRfru5BhylR1rRBEhJp69skbYsRnfhqVHbAO/vQxqctPUqQ
ZIhVZidjc23lKjFU+lHpLPC9ZQ2ZB07Q5ZUq9WgGFz8bfKYrZ9NhYPYCJxiQqnO9Q1c9KX0xX213
Mqi2MrPkOTM1hkFdNk59NYuCqKzxMwp1QlNweK8bqVYLGL9k+AEcKKg9Q1TQb4li3SaT2aa+VRVH
3K+yipvGyMcsQ1bh7aoPy+SyYY2CGm3arQCrC84gfZFSXIHhw03nlZWgKZuc3/n+lf7qWAPC/jqF
2NjBsL4Ie7F3J6An9Fvx4Srm3pcXUNw/W5qg2YDSuxp5lPd93Hxx355M2Disa32jd3gg1i+gudqZ
l4NHR5rgQ7i68Z0qsrXbyKbrFpFoh3JKBwy43FuCisGn6VqguL61DchWR81tOjz6bmqFwtZGdkcZ
MsTX/7xUqUZYNnPBMkxCwiAksaMhYwfhpNUVGUx5G7oYtOOljSFGXngGnt7/xfpzuiOc45G8t3+U
MBEU/gG0hSJaVRZcKrvHs9qU1r76dSJwVmuKJ4r11NtOqRveVIdHRKec4mGEwuypkPGYGSDKgYwE
FvPuj3o54b0cAOMA//wSTSL5c0BUUYPl4QviQ3Y/BflJauf24yC/Cb3RYlCfz7SxvIeliKdGp02d
axT7tFf3b3bGCQ9u9m3oFHFH3kZEjzLnRwGcI8gXrsLBX8qv40wGf5lxdazOmFuSx7WtTQiBy2ah
fa2WVucTN1CnfYRkPUlbBfFlf1Y2x8afzxW3NivZ5pGflFigilwzl8S8Pmle7myJWpSO+vQrM5RC
2EEhGb7C3Nzakj3HCkfMMM4OBJ+KdMszeOBYFPQr5PmZT+GIRfMoPkel/IRKS+hCG21u4Gs7aclt
3dm/rP6BWNGlB6Nql925PYlEtDGkJHFdvA8yV8tUwYuX42RhXC5Q9ALh43okfVk6/5PwEZ0qkY3R
lF+iL0t5+M6gHp4NvlwoSVZN67nUBwO5Khn7yBSmeX9W3LhvcsA79aHB9nWqH0SaaltvTU1e7HhN
PLK21pZleWUgztk+yfobgrubRetnvnzrWWoz5IfBFvqwPSnhh+nMqMlc1YAnGflmeiTYVYI1Ok5k
7hv8U4lF70KODLOPzSHMuCs6MbehtcnyYiGqWVW2mDqN0rcwob7J9QO/CYIqU8XSI73WZ9KXWPWA
S8MIpOXH5d0Z3Nzp8zxMFz43RPKEkkQLaV1K8YolhEIVTwy84XOmqb/alWSd1wwvU08oSrHm8vfU
pDDzv9pQ+O/mZTMLbaKVoLz1K4pNx0SrHeBnx8uBXHvc19q9nIkrdbgb6691f4tPfhUokrdZHXai
M2xos7TFOZnSNx95j837eI1na9vcNVhzfIIj/I7wQx4EG6m38BZmX0y/pySUDw6SBgI/g+H7uy4j
qF27gTNMeNEn9gCIB8+qS3rB/TFrilp9HNwPqY+oLfUzY10rWE0P1WnNm3Sxcu1AdasDw8twh6u/
BYKRsr96rGDE7To+8NqzoKeIaJoTCmdFeT5Jou4dXAfVjQCLh+wsEkwx82i3ZoD+Gt9hIRuwPMob
jqXfPCHZFE5IriV9egJ1C0T6VImZt4zQ6lfC9I82hL5pIaR656jF7c4QyZ7/tFdaclhXNfGIMvNk
uGF/Ox72EgwYASV+k1Q6gIvpu7Amg3+TST6opvRrFBjZvistEcuYjM14hAyfr7y5qKhXKPxbqydG
dA7fTtfXUBW9JoUahWb8tD8pKVayPM71CHP5silSOPQBfApUJKN32idNFWj2WD2evGbn2N4arMAU
Du1HHR3O/xfNkGpJrbAqeZsIPYStFp+0aNijwBf/hKRI0ePpBxhaCSAV/aQg770XVH3zKJE1ctG5
Ktj1NzDLiQqvr4SKmYjwC1HrXaMI9/F+RbhqbweUXdZU3YS9jnfaWR9jDPpyfoPxDWd/pOqs9rbB
wzZhz6gaOYKxnn0dcfTQukSV8r6xVG+lhrq3ipNN+1DUBChdCtqfHoC1o/cawDdPEABQ3MAyL3Qk
wksNjdrFAvZfUsODSc4hMX3FbEpcFVyrscCOHgRghJaWPwqbEHerC4ngcyIhql22LZqhnHjfeTrO
9+oGYGqTJUY/DxF06Kq53GM447/cTT9wIxv5aHzogo/7wTzf6iXNpTrjodXSGkslNjy/g+Sqdejt
DeRGz4PfGki9+TSq0mXT3kTD4SouxBD/OISznYXunJYnSItrcctCf4FinCmXuvs4TU+pFKNQP2Dv
WhG1vareiegwNd0gfdvkpo8GYYsy9dliip4xJCVq/RJ+9OQognyU2a0/T3YtR/V7Wms3FoDW76SJ
qfPJQQtputl50Vp1QgaLTfs/6fzbILa/3v/Gixn8TzW8R1/81ynRI4iEp1W8++KeeaYrvwZqSh2f
55eePzZBq19+0AJFIDmqdr/tdjPfazYHtLCwMVvdovt2bcThXohtAtLJcLiAC/2+G/+ObSKW8vAc
qzlSNUThP8xECvoBiPGohtil0knAEGGfaHegbcZcK8QK/F2MWKBtrS9S0OwjF5KxEyOp91CsQ14S
nORAyJL3PpejNAivSBgaO37YMsKTSnGYl1P5hqBf+lpPJeFv51tWjLq2aZy8BDvLIcashNqg5vwo
H1G7JSXdDNAOZIUYNRGzP6I6LyqxtgiXDGx2TMcQE1nJwq2IkulOczbe9v512vu5w1abvLMTfcxY
Wq0fQhzP+Fg/xx9rLx0gD4PhAHJvVSYpmA/P+jdzYuJS9piD+9h8S0XLacryDkErmlza29tV1E1u
muBzMiAiG+JgoLQvf4EmH8G1+UosU/EiD5rfSBDq8uGgrElVBr6d6cKI5Lv4sJkWf+TbHfR/9Yyw
iz5TI9Mz46FA2doZLAwSyJPfGI2B9p85b9xo9xq8jUAEH9hS3pDWnqQhu+iONZD1iI0aG3ERxmR0
K6TZAiscxOLt/bUWA1WcmO+26lla+aySS6//+vP+EVSyY/3BhVfyGBZAMEIvt6RcBZrV0wHuEdqE
+DM+utYB0bcW9MlOCo3xAlEmP9vJi0K6fHenAyQV4gF73F8eQnSMWT6qxBElBad64E0RhL+CjWuI
73pQ5aNnovuqZyz+MT80SDh+n/7gAYmXsiwg5sJ7TGnTgQl2cmG55f/eehHqxcaXQJrT/QZS8z9j
vEOhmKnPlq4PAARE2CcgluuJoIz0Enixgxaolo7Ceyqq+TpJp55CngYQ6Uh+YblMYbgcWP6+xwsM
GCt8QVvjwtcOG09VtEt0JCY4Z6SO7xpqF3cLlvgbWl827hKG84VNhL2WqS0YxU0n3DvZxBm/9syB
/dzyi57bbbMaj6rEKbtTk+oR8SKCDiBKjXdB1JYBBVqpEhqv+DrtQnfwL53CSlQLcynxgeulctTa
V99VaBOyFb+kQeSXRjK61ME7RUu2Pk9/n3B5td4OH5LDV+/8yvSKQZW9wWHRtugpp9m4miTiH2Vn
4m7tXobG+wWYv2v26ZaVAMC9PuNFsqd2qrH3Kstgn1A3C6LVL1NFnUsPWxY0STD+L2GE++dQ8nN8
mJuQ+URR7dzfTp5zhG+1/w6BtECSTByyTZWlnkqM/ezH2+e5F2x1NMaXP0XscdGSIIoSiFJBqGZ3
h58LVPww+vxHPiCobpa9GMIT+W3jvaZZU365O4upKEPDq0mSQiuGcgAyMZwSoZcBBzA3Ky6ySM4t
9SxtuX05NGlSQFUPHeltNXrTR3nAseTOSLMTh3kv3Vy/jBMm4MFnD8zp9tlxzUp7O46iOevlELCR
dto3hz2JsGm5y/WxLoRsyHAjpZ3I9pLlrQ2/mQd+FSizAjnRqwtsdjyr9NDgw7kajAASSTVVLwt4
NgGbF1+jecAFc8CwyQB7H/qie1Ghg8M3+Ts4BqoiciIiX3DWImk6RCAd7khVlqIqWGtIdNAKrGWt
PKlgOk/mBINf2EbhskP69R22VEp8Kvd0iYavYu5F9iRi8HT39xURL9+00ZQ/p70UjebqhdAB9m+L
6IPyo/JeOl6/Sf9iDWExcZKHdvaI+9D4cmmkQLTOoQVbRW9c9iJW33Y1+oI1mSCSbyUy3c+F+Wvg
mmJs0/D6b2pbzM8K/nwpzthB+Kl5RqpfZHfCa2cnBSwTAMjJr6ZfDOWfsPX2BNCzoY1Yh8mtBgAg
PWshhqaE6sCcYc4avl3I3pyLK220SA09G37/ZpZHDKU10fwrGwr9IPEOX1UAnvZo9eSueLAylLgB
SHQjQQJhVeVaVarKPHf4cEjJEmW8+xLbfStZ/L1CFAnN+03ymARirlM87LnYZ2+yLquc9Iv8bLJH
MVn6vJrFqH1rp0d2fB5sA2cFQDhWeZT2XrQNEvDBgQiyNRoiehO1NslGGPxBaqLCva9eSKb0WfvK
5WbmGqymPj5UfnaL1s3+COvaATYwqtQ87oY+EFb5M4zE5eggjfWta2QMj1WQP9Dh4tXYB1erojAy
m2f9L2LXSfdivqN49gdS6KLvQEo2mYXlikOFyA1JQOSdW86mkm8yl2E+J0GL7LCUtdSGFPfPMGmJ
wZxDLHEmeqsHS8nsDuX11ytt0DDrDOTxBFoPhD+sHeV5elEr6tbK3+iOPn0/xmTgBbnCJBUx+1iS
POw3Hs9/18lHha5WyMnqvpGFd+2g6DgaUUF0hASWCoky/U2V7m7Idg/PfEWaIRMDNEX29Tprtq5Y
rSWeAH8/3f7Z6UgWSiSbVodkTz91OFLhmrf4eFvq18GCH7FN0OuzMVrsSKEGVqxkEMehMU6wCaCw
YT863iL78ZQ1oRiEGs9Qh8moP3LFfisDYwsNWOWDdUjuS+KEj5tZhfrdsNfFJKEc2ePlt/hLSopL
WDJtpfNoMDH838tCCVw6VmzpFrBpKnid7VEipeJhSPPKWZEv5rVmTwr8qFsdwn6+4nBje/hcXOCv
R7HNBt2YnWhWX33vSiEjjvYiiUaYQgDqmfl7i1rms0+NH8af9Rgin9Xo0/rVogU6LWbcV5NCH3vQ
eWdKOu7lGDLoboZ+SXSvQMJ/XD++uhBVdobimro7pzZaPNURAKEf6sYyT3sXpSEsLjk/eezDHlsr
UfsHSL4Kwc0Y1QkyuiSLhbovGBi896kNdj4ZdGMSdJ1UHKbfHmKYNeEY/HCNlC7Gr0dtW9FXJa+w
jakJXKoPMT9t7vT9X/vDFlDdcSUVFzdhiUlAts/BHUsrweNoh8L468RsoCUbmL4+z7lZtmrnVv01
Y33shgzp6a4ldeS5ku7gWBei3Dhu9KJWhImjy5eg4QNVZk5vdbXAcpXEkOueJgTMMF/qlFCdaQ3R
e9BkImT2k/pg9tmR6fAwkbPxrmAqdFnJdDqNsZHArrItiI9TV2+Qls/1JraYi8NSGETYxaxB26y9
0o5u9NWWrcto7t7sLJf9ji2Pzktn8n/PMguNDPfvfIs7HbYmH9lfFcU1NpkbbfPwIwCeWemPZEfW
a/NpDIfIzeq1CyIHK8Qh3YZR5njp8FoLUG4FdwQiYPyVC+pQBfclv3S/CKvdEaTWshyDM31S55l2
nlHAYsVL7oXFaXUFfWVrouVedeGjAIQag3x7oKqnC+XedZMVEhIqzNBQq4D8pvkwlKqZ955cAttg
y817JIMbJi/ccUcGSFXTl1dxgj5eYTNBxHaSK+I8MXntpD9CMiGzJ+rX7z29eBGTyfuMO6mcYHlJ
mcE1aJTUjD+NhlrRMD3YI+J7//u9lUcroS2VB4t3lzuH5Mw9b26oXLnDLWEs12cboEZ2WjPekzas
qnWt+MPJcEiWMXjK6FfVOZ2mS8rVnHyPeod2H0d+wwkfV6bzaiEbgiAANnggYZTBq6vURKAB7+OW
mNHKeJ3sSnrEGY5okM9VCSEx22cIciACfAViVorecHrpimebRgAy+/iGs8p30aIRkGzddGYzRfqU
YpHSfqkXJBmPltR6QqPvVWzrWT0+gORVsUaJsCzLn302JsVYl0GXArNvvgBCaFE3VjnPqw8ylIm5
mOmULl3Jevokv+C8q0XpuzplKitfntrl8pG0fZbgvWa+sJWsmggBc+zqEZ+vt0NeyiDS0HIKNl8e
QH7ysBQBrJjEcTMUtSdy78HukaPzOdFRuI0XPoA0x8dtQzGL2W8fdl67RWrfv+El1HP8hqCBwjwD
NeLsOjIQaHx9Kw+EsXQ1CckbJnvQJ89NyVJ8Na/gntHK2afIY60A/tQOoYzAOcWcmdwKoGAtn4cF
t3tYKuIK/WT5zNYKBKOpPRqYJiaQXAOyHk8F4br1aDiUOaHDQXv6oQsZJDBnt5+B5kpjHI867WX7
zVBoVy3DMeioGHqtRKYT792bkl8LdaGyw+g7ie095GU6oef5J5y6MqEQQ4MgjHiJelyHstnn4uZK
eVl1w+FKIYRQgIJExa5X7UbjYM5osZCr66VEfZZyfWrU3U9MfEaCtzmQSLPPZt8qBGzS2hKWdezb
eK/bd74BP9q4hckJlfMzbQ8oWNvrmi/r25XwzfwxWNJtgpa0vhlOVSmgc+ZOypgJ/HwsKh4r/Psg
QMPFn/RIRDshtHpDQbZOb7If3s50blpA/s9nfB/8C7QNtsQoZw2mtGyi3BCK2g+b4ocNRcXW7Jp7
NX6iK2d2UwonuIyzjY5iesC/z8QnnbFfJW3dqINjQOM0Z4rRQiHg7jVJ51aa3M1I9mdTYc462IXz
kUJWICXxkAZgpRrxgzQIjg1BkyfRCX/D7HgynZmZ/jVBqbcHq3OjbrtcH73JCX3/FlvyvDayeY6f
NlIQbDx46AVqe5GfPctGDuC6Jivhf28Put0EM/cXf3NSd9qlATRDOu6DVVOYX+yHL3xz+PlHcEjx
KIc6pI642+eMeeDTeEyfF4imXguWMmSAcNs7kxAJzmddn/e+qAh80xuPkjoJc1UNqnsu85/CE17E
lQaQg+EVYzJ1cHbKtPTazedcmvYFBiZNI0yhY2SJ7X1FySKJbbp49gGGfNk7oMxsS7PkvWPE5SeA
UVXpc9ZhX6/fxoji+hpoTKNL09EqO1toMT7W/6znv61wEScfBl7cRnE3wYA36sR2/HVxSlWwz09L
0SK4AFEFkNKR4q1NThD71djvnNRHX0oylM+m47/2Bc5PCg2p6mSMwW3OaeDWSPFzyLGTDB1wjPNw
HrwDCSnH4NOqyRKUxWzFScWF4U1Zt8JPNEtvG5JWEZQmdZ4kZVKqKf5iTR7i/khi06JeLQMpC03x
UhP6f4kO1FpMpw7aArYr+ygeZa5QpbE9WCASyZedEUT4PALJ2ge9LwMGU+6QSLuHL5EoxR00It8T
ryyKEGB2EROfr7hNhNkviyeUWcrlMiUPNIaPAHSnoy7djx1/z+KYTfIuZGTTR3T/4izQXrAGzUal
xEldYqwvleJZ4B8CNFI+ibIAEuMn4BuALXhhGrq7Zc96k1V674haHFZIxpzIOFoUCLoVcwgdMm56
8wue06WzFwiIg3Xy3u+PzZb11Q/ZH4KFQHStcBM9iMDlVEl44azxnpPXCsH29db7lFzSIlYTDGgZ
qRVC3odHMHo4og39lLY7hKxQhm2Dypo5ryclBC74Az7ikJhpllasP08VrU06VZo2skFqqJCO7GDr
GkP0AikfgRQ/lVRqP0UyGMZ4S4xkVLLcm0OjsTQP9j+RnEyFke1Zen8fJHhjsnKuMQthG4vO7Inz
7aQf8FfW7hAZcy3QRSMCrZHrTY4yyMA9RR79yHxQ0enR02nhMQe/bxBCx1NKS72DuVDsHeWi+KtJ
lBt6s1WN74JCpTPJEQI8YU0XuqLV15vmFDn90dUBWzWImQxTcjWQoZD3aBt2o2JsO0QQ0/DjPW2O
NvIQRDFG5eAsMLWCXzSfWHIhgJ1/UvsYEHCgD2FkULm36wz4LGisSltfMLU0Hyx1MDAsn+HqfTUR
yqDKBhJOBsxcOmJ1WwbmxNSykZuVHwIF8laS4M6Y+r9Mn0yqjEQEuOu6CfPDsxcnkqczSrbItvM2
CQqbj0SXyu1d9lVOsRvt7AidjpooZ5CgX3P5p1X1ADktWDzuwNF+aXqJQMUw2YPKWVEmBAJkxg3W
Zy0o6LupVQq5ouHeGn/O1t5VMAGNYj57EouuPgx3shw909YNF1y+YQa/K0s195T/HK+5ThMQAmVh
qbdkuFwBTPA2Pxs56bJIph4bFPOTZYS3FPvSDCELXA9YS49VyzY4UbCAuV3q2nzFbUJWhioEgyW8
7Ac1nnqodUrJ5Qdg6OF2tTuM8LZBo7HLeQfReMl5/t+artCcwRp3anm3HIjkoqLutcM1SjxW1iyN
QdTSOiuZ+uHRCMSrVTbMy1WLbOP03vDxkFy5DjEisyjimaGV/KsL7KK2/sEfDxhVLNc8SEEu7bMb
vPcTnZytfATALdeaU2hMe+EjE06cb7mq1PVuEhRBGmh7EFBh7rtvMIbV5/Pa9whyvMQ6ZG4MmGcz
VxIsKNM6ixdduKxkf1cmVYOELisCvG1CTDALp7fPP5u0XgqbURNISv2ct/+K+o16svg64/ZbHqER
5FGYrCv3ju4f93LSja2SkYVWaVmXDHqj28Ic2clw9z55BpG3ieLl30614byOWcWEWVrh6XE0RnfY
91gG4yLeOZ0blY/qMtI248hCzD136lO4PwNLIX0fivtzByn1yht0wukMuiLNujdS+6AKikbkZxqu
cvb+EKwqOGypA0AweXSkmcOse4I+sPyyWGZAp8P7kzMEXKYQWs0FFzn1nzXeHQQmq9fp/bpf/OoN
pma6K42XqWUxeAn3frFGjgVoTP/SRypVAVB2AnNhLm7hP49eIPfhVw6TLLFlzppiEENlJrFiMu5W
1OpHf1fEnDF7xbTHVSGfBKVuc4JKUswWX88yRO7fsb135KmNiVX4VnwumHQq5csHFS6wKwlCJMXZ
x+yxrnCNiEPBayYmJhQE/M917LJsyW1SRB1+1lXLJbjsdw19UvSZgmSv7uXftLug8fA/T4fIr+1G
KiqUWwMNnup7GyKxslHtsYOP7dGZeL25ZrVHXrf2t5hXaPijs59CZhJHhe8EHgY5YHn7Wjti8B/F
Zi7DYn/8Xm05ChTjnY8iTqK8/atbCVC3B5NGYu05usjENR9ClpOEt/gmpqcOYqCjE1zni/0NPSRn
ecDHZ7h9bf09gKFn52VC2fK4tTj8kFrWbvZ6y1xXzRGyPwJ4O/Ck7RFcZRjplIlr4Ccs5BCr0wpn
zUACjNcSFqh+CrMej7CEyFU4F4/XzRjFepOxqIB0r43Tg7dgb6/r/rDW7RTDh9Ssl9U5/yJlqfXG
d8P8SLhLNLtKIy+J1FZh+sbKxFM66eFvexKwJowI+Obq0TPE8HfdOaUlAqMt+DdTh6mlYKSTbmrp
twQyrB8M0si7H2Ivm6fw8i10EIfRIdzFuSg/57eSzdbLatK4ea1iNkC+3BWpWG77JxkWFe4bY3BD
wxKN4XdXDPTVQG0zINLZZb5IkPSFQ/5O5jCR+EFhzqxqttiZZQY+ZiC/B/Ps9HXD3MzLT5khPor1
s7s/RiLJgdFdcjOWtnotLARqA3UUayWw0GPambYkaqhzGSyZMGrwEKJCN3DlHU0ueObT/Qc2DrL0
leE+MF3IFD9Zgb9sXv2k7d0Q23xnUSoVZ3KR52O9sRwD5cHOMND7FlH2QHIdZx4KoKuPQC+1OPI2
ozwrpueO5Hw5REl/rhg7FvbvQ2R4xtPQW8i92wTTUPVUxmI+dOBhIbM6DStZxo2JB4/6SBjjRoci
7QgIHBWgmK8kVXMt4bHYpsiSrvkKoS2iD/RwJc2QOv70IRWQaeehA1KLH9jRPuuKhYcQKik0/ZJ+
3y9rBPiQXmMrLmmojY+VFvTIbtsyU6YkQB+YzI31UDzVekFckSDQyuhV9pbuhcxm+/lSpqy3GsBO
XdM2/yULj4aGmL7jFSrKU/Koor7cdIY0aooS7Bh8k1uOzKMTl77VK3Lpf05pylxcBV/hPcXgen6v
Vmu0btQvb3Bw06Pv0SDI+2SfbEo/ceWJTqM0fp7LwJEBCE/iVF0n0Q790DErPsBa7vRxXDhGNRip
9RIDG4kBD4KDcGiMtO+pbaTzMhoeZhBFLqTEHTxSXlzclQLcdxzU8GQNzRRglT0TiJgzKCNGDanw
8JI87H3vJ4okbEC1Y8dt7FZ8LkpMaq9+7CYmTetkOjPzO0VBMZxQ6LRVljGS+31uMl7EwvVAIc7/
pCvK0HJgnbkFOnApOKFDuzUQG4uueNSdK56p8dLOzHc69FI7a2n6ogCPyMh7EajUC00QrQB/isuJ
re8aXOfNGmCS6p3rnIUJnCMbhywRAH00TlenRmatvBDtX6RkkA+zjUgGBc32FQ4uRVq80YuxNlMg
Ukpv8+KYbG7cpZfNHjoZMCjdHFLwsPbLB029/2pUMfShuj5ZfHGe5OqH+GFdPsS+sUgsImwyAol/
dxr4WXQkJBYWo+yelqrQgl4hHqbnw+eZCs7d0bCmYQtMu9zYKKE1OM+ixU0lUZSaesO5TByx8iBX
tPRWkLiQ1G165N0TMknOEyV17hG5itlgXVnKKpxiQhWl0bKzarg4H5i3mgdGIZuLDt0psNhrB/Zq
ImCeqCMhhLJZ5uhpJY6e75hE3EzdiiV/gn3dEPYwPouq+EWGsaIgpZyGLK8P0FE7CJBo3/glfzLv
tm4Z4i9R9oOGfWXTvLj4n4u8oq02XRQTDKsnFiRV1+Gdc0VkSsLQ+StGZib40me6Qy/rq9nQhyWI
Kxeq2OWA4sG2OS0QxyaIvCaddu9cKgyYJTFlWlH/FrOZgT5uFCUthEaxTDNB2jQl/li06bhZEEi5
CC8Vsy8ESP1IzTTHjyXVufQvcCO5r/lqHWuVCbN/AZ39t4y6HDiB02s6g3/QyKKKMvXvPcixcElW
Pz2pPr2RN2W10vBOpnBD4SBf9Nc5CH2tXId1RfOqupXdfm+cXvosfMSISRGOZgmz+xtIqUbXoqkJ
e9fAUVj3aPm7Iexm10pggrerVH9Y2LRaTgHPaqI5y4vkNh4Wb6QrxjPoPYkeX9ThlKM8UIQLBURx
+8pSODkHU0yxZ3NdEAQs0GeR0HinvGsNsAKThcWQxNdn0rMdbkzBK4xYTN4h31TerW2CiozPOLA0
oOOiRX4uBGRdzqmLolMyp9wpqnDR2iJ/F3FcL+tElCm7JBKU4uzNgmym8AjQDy1K+zsf6HF6x1ZO
caxc0N6zWMWhCEkIQVCL00NOhN2cofBmyE9nWVXC3x8OUedIx30SYBBhkwPS86qSwpCQs4vkVqC+
lxdOL0Q02aBK1k0SlnEvta1OKv7ESFQr5+2fgkGgsa9Iv9vXOqph6Fg8ADMCMeR0TRBctZooCiO3
QLFfGEzEkqjbvjIgmBMTjxnn/B8K0R/s/dREeww23bVAD6htNTsiouy90Ug1Febn6i4Opmeszdkk
TBuybwal7Ncd5VZIMhK17KpZGVWdSZs3lGF3V7RT5u2mH3Nq6p/jEOfhakC9GCoTaBOytavzoRIF
VHH4LpbCtOYajE2rgVoW0lVho8maS6h0lx/1FykJ/UhgDUt0kz/CfeWi6NQI9sS5yurcXZiFZYtD
4giJRR1S2RxcvSULQbuC4IzP9Yh03jCZmJ7M33A2maEh+LM3eGJB7jYrO4y0OLNmz7oU4GSi6UCy
6N1BJwk84XLU+Sw/BHXqgVOxcJPM50pDPkEKGFiGo2ZXGguHKT2vbnxCudb5+Idjgyi9nca7sOOZ
KHxaOiixJt4qI2R5Mo7x1VnaIsW501puOmyjTAG1QgPWIm9IPwgLv0L3KnISMP56Sp+C/ZHhkt54
Tq9m2vHrTZsvOlVNjzZHFRH24z4QcVPlAzWx1IwS7hUoWxjdfSfQNcj1wuqQg58N84BodC5hGO25
Z1QyCMykw//88eYNwpL4nxCOacfuW+H3LciH3sMB8JM3AImM5v3ldpPE4F9JpUHgAKmqy/VvgYLx
c6ua+2YpRVtNCFz/lMpHMcs+Q4BrDlbIIHbLGRPZsqC+uJ3FwYuZEkRYzPtwdllD+qpUjAIDCdNb
dtRe4/Op/YpK0b1PaLPIQGeV95sRHClc619XtSbrMMESIe+Mq8TWqVPiTZBu8tiPWNpgLTHZ/WU8
veT9GcYTd1V8ih/0wqWYWuTfh0ag2EfUA6+Ay2vrLGmFLNJiCyS0Xi8Kq432/NcO+bk0mP3GTyJ6
X7OOZVaJunzVao88Go8aw2dChAb7V32ERe6IuRB4bdd+uQ4q8Gx9nMj39lPwWhlf0jGL5plsxrlL
vgjITdpvGyg1CJfSyQXFRVmOSygZ+w1eMO4TVehcy9dbJudqS45sJd9wlJC+h3SWgV8AxwraeWvD
sRBMZYSuJ1iZ5Sk9AeBECA6oZ1zWEmk3zjx2Ed4lU9RYAPxKwALTpNdN3fsS/+btq25uCv6gqzy7
8D0mWsMHXSpH+1Fm/YYNj/SGod7yjBzh7ByKf+QyC0nmr3nZg1/LYL+2ayxjNgwXzPWWMQoH/OHJ
NpWYF4PhvzVRs/q2H6BjbwxceWBa7kFL+YMoSiwUA44FgFcfaB3/W173JdndYruhgRaos3hqyJff
CQNgCpoiqZH9NiIDMGJg+I/3rN/Pko0OCeRd7qz4kpMTdLJiWUdQlsth7+xqwwrCj9zzmo0+ciyb
eUD7859XvSjDwkkaMorJes4cY+L/RVKuq9qDpxAub9rWnd/3wxDQVXUfbRtDTF/k7mZKNkoLTI2l
AkTKaf76k3RVGocC1B9WBKvskNULVkBj0Mx+x3MfvXbOzFzV/jV7JwZLdNuGW/ImC1dRjiX6byYt
e3soUGzKEFPBdH8G3Oc5/1/7D0ubcV/CxeJOPWPjqxtb8uOlGPsLhLQoBjh+KoArynHxNaFotlSn
aWAw3+yVYAXvQz612lwMHm0rpUqCcTaEX5k2hPMPm1mbgNhWropSgUu2na8dwaGbAxQefKraONVH
RrgyC1AQ7giv9uKGJ5wEBPZ79hkojb3tBA7kMMqh57HCglXXZ1HULW+Qfq3hr4k13K4NZ5V/GZCh
PNhZWFdkVBeJ24KoFVZ2EGLm+AO1HlwDd3xHhafw/Ji90nFIlTxkj/fRaJovki8t8P8R4nW/Z2n6
eQAIDeoSatsoaz9juDfWgdY65OtDO1W3AFj0D5CzAzL3PmHFuhM1rgSUlLOC1HlUF93BG6t639xH
SlikLZgLmfOiKfNkMrkx2yYBdVZpn2ss2EBtTXniB+QSMTpsRk+QfshVgY97rRTsL+adS8HXu60h
MYgPYoOt44zaZdYg4Kx4/F9mmc3zhhZviPRHayJmcm/EIkbhO6cu/aQnrIEksYVpbGVkvoDMBp2x
I30ywHLPWFh4WByaoq3O/+7FBTJ+nXvqCHGSkhRZEXjlYQ+hEgq1IxggUZmGlJrs27fPMpgPbQQt
8gg9/qC/I56EAAZno165z9wUmVmf3gDpDnlZ1BKgAXvy5Y21o2WrnINYQMPxrh/fUU5Xo/Bv1/h8
K1Ao+zbjUf3KpFG+u+jV5h+oCKweZBMObVEfpfjWIG3erIGHQZvGUIpAzYFOBOVGAL1JAJSJELcZ
kyruBvumtSckEpCpRMrh+RFgyBM0N8KI5NFrqekcun9nSO0sKAYHn0QRbmT2J3Fc/CpLKGxRN54a
QA0wIMV64A9DGGbF9YO0EETNvmQ5be0TOAOsd+U1l/xhiywFa75Qjjc9ZPkvxDgU507v/o0puy4p
EQ8GUD9bdh9YL9/mpIu7D7cEoyPXyItEPsgz1UYoaWRtiIGAT02u9pu1tjl/mY08VxpfirdMPiLc
GWzAtp79YLcHTRoAO/nqPeV8TqvlwALIDfs+SfFqhji0bUx/z9zaO5Q2ybfS2A4j3eBiqMz772Wd
ptayJZ9BF2QqIwvisv7Wms0vLTlMHsANR5MPsaJsGljbPCdLGohaTcmGxStOcTzO4sC9l51Vx/5R
pTc4AZElQsdY7IJojwqbxwu29wfsH/4CDOWp5qLsKv51UXYCU63AQgmsvVxZ5BB/Yb73dOs/j9cx
bPEn+4FYHE/DYmWBMQb/7eNRRcJdsdvwdJi33jfnmdk7xbRoNlrBBrkO6aNEN+0H3GpWIqW/p91I
x0BTKrW2mXtEIyu6bjEqmyKljOpdyFDBp47yfJqMdLPLI2j2k28TVAjttkouLX3Mlv6ZSY2gAyhB
DzFUSW5eTRl5KjIf8C433tMrl+GJ/wi9WaRF1rTD92Nfkb+zwsYWMcajNvgtAPxPARYbFpoDAut5
fDGjnGuYX195rDZBSRv92sg1FRgBvvwasQmoxz0hA9y8toqVSe5yv6Gc2N5W//g9LWaq1zJeLhLL
jwABx1rFjUJjnPf5F/21UzM9nvBSyMyqlNeGcldxKW5Me0QsGn6Nlk2rGwydemNL8htL2LHU1JdG
bBBgsCMokaMLbvyHraPjKEEKn2ZQuZePZOf/h85GvCE2u3sNUnJwNGqSn+AQF9RidfzUOz5/uKsy
8UPAtJ4NjnfvUjQu10irmaQC2miWv6YZZXkDs4I2WmDm/0+bmoIJ+Lq2PqInfXGOi4kxHoBsMvWZ
GroqLvrd5ueEVd572Y7UyPC+CEhSm0yUHhfivExQZ4tbg0B36FLS/q3RiBfHOqMb7wC8KNYuorPl
1nBM1Y82VOQwx0lqhhQg8/knVGz0I/ygQSodLlhTI35ttzdfN9g29+gfvV1uwxtpVOnIB0wa2L4a
j+Ghb/mZmkh+7yCYm9Gyk1jhdua2dtTFYvQwclfdp+pOI/nvPg4yaWiZz+cAq5j0E0vas+C5vBvz
0PUUvXRmwLzbkExHUL9hrjHmq/NFXX7Vuq8/8+nGaMkYjXRkZN/itc/lWMe5tr8GperVOb+O4mVY
BTXAAqTV/d/7awXt1mzs+AxLqO5GqF9mfD6gjfKVke53XcTv5/RwF3fhSem1oNBsGB5beGlkCInJ
qggkUDT96rp2Yi7oapwQG7jVYR97keCQCwYHoKuQzzyLe16b/TPt6aW6duyrQIgUMUmAnNyaFiEH
/6zetSYOXjtBcFXvOz6FNFXa8Q6G+RktIMzzvXbmIuD30h0aMT2h9/LtZIFSCHxGsfDCIoG6mD1I
jUVgNp54cu7P+6JfgHfLYfLED/AOIayW5+gDPDjxNVDQ+khg+e5WxlJ0fbgHpiqEFMdQv0YrJ3BD
xZPdQEh5Tllb6ESdVwk5gVJGNx0t/vP6onWmRUZ+g9RyozkUSc4ACOlPXiZSM12GicNlixEOyba1
4hJ6FIf6q8eHUbTL2hPAgMS6LIW9cTwVlTm81sQB1omZaBKZmyI/piOjJV2pYxuegu+KTAgLr5Xa
B9JVEdwuwSlxWQUE0sCW5868Mo4mHGFychRHjDnrZGKSM8yWFpvYewd6VSliONOg2C3enI1yhOUI
Nu55xigUx5pQM62vOBRzLp3PwNuI0+utLSTFYlco8wnzOxXUudBDGbqx4UPrFKR89R0/VdLT/9Yh
eRJ8pf2BoRBPTtKH1tIJ4O/ecD+9Fbv5qn7+NqOp8aeZzAPN5eYJEZ/upXK9Ig/SGQ4XxWtvBXPq
3rC6OK1Ql09fZGIrUc7UC6GVAN+wWVi6WGxgSYGlcoKTp1niasa2MjPGI31IVl6aURIo32oU/Av4
mm4faR2L7xmdeDNbxMpZtY6mV4v8eXIMq6oPvOj9dhNwoisjzWCVMg+7Ts4vf48lo9TeA5I9K2ti
1dFGMR95L6tukxHiugVjHgsk0a8+Wt0im1WZBevmEfkW46U7GO8/sUdrHqnNMtke6UVm4+ag8Gh5
Yp9i5/lSC/E4XUXqGw86BaAyob9nsXJfvhExSzrk1BenOPRABTU7RwY2u1if/zhzKKunJoG7nJCa
ox51X6jxtQrzisQ9NKNO4xzgbUGHezNK4/DjoiFxFlteavmNqxc0chScKHbTCAHlSEMTVkAuXLFq
A8WU943oeultOF0vnjX67GSURVgZlxJzdY5gqoljhnlkkOcXPODHCcaspSKkQf+0ZZkXLqldWyA0
zSox0groyTihNnZMdrzUMNvPfLtOIe6ZzPDanlTdfxGd6bWkCKmtgURl2tfOoRTD/ZlBQHeNkCab
zYaynxdC7w5TXwGkxfjEoq7aCGqf9DBWeMYjGzf9F44NrtUNRL4eywc1w1u9d/iP0wTTshuqXnDO
w/E5gNE8GNIA23Emsi2QU08TOmX4BEWBAxWVQ2U6aRJoKxoSkSNyyYy6GZoc6NwQ5r5sdlywTjd+
rtn3XRLT+ySE02fC8/+0cGj14AiHKRUc1YzRKnJ5RhUHQEclaM2d7Uxi1w49Rws3l/BOs/W2mQEQ
hLO6PxRCH3bMyAVFTLA8MdGKbRkgqjiMQeGgxwmEiTQEaIp8DTfwCUk6deelsJ/DNkJy0uw3T94I
zdY3BOIeLnEc/Vs/uXVjzHT5Ns30itFrscT7uXIzVwB/Amn8pLpGwOY40Zr/u0n9TCH+Uge9cIth
QtIWnyAJK6Rk5hqw+EKUcmuLLIMHN56FvJ5ied+dnHzUuRulqrqQmKFMYUO3forOC0rVA466JbWJ
4ggSVnrGxYWhWkSRKP97OexL7y1gZEme+mz42HXimFiGcfM0YxWB23ZWHuzHucb/O15mMZZZg5wM
YOEnrlj5BXwLGuErL4ECCQF2XGXqtrWr/4opEh2qOi8qGgBOoxyHyOP5t9qMnokRunHmUVv/QJAi
CbcTFyPgeMGv9ysk2OL5RxR0zbmP0BOo0yKPrLhdC8+4R9pnSUc8qCecVQRpMDmYFpjy4IxQKcli
kYlYK0Y6KE+3PIXwlLzqATiDukA9CDDbQ2xD9sjgGaJIXPPSmj+8DgEDkxmq5g5ys8lvWKTrWelo
wbMrgHTztOPtAxoogyvnkUtsuY5JPEwomqhrPD4vTcH4SoT9iWwcnLL9qfkg3RshaLawHnmAC5ye
4XDz4khfIDAYhLwr6yauSgnaufsJ0B5ZpjNg8LnGEyiTHzT0dEHPdhh/L7c4L1y5mqI39rrqFI9Q
o5yXFZA+xR16cOSz7ON7YRguB1caqMPxsrf+mxyWcdSn4CnlJOuNds97zBJekadoJYROLzta3bV8
/fw8adRzKWUIkiYnthm1iKfxwvi8z5nKup2u794/Efm338vGewLXrTwzY2/j96M6DwLxFu898tJk
vmam+Y4VNdo2wh7C2+P6/C1PnHyfJsR5gL5yg39ledz5YEWimWxjBXXi9sb9AqRStd2KFnIHAYxu
x/8jw4w+Bhk+LQNRODqtDZw9ENTroFY1e1jQD4SJQ5KJ4/xbU64ndycy+rXiqut+FUbZihDLitCK
1x7vWzTGuQurOXo74EwVPL0LBjeIQnAqmbEs82RYlcI1kjDVIVsxmo4dzakIjN9kVsyjMfi67H7b
zTP6wo3o08U477FRocAPOFpFhqt6s4HGqbjNvDPGJmh2ale5IjEomgZwxBOncgUiVWyh2NFNe6+k
HfiyOj5qhmFL+HRZVBCk7d/Ro8BNUfD5f1X2pm7mmXiiF2+9a2R3XOTqTf2wG4poaccbI0UW5J5l
nLU1ImK737w/DkA73GZUIYciKel/hLZuG0KabtVp6kzyhwaKz5wpxnVXjfzRwXESk+DPr45DpprN
bhaQrMGKiP8SFc2yhRF85BUJcrj2FJJOI7JSWaWlmrX1dh8/u4LHfCW7UJiLeayJ8bLhaNMFTY+j
aids2OPDoKJ6Jyh/WMrvT/jeDoBHFCZb6w+8XRcckBhCDyfTaxEyo15ExfxCsN8RnrJqmRG0/Gpb
h3HcKQdCA2eH2CrXgR7T3S1zlTktRAyfcklAtsMhrrZLEaS2+v18OhqXgx3btLJPyMN7uxInngmQ
yVRzd0hjib3bEs+f0u5Hf2AUA98kVrZyVcg17ORe3WBa7gFe6qDhXsFGV03blSzfXA9U8CIBvMAw
rJmtkbLDQnwXjwZW0l01uWrhI/FJpSWGy8ySps5aATw2avc4Sibvl2mfEowEJMKIb7WjnuXawaCB
3VRhjey1fMP31oIBMJ9wc+rN/a5baAwrctQVtAQ1viVLB/6X47H9y8Nlg1PRAfYtRs4qbiN4IBb+
xKYBsX+QgxtJFOayyj/6/3UZiPYB6pjOPrMaf5NBiwDWa0gBT7NUvvioJ2VetvcmUvcv/IvPi3Lo
oFaaYAfBlxVF7pXlRnTiBOpgD4utp1mMuhR3yXeOFoHx6Bgztvy8Gcobhqs/x7y9De58U7+LN5rd
rqkVfezjrzzClDNgGWTeOmPatsUYEWpLFVTGJFUEnMGmEJKmZEgrsJI2ZulWRSnJQOhsJnamVqPs
vJU8YZAI5x8QPCJjFitONFrUGL5BE2v+ZPRf35qBn8RFAhKkaF6OiZoXohA2bmbe5lwOph5NSBqH
wuaHIX4KYwrofyYe61BVwdWIz78jlu7Pb3U9zBL0MHqsXrcVGiEYdgWjGj+yEz1viHy/aGmzN8cN
WUieX8KhDI4/5fE/kZNcRcdO7Y9DH3FEuOBLIiMcBN6rcNxBu59/n14LJiy8DsyomOiFD8ANY9Ck
Oq4YiPfKUVau2tG93Sthl7aeejvkVZl2qNCKVxdgZgADvKNqebMaYn9GTizXtlcdtLkgb+iPCc/u
CYTCQZNKXQ/Pttyjh6l5lfKUdE68qcO/cv4xgabNB5l3orDAr/AY+26V4zC32qUrEE8A2V0MReAu
L0RvrDkE7HMGJGuR6C0gBM1KRdneXJ6+R2ZBdiIyobro1u31TCuNJ5XSNDobhX7hxA/yd38SiAxk
cYfJNWalG43cxyt7BYTmLkyS/psKE97zS+obhCzKZfS6Oh0J/X0J/lg3nUnI1M0lQV43lb6vXpLv
M09ns5OeHtdo9nmjs3tLIcfurZbUygfdNXiAQjfLNetYXZmFB2fFT3GSIhMc+R+gb6ALa2xShVeg
wmIpwFqhYQVWiqal9T+w3y8vWu7XlD6POD3pBcvY+szVP7qj62VJF34/niOaybMn8JJEkxafc4HP
pnmpdXqIKSg+09RSG9SMDEoFkODJnMa6tObI+gw6AHLZbxrXdFQFr4vYkHFs4e4m2eC2m2PG7Ywb
BdDjPOKyZB/uUu8UE+b0MFvnKewlD1oAtO0lO+cQHSfEgKvgR2KzgYPwjRbcHqERjrobgJUV8vg+
TIhYzUuZm2N6aLyXB3+Vh6kyC1cr7UETvFjmOoftNfIE5CBVhcicurbU2iNO7mgd2WkAC+WmW+j/
0NWi2Z4y4qYk9i/HalCa5POPQ7DrcG8aw9l6TJbWOg384ACa/vy6xQAx6jMpVh8TBfxWfwHwX6uF
T7JF6TySnXeSQFQduwQfZ52+Tl1nmMW2DL5nW9AEgWL8UpnfBWqsHsCHoLt9cvpe39FlagqFEFbN
MVCUORLvOK+uq/T/u8kAR3/qYPpQVchoRZr0kxMO+OJT9RzMIFwsSJ4tvrC9wuBbQYCi5EaqVpFR
GL5WGdPI1yk4VS+GiUcq0FVXVeDQYwqyw+znBPvn6S9NJ1IEyTy7wA7oLFurQTl3Tox/L0B5Aw36
9RKFVil/TZYp0OUt9BXD0MNrMH5nxyweEtFl0vLcKxNjVkXm4TUGKknXRJIzTaQADbP+5ojNFWFP
CwORkX27ye2IWvhTp/40y0UGgBWJsGMhMAEqXRKWgCCkjiBQ+mh2/dKWehR9/qPLg9cxlttAh+YG
CvF8bZva5jb0OfT4cabyT/YFEZiojPVWb10Setd1naMyvGr54/hVqOWwMyi8XqRjEgBJMNJQzT2k
Cgr8ACYt21JXV547oByarxBM3PdgI+eFsYXxjoi2Nzk+E39F43TvHJ7qGqlpwMh7naa8VYZJstGn
0pD6Rw1FF9AJ1ZCDux+KjSRZzSN3mMWRfe8n+oJbXq+ydmgovNgQOXRH0dBHVm9pG7sGL/iqR1sC
kaekgSj16qF95LovOVFOkr5L7AWAzP3JWJVytKbBqgWU7/qrhvu6WJ0lnO7UR5RlUjDfo1yw4t20
dQOiaRTNYNGRBTKjiInyTqWd0a0U0vw1Lu4AmMIW8vtC3DGMGBo8vgwelspcaZtJ9GmL+nIlIYPM
aADh4hlw3AcswQD3fgCjPepfMgGQVcMxtGdvF/zrdzG5NRw8XG5KmCu/ymxwd9XoVzYiQoe1lan9
h3g5TQt1ep4/88XgEci9TaHcuAvVc5YN047ao599VWjSyp9e8hCjUabtriD9ABGzEf+rM/z961nF
6K/JJ7UMY2DxfB3VElGrkrfK0H4b8AIrVTRdT6ZhD0lZZiB191KO9xbS5Xpz4UZcz4uJhsGp1Ijn
lGuwwtBAzRUPd3JMlxdRoJo+Kn803c75YOLKRKtXtUw8eQmDW0ygo/KulE6DwqILNh3HU7bf46RU
2p6X4lDFfmqGpaO2qIgHYKIp+3LDmdbUb6yJ8XPykwDzfK8rlj+O5o8pND1bG7ht2k/6f3szLweO
jow7RxpKxlWU3uoq3r+JMn1WOu64IH6IRB7czNsWo1rAGrjTOUq0MyFGFZKzkQ65kRqMS6ANmXtY
8bA2I+Bq93ncYzBlRc1JU/mnExeaxY629uZEjDHmumfCmHI+S1voGDDK+9ryDZD8mYqKKyovJVTz
IuORQJ8T15x7+huCi/7qex+/T3UUra+Zx4DHaDkuKy9pK8LSqxpDdZ1hUDSG7VMxdHFRVw5oL8zJ
EAyrL2RwHUcziwnmVTJBlv2rFV/NMhqHsFO1bTiAJj69F7MUcQ/sYlpM2SJVcGC3VUNOdVwufe29
PKlVgw+xwCC/Hs3lYopGTtdXOWwD7E9RjXOl9fPXDq2d4RiBDr9AckvJDdnXgazlrKcMdiT/4uAQ
dioA8C1wVc4/bwv8BJDYA0NoponbiRlIfFkn/BZt/xLyuoD4YIZmnq7LLN6y20zyyAI3QH1QWeTf
TzugzJfWrLmVkikBm7g2GZw5tb/Rprz4k+UygF6VM/tDuSGtzQb0IquojNgVq58livEaamFfVNAn
s/r0u/TqkNTspHNAGdvuPIB+wY1qiP6/HS200bqskMJMGcWKMSRZwg//GTL7ftDUOVD3BReaqhRX
1+jadszbCv26df35gXashpz71DYb6E+JE9hNtZ56ObxJ+ih9ITaVotbCZjT+Jy2/LVniYU9qIzx0
FZHQxjvPkPCSg8CpjOM5qbKWZAtS+A6aP6G6L3167PRRpBbG7ng/qOSoTgZX8OtfAFpVaxVW7F7l
TvCkKIStToWDY38RYv0XHDwiNH6VfG1cKtqTtnxKdELyr3Kn/j44oh8j6PwKf/bBlLva8BGlIMds
QfvLdOCtvb1RQvNDVBQIMqYGpYB9gOYS5XQ+uU7nbR1LRrn1gzVNC6QgaJdYeb2NdtdaZ19ROe6E
O7Fc+/27I5DoF7MpcBUY5IGCgRJiMcHe8NaLpLvFe5Ot9HscIxLfUNdTd50QTQYm6E7d4mECS3FL
8TTTBVMBq8KE34U+kxOpOs8AZ2nngtN/WIQelY/trVzav6gQWQYnj8GFnO8ggaGOL6/ZYL9ji0rx
jwks2ANxKHbm2lN8y27G86pm8DCDHvP82h6yGXogEtQNW5YzLsRnVzsY1JMiO9EIcm7wzJuhVGX7
SDr6ZwOheGPGzfwyaju1/Vj6jIBbNF6JRncvOWmaHFwlcK5Uw7oI7KeSrYajdrVe1Gfdv39WBp6q
t9FjqTtDV0RonLKqjQIRhAe7TU4Ndcp9hTmSRGZWcCaRD8GExrQj8FM7us+8NB/6d1ofm/MeoVV6
kvQl0ieBzvjhxHhG6KDE/0kZAbKSIlzkAbZKalugisndkNWOYEyTLv2wKzMGE48HC17nXMmSKUe0
QfhgGUraJnF4V4STbLDcGmZL7wxK9Uql4chbHb4rAmPrMIqbdEMh+jncV7jaAc5+NFc4fCQ8PMri
J8daPNBtZ6z9ysdU3/NReYHeFak7IGsXADKUi75zw8kwdxxi0Vniztqyr2QqTC/T4RVdhiUGeh5x
711VpCu3ICVtGojBgBdYBfoFm3Q2PuN7XcHki/t+MNulP6XiuK8cwyMwOmIGCkeQlV+3PH6rw+yE
IrJYjl3fW9PD5wZuAHxFxusxHjJZJNDqZKnLl0ajCXN5LjaEH0cd3FIswpDhjagrZVtqhwhvJCMg
g0y1pEo/aj4Tp8FgwEpua4Y/gHTcoaB992lJWNNFfhOQ2m6jdEV8wA0ZJvslvh+ty9hVUY8Ct07L
Jq5V4TmjhqEkvdFLNQpkMH/H9k6uhJqischkyV6f4ClGPUIumR/zKouZPRErdNp/kSuR2u4YfITQ
WCDRyiACr9nfsL+/Eub+OvmTwlkkDGitBOYkS4MJX8F2HNgxIRvBCEj0HLcbU3M2tSwoROrm+JFe
9WCItvOkCnHzg0XdoPGVkP9krBBZ0TmN68sYx0P2KWjjc3fydnUl/nYgTZp8NYcbIiYRgRctxz76
09N82LrAlK9doDFwCaajXGuk39Igd1bJ9K734vjJKUBgWaAVNCuXSo9mIKsziw2TmGQ9wf5BGzlX
b+O367xNOylKXJPSnT+v0LfM+/TZM5lEru2WP0MFEtZ/YoOQqdmJ8vb0uQjG6+YwvNPfLqrPoND9
Vt7SNFyQHgJBFV7D7jiLO4R2TMp5EkPTC0MjukmV96uUQv3fWLLcswzD9KiDA2JiQHmMVwTp4f1O
X3/rrKzItTiSDEU5OLZQhb12/O1Fo07Cfw03dfxqsrXBOJ/C8sJVBqdCGokFhgVutX2W8hOSBt/p
5GwIWu6n1CLvd8z2HFZv35BwIxyubWOCo8IZ7JK4Ob6L1WS0nxOJFXpVsM/bIws9UtkeljJwjpdN
A02iO5Xe4FGyHnKCbQ4yTRwlFmZEai2y7f78p1+S3OEZYLP8609QLtZb6k/C8OyxFkAQc9q2n1GW
kd8ckDUpqARa6xt/o7pvbId6hdA62gRS+NfV99e1ZWOBByq4HeJmgmaMP+MeVh7ZglS4hlNiOPg1
+q46iU5juxFSzrZW2UgVzFoInA5OE8JtGd4365FWm5hqUDjoSd97MKuzYw+styvOERyv/b0CdIdh
41AVdYeHCuk1K6eydVS2wyDJBIzY8kr/x46fUYPgXXNKk7256TciPD++c5r772rAqz62vg8ZHzEe
VHB6iepzT3EKqNbky9RQIHO0qBksnAvqArqysbYxiuugC7fwuixPCBrHT5LqZFVa28+HV/PKCyq/
7Y/Znp1ex2Kmp8pt+raq3GPGY4p2y69n0FMeLchD2qR3AE7HrDR01jyZrFZzGQP/5TD9BUzzrKOe
aQR2bLF/g0RxGdLy9MNRB1tyt3Fx2Inq5l5AVu+eUm0LcSyh2Qr2su9bGZISne4LhuCbSV3LEKrx
P73OMRKj9C4FyfkpR6yZswRYVBLdoQQPXjKM6LayHw7CXypCksMCTb0UJ6VZ497yIHrETF9QFB4L
d+gf4XbKAq1sD7nWbqhxSAgiPWUpUURKBZjxvb/LGf/XFOJId+VG81PD9ijyYAKt4nEhkfu8awbu
iCe5Ibtckn/Dxde4oBJCyvN4phzO12s3VjkboElB+lXr+OyKEcHXspyaYj5QAC4QuZVKjI+kEIfF
dDpsJv+GBD10vqagUQPpPaTJ+8QiUoeM6PPrV9m1wj3aRIGXlMp3XU5gjE+DQknxFq3HMCDQWF54
z4RPM7ZfZ1ZvyhoOe6P8gRx6i8pmh4cXWlNVmZncATdLDyAwSE5fVxedRi7m5Qf/6i9K0n4WOJ/d
qNbX76AlRIyBuu7VFZJXM51gWEhy9a6zMORI3DOx8i0qTRtgp8SjtzLAhNJ83B5AxHoIuQ/PdDly
Amjm+H9PF1m1MzqCWjpTrveInfiT8i1KMcU8+M4sq8bKULqhTgpvr6nUyfMK4u4UjbFm96//ECOJ
3p1fR8P8Y8IxGaurzu8PDyTcnARMMBh66yW8ckMXTinyiHVyhV076Xdmmt4KUxuI0pY7h6QHyIMh
BIKKDwpe+H8wsMertDCNem4809DphxNdBTht1pkiQ0/MI3x1i6YivTj3vmGRWst9/jPn/i3b48Ux
G3Uziy+KCcXr+2eibOMjfKMrusg27EGnrFlVlkH71wv/gbEkhRmlg04Kh86IYJVAEqNrCwyqS3Zb
HVASTX+zJkyW+cG55XnyHilGgwUuWu4qHro9e57Qaw3mNtG+MLymWD7DkQPj20HIiT5l0hDtu1TQ
fFVxaoStFL1gBx5ZJosofNUJNZg4w+bUnhnyPHrJ9kS/PbeRxN1BYIiUZyCyEqH2EyhkCId7N/YX
Zo/qCIWjyahc4ecSZrcmXmFtxW3a8gX2RCqlQPuyAMCDWz7hacUEGGqMPv9Lj17KZUjNp9uDRX+P
hXIPkrc4DR3z7WQ9xJ8p0yUli2o45j3DbJgipf5GTo/FvAwgK9Q3y6xGYslTw3KpxAM3phBrMUrU
r6qj437wJQgoj+lfL+7mnsPcy6btWXs2FmAS5z7FkrDRtiQHNeoVVN3uBWcSqNh1bzr3MhiUqgZw
5W2I5Edp9QVgt0yVZvmJe72d2hPlj46Bv2SB/udopIQq6nBXq8M68WJrs/MFHSapnX79m+VoGQbS
RFbJoXshZzIG3lZR1FB1m46Ynz92qI/DBAER2qUbntx+HKMWp33gUwwc5aw8IElTfqp8WpWDzkHd
x5kqu1TnVjqPx9eJ9IFvomS1YzhBKFDrsjgoyD6vvHNPqoFQ6/ADeRVb4FvFz4CLW+/Lujt5/nud
eIUdI7cHf53tPnRm7okttnjaACYx58U5DHGzeg2GdZ+RSHApEBbzaVEhvVtSy9lXn/IH+Nk+R5ii
085Se62W4ncI+A0UWEVmM7WCe2Ya8az60SW6xbllEp5XwtL2ua8LOMuYZk1JDk1OjoDd837NvoMa
hsXvyckUu7uji89zcHrJBX6IxwH51xM0bZAtUtbdtoBioaG4haUYOZxLc9zqp0faDdc5DuYUgj0N
73ht6W/po2HNsZQUdbHtSC66JbKfN80k1qwPfv2xfbkIui/dejyG47DX0yTQn3V89PY/2H+qfS7a
ERNO/g01IFkTOWmxiZd58OuUBdglDDdES+Kg7hWUY6yHfFd/GDbtowtl0qI3w+BoISPn0/ZfXuoi
iSmHTTaQR/gu3xm5ZBtIQ73veQuv3PPqteMCRwsGHlNFq4WRM9wFNi5INoCgWNX+FC0FQxymwfsa
zb+cgkF5kxqqMm2gDnuFRzspSdo9/f37jYLd6S4BluHV4Ihy593tZKkZYGZJ5yvijj3eEY4dXdRU
H03Ua3u8LDfNQBy+0bic94LYZnWDpsMVTzAJXP5dMwdwb4GkSSIiwLWvtaphm0uourG7UkaRpisF
oF1F/4SjY9+Wbro+e2DdLUfbxQwXRhfHsO195EFkh/gefHYRVKJDaPhRVof2i/DOGIm0lZHkNRE8
1vbQIMSsj+NEKYWilGxQRhGDB6fjl/0FTSuetzTV76al/ItcKLemxkjOUzXmMTV+MT4HfhRTedaX
K6AracxyeEm4xcz/97aB7VeRK5gzEQGfeWkB5Nkr8XQTftzJWFXSgy3MM5E4kbbgGdLZMIXzpWSF
69tkNLn8BNNZWd87hOsIayE/NS4piqv0kFaNtrspgLwjk3BsJ5sCJ0w8FjZ11b0GCEa8Nh/cwIUX
vGtAsQ++rNPMlE8lbF3RoIUJfr0sblfE8jSqYKDw0PcN6b1EbJ7qzrSFIxEvH2H6sede7sjfsufd
kUUWQ3XzQvuZJFoQ7HOksR47dZn0UmVW/+NJ/I0aF+fF7y0k5oa4ZI4zOjiDWUzidCI5dHgGz2Nk
zwY6KLLRhQG4tNxGl9mOEtXLtKdFy0UQN0+U7SDoAFIfkPOytbBIwEE65snmV8Tho4z9zUycTFyF
9mtGjcC8uN94SpIO4FbGiBDeZFO+MZvxnWihPugcaVeO9U47GQInrWj4RNR1TX8b5ClMvZd23cUw
7sDHNgEwsjT/foMCBunRoVccfY+9rgtSjv3noiGUv887t036jeRT7weZ0i44Li6XmcllCfu6wXSh
30WnqFiD3pWstU7QoWVkuvc0nKFpp/0jqUkV1QLQyMrST95FJ8zLV36f1cvbt9O2cQycPQXJtfqN
8HG2ixNNFikVUDK5Lr3t5+da4vACWcg0HVxgGFe1qFP6MJ3YMJt6ZrZu1UlynghVUv1SyZLJS/QK
SrHYRjPGtYcRdtjBaW6ekkxTu2tsJ0agjk/cyMIjUq+BJ2UI14/g6fHJ04UqFh7/6bJzryx5r1IE
WSun4O2IlUTd8ysmc/NpYJ1dMT+FUCuysZpYnJVba0LXgB9940Zgy5uN9laXkD14z+5qPkDBGQ3V
UmkvnfRhd7pTJ+z+oDAyg28M/NXp6oQFav7240mlju/34vuJL0xjUUamaTMTW2tg4kUYJtvrW87I
L8HeazzNN2wdF4C3sJ7nBMU5hFxm+Sj88hIrNsy1FKSsgxFNebG16UCdx7DI8tCvVOEMZoIqtPsl
yM5V3hDpmvMlFZsAQmMXUil2AUaAgaMjGNbXEobKQhS9S5Z26H2eHuf/4JKdZZwwsvVrc4JuiD9P
TP3WYchqlYH1uYKR2jGnw7g2pedl3Y1fJuGBmf8nSP1kTVM+P8HJxhuoIBjKfU6nZac2get9C/Uw
EyEFVyFaI5gjcMHhk0S6LjX8YQZU40pa5btbo2de28g6wPplsLM2nmeIWzEeE4q6zNtuqbRuJrB5
B7pE/i8Mw+XoRQQS6tHoZkM85iV6FJ/XpYMUNIncTmtdoXMel8XlgcUiIb1WSpc5PLdlib5/fPKT
oWmFuodI7fiXbiS7X1Ef2Vd60CMxWhJtr41s6PbxdKctt7DcjO8eclpgE6Z78niE7W7B5PTyuFdO
ues9W49iXZjOs9HCe6vs6SCnmwBhjl+lYGK6ILefg2ry80tSIGn+67UHvznAOCumHVemQoGcHVMD
o6S8d0ObLick9glNycoGyRZAm6hXZSbxIYE8EkJ9EWFLoGst2XDnOTVAEtyZGY4xczAPxG7mNz+q
a4pfgrWsQjxu65LzHnijdRZe3h8vREWXOgZHUE+5+dru9O4IKabnh+9NtYJTr/azE5Q5Uq4l2QML
VAE0hOi6BjFvLCRVz6M+vVH69ZwR1VKPEo3iiLAAVs0lOhVsYksft3fRK1Qt8BNd+BjoqHsk7Rww
eHn3QHSn6UDYx9c3LHxzOHpEcR63PCRYQlI2B1gmdFlvYaBOhE6OhzDEYxGDE8CTsLKXM1DLBrlw
E3KPbc38rAjWPBXRrW91BScKRODwEajZey1sGAjAybTCunPT8oD5pFZPUhIYTbAWGv/JjDGLYi5V
zG+n1cu40XUFgcvvBgtcWK4hoybYIWJI9WAt13h8kHW9WQ8RdPpIkx3nwro1G1mCitBq9DH3WGPb
/8qLOJAxoTYXzw0ValyeDjEM6AospFTxGvMYXd9iIGzuwcop64o1AqgOE48Ce0RfwkpT3dq2AEZd
qR8Rv5Xn2TtTMKvyvPlmnA+ceiIqyUXAHLTJ5N3JTE+hrUpadXIP77iwiLNPea5CmK5gZy56OD+2
xCrWu/mZmc1yMeduSnPJ16R4hMi5tfDPCH0mG00COHVA8bfjEEWQgoHAUZQ3FPwl8W1RgP3YgTMx
HDF1PLAIskmQuhqVlHtO9manOz/6Qst0Brx2I8LyuweEpRkCu+3DRYEl4XZVXok0BWkKrTQPPakv
PUGJk9LIM888RlzW1i7KHXkzUs54gujoHfr6/t/TH4PQS2/LE1cD/M7o3kR7Lkw71ZpaHV75pPgE
gD6ZJ4czswgRscMeRF/bVlL4GZyK1Q8ByrKRhDYH/JQMKnSaJIHjCqyu6khCYiFM9dWcLnYppUZe
bJFFh/oljsn+E/vjJizmqaBE88EblazqOa17TowMbxadT+9gm4toSSZh+saKJQcaRmkpgfNrqzg/
KbNu/aoDG5tgJKddf5SAevjWXT4XUGn/Iw+7LECGHCY0dJhf+jlrReSS/OI2zgjFODuyd42OdFpq
eAlb0MAx/z4y7WKC/zijj5S5AR2uqXYQQW+TTu2jjuV3RieHHUKJ6LR8wmo2SpKtvUopTqf6DOok
VRlSGePEPgFyYqD6LP3vrPl0RvGff/WutykSSzv3gI7OihLM+hugxm9j+J3FsNUQNqYn1umJuFZf
rTxbLKkmJD+uCt9aExmylrwOnsOQm5KlScgT7Om99EQFDXQNKy5bLHUd/UXDjZGYz3yfS5QgtQSS
ETocG7uSxK7xprE2a5QnNfe71EPZCpccSaboQ54omSNTGPhnC9LoydTlrssheIzzNUNZu34Co4p/
Vq9yR4cy/krXT5lakcSUdjlV5amtEsKRLn8XlN8LHwvfyeieCK6EhJ/dFt+bBTwgSTOqBWXapmkN
30ZfZfXnAZdS5FymVBL9XyMtb4v3d54AaoeRyZJ7Eg+abIWtyDp7oXoNOKHqa1EvOpqFAigGNXJX
XvTT68JiIa6VN1bT/s7XO1q0f8zuF//RmXvSXTdkYoX4uTIlEufwjyQaGPMKEzVf6IAVvvqyT667
1tNp4PYwiV8WG5IcYpDPr+Wzqke9MV3fTFsHHTc8z/ZzcsxQRiYTETmWqFWBK/PpTg+9HS/JRaN2
Y4UqO3VORdkgTRt4r3mSEOZSvsG6MkhjJmt+10b7b1QZW594mg7BgNz/v+3b0Qam+1AK+rh7YHQm
JE9YDrFcvps3/MpUyKDyRoARIPjNwb/+ilTeRK0nr76HF4WOw1BSuPZiE+EWHDC1TLjBkXGijD0P
IvWkQ2nhPuYwnZDm8DTj0m+/sJV3BOvrWWAGyZXe9gZvl2flsILnMl6B8yv/q9ByVIOsUoHgz8gE
E40VQ+j23g1Qmz+dDaVR838UULWIk/OcOOC+bmBhmK0urCQyHdL0L+WXbz2+AYo64H4ee4CdtjoG
d9d9Yr56bpE+gqI1R5jhaI9SqbFWT6fnxjPJ/3zaLkHr1bQH5xolI5LlBJlGq23GtPfgq3hpJ53R
dwDnA1wMg3l523xKzjp1l76ZDy18Mhm8i2fw0sNdDHsDklIqh8Clv74VEaHY96cRYLuUpcDHqWfN
VF4ljb4Y8t33rKBN3FaNM9cCLc5B9EJWz7ddJKsG2a00RO4aWXx3JOdqzWJ+toKEAiIdqbaxtyvt
vtk0UMq7RBFgg/jNp2AW+Tr2T94ZJ10AOsr7j5qE1eyRcFpjz28+C5XNRygs8MJJBcYlde+Zy0av
sUgtYPR7Ikt3PxgIHprAByjXJ1ISt5pc09WBdW7A4sSt9gUKWc5mDkjRfVMtGcSligj1ofqZPj1V
IH2u71dx5ZPUURoDglhTjziqCw0DVq7Q4EWdkQpfaaxAus7jqF3sUl/VaPrAjoB1riyGhNXLkFFw
DnCQVzfyzh9DQ2xG6MYvfBfdcO7Kij3l3ZRpaV7RZ6xdkyIOIbddW9BFadDiJ0/9TjHb7sFCjRaj
kX+uniR/M0hGdMnI49fwFAsVMKIQUWx1YNV3BBuzlcHzIuPJ/vlvmYJPod7xID5eNNcRtmHyMJ5W
Utsmp6nbyBY6YFLaKulkzUyqrYHMtuV9NcDfsWSy+S3kLJwyFJ3rQmyPp5O53+nDrDjvkRghJw5d
do/csNE3y5n86L4w+Gl6zyiqAweoQVn7Skhc4q+vybuG99MdPduFoECO0Oyqj5R1zi0pxMMRM122
H+ZKWMtgdqm8l8sevfktRKLNnj4fBkBdZ7WudRSiQlTNjpJX4m+FPFgbeqTvezTERQ5Divqj8qKL
RhDUvgM6pszF1PVvraDbf2KfrcUE4jjlzn2sfrXtZ+X4HjDybumeZTY1SvPBhPwNd9IZAjCVmzgl
8x6hnGVU/kQ2QIKaid7KgQsnto9ewNiSjLJUoAp8E5FYp6dij9P3i0oyeBrvrAcH6ng3tIRCUXAw
T8VzZ/dDoOPg0joZVJO1j1gAeFjdpAzm4GndUfkIUs01LndZnicZ4Gd9W/w+8iUOrSujgy5fUiJf
vnL8DmDQM3uPF4JraA92Yr2J7r8N9PWzxC87XxYI/y/iEko40sRWZq6X3WUkFG0DaQEu15P7yfZK
AuR2XSbenfP48CqsHu9i8ORXbFLFM83swTfxZA0nc2x0BoY+qBoULbqFYoYq0mOK1DyEwtoMJdUt
ku2AuuWHQUUIn38RRxTlHaI2EqHxh1/CduL/aYOcfkX10ohGMFZ2CbexiLE8rWU8HIExvTd5eQ8J
J1rtGJTg7CqFdoflHutqW1AZi9s31flt/aEeWL1Eqj/a5xGubleY0jL4DQuIFf8Opn6WyTpoWzD3
9mfC0DRYoUGrUQx4JqnF2bNrjEvl4BVQDkoD4DKbXrxeG2VDtnD+A5EBzA5hPWaI8+cO/hA0rqxJ
P5Pcex6WNquC53zMIAwSIaV55vPbULdlSVMO9yV3habhEXmLX1ZXmW0w+CHlb3eJ8kS1c7eGVOCd
8qp2ayIxlNDQGdZN6Zudt1ljFJ/G2ECX2xji7anlI/vATHAXT0BXi3Iu+iBaWEqNzzqZJAAHD3fN
qP8/V+Z44d6YO5fVc/2R2XM4kCrnZVXjZi7dlos0UdrGNMOH1JxvFwXQGny4OcaGw095CK6P+zVA
HtD88i8n/Lrs3TMcuYIwIIQZu3RlfUjCyHJ03uOl7Ii6XxcMfZaV9KHP41/OWZ93zq7YYoPb5LuG
dE8DR9laWskplpFDQs222be7RgWNEPphMNydwgsPsyiDp+BbUsfH7kmkfo9RDJGpBVJw74G1g5wd
odvCCLYf67qSntuDpBbiQttqU3ny6sSos+p8LzcCw0qU5EVgvX5oMxK68Wv2xzm/UgPXTtSWu0Kk
yvxdxdf/OxkQLev2ZmYVqr5RkTU+wvCbZXSwCGhiUVTlMsG4k+OXvVEq5rSAYkhKau5pWLDJtsip
PhwGCQnI6sd4wjqwYd9ZOuTjJj/pUkBWxtDEkKNtcGlzl511XBAHG9I4ERk8B+/ss8V2kSb5en3t
t0MPkpyJOYZLobicHDBV3Y3ZOLtoHT14FYcE4B+g5WtvAOgB7a8+VV6V+tYP8MRaRiXBLTOtNmGH
81aj3ioYc1pfVwyB7ajWcgyVSYhNchplV17ybfZIdJFikNURX2UzIcev3/JhxLPxVSygeVOjI5g7
UGnFErbJJ19WAAX1uUx8+UPSCUeN+GnWVV4auBzP1Hhl2bPzVdOkdmoB6fRcKVD1dKlcIr/hrIES
ZKhB+kGIJWL2HeSxv8abXmXKA1qa0EsGZp/FgrSD3UZAC5a2Kvs/cZmyDFQYecGcyIKoGijcyCSy
Y/dY6I2gFtVEL2ga8X2ka3euXbmkpQp34f00QyYTizwIxdohvI/G+8YI6OttEBSpQiqWxCIu5SVP
/PVQMhOGlTjnmkQWBlNswlEdbfWyx1ZKZ+CPoez3ig+pDRVJsdytF5cMXmzSTYMDVHlHIO8QuIEe
yDomx+qMjpr9/43QjKxDqavQ2/xgamWdvJf3Ny7raCjwP9+aEQ2WoJYbTft5XQKLbeyWAeaaERty
t+dkLQFag7BWD2cY3XQhjds3Jv5zl2lj84fHAOoXJ0LV+xA8kWSvOIwVEuGvjIveY2ZiDW7uY8OS
VI6IqM6J2fpY2+3xx8yibGIi3u5YIVkVt/UHn8yrciJy3pyfSyA2McfCLLyuGF0EqyDKVvQeWGXe
FWLDt+A+VLshguvQC8t3uw5IdSvbnBw4GMo2TuievvuGDAMpYjdlYCbMMY1BzbAiW3qxkupkA8m0
9bJBQJXGoMopVK82kKNywZeHQjYLx8u1C8e30y3f0bg6tQeg6EAmD/IWg+Gy9pSG1AdNR0EnVC3U
EDv58w+Xc8Boem/Hz0PQWMMh5fK5kxLx3ZRJcdMf77dDiqVK5YAAJvJUfwQY9C6tVYPvIHwLrlEy
BBUJmxMYbZQPlDV877i24G01eeI1wON9VKpK7LKUjwOy1v5JNu4igovI0FCrMYAEirGKIkC575Fk
fRbnq2tSW080qgyPwM1OxMtZA0utbXY6BUIhvIILV1TS7Y6BKO43GNjGOKxbobFZ1E/A5bCmJcSC
KIHZH1FQx1ed/lbb0UbMXPPDyz/BjCJ+4WgXuHKW69Shv3Sem0pVkEGHVes0xZJsqkAo+RrBmYEy
IMaGemUTg5FgsZL60OkMAxVU9KZ4RaTth06ST0M8zWRb/T6ub1T0IT3tjT6unc5PiC0D4Mpx3vog
PO2LG+uWawGqvSpusA7vV9qFUQpSWEBwcLi5gAWhJPtxkD5BQOIrnrqvUKQyxlrTWtsS44hmtrqo
CJqMLYEDT85mOhD1iWCn2Ti+EFqDyl8Au3VCjHHcl+cCg8N8m1Ryfb5esJ09KK0Buu3oh34ilQ9F
my/mRGwAMWG2jzjys6WsQlaOLyuRZSwKSwmbQCemKnOGjRhatKgM87OrdkmQ9P2kHVv02F47QBtz
uzbwWky5PJx9/UDeHlgnQE7CFtLekd4lPU674P2786sy7ovqVCP/WrshD/gCywKawaAbX/1PLHSa
Eb0iN+7Km16qqvqq5W+bq+W7me5rpNU4rSoGaXGGa35UCdeFmV3rwIyv4QwRkuiUhvLOM3UgndWQ
/2g07m6fwYs4NhCpFkrj2QfQ1gNQ+1PEVQj+V02KY5xgVSCL6gJucqo6uANq9cbUh4CVAvDFM461
6+FthjRFLvg0bW+vbYCaMGepgSYKB2S++qeG1Tsx/2K0SzIEoegnSdnfurBeYj/QcVdYCk1b1al/
LVHuMKUihvVr4HsTXebg8c5ghSZjk4W5F+HZ1qwZGyMJweWK/e2I/gVsMwUuGo6EXntXNUhwsRvU
xdcMmcbgsEItS6nWo5/GQ03Vr4AniJGGeyEa81UVy80A+sZrCMY4rIL+6UOrQ+vjXE2Fy5cH28Xl
PA3DN7TTsmbAxnPghH2qA338cE6MxI2lJhlo+eEkcJg/AGH2A3IWBNygeVpbv9jgwCAVGz9XsaGn
SU2aiUsbJR6yvVMzRtTwqZr0DvPcbmIZNkyZ5eNwE/m76oVAqP+K8DOgGQ3THHVnkkW1yW+X66If
KogP5o+vYOhkbYO2oTHBgQuaBVngtgHbCJ04iN5YEjhMI5fhhTBf/ouJxU72c9F9r5lMtO8Bzd4D
b83ocOVyaALWdmM4B51Cqk+Y52ydKsYdb9mmbL2A72f21eFA1gbbai3MrhJOVM+MwM9jQopx8Ixo
VWaOCgf/lSQ/sAkZ+8GfRC1o0VxPHwfwtp8WN+O4wgy7bZnZLucusEUPeNEGpCLsKZT/TI1G3SXW
u/PPyj2LBrKStD8m5BlyTEPTZC8e8vuzVa+EN7sPnQ7u3sKizMnjk2V9rloFUXGVg7an4g+2gZ82
GSf0A25sUogILMRTct33zWzJsx35PecJf5ahnVppDqtc58REPZrb9rMd2a6i2kjPwaKlDqA4v2qk
COIiFNyOnymPANgzK4aXsXxzhPQXjq0eh3g6OLBIek5iIIhf7pVTqVKXjIpCDMmPY63BjKC83MzD
0BuMsJG3nseTHwUgglU5tFozYTKmZwmBi7IK+fS09PsOODCY5VXRsK+KEz3n+0tdIndNAUDLivk8
9CTW4o1UelSnIlpsnZV9s+CXKJbmPom6BEa2BNE215xxdBgGAsL878G+NCT3e8nLtj8bakiDAnGE
vOd5SQEOsqRyagyfctSGDHuqw6Vyfe6WN8zFPdNcNMTe0GH7QdrZ1/qMUP9JwUkD9w57+kX0Cn7K
+XIlOtaLOL2A++hOGNHdCmTVh9q8cs7GHARU8Kn4up7Iu5LeVxemTP8U1IY+hN4QIB9mYTfPKsr2
nGog+Cx7mpl3YhEzvN0D+bqjna/2ERpjp7NzrEYAqnVucTRkWo33+F2JrHPIiYFTbWBuiSOh0LjG
4Pym1XwCqvGyxbGjZdUeh9RSgp9j+iV8to/AfsVHK2htDAKUHIRDCcTyEG7dh1trxF4A2KZy43k5
WT5tmO4v/NuYK+3tHMdYkJM7uDqoZ2fY6dv/2WdPq59jzGnNywg6TSgdPnIhIoUkYCHwwNItXpPx
NITisZ/DhuIBslksQ3/qAQUulI34gx84e8uF7lLWSFQMDwObOOu18nM3oeCHvBkH17CB1ouCwi45
ujnNxRbQI4yowtdglgrFJmr6995s3wXEitK2kFgakdE5flk1qzgVNOnvtZfAV65he8WhMBeudBB5
x1dhrCjAZ0uFv4fb0L3nKwEMhx9vsVj1lavlmHjQhwvHih5WuE53EQGPF0XbHJqKzAybge6L7S0c
J/eas2ASZnNdIVBmu27BDWGrTqqtFaMAVhqdj5ung3hzuWJ+OO1LUVUDiRRDBXexYqB49hVkv939
/9bkA3hUT03/IiuhfhHq7xlOexr5jZSSjRy3yrBDCebM6Qfw/8W8OJMjriOm1ueHH34JsvAeWURO
aA17hHPe4C7mWdzwJGttR3Q8/Kkna6f3JJppv2oMaQpAETsWY0K0pm+2+Rls/Ubv8iwnpqkfRc7x
Cd0aoYq+nZUF14MhYApWgDqj5igeeW5eOp8pOVnteAV4N5gNi20CxbpNkMmTRCts8yUk+V/xOXH1
YCh924vulguQPoWSWcJftHuTHxkF1rgxszjrxW7w+cL6SrUQjhWcNzKTtn3d+q0xyqjhDHR3WM2k
i2LDbQvZNEjlk8y8ZNSZLVE9IcftAEuA9hwFh3b0Tryrf9qNjFw7fYIpdTFeXQmrGHOyWNznJuzs
+wU5/FxD8ocZUm8iDL+nhH7A2L4nLo9pruzE7nQryGC1h0SES/2rAmilFPlkKLbwA0qVwmFCTGev
GMXLeGaWav8XBjnSJDR/id1BA6pKvZu85FyDFkj9veySOppxqsn3RZMb4tNLf0jqXo5h7YPXg0Dh
t5tLjmQADfheZhH0W4s35iMxyIc+DcZAbjKl83bSk9D7gQmoYxUR/33PsOz7pvxrX4ov2coeJnGl
UKffVLl5UyYWXCsXRAHoY+dwIDs/ROaqCfZovYlW8nBYdudLwADxSfcv8X8gfsaIZK8FzEXTXece
l8HSi2pGTOf2nJzTvWcFFOVgIw42JqY5+al9FbdSIoQ7YdqixVdvGbYeJYxnrF+lQ3CFCRmS4kzq
q9Ir3xTya2SnhPul9DgJvIoVoEGRTBareZCqRyk3fCLu0xSx9WVOG6DmzPLBcjr+cYdX912eKBKw
oKmmp8P51Cr+CPrU0Hqivo5mNfUYkn2g11P1vEECY8FQUxDMhkAw++rs5EaxOuIVGb+clvRE1cg1
DCjY8Scqjn+wF2put3InJdy5d9MzMLYLjZugelInbfC2UcAPFGY446VrtNnYx1g88YZqMEx98JaD
vONZEy6qOZS6jQMPQS5dxf91Cfr8qFQw5IhEMSf6TJtq/5IjLgHYlD3MRW4QR/3LdXem+BOw3gUz
cL0VN3C/Yx/grRV1687IFSY1MhfLfD1BW9rDwUOl2xUH1AGVEqITiTGR3kjapHxRD9D9jlP3l6rF
Ss1lQ8VvX7RR2bdQIX9qBBrXt/g+QEBKmA/4PAyT9jHsHttZk6qRUf2fJ8qtONDzUx0xLI1iupW/
/L+4ixN8uA4TNGaxiyivWV/w3YiSy4iCK35pXk4o5YkvYxN8N3vNZ6xiJeUoU+37gXOZuspkVvVk
/4VbSLkAAsQ8yNsVl7/P3GoawHLB886KUIf04o2vhK0apDGIzfcqxDmM6Rcz1EvtkufaR+2J3yF/
tdUDSspvi41KVtdGECvtnQ+lCtGNbM3kYs/wHF5NdmLyeHn3yAu7pcyjHoPTQIfTjoLlWpzZaJAz
zrXWqfNn/vtViLii7064DqGCchI80tSxP7GDjUJCPdo7N6febZDrSmEHWKPtWW7uXf+F6Hyzdl4J
W8Fjei7TCL8yFXlDBug4El6AwRA3CBdTU7MrKt6kFfz2hoOsvrb9HMta6+imUuRaUgUGjQftW7Jc
ndu/eLG8mvh6w7RUG0lbKXIIyR4/GHvZk57LN9g9Rgqp0vEGBwcL+Ac3zWQZaBnpxiJcCQqqwFUu
lv4p5h5hQskeR45eQEcz+zrGwI7dVWw2n/J8OXEpZy8+k+QT9+m4+FnmBIVqUjGWon0AiUHSeHFp
sDJy/SVj4HGcJbFWb5q/XDf/Jd/rjfSI0q3ShoFKqdJPzVYV1ToAeb+dXe0bwwo8qZpSn0aA935e
x0qlOqEkwitX27OPzbbBDLOFg9h0UNEE4vTR8H0QAvnkfhrQI89MGMlRwPUJuliVSiQH9Ae0NKwP
XgKyuk8DsmXbrhD7bsq8zA7qJAc6oFYHI2Y1V87/J2xHFxLbpJTlD8YNrr9F62OArLoLkY4hx3De
P/rvtb0XwlH3qgtnZoHYPlp7ajqi1ARzeNio201BC4s1//tb8JPLWBhgLgBLvWLa/NWUYW6F0Ud4
wIkwXGOljlrT91rB2E7oIK/q8gwo/EKrfaKtrqVP+ZILK6f76G/tdH4ZlNe2sxA64y+Srk9f5DTY
oeLvO5oByWBsm689bF/xD8zTJJZ6+7aM8tlHV+2g96lBm/JF8R4pFCVc9UpH6U4vkRQX/Jah5Z00
GOGm1Ss/AFhd8H67Oan1ni7hkYIvge0Tl0cQDvLC2DJYfeLYoIII5/c2qqDGpyxMb5G9sOvceDO8
yU12ucnkyvK5bm59wxIEQXfWzOMca05ZQIAU+hmBJBmu2PhJH3xXabDikZtDP/AGhIdanj5ed9jI
rF9mWfmS6F5m87RMaf7NSzKzmURL/oz7XHXogVbEAZfQZEMPBEbLnhPC8U+/vApS/HxqXo1ilGxd
URgk3pHu6+KnyUIJ9xocdurCcBH92bBvuMDtj8EM9Nh6rpv+PVwcPD0fdISKhOl00ug5+7x56cB/
cnQMgVPzwEbeceO5JLrF2VRtbDAyH8HQTj1wKGi604nVeA/sqQVO5Mc26IfWnijr6pKepGT9RS13
ur+AETgVBYbYsuyHUNgTKK/r4CtpxVaS0jWFalVaToPWsCzwpVmEbLS6OLc+quMRGAzwsU7PPVnV
ZzbRqkC1/IpG3THVUe+2bi2DRtPrqnyo8CS8i1KbxyyTXdHOhWmXbS3mosErnTkgzn4UTkqWNDAm
SDfMiA6wxv07z7RgRCRmZGSTSpXoMO1esidJW79CIo8kSYCPQCtfM80gJ4rgr1IHj68U10Gm34OP
9PUw7Izfau+D9mXsE8tbRqXfd1vbPqZibChYZge3NbTzTW8+oFqgvRjWwj8MA70ZzConyxjobRCg
NeihJOngNqEicj3CsqLNXwilOUWBD7d/dpcqC1tHEbRAq+GdlggBDC1pP4UdKIco6Z/JXB/iu+1n
zK+JDZxC9Qn7XI9rJdtab2pJhBqnRbDeJbNL56WhedjKJlIbOPfni1UnDGB7nGmZ7RVOlt44ea//
i2DZuUXO3ahwOup1e+/alGZtSNh0iHH/K4Snyo2lxdRI9jqktp4Ffcq7JDbi6VT0sJ7ormwvZDhf
e0/6gaD042AVZiwpzxXaj3SbFONIedzYIIIEsv3w8sxjhPVEY+9UuVHjSM7JICKA/z6z7kqAb0P0
AjwPOPPg0Kd/Ql0Zg5XcsfkbLoYakJRb6HlsGiCqk2+yo7xT66Q9Ef3GRASgWFqGC0hnPS6zgupT
PCDvqSenWWcDV/RWae5pRXKRq5pA7VfPKm8O4xoYiMUENP4zz3VrppTqP74CAhlqp2l/0UQ+mH+9
NqZhoT+S/lhq3nFMeYZ3XOCDlQ1mwtCnhIguquuRG8RB++v8DPv+ERtis3CZduEzo8Xhg+VjKxHW
4EfSmFauaSYlyDYeXFvWxV60omgosjzrS3ku29Wsq8r/947StUgUTBne18w8CUgZH1HaNPIt1ryb
vd0twm4fYPJiR4tFmnoudIc2zGEN4fj2E62iRs2Dyj0vLqMURMRr+y9e8bxDHoOsygpC3jV5xSSZ
Hbz8usNohAZ9afcECQ1djar3wiTvtS92iBc/HFDPhcMo6EjstynMfys1dEW4yAPmBFB6Dr+EcHKP
h9604SCWoTm6LAUjrLqw+o8WRavJhQSTlKo9cZP0t1Yh0JedzjNhLJ1/dry+8HjDM/Zm9EQz+Icg
kozBUnv51pV6Zj9kSGa2ZuPHe9c4J+OQKNIl84GfA/dw60HamY8s9uL1LnXq38yQ7Qdl+9Wl+/ca
opaGunphJFz9rnVVbXF2AiiVAKMT5hgv3kJ7JkLjHKymqHdB6Xg3rj0aeZxGFRp27vGfzkKN7xAP
I/yfgAUAyeZVAHZ1YcsI/lMXh1cNpqIw8wPS6S39lDSJcy7tN3cUEsBSyJa/6qp+eLi+VupqS3rI
+eZZ/DXgjl+WVBJ5q9nFYAYAZIRw1Hp6yI6VVZTB2THUaK1YJ27/6VA7fCBGKAlldlQshxfSJpGJ
Dni1ixwMEth7ggHa+rfePnSx0S1TwbEeC2FJD2P9j4yekXZsbmXDiAAjxRRwXUqtLC36EgUSDVWo
1vufFR+piNnIW+p9MaJMzbkY2s+E90FgKgVg2ysm4PpLDW1UydDX+ut/IOacEjjMVr5o1/DslEZC
7x6Sf1vw+hZ8NakMErqJUFoFdqwqXGJ8EcBLuJy8OXoo1RsH4mn4ggiJKn+xJIkUoNQ2jatY5uC1
YWz+I5jn2QgAXl21ClmhKC8jaTYtYYBL9THVuyPUx1Nq4XK/jljevuaNaAWSeo/mo3REza3J7nqB
+ZlAkRdTy6rBm46jvj/M/HroTkjJS+7FAuDZ/O07bDBAVC2Te+Ui7SLLZpwvrwdx2DR/alWAnSgf
fLUvDr7vr8SLTwNG9UGma11VZTeXUw5pJFVXoqsDquEwqgLAEnzdhndfiFYqqGUhmEmy+7dPb/T+
9yAf/XSWK/W5pVscxf6ASMHofx58/EJ6e9MogLvuCxjRaQC1gAqOnRpwsiKEX2jOtXzZR11y77k5
GWJWlreh+1dbsTU1TUKErL6Z2dN8Is+Cx61l9ECbBmxNmlTpR40mARiHd+Hd5aKMRLQpXG+sthTr
xOh4l1jhAwbCJyuV7rWgOq8aXjyZTGVV1Ju3pCb4TlTIl6fdv9ASurIl9BAFJx+kYExldUrLysV/
yTijFblyG0kvZ1W6tnyGE8wpoEAvImmOnYbB4+Z1Oc/wDg7LwmzVAxNsVp3rxJMrzyHVgW5O++LR
CXZxGGCmahEBENa8xutX+SkpaK5EMlTcdTqmBu9uL/dfzkY+HWNNlLyzJSbSooafDS5eVEEXJFZf
d3oAHIwlW3DSuva3dQ3cmI7/H+f/Cduw2QboqC/u2OnE60TolLFBt9zulSNbR8vLctMcaZaSZ2lC
WYrtWgAlrQMV6F0BFdb9X+Qf6oamMjQ4u6HzgaBCY7USdI3WWt1XKFop0zaIwENUiL9PO5QDly4k
eRqVEoEebcSI57dd72trZJsI/t4bphM/XhlfcmYXEb2HyXLDRGM1XIXvxnF+dVR7JBJLYB6vIwgC
mA/onubnUBNoJvcQvvP62wRhGC7WoCP8rDT87VhMuK4b1LrUO7TAQbNC98b6XdYJRg9o7lhu796N
Pasn4531jvHQtJNHQLOeXjcJzXJiE5W8LR8IBXf6REYqPg+1anXToEG4GvJMsxk4qwZDgqcNHs50
/fDBCvTcvNVTJKU6tIvcmqaFOrEHlnr0mKRgqFoJRXD4eSD6GjScR4dffsH6Sj8dSTrtyLxC5XV/
e+eKkq5mqjsVzQ7n+mmRQ6ef0k8Xu8CoUsldgyftmsLgPbOuGraDsazWeX+thN6i8DRZg0MA2MUV
u46T/u9Hpz0OB0Blvkp7MkG9NJnQIus2WkRnUMttHe2y8KUNfsUep9A1L1qU6BVZfV3PJVXegH5C
E7zhqJYbDZ3XhyJflsAQnvKkkQ8S4U3s77DQ+83QXxELwvTfHLSFh8KsvjDsqLBHBbVhXQKQH3OI
IgudXp6eTfQPLiTHcFp3/ehOXTqHYXJ+zHImwLwj8hqeY9fq3gbaOtYMxct/CpAKpCf7FY7applB
6Hx9YsGaYH5gcHPGLBlckEs0MngFzbDbwKga3IFxxLn8U5+yPe3j6Ezz/cSoYuLpKcHFW3Xl1Hbm
hh+5pOjBUAFPhyOF4pCN5Mwv9A7RrZj0/ySMAkg8zUWgboB4kNWTwz86WaSqLg1r+QyJmc/J32xB
jDl5v81aXNh+70yHK7tXHnzGifvHRX/oVni4aB4H29WZQYpxWp/KSn3A/PAuFqZk2nmU6z2NpfH+
6SWmCIZyiaB/dp7qeIR+OeqOqZdwlgqmYjJnBledH94TI48Mz2ic7yIcBJKn3Xy7zZzZyCxmuoic
pxE9eufOi7NKE0ZT6LC5bzF8nNLCCqc3stSZgjwNiAyTn9JbXD+lgS6XY3ETQ94DEqVfpxa7fi9G
5wD0yAM5TtHCWjGFLhodHQk4kX/mwz4ZER8xqmOh6s3+eU/MFU9D+lJE4u3qW0l4C9wExmuhtE5v
IDP5bCf8Hs5hTp+prq7tzAm7FHMKueTYgZw9lUaXNXtvH/GgsrdKYyCVhc56xVnmoN8Es9uugrcL
PxHF6X2i2Oyrk8O9lQU10Mih9V7So5zVBYV1bHSlUwGZOsgCaWLRWKtsN+OwMJoMBiFPr5iQaTFE
DaIoceMeqQG5uLQvT7NHzxxeDMt6YGtjNu+1DdiggLdfJ6prgcLAbY08qqiWSRpc/bkMlgRqEA3k
mWzSa/mpq4G4lYJHLe4wmDA2B1arVNUXh4zZqCCTU0GGFfK5iCQmLTh96HzXBd7skGrHkz1EBQ3T
L2t6vkQwEwIYc+JwKUNaqx6qYLUBNgVPzgZEKPZjqDtQC+iBB/KCuHSzk2yAmSIQJlAJOqGxmeOx
ASnBM2iQSfCcaUG8QKDVNj3J0Jbh4kFvMyKWUyJDSWYwkME7WhWggBx+thDbqUBYdCBvkMmIBhUc
y8zPjn3YDYHm2U9DLEtm8e3It/MYcjkoMaQHhiao46wQbGZCMvyD6XZDMR2co7C3RaBHlZBzfCL/
MBW8O/PM8dNhqd66BpKeDLWDr/sHmC/BebJIqq1Jt6ikked51tpFQ49EqiQ/pCg7emL1SeKdZtHQ
bGw9aYRJmAcMJLCI11bF4eQeAJdBLBzDjLldEzNaUxBrv07UcOI56a/hdzzWzg2+5umvKLBE3Oii
lHk4LXYGe1uUqTROXZNGDa20oxItlZleKX0recUKsfHZOwWqfvbJHABYLLws6IytvWobpL1MynaK
xtU6nb82ttGYsR2HZUit3s4F2N+GnwkfLb+sq+5qrbwCjMV6bk2npEA75ErB43KIEl06CYXp6J5V
n/1uTuyIn16g9uoMHU+xscg8HSyRcQ+9MJbNQde7cScPVoOqHxFcOhjjYwIQkCU5E6ms349XmOpI
sL4iEtsNsDU10cuROw7rlfe9uQuxmgIHgebFG4H456V7m284ILNh3z6ik60C5cM/U98Lrq+4akoK
Vr+WOZjYsEcRPGrqTPE36FM7DF4U/waaq9Hyh0PeJ9rO3gfXlyNOOWA2c7H1na7Afdq76cWL9ez5
+5rJAgVagHv3v+DsPSWZrT9DwkHeun8d3wW0oImQCSCv+oDJ3Et/H1xGadxv3Y1ZXMrsRsaWJ+P6
HIguKtjZg4IsjO/bmKX/hWRvJMxrty6e1zZMRhOvTPiqieHzH2GY/hmp4O6IaL6KC4hmeeQh0Mnu
yxK8WiSt8JQ8HTpT4rZ4ABasIYTW1kRky1sSfMo0iM+H8k/Z97pKut/YqohAvZMtBW++2HEdQa7r
G4utd8fQxJHsntbLUF1oJ3DgQS+/zaeB2AMaYv7B05CL9DzmHAG+5lFO2BnpexcxhIAxI+QYwt1G
J6K+dIsV8JIjXYsAzeWtfUJpK86XiVopyxUotbtzlzAk6v6PeklZ0zkmQIZgoCdIyWbhbR3rm3CO
jS/0K7gGrmojUsGegLxulZeUVUEOxsiRKkqZIn+fs7s9kkbZSFL0SNLiyl0dRB3gqdNxsJXDIZIb
oWtQJRME6I3HziTI25D6JZmr24CezGplngM4mH9zrhadYIaYea0dkChIu4bVD/52toaQtQ6RIodX
rOtPbmrsk6RUq6RAV9ymjoUPG3Vr/CIE+gaeTIUbTEx8SS55nLr5bGvYiZA42fBP/4IT6/GYaUof
F23pWbxSU14Y8F5QFRf/NEJLocfIwdDP2jNMp4mHznSpoRhvcoGWPWE+aNbfoqCswqWiT7534Vdk
EgXNMFYghhujTgpabTd0/tjh4OWWL64QINKnd8e6L28NtZuaIgYwyiUDQ8PSrvsityXxOFIwAKba
YJyWBejuA6wFmObvYc2701H5eiVRlvYS8JDP0dyoG5kXU/I27NRhk4w9PRjIfYyM03ZDLOa7Nd1p
Yu5zC+GI0LYPJHWqtf6oSUs2I7/3uB4u1I/sjnhn86QzODCUN0FX/ht2a3ddAhmy63vWEj101Ys6
qXEdD1sq6BrE206duGILAmUtKBL1tswWSxmdCJ22y9iGd9ulOJJVyOyntbZ4em6dFzuk8wwj2SG3
EuqHDb/zKcmVQWFeQshv6JKBYUlNwc/lre6OwTbUDHpV3lhx2e42wvVKElgnwF1Lhzq1uNnCk1Gy
oSRZAUc6EPcEQFG5iDUL/ccch2kEMH4yDaF2oVQLMMUPPoYJscpDlWL8ukN6qO4PR30I6Z3vt6Eo
dbOuojAXi9CM7TMLJXZVoipbbQ7FNj77F4fBpodCA2YNwukm+Yn9vMSDzFXJI64C4LtZ7zY3LsOS
sBfU24xJlHgO9vsygLRe1RJry7aeuQmyQvBthEGsfAERFpBbEYQkRnL9ywtxmn+B6IVRD02L/qlb
yggkogSqpJ2RxXmWhw6WfCNxAaLlvo6VL1xjxVoH8vDPpOgpVUks05FmgHrmfcwefXtVUKtNzu3d
X/VsSNVNsttvP6GxOSCQusAAn2DWf40GK1p/Z0ckTCz9MNhMk+JcfWjquzq6yBRYTPIIBT6FL0aA
ZcEaxDxcZjykfPEgX1t+j8ImXSy623Xe+pzH81HdungtG6HU2z6njoWcuHtR4PocgSARjVhvkMEO
WItxVh73JKTq6RKjEUcixS+xG288RyloXGRG2Jh8cyVKUSCAAK843ubg8qe5pxURnhulpqlA6IOs
B3lZo3SRHlwOlOEXv9d5mP6mPuxVzI3fyNhffi6YMeClsKzoB1AL4hPv07oMzzVPE8FNjWLQlZJG
DC353aZl1fhGTtcsRxVXgt/9ZfCrE6lzJEBrQYng100QBEmOtiHPc9X4NW6iZ9xAsCNGrlOQwsFD
MsoBmMO3Fx0oLDuS0sGBjzd0PJhnMNKjFdATh1zAT7iTxkWEWj+Gia3BSwPewutDefqzecqDIyQ9
FYxxNjWQKjabkWK25S1D7R+CAZGjLP9s7y5WW/h1MHz8L3KxGnhqBJiALJHdnbYvizfv24RsZVc1
Yc9h6ERWPTDcuZyVM6wTIoEGjrO2XbE2/Q5GL4m6VapLpu6GPn44H6CV54c4s/R6lPyfti5v9yvk
sCkBt11pe90fIhRgdj2PFd17m7vcDluyfNvluHA+olaLQe8H7XCOKDoTtMTGHuwUmVYTVwplbfSs
6d4nGrk6Kfzdyc0xMNzxVXv8X3+8CYw3paUwFm+PZp2q+RtyC4OZwfMFbQk1z2yCeLWYR/+vYLqJ
OSOa906dmsYvR73h0GwQwrrx9s35mPnkRKvZK/ua7SjG8b7WDl9tgci8LnR2JA5elqkYqqGrSHS6
1zru//U0JJ8HYc4uSldPzg2q8qzQp5xzxHKO4hJLNbg2De2eEC6RGUJCbuzr7/0tK6gFLFGR+Gs5
dlJ5ftN1hpmJ7/Ub7bBPAmmBIG41UuKCe/g09PYAXejMcMAHMHPRLKfjdoxrKmUe1fyySnPYL7Kb
MR8o/+EXftbNtdWLyURVKCpjAhBY/onB8/EQx4qL2ECW+memr3Nx2Q2vwr3h5c1gN6kLBBfT58an
2TFYA3j29Sn4dpJvu7mMQkj/O7uxdrrwW4vo35mKMjNaku3YYZ9OcS4DCUbgUBda5yCYHFOmSViE
9Cs+Tf3gvvQA2IRcSnPE/WaUnv6+6cog+TM720rO6Q1KVFW1NxS0jQJdgqs/4uU6ufhQuXxFVeBb
Vlq29Gk0gHJ2C6VKOEA+cnfmZVGmCYvpjyV8THZbUUixharQbt7oZvQH3qyjxF+YxrfY/18kbsZd
GREV2cWQUke84t+RG8dkg1MwvXcouvUusfSBoXfKKVboiP1QJ1GhgSovU8BcDFmA4J2xWcdYCVy4
SSsYP12Tv1sZBTTY25u3R1iao1rRU8h+uRkOx3HF23BASWmhx+XC5tSJxkfTNIjRdLl2zqg/P3fC
tYg52f9MAAMMa/SwXWD3mW+0ehZfmssjLyio8ZiPmMoi4PCcNnSWaTaBar7xCH70h4t+Y4sCmVLR
DwZGVWq38Gyvh4jVJD1ew70HOnp4+g/PV3lbd6z6LVegNShkOy4DsoCGHfy/o2vhom4m5gqJh8op
vPuzKqRLls3GzjXKVjtvm7321RfDSmoWpJpdKMg8Qqd+n8wSAZne4F1O0z1s/NO6D0tQVBTRc9ad
sLzRKsvIHsoNfqQFSDG8v2+8X+5yW6zoqnJ6htsPVQretbhYoSkUSiV5HEapQTY0t6Z0I3VftYus
FqS8tsHFy7wNPlWeYmFNuwa5UgO/o8F7W+4yLWO30xzcit51R6/m/mK06VhHpy9edThDwF5vj3Fp
1r+9DHkFWiJHL7IQQg/gIma+mPaoOWtz4L8JXVlQA2zkrVVCXclx5Vt3wgyYegQU/aybcj1g7Hvw
QmSPRlZDFXoiiX5+AIisPSLy1wSshmXWA9x/ha44EMl4YPhjUHVsIsJ6TALdEHRArYzBUdbqmD6+
FfTD5ST/qGhPNQurOzR5KzTbPhBrmLftiaPknHKjt1bfuaVlGW14x7zS3c+MCqrTS4wytHjEPGFw
CN+8jca3DUEWBkpz7f/Z5/WEGC/Hx1O9nybY0x6Jqk4vFdo91u1+WerIkiZO0GHF5gos7xf2hOZC
FBKoZV0wojy4T8QA/UcPvudJbE8LJvFSwTROkPgtlv6vUbJcaZnwcAS8HcOHDqkxwiF3QzmWs81I
q4LgaYnSYeweTUTOJ4LccDtM9gZHubYS3qHrZq4uoAcph8PHBf0ORaxrXyUr2PFXe5mNBqrLMHpu
sBUcW9d1L/JGfoPyi6qemHN3zU2mzEEbAWmzdsmSzFDsJUm7r5qBSRjS/rNS9fRiUbtm3lpuY1Ly
AHDuub6CgPBM94jIKtHTSebpZ1efRRkvcrF/6iudRT7f1ZBLSIiKYQ8z4ay7cJ/nTy/jmECqQHmD
FGSz2+nwR8wy669CnU+u0wCG09oRL8qBbAHL18+FoY5ElVL5d20KyUgcspSK7x3AOKn80bT4yAwx
3ic8+bM1nTXIppAIvCFieA6um8ubggypPauieTjBkctkYGwLQxWtJrsNj+wHKzCx4K5661Zwj283
JcPM5OLDJx3joKnCXKFlQ64Lt0uqYRd9hdxvDK7NofShYOM6a6v1g/wgg2SM6Nq34UMK5Cs0rRzd
iinR3IcAZMjWdnA5/oWhFq8biYMip0HXEVzvvrXWW0lQnPWPEo4K8Pe1WEF3agDv69jzkauBGqjQ
NIC2JVMbBQYvGIA9gZ7RVMRDAeaNiFNR9U7TyETAbbBXHTNhaq47rOzdnWCdpCloXxrkpEyOZAm2
qrdWX3thFkvtJjvPElbdl9/sO9SwUCw1JtON3tcsssjEFF3IE0HqYiJ2f49zWur0l1oYRGdLIiyB
vVV5n0/wmc6d2E2Yr7cxSCgRgWBs2NIxLk8TdaH0CuQ8gXei0WnL+9/tLUolmYCgRAhNvtHsw88h
aKl6AZnvPEEI5xyyCVGgWOa1i0RKxa5U3cfN/DrkZlgCFUkKLFhOtzR/J06+W9l/7lMxr4sYV6JR
eKRYdVbn6j3j/a5f+01L/TyymrEVXUvEjMPLJF3etrlU6goWtjdNOMlGkHB46GqRAvt0g44bQnym
k1tKLK7u8CeYC1/PVDV+V6ePHKft64nzMN8SqUlzkO/fKgW43niE7HC7w3Zg5YEYkqF1/kDDzfDi
nxxmycm04GWTIa6QEJa4NJ0U7ed2c14HtTIibObwzn2IqE7udaczMCT4msX1VFptu0xlFTSffEIa
RiXb20Nz8SvzsvYL+rMa97dm6vFX5EnMArjP204pBIcuaqCybWl/0n8hQkkM/T8jNUIR4mJPkV1K
Pek4mcOf5Fee2mWIWQXnmNV5LEfBP3fUkbKCUOYKyrnsHb2OP3hpOnpTZclQmcWRekKL0bfAjuGu
SaRBfreAn5MZG4Lnl1o2drsMhtPazXS6LBUvFpT9/TgvUj3iAGSqkZFjahbc1tzQ1ZlDY5UL99jc
uNanzDNFq071MzYuKHt3soYQVsMX3xkcaNAbXQNhcgxHQ3jifWhgK+a9e0Xx49uwnAtUTWK1Gk1U
JpuaFGtOKl89Ag8zbUBN+lzZ6QhPJU6FUUUL7r8bjRYefUvXPVHFGMNq0OOMQPZbHksQr4EDsYj8
u1HwOUzo3ZAIEd6MFR195ldmq54LtEDyULYDYexgJIo8OoO2eum7JWiNArDLFgqdcoMbFYI97UZE
o9poN8m6gMjZlD5e0BnO3WhqLNSLVVcy4K37F0WOcNJoIhPFsWHYksqyZ5cqPXu+0vkzKGIRS57B
sLBBlc20N/BrahuTweOwxiLhJcUf6b6ggmPqwZiqToJ7sDUIwuuzDCD4a4kOQV2gdOY2wEY7Ij2h
vYXDH8OWIRdwAGGaGgVaAPD0Mjfq+Jt7QF8EeDcAdYRulnVLm6Uzx75I9JvmmedIvIwGWCb1MCwp
tn/6nKzDLY2S0MfNbZCB2UVWljgfRgPICA/v2an0ZcyHmhNCaUzSTTBJZICrv0Qf35kvkBJlX0QZ
5wWLA3lVuc4Vd6dzvIBD3qU0R79Me0cl//IZ8mK1cbq0Hu5W7ewI2ipnOpLqB9npEqBOHmfTpQa5
VzWE4iZcv7lgDAggQxeWBySDSVoy/lIQ77IlT8rFZXwwzOyWEVqcfBVEztW7zrzxyCzf2v4W7SBY
FHRrD68hNIXAjSUoflgXsz2PgR0aLbWohWk9KMw3Bbyw9UhWrbc+fjAyucRD8LVGazVs3ileTHXQ
BCYhLJZIPOs1hnu+8Dm2XUUHueTdfuiMuVfkn2RHX3o2Z320lyOLyOnSDsOnfU6wiGUxyjKjAfHK
+Tw6PXBnwPNV4H0Iscydg32JMd+d8hoSHHJl17ZAzSK5YgX8ittujlZurxJxGV8Kv3V6wWlevcmy
nnM4B715TpXtPXNKBIWRgCoFLHbkqYcElEx1b2TbY9IJMjm8HeUx/2zXk5VVUqu8hX0L42xDFe21
sVTRoirsPYLY5qUyNM1VigJr8SUsf0NXlgq4D5MfS5aG2bwZI3Y7AsGpxJLFBj5vqRCZwTYHXImd
itLgA7glWCgA8L/Yy/IVuM5ZCorQz09bhk7kQNZq6ZBClyJmdb9XnuPM77k7v0B6u91XN4Y3tOJS
RJ8ZwwAC9929JVqSLV8hIdDlnXKcRRB/bl8bFJ5Huq1Ck0JEB1DzvD1/yNThBxUpBgMH0RBHcS3/
ePqJcCPwYwPChRVLU1x8lMLkteXSId8HfV4WGiixH6avvg7JyregnLIB/Ofc+woDU0iVteksVrLG
Z6r2caCQ7rwt4JDlp/wphH9o/ZGdwal6nDXAylp0QMeFrGL5L/WRoQw7rcWcya07CkyMVnZ/j/EM
LYhmC1cV0gtPwQeXb3TUc1VOk446/FZ4t3pkzk5KGt7XP1KilluTWO5Q5FLlcy2YcGZsnu0L1lMj
UzwfqE+ocQ9k8Q0ALo1pxI4stUhdAfrMBPzBBjNiDy3gWE0i81uolqM7RQ3kqCsDk6fuQOXRbt7+
4V21Okh35GNKhB0pfkY8EC5TXw0Fex0pwTvR6apHjcZUBC1yizb2aNnFSgktNMfxiN85AK02L7bu
jf8V+1ZqjiwQs2BTRtc7ce5Mk3QBTUu5hWK3wakAEcb4jYN0QbvQcomYDLn6vJ5vUiwIHG3bAfYO
ia/0s9Hwa7Zc0XA8IxtO6acZbo0oUrCZGqXZcpdofq0IPBKULAmmimeEJ/l5OiqVEtgSneBAjS75
cZiHKureHtiRw2xlQm2oqr+jKq6pb5B7MQGciDzkPDhsfaZbTwPJaDmGpKlK7X7FnYLTXNpjc54t
A6EPpUJokYZplA/hE48UvcgBMsSYwa1QDGan1CXtfUM01U+WirauHs+8JpJ9BlCk9dz+nwVD7OHP
IsRHcwhKIP2y0Vt+wTXS2IvJuSp1p1tOL9PjBMysJOFxt25p5+ypozoWSpL2zLkLEJ0PxGXsoolS
rWvWXZLqVDPb/Tg6d+X+0qxy8Qz4Am/o8R/A2cFt2C0TAWYn/1ZrDW0TC6D/YmdWBKyVGNQ5CCFb
bNvDY15G6wcW4yqLJ4++Hb8VAv4kUVSiCOf/qHIEy0RRx4siwDAnWzQ8FPbTc3sXnv+HXkDkR+kQ
KIYpxU9SfP8NtOc74b+E6yXZXqIeuQIOOaHX5EvVVdCRO+V8tNrmGMspgSd+hwsAHv0QTl6BN8qi
zkBdb9sNoY4AtFAk7DrWw450DDDPGDe2VBopt6MrJJY1ZjIvqtsdThz2tHiuCBKCbD5m1AziBxgi
v43hju60SCq+sYFs7q9clEtx7T2pRFPQZZTOH12G9TrYIzoUtLtGF94bNd9anWEdpxfBOzaMibzs
seKXeByAKZFE1MZGGSwn2vYkM7xAPqD5FwJiH1t1j/hEdWqkMzuxA4jHSjaqLJot+s4wrjPF7NJM
E9wu21s4//KUEwhr29W8/o+EMhTQjqh7zeIkmPW+zV6iAp7zAzCCoCCIhQB07EmkYeQmZpsEZuk2
D7e36lN5ranHbLHGZROEEnkDygCxHqM8ae8WL5UHNwKQCx6sa53xkwHVERKM3M1p8YSfK8OYPPqx
QD+1s4kOA8t/JG3ZeTONNXa4FKsqkYrR1KRPQa58C0qxJHfFEUDO5yg47D/WengCqC21nVlcKIQF
nM4JrW4g/UpM0QAC8WB+mcuez7qs9mK113DJ803/eEhB0zDP/FPj2LO8nmyKBbQS0o6eNcuDjrtR
VUTP4zgoq7WR64LU3L9C30I553JxIzOFKgUjmXVgWoNACLKTWye3I7OR7DdCdcpz2T+8X8FBpEsn
RsX5Oqi2xMcOmaA+vaaXhbo3TMZqLuJh1Pzr/Ih8N2EsZF37vD1zJMcwZCqbONFogIVajZE8rcuF
KlZPfR3IcFdZMCc1fLiLYCxsytyssjMyk9ExmdmmaoGv5v0ug4yYHZvwSH/qpAOUzjlBEjqPB8RP
9qQw5txkaZi9mCoreadf8eAGaI1uSZMMIW2g9WLrW2S7Tmd9OBD1gzErplOtDviIudqci28FPduE
LZkf/+UxsXSgU/aDK6N061tfRM4YY5igSRHuVl8yhjL1zzAyDPregMXGHAOHqIjdnNK6e3mti0jn
b1iv/hMLJG5nMredVT+/2fGlYCMi45eIBBvjAydKiwrf8ymqpKqgmQNwgbWI1QbHEQzhO5XpD+rH
2nRxs9sFqYPSFZ2VWI7W1d8WVWnYqdBytg7WsO6G4HC9G1BYWRn0kkePA0ODiYgLJGiVZmH4a0Fv
EzHJvAO0F3kIusWybZDUZEaTwsbUhybjSHykK9xilRVTHyR9z1C9yUu1PMPIYNykDBzv61OAueyV
/Mv3B50Y2mkvkid3emQZb7wFt1MiTmlebCYNXC2ahXVqX7p3da7kex4I1jq0xId+zo+Ox4Qld9V2
ybjeiWK9far7yfq23ToQ0V2iJZfzGZHcJ7VDeIxMl7A7fSLq5rJTrumaQ+lMj4C32xSdFOv0/8nk
Ep6QVjxmqnonF84PaFk3nfTw5p5vxR0FySwotuaRS6q7j/UVwvND8moNQMG4EMeilqp0ZoSSjE8c
50Vongi4k9aOneyKjchZoHSRMxeWhBViANuI2k+U/8huG/i9H6aNmL8VJohJewsDuYMStSrkf9SR
0w4oDtNPWXJs9rtqqhDbX9AcAox14o3+Pax6NhUakFdF5fAArtWbqz0OLWVnCPaIc0kk6HLG3fsA
989+D3nZRG1kp2vQS/JA28RMAx4ChA03AHPtOYDXOBXjBZvy6r1mC5iDmBDdn+CkrCge4Uo1Drmb
piX3i4zbnETnPFn1dm4rqUpjkSneboiAdoBDWnu5VRLfELGuZcZxFmUxLQosZQgOMj0y6rZRTPwF
7Z5B1o+AZZY5mZzeDQ5PRLbUHRRcToXGTNfwDP33braEnSjSnLU8CLqeOMnTNJa9A8S/UZ8eOI/6
tMq6eEqmw/E8k8vtzcxzvcLQ0Y+i7RsnOQr5stlYvtuGcdbjkQGirLkpF6netfGukmU0hx6qAMMS
4tuW2gy4JjflpymSc0YlUObaJdYrggawzh6ErjpAVNIId3m37rFOx9oDlqKguJ1X4rx5+sH0p98x
NcA5lhY8FURhWnVEIYJgYia2ubop0TUU4h+JPR9tXuaOKOSX/aWiw+YnsbepCFLZggoB5KVJ6Tom
KTnHJBGXTwo2AW2RQtpHN/pxtpXZDWAj6AFY1MXWNljEYdDbSf++POt8pJ6kO1kOWg2AMOwvrsCy
/muphmKpu2dmrYv9RLO1BBgfKz3qomLxIQ391r9d91mYj5OHsoU07ZxnoBycvMFuNgvtouOeu2If
se6N7kNso6Olyk9qFB5slWDvE29jT0cLumKAFfipznoUSuc9tpRMS0eEfszrdFQbAfDZFRNikt6s
vRTH4DXKep4aA85gZEaH3ODxdBbAALgojvKzbEQ6A5AyZv0PX6mtpwLta/Gg1o2A9FamB66VeN5m
VPeuFIPGWWA/PEFmhNboO3hpkDp8QnbjdiAXk5o+JjIqZ0bUX49bfMhC4UQ0VTCj+Z/O0Jfcm/04
BeH2ST02NuspG3An4kJGR9aFo0pXmItayrdgWJ8PHZDKJcb9MnXefFGVxONLf1WWMmw2NbQjRQpX
4H6ahuEH+E9FjEcLrX9OLv8UGVIe02VswPAKGB11it5ZE8Zw5mfWgRalNcUxzQbmc+rZGy16qgrz
gwppPBR5c3qEk3nXi3ymmuMwxylq7Lp2bnjL8GNN2pt9AKQ2qgj6Glf9o7o9WrHmWYrQH7cG7xOP
RxkWA3smSnpnWHQDxYmo7ufS3xVbGqzp5MzwOdV3Lw1lVjXE99lXBksdBMvMQ6B8K1DOPj6dMPpy
BikYSx4mi36ZWL3+dtlKQklb+pQjNz8awlgZtpucvjTZLu5ckthdhNjJmrrFsrfYE9JHjxRrK9T7
n2LiwgzsdmadNoHHvoUXQJ+eeTEqCpb/Lur2/wrfizj0CceFyYJ2bUgICZ6MQ8oEAIoUxhOfDEyO
N3uHLrbaMp+8M/dfuD2xh+9JVJGezajnaGoLLDFEkdHdWYlct44cUcYt8R7vSE1hGnh+lRe6IpsV
McdCYUWwUfyAC9vhyeV5fkmc8iCa7OhnarlhIOTVe99yxqzP7ty/nmYwkEATlfFkGBGQHfoO0+ct
KXSW9/MdF+JXkHoMbB3OJOfHXTqRp2Jfnzzeppgy1U+LWE/MpKYre6xMSloBoyrvjCJF1ND+8/jl
nH8QkyW9kVcRY8J1r6WlguvsPsx5qTj3xUlZayP/DFEGMo1SgoKrKaj6l6Z40LtWBvXiLjTWlc5I
nYFmrBqiApVg60NLK+hsOUb7+3KXhEUWovlv5dlTHG3mqJjoW4tgzt3cdgUYgfaRDnBeD2WxGABT
Od5TwxyWRiG/v5j7ZhVfZlyb2JZnqA9WFmPUull8LUfTBz/vfSdX3MmDIVglJk31hd3JlRjcOgnk
s5ipp+3NZaVsxBTtoBUIkAAdkt9IbAT2+oTjokDEk/z6UQMVqehMBdHoF890eLrP1pbKyR3S6VrE
jdQB/bjTmB0vIbAJqYKvmt1p2q5hOTnmKsFIYH9BWlU5ddCWKsOqhm9slJrXLg8IGzOXjvJ1k0Yj
gA41Z4fz5tpxgZsiuOiJ/jaVCZUBx+CEuSpCkYokx1TmUg1ETEXodF01hyEWlrsTdxYSDjNyefye
XEc9ql7Eyl70xij5RxcOavthEzwtK9nbrrGJNjV6N+Wa27JaseRbvXQdwEeVei5vyalngWKh1fRA
MM3IO+TR+fhDjoiBErYDU098T/OR+ehsqh1f0fxfkVtRfKCgiFBPT8rcbdir4YTEg/DbRQYWeIzS
ZarpX6tRc3BwCJV3LkygYQpb07HHA6KfSqAofTBXOvMmDGP9FZCXyLl6lpcQQGfTop9ddlOfArjK
LL1JizvZRQSyV6SMmpXs3AbQ6N3mWNfmu4m4JH2QY6DaVWbMGW2BShnXqP+8URdRGDN/hGb1IXlg
DYzklluh70tKvFbL5GGAX6vJObQLr3IEIoz26m7oT2nYXul6VqzMMETmG0l7lnNku9F7de7JdeSV
1u/0h6heTcRaeUJyTvpTBaobKuBIbBzZFeTiuiK4EilRlTJ56F8mek7CDcAGzHaqTyp8UB8xzIMX
Gy604K3b4C3oiRpsNFcx+m0UaZN4WFjv4Ggo5R8VR7qyIbf5QyXVatRj40BHcvaXtuboLCFhBDaB
7Xiw6Q1JK8B0BYSXOulh8v6OieJq8ecIwEx35QdjxBcYpJzp2Xbh7uESzInegfOEaaIOBlovoEHL
+Zv9pNlINtSmLrxZPDkyN76M1DvyWCZoiF3Kty+WBND/j/y8aENKl6NK5aa7JxgM+wZKlQYarO4v
kr/chD93z9iMxeKBmfi3XX5cmk/vwfg7jkEfM1/Ga5X79COBj40X3EG2F556YPUqUAOEqXetyvJt
Lr1mDjhtgubb3ZvKPXzwU2mIeat5u2++g2G83FPf496hkiOvErvBI5LSGnvV+6M+mlgy5/2Jd5zM
tIN09w4YIlYOs1Or4JGZIe15vd32nl7VT7eLe7iR+yL7T0UsciN8t9jdGsR/KNSZXXar3DVaKh21
pFxiwolJh2f+LTx1so+CcR37HWrz0ZsM/Ue3Ye2kEM9H1laTRwAxyUMOHTEkM3bhDwPbpjPtxIiq
qnqWjXbz9AsdUyMtaW58dVnQgdq2CBWWAHqYUewVx/HriXXbRvzHoj5S7m+z8GEBiFX7ZELzchXq
6Bk6lw+H9sGuPkqzrVGTiy0Y0To/h3QWHI13yjrLaZ/Gfig5UyJ4ywCM1VPxI/ZjtxlcOFKc9fSE
pWCqTRNm5XZgAPJPqC83g2+P3xwnu+12gwR/38r/EybH+X/H5z6KWmmOst9eXBQclMXfRnbONkOi
W0PsYuYuKSP9BgTcySilqHxuE5O2ao+ANq4vT2gZWuypggnYzQ7rf7+8Ns1K9OYKyDQT+kpYyH6E
7eyF1V22H4NOZjgGRGwWrRtXo09b+J7Pt3cP8+21g6+aXU8AVDdc51RTp/ceJqjEUUvlQvE7GBw1
gNk2X/IePt3qpSSfWYFYQiiNPfzSmqQ/fxhBd1wwbdYQfJSxl3F89h05+QBt5KwXQuOTDAlCri1x
Nc3aE+lXYcnexOsANwU1hB9a168aHkBEXF4MNcD/tvAa/pdPC4lD23L/UHWF2AugBk38ipQt8nud
vVToNSRvWOtdJ6vht/E0+83B0IRCs4hCCv6Z/E+1mJmiOB/unK0lPGbGXB3qh5XkDDs5F35V8LaY
KTV1thj1pLP/EnZIdrrQP59CqItEmTIHwnO1z+GHkauTngX9tHUI2PzPGumqvawHW1whEogB3ozx
gZiO9nzDqPfnORJhzztdEBTRq0/moYReFoT6RaWasnVBMYbsAiOHKRP+WhdGae9QLlviFaeOP7py
zdJeZYXfSVcJsmyWDPTIjvjTELGD9YrsBUiGrSeUdnyiWHODBaj1BSevmAL4N7hApmusoQ9ZRDiw
9yyomTS7dXVnRd+nPc0Pkspzc61u+6we+rFzS6SGo6DmdIH71cAUmKgz6vcZMwodJ/xLI57yhHTE
wFUBbsNxcfGLx7EuU/ckJegjfk1H0SG+eUrwl7EzvyfdnOj2+zhmm5OYmJ5nQXA4oJP+w3C7eSay
W9yhC/qFDwUjqL67oeyp/U+Oq6gdOoM7xi2KeaLNPoCsUKjowQTVza0y2c8Zg+E/bwdMV/3ugwrM
twFH6fpEy7uAfQtIhdJspzNo7qB6eCjtuyg5zur16VVKUqsI8PaCfBuJfBwXmSwLwWhrslQA1C81
Iola5/CLVmjt0rEaw2pVAzkEyXy/0xvtKBSi6eLZTnj/oM9TDNGNFP3Cr5jfxPXqQBzRnzHIk0/3
CPDJcc2LFJ6FnQUjVRy7EcHsKtnh6B83lyGPtIJIJInWV1WzuCASLvlxUJfUzVDa6Q1F/MRedeA9
IuKPmt8D9Bs5aF8b8oRor7vrC9rPcL9GBdaywfIqnWVuGLstVY/QzHBbWV0cpVEHqKRGpDUvdq1M
b3cfi3YmzTwh1C7Ge4+DpV3bRADdmDGEb35b2r9ZrzavYTA6BdtHPabR9kjmszkGWDRbCTaijSwj
urvIRb25FTl2BbiisVV07OFzXov3CjSjzi7pvvFlj3KMa6SjawSxTfPuaBoNxGUpwL3d9Ves8Ps0
9iHQNGJaiiO8mcQDon4xC2JUdm5TCcoWbOTHW1H3vYyyx2Z6g+RthgfFrfoFNErVDGmtPGcto06T
+xTjUBLOk9OaZmNhTRm7Dns2oJenTJoqLR6hvLyl2ZnnJwqCeSGSiPJ4So7R2KJ6ePODBuP913ue
V8Ujla8RPy9jCrCIKiYCcfnr6UN0xdEZk+q+cfWjG9wcErjyRN9IjqPdQkBstsXpQEBYWF0oFwGr
RKyJcQn3mJe9v5yA5S8J7ZSUBvR+5BpDRQRRVVQJuCLQEgNWZkQZCQIF4taZAYDW6/Rh4hyehq1H
C0DPzUvdZgbfSnjypqQOLNITmn+vo/Ky4VPLWoracs069I1vFUbvayIxaq8M5aQ9RUNpJOweU3uk
e4XkRnjofmi1I+VeJpWoIP8QBjWZgJTNQoSz/tA5vcQtT/EKFMBoxy700JrfU3hLjeIsPxUAuOil
ZlP7LYSxOAS/yuVpPVCEZW4Tb3z5zMZ2zNAxd20o2KWSD4BVAcMPxm5+0F7iwqKUgWW1yJHJadS3
lV/DaCtAxA95xneG8fnbs5mRST9nd0JMJC86kS1lhA9OuPDzc3atHDHe4dvcs+xnTUsIT7gN46aj
/RHAST065c1+fa0hMnRx7XOnrgGh99M1jmz/sYjyppR4UD0QHoFsJeMfYQPkyg7xwX+BZFQsCY/4
HPVf0AmPfb8z1CC/0qFl9ij2qJYmMVY7lcX6wUSm2k+9vp2XtJW9ZVxwMYa3MbZuq2TKhPn/fHCK
90eswVVh8vr65J8U/iKZlU/S1xa+GWYahEkr8E/bhJyrpW8NM9532epUSLvVcJ5m7sJoaT4MbZar
S2bnDuWC9KBn9d/bOB5pIzea0vaYSeeubsBdhvMk9suG42rjX7mSaQC+9rTCV2Ks4cLfnbMMc3OQ
eYYZnQXAxX8/G8lYf7D6NqSA9ccu0HzESvz6fbRbec/3CdOY2bK+xr1h4NoTd8lVgM/shKF80O3s
LGx3OdxZ8EUp3mt6zdzks8HENLOZ/Ms0fCY0mZZCo23vgkWw0IpCTvz3xwxw1k+G7SikZ6zeaW1X
FqA8APR3uY0U1thSGRnWxA99MhC8Uz9JlQNZC7sk2/FKsqxBS1LNmeOmCUc8swhPyilvJt0JaTf9
cb3b8ty35dwMVlAi8nXAAj6llC6Dp9rK6CCYAK45moaga9gOtPwXF1gJflVNLFPvUFaITbr2RCiE
GFR/hfLLDQ+S8m8pxnoBHg9oc9MQhvrEO3jl/24lwJlP8aIoZrGvpnTFiC4QKyDXa2NdKayCcDJF
rU2arE5/9is/5+YlRptIrHfkTmsK+24fg6ivbRzbEUzaRkgtA3+2TzmFrEw2A/FIdqrlG2sntEXo
KW1Ttxy9xACtm2jmpmFcs/u3OR0KLiiGE0CFnP2by+l7UxMwoXSS1ObRexpANWIcmXg1t7VmjE+W
9ytAEhgBb7PZgBB3ESRcY5eISCEosBTqycOyApJQQsf0uHtA8ZoyrL/bnMRjfVJ0TCII7Esi9ais
9mE9BWM63l/BnxLhStRctkplhRBO3KjVFHMvuFOyih06tIvSKMM30e+qvut4d5xnykjScFkJQL3W
6CVc6XbvzxSHOJlP63RREcLy9rTYQrS8wZ8SqA9nAe80YcvBiF2IuQK4noCd/206c1r0WamJiNsO
FJt4pjJyo7UVyOUNgALWTwftfGy9e8KNcED25QwVjva0qcsXoxf403y7ytvB8krgQlpjGev/7U3v
wUKjAqixmtFUbbzHojV8W/9C3rPHlhxGTTmX9eFCmsdEiI5uKdZXxmaAgBIvISVoOxfpa1lCYJnx
N3sE+FXY5n09GfyEpHTIj09RKN4RKdN3AtMV8n14YU5DG3zOqTXYa1GZLV9uQL0ZSonoYjBUh5ua
fdswfUUktIOjfjWkTE77MWxAXdMJdTPplrVILlilNmWYemDm0k4iw6v32JtMcPs+Ewi06mVt0l+J
p4nDKS56u3c7us99LJ6Rh58QuY4j9j/NrC1lZg1k4WAdq7AUgdptII1zmnlqhioGgMecAXvbv7nU
HhM6lsdBj+Oaz3BIL9iVyQTQemEaiVETcyN5wDQPvXDFjHfYwt4ajju89p3C+tuUQ84P315xb6nm
aXXwwJUoActENs3tiVna0j8hExismD8xHbr/nF4HiZzqCFw46BPePKfOHShVgIrKm5aGwA/EC4Dj
sdMJ2kq3pxa8vp6ddJucLb/T5IHdMzqnIiNouYH4T2j3bdQjbptUMhg6DcrNLbg/sgUHG8sqFdEN
wZBWD9zpkE49+3+xY2BVCexqHu+my3SwYxU4aDTVighI5L2L5OqRj50ZE2mvGBqOmpm9pKYV23po
/3v/wxZf2DGDPWiyGoQZJihTTdfv1xyHm8sGdMf+fZwzZvdmCG8W7X08qpWIukDS3QHYFpuPqlX8
1Bt6NdzM99GgTKQmgwChZ5+CQRH/xS2MF2xkmnZQBjnYFMRE+tfC1gFeJqb1xm2ZpycjfIIz+4dx
7+UYKMy9kDFe9xqFVBRIDqinuC9mB4Kipvdaomk3cXqQQVx769S7UzXT7udQr9GNyGAnAHNu18Vy
dTTz3OgpcgooEQW0tQgWL7EgXs1/5jdR9XGnPrIMV7ntemtcIRYQyzyuw5+srHrCvWl/S6e61/7+
DuFYuMSFdDAxVEy5SQdtLGd8W3/nNruUaWl7TJwC4o1RUToyjnuZF5eEPzsxpcw4XoL7Jo9E8WHd
91zbjyD9XfD2cmE2pe8ZwHRgaUwdXv+RQMwoXHA2bjRoL27l+q/pjIko/KGKEHwymuKfeVyoGEjn
TDQr/XeO9psh7U1Qu9BI9hQbp4qjQvl+DQE5h7ECthhg0AfYACmN3vmxVyxb9DFpqpXzHFXDDrFQ
qUmTied9eGOtxVIkI2X6Bn8Fx91ZijeqEi6OoYJ4zH/Mjg4x6BUmj46RW/ERYTr0Ghv3dtP/Suj3
k4RgdXSc/qVt+hRvYfPmr4XcOrf9tQpBSPkPaNDrpwNoWeIfNOWyJMGrEuUNuXsWAy7T8MSmwelt
lzgGOHMf1GhXoFmFjOi2sdK+PpHspi4+SimcHMCf+nbKMh2h4zjZb+eDnxTtuGZmJvtmXTcLVdVL
Sz1vWXw3LHdpx49whPjv21bIZMaJ6DyXvwfCSnRkB2S6t+ra09HwsiSzjmqJ4zx9EXEfMQAKT8jE
lDTkjNShFop5/k1491JUqZeowPLrDSReBV7R0vRcwIEW4lFJZXIIw7feudU8WBTmhRcvtE+yeN+I
uwvHyXUgEOvvdUYdFiKvsvlXYTIVGYds1JNS9DvAgbKpQoxm7e2l15UWDDgHSrvtDVn+a4DkNFxk
KmBLZUUmQ//ey66VbyRu9Wf2ygsi0BI9Xk/LkKoSUjvABGKr6Rsm8VZEUsbucJmc9oDABZmlS1Ir
+oCHyPcUD6Z39DI19lkytYP/lYD16F9ky79mArWa8l3ysbW7likN/cHxuvwUCo3ex5EwPm8m+NRm
N58oMRW5IwYurSUz3fYnB8lgSn1Om7VRZyIrR5ptf6XM0RFFHublSzWZwBbD2WA+j7DRxrSTbwtZ
cixDUqKs5z7FyQcXbq3r9FeNuYMas7TE4my+kbkZjTDnzuXIBp+7s/GHSVKHMaNF7ylZ7mXKHffy
p3BOkUpZN1mWPar947Rm5hqMGG7zqtg8LFo/7Rbbac4pcq2McssMpWr5lmPyS7kKUAyFD69zYqY2
V3n1JtYq/Ea6wzHpBPqazUXsctlwYa0CR7SW13Ad0S+zIRO7LVza7kDPSkevjlTIoxwdn0sQ6SuT
zxW5LRWelPsBlm8oOrNrNDsOohZPbEiKhHHU3h+cgat5a/dCYK83A9faJzYmdDCrFAe/wqgy5fwY
uCBwEJPCH4JBQM0nQdZPt+XRp2w0VI6os8OOelX0rBB3IsDX7PahB3wAS4qRqERBi15oyhKbgM4p
LVyRcgAUo12Fp/aQ94y1k3XfFmk1d4eC1K1ICpBpnuShYiXGL+lXmzLD/u8Pjjgx8/3lVriQKEdc
rMU1G71d6r+3KQbbKJQA3kJ6Danp8Pitbz+G7BGxaEqSTvLEuRtM/zgRXLraWiTXbZupqPWvw/IP
nWa5Ire/sH5V8djIF8pY8voY8ypY/o5BgAuGBwQOz+qWG2Oi4g/YHNwt3yxE8VOBk51dFw01zP4n
chG6G8f9JvQjhH7CegRljSqR6s0lad4zjPkd3kFeTx8BrMVj861TmEEnI88e4BtHqtzhrGb0zEld
IZv1MQaPopC+ChhTk6gfhJU4xfNGVnSePRN5dxWCtH1kmah5TGNSJFqbgoUnp/ypRuDUox2lVr7E
/174V0/soSTWw8i/Gab0UoDKM1UbWo+3dkSof2OkrTUIev0jEYA0nHNsoBQX8CUI8DQmeg6GOX2e
FHLpiYlJ5j/XnKleIcw5yBQSld77LdpEeHJCeuBqVs5o6GngGQW4rfSZK+clAvtkezB3H9A6id98
F2SwQP/ARs05ZXZFbHyXH4QIf7430cLztsr2GMSTyA+j/H4gWxWGnT+06AKgCpzlvFfhqpHOR1E6
bKMTMhz1Afj+6lLHpdF0WLjnwPHthnWh7N0Qa90+XprlukRfPWFNUNBEGBGbfXqBY2JTMGYySn72
EISrBzBLHEg+Gpv24gVbTHMxqICwrIv3tlL7WgqKEh0YnH3YgVe0swb0y4vbxs5Y/o5q1ZlsChbu
6qzckzz1RVPDzy86n2CDsyd2TnsHIYKq27FccMaML6A4x3J/jJb5a4eYL0Fxf0M3O2EUjJMrBsmN
sOgbJjR0SJmcMlL+7FaMJdqSIQ3hcRNmtLpIiZs7DJV3BSJ3NQi8OiKJyUSIGI0B1aH6OK4xnnpq
8CLr8nTKVxlnoMw87eUEK8B3QvWAx2QPnFQlHODVqyz2HdFYfJ6VpNZUUep2DUQ1R7vW5TWobBqo
Fvs1CN+exyCy7w3k5RonCoq0jiafJo5bUIjBZWGiP7gAGFDyuH6KEjQEB4p5J55eQh4977dXOpDk
gTLtG7lw00+j5EB6RWGqn5JWWRplW/BO2wqO6kgwkH61LGwH948DTPe7D/kVIdiHYTkABuiVFqRI
ewe5i4Mx+Nq3O6F8N8JA7FXqHz3aJ9XTHM3AUQWVZ6XXWvDBhZ+beBTgXi13IwgiZ/FLdWozGCxY
1PESQe/p1tQ6mvFlIyOSNsZcWivLisZKQYmVkhoBZELU8DFCZPnfnLWkmhD2DdOYDWMoE1tBSi4s
L/RmGf9usaO1IwotuGu85UgMSMaVzwWmjEILQ9TQgd4zM2cPIebFPrdCn7Iuy62pKR2TFzSqhzZj
lz3sid4AJWElHG7iUMLfc0hp+phc2euqnvhOfIKGvKOFxvJdCl0EvvS1gpKmA+gQ6YgSRRT4hDk4
r6a9pYlHWdTYxBiE6yKy80NDll2WvodSp9aVJuTzCqXfwY5oxYcg2xE2GWl0YDqjERKZ5b6rAIqB
FpCUpxOWVI/jJRfuo/kt5BIDsCKQbr51ksGEIWCd7Ki0t6ewcoadEOFg3dzQ/8X51ciuSyx8csRc
6vwGut5ngTJa8tUNCfZNHhEBQ6pYJJzkmf8raRC67xTHp3KchWdmX+P126rWv2G+HwdE+Mj3VRwE
UGB73HUvV5xDU+fG5y+A/Ea9erioWqCcaAzpsPWoRIqARQRYaYj6/o380B+4WLZbfxMR8rT/koAK
oBQuyMcNr9c0EQGaf6mVgsQ0tiY/3HSRvqUiWzZrZLo1zNXKjsFCAGdf8CTLHKFOl1iggh/n5s1k
Z75R69Ve7gOorUOtsvBQQdLhW9jEJaq7efDkxkLpNgv0FHpE8M8VLt1J7MmGwS2SM0mREWDOQbl6
GMEWmTLCCCKR3hZyKgady2KWmb1c76ISLyD0riPq84pjixnKjpz/LhqhWDZD9MbuXb49WEE+VrEJ
mBvZgrDEK9l9BdbdFw0ey7R9jo6OXMfQBfXykRcDfaHxIp4AIOR+BjZrts8dyXYhJE24kBlzzrsw
vwUpk+vdEMDjlRvCDmAeGlTpNpr7OsgMavErw0OYk3QnS8q8qTPp9toRY2VDyqaks7OcLnLajfwt
yJw2WIzI1FeIXT1vX6ZLczbihJvTzgFHKILAvLnhCDuxbN5mRfK3qBm6yV0Y9BaK3GduqwLyMq7H
e07VCd4vEK+XFAsaEG6EGB6E04bCOKKIQOAp+z+OmYt9g+t5dv+BQforkuKCHtMQs3w1bd3RxZ4Z
dNkQKtx5eJphvdkm5FEaH+b4n02lW8IUzJh6fTxTiqX3E5g4AlU9kl75X8aR2d+5mz3A7GPe9ik+
/Ui3wIcyjqNhUBomA7DGSApiJCHUH2jJuxUpDwC0Iq7wyJEuVSISWRsvpT0txNqu5E39jzrTzumS
9JznC0uARHs8j0qWfk8oFQfoFKbhq0p9UiANr6/3zvsKQmCKp8xmqdYkIyoJbFhPR+bMpWUuzRCu
FUPxAPp4u/X4r26d/Z3XG+sucmT78Xxv5dTpsFuLcs8dJ6i2F+5c5eHR5twKt0SUNjjLzGUbbfOj
Ce5DTsMaVbyT84Dc2hkL54bDmKNZMjwrRH1g7SVMr2JZV9/3EQiBozimmaso/E4hRRZbGITNxRvY
t3bXAs7AEClBnUxrhTcBlTqyWNtU3mDfMDpJElqNh3Tt85DHIjQRxGrWZO440q+n2Wn8GryLsgQp
hkeHKUcDl4a1p1GYOnz/CSuJqC/6u6rSRWOXjOuviVqPPnFUqk0n2AUbDW4DNmhtya/V5MIlTyb1
vil0M1Q/YqyiUtryHV3GF9Fd1RzyIcNfK/64Asc76aOeWBzTBm42R/u1sXJcweMEezXinxoi9SFt
8M9d+IJm1YfoV34AKD+oS0W5COyFDM129F74SqPlc8rCFr8CaYEFw4SPdoIVw5Cp8muzHsKqds2W
DA39Sr8xL5qCTGk6iZX9mFsQlDbK9iSmZRsAA7SzsyVwIM/KngCwIdFcTo5WtNvrXrZVmH9Xdysv
+nbQQE6TJ7AuQfXNNd2D2bRqCVogAmTi23mgX59Je1kZVLaYp+cVkFE66AfPKboaNNHXzMA2K4/Q
U47bkSrf8JY+qpZi/V4pxYiWvFSlnfcGx0j95pTe5DPPiMrK4mIwRVYuv737tqIApsNGYwVDmA//
eqLJBCTlTgxM/X8nNA48nNfBFVtvZXslXSGBg4liPlDeAeZF4DDGVsxse5iqH6s0CVyxFTg6dlV7
uitLCCqt5YLhPfYgyvJTNq7/gBbqTjFbX9PQ4Zfy4FaZ78OLqnEd+sirt5oA5BEvYrhQmjkLotgb
GKZDkD2YqYxieXlZeU6ZHZmaQH0dRBj7qaJ3h0CLPoAStnbqCnY5TeLP73wITAr+nBxsCWJuNi2U
oYkiNdt1FzwmjB9MuKuToDy0F4CiDzpaf8hkMRX/qj3YrEl0uPiquCHF1KeEsFRhCFM21mEwJJHD
AyizVMikm46TgCgmVtw51BT+b3R5bB8yAn22YFjkpug48mUf3n7Vr8vPK7GqJjdJo0XR7TZSY7O8
vBDs15BXAgPhWa596QS3wR0R0A3vvUIZh88tiWNB2nTxW1G9OrdoA4mNHlwaDU/THY+WpqHI6JLx
SHZHekwMVFT0k318GQRY3oWH06W/8WVD0JH+GjsIC2crKsuh3uC5w/1MBAkYevTlLPvx8YpHIQVP
IufHdIRTm39Gl+UJWipG/eupT38LvKm8MW/7eCAwUEkOEEsASIOBWBeS0PvLwYUPEIeynZjG379r
L+9dg3CgNYjqER2A6LB/KKG1Wv+W70/VsDSnxvwW3iKy/7ea2XtAo9GOwZKWTzNRw+E8v6gnBrbf
oaE8FW+Dbg10xhoUxTD7nml0K1XrOJyBVE+t7nI5WlMXaQ7hohWRm0mLWgkAGRflx9QnZirCzeFb
knqdy7oa37gzi1sPqfcyhDPYPSpwa4+hhrGOiFaOd9plgNSyA3hr1Ox38Vl4fKu59FujyIueVuUh
lqlYcSuh99EWEfwSwUs6GXCXbY8klQ5B/BIZepwZws9peu57uzR+PyFgWcn94gfk352KOYWPIn8k
c95aHylEzQ3YV39yC8OJpkZcLFdI/NJsb5SeOzj5kxDSoLKwG+4MBsSmIsskYnw1e6x/yf+kpXeg
laAYRzAl7ZiTRWGA/wGAio5r4BQgNBAPSc0KVgIiwJVPZiONLpExKBXRwLzOgRhcWFiPcrSqWI6v
iaABUUfaiFqu5YCSacWC+0RBW8M//fNX4EDoq7IFoeTrdBx+YcVE8TtQ98vm3+fe9tpYZYVuKEp5
5QDpEEvcTDja09D8j63RJNt2zqHA65SQo974yRe9VFhMyx+LmfAYGGoQB97L3H4MW279cYyQ0xbF
RsujPUUCieOXwy3N2KeaD/3zkxJkOkV4lP4dZdUQQ8RstFgwq2patFimimdUQJNGM+nxMw4sKVtJ
C22n8rd5ja0ff643JQQioDd3vPkMDrAADzk6+W08Uh9+S2OlNtnIZxhNjTrzFvwLKMxHaLz88yXI
ZYIsvjYxaOB/ILLqO+PhHTfWZq9eg0CCK4iaVEpC9d1DNUYH1Ry8PWUPISwDEShNvgtTFrgGlzrP
Qrqtwms65ouJ9YNgbFhHHdyYXxrXO8h4oa9k4cUDvNsucvE34AK8JP2w7i61hQuIwL4NmVF1eGfZ
1eaS/fkdAUdKF8Vx8cvXlnFPOBZn61KB97FBp6LuLvv6SCLtbRwS8ElUwmfTAC8erEm3u87HjOHD
V2cy+5tb0yEzL4UwoYfKHADjiIasNN0XEnSg+7MJzT73KhTgWYGi8KJdqvdYXi0/yCv7S/gTNCDk
bQ0U11aUpaq7mpxCr3OEU+uZuuaD+Cs8PIIhUZvheQAM1I29YfEhyykpAV3vKfmekbtXZ9m4BY6i
ZE4wKGKAwysgEzzGI5XPMnNzCdX1lqiNeNQv7H+r1pV1Pqh6bTeI/gAOGX8WRO8aKepNJX7aBwED
/TheJ7CZ3ApRxUOp6T4ghbF8VWgnVrF+4eamt8dZkBdf9V5Atv3s7EV6NDLKCQsJ74h9/eCdOUwM
8rdwAbY2c81SHJglaf4cu5eCfEW96mOixre80q0vwifHJwRPjbiDtf/NcSBhv+MkkIGtCYA2acL5
qGCd4AjCzAaHBl5LvV08Q7ldAwsHqE7LuuCp53VV0U++stM/3kFJGqNbw6nXnUaTn2KVKCU/68eS
lQ67edVC4HUXEZjTz+OOmGMd4kE3twu87TrWohSw2JVcaC2j8zvxgyRrH83/AdL+ZoRCTJ1O0apw
Mo8Il+BvTSEyx/JvomHVqcL+qC2bwSFXWxIrYDQSg5xe7bLFxLetthoET5mJuEICSK+jYWCKLI6B
RqrRqL+LfWX0HhEw/9rmx/0rWnWge6o7tEY71B82ROQoViLSgjOQXNf1ZwMQJqIGwROZOWe3tQ1l
K8Tf+3a7I02HIyEntKKEYZ/0ijHkMBiOqTm7EPk+XDNl3O8Q+7qrdajoLo/MVkxvy8HfZ2ixRPI3
7ODy3mxeU/rjx3ayeayO2wYBelhqKyXNph9LIeRNYaVEwzg0s4lBDvR3O3ccVGLwV/8taek2xdYR
P+l1Ypvts/P+BCum4DgAHDtg0K6E/aNfKW2oBiRAuqQ9i3+PpD5XLg4NgvnP5qPbd5VbDkGz4c+e
Glw1a7TsFxQOFOciAtPTTkUt/VIMfLfGfFh6n0vur+eA35dMljpStvdKPSYNi4HcCD1K9uMOrQjg
IFFpTDMJHoml4iJqYnTRq3fNNrGELjokOX+y2XgPTc0qEQGaAPcbekgP7ECecXEzgMACIJJvNwdr
V+JN8zDDgRWZBtoSFRgMHYwzSKGSWuwHsibB4WjUosgTA2VMT0Ps8O7/KUfjuJzeAlepmRzyqvCI
R3+xWjxin5Eln+0QdQutlaLGouxKhbe1pwujg67JZ++9EvsiCuOA0TSIAHXrrn4x8nT8BizI50m9
H0yqqYJNLJodhP78gY8VyOhJmpZ3hm6d4hy4Z0JNYboEwq/4OdoOsoRS2cjnihHCPFF5W58h++R2
i+CUPs9Y5AeUpmoenMu2KBbbGISWZ4W5mwnwiBV8re3ccBH7ShJsG5ein91toPWCyJVJ5sLB0UWh
B/7CUlQERp2tKmyWbLu0IXsxkR3laCIi3b6H8mW4ytxt1uGJGWK9bxVrA2FzPjfzWwxWFPGDAhZh
fG4mdV0612ljoCbaM+c0oSDszeYmmLdwtbvM34a6ilQYWtZkUAEpzLYPS2AOmCbhvvC0K+IPhrou
dLbmR6ODx3MdA13fWjMUnqa45kP2UijplL3JXSEbewI4e+vPNb3Jx5TFEnjLZcQv4BGwRLJPRhqM
a3TqxFLosqE0h3sFAdL5nwpyX5mY/SyVnPxNr6fni74ssJxbbjVAYiaUHRbcJhgSCkahCn2ZYs0H
CDx1ZqFjwQt6aNYQieMMqMkXrGRYIZMg/h1zyxm8NFzXsNF7maoLlafsLpC2em2RCNDAaWdrULIm
9pAjs+1wywgDghyyLg2bpT+kLQetxSTI+o1QQWHxgRUD2LN2QE+TYbqVn87RGSUVxXzg/BCyY2le
mvMZjLffMneAlAeXXNWHQgRlQUNv/GoxTfeR5fo1LEOfRjJH4t61nNWSGdqZhtovGwi4PwHDcTW1
GhiKpLVU2/kL7CP+bQiSmLw9hVp3EhbT77iMmNNVz8iGxNYdrXYVcDgA1RnW0bRsRgADaQWkYK8h
CkKYx4/Nc5DZtaD1n9+b+kOyTZw+TIcuFfr678JCM9OAL2EM9v53QN+0kdiNhedodduiloA8nhJV
kRWJIyDubdrV0tqQJoypDDsqrjhGDhpBKdhWKKeDBEZNBv/gCrYHz8Hfg/hJlGmflLY34h1mqQuO
nBs4uo0dbvtuKKYQfjyS7V3kg+DwWg2MBW6/ocCIyyLsTF4W8XOAk2t8gYwdrXpRljLzRh4meosI
okU9TCVO024A6MXUF5S3IcfG57lctXnkhvilGwAdT0cQwpYu9DovNmK1+VcrLhCxKM1ObHLALEPP
ub3XXSK1UOUTcgtF51Z3ec9ui+QDBbZcaKSidGloinFSvtc6+uGvGzHoZ7xfeIzPgoL2fe8TYNUV
cNrKjVLBq+BuRmpKp2CdyYHulwxWHuB/r41/9D/pzzQp4Mm/HNBYDkZhrUE+ZH4gNLDUBkNjb5oh
7N93siKrQcKz/WP0qj5WJuWSlYSs7PsYRp3bns4DWFn4g8jK8XKYPdoR+pGtqMUhCAtlTcmNuqT5
DVoCKK/+2aUukhi1dyvEO7rALKaPirsb+FitA2MtUiCCWCQ8+ZjmWDv1PDqrGRte4YjQg+L8nC/H
u5sQm0/a0YNmuo7/wTbacbHc2jloM/H2vTD+6oLswV9Ytx3OaUfUYtp+CB4+c/8SMLAesPziVTiF
NZXpcRTSL2tEj9lnEZkxaKPaie9SPg2LAwxnMHHLiXl/raqNuJ7/XyoCMejm92FbaPskkPG43PWq
KDioFn+jaZktorb3sUAvlEY2coRBZUa8Xc2EtC8IR2h9UUmTJnrtSMhVtaswJBiU/MzvacVPV36/
3yH1vVfiX71gT9q3iYpcV6A3MQVqYnEEP0RaZgzjwdTCwdaKq8M3mMeD2gLR7Ma+hiHAbeK2phGl
+a0NZjtUcIQXx/DkkXOYeSb8HXkxRQu8VERqyevA5H2NgkT7faiOSDAFBnlNIzY1NtU/1fOH6mET
9QW8or/TAExw5V8EWrrXNODwZymKDuLQc6jtEC0RilIMKyU31sl7e76mFgna5Jfc8Mef23Fr5/GI
FGgrYvpLteO/0ciAVmBRHE4ADGWbkAZHxiPhqlazm9t7WdzmR3++175e6gUuHdrYQnGsmdugMoAp
d08DtkYDsA2+gtSVfT1buhGQyLrraCJCUWfq425Jn+OA38yXi5uw9RefGgchi3oEEe0VVVBWidX0
q3vN9nBcz2VSpALTTr+DFjbzZB5pmSBTgqm6Dv2OPWFEGP4IppqWwykqDHPymSQ1izqgYQJlBSCp
RlR8fkVfTWgxUUhTcC7ABk3QmdJicKsWjHQ+8XDtbX1+BojDJDDxGTyxitaeul/XeRtT3YGVOqVi
kpF2658Kdw1/bKHsRDzWF4qv/0MC6Yb3qRFz9NV6u1Uv7l0PQVXqgOfltkWlLsWI/1HsbOUVOR2r
LjDqW/S5NTLY7nJXEEHSBhwqONNSgMvHS5GFOIatTDh2HHNjZxQ727y8upAEn4rHnQzDk9ghw1iw
1VfgrT3k0CX29GOVLb7V6HvDF+Kf63s4gs569689Mkwg6XwRiRHfYXitKgmHq/yOKeuzg24T4bjC
PuzLU6SI07J4OGLWOc9usYSn63OzR1CJ1BTVhy4DLdqmC97CM8RUurzkhPpHYO0kRZI5YIOOmx+q
KYn5OLELZKgTR36T4Eka8wRBN9VULoOIUfUYZxuamW9CnOafRoHpin9u5bFBK5bGfD+IjFDkKzVu
kwK0HaabLTV3WGu2dceG6hTbI8oNlX0C1+C+66evZjO3RlprA2PGNShN0NQNE8vo0UUFNnP+Ynof
cDZucxMLhFsC/nmXPq7pyzDvOJ9UDM/rHmq+w1A+qRZ1ojpnejSExM9nUVgmxdWgiKhYNqqM/qxA
HPyYbv1k/a9Lh3YON2AcCbCv5VSTsIH5lpBjrTwYKgqFNuUyKRMk4jQm3TDtLoQjv+TM9P6WQTfA
GrzyJ5aK9RBiz5gQl9cUDXIqZdJmetlfZNe8dbX0IZrdlhq9KtY4mSp5ja4ftCkZaw0pOaK1RJPk
QwX+O7KkryQ5kUr7tqOsJmRYJjeVuk0VXcVfYvzaTEiKIQG/puw4BjWLJlIyb2avKQAiBR/lx2El
YfCEl9dXFdydRFrPyabnjTmCFbtCPtVDYn48S9WeWIjntzwRE7oyP1oV6FJbwyzAoL3rxCvN06Qz
OJJMghiIhVoozuQsVO9kqAtEmZyucoL0FeFgg04HhEjQ1bACJzmMZtmzhmN3LX2W7O4khNydnnfd
GvTD5gZYOpTcH5pVCTpxajjAvI8LGs0bjf8npoU/hI6i7ljzVQp0AlOafutULv8ZSyZpUMScaFXm
IeVbH+EL9TDDd/HNBvVcf85EYWPGL6t2UrHmWS55RNhF+D8UEMjwoDrhPlhBdOWbymEsqM1OsGpO
nCobP0Pz3/f66b5dWzcErGzYihvcbmTFnX7B/x8budkjylGkhcu+6wTQ9M6z3h0HaPv0jzWdfsw4
OhigLsNaSkKeqZjFudWOROZbOd5pSP2gW/i+YoKzZkkgQooq9AnO9ytSIrVFuGv+IBGsnEOYOvXG
m18jwygw2DIbhkrYcp2Fkrx9+h7KA3o2YBdwdjMAfD29qr/1Jta1dGPYn07tfCD2LpxCwtuD7m1f
wny9k3yt47LoIV61SGOd5PiOFCoQozrC8jB2XH8JXQ9gP8ixlU/HbGmDglc33AY/z7xop4QwWA39
xSCPhqsiFcFjf07irFRoi4aIaRYh0Sj71e9ZJlkF4Vm5mUIKB4BVFTLg8SH0ikCjYN4cjGfl2MSm
/Hbj4uSnwcAoU2bavULCX7vWuePT54x2gjOYGuPzBsUnRKJAk5WPN1yHOGChMSihJHO0tsQhfVOf
sCF5y2mZZtk2lHzOwvisQZo22eWwSCTqTU4TnKcOFzvOY4snKscEKSYVPBzd8lJTFe7Ip6ueRdYm
nRu7i4mmCiilpNj6DH1XpahHikFAK82LFF8T/d+3jX+VCkfYcVLv4OZMcy1fm2EJOscg04hcYhNJ
yTOaRqCzb8n3mYDQJd9FZnXayo0X+gf1MSiLC3V84bX+gDv/vlGBWNUO4eTpc712YFuZgtb48uUe
5R+wxZc1g/8TGZmGc9S43FYQh0ToojNuEtO2d7tN+x+Wqyf8Y7vS4mSJR0NujW5mqL8NNtz8A2LC
PLGdTLZB5qnnsEJutuDoEZOtDRfZTcch1eGOFuGQGgL1K2yHz9Q5xuyqim9dj6S1X8GWtusWxRM4
m7gvsC/ZlQgYF9QA9M+i83Xq2FgkveoD35pHKlSXXABlwHZOfK/7xjbM2GWucgzihDf52N0pUqKC
9Hl235n8ZqZbCMdOF6BRwpRaEiwZSjciLJ+dME+lUXBbv6+nMU+55jFTj3hMK+1p1hxnjVRZTbfa
P43oxHiYzg8vcdM5eq87TT5vsoX9vPf7p9TWU/f0EO8I9qZOJDm+3ip5C3SuSztDx8mnATAKqf+9
4poBi/g1ypv+d0Z01eDBwbDvp6O551qcIgONLOb18csjXunZJBSYHXcKdEZx/JFGUmHeNVYt8ags
RdluiqFeZWp2RLHhyUYCp4F3s1F1HTXW6/atXFEKqTpDXXe5PQLU7cVuoAvR91rRJzXbvFPGlThX
0THRRum2kDH7Pj6YkShcZIwoZIRsDCPsK+cFzvEBqa1tdrT99I3QG+d9idFJN4YFiFNoh5qUNLxZ
WIT0TYiMn+3JWsJFaEy/EWoDLtdFQYcMSFFpJxjhwUa6KQuua8+/63F0E4znNvRYgaADt60hlEvC
gU80QRQu7AxsuN285xKWtSe6FV+/UV5/JDtCm+dc3p8P+yHxueq5Fno6Xd+lYTvXFxeof/oL3DUj
N3aP0UPzwqFXixy7r1NYF2dQQzYeobLXQHCoEyx/ryERWAXzdb58ju3m40hO0ccPzWWWckVqm4YA
tnbJbdJsBcVtzl8WEbs3OOaEFGx8COHbAj48f6T+KIb0H/9hFOpeunl8t5CHF7ebcqWO3EihxQSf
RQwi41Di0xLoY5WGQrnrsLq2lRyqnFlC++DgxIadWUutPpK0bvr8K8fi7GMXM/eqiNzK6GxxTzQH
0GjzXY7UkC4I3u9LmTmxqLKAzIRGqBEID1vxkY1VAJT1ZfGDcnX7joBv9kVCo9PLrzNFcV+XMDd7
41vPxnqD/fEsyB+i1uYz/50YBlOb8HxbL/o6fnbxu64xtfMIgh+zbBclf4w7jKMHeDU50OIrMIDi
JTHX7N9ipU4/2junvihwIFimUh8P1sTUVxwgjzEzq9aQmKFVMb6T8c+0fgI4WGLumLohQtOw6jOE
yschGw2+abdaWlZvYzE5ecUrs0oFBZ+Alm9bqZYYfObeB59EOB1I4+aSWQisT6bF9+kCezCYivXT
wY7kTsH+IvImhXhC9tjYHpLy1RHhRL2A1ACa1G5Tm9502U/GnGp7hPUKlWRvXm8HsiZv6alFPbbG
f0hepvANXRUbVNsvDR1nCmf3aNinw3VuSsd9uSTRxjSfSNf+gXLeNSL4UmIVVWJGDl3RNC6AgnKU
0oI6rv8yp+hGvk8dlpbRZedif3EkHtjiyVgKGLerRKEYRZHR+O8+j81k6kxYucv435NPFgvCeyQQ
FtgLEyq+AYEk6F47bt1UUx4unniZ4klmRCusVOGjOfoZsY8OF20Wov8m3MjXJr/pTD+uOSPyroBI
i/9xQ2g/5j1raE9btEY9uaqEaWABTMLhmCbHszD74a7UzP94VcnBvBl3TCmP3cfNBrYDycdGH7Q7
zRKPeCX0WEW+KMxNvRrzJl56K2g8KUWlrd4MSVbUwDu+opSIXy1tWL58jILiPlFcCIyGBWuFAd6q
HVvikNV0jSc5XN4ovBr4xrCazGQcCUMiSjYOsGcNR0t138c9mwGBluFtEpnYvyrCnjv7MxWr/TGe
WauxAugAtdLho3JI8NSC18LM2UHJ7kEoSlvJh/X0EA+AcUdWLPT97KycjREkoe/HCIAUYMgEgAvf
0sR8BycLLI8pi2hkv9B+waaBbtGGyfgXLAzD8ddcfm7/nuRyq2eY2I78xOl2sp1FxzSOCvNsPq4O
v1NxkKrIOUm4VBtghk1Inhn0tkwsHP2js+zbDUsYqKX8VQ3glD0YeAUaDB3VAitYBa49UP+1VDk4
Rl0pw7CQ7sKG/0IsssXwvH6+TfCE61ExBamURiJAYJH7vKJYIyKIBiojw1DlQ20n9tlz7Fw8p286
TMh5lnlpPAw8dz8XGkFOw4lro/BgK8KSZixQ9gxypGSjOjGx35bOQtOr+IzRoAn9HnpT/enIEuGH
4Hax1qVOP7kP6G6yyCLaWnADGhvXNNKBrzrvdAFOrBgdQ2StpTlMt112LtAIFkvS1zTr9T917fB+
3RaU5/yCHbXo2izoYX4nqKN+ZYFvf4/ZvNV9Hxa0SzTxMRyCYwU3cAHzSdcAZL8t7+ThDpnV1b3V
VIeYGYZ84GIQxgphsEzcAEqB521Ves2tw+SgSQOpfsjoQg2FW9M/74HL0Dhh4aWv1IvFBCw8MmNb
om82UwsvSr87z9uKwLIP6zz36A818Rq/SbE53NXDV1vlbxFWyvBWFOIjJ3O6wywDngJWF++mPXvr
nwm1PtOgJ/gUxHQkJb26Tv5Cbl2+4yAzKbr/YNlcNpuV+2jzB33Gz15mUCBRWU0hJ8OkpGRoRtwF
3mhecle5pGQxOaG/axYZ7Ht8Xz9rcWrXzdsq87JRCgQNB/0CZngpwrgvx4mw2M0JbUBQNDSvzIzR
GW5d6/SvvnBbFP/G+omyU+AY32P2xQcjvXpS9QrxL1I9QIgXuloN/THdIYnJF1BE/NL5naP9xvhE
BZ/0fsdOUv9Ha4Jh9z2CM8sZ4jLHk9IGBPYn0W+0qjTsY11fs1XLQ9o4AjklWCmjHfokF2cCFbgO
M2PTbzamswMG9LYStTrNL8ZUPkiFhGh2m4utY03niYq3rNex20cdQrOD/yQx0cLEaF0tBVtOQ9tl
y79YyJnLI8McXvfnV9IFEG9JGP2jfXmwn1b6mGJICKY5gZ/Ip5QtBwJcqA0+B8Wi/O3ZaB1IskMM
LLa4JzDIUnk19pwiH/nq1+Cr2WS1bLxXLtLXN6BVrU9kIwPTNU6ObG8MACmiZuoLkUOQ8MvjJP2l
Nk+D2NhG4Kb1VwKATqnKtrnHZ281rS6WHX12jvrg82bfbHmTrSa3vIEjIsCrzBxM564wlHuDoNKe
5+kVa6sm8OnoKhbJGrOIz7xfWXQzlsEX80DwdtWH+YsR3glypPa6+JqvlViLdDLiy672qNX+lOU8
8GqOjz9jUxa0irp/7FwFJi1FVk6IJ/hb9D6OpuPfpmV6hN2X4MWDbdbrcaoCKg4l1Mr9rgmONH5J
IKOj7ZXndxYD3oppWTmmAdkc1Lg3oLF6uqto93luAkDWfRUOyLcF7egdxDleoDFlyD4dIqABn0x9
i3jSwZOEPBPCOpnGE0H++auk543vHRoruCOXi28AlBKlRcHfgv36RDAggC4o2aDSAcZ28+zBseXl
ykPnDBsnsSPDHDhigm8c+nfub0KU879rzmRdLldyl1c8nL7ubBTONTqq1nxerXWQii7HC+24vut9
UAKbZ3vQxi/HgKGUU1z4o9EF6tFCPssmpiV0s+Dt5c0lP9BHdxMDTsiBSbyaAvWW0n2FwUxakHiu
ioGdm9g5vLeqRfnd687ewrHdFjYjiWI/N+ac89GafrpKpUPfrFhACflv9dMgR0gwcu2LaBDSZ6Fm
3Vq3hRCymEhggvAJ4KT6KlDCMC5ZYJIdud8369mVM9Cshn4+nKkte32LILgLmKgyHeZO+dYQbUAp
R0D8KdL1sSaMb1s2JJQHVMtVZqCuAycGky9Nl2pLxS3/ajOXfZtouaM/hwUK7MFOwdFIoz1mKQdI
deUoaciKa0CjGySAuEZhYil6zz46HGIljqBA/xB1m2LzXuan6joNbnyQjLcjtsYcqok4TkfOq58v
A3+GrqeVJy+Z/32iJf8SYy4tX07rq0I9uhBO8Ui49uVyd6YlTB+RsLCdopT2xsMZhvL/C4S+XFCm
tSBrWxo5Lu5OsN6tKMt2Ekc1ZCe2GI+PKpZTyX4O1/ZmotdYV4XyIywoEKRGWXqudRoZqNPX9QCS
tCr3F2s1J+J5A7yXEbeKeNECYz21TkwOKCH/DG8wak+9wzlEgJDP0boBnJ4nxWQ1eS9BWv/Fw7pw
dCCT/HJPZLC6M93U/CCDjf1P7FbdS2QRCHabWD/2Qz6y0x/2EeX/S0+6CAXlCv9j04gTLkoRFXGy
qgIsdmGP0qRm/WuT++5wzsKkASDmNK5fVpuL7ju2MS+AISfyAwHsUkuFfyRiWZ1irp0NrOCheUHS
rOT+cP9UYHRreWS1Zcxbk8g8J9ru8WGcz+IZJLttrh+bW6n15duUTJiP+WW1vYiSg3jB4sPvNVeB
otH3vr8hY7AIFjwkflUtZLf+iyz4doAlbH0dDKlP4YjR8na7DwwVbTlTUEyeTq9Fsq/iPyWJNxDf
tbktKldIUnbl78pyjCnzrujLR7dcRqjOJy7o/R6CWChLkVIOaFl+j94rpVzbklKjG4yGsS2AhXUo
a844ipvMEFWs5gecxkByTnJhYyXZcBWJAfAL5ZEtsBPK5TdSWMC/ya9RIp843sts3Ykd8b/tWLXk
p2Y2HKvzOYqUeaLF/hrMgJSz5D/tW3zp7f50IP9ASEhtg01JiZq3qvGBP606InWRAkZEx2e9euVC
5+r32QBvnTKtetQpqOlgABy67rHhbn1cof8YFFfwtXp5qddcGfRulxymYFqRq4R8d2ICZ+MWrE/c
joVH9G/r20wtGCfPXrj67bO7YQdn4TUeYJIIDpkFJ8KoF4OtKi3vdja046ufu0j+iQgwVLdJbHZB
lzmdFVHKWPeQKQtaqts9CtS1eu6Bmk/mRFCRB3vTZSQdSVt+Q9tWm19qI7N0DfVR/llmWqdazTme
Z5/fcckygqXrZxce70BzytFHawSrPwxmTA4MXPWz29n5WHA0L2LlpnTZjcifsFrekrPijit00Q5G
4uLG0AVNWmPsvs/HYWU9pHYkgvnWMcgzYK0D2JfQ3mFri/o5+heBuBiuywMfbUEt/gvhR/O+Vw9F
nI3S+w9seD88MBOlSd6AmDBAe8QLbw8WBW8Vc5pQJHqvJBhIJZD806TiiOw3MYnrjQMeFJtyvGjs
q/E1Bg7wiL0pyjxo2Lh6Yp0qwCRh3U7MmngYrJAGucEAedryjO/F901bs4xzNLDthFxXzgqc7roO
sb4GWT/cTCnx4r7Bn3s8mVY75AdvUOH0eTRF9ZjbXJMSSMF3yJAawOS0d7IQ0UXdl7Ec6MbVJCfi
0WhBFEkrqYmSn8QbGtb55veCePS3KOtzgrLDDh3lmMJaVOZt5cWLULT/rTw0fnhkjFy5W+umU3Mj
TIZKUUoSodFE7i2HIoATCEJZYdNmDeyLhqAnJVCSb3ypp0qlynRpcHV/Wuxum9CIXO2ckviW1A44
MhYdhBYAeyU3W7k0Dx9/2aVyUq1B9ducFsGQKysZZ0mEKX20hl0kOPTyvJrdpHSgNTF+EBb4E3VK
dvuhtvQ22THuajBeKGPFx2vx2BKiJIK3qhc/mx6tqho1Ic25yaibKb4X8eyrpC7Ze8rXoSDhL8vt
gozopG0tQbPYKPDBepKIR3qVKAAHm6dDCg3xN3kd2I5sqV0Ll27icI82TUZxCOrnvs2lj90Tlpu9
BU/7wFcoxg8tWAyZO5QFMVi7ZG+1gzcHEtKcAJ+7b3myNaEufaIJxIaeA7zK6fecKVN1HmR7aD7w
7g7UM6aKTGu0/4cRiPoD3KRg5ILz6TCJvXNeQeMGN8qqP+2G/7rEiLFi7ov0MZFOKRF39f7b9qou
lH9VBmFbkw3eQF2ia3hmyRHsSL81Vzgr2Huug7tu4Rp80WXp3Dg3ChdsD+hBr/xydHBLLRJ2Q0Ce
hPr6L07N2onnbp+JnFss04LjpV2gwwYHv6EtCSpQZIdbvxTZQ6qU2eGcqc6az7jn7VMDPx+Ew2Jc
75YJwLfUv1JXOlfwsrMx3mCFRNnjX54cwVi0xmN9+J6lgrJCLoUhRDLcKGLDzlviufbMXwFuEPPu
RzLAnnbHJIvVbLJ2+WcCWahxmRtKS1JtFjLX0x8ZBLEFzKd9TAjC8kepM1dJY6EQDoaUQsAiCQ7Z
V/94etGvCrkPfM1S81tUJyzgye1Go9P6LAVeEBZcpZPWL4L3PeR3nUFRm/LuhoZIwYkYoByDCxJE
F+alyO6EevpxardDEGWsIAle5G3hQmvrM8hFIj3bJl9eiVwCMCUVDPt9bfNgnOFxKGi7gt2cp41l
hNPqeZ9Pk5Ha6K6f9xyJwIj8OcHSZpfPy84uIiHjan85C2pzfw524zo+9XmCDbCUmmN0j3bs1IhQ
O1ILGq3wu6S11kTXWqxwe9xI8+UjtC2Ko36fJ3HML66ChRrRSULDOYTQJXMyeDSoGBKuMQSqtEo6
XlMnGMImkDFDkyEdZaf5IKExs3R1l8lkX4n3TGKLVmC/CnqPKl9UxIewfTNw9RhsK+QpRgqO64jI
Hh+B9Ohme9d1C3RqafNrwE+EYM5n7H5MwncZ4c0ycehKpn5yM83O3Opb/+ygHLhj30zEXwSfpDuB
6MVBPjEawHKi48WMKC6tuksf521sv6jsVO9ZlSyZNXcnyeKK4A9QZekzZ+nC32/qRj0a6wFoMRCL
KIo6Gj88hftLKNN8QLV6iIloc5KivtsPKGbBU6O8g0yYDNYeM8DiflapADA91yEOgGRgBHYoBHCe
Zzdxe4T50vJ9k3mgwGgX53eQdEBFQpZRTzLeXKTKuZ1h5PPYD00kWlCrieRsjBH7n9e3uBpKpRp0
W/F6g20APKijRjNsoo5L2TVRJsLvTw9pYN0760QTjBrmhgBiXaRmhLNobvNIokLCi2sqHOSuQLgi
T+x3ETv9hfCNPtbL6wX0NgCam1mQn1vnMiPmjmhNt7gMg9RN5ZaMccojXLLTF8ashgazMOI380fb
FeGqdP2+5ffSQArvUzzAD861SLauNq75Ek8mrAMUMN5xpTAwaCTRD2oZk55r0KkHP6vOwLmtb2Rx
34gzNFptAqfAlW8Kq6xCIY4j696H8N7QjajExWlz1FNIo7Z3HVpnsnS3M+L1UfrF7AtzdHg1sFPE
MEK828BTj91Z5NkIvsEEYUfqD7RBidbL/q4vTuy4uEo/OkHENKJCqlP4R5kO6BVVFxg97iE8mKiU
zvy001Vm+VE/l0i+sKpJ+IAV3wS1u3OjR1Y+7XTcIyJiGu8DYTWDmY8hRn26BSUmHbupn7FSaGBq
LN0Z0ucGrWJPVOiEPlAsXt85/RyrqJMq2Kl1RRSRm5ElL9wjUzblUpP5XCS9JntNGD0XfsE/2rXr
Dp+omTY+BmX7kfUj/cWGRkNkfj7lXlWcdNg4YVca4yvj0wdgzknkl9saNalXs7W9ni7Cz8FWJH0V
3GphBZUH9nI6M/WiB0V1MBQeGxMAQNZzmLd4bmvWUj5Pm0K0HX7biHIBnOsMeLIi/yhGBDr+IM3A
bCWTpdOBi4qIwW4a4ferIHrkKlXcE0WaivehTN58VrDRn2Fka5encoooEaF+KRiwdg3aMHuDwh4x
RJ1XiWOwY3azMrdHeQKRZTdW5QJLdMCygZWqM8IntEJHagkBXw9v1CR5L5+C3D9KJ+l/jIIQ2MIK
P+Z12Azq1ZIZK9g4WlrtTUpYVWarerPJxmtrsd/rfWk7ndwgpQRyzB5kdrhewBbDEehdMFp8Zo+2
h6PzEhEoi77R5hr5x1hHiXiAwmG4zO5UmS8pBAozI2kBDZuBwlevXojcFewXirUK4uBSoN02/kz3
6j+cHV2uVsrH7F34bL+JCHclGOYdnWG+9kR0jYxowp5gyXRC76PBErRtGBfU8enZo5g40K4nO+B7
4tMLOL57gosXNKUjxvK3GzgkuX+dCvSuPusV68DaL3mUUu5J2cXf6PsnWE04gse+ExTlH9pFQmSr
nNXDGvg0XGfQJzkfsiPiDDgwKqMPimt49QfrIlIpksPYFCu8hpGPcwbNTdd7do721kw0FyaMJoda
qm6jyLq76YCeYi4L+79xmCqF8bSxyxDyqB1zag9VbrmhN90/MZDi7R/KDg7uflJNnMilOH2oh8tQ
aN8kxQzENLx5xX3u+1SzrsBMvt3X7tbsS/v42LHat1WNSu1yX9yVFsNoQHOAy+ZuPriYwxorRah7
ozLib/uCPn07myoc8bXuPRf1tiK3XhnT4ZEXSxmy+6YwibNo3DNwKqDpV170VLKAhpnQf6GiXLGm
4iERIrKr9mAgd8t/GnKARN0t+MDWXQ9k70INDodcjQvg18nE2lPmNgo2G8GeylBEJCcoM3pbjdgQ
dCm580Lhep5zWO4UEbwTSX/51fJ4N7LocBWoC46Z4OcJqtJPGfqxodDHAJnTORufgo7T6tpX97ca
TEfEPcQrOvng90cygjF7CtwvavTuZsRzF7/KB6ix4YNfJbjaSMh9djbNDt+8QMXgKTFvO8KZWyZv
lwGcxQKB5M+RhqKoHU428bjBLEPjrvpTjrG+O+uD/FHyzfTuUot1s85lJ7gMTwH0ynqkzoXE0/o9
ubwCE5MTImSDm+7xC+EPBC1VQGdK8wEjqS5cpmGan2oZgjgHM38kGqN5fm9owQes3ZEC9rPJLPjO
yiJhFd5ReMK+0OrCpDh0SZWX7MFWg4JPnn0YerGyy3cKvpcjd2d6OPggWwymawdAq+9EtZJEJ/yr
4fNhAo3w+hCwuYRpOklpDwdjYbJ7krsijqAaJk7HyG9PWLlxdjKYW14VCqiiwvGlNj2P5i3gMlQ0
OHD/bbsAK1tLY6d5EkqxplQs0eI0Mu2G7htRgya07K9HkqRO3d4jFLvJ2oHUCv5iTos233YJaA1I
fkQiSUkC3rOtZSpctfpDkdb9ZgQ0jfkvp2pj8eOEAk4MJipCTM+C2fV/noTFqx2qRTxyna2hgIcv
HLSSkGLpr+Ch4X9C90fr6iUXMTlymjexiTV2glSCrtIlBZLgBndp+DJRL786tEuqkJtr1U9chZHr
IKYiN4C12DhPLOnACRvTA1egZ9CF4eeYyw1pvhFbzjq9vUs/YSRVm64fjCvVfJQ3/woS/jGGDuLM
HQCaWI4m2rTVtRTyqga4icOW26rgF7L0/nsCdKXEhI/0qUWluuvn1WxPW7ifmMXg2xRrKq1q4WXr
tknx2YeqSf4sVxo122kaoZK4dbCGiuwrRdLrndHCUs6LitEIgZtuE6tkpBVHMAYwXDkQhFGiaybx
83Lzkillqaf9Z9WU6XObw4loJpcFgtq4iscXxodZj6LeQ10yRTKzgSKuTSNbt9wu5Hgss5qt7Atj
h8RwvTT1ErIC6kZQ/qTxAtal9XuY0lUo0VMMe89q/hpvQrkElA9TGRgPwdTvDvE1N6b4V2k79iJ9
/WCshHS1cCe48d2f4A4HRwKUYkLOgIJmf/lB0JLZ1jf4qETBnjrAL8JlD520bsgZC+J9fMD/m46H
SgQNrhlR78IdePHGkpU8FyoerEOhU9pRrOtPDxo+Jh1nMyAvkbmcFa0KtnOtQ58e37X3J4Cd6kBn
vaj7Wu3OOv3YdLW1g5q2kDRoDCoUbuIvtZGlkM/wV9IoU9OZD+49uyqleI7fp0Di2C0ime4BeLh3
R1pT9hltsW545t9mnC7n05loYO8MhpO+PmNPNC3Ua17KjpaSQh5BaJET0q6ELC9EIO+EnTCnZpsu
FhkSnYgqfJZy6eRpWROVir52w7VzNgFEdndu4FILGEy3SyJr4wavoyzFkuxhTEyypWJinlkEjjL7
KD125JOJgo1nOxsY/y9/l/If8+++4HnKMPdspCCIcNVlJ9x5wKF4xz76o/By1rB5vPCOZppHVj0h
ZpUfTY1S3BE9zsGGfYoNaHeLkgGJ4SaM9lBWPl042kzWf2lw4/qYIL1BOGlRxVIwtEjXWC0p9Tbk
ybONnXlIi11xHzzVqBLcqAl6v3v0wWsQWPaCcx3zkkXZGPPfWHLGsXrwyi8wMWe7ZZt4YwzvVE+P
brlORx+QsuF5plPXiSkYgCgh6bZ3y3ZmHYGMN7JKngH0lHuf7eslPh111Ot1aUKKxEqnKlovxGql
4b0HtwcrfW2vjvxmHlAfzrjfbUMwCFydj1+RUEViG5JVvJkSCj+wUSRm0Rf5Y/i7yGcctoIAdOZK
pfaRhrk9ulsnY42feQkZlmYbw/FstLxPmGDQtirATbuBvZ8nsyEXPnJYgw9GBW83uKHWSaMIcco2
IRftUosXbAE/seuGWj36AiaKcALp01mE9hBDMSRq6LnHSn/3srwsXbwV91kyCLWu9zAtDe78Ic9L
qWfSDirc4v3uXzZ8YKRfUqZ3Re+2bYxdJBDNEBYimujBmvKaNzsA8TxTc9eIkCsAw05ZUyIAPhoo
TT2rbJrCqpm7QYrj37JNTEqLDlUS+kxmNAiCEs+N8rvYBSN9d+EdEuLUgNCG2i6LVu/SUTzz0S7D
PZ+HQhfABTTKPMWD2KskKYl6TB53aNi5N3YNP9LCrzyZGeICgjaAECL2d25ds9Kcby0V8IwWuW08
fjy7hvar8aonbm6yt2Nr1m6l38SF7FWt5/2cChVShhuoA8yJpvEmIkJ8H9k0byIDoBRy9LfxPt6P
z7PotkJ2tAWlDyQ/1vNMzCHi+hOHiC3ZFys14EYmU6RbJBfBonLDDe9DfaVMvX96h6ImEPcULVFv
JAQYOZoFEA+u126GZp0WcVI+Pd83Grxs48ae5VDzJZHbDCEJz68gGRhmVTGnD6lP6Y1W7QSL8eHY
YHn7OdQ5fBIkONeA4FdO/A7obZGjNmWWvipPK1jAce8d8PVNAxSG9n4zTmzCb/60WOnfxYRPx6Kj
WEK4P1qWr+8aSr09rzas5QIUSaliVA/LvXRU1BjmiCqgf96rmzzx261QH5ogw+4keRzkwvF+07DY
ZKqmnx0cfcQorY1R3eDUHpVzFeKlJyzQ1nbmwIhS4B9Rq5792jVlBgjeYaNSPz0JDMHlpi4+oZ25
lZErPWz15cQk67E+qQKY5jHi96hIG5GrhxrmK2s5NoRTAohP6redJzv/RkRo99asSrw84J3KCTkC
py6RgBbTepAecUkkzl/TLmxltaZHl0IU8iLEA+u4nX5bmuE8ZfmDD+U7i9sCoQtUi5pRSA9XWLke
2AAxXb8xENTwU3hUp+dPFYv3e+i78C2vQZQFN6IYQ2ohRnx7kOXEc0Get8P1emvsxdDUkiQiUfjD
5w6AiT2dbiGOFzvidwPL1oEZdkbweJiJ+ahPP30dF4kq5PY+7zjJVG0kZWeUWGgOpHZyRjAe9bN0
gkwXfZpYWZJDG6MHs/Ss7yJUUgLk3VmRWZXdJ7v+csKCYbBgD4pagKAFhf1ihD83Pef7oOoYc74V
h+ry0QCHg5xEYeIfONOpiaLz2PZatvCC7S2cSbvz93rCvDZfCFBN8g0x/7/5A1dkHouZMAKUhL+Z
4jRoIBIbvtFj8khHTitzPuUbPlKcCrs5qUWGjBKpKNOA+jjveIRRzHkKH3mDxmbbL6WLFjPlccfs
Vp/ZifWZkCOgDYUywlIs1AlqomGrTLbXm56Mf1pr+CWH86jj+nWjfdlQck5OqnP2Qu0T9uEapoLe
SGuRR1d0dMDqRwVdIt8EuqO80wSF54LhJ1L4u3UMRNBfXZuAH0EK9NVCYE+webVrvXYN1oOBv+Cx
Exq0aE2a67sFHnK8EqlEtxCBkxDSkyp6ajFrc4JCb6IKN3ytD2MxvX8C5WXLLECW9oZttEOSxd80
1zzGNF8jYZZaowyPB5ABEmizrvgw1yNS8dL1y170njQ3tjI+fje87FJz5MHr45zsjLYHdlhO3rwH
p/5f3W2JdnrsmM42Y0c17v48nNgiXMe+KrXQBG7Y/yd37aaGeTQ4YjV+T5YO1jaq2A/9gOOwQ7R1
Iw7QQ3hjPKA56mFRJhGo6pF9LBEBFOpImbUilfw1goMR4IB74JqeyPmHFvqZ7g1FFslEtkcSvgg3
NJCwTBdWjjePcTCvuGmYVNEQ6YyQ+mLW4OykLvAz3TMFvqTJDvQY6DSizqhy2KrX3JjK0gyXNBv8
TPZTTf8k5DuvVwq6cy1L9ITevaxgaVy0y97UzgpI8XMWsMzue9vcU3wBt5XMHz0GwvKZ9WHOXnWD
RuWEhwBO0KSgL3hDuGztXdqdPMhq3KGXN66XAY7J2G1tZPmykfUtGrubrbP63mpHvF+Vm1MMDVJ0
b/XL7q7p4Oc6TscxqNmdCpovJoync/WHQX4ecmcF1odZit0EL5ovyctmhQA8TzmLAr0bFoKpmhhN
yPYojhJbaJ/1iRUsVd08PMWFlf9aAkQJ0oQRNdqFOAnEgyHoqmlG7NH/24Q65fve/Nn+woPmMU8r
8eUJXj3a8Qm/02E8r9ET8OrKWoeL+CnR1deMgjc98G6VnTCEhml+M3cw+H8WFmRKzpdMvwxRIc1Z
RDYcYXEf/V2toVp5k0obJJcvH+eXYN5HyAApqds+fwqTrqiXPVDXPDQ3ILFX+ajOS4NGXiOUU9rW
SDStfzvQpYTgDFB+A1tJ5XoqnFkj8+lCWy2rH2uD39bd7AVOxKBEVCzQzArBG0CiFs0CFE5rqD76
DRSq0iuxJo0rzqtbqnMP5TmXsut+r7Ku9Z8IUxElARLk4/WFBrMXJrZo8MMEWciM8aGuc6DmSWZQ
VxPOIYPlVpAInlkOWu5UVDF9ftY7JpbfES3LtJuuBt8VcfFODGwhJuCsHae6VSiN4L36PpsOjy6i
UX+LwVnGGofQTCn6CEx/M6gfxPz7bw4bXRiQxn2mORC1oqRlj4BQxYoAD8562Cm9FumnbqP1F3Q+
/+8YljeQzIn4qq/YFKotmd1zztjq7AXEqJINrKiLGzPxpOqU352WUrKZ1O9pPS1Ojkumcygv+b+a
T8/uNga6XtfvDSjzOb0hO/LvphT1YqPjZDIZ6/kLuo9nlrS3+6nguAGfywqt0TJHnfpl4YTggeO8
UDykYrbs/x9XP9OahQAZOu5L/URbofVPNzCNkt013laWtAm3SFL5QUXOT7OVbWK44WwcsrCo9yng
4X5lBu6ZZ1XJuMfB3W0FzQsnOjybE38vHj3Nk8ZtoLmcTI0eQmSCrQlmC/dVkFPnve2zo66fbmLq
4OJaRZzADfd9SX9EErQaxScJeJYd4oLZv0G1ckmYYS9f+4CM0211g+GP/YOBAMCOWfyvTUs6z00R
d+uwGO358xUySVzNg7SlG8msBUMjXR7IEsM48RT2BSNAICKTlYFQknmiF3yzvnCjxRl/NDUTGKIq
WBxEbWSEaMNISItHIs36YBc/ZTZpFQjSh8cyGH7pCcM8zBySbxFSXhB22Tnlio9oQy1vY6sEg+ST
Ki0OG/U1WzzjSFbjwsTBaAFr10agf/Xygm6VxsZGsPkMp7EHgOE8AQ75dYL9pUjvb+L061rBprXk
uBlG8KpTk8/pfvGq+qnwG8mMXEiTqAn6ImVfQh6oRGuSxTwfIPlkuLkRp6DRrMCFY4ait3Ad9qcQ
Ap59XFgqw0AqL2dq/6QTdXuhJLTCAKVVm/a2CR7jkUnYlZl5kztmHoHAna01zfi+BKG9hDlzhxRt
F54WPAepAW/tFIIrk++sbquFghYvFT9rvgIvufFxXX6X/utX1tM5rknqRYdqcjfPS2mmbFpTwGxL
djJuwIbi2Rv4/fkm8B0x1Bb//aULUq0QM9u/8r93byKX1wa3RNowmbsRT/CYbkdx1myX4DFRjMSJ
nW/36/sAawTjrnhTCAhem6TVcPQvKm7XoL0LxokecdaLowACvCl9epYJmLChhcCTatnyNfi8tL5H
0KOoZjLckeMYzdv7o9ZzYBtNntgKMzTb9yKeI0+HcLa4Cd1fkv5qf8wlIaT4iaBm2ufqDj+DuNp3
XoJoLOnjJBklJH6drdhEhHA7SVl7UHBzJ4qmUykxhlUqRb5QA9kFvWuHT8z1704xuK7DqGiB3Rqc
PsXLMz84Uxai+3ZdBVBdZQyA2yVaF9ZpOODu/fnIw94WVHRSKnBy6LlyqvukJnbQ1Bg4ANlNZPUq
NJ3BpRhtuD9lkxm+kqR4rEJDnqEvUiAc4/OqWrrchIqyfsmgBS1FnI5J+dAesiS8dXFFIeq6W0eh
aeUVME/OgQvX/2pjmIISaVG5o+3/eu3uFliuDVWApTBEc/vvj6SHuponc3RsSjRGSlH4T58CsiTX
snx6Y1NQrX3nXKcZQU00DDWoyR2tTEjjhZJbqcUUg+9U6RQ/YLYFpDvy6Dsv4HnjHlGgAA/lkj2P
XCIAduAxJx9irO8mOX7xAHGO9HESKz7NxdhbpPxJbCkAxDmxUVkTNpByGapz+H2kKFEp0bnupr8C
xYqfKyxcfvuBszZotQpnuDQVk6XcdCM/12qee0I+qV1DLgEcJhgkPvys9OzhASttEkYttl39zZto
ccBgWZeUDdJR4SnIZ2trTOAeVfa9VkcMVsBTUUJ6OkVMv8DuSkdBsq2PDsFU0IG+H7Mp4cTNV7ja
BloWh6pvGS7P1lBTFTMgmwkq7TXK6ogSWXckkmPF57MfNeukdqaW15FAryJQ5awLrf/ihYMwxfcZ
mJb+gmgZnpLiKukLw4VuZ7ekSX5HAIDYLsdrqFx8At4SPyOhk4XpDMYhLTxBHJVkGKItfju2gVrC
6OIEMYX6tk9Fuv+JyPnIHBOmuT1EXJIFj5CT6tE850Kc2UKs2Ni34kDUQCjUS78p3izl73jg5Lcw
D5hqT5qJt4/henZWusPczkv5l+gFAea6x+SkG4i+I3kCXvleyRqL7DBDd06rIRA1x8r7Mga08YGJ
vWeEW6RuTc1ZPibC8AAGrCPMS2ppirwgu6izOERTgdglzsXB5L1Baw014yTJHwl/JMvLnUAg9Egi
G7EPOmTsPF1Ksxjnc/yUqsQPg9n6bRiVJTpHD/UY+4nvXosYG+5UZ81PO9Lqwy1N2AWsGbDwyiqs
7vyKyN5tfHsonK0k7RLnMnKzKvO/E/3mmJuJnT47523J7FR1giDbPbTQqXoWQl8HTF1ZdS7Jy5mv
1d/cugbcrYhWgZ6cb2dHmMIXHDdTARzDpvJjzd2AhWhzSZvar8XWtS6RBtyb7yIoy5Sj430fdwpL
H78kEV6IJBASKYzDJGweODx5n96X3hi7dd9n2sN30DEXKuepIO+8rieQ3mGSXXHw/4ztkH9kyAhb
udSzmmJuz2eQLvWKQCTZOd2P1CfDi4WtrqSO3p8JvRuXz6M/JUX5Di341C3pVXVdHQQrD3aNf6L9
M5mB5jfpYZxL3eBdL0qdHEgUEsRB/f6scyDmPAv6WQ7QqojZTMYWAfZLDsFafs4w07X41Jdi3/La
AVW5nBGCmKdwc3pJmjC6s4NuLaJiOhAVowHNBaxco1p7skQcvVKJWy3qjug5L8y+QajHLYEu/Jf/
FTEnvtsb+IiC1keyi2L4yf98U50rdzmGnB+JQ7tJrfolRBOJ97ykHnlpk4HWAr2mAFVcRKbCscXG
bxSXxOuDyzuGcf2p8nxsw0fYLGMxwxZTmEgXdoGN69jeHJ1CIyY7G4pvd+OY3MGf/1c5Tcw32xY3
uhRzsWjTqGDaevPQ6/ahTHOHAUmoKOxY4fs5aYnObZU7RuE8rc5X/LD9I9AdTx2cs3NQGJBH6WcC
Num3Oas7kbPSPfWSa8U/uk8WTxAhqV4cBbj5/0yl08IAkp/oYrI5V0qynCpgeg34uP2J9ci6cX45
yh6GuTeRUOJRFLu7FrwyNCNqTremSzTFeYyvGmsAnXUP5oh0lu3cnrxKOQaz7EdytELSU6jCAdtc
xWW1qpoTrx7LFcwSjhQbIOou/t2HX77mujHIFwaY8jPRTNp28E2KokzaN9nJBzoV50UGi9O4VQII
WzXOapv0YxkgJuEHdse3qPNGYUPdbjOX/Va2ZWir3+yu9AbWPA+9qYFxtUK+vP7Bw57xM0+Hy9U8
0RvxSEYGO+vbylqP0/LveInmKmVzuixlHMZpEbd9G5sJB9DaTzB03FsRFNNo/vJSv7U8XQh+xtvP
cMNDMihSjzYv0qQTZE9wN9mT+r/l1ZcV/QmxVYAwt9rpaNBgFcU09/yaTT0gGMNehlpVy1tn2Uki
LyA/U65mPmV+aFJ67s7MjICpzweL9l0shr4bO7DUQxFLkNsdfdd7dZ3mMdMfIxa3XwOUlgvIsGO7
QD4PulcqcDkLEtM18HghzkP2EKrqLGumuBLGu1ryq2hVvGkn6sUhBLoT5TE60YxklqWpf37V7Vm2
gz8iKJKKnuIw2XMcokQgROgvWIF2d5lCzBOtNv1lWbWUojY7X2mHsYhPSkCYA2zgg0nTu7JZYq3A
6NfikBNoOZ1/ECvAHBMk6T5AmI3uUZwbWwaNfnCrwPHk/KxTSRnJbpIbgwQV3E9Q1peH5Ql015sO
lRdE+WIpstTPr0pWQJh9eRgLuomwho9rKEjSwzkctVqMEI9S4xLO0xVcYR4118kMGEm3gOn9F8oG
NDTtkCAvCJomLZNRf2k5uT4VG9gKrIabwkTokJTSVSa2IVqaDnDmRcDmEtIgHH0YYYglRGWuCjTZ
R7vBC8hhUPE41dVPIEeV1KaYq5Ail128znMDv4Jwf05VGMSrJR3mzHiDwNkFIOIQfFHiLSYGLWtk
GzPq1mS7sne8AxJB2CIImQerSkWnx3L9H3qg1zWxRuf7xQ9CScphC5xnC3tDHEGFvFt4W2Fsi9CN
qEzWspw4nwYxVD3rjoYo0YXBPzNRBKO/z5AGN7k9Qw+MBBlXwLEHNwuGOTW9dZ4nsvMuNk5dhKqq
dwTigpiu79lAGbqVBJ0PwdjHiOp9apcCR82m1CklmnpUCHQMbMKAmsmht7QG25NSbA83Opv9srxk
yOcidAQmeRPX2fcEB8HYQG7RqQiYWTvngtgDGO+u38iwm5z+TZ3DmGbhwIBGZ58nq1kGGar5N+Y3
jB/eHQWKaSg1ie+UbMk1YLvoBpADqLg0EcL5IMijFL4d8Te2nyM+YrO7f0IDOmwxFQXGu+6q7f+B
nMMrHcXil3unbQWma7Wx+pKJqs9eGyDtp25+lHN1dLtejnxitVpjv4F4Ojn+RLNMPcOS8g/kXs8T
/664HEhXWmqnJU0AYtqJkKkoutOy31ZFc8QyOqzaDKLNTBEc7UoJ8EPK4DLYDcmdZRdWZMqWN85o
vQf+RVTL6e9QWLn79NzcHgatkBxpBx1Zh8qmx1FDj0MEikAuW9jexbrmJ54r1tsJg3Fg/SuatVcM
wQkVlXMls4x9yMWwYJIVT3Z27MSwrKI7aX39gN1Bbnm1yYWD9MJbBUQ/m4JlCrRHTgMGKfHGq/Ou
jh35AecOPgKlqnrxC5+mNZK7ZlYtZGq6BdhSdl/h7SPC2G9do8A84OYbmRengYk5ga3Bo7CKKR1A
fZ0lp4Bqbju4U3CBEU1foekP/bS4xE13rsiziPT6y9Tj0wlip8O3bmJiu1lq9s3qn/uuWFevfCmC
YCrvNbp0BCt7rlie3r2EVT7wZl0JkEYnea2Pj1/LfCY/MQYHyBePH8duygU25cyBvvQcL8e+trH7
mg6Dhd+jrOBTeYJ7OweksfUPB7UD/NLMwhXkt6r42MB1AK9aIenoh/S3higsI8iJ2X3swIBtskF3
nnZ/mhk2wMj45LR7NwSYlQSAWwKMpzSOoBqiVd/N9+eDHTN4cPuOAbZpVKlH400kxWKwfqCbWz3N
s0d+v72IsGRWp2kKF+td8ETBjXz42+EQsKY5bO/xLNYYkYI27gBMzIkw8aY0szd8iq7gfo8cuYNf
op/PoYhxXWUUPIpYQA3dd7gdiKM2bO6YpfdYW8XkEDFB0KAB7OCQy43k4j9IrQi/qfTHZmPwgnVR
7vSllUXdq2JkhHTXhvKRrmJ4x1PuQN19SWrvhW9uAyRmACriFi301HkSEwJyoR43BwI3oSELnv7J
O32T5HZQHWinDEsXhMEk+61JM/hdP+tgGHfxl474aHQzep6toaqzz7R8N+g0Q76VAMhlTd0Q3XPZ
MVsvUmKSlMkNSCKN/GKU43kcRPZbB0s34i6FYgM5/dERjDa1ETXTLPVWl/lY50uU85qvyhnD2VIA
1dxnmx88PFHwPvl9qligcThmCNFEbg3K+MDCI3d6puBEsKgwtkJRQkBs0H5TX3ZyK+yY1ovHGiCJ
sf/R2kzpNFZ73UayDoHlfSDac9NcSJXKUWxKyL4PH9GM14EyF3uv/5YRE02qYxFdDCR4sQAOH6o0
0fphwUa0evmWc2JUqbF4VCse3t4PpqI1n2PPe5RZcjdC8IM0ONH9u55aW7mbpPWf6fen3wXubNnl
aDAHOb2TH4LkJqsNn8SApjki2oo0/n8gJTqqifxLbX7CdukvysMCcEnN63Mvjsg7NaYha0CtLi2u
VDAteyog1w8SYF8OaN8O0CuP1LILTFy8/DUGDCZp0G+M2J+Faym0vg4Jc1k5UvmCO1afdly8Cv2+
T3zs/X8lQxVRlwqXPFd8ARxNDk08UpHQ83Dsct+JNTZExJurlBhkX3h/6zKT1BB4u8Slcb6zLtRE
Ec61/A80uZYYTN0jQtMOTGo5DXtfhXptOIX8xjJvGgVlsCsbgEzj7lXUQQUCOvFdl4uzPOBl9sYb
Z/+Nx1DgNy2OWeVRHkuzS8Dqtg9mIOtDyapcAgIBrjV4CdYiifgacB3tdOAPCl+cFKv5cBN+IvEo
1dnGv3XfP/go5oxglnLDd1yQZfyRLM6J8MS6dBuK7aVhmTjDVMIcEiy9Hatb3ESpFzyA9GU7KwkI
DkJhGMBL2Hv+5hqMBcp7A26crkghqyUsyLaVxe33nc7UiMiWDe70Vs/g6/EZUF7JzRqxFEqIKGxG
D188DH0JvhVHFTASfiucJdlm7CFAjKxTlomv74cXTq7dZNUJeG+6fIiftAaq5sAT8VIj/aIFSS3G
vr5gFESei5qYmVpmzGPu0RYYymAhZlM9Mv2w56MeFEAEwx45/BEH/T302qXu44Zj2hoSLPmNq1uV
TVeWdQRMoVAZs2D7QMryjm8B87IkNR+Y68v0IKv8FBnJD0khtMLR6gmBi6oPHBtC2p6LXFiG0n4c
aKiKGgH9qLuK9lyIlEXHLw8bFOnjENlhIuDHFpO9R9jjKaRNUtR4uizXzrgwkymvClz0K8gt1Vnm
cir16DprkBky8/B9+vreLakeVI+ap1E+EnVUe8iaHi5RvOljqlg6cgG2CmzGntpJqhnaWQHmo2DA
Lo27efOi5KeLHvlK2xrkJEl9GSRmbiFSzCLAJnNCp0V89MIGDNxHn+ZUrI65B6PbSfoD9cBUqyTd
4lRKzwml2z4GImTDXY2noPvAiK7vAclLoNMAc6PSycWNAVcLyRBik99/CwxNWfBTo3z70xyDshLk
0yzafOOB+gz6Cjo3iWSMdUWTRCFIJVSB2HkBWOsuel+PrPIFA3rerb5f6DDUkvnEKknFlgEkOhUi
mYMKbVFehnksTAKpxP266XY3TOWyRlueiP93nLCbLdRdIPZ4r+NGUDeuy2hLz3pQG+gMnHUu+EDB
68ZFym7vCoaf07T2Q/zx2elF+S04+kLkCGFNhUKYwibgRh+jxexhn9iaeafyZrUTwIazLDYvXZoc
kYrB72bdyi9QjnWgJUgsyLJOthwwLe2hpIlv/TLRM3zFbY8la0TdzZMiPXx4munnZ1ulQLVvRo8I
jcgzYbCsmV+3xepoAyZUSbldjC1LYrZGKa8ZP7HpgjbOWyuWw7p+xT8nVxa08UmkNTr7XcZ6HpCC
KUPVMzeyV1KMaZwH51ojrsp807MNpDyvxR2V4nQkJsp7FmveMOmEScrps8OX8Xh0GJ97jfnKPfCj
jacRQmWDeFQxHtGh6x5ntsfPfxfzreU7tVwfaPQ2wGNpliGv+mrhSqhHviB+k7x7SBu8v2VfCL2/
jYIoRWzS758j+fnfBZ9eFtxEmv6TSdSzV2HaRViZacdiBVlkRgWzJ1Tuv7yLLatojhPX5RWpeTQy
+zYkJq/XZmNfOoGkScNz7u/3FwUCGm1k67sPzLVD8uI1Wc/t7eHg/IaBsbJ84R/bFgT7dADm5Too
ZvWvjWuerH2evRNxXGU3Col+HYQxomAU/EPoK37MVCgF6b1mF1DxHzn8FRIZIHhc9Aq0ft9pyWSc
VaBjGKeyO2wR/pS+GixQbcnJRChu/TewTmLf6myPOfZZVC4/1GlSvyBuwhiyLZ49Q27SEqpszVLs
nNgHAPSclHiOS9tJ6NLgWqE4+9YxEF+/3x46IeERy8gI8IFFL1hdSzWSU28ZLwtHmNHfriLV2j7H
Lwf5akcsj1mYYKStWEJ2CxqOROsijbJ6f1m5MLEqk0BCIETk7aswB1P9uEGEt/LJKPy6M2mdlxig
K/Yehtofk3iBrbWKZOhDNZXYIUDOE619r3fjJrokLSJgQL941vWV2Fw3Kq28Dy9ORtTXWFoDCj+V
hnUugTvCwgcTmAe9gTGGP0SwcSfhRYEsi6Jhp4XFcx0mLVlverD5VXJ3LAiglDApsXUSR8eYBA4i
VDKW4qrXkbbp7b3Iyj3kF6y7VzkBY0R5l/6M9HiABHPpLQzIS1POBc28VgQvxhcM0sUa+U2urnKG
uyaO3xk9aN0YUvmp7AYOWI53Vj61LHLCzwe1kj/aqxCWvvBElKTz4KMbXuNwWce8W7tngqZ43nBI
zOnuObvNlkB9ynU8Q9lMS+I/6XThW5fEPVVJptfv8c6iArAyw1kMVXq21VIxgMyMWhtR+RDAR3ov
K/NIhJ8GW2IA8Mu3UyY/dVBqQQkzPxPViODANXzdBbl9xdNoZWDvXkDIExoK6oMmr/x8OOt+hLiN
buOemuyBAQmR7RGnFslxrqDFjBWS5bUz3PE/SmOwr9NC1VKZCzugbAkm3LxzunM7VNdkTpeYwpta
diqg2hCrpjxCZ2c0jfW+n2FdrVxoX6pY6JQqMnmZxPSuQgQS75HBPcb4+upWRnEeT0GDjXe4MfgR
te/LsncJZm/XS+EhceOaNq95NeovrSFz6HRknePvnTngapbzlMllfhS6JKiV18pv1yKz99G72402
hfijY1Qk2Cutb0158EYMfl6022PglLrh5UN5LoJl3DZc+4Z8Qc+IZZSgSYEZsqLnyfyC22KT9vzA
j/Y12t9K0+dC3L55VVN1AlRzwkECPj/nI6++2UCrGjt7xP62qTwY8MDx04nmJYxiX0R4nznyleoo
AYFe3VZNK+QNcF0KPDF85deL9hYeM14rn64cu0b99RjJjZF1haA4cA9FNqLcn+vwdEFfVhBv00bV
DUI+G7OAb9anLgZcmh0Oha4g7545l7VUlOPFhPXuyo9f8t0efRpy0PiQs8En30sHg3DXfavOcpz8
GJM58xXGejuwW9vJ5SzY9o/cnjC72aJH2pi7yqF+4zui0T6VvNl/U0AomaAP0Oarq76Ev9X9l3SY
xGGl5Q+3D2K5aT3Y8nySz3R3urd9gY1SXxKu9E42vhnYooFneUOdRQPyEdG52U/VetQ8FLNxFzKk
wa5W9ZXC44eCOjeiJyukWMle5nfHIfSyGDVspr0lNkfIV0ywN27kBjBVm6zju4zYteUn1/nC+cT7
1SxHJqgZQHHbw1mEcKshvdavuubu9fRTtYBhWNJwyKPlJfH5nJ0zFt4EzBXZNV86ZGMGwrPCmFBf
3Q6fzf4KOcd/224E58S/zEEHXHQCbu349HmqhsnyfsWBD8z/FWnkgOhPX0MFg3yPHoOtONQs34Ng
b9w14YT1cUOmoHvgnJV3TpHTrv4oXT1UmCKaXdDFDgqvugzfH9U4afuXuPR9+d8px0TAmT0xer6D
xvGdjxSbVkeCfNiWQZDHlLz62B5vRupHyd6BcFOqe1JtW60ULPUQi0AHXr2ycK8yGS7xL7s7I4Yp
kWOVv8l/wxFTmByr27wXGnwNvMtvUFHS/Le47sFTYgtOIv4azhmm4vyw+iJzfIBLDvD7ohJJjckQ
28cRvaoz1yeedo26yAnt8PmhXybqREYueGA1j6KTozRAx7aBSodCsR3+hCcxCa431mTSmujj2+mS
9BTmUKimcr+wER2bLY7laVHWRBLFcBDedIUELlF87nf3S1qiXo8b+E/NzPv8+iD4RwvDQInH+W22
mlcUuOeC/bz2wrCqpwV5GP231BPuUdeFxVyH4p9gGT+3NfAil25JsOQCon7JsH6Gm/vDwzZp0tkV
aZyr0zvmKdB6BkcW09VkA/XnnoCQB3INqfXYqtg1stgnUnh5uzvMiylIaZW+jI07UppH7VGapBvh
2R2wtBmWlI130AfT7S1p/D1FwNDBC/QNWt3M9NU/Li1KZ6igwtDETpGGTLMdx6TQtO9ezatcauD2
p1denLOASQT4Z7U6NhyFixaC43eCpnAsNjui12O/w8awwJV71ZiuLQCfdgIjrlKY0kLot7R1vFT2
ivPnINcWgA5Sqaoll7BZnW41dk4JEhfW0DnS+q+cfC/Cg4XjWYiqPj2lWCN+q1PSUgzWoz4dTIm+
d7aIK3c8t5TYsjpoYnZ7tbcWwZmDZaEryYBkaNTBjoKt/2qFNInIuDUReEVC//W2JT8bWqinEj0a
QxlsssrvQEOVlgtdWN96nBWUhdcidwPcbS7q39NCgQNt/ug8ZiHCQMBCOXBAjA0DOqrJ0I6KbPIT
U1IaTZhrm84EJo7UIKEJqCEAN3QBq3vI0Cgpd8KxpfU30mGEZTqT8kauSC24RAvmB8gZn7jITPOg
gyyXgxl3VY5weJHMX7lt55pD8bNJmu4xc00n1mwUVFJTRyX2Tl1TnEOQJ4jREW3TvUHalqmwFEOO
sP+oFMlTT8XehIArWOy4oZ220CdC73yBXqOM73mTaf9NniRUymwxlC0EQtxCcK6GF7Xtxe9bo5Kz
fVPE4EPd2uNrHFg5aL6n5N8tMdXi8eWFwQZJTZ1zONz9P9nWwHbApBZSByuIlaj5/Jwt3Q+2B630
WW3i4k1EDBu4LYR1whjnYIZzxwWugOenXH57+TK7nm6So4pwq9eV9A6j+jTxmiwLPU3pCTvabJvE
1w0tQlvaG3jp0YpHJRKhwU455uk/sbD4ZrlCQtLW7EvbbM9EUL75Dq1dvi19h1Sbz8FHiktAiq6j
EC3sNIiXn20pwyZUmisaZBL0LxywNz9tiaSshk8nXzx3RRHX+32wpYK782BVWGuioU0L6p1NCyzQ
W/p511lNV5Ru9hqVWqaasDADxlNoAHaxOhTOMqnoJbdisRbEPPMKy3TkD4wmF2/mtdbWDEWtUOwV
p+70tqnA0rWCNY83jgSlWoadRftDb6QjQYTOne8Mg07Cd3qcr68ABrbrzIU3+zSkSkJbX62NQCUQ
7lk1VPR1iBr5KEscX80gnXaTm/gaQMOfsMkGLAIQCDula2oO8wU1sC9dRH4p3W8fqpsayPzkDBMS
HsC3UwXT6HWgSHHZ3VQj9ff748fvwCxSnmhZx/qNF+c1IOh2bsPqBUivQkYRfgTBChuKefU0HRI9
KGzEMVSHI7jC0KQpPAYI2DgmwVMhZzSb9BTn85f2eXTCFdZaG8gvFhV32o5D2aMwXrLtTLpy/6EA
2aT7uXeceIhyyHl2UtTwWKYE7nm7lZoWXPA1hd45lrMETbLOzrZbzqy+9cG47yjEm8M2rpz7Jq6S
RQItvYc/gEOKuvUNsuYociKPibCRokh8Dp8TY7mt/1ykYxpkuEzESogxPVRWzi5/wcBYXnecj68a
PbJZfMWwbII/QsHB1z61DoY+MCM0m96jcxaHqFAPjtyiF9mZRrRAX8Lca85rmv4aLcEjy639TrZu
qubYsEnivW8H1YqmOsF2d3upOyOh19QZD0MwM43sOjk0XoxhYSYl6wV/aPcmYxdHAKBJw5cDRUW/
zyzBF+J9LBuu7+hZ6u9Y3B1SdZTEQPKoIDBbtwEWpHNEv7lf/3/iTZ/0TfvJNtb4n55pagA5LYF0
RtLRvADDQwpQTu3H1e94xOdWlixZLlQGX7bScVsmcjI7YmA+j0T2SDOYU92+NwyZE6CMATo+PlX9
YLX+reCBjw/llWu4CL0kykCcR7L8VYkrOJUPzznF2UaYxvwu1IrLOKNUakybR3rrPBfomF4b/Tvc
r1SywWKdUXUibYdmnfvSubr2o1/MdD+MAFAeRCWJAHAbHY/p1baHzCHaeIXZoljmyFd+7C5X0I3A
NJvZLLBbBoRfOWVCVcKVMKQc367f0+l26x+HS1D0UWPGqjHj+WpRv8baKiEb/SxFCgEgUokbVqrL
Vu4FfE9NNVtfyVX1xk04ZzRUgMMk6GDBGbIZYeFyeqfKlB02a1GS1X9DR47Rq21NZtm6GHYYQJx3
Ph/YxK4oehLn1BcPJT80OSpXqq7rFWeeFn9F+VfLi6pA6G+YYLZl/XMl3W5dZYkwX9/VzUzT4lES
T6SR/cPZyQ+I6p7nqlFtwsrXuD8ogVjaMCz/+ufeBm+8ejMqPLMjMbkYDr9rBtZlUPJnmJ3oA8cp
fDTlrtE5QHvgnR3CWPZ8DvM5ef6IXjm8AQWoTV/0NoWSKJT7aVIAnfERZ3t/Lb/dskozrk4WLHsK
XB6WtOz2yt+XpSnnLHmGi/LcpNVHhvC5xi9V4xRPmLsV+uzykrBG2d6mVgolwQWUnBmUt+spesr+
nj6HSRnfjEAia01OuBMtdgxhDRj42G2lyjLsdooCUR6/ugJOm0XCyLYOMNq8WgR2IT/Bb37cRbU4
yWaZz6RfbaZrZ8DmHYeGUnqRvZatzrgeayEL+l7eBBucZNe0pwTdK1REtzkxgpYMAJdfeKnDSP5X
BaNJ9rK7309XzAS+YQ3y1TaOltUa8LPx9JkRsgq4WmNkYtRtBLp0qPVkDW6Cc+Bzs53AEbdoCJhT
E1mhQUCcT/HZ6MD7bULj3KyMfxzCyDtY4QST/VuziCL4spdLU5paZzZvoavdhogAeIFMA3eLu6SN
Z+T1u2Z+0vEQFD0PBcfU+K/zjbtHJ8JM7Ef3vPxfMCokUCWwd4EEHVMh16Pk1UUj8YA+IwVSYdCs
JSXLKzzC578VACWQG90PPv4JzCx/fmf4o8sLAOlq1+q0IcjMqNE0GpmCKmnMEq8DHGVLUsLXEsvu
eEaZ5wxhyzsEPxqN/LqJveyKGDl/OP30MpA5UJD5/4EJfNh6Y1fOspq/hIE5C2lLi2863/zt0Ilt
iFfNOwQORCchdZSNt7uWkgsxav1nRBxRH/2gPswAweHc9/1uTf8mOmA62OBPuVmoWNz2jx3MODwN
ve0mJx7fMbK9KuBpKFeTMvLDLk2vhtyCg6xt1xlEwhu1pfz1Z3dZJQE7PVCB2cxrwcGb9pX+O588
YYH6QD1azW3UVyDh/hW1c/qdWxAgodJFlBXHUzGtgAYqFplC492Oiz2vBksIF+R7qj6EgVR6+9Jd
QPJfNS6sAm9s5t5TpAuJtlHerTJQBk7F1cJRu4jSUYp6K0D9u6nGcbii0pN7We8WEyHTHSjckGRb
RdOFMshV1Piag3phiYX14XGbG6H9XuH5HowxqpZCxPLvokTJSsy/ca1joHVLtGWVn4YC9MQi7NQM
+ZadHAHiCbC6rLeYdY19O+62/H8NU+HFHMDPpayiV5M2gTIZvMOglFHiLfppyfhAsQLGSk4hzNJT
VW3z9i5iTJkEzMJJbHIYwoEiRqWR2+/pA2j+8yvdifRzpIi0Sj4wcN4deSAk1DsCeXoEaxmwHL/L
wpxTblyBLENyIBHelaP03fmYu13WNSgZwjowNLFcZmndYVQoTsBDlbnxjshvcpjEHCXs9XiaUHtX
u3ZZkCLcEqusu42rq5UxSQPgaL7TDgkT7aAHiStycT45dMG/Gwph94mGp0UFFV3Gf96167eGO0Rb
8yQZks11hduUt8gMeE2SqsG/FsArO4F4GWiRPcvFT2hYvoRvnKeSASc4lXRyfikkRKaiQmbKmABp
9G2zEwgHM3UEnWq9WVQ/GEDyp2C/Ht9e/1IWZJJXYY7wLfXgygHm5Mdy4CbxTrO1mXv4dCOIsqX/
I73BWN67VEtEx9fUEohRtQE2TOKmVO46lZ/tjgyniqeBJTGvQByOgcIYCvZxpRdeGSRxHLBFTNbW
GTJszQmgINhMA8YLHGvRA9WrgzS4SthtckiheLRCeoh/3wPyIFS9oSJI9nQrl+kx6ToImZ2NaiB6
606d1uH6j7B/fxElMCrn+5ISbBuCg8lU+cij9pS/R6BIXCE11s1MBeD2K/FbgQS5urw1/5zl+Xho
bjRE0mWKwnwLpl35i7OVBLSPrc3WI8I9vjfictTJLWYca1X/lvGa2fLzgiQ9YOCRGB0SDpHbeNiz
TYGR9qhZELFMJZQbpTwKO4xTQqxlm+0vLDs/J7dk9NA3BOzHFJ+omPDTMaiBLP34QeJa/UjgyNmk
jgFsP/27JZNY523DGA850o7fCLQmLOTBBSsGDEQeYoet/R1DpLr9SnadWq0LEDGfy0N9p7UqovhJ
0UC0v0cE73hWZ3qjRhsKLi0zGN9KPMR/cfCbyeqY2IuWrFPpRocx9xOkvvbN59Bctkl6G8ntFMAe
xveaDppRYHs1WLjdXe1chxEdjZGAzUVwtW3jzcylZy5ScahcXndySFTaCIXP7gePLWLuGGeYTRkq
gBQSUBKLehNs4dpy03kM22r2o1RJMb8Vzzw/fhklLRyz9ULseUo3gowctsOv1motZ723g8yQpKj7
2o2W/IN+xeYahcfGUN3LG5NANHmr5tA4VxJBzBE0jT1NIEEeH602vsemaYIIJgYzfUmiywnJ4www
41X0QXpBPKq5fpbB50pewxbqwpUZAw/xX2qzMUW/h+XcWnr/xjtd2k2sWwd6Uo6yOyv/GtnQMPUR
SgI2Cyo4nM1cqWpRYMy5RTgijfu+kvA3uHH+H2NqAFiyIiB1cfoRhzz/o3ZSY/ImuTVUccqCFsMK
/FX4y+GoNNS9o/2MPLYpogsmzV62vFUcrAuJdE4fQ3mU7oDukdJt2RxCUc+6IGpTwCaV/NstTwxa
7BlpQoLV3kap/5aZZw+M3lV34mJciRPZvheQ4PiMGBHiA58zXwiemyB4cy9Z+imK1LDywdt5NEo+
aIZaOrl7AJn8IciSh5TZsKd4shDr6o1Yn12JOyJTNuaPf7EPn5TRM1MRlWwpe7TkWTsPKWIVkQjG
BfZQIgm6hZiJV0VZt6+DOFL6nTMX6kWukIBnhZUVu3AAtJqR43TeigEIG5m0KBvB6+8HzXCJp2LB
32Q5F4h0VtxU0u+U3kftLXkOHq/fBMEDS64A0XSkkn1Ga3l0R0EDB6GDxFlhNOgaCqrCOnmiD2cP
u///KTul0nmoIuZsc4eabR57jdnJBe0z02GppCIXfOTYgJZu7qbBrr2+jwO+rC1UjauUuvvQ0OS/
E12lMUfbDt8KSgFLwkf8yhguW48fBK3Sg66OlEQRRpOIGqzhKcN+Z+o4sYfGnZ2NMThjgcaKmpTd
AoYPORItFpNJTHy0MkAksP5S72LbEX6/ZS1Pr/xHqsxvvI4n9b/XlEzK2ncZE8jnfLC1wm9ziczK
o4kAlPIk5DNR6AzMwuGiQZQ6ujQhMxyfcbcLa6UpWtk40y8B794AjNBvwnER+sJOusoJorYsVJYQ
Jf00g8j8vFS0JEX/nhsXs0rr2fJsjAcS4RNV002syuryzPXCfuvEtDAHA2B1TEdt7v4HNWLJOJr4
koCHc03LXs0xLZTUzYWYTSG+KxWKTWPbsqtIzKCZM9WWItI7zIT4r69iDhgckXEO9C9ZpNyv7EaG
iqDdCG5CWMoFHuAabMnL5F5OHCe7ym4loBRXR8WVJOKHgM+JTXjZ5tIaAGUTD26lv4DXfxbwkgFr
LFzAoS8rEiFsPdVqdmUyzFbDe27nKNj2eyhHgglfAVbG3fGKTd7wtOHa+1C8ZsDrdHLppCRgaxAu
8lgnKB0WZSRNdObQdBahak7G+UEHyRnK9QBY3Q+AtYrP3BlrcWNBC6/rUAw+2D9gI4vTep/EiwgA
xXPFmFL/3JMNXzczEPHS7bofCZsD6FtMqrvG+gJ4JsLqSw11VlV0oiS2f3+KqZfQv/DXG+Gtxeqe
pQ9iK+Nr1gnI22JV/kPLUFrwIhjvTzwn4CBWi1YESroe4CxJYViXp7bKc9nJQ3uf9tdNN+5vSFyU
nV2a22v1Tg6wRDFJvFYapbDXySK8ZLETxPOhEKDvSIlTJDisUZSq4afgmr9lKrPhJ0nZRFY6Ij2w
I3dezHcNcAtxHd97ORoI8Ds6IOWcaiWrPCQgHMwkqC/YQ4Sq1jDBizsSLc7Is3f0vH4BwIMorJVp
a+NVckxQps6K2YnzkMuvRCkNiUNeRkkP42iE3NnXkNI6OKmcJIsW9sclaYFKwIkVOGnuDzQtKeHz
4xmhWFBn1C6jLFeAenr7PsI87tE21MvbBQJQerkmFyge7gr9ol9UJbG1nz6NOyFiTWuQk2yJk5YU
5q/SjODwapTEd3QNKoor362+XEddb4xmEJea8kUQu3Os2ny3WQRXJBJB0O7Z9qh/+AHw5UQVtISh
gYnej1NG/7JGf4a/P/vQSM+PCQhjlJop/lh40Yb3mUi1zf+A2mofrvoAJmIQYlMJeVnFEUS5JlPg
uAVVHr3vylvoL0eDmxtTNAjUpaRQkAlV3tQ6XUNs+smWWQe5ztijeeRGFiZWe+hu+j7KpsCuRP6e
+0ChvTeLbpS/odBUfFSWvez2f52Wz4GspWNrpUlT2o9wKorWmeRZdrjcryzeRBNyZCJEVhl2iUQh
ylQk05KBozpsKrt9ZEolPEQ2t/2PPavT73id1v2msWpe8X/fvmnpqmnLlxCiVa9XqBZnYsuqAWD9
VGMc4md83r0ynr8viYxusA4Rsy8HYPaayOi38LYyPElJ2B/fxUsBwt7HmFLUP+Kla6a0bkq3v/r2
pkIeiL8hCF8JKtRupW9/Pokgln+6TWlfa3AsAvu+JKnGUBQ6593izYxPrwxEf6dVqMLcaNYAe6uE
d7lu4LY62Zo4jSfutCmQ7m/hXBy+7UEAiExYWDJ8zDQFWAjWRzcUvJAxK4NP5lXe9NwUZb64ypTc
ksyjQDmQrsO4y1Z8yADD/x0lz5sgS6Hb+h7/yHF9u+0fADz/9yYwGk+7k3g3qCSR5PGi16aYxrhF
i/zAjf94S3r4QPSMLjRYQQlzfmFI87T9mhB7yvySatCTbe2RlEp5vzR0JWVYmg8oAcXUtyQk7yZ4
vEnCSEHQK7CL6QdXbM8vxIM71kFgIQYzGi7PMdGILfQ6GBzu497usR21Ctg8eTsbOMV8thyoklQU
wxwbiQVCNOEHmO/4MmkVw4AjRkUTiIxDSNOLtONE+PgDZXajFVpHtUN6/6hPztxQkSG+0fE5eQho
TK9A+uz0Yu4YLxuUoKLDnvt9ma6i+fSEMIBHP3gWn2TVUGJ8EAWbfQeXIgVtC20Zupv+Ags6B62f
DJ53qtFtQE0BogvqaXVZ+g6fu3PX7rHqCEw4d/809Tg4ICa6NYZ6/FcnbK2NPV3WsjwJ20lE9+qi
Ao4NB62H0HQooffQ4BmDYilESS7Z33wwiwvtItsUDUoY+ZvJxLSS6rbk6Xu6hWwaxaFJGzcUyM0G
Kh/wdMUaQahhoO2PRKIjkjZ6WvVAeg5jritcRoLmANf6oCZG4yxdAkfJfOkzZgvt2D4CtYh5XTmQ
yqGNgMr+L14ux5JJed7iW1AZVwZLxJaznHiXqMkZ8XLDQWhHkq+RS3T36aBS38rCeahwYB4e8ikd
4lqqM0LByGPLd2VOtY6wd4T/uuLaH+Qjxg9c9vjKKUoDzYQmFbYwDDmUKP3CiEUh6I9hAUOMDUxq
4O7bYz0erIbXJCpB8Kk2zVQV0L2OZE2BBxESc/i4ljqitOdVQsNpZLqnG0pDCEtMfB5RhRM6Q0Y+
JxSVUiy9WMOkHt88gvo5vhLrsr8EMIQ4xsl39iDS5zFK/insK2rZjBDqdBpiQTkVRQVVT302zsCb
2oTcEYg3bLIUaFO5rs471z4xX28xCBTTEDVUltHdfTQge8MxFZzFbwowPF65oMoOeccSCnimza2v
Sqnzcb/9SCxLBy926J/Bo1ftcHCL8ah92lCezuwsoWCGkdAQve2XwO+3MkplyMa3q88IfM1atbQW
RDbGx/eVTSyZ4e7VWYUzsvmWtjtUDjt1XRMeImHSkC/8WIKll/kRERUE+tIGZodQmpYK/+PQuKEG
9/UN0t5nKv4/iGcNeoidjsAj7KE61QL5mKix4e5V+viOR8mq+CtiRfLifUAfom3uxUoXMGt2Geiu
+rot8HE23k4izMFs2L3NHQuHgzOob9XKb0y3q6dzRDDujsdurFLnd7OoiVEo4gZgs/mCntSJqIMn
81bmEzuSQbCVcWjQv078uVWTW/ZrzNJoaZCr261NdKvCudSFpKQDKCMdaR0unt8JeFUB7NMkYeh5
RaT1b/WSwoNzdZnZkJWWYuNZPaYsnvYmb/MgzbcNsLiFbW9TpK3yS0TN/jTFGRxAiMBVcf7dlPZo
ttwJVgimzKzxx9BJ8iwEeAoOTBGhNlKNI2ggpu+Fxd/10yAacP1EAXsb0LbxNTXWPI2iTJkJl0Sg
x7qN63VqD8/ph2I4UjJIL5SrJsY1aAIXg6uPWZaSSpLl25Sov3IcU1XMWKeP6DDo6eYXZtM3uH1B
aq28t46pnvfD9CpFT/6o7ufhUiSLhx0iZ8L+j8+/lRD5O6bK2hvBJ02KrKVT6QM9dK3g8WoivVtQ
S6uz3TcQsiw2kuxIiHg98iQpKfWfvJn1d0Zj+oWHAciGuNeaQjqIRIj1dPaHxSev9xeF2OxlG4Vz
vZySdQQhIO5Drnj3HCAQpgRrN/oMqSVQoCFOKc5GMRCUtJu06ue2BfcEBo+xgVtW8uU+a9BidOss
QKIfXALYS6md18/C8cE0v3OrRDErXR2R5gVkL2ni/IIzJjXD30x7My/FfG7aaG0XSWL9qqVWFHc7
9bEYtg/oUsg8I1jPZV/7PVvG/L4SDrIvlzJFAxt71pfpYhi+Cho54lTJhfXlOUVDlyZBArili8BA
I1p6nnAkL9NXNYErIOlz9R234Ww0AXWBXXt2lj3zVV2gAwRpzn02CMbgr88TmjD6UNkQ8ij0zvQq
g42TD5o/yuqbVRJzP6FvoxM3DN/DJKrCgfZSkp9Fg5wwABUrpEJrQN1ly3wf0AN3B9C++nePJCc8
jM2dbKTYaAUeZNUJdw3N4gE3IQpiWpHKUJqb3FCjjf0FuoYCmFnwRfM3u8sBHrHvpguo1hbZRiBy
RncB/ezllXrnDoiIbLrZto2swZZHxNthaAE2P+iugn5uLEi6LbuRF+ow40A2VICO4mw6x4hC6Vfe
tJGMsx8qj5+uP78M1y5tA3juMtWfLVfCVDWB/mAtW+3tvdv1lXSOXFpm3we+i8N2Jv85rloMjlIV
O9UAfvnN4wgfsUAkZO/hOl8FdSYGFtU/kMuZuX+ZeiZghA2fP/p2HkXm1ZIwBrCU6t5i3o8ZRJJV
03r74ZLtm8P07Jym3YOY5OWeaPTkZcEIsni+rIf55jk4w3aiuCzguk3MGWwgxqyCH6LA0my+KNm9
Yzqp6ObV2VT28AqIc0npMqPt+Z0LR/aIUrtM0SfJSvqYfHBa3kBIO+XLZO+qWNcorpEjJHCu2Hrb
mwG0mpDEr90xW4kyKFTXxIvkAE0jF4XJp6EW+yZ4UnQKKxtikSCSZlz/uOyhHRoI3N1EtoF9jVFN
yUrpLpqnoZTnn2YBooC19Dl/ZfaT9Db9fpCMRRyLUaFqMUKgpbu0aKwEFcWsyizI/dEFAcvKpVfq
6jlfWAOa0+NLXH7BlATcJE1rastFtn16C8GVwbLhL6zBFE6Zl6pL+lFj+Xgi6LYKFi84+HzxORw+
/kF6hhCZpjwMlnTZgSEY0wMU13nt8DkK7V/ft6WH9fFWc4Jzup+0FvO2LYRjvmLUYX3C6/w83x9L
88BZKvAH98QU6MWEshsaTvhZtN31ajLKI/jhy5jaQvfnjaDVEBO+rCJ4uztQjHE9zYxSplButmAN
iN7Q7PSPQ0yeOHHoCo356Y6KxM04R9bKUQe2PlhLCz2eTATZ+ANf+ganPDfx88Y+1zQeZOpIC2XA
8gFIf8CPNgRz7Pyx9c7rSPjloIYDW5/1cS/BZC4sCmi7/4c9pthKrXV7Ii2dzxThww4JOV2Bz89T
NOR/ckbDMNAq3y94cqhDNDxPp9Q0ZHqFPXLfFGV11/waKywBrrxMly7ySQACCBBHQLjlHycycyOg
TZOgmsq/7MxwtjIt3KMiF1kdEiaHbXzKxZqnANVETLrsCy9EYpQGPOw7R33g1hbctDt8vTiTlwSq
PI90A142PBqPBfVnsR50sN1XN3qQs+XaYYc1L3++KUmBnD0VjUBcHmnneZmUWgwvhisQa8K+et3I
FqHrLrno55Yf4QclUDvFp8Nkx+CDsgc00Gt+k9PKOa9n/mufQryAzIJqVkEi4jJPBRT0pWvjPhjt
f54EzQNQxrGjtbITxy2pxYvf7wJ71sA5XBjpgHgOIct3R1FIhSk/3aJwfeyZa7OBKJttWv+kyxtF
Drb+cttrTfKLMVq0eeL0KD7CLLjphMFboLCu5o1Z4+BZEwmUqek17Bc6FEcUmDYrkfnaGC5QP4s1
zhIEyQi5ZYSkK/6SZl0XeviSRa8zu0oMSv11L53WA/mH0aIoF2wSAe/Fq/tTTIekL01isHcYapfc
oZYzMOAYA6RBP6aor6NYRwAPHTsbWrgOqzOx2SFR6bDYaXQM591KRtzDfI15RsLKQ0zrY5fsKA02
q6mM6ZIUKKKMjq3yL8IgfrYYxu6H6JogczcWBoFFree+4xne1USXH5M7FIUP0V/znWxTCXbJku69
3TcAp1rwEEqiaJIhf2Qc4AwiPsAH335JwAMFH1tlYResXkbw1k1McbRfyLMEkObTcQeK/is/8Ido
QF/RUalqlem5xtH1H9vS2dHOnpGkOJP19sCIYBrMTy2q/+E8W4qJTPmdd7omVI8rB4y74EPZtbTy
Z7xQlNr2i36SGToa4MX2R8Gn6T/178Aq2ljEpaldfaRd68j0wlQnpUgnp/Rgt2/I0tyMvEyxQXq2
NtuO3/iYBaxfnH5FkqHCh/Dh73scxIElL7cd4lfkE4FiyYWXFG3vHr2moNTBzOTi8GZBC2gryM2s
Enb7DRhYlhi3EJXBpZttbORZW8brF6g0fDjkbIy1eo05LGZm/jmr26NQyUkxasiL/WnSKzTdII1x
7ucX26IumfqBB2uHO6HPulM26W11+oMsI4SrU91TfvvXMZbhRpt0qoeli1FUsj0c2V9o0ewjG6y0
fW5Ur73929/g+G3NsHsKrRmuJO6HnRu3PIwC1zQYqxRiLXSp9zeGR18WjOP9efob0t/87uMfjrue
9wHbrJnuVPhg4RQ9C1HnGmYXJTYIL530tngyq7AeKChOGx+WQs30P2JhwyMg5qFal4SWb7/7vsJA
rxdW2XMg1OGgDDIwfhw9KNtUmX0rVuMd1COiqgrYSoQYe9leMQS5HH8Ox82BSar6LuNFnJL/aVIY
fDPCa5dPT4/jRv1kiGZycftdHL9NatPhv5TNF/n5Fhk62kP3I/NGyBv3e3aIfYVNUaODsuUPjk1I
l4t2ZM6KtniSFWPNUUeM3aZhBCliRoAZ9cfSugiACC2B1WtoMGrJOyDIsb3cHxQMJANM2W16rs7C
Z4uWf8FgzlEINODifgyRkR4bPpS4WaYTSo2d8g/O6LJPYHGekeTnjnUt24D9X2tpomPl8klMao6k
39uZjR4PCLMUOZPb7lFKtmZUqw3mjoTXDdVFOhj0f55PSkCqh/yl346dfOldGuTv950spgUeUnsE
X6eSt1kvxIfqbwKQdxkuX0Hd18CRCseJLxI7rznhBs6N0ZvnGXBBdakVq3n9Q5fzQzJelKDqKYMs
lhy7K3Ui4XthOWN21Nif572dHJkPC/dzGZi75worO5tPo1qnY1mQqea8l15eLBNk+H99Yr+VGbel
vvOzmFxL7NeXtjd9NDj5X6kVmPz690PKIW7Ir1p6XuFlqxezNIj/i+JA3hG5cK6dohsRrvP32gw9
RA69uowehHJktZz7eqlk0+J3IDvDkRciptKCrqNRB9XNPbebi+ZAX8rHR6Fd9xf2M3tu3bttA9sm
0T5G6Sy7E6IkzPk9aMO6YkcooQXdp39a6Qz6FiSH8PgV+mzxj26c41tY7rr8C8307GdlPfA0+GxS
k+BKC6GrlrXDIvClaFxbtXy2FbdrMSjYiBWci0XreY19jOQ2r5rRc/D+4cVgsLQvFIf7OCGUK+yC
VsdzJebXemlQogK+TLusFXp2YS5mroJhya1uHOXlcyh05E2/8yXweeNIayRKffamPbDAQCtRmrtN
PdnMp9CnA088a3nh2KKUkvvXrlPMtqNvN8czuKZNcsgrBZPwVvW5Q9+hKj3Uw5T1uR408c4B6Y2F
AYtV2HuSRoVomt2QkBhhhLxX2NZoMTLQiD8Z6Guft+TNLDbDaajZSQtRcC2qNPMtuPQM1qCy3AOm
dkNSFAiFne5wEBXcw85CcTCE+VaTTERWY5BIHfRagbA28fGlLHl7EwlDg0LzEh1cr0CN595bCh6N
hRF5M5I3Z12u4thUwAGHNFhuzt6aoq109c+8NDOSNQ7Y2j26IInjcYkAHhM7ZKVb7gbvpXNiF61a
e7FUV6qSBi3ekA9IUD+ixxGwZAMD39n2zOWJLSj+QYECBFdOXu8vViANjEFQST3o+ex0sKUMWmIW
9KKlB2Pm8Beu2+sK3s/y45zGorYlhmSDpD3aeLTqAcmBAZBSjhDgOB39Hmb8lPXrHNvc76m5QHvP
JAxhRt9vYxHjTmGAI1y7pComfryqPRENEnQ/Sk1xUfKQB9RKHlYHlW6VCfosAHr5UkW7s4seYUUi
W2DHpXKU7+w5d7vgw8qE659LscTp6+vzR6mR8qf9Cw5xq8EQzNqCxDV6qQxuhI8l4peQ78VbVTOq
X26p2yt3x9NSlpklG9HsqbewD8t1acS4hByUvpA6oaCzCf9g4OZiabaVSbwFnyaPvpXvU+WgnHae
nsc8OIs71LrRzzb7omZflf6tg8NRPbG8/Pf7KpMdQdJ0fbXzk0z17lm1C0hwDSvH10piHS/yx5SG
iwLrTTQ1MlJIgGmIYvK23iNMlWMdyFMuixrTQy9bWqmTUK0pYi40WJqz0yS66FNIGiHbxBEJJp4N
QRifDH+U70BqO9BlOosOi6C6L/k1GrF+oIAG4Qf8WXBhWSgh4v5usQXBsMxS+ZDqgR7fLl36ScFt
BBclGRN6dhYhZ1SeN+pN3iDpWYFuevCf3fPrm3iwEqxtpx/3sOCxtgJqLFIOnqo5vhOO4rJn5wgj
hFlEHzqu+pswiHZUNQNJ7zGbuL0ycyZ93qr8dhxdFGeIQm/nKzAagNifwXoReW8dcjO5gssFlkqZ
t6TaRbcoC1IaDMKcVF6dkXQY9keayuzAEfUR6Dw3ZuH0uvzZS2ncrfN76+gi/CIDMOzcu+QnhZ0o
LQYdGGMnL07dwsBi1WM87nJJgl9TVP0fQclwPawig9x5B7GaVxYhFCi7jzUmhv4LDjJxKsgiFQxK
a0Rn8LuiKC5hVZGaIJOt+1VubYn01UZCfwOZS2pe1uCh1o8PthuFp4DVS3M6YYnIhu5tKI89arqT
98EjPLMF+rIyRH9GP3+o/8D8hd7j3+pJI2667zQxzAKYmK3RUDysjXIo1oNvYG62Xnfy6vlQHCHn
Tko1Ljk5DSWV3G+1s+YQY1PqWK38wEvyW3/9meD5xTMUgB/z4EQEHZWakYRj1Jx6Ai1X8nOO3+Ht
i1gIYZQ7eHFfhks2OH3KG5E9bC02+e2LXz9c2EvqhmDQqcBHyw72KLQLKGfhvNSl84hoPFBECoF4
2/1lcGJD1xCFsr1CB9rgeBGfFcc4XAALv64R3ngjUOiA1xDQYtEua2tMeaTnj7pkyg9JV2cBrRXY
DVISmuj6erP+kxn0FkbtmZr7K0L/2sqci0P0inOoBOSdwobmDtzMk49ZvQGPf5RQ65sKEOAfW+2x
mwBSZ/ap11Hh3U5x6T3dVf+AaTtbC3YhcgVOurL2eF8meQ1mo6jsjuSe3jFiOstQRloIZEI7zAP1
NZnXi6aY1CD/X62yNJQBsAvE1oqZIngTsgBhIAhPJtYP7g8YjswHY5ByE3tu+OeqQeTt4So+zIjv
3JxMwDugTfKHyTyIdHzPkPdWvcfswlXZlMcSBsn+SwaY767xL1K5HHksl1vGyUaHysAu+1ryRcOQ
ga/o1i5JpUHzkvYJYy2FxOGMdsowTcNAc5FGaSmOOwipbinfhTCoVQHrs2Hy4ixKqKxZsLTTKEME
8bR3K1ojnvOtcqJd/HzLSPc8uqfaooWlGnsgr47KfD8dTv7LTt/n361TNSqyFwD3xHVLfDpX+c3R
2b0a4PLmg1JTPbJtbwxuXc3kkW9a1P0AiYEjx3MSDotu+E7W9MSHiSh7tj8rX2CSwL5YcgaNDpG5
sNhAaZdR9Oave7clpQdA3VWt2O9yByBvjTwwzTqnfKDshur8mrfmjFmy1nKQdnrCBBY7+0vbDGGQ
NROHj7dh2uJ72Y5Li+53duihugc+ALTJ/wcn/Iz2lOoiZ1RgGOSCzZbbAy5L6RrCdaBT9jA0dBX5
9Sw4+3J2vTCs71N7NI3E/NDJwXxYVOcA/dIPZsh5TH5AVp/291N2g2fRUYZ6XUyMjgFzK9G+m9KZ
+YRnU8FqQRMXpuXXfsRzi1bE2ETd06qzLvcBjtvtrnrYY7hZl4qDjAeGeu14LKpflDYHUIxLqesV
4q6VCtZzctNcBNJVfYMVaQjomG7Pn7fOaCUD/c2z10UJeQNXFtyk6NVst8bHKEam8PZ3Gapx/Phj
WyU/pxY35JPLNypnhjtJBtKdvAWu1r1o40GWbfz5IKSrZ4Qj9UHp5FO17bUnjnJm8pod35CS3uYW
9JbYkYRLsUmT/zrl7cn9g0wyvrowOZjcK3GFuHU108XDskl0y9bCylca7dtB0NuboVx9ThGG0RXJ
SVVncUqoL4ukKH660eJyAZ6tSzaUXSm3bcQyo2mBvHjhgTsjD+BzKOY3HQzKhyHxP+OMzYJd4ulx
rbfvRsq6wCmi+Lq4UfZNpBsRKdKGfgyAd4WJwOS+le9i4eyX/YDNdT8i71Fe0pmRDmZQP9g2M53R
qSw7KENprIEYudG2p1a0vuacbXLWf7/6DZCkqT4+Rw1oacw9TAsyZ5xAH4LSDgkJAm2pW9nj1w2e
dEphB2h04lbBFVLNLXUxBNo+9cGXvEuaOHwCvozNSHic5rEIfXPAgCM7DdsPA7bwVyQXEQjpP8H5
pZbXwbmTTi84CZZUir7jlzvff20BkiQZNk2ICZJgIN2wih2bBM3iRPVxXqKM2lWs8WVhkn3Z1DTL
L9UXQPrSHl0w/DP8iLbrIkDkSZUbYUOmB7tAnnjnSDnRZiR5BnmtaYwwj5oY6w6QE/z7EIJzxFYZ
frTDP4OfZTwzFljEoCHBHXGKEIqjRq3MSin1r0c+DqFN4RuYnY5kl+fKrgPn1Ge4aRsJjhfiXl79
JC8aRzHuyLmSdlx0YZBPp59SGqQUwttVEyNvYFvTDFzHeQ9WZ5W2igJ7oBLhmGXgcfbYQUsjEHD/
OjXuxowfZwxjvMUJ00Q/WRHeIukepYFkYD00F0gpFQVUOxsLY0nS3bousql7K9tfmU0l9yHtNi0b
NZlutuM3qYjnKeGrCdU7xEgN/tjRnOSQbPw+GcKJsXywz4NFS96JvbQWviKD3Q8gFSqUrEd/aUN4
uihG43CaTLKj8XIslR0i/K14WKPQ8gW+tyT1wCuGOpoJ7jo28Xgv8psQ2ssrBaZt0jt310HVkRpj
2+YMk4a9Ev+xZJQMfxf4ydcig6KUv/DOIaToIGxQWp0QBxwpsdi/I3W/Slimj/2RlCW8VFGjjZ2C
UDv71LzsG72W2DViSsSr5WBRlRrzG8OVdvypuwKfp9wUEIZsIc486Tvn/ir71cqO2k0en2AWlT//
z2EaElN4zjQdIS8MnW1CacO1S/cNZOsPVTodY014MiWzOQzSeByoKyPlgHd90tE54H5J9Dz/f4bo
nftPp+nVJQmD9FmRQVRfXeP0L/OA2GqXeOwDxvNXisf0DKMrWthEduqLnjQwAMmYqHjWTq6XgmX7
AnhdtGsH2JJ7reh1CU2MQk1IYGnNCew+/XlpT80pXVsV/hEHWg4RHyOxWgljPHr2oOReiswBpmYQ
PdlpMfude2gagCB/qoRc7PIfMEUXK4tQSE4QwwAi1jvcm8DW52FzVZLlpaP0KRjkzWHeJ3McE1r6
ug1H8N0Ppfv88EXEvnur6agvoSLCFb//e7F4VgI7QxasU+3El2nb/qYMgB3mkjxMLFmybrqLwreg
ptBqT7sHOo0d/3o5xNcip411Cls3dBRFI/qxJhHUjtzU2/sjxvI3o4DPbiSPGp+3KaNoIlAWhQsW
KWWUICjmJaphZUESWDkBj+z/iHkE1ssaz+/lefnBXbrHQkYM/ctNnGFBO72GOc5FbslrwSm4XHVA
pasmwJXjPVuhzPusTzJBgNyQDXSJaZCBx/F4Jes2HPcT3VTPMmImF77DoRAfGFuU0gZ7AbiAHW+i
mDilPr/HJ6dO8aOdKgxywrdQdR3Pleym3bnZs3+9ughYsrj9/KZIS/exvU7BdoKU4lope+2OfKSX
ARBccMTYsJp++8SntJK739m6ha1MFHBmKA/79gX84mUPBzrGg3uD/JA/XRYuTDAOjnCWbO6Aag9X
utHfLNABGOeXk4WdHE2GryN/BeL9Htk03Tm9lXBuXE+47MUtWS3cAvq95hnMk4EIioIvRnQh2S5B
wcOUXk2G+hiKzW4kOQgc9IWmLRgJQREkTlsJsWAos9g+gJP6Mt0UAxTQCzWYB8JrOXsNXj4uUJzt
M67MSLF5xvAxkOcw0ndUMxrcLshjwJ6WkPYbapCjy6PEW1lzzCtySGQ2LtODngtPsQbcwK9PNJfv
oUvz+wkbQUQUsawTSOaxPAi4MnDeR9/8IVZIn+MYObZn/3NP1Ic33sUx9csbDPjt3jdTmBxIAJFQ
x912FGmngH13k7AQ/RTXIl3Ssxc/pFhzLRUYWelgu+Bs4t5oQAKAjjVh0l2JloqhzrVySFyu5RNY
kQUdEVG0hhnLvgzvpE7dZRl+wEGeIWiVRTlt1PpAlK6nohOz4n23pcrol2uZejIG0tr77hTZ5rqD
6ro+3LbOh1eyk7/tVKi65xrXhq/OKGsDVdposOUwvnq8nk8Cq7L0pOaaYvYWpXyg8p/ZnQnL65hs
eVFRqJIO6rVYeGLQTaq0oZ7juc5F085ShY6Z4SW5DTpDmlZ5vTH9JmNV6ej0FrSqldlHV3sc8r2/
XaYoSIXzpJaK/p0UzKvdi/PO5a5knESUvcd2PtzztvLBnFfqYqVEoUas+mhcshqLfuLUFPmUW1JT
x+vUaiInaGjOlttspFHDOsheXoiXBpxzLSTQI2zi9zUg0rxF4ljPMxMlfHzqP86yxFiQtaiF8I7B
xAJ16yodtUX2uaSb1+r2RiYIzVUCRjm6mcSgp/WoS9uY0z+VYSVXPAHDatoM4b4M44VX/WBEs3Eh
WXZZo6Y//iHuAexSKQSVoyttynTA7D2Sm5aATH5tVg/dUBMz4+5Dzg/DaVzGiCKG1kK0fQN1j2ia
ee+ZsweVYAq8roL+qGG5SbWsjbUOyg+VufIlt574W6DaIbjOAavCdYjHzwvmYTQE+yp9MUsMaQI6
QDc2vV1HuTQVurEZrPml0w4FQhRcxlgzWq1WBOaUfYRPBdcgS4JJh39szY7jWJSU0ZQvbfNg/GLV
eHQIBdV8OHpUesGymJoOxfX6RjEa1ZNpccjeDbWDA9xQ1mkdjePJXSjlnkexl1wARqM5bVbAqr6G
zlwtHfCcss99jbpQ+lSTR1FZxXJT4C+5XBwR2OxKo4XVpBvUzJuKkVrW1XlLXACztIlmCAAOiDUZ
NroQRM72R/cSCXDYmVChURX1Uuv925qovsir2uotXrNNHGE84gY4mfjNecGmrmnKpCpYgFktIzCw
VNqtXLF4qCo/m9Ym4/AVBpCidfA5CKtMHiUnQrG/DCki9o3NK7zjvQILCsfu+b7pi0ZV3Kr1tEc5
/rJt5VmrbpUpL0kJXF1cq9Ee7rlbBxUpZ8kkUsZz+Ax9g6joSdf/vQHsrUNKvJYFUxudrr7zL1jD
RH5hoj7KOBABnotgxyFlaNHy4V+CqpKEMpsv93pxbQdu65cDw1K901bJI31xjmoPxjtdoGGMKESP
Jbe6rSTZpwkQPvSoGmBiKeYseqFw2sBA1LgkD/uvzoIgM9F/7DY4Z9cn/1u4hBKTbSuNCvm8+6y1
sxeMIVxA3JJOHtA2r0mapeg6mpmoLPcIh5cQ14h0RpKMxeCVzND9D9XnSPGayyhiO1ZweDcgpJOD
oCFKGdEqG2UfimE3fiwXJwcr6oRA6r7o6jQXaOeeF/iYQiG5mea+GVlJjf3GY2dy+VW3C5jRotEb
50q3gbcLx2rIEuZvSthkiesTjS7BoQ4vcXIG+21TKN1s9m/jZDZPW3z5qVt2Xjjgk7yXGTW3SQ7r
jRsjTwOmPDyKn7BCZjZKc46mo3wgR/XSbUA95efPqNe0tBBfs2he2nngqWcrTWHyTDdeZPXics5o
gjwI7SrLMXcP4hkLTNbZsL32o4mya/eYu84ZeXUlZjtca5kl64+dOjBhFNVSukbCpcPa1KFphHOK
L02FjpVyaK8YSGJ3W2IQmgOF2CDajeo9LgIYRQPhy13j8bYbIHI5xBFEFh08VbPasirQU++O2swD
a6v6M9kUkXibpgSA+8hrm6rMPaCihFa+9R22T6Uk5JrVv26h36Mpw28qJiTI1ebtbPd5Gk0JC86l
im11J105ZF7yyQTHrjJbs0fF28SV6tQY8i4FjGwbc99sT0bRpLEeSCrF3B0vGtjW01Vr8jD7Nzwy
bOwNFgI7oaNnZ14D46jV76EdEQ7lwqUV4M5rwudnp5l2aWrF1x4IKW7bi6LAH1ZKv5u3B/55wOai
BlKgDAgFI+JJzQ0QE9d5JoEZxur6CgMZ39g1bPw7orp64hWH+OZERT2F6To+ox46xFwhcANlgtvs
gWaUvLBh5RsD1W8P3tUCY720c5svBLABLNsG/qLzhmKVOGl0S7pvnEfPJWxPz8M26VEfbpSXsZv2
odA2uUl/U3WgGwHRh34N+CPzQqRIPts5L+5q2lhlllxzk2PSAX4qY43BbIdzckkGHReKXH3m4fIs
/xN755X8E9cl4PVnvAjv5xKv9efEkJhYEM2YMcppu/F1rbsJ1Tso49xEv286t6OC+swGUr4s4QUN
YpRHU10LpQJnh1HoSRDPejCT7Dji0XB0fCbPVWBCepdXK08F/FAqD0w4t4LfNO7BstWeDLIjEha1
7C4gzlYoUBpsaEc8sWvCiC1mbUsnzgo2o3VXC4frC3ZMaMQM9Ewbr6MSBhBJx5Y1MJU0tr2K8eO8
hV+kyxuPxVyCrtKFXGh4v1yCMNnlnSnMKmqcI9aZMlzPwQFivG7pAD2mUHTKEA+Mbon6iXENEI2v
XctYyoPvWyi+Whq48z3N9JqS+uc8+HEYeMzO4uK8p3pphQ5sHNzJd37mmup/btv5ds19t5ghgtfu
16NshHl8gTH3adp+UMn9edDUFh4pPs4+JhD44ns0YFvVsGEqj2MbwhhmLruApdSXuTlRSoE1RPWx
3ZT0WLP8a6bJu8tuEDGWwW6tAnNnaApbi8UV9c1/vc5ZFs24VkbYn4tWSLNKf0x+alRegA0fHEIc
YiVBrWnraihRpfDSbpubgHZ7b+XveA1footZfg+xoNgJDRXszlzhQPgiI+dV5iULqi8S+IVkwcpm
dS3z6SLzZIrAMMcCFtGLpuZhAyzEf3HqB0EsgTNP082x5rNqJ4Nyb0YKLxYQX3JztXi+8QxlahGa
CFQcMBIx6WybOX0rDCVQz+IjmFzGPqi5BKxyzv99+2hfMODXE0F0vy73wI3prk/Mo/RcPYT3/zPj
3/lhfqmnLpo/NOXEeAM7pHgSGG+bo/C5chap6ektYth+fc1c4eOrZkIxAOcyl+6REDI/8XYMQ6Ph
G7EXsQIUDPaU4ooFHMddJdfUCglogmDQVHRZqi/kIwSK1a/Wrh08uA31NENSQdM2mxk9DSFDTw7M
jLmpOZZBjdQt94Fb73Wny0q44ID8vvNlLrq7OtZfnvuCBC9dXkLVEA+rwiHIWqAtYiQnaSSh+EyZ
W/xaCLNyO44fKJo047qRGOcyWaT99+4XbLUOnz6a9LsPEMF0cbYarkFmS62/ZAqrkRY5AqNn7uKT
pQVsTPUYZUD7/FqFNTvxRSFuJP9UInO5ujnChcMK1vojW7AAMixKw/fAPliUe7SGqH0jx255540h
wld+8qLOt9mgypV21M6sPCHI7O1r09V9nG5TVrO4FJ62ltjFtEHwGqFB0hxcmPvutVAtBrD2koF8
Qf8GD+opw8tRWSKOSnLAkLF6vYicHt6KNadEuMyWEvrLogUwVaU22HPQWZeSNpm1GDEqcHyAkxPF
6QPrP4wpO8DiE4U11pmTq1a7afZ9z8z80XN8r/1Ju+oAXc4MNfRS4dmMbLnF5F2tph//6bgzUCDB
Td1MXC4VPcfJdLBSHjpI5D6jp6TH1kyjL8aVH53GEmXMP3c8eLEt6jeIN7taUbcbioibaI8o4LFy
qNxcRgb4ABn0RtaaVd7wZcAsUZi2bAJgNj0xNBR4lpQ7xTgc2oWyVqqrWzrFiiRl2IGQhE6d5kdZ
CrJvUqe2WeWc9Et8WrBp+FXDv6YD97Q8qUAyC1MvX+A8NV3GxuXfHYmBKtsHX2c7U1PSJlfuIngA
VohERZMJhjAbsAaOIrF1JeTGuWTg9ORdq6IxZM3cl87tcByrTrC+NUyC/Yo5HNkEW2kkLgWuxJI1
MzFFLf8EWbOwPoQIwPi+IG7uIZko8VkELofVxvIwHyaltKbuOAq8avfuGPGg7/nx60P/xRlJqwK7
1s4Izg/fAfWyLgtp/+/Gkc1luZJ5ekBbLdBUGv66woE+2MSpi6Q/gaH7XylNeFtgR7Yuiqa96s3L
QAkBcmqtj1E9dPUCg/NmNL1vc0wT9T0zXQaJDrk+iyn4wG6Y5cBe4Gv0ZiJ6LGQZs5Lb/4cT8Wkx
7jJgOKTuMLfrK4GYksPCZTtlXNkIKnwBWBcxcwLpjDqBI5cm7PBIMC19uVrDuJzz0F+oKEC4FHLg
hoH3+G+RNW2pHfJTaquFMfk5Crz4qq9Lg4W2sbyW184jbB7UzpH8hA96qSOq5KomVIuLIfqSHHY0
PgRgLotlSZYbwYT50+d7iFMdtkrreip3JU3id7pz2cE4dtmSAvQpzRAAlfarsy9gJuCFaoLAAC9e
2t9gkmcv49qfXXz5nX2IoKCGeahteUL75Hr0Vmq7j9rq1/7LIDdE9Kp5Z2DHsQfpo91AhQ8Fq18B
YJfVDTgRIJseb0EwVNHYFX80l7ikAc/0LHYFSuVT4LDG5HxswpKjJD21mRIzycgdmpiJMAHxwqt1
VV4L6v4FFj3HZ73O6Vq9i+0hoMuMRmxwoWTI34uzfsVcKbsYizjZfGiqm69gj6N4EVu1vQsq3irh
hJDLd2PFdRbzcBshUxHJ0Oz23KfbTv5Id++WPWbj99wo8Pfpw4ZCGPjbKE5emwKVjUea0epoAY9B
+zogzewknrX4fdShkH1HFQWLz5WGTD0TR3Xzxq/xGtxjIy2iqqPors8OHuhqAsY2rzpXzbgf6bC9
2ULU8mT47VU7+SBptdLmolp83qHh2hL6M4/m7T8VNfDveIRlFTQ20y0cw4wWdIAqm/YYRiaYR9Mx
BLwKkmcSEOuokInwSgkvO8LMBQ4kkgyE7HwvdetbcRwKO3Xgberik2JLHR9c4+SJUqhGZHGCLOYI
ehotVdVYql4nZ/A6Z87bYEEmrFnQD9vyOR19v0gBC2DlkYEj/LQIrKik+VsAuU6j3kCdq8U38t1F
tJHjM8Q+75ADodxeNQYMCg0/zAgjQjB/7M1WNnzckbdeyZDgv2la8lo17M2BZ9bBd2ICapaAHhp1
+nl2D46lVm0qY2M1oGQW4uLf2wF56qj2xWbDRPqQ0/xhWS5y95JTAgGsKvnSqbcYnM8KrWIIBIYT
wQjImvcjKv2R0/h7JEg9v4kAtYDju6SJwxcWUvYo+KA282P1Nj4eLQU2HwyxexB68c8UVBtnVuBd
eY2B1GIKMdlcD2eyREf5JHqK9GUUxELfx4/Pm7knwnHvrlKLS8BhpZA7MiyD4/ZrbA4ScL3COV5A
YHSDPYtzSTbqlC8di/HAE4O/kk7oorWEsd9LIsSUgA+0mNcVFc/iJbnru1rAp9+00vHfImnG9IIQ
ij7Snnq8FYoKhLQGQE7C1RT1nOS1ZKHz8fv81blq2KIaHiRBUebgk6MoJbgWDvwklNC0mE5vfHNw
HNo9iP3EEh9frVJE5W3hUU/CexOoRGX3Se0lOO8cLOvjBgQW90Q1o1TyGIF2DOKcB+oIz/p+bZfm
sUaqJ8Epu9xKtm0UJfm47xAV8Ziq/AaHpILwSacXCpBgTJrui/z3Z1r41ENMIaJv7m8edkAeVQpr
McKQCBrTGLyNCbDs/lJh9LyFc1+BCk6+UfkhQTzNRKmHt2FX2h1ERFxotYhg3yqB93vYsNEBtxn5
lWFSF/cI4QPa4N2EmBT4sLTwqCpUQhG2bhxxM7Muj6jE1/4TPDXgVSIZ/fXEBN47vJdbTtkXevST
5BguQB3D0Ci2ASNCfDn67AlszlGdz5rP9EZCACm1SvF02esi+Oq6bv5AtP3zNSWBPIBEgm283ANJ
tbHgYAIJLzR5G9hB661kbVTQGh5JBvJzNQ6olPw5J74JDvabDutYriBYFdnWcejUKv4okRR0T+h/
KOUcbsfM63MaABpiZeyHn/ft5La6SyHYSk6GMvq3vvBPfpGwPn63SSpAIvUHNuKDSEzKbQdw48YV
wORNNa9IWvZtoUjMzTGIvLDM/2z3wAJII1Gh+Ri7A7m8MNwiuLMfNG4PuFSshsdWoVA85QhmJnjD
6dm91vdef/DXpa7IdkvsFB/bn9oZ5ySy4O3cs8Q+vaDdRmnveB6HIoupQ29wZFYQiQiVA3+uRQm0
x+DGVy8KfOQVP8gu7YQ83scx4SSX0YZfqVPJfmz+ARfscWN+dli3d+yEs4DCgBgLbt8vmffE4m9z
97dYaRdhBadSIZJ3pQskDZKQyxiS6+RO5+5XbsKssOhCKzYh1dd8vV/VOm2IsPl2WFVHFBtUTNHX
BdZ0BD8LhxFJDv9WKSH+MySUmuBKMRqJdda+6m6BLvVNtO9DBkvLr8hFm6jJK7n7niK88L6xjBoK
zxZ6jfYlXqXiQBySVKT9y6qNuIjAcJSks/gSca6Mej9xB4B8Hmm4CRiQSNIqOgEr6NBvLGjWfq1q
/Gzp3xeAqi5XuQa8OE+0K8KeGXQj1VqaDKO2PnJ7PDP/DuP2hngqpJB4GW9iUJ6gAXAjaTqS8f0b
p3wqKvawpE0XUe7VwobC/ro3xPNPMWIZfqq8oko1ThJVXU7qvMDYuDlC8qpmh19eouebBKaZAZpG
5Nan2YkqmWo7qQvk4bbYGyYOf+AbkcSgpqbMWhFcok/IhPrDPuFRASBErnJsgk3KvpYb3MO9LVKp
uvb1dG1NDRe/aras37OVZ4kfcOEtapUifvhsTLWJ3YYO9I1egD3hW0cwWtDhRqY0kkmxgLaP/Nck
SI2Ld6ZxBKew8bmYMmz54JHy6jzKKZiLMyya1f8aGpstYKGo5871oB4DpTxPZWFbu4uixa5L1LFr
rddiT1tuztPcmLgbv7D7S/i0Sa/LPFOXgAuI6qks1Q8uzg3D9/W5N92DquJsbs2Wp5IDoZlxuuQc
SG6iQUjIBAkjR2kBZuqkp2nT7wFGkw4eQ2vD6AeEB+0drvCNrjGpSCEQraRC3/qfgTeJBTabJgVf
bWejcaANIaYEvXOkdqqC/U/tnaCIyCW2oCedIXIKMIdMLAsApsped1dvoU2MPH/VAunB9xbriTeT
gnzu70G8Li2h2pNdowLN8cxYk+5tLNkfRP5lw6iefCCvbwTjpS2CadNbhaQ7BL1EgR+AcommDQOX
X8uDCRCcy6GZGgdZroOg1Tl3iM4+/qEzFSy+MRPgyNrx8I7abk+AWzWYnsZ+7PVH9HU4lyQB2I7z
qHWh9PaghXVRhsT1x73X0Jg8Nrhvp7KlXneQs0Y8TVyOIY8gopmMtYhl8ezkhgM1xlCivaAn4JPI
RGfyuCs0ZgDiqOBGd0pweBT+BAUmJQEBqT0R241cxUA6atugFMc1BI6jUTh0BJjFtIrLfnpM3r01
uX/lWmnKbckmzZ3yVlPPvG676PPajFxAb4TAGY9/rsGOp5koszs4g5G7yz37i27iAuKwQopFm74T
OHh8kw1WXgtrSvuBPaPTBniXwKYa+VMPSJ0rfx9DefSFyJQRLrtjbFn9+JJkBBKifNbM0N6TZfPb
qY8MS5qujIJYa9qkotXGTpR/kTvuMU5wfWC/7t50knzTNj34LqkwHuuabQeOZ+2Md/WPHoR6mShS
dZ76NEccTmegkIPpivx5iJ2bp0QN59oBqG3SMCKHXOhFXckadP6/Uxjn0bct0Vq249PqHGk1sP8H
b2GpXhRE5w/MXq9gOUUEQcYM943V0EN2K+dy0uTt7l6iByI/yEDJBelzThfeXA8L/EvNb3nf1pyb
f7m3xEdAzq/rpPm/crSlwhRvFsgzc3OITQ+Gi8w/OIPPC51tkRRsgScvSIyJEunwPfjnGZFKozNu
/ht16WCSDFCLJC3bA0aIndoXnRhgL2vQQWx7LKLmh7UdDKsKIXvzvyVK9yUl1M602/ir6EyQ5PHE
nd6or1yEorRRw0RmBheBWavfrPAvLadyhiHf6yDXXwmK0eDWnnAwSf96bqNd5Hp0U8knQBKetMsp
6wl3K64E9jwn94ZRHf70PWVR8bg+i6ldSZ9k3f2kYegAMMGdw6xUXc6cVqhaY5296cxqCW1+Ha56
vHTSz14Gm5JNQvzfr+t+h8PzSAfdzsWbUsPzij7D1uv/G6zJOg7lpOhCViAZ9KPrLHq8IYgw4iHo
PsJnjxm5wN/paueAa7c4Juyx4s8ZUozQlZegoD3ErJxrfHYT94jXWsVF8tFuIn7CNQjuyYhT95qk
0Px5hl+LX2q8SoAlwbA5HJWhpE9iYtmu21hLRyo55uL4fFbhGikQ8vGQ5bc8/uTLWwreT0lxkOEo
whVjECHMB2oZq1WReU9NF/PnJZOPm1GUWUMqyfGZdCJQ0beUccGIG/E6Azwcw3t4Hx+xWJe7ecup
rfPUjFa2+u4PvqXe2BaM30pkltkV4vxSH3NK9leKhXnFyq1ETBn/Mr+QZQmvP/nJn6773WhEic9U
dHLvEQYHvPO1+PV2QKa2ynMEKUkVrSo7gqpqJizRTCCO3/Qzd+GTrIsv3LpIqB3NZM3BK0diAspB
BCJMksIm55meM0K7q3KRuwidfkvcfD/FT3s0Sur3LNFFN98Impg2nvLrt1re199S7YdGAy0fB1wr
wBa9V7tjylWNfkHF3NgDtfuBrM1DVvs666wo8C4uBh7ETPXXzHTENFZRijLGt11KD0ZPQM5f/EEK
GzdkqPwXQ1xwY3CB1jyCAsToVw387/qIw4L5BZE0wE0R3Y7F1D03PJ8T/zvjhW026YNekcndwyUd
ytWtQ2C4xSSuSnGumnu4tXjNfQTKXUc+531F8jjlKeG09zZFa4pL/hL/iOPPj7EusjEtyryTJZjD
wUYcNlWFTeeBXsh3X9wQUTMXu3AdmSrTQ6M8o9q8yA7GUtJpKfO2/gVaJ2fdKukZ3GwPhfhYgrfA
5m2seHpt2gsCABW0dn0Q4Apv4g6EauiVjmdjFAG5BnLXoloVSSfkWH3bw3DsSLj1r2ZDPW9e0PM9
JYYDn5GPgylGN8qvdOfX4W3i/LMT74D3F8igo1mAQGgik8eKbdtupXw59SVgxMJUR6N1/JP0VnYV
PGGVr45EXRXmlviow6QmbFOIv1zCog1WXZUyDZilen+Bt94ot/7JxzvROVfr4f6VuOccnnDhspmp
zZyRbpRde3VeivMoXKCx4aIK7uc7WMDOa9DZtaFdRkQAylkvPeHNbaJ92IsqkHF+FWmD7g7wwiZ7
XBJdMACH6qnUHbEAmcbX87K5HPoQ4uM5va+DYn0kqaRY5jPCO7h/Y33FkBj/6M8sYhvRKxG033uK
yb/zwparCHZjZG/CUv8suIVw20zHHdUZX3ad4Z1Nl5MdvIN9switwp9esz0FeW5Y4lIhMQBCsqne
Qi3WjG8sP9JMz4kTh3S519q3qINAbjUtav7ABbLMygpY/53owoKhFsq/W7OUp2yBHXevAO45/WV7
8qT7dLJgGuuQvBgsBNkZRTnNieigLE8Gx5m+2RVRZssBGw85e34DB9dTKPOlSHQ3GViSLRQO3VZk
v1QkAbTHJVbEzkQHyqkyWa7UJqRbYVPm0SykPzug2W3ztC4yC9oVDbMI2N3sSJsPdJCyIJJqDWRG
wAvv/m8MkcxLvmoukOMVMOI7eLcnWIhNsbZRGFZ50GN51iZNJhZjuhNyCkpqAlzwSTnFAt4q8tE7
d9JsWCdVJqZi1lMAIHA9vMPMdaQTXl1wSkNMfygp05CCiZgaqEjj4nHzR6K4qHJ4pkY25AkQerek
oAzLzgDK8pxdeyKkmz50Ldah4ehicqm0kyYeupV38Fw1t9QHdgTD+mI/m31QvEcBiaycig6tL149
E892OekazN22E2Vg5SiTzvtuc7kto2bl3rVhEwnUxQ+82fj/qUK3mPZtyJCxzBhErgvm3CNI54tz
V9oHLY2XaP7lDKjjViAl+aacmyVOcJ4OzI5hKx67p+YDJT8QG895H8X4yN9fzrZZ7Y3yie734++U
6AJwo4UFLbPbnDRCvSXpX7lt8NJtlxcqykMUlQLdp7jJnnVs4Q8vxU1NxR+l6Ka1sj3JvCsltShy
Et6YYbc8Wk171TZMhW9VMB6TqQcA9nrlMqA4e54CU4/2RErQbsEHk0awL7w/J4cdtg+TQXq8aZ/g
rzRQek01hzka4eVhm6z98PplcL5kPw448JGoBxEvlbF9aEzd0SWsxFcB23zdLDaHQxI9ibqcUkLk
7MKJzEJZFX9pKwI3cS3H7V0ncGtY+f9iKgS3rNLYH6UM+6Tb3UhS8cgWVQBbvm2qFl+gRktlnWGE
CxhfOsUAhP1lYvPYQzm5Z8+YczDdNCO0aL0L953PhsDcVe2YwrDswkWgqI7yjiCqGOdDLAETdK52
FZfxBMhnkHh2IxQzvrQmPIi7Vp+HYrB7wD9FDx9bzVaNeIYYsvida3/FR7Szehutce+i+AqTnT2e
V4YjqsnzlLKydmyGBOMFSJeiX623jcW7b2VK4tAOsuAxYJe6pPZmeOBrzZ3nNj12IvZ3h/fGkvbR
Z71PrynlnoM/rQbyk17krKkkYCIf4Km+fF1CJo9H0hCWze+F+CZRCtS1apzhox+2z8zHTIPKu78Y
hDMA0L/SNg8NztRQdNLDhcjuD/RQQWoNHN6oWhtdLua2sZLpTYE8Q3AMn/v2o704UWSlt0crngU6
q2flheVLq6mVuQEB0buuNK/Wvu3cNg+sJJMlwU7ZkrgcP/7G25ygVa3v7/fCZlXK1ZkrRcOX+Bpw
wgEGvdLthvkNgfOv8vRsoOOuMJowhLDYkDirXbjvvm2AHd3/+EOLMwVEEMaLzju0l2f4A/KkH+NF
It+7kImRUwC1W8smZ4/lXG/xFREDKw9hAFXsagn1gviJMpw8b3WS/8zg2PiNZvVzsENFufXt+u7l
Mi41N8CLB9QnB95SuCQ0pDrwOgBfzri03Bm8pY5JnOUGJ0jL8IizkAlf8EpJGNfDSOiY8GcLOCdD
m+0ES2E+3CquHMtIOBkLE/04HzS9xaIc5qFo17Vr9p9ZY/Y138JcRbk3kj9r/lqUvVWhvvnbKBv8
MOesoQ8Tz4lIJkUPFy/sFxOUvZi5ENRpLjqdFpKR2z0n6I1K+dS00hW4+jmjA6ETsiBjxtYH7XR2
iIZrMyTMvFo86XJijfr/i9LThD7D7gBGA2feWvDjFM0CZ9j5vpTNo2KbnmgySTccX5fYoXyu6R2G
KpQS+PUPQAludSR9qf7J4xBJ7XOjczlWQ0IHNusmHbWmdyMeWUwic/PYbuVt/947qZzZQZx/kEfJ
PUEohEPOO6Hyaqponu7iULJbLbI5Y1cwO+82NLRUCB9OIH+lcZTi1A3raTW8R7+hLZp6Dw8mrrYT
PGZCdEja5LLFmtyFDB7c4YAs/MnCSDN7gCu4ESLtcY3XruiThEpGL+se/y36haLk4aQJJqi2CXFR
39BE98a2qBD1bK9B8IjqiELKRUTFMSKknDHLMRBbMPzI92VRvjhCvb6yBeA1Qb3yjXkNrUFZsN18
zl7InTkrbhMySFpaNix2SXzMFb0sm13+FOqcwfnKUtZ4+Uel0M9Y5UFW7K86gNJ/qIDVtGUMz9vu
Kt9ojgdSumnnruXj5+DHdw9L++vUN+ybedGgOQIq6brwOyca2zEq6CDakPLL2JHRwlTkdGeBgM6A
FVocVf9UqOwtkb20tSWjRgML0MEbhqnUibtB5+tCuvNay1moNmRV+HVOIVCNae9FWK8uEUmfCyBr
FKqqkU7oStxieHEBsv48N4tq2dDibxpM0X5yzSMP/YSJdlp9SvlrMVCeJFPcjzb4w06pHnDzNOp9
hTLhUCbYVP6hiw/SDKsmcPpS3Hb8LaEoZqqYcMrIVMoJYlvDyPxOIV+oOG8wlnKyt1m2b6mHsgZ3
RpgYN3amTGyGCIICkc5mwX78ntUXOz9FuTAMxFsw/EKxrjLeNnlXzT2UJSzmv8COSqHnKybgHvga
baYX392h7xFc+UmrTZPVWEanMFSg6kDRDJVFuXDYOsw6/rwP0+6i4Hzb7SVzVNAThqyUfj1JPGWl
nat1MTFU4mPfvUWxLxF5aAgQZyAii83wZKe+hzy8doG8mMRpXcefsC4RMop/rsnGnK126HIDpUqB
xtr+IAa+a7kpmR71Kq43ee9nfQtDdKTnepspI/gYV/ssOlO68k6a/1zs0y3eaZ7j8GXlH9cQYh7U
IpveNLccgBMwXcmlFObS+C+jhlOg5AoXqDn+iMwzGn0KnpPJnSSvBJp3/C2xIKuXOT8EmnKMjMbx
atbtUqUTq/OYgplQimhIX1Vgx6dlYGYKWUPbDY59qJECP9n9czjfYHMYFZSldLR+MgsSIIeVe1ml
ltrf0lla3fSdgfcyPw7Cyhg6dzge3O30UBlGj0ABL0Avf9lVNNk3WPTM+ys5F2eg6cMv4HqGcAUd
KulNsMiReCcoxLot60ABxhmAgAOiuY9RYT9ffZkhoN0f4deMYdjousvDAd+PkdxD3PF5bgH5N827
irdPEgHdrhnMcotfUaBdkMOMu/YcR38GgLm5/5Xqj6ydfvRA4M36mXpeuIGzYkQVHHan+wWgDIR9
V0j/40O6p+dwK+Xfsibx8XbaO8Qemtolv9PZsxhe5/FNw+AtcUBckBwJcQHwG2W3gGEQmLXiYqKB
ra6upqxPN/eBvrSiORKbK8/4r7gPCoRRBh1q2ddl7FNsNmgDdBNjcHWA0UY0JFwqPuypqp9H02AN
JJGrN7Ol2FiRpZR1eoyQ6jGMn1hm51E8JF9ae4W0SdIwErxrrDW/TfbPbJYzXA9wlc9IJsndb24s
dS4q+AjpjnjS2TOGZanqXw6RvObAmk3V86S9Y/1I5INCaZ792ihOiw1xu3QDaPa0Qft6WOB4SR1n
qUF0/xwg2Ec/pQPDpGncIP8QVQlgpbfTqgO4ZK9Mx+BwauFyrlYOueLhC4/DycFJftylKImrGX99
hFUc6siak7BpdNpnFTpDQ40GbbKJ2FA6Q28ByORE+4QNLv4aZzr9fFwQaOYxG45IImcmME0+mspb
tdzRUx7kh5zguSsRq0+g17XDnKEqevGwjpYNu5JU3X0ScCu8nE984KoQ7fi/5tlUZks5BusiKAA3
ouC5HjcO1OthIxvCCFDuUjTX9QSwpWJie7Kc2OVVfO7hGoQWLySkmdRIX+sn1DezI1LQeBJusoMa
pZXsDzqm4TtXzjmkPGE5f/p4r+EIb3iH2gUYMF7PFvAcx31KzSbmxyf6ueB8FmZxj5TiwNn1mZPf
vIyHfy+eX+9hwPdLpl6hM+mfQmCInQ9MMkCjXjTeuLvodRrO4/JFRiIXOhJ5j0nlDlrbI9jJaura
1KuzJ6fFE0undbUeQOuRpxeEhRpILKDRfqXSV9ARB5EJ/eFNTmiG7GQ1kHVPj6NZ7LlgmmNTs/Tb
+43joW3N/MMKT4VvCULVR1N+DDvmr2muVf/wASdRAhluxjLsqLVdXI+vEGhUWvGXMFLsP5wliP/z
AG3aaDUVyOJPl2msw8ElnhTROppNxkYFLxT8sC1chCqD4r6Ol7yhqNpIbRZN7QgiTbdqrvgTvjSr
fEsTjtZqeaEAYDfZNCVWeEBVwVANwqcF50L2lbwia5jjUHsFx10ekK5EcR5SRi4yLcJPanAs68LL
YOdhxYqU3FqrDlKm4AcoivDGxnT7WMhN9Ud6XW8lR1N6CGQt/CVEPhjqr+WCBQVO7DgbGAl4snQY
ptNBMiKfmf0ePwjERW9WVGR5Q2yVMgAUWAuXLA40QTatVtHnxDEOFCfIn+FfA3xPcOHAeLyVPzXh
ZA8e2KR427a9U0XC0S3G3eowZbnyWqh+dLnIDQcHTJtn5sgM8esrckwalbqLOND4Rhg5AgRY+VRZ
ad2swmfyP3eHPV2kah+b45m9wA2n6kOmweALIbEoFZ3EXLnQ7unmIo2cQzr4D6opeNO5dbfzYPSd
E+4eTKSSbszC2q9WUMtMC/YOGTXr/leW8Rg3hfYX3GaNFwwtY7sgKSNu91QZy1enQq4aQqdNO/OT
zw3bvcxaxwGhpoJ1l4G7kP2ZpiAtS+Gdg99/Qx+aseTI2WIsNjHMQd9yF/uqYphyuRSsNm0w1p6r
Gxeq3tWlcTotovhK8MaMChdPhtyPkEyDJ0wwzyY4vbCBxU/0DKri7maMEMPZFmtFFYNoE/uVBw/1
gvuQjdBhzneUw75+7U50rW4noE/tXWj6+ecEpLgIPlyHMNzXz2hBWP/OlkSbasq11pAQv5W0hexj
HJPY/GSi1Xvwf9mSM+dV9EcpO4q2j4BxURGDx3EU3KxBwXz+7+QgTCKXTQd7fI20mKWW+WTNyGdM
O3v0ahVwd0yXpZsyawkD7RUraoxwOwcySgeX/wrAJKCImv2rJxuj/KQL/DfE33hrac2IpEmp25uX
xrBwL78/Ma1j61sfU7WvlP7qGDqBpbq69wKDYK/9h9JtZgb2ApVhOedLGDUfL/qKMW7E9q/GQhku
j7CVJ6OUfZC98ROG87nBVUqdXevmsx5EfV3DqNx+j/XXaWV61VYGl73BRg0TqR2Fd2CGkTm/PpKX
WI/nBtmfHtgcmQyYO7F9hUg1zOdF1tijhmIzChHilVaV/qS5gUq+PM+h/x3Tw8NJERzEKSu0D5nE
KvDPussFVm61JxWBzT5n8uGwkm1c5SqYZRsuBdC6mfQZqMPeQtcoaB6XZnHVZ5guiCsNdrojoPfx
Tyv2N5uKYqSYsKM4hJsaHg73849KdPOv0LffyFJgN7urDEZXRGdnstjLoQLBU179uwUKeXsuwgHv
cB4ep0KgqsbqCx2nDQwcwbMYXt5dt4lhSyLl8oDg6bu5FnpvNHGiLuMawDrXWn2VHF3zykpubVvB
a1soFsj7wyWd2XGxPaLJKG7YfaYFCRLwfy+Jtr384QoLih2iAcpcxPB95nmnr/wKoZtTdLPVAgLI
7vW4RbyzjV29QIJFubTO3qG7tHHL4v6J5fA56bs8OwHbwb1y8x2/Y3T9vrU29eWDQzXVmdtAOpW7
yX/xDISIIK3b+EuUWwFujvgZQp61N672uaTNMUjq4T47cw/w8EsQ5CF/d5xTJLpi7dQsViTs1sog
mTZR5rw4bH69m+7Xtwx2km0MB98PYSr1jLLg+gOf+emESFcHVk8OJenNx6hn3cxFWZyzFV1IcV2z
YoiTllAXPV1zq/feGcSgNJN+BvhqQcWMmzooqa42UuzWARHLfECwEqWY9zVgiq6p6NLgvfK5rQVK
lX7YxEI1jqLraDj2RnwZAOZsH0L73GXyst3m3TrnylFYrOrzEOSC+LiyRU+2Qc6AugcWUetSAqm1
EsLW8Y83YScFL9kY6Ua7UIU8PlkjHMekj9YSzD3Iz0YTILWS9zW4xeVBZ2HT1AWqTXMYStw8SZeK
5Ox1E0GzBcrxtXkn3pXD32tb7qpO3o8HapAPKuvW++J8v3d9+KYPsfekK0K5aRRNJmpTJlTeauzU
PT2rd1FSraW9YiaMAXZtGMC0drQ+Q7Ox3nqaMsyZCbCnUHsM67UsxCnNcb6Ghoon9JucnzlVeqLs
cgYulcvHw88kV1rsXYH3ofweQDvuLEsOCINNt7IsW385AKdowxwyaF9wCTCjsZ4w7D5veekuaEmF
XZDOlivqJJNobUSAdMF1Wok0sovWmysTpAGUd+GwrBWx9zu5huaUk4VcwAvMTl7sDVcYns3SBG6f
8H6vjqzR0P5MsR/145KfILMMg5HIE4L7XZPopCHNd0YVEUTlNXb5HF2rutteQbnD56pSPMSRCYs+
gIF7dKa6RMmkccX991zQNaPS75P+rhFehaUXsCSmd8nhCuXCBmBLgZgL7u+79kr6SxE15emW7WmA
QN28T1kK72ZV4MXMxhDv9RktXpeJUqNxxx+ApTKDlk+aS2jHA8d8d6EpYPZWeqCqT4Y7qe4eoz3t
3YLicfqmIsEJqLjME1hDKS0sPDSCmzC9PuJhEpszI84Krrz3Zefu8Lj+QfOhx+CJSl1tR8WB3ikT
i4Z1RmXcZpeG04sGszdefDxIxTpXFXPm7njAZKpwv2rWvfZ1zT0lClysFG5x0gSXqcwgAC+nf0yU
tSsiDOsIej6xMgQkB2cuhLY7UKBA4naCkxJvGtTyM7bdtC2YC7xmah460RBbdcoJn3i6avERQmvD
UZEs65Ps0ENPEASLdikDZt3BI8kSvnRVkf3PdhmdUcopDXC7w2uwfJxHinE9T9S0u5kbmDriW52i
1LHUBm6vryMmc8z8kzUGccG2a3gtVJ1+DSWKdx8RXPmSOcEegcdijiAddPWsoS7N8Km1G2N4yszf
P7FOx4kHhC7ztLyVNznF5KCSMDDVyHq66SRkRiM/uz/jH6vNhu46qnmt7WC/6JkAdS8R+He9JJx2
sqtUGMH2aKNcbN9CFHZp5HaURZIZ2EY3LPJCOZPhc7el5B9t9YJNK5AbA2BFxSma4R0ytNbiXozN
+jp54KHOv6dC5g3+XaFN3d7FzKgq2GOjsquYp3Gsx73TW6A+p+aMnoZmSc9xg88ZvpZaGNgAAnlL
xJMDZlEo0Bu8LxM6yMt+Ud40egEbbOHSleVgWrNJQzgNgY+UCEk+dLi9SSO+uEI2hAUKQw9jFFS6
oQWnqhNm5llv//dHMYvvV5mFnTYcZ4MqZzx/YeCg1l7T/6/SSctz49xdlrxfqb3BDlvUjSTL1+nK
CAl7zC7gEoREWWFtu7huH/B/SWe2EHQEhIkFKXDPibYemYSGpGR6ZGby9V+lafTRg1ytPSes+wTm
WjtCniQ+P3lb8UVcIzb8J/PQbYuwwsWhBAzXwoPE/i6Zx8Aw6yVbdlYbmEj+7gRsd9EUBWQzUOru
LHJ9CX/nbxhdiE68h4XEHg7acJQ194/l2I+Drs004szaSQy95vvAVXbwb/jM6z27QHtrOHCAVr1G
xuD02Lvrx4xIuoyWmkbSy42MPBxTTFIYYUpekzSeI2h2499QjQJoGL/sOUxMHuubnyTX8A7vhGtn
h9X0IoFDftJTX7Ga80qqoF8Yh+RS8Enhs9lRllIic4OWagfSUMns+4AkXUjR64JRhlzr5d0bNeGD
JK8GojahtujmOHkNZuMRqmbuSSYAo4tDQbiH0y/QenHzbyGeaarQfgKnhceeQI0EKfKyNigoQKVN
oawtGk/pvTdvlxxA/AJrLhq94STf1MAn90hRHHZsJYLbHXVDmZbv7WD2rzxruEkriOiVghWtlLTn
zy1HYn7xPXaFZ0VKNbbFUEDrKfdxHMp4pab9GlxIdth8/LV+h6aL2GuP5oYMxSNvNgG1GIWYVDSp
DWRaOc0sdbrYNLMpJ0trGePTlpEKOb0PCnSuGBMc+UDPXvBEWVeAiTXVz4o141dWQEg7NqMOvuvP
r1Odwe6dcmWo/SwNU8AWnk/f4dRn0Ar3VX1RsPY6OfsgWEZl4icJFRwZbvw61C0EDxRFJ+kMIu2u
5oFqfk4GgYXVBz5JABjUIojBcxoauzfN4UaUKV+rvufYUQ/zAv3pgCMng3VGGlmn/qYB4IWGOlnF
WED+BhrzdoMilPsyHYklPNUNjte67ARPe60RJx9eXQchvHVQl3WyyvV5aEeBtW0qEf8KCuPtEs+q
ntyxe8OVNtYigWSfXxJZGZy4KhH/xW87VEkXUNUo28ZfHa3Z2nn49AkPcmGILXbkVj3iKu34da5z
2/l8RiSubXdwLi+pdZR9sa796xHQ2kPqohpz1CEXp7cHffKb1P3YayO4CAY4LUJcb0F50TVwQbik
NxBaBys3O5VSIODUox/cdSkQyrO4PGXVu0g+suaxOfnG4Vi3okrfk4DyfyXVGgR50V0NHUMpFa9r
X5qqBxDlIvHJc95isdU+LJgf9Qt8Utzbyj5EtDq/Zo2Zup4rACSnC2K5BW/1GjZa9fgUeZQGDbQE
mY+hniQZjIy3rHeqvZRnywyiJ/+o6aHKWRdxP1iCbpVwGASORi59GzvYlyNTw2wWF554STYll2fw
rjoxpfVf+5evyI2wa/jfQ0w/2Wit79gh0wlpnuDezO+LbWLnEu8W8Nzjl7W79ggam37/pNlpTfSu
T7MkzQQBB72Nt3Lm5tSBZpVyZa5Tpa24jPAmdlGljJEUS0wZHaJhfQJ8DnCWOdZWl6UiYAJSRLWJ
EN08v9TJkrMEzTDElOeJkWc7Mo/6lQ73gsGtIUqORXSAO+f1OiPGg5oDneS3jK+HWCR/ydzTPMte
FG+S2s5HW0jDloUy2E6zLZih8aUF4IuL6PlxZQ2sWCS7quMP64HUwTQD1IdR8Rhi1HWsUaFBmd+i
nykFDGntZfm0o4cA445yELThC9Njk84lytxE+ufJm4Xif7VaL+9a/tQbxDYKB4M4CvM0AiRNKy6V
A94TK+aEaahV3GGOnjI4asDbTgps1m/g7qGJIhBofKpd1ks5KbdM1GZPsUhJytSoyr6pU4fTUjF/
ISCr9aBejJiAzs2D+7ywDCmL242s7WIU/8AVlWtJUKouREs9zbCYuc79b0kQIwp1jBrM0nVPqVLd
xGWZ7SB0aGaQpLSqxP+4zjfqKRwnpyV2ByEovuOWzomcgec6tsiNyngwHY9HLQ4H8KvslcLvFPn/
vxXtypRwxBgmVUiq0g5S2cZO/S4IDLS1ww0eXG+Ns8pX5ejTybQ9auARFvTTzUFYxChpIMap0owk
wDVb8lbuUS2BP9jItUWfxezYTsestKC57OQnb9raNFf94nyt3rLvylp2HN+/1DIUyGSFpfNEZIfs
byWueaQcxEyCVwYbzuQ4JZEb+Kq2KD8/LsPjQ0l316UO4T7xyObxeM0IiDlX0gzszo3uUkKGyqAm
hTtdVprkjFYKlRoXn5qMg6C9OcscpVY8ly03ShSEMMmoCxUTjrkM/58oXckFuQpLFp4xLJ1rZGGo
9ZW+hCO+ld+2jTjLeQkrZcOUn07DD4FH4Hrv+TGKRbBMec6xMN2FcFVITnyouW744rgD7k+2xST1
hAS82Cu6xedRQ5fCvO3AvnRw2rL/YohypRct6cSmMK22SGxFJhSKKc+tuZb6tHfLPAsO1EaoUGCY
D4lUWORcQNlYYcmrsjKqXSGe+OTYgE/kHL6toFFhhlF06jrN3KgD1AV5VAMg+PZoCVY13SM2HhuE
XB/J12XREcX3LqauOXNw43UXNQRkHThCsRQjnHMAVMu9LC94Gber0+GFtypJNp8sDsxYo0XMlb0x
jOOcnWwLiS4N8DitJY4DfKgIl3oNjAMfOUCecNlO+eJB8MX4k3/B3QnHHeM9S6b4fEl7r1EcYciv
GMZHpzxmy20B2yKG1JNPClKt70lDPgKU/qnL1m91TFNfMtg8bJ/H37ybv9AUtKRZ8JKgkncVQbxQ
6URzLC9glpwTIJ1dMkKmwSU8hOntSwVMymY5C9Qq986kV1y8nJ7PU9qCBtgfEjTDJtSOcowpjQP0
xRlWZO7fzDPOCj+HM7WkbvNy5ki5pURPVXjE3subGbL0V2oiYkTuSomlicboOy/XkVR5wgGkQrDY
X5pnPMy1NDhZDtZxuK5m7aqskRUiFoohYyqppnZsJmiQbHB1tsqBGJ4r1bVp2x2Z18dmjIfxcoi0
UxcAhNfbW8h5O0CdMp3njKGhg1tvGw9lP5Zmzmjs8R+Ow6pnbYDTOZuZDNSyMUIrlWffQvfDOHvb
KB/B5qNudgGHv0cql778pWsxP1H2VQlAJ3N+MqCGRSzc0g/+SXPS0oszGCYCQaVbGo9GFx6RFYhT
/cqzNlUXDpl5hr35Y9DtpQ9KhwczamkW4sK6BhyBTAa9bv7Eum++lee67qQb6sWdjF7KcuflBSCg
JrtpOeair6YyD82K5/Qsj9qTK5uHIimCEvdP6vhEt6Ue/7eKbj2OETdsetbFi6r+woN2lGhEX0e7
wrLYZT9MFdrJ6YI4GbjnIZpaYfCBi7AC+DLm4vo9Ag7e37B4k+gpSPr2yC2dbJL64/8FJNWjqUjH
anJR4YzI9lyNHz0sMjsu+U0oOQq5YDJTLJApcwHC8JL4u5iYVDOAm7W5fYZah9QkrGv1bPjUBw2s
1w8zkkFCw+6m3I7X544yLJa1TqEWUozEkKCpUXycUpk3W8B/kClBrRLUIh3mD0exkVLfZwCrdRbg
X+pqqeOcLjaaDfV42e0g0fiOg1yxNQje4OnY13w2MirEejGcPLm3OLohNLdO77Ph8IJJxSLw4Oie
rkGFxV1RWu+HvMwmdvZmQSowDfrv1J1ZUSHhEZHF2UBkdGMkcblBNjBRjtoSDbfZGyAH/CmEQrRV
q0sklXIGgRoGwWkBgoAw2GG282ZOdxtOukvYKQin+W2T1kg34um79vQJpOPZ8ooZCHWkUOV/X6bY
aFYC43QTDxjvCuGxGNEP6MDW3s5hO3nMkRRrCRROZJA7yhg1qiiCGC6DBRqZQjHx4/N2+6uReLT+
ONvgLUmk6XHzpnlltckPmiy8AO49RIOkimccSieuMv7jzaAg/9ZWN30mBnaLbycUIP1U1bGM+PN0
VWg9xAPOAgO9GxurNQzo6VQJL/KFZDx4ylg4VE8qpAKrcW8LsBGgAA9d3h0ub/5ZIVkazsVe6dnu
p7mivFEJCMTqDwDHT+Ukkr7SG8szWFuHi+HwDeRiFa++RIzYAhAp5NUPqZ3M8NxMGGO6W+ph6/Zf
wm1NiCDaLBCpTkuJ8e5pIavhTh0kbTVyYfQ4qM4/3uEbjYz+Umu+2IvFA4C3eMgjg36qqawZkF6Y
zIgZzjwBmJHrpZBmDiFbdlsU5lQ+NR+OwyZEVDu9GIHu46RzHJPnoHGGJ5GcL6CFS7qS0Gxl6RSw
oEZeMtoABPb4sF40i4cvTeLSmKOGBfAVSKZNmJj6tOJIOD0ug+jDvShxK2QiqGpr00UXcQ8KAqCI
6ogyZgkEw2kar02SIOpHW45TZ67HiyC/KzBs9b5GHzhcBcOBR4e642K2B8fEslD8bG6dyj0bf46c
XBGEH0UkUZIkApyTnX+YxHI0moyHM11v5ak6ylqgJYTiAcQzy28TzSJPlXcUGcZoaulnbqxep75i
8Sfmsl3FcCEx1uDDKnEv+MC/Dl3WA8kVJTuTmV2wpSMwp8GWQHefGFj16oEjpk6Y4JKNiOyQs0pc
7ScgP8XZBNnTr4jrrA63RTTp1fpvNfnMXkU9Hagmt4yTavhvzy+dA+O6tabPnqlTuW1GnNH5LI1w
q3SPhY84dEWqe7PVkmxTnMxHsntwk952UqlTyUE77RJcUe6hnls1jE3yNd+BE6Fl4zuyBBuNTtUF
PjUnyqeRVqGqW2Gf6GRxe0CnLkzB57aeL1Ov/9Dhb+ltoDQ6g/HBP0tL3gWp2i8j3jg9nWaITdDt
JzmAUsRzxxfl3pm1kzaqi6OMmIO1wUH6HPSpULW1M/eWjiaXT1lEk0nuyzv6IGOmyE69py00sDGW
dxEGZGCsyRhGBzPbztvaHz0VuhxR+Y7R341TSWcJ1zJmaukhTflmBarO47ozxomdXogtaAQOP1E2
7CmmR7w6QqW9cPHZsFFuqgAuqx5DAxk7AgqMnI47/KRmSPBA81IQJcyq8yKn9iK9frtsDs6bwOVv
61oA4JUs276DLDbFWZ1X8QiCGZYO+PYjIUvgpt09CPeJSWZYhfMNGGlGB3ewblDsXMX5ML4GI0pG
oEKETxtwMsOtT8cohMPrsGhELoCqauPYWtHknLUaN6lZpgTFOoHUDI/n6NMsG8ckwn041mDYnbHL
fsJlbZcBcERmMJ9eaqcQTyWgtanugvllZ/JKheCMf2oauS6Prxn+o26ADDrLkLRcoyl94A4NtDZA
rCIiNAw0ewjrHHws0XOgvj7MBH1yuXAFEM5sGNB4Aoli/LM0S3zRJtnPN+G6vjXo37+F62ILz5xs
alt7Cf5eqNWn9LletxfmfdieHMfoj0xqw5RXhfuz/IfoDpXgtrHDzXy88sJmBGzxyqk52Tqm8P8Y
jubIbuI4KsdhZwF6YqQfjX+dOESPUUKxnUSM3v86keDkxeBbm2QJulPGukbcHJn05y5guOhcY9K4
iUyqcAdgc8MeNxLxyxlbV/XKLpzzm56IBDIdvjh8lYKksjHyAbkXx1x1VZrfNKlcQPAYKnBtnRhV
xiIOeH6PZFa4Bp9yabyahlfObpllbzPs4KV4E5W/KZ+cJDIkG6a65bbsIHzkhTqEfFkg5YLAcySN
9KT39fhwNhxbj80XramaXPBL6qA7YQ3AeF4a2kCdh0uCUapgoID8DLJgM9AOlNzB63hw+f8PjveZ
cyTx7tNjM9SsMnPSxl57hhxyxxUoBG19SKMdK9V6sWRk0RuWVX/XLoMkex9GwUxSX/s7C1JMqJ2P
JQK23yZ26bwvE+acRtmk191DWeqGxgGeqQqyfDqakJzVo873aHeCY4jzQX17+H30AZ25i+BiRJQb
wnGXb01JbzEpKbns8PXgDnaP1cBd1SIK4RxOOvTEEl66MmJkTd2p67voSmUpjPlWSvldrgeS999M
h3Ovvq3/ZgbCgN+TlvaMZ/uSM3Vq3hIYgfTg2cW5CLUPhK/UodWSejGw8SRLNNIOSNaP+SNLS/3Y
m4kAJZe3+3Uu+owGnnaYCd2glxVUN/h/9lksWnn5PFk1llnsYnLYFDW9s3ydfJvLaIvuxHWT8KCr
dJsiwGbrMmPnsdsAiNujvzgOrvfru44W3ZYqAhv06dsf1D7klUMeCX9KWX5JZ3kZJmS/PNae5cRB
80qS/tmyuhIyLNKTDgwcEX1OX+qsjm+SuLfDiCJndho3r3RbuJYKK1owILkuqgU76OaVrW1EuBvh
opj1iRcHHtD2n6ZMyVDRQjUHpKGHvDhBKOr5QYrwkOnCZdPD3swji0wdXKQZ1rNLzOohDkkioIgo
id10UFBDzZge8KRB+mP+nbW6ELfq5qsEoBRNgEfyN95zDUR5oBsmc/tvPXbEy65HNd8CnEergYBG
Vxf4Qv+qJgakHK28u8ICC3P6AEFt0cADTL7T+tX8V2jKtpRHHLhONkkfH23/JHRayWCpqOitL5PF
Ortbf1ELAo3nlQh8NbLBAU++xESFft1jv7T4f2BWybuDvAMN95SRp+JaObD4ktk7o1PEQAe5Zs4L
/A/5BIsV9tY40VCRgjO4hSwGMs/ig5rOi15vBHeTBNHt76qkZtuSZPXhUaDQdsLULEVpsMNDDWEe
m1PMgG/yahCThu7w3oKMmoxYkerMx5hZhw+SfONt1/UvUYN6aZREDxflIO7Zuub7tXLQaaQvUytA
2OuPeXR3psov0G7qVcKhy5z8Llgdm8/0v+IMvCToR+87PHfGwdvStSKOWkIDp0BRf392gkPpAyYw
wOvjjxufDKFt5orbUgMzNtw5JNua2cMh/g472yUAbiRqGXfoTzEbcQ4HIXkU1pC0iswTRsTJJOO7
4K+TYvByZYNVGIa25uHhCTWSMeh0zMVHReIwBVgHUlIMqpWQedykKq9C8b7R2K0MxyDJdKA3dBlc
+DmuGMesYgdJfhY5g02KIYz0SI1JdwIRjhjhSgvkbRmhiWy3m4YXZKvo9Vxul9DoMnzjRxtwvAg1
HtBkZGcxOvgsf6SO8ErwjNB65eesJLFe8cSXLx1SRlPGBSRVmkK/CGSBw9wagLRLHeBOOzu/PCcU
l2qjYLEDbchQW/pSqy+scViWKFWCGo2hfC3DKYhzmWedBgaHo6ol9mS6Ump2bDFSDzlcVAR8qG1O
0Hagp5YEh/LMmv4uVx+CZX4LuL1ROlfvu0zbryyx9zLEDdxXanbvsQXF7LkyWsfxemZen9vwkvUf
cGQVuCcAzZiPaa1aDUe+zN2BmL0v6pb6n9LSiyUw3cVOjxPPu9GU/6wx5rXj4dWZepBjq8xtPRJ7
kWS76rgHo5V3Blsq/Vcu8oE8RSGYkyyB/frX8ojsoiwi1ajls03MqIiIwA3ZFnoayvKB8eGL8D+y
QBcvuX2rkg5scjzsaGAFKC3vFcFuIyg2h7qqlS6FBSLsstOrC4jLnRUms72EV95CyPA5gv9Q4Ze8
nxeYS2OPZNTb4qqJSwMdaDgx3O3s5ws1W85yyLaGAThWRZ7doCzvgwItrNvSJVwMX4Zy3GmAuSB2
CGj3KtWYeJFYI6X89aaXEu9uyR4mMhFCh1II/WNgeMqEWKR1vRVga7zHrSLJ25zE+prYI7cF3ldK
7E6Pw1J3T3T+9SDKE4eSs2dK9c7GGS7gu+mPZxHQqw8nq9QPmF80WZkeFC0ss0HAd9173t4L8N1L
SOtCoPOObWx5whQd7dTV5wQy/TNCp2yJ/m0YLYg2K58eqCB95Fvt1lSNavebDJ8crtGLXeWbpWLb
mnECA5QhePg5jifpFGoEjrdKtEXRZ7EOcFf0YZZqVs883OJ4t2kElXxwiD6ugbKCvdYjvNMZErsi
R+ZRmnWEoLQJcPU4MdAlhTjlICe0wuC5etriDIebE7b6f04cMp7EE79r2St9t/cFd6czPu9ghOWM
0+VcnG6l5MH4GGrVzUzkf4y74GpahS+naAqtDtCT77nQQ+Q0iPrisVYKxhP132CM0hyWBvRl957B
HCYDGFSUr3JyeT9SiUoz5BfKlZMu4DdZ5JxHiyN1dGdOgN4V5rOI8v/8oBUdrhb+18vitFpl9SQm
QVk5vDtuaumeP5dRQc0jpH0a9ae/MlkgDxRACmdFiHkrOGk0RJMO1q1W3VlJ+ILqFgzo6ph4T8SH
eNR0WLrJEgXPvqs0AFw0I/FVzuNxxvtlbV4lIHXS2LJiN0r1oZabLikVv86r+M39O8UKdaJA0pix
vd1b1i4veigIvvKJ+R+XCkKnU8/iycg6pAJee3pXLqO8qeFnQgsf3YkCBWW3OSaRfhEnB7H50DtE
L7waju9gLL9Rc8sRfvObZqB9kJrmC5+W6f5ad8oVTJOyY7l56gS7+hd37qKqO+uGWn9m9aUpM5/G
rxPvD9Kw2hA4KinL7FhAT7SdHv8i0yLT2YS9konaIqhV2DctUyHaeuibNRzsNLvRbu8SQ2+dZniP
yUCsszIkWaf7RL0sZ2QLRTOpOXctt1UZuMirfTjs60rBluXRq9Vx2dp83sN+ncCD1ztyWgOk7wRa
izjM/dMKBK8CkcWCaYHxALvLrfmykU1VPgwYbxZtr1r1d7dG+EgUZjfm5TwH3PXZldcho4S19Zhs
CGbNfB7Zf7vUO+PUK0b7QnEpJCoFXUN9q8rnvBDfh5+O3ygA0eL8WXAdNp7he3XDP5RG99ktYAiz
QcS404xgwebuShCYZTxCMWLMUK8CStMHTt+AouUuhLl/kzGj3RgUD0schzA8D9oaMSnQhLI4EKgL
nyOtZ7c5aGkIz3X+ZyGGDH6VKhdK1lW1+IsnZP5QB1PMDW52GKgr7NOmtQRzE+yLIh0zFK/qTAd6
CocqDCnODPR1DFkTgioTnnEev8OI/wQ/3NOxFctjE1tYNx735L/TL+RmCWQATZoiyiMGkyPbR7IS
kipmz8WyFwuJWCn/uTphSjZymdxaW2j28QBG7OBtqQNEZcY1+Y/kfbwq1ftVEZxr/U5ATfq5aeTk
Bk8NPystun38ynGlg/7rn7p1bx3EtVf1igmQnTq4KgR2QeJ0wHmfkt1flFYjkrPTvbGXiX63Oz6I
F0mhgFFHOCsWBm0FGfxc2FN6LplFonQccFOaxP55YzPcW4I9Asdz2mhiuKAm/CK7Php5ztVdrxfh
d1pQYEv7e6b8EQlvJNV3LfDyBFPf78alIK0q2o+J1ZEZxAKOUQiCIGunkbtEWoMgWaUaC1X/WT9v
3X/QgNyVWGNhMpNGkzHkIiPkinUVO35ZRsQpMUsHBjomP28OeUKFsXgIZX2OkSrjD7aiqfAGA07f
lmpR7TGoa/fvASaqilpAemZBkbDZ5hk9cOmHRixjDnIGFLgNSsmHtWlefwfy57cpCYfaEqun6zdP
J4Gl7R44qHH90ytfvYnQlbgKDAaRDo7BshTRSzrdGjnpDdPbNJRWqjcBMjnunWsZKQauOkxjQEWH
ZusuebeVVfk8tf3A9HpL79eG4ct8rFUYfsRehS7EpPWll1vHAh1U2NHQqfTGaKxwKaZD7SVEqtJw
qHT2EMVIYAD4jpZas3Qe2xG58SHTz23oP58jknHP+ISkcifVZPgXX4bGvGXQDcbwWrR3bF3sx47/
8+PceNvwg3zRLcjbRSCmIhTF8DhgNmOsNvtN5EzJosOB8qIOSfAswcXbiQmPFQOiAtVCr7s6/YF2
p2ipbTSNueTszY+esAXF5oznQK2xYfMKJmdBMA0P4e+xMCrBMLxNCD9PBRbjDSzwp1Af9Gy3ezES
JMQGKnERLktqMsggpCDXRMoQEPYEv7ejmUYEFcnFCE0QoeK26lcHA4c+ZRCIeB2ZsPONzAPn7Kgr
t+iQW5K7NT91ukCrUCS2QBVB5sC9wE0TUeuWT6vloL4Z+/ngMC2rkY1M3FtGbEPrWikpcfTD3P5I
q5J3BFyBjHIZSdOUMi33LrFRdSYl6GlcbsT69vsZgeARdrmf0rin9ynBqX71Q296Aj2o7hcKbXTQ
rzY2eZXoW50O8ScNWEHiuDirpxyc5Mev6dg7opcRAtWu/iSGdwRZPjPcMXXKDcYqQpN+FdBPugNY
ppQMbtI1bPgNLOwbU2HSfHDSrDkxzrAy8aj4YjqyF8UJZLaBs+Qhd6RDJWNOfvZSF7JOr1INHokO
Rchn3/L1dGf/Za3g5owMePF8K7FY7/FWJutJNEaQAhBc5gaY7FabU2fL08/BaLVojwyHbKqc6F7r
g5w+EY2/xPmQzJLzfksQFOoLJEZEMGEvcMM0j26O03mIjM4i7Oar8OPHSoB7fTAI3vkYA1FLD/Or
quB8+A1jEyvnJZ6/hpvXvEIlMbp/hcXMYhxa2k9hc7nr/CN4xblTjKQ86H9OddKHcEL/3DxMlYyk
ZhioBm1Meomes8FHWMbnCdkenSv7BdC1D2WA7OazuANDKiFdJqkAfNoftd9fj4x6DPcdSAqyOgBq
W/aeMXg1zw062AIKak7zMuSrNX0+q2+JgwkarJpnBBYECWT3rxv4aFcZq2xwv5vZVBd2O4uMnNzT
wOWTvr1UmMNhs42wKM55gYz5as+JlcR8NTwVa/NNPXavtE0uLJWAlAAjNfplulOfqUzR3XthgKQJ
XT5Q9MbQ7iJOys1lBAWmduCPVFQk7POeE7jpolAWCya7nYsEcmjU7W921lxuJ8hWJmFXkSG8e6oq
px0/sOzWjrIpTJwTjRF2Qr+XBSfXcWZ9ogLjl28y1s2b3CUBX/HcsbMdvRcQnpmeV1VDSsMC94Ye
utESuhT2vr0DBEPlPQFxrs7KRZor1/Z/8+w0MLcQC/sxpgFZCaZ53GmNhDPdIbQ/HutrGvYHkfJ+
wL7Yt8CeNyHyUpo5LEKC4F8GQiD9WbiAGIy7BK/tgQMtYUhghgdXdia1KeAhC753q+xPa1ytWLld
d+ft6QAvIecyWYVa9r9ePE7RDuIxCIY4ujcSnGZ3yc+0gT55dJcTk/yQ8Nkd2uO0puLZ+RlYRjwD
HbiKSe5ViOaBQK7t7UBDx3SY2YnKq2woWyu/Z3sagc/CTputBDkiuNXzWtjMRWQAhTFTCCM3Ms4i
87lbYiyxx4hzS8XCqR7jnAUFEWr9+Q7LGiZC4pd/yhilo+4mEYEiGqiN23EUGeJqE8O6r4kO2Rjs
8RV1hOHW2NVe+JPQ1GPJizTcnyAWADxHUIiXVLWM1uG3IAXKwvr+DvKJeQ8rC1x5qtehO7YUl8wp
/HlNssY9YsoHaVZlI1P2f2xyjsLhtU+A943KoPa94J1efQ22Q2kBvNYQ+zLXCypb1mOGO3FjtZ0S
qzxGXfitRRI7hmhJSRXMILJhE4J0p/5tKPlcOaVoZI9dcp+N1cAJWt9mJtezcHHM2h+PzbKU96J9
j1UsuiHAaxriu9haNo+GCe0a3QD8VQEvKVWMl34O0vE3y4/s+/mzClwVvH3f5UPn5bZn1JESMCIe
XE+SA2lEYhflw5/pik6XZs19t8FSApRTNyihS9kqLIkyVfgnleEwqosk9Ek4u9NRg3/KALKARel1
HTV2WrCDv5ONbecon4Yz+bK9aGHFApAQVx9YViEudaOq1QfNKCcgoDLg3FQAx133i5Iv7EmNwurV
NFgIcUdh5QyMuqrRUIQt9yKBzhRabkxwb9ZC/gLguM45ozvYdvBLi10hCvwsNVg2mxIGw/9kDCq9
BGJbhFfQy6kwJgkKwYmSyvpMljOolBFi9uOneQrTccpmsOd1rxdZxj4cpM3ysAAHLv4zsrLdYmx6
4pxce4lzMdZaSViCT4KbCxwErEXUvyy8ZLjCD1Nu+D3ndYlN/SpRemYJCUgGoxLMZTnzmIb3wWeg
ZFRoSSdT8neZySwwAViEA4SCPROwI0R1eINUL6POstQoVt5bgSjzQn1ubw11Un/t1eK5jp5dLLcH
FPTCZMn/zvliKBOcntf8cOGXWoSW/1ZvIe6noHeFZKZgyB4GF2piyELQQ9GAN3EfkrcQhbfklJWE
UcG34m/lDZE6xUn21tzz3u2QtWPBVGVqWWcCxcenbHFzkuwx3FqSh63gQmZLrP+uH+WhqPnkqYcA
X1/lTu4ZpLpX6R3ibeiui3L7QEePvt9ePeSONrDkiAGxWYRfkrdc2b6yGmzYqbZotVbooJPZqygW
ohc8dZKIND/tR6xoIwc2UsOaGGSoPDF9dS8yTTxv7eHyag43pI2MlledljZr49zrmMEPdEsb692i
RsoiL5ye5fWdh6TqmO9RUX11DzzLsC16fDGNqBJn+K1Zfp8UDHQK/vTdeOya++OBTIUkCxS6jgpy
zqjsAE5gb/rssW/JU0OTH2nJO2oFc7b2TSqADwrpz+jSb7CF5uxSFLQuzLOs9VT4/YxJyZ0uItMJ
yeMoJhbhoCg1/1LFXFrSu7YcwmSh0fTzeDoVsum4SZnKSeKf7pPTonUpIcshr7FWc9/uHKZAYa87
xOgRrlvKsr38ckD16kbsHivy5vnnWMBjvqdxVZRAeHG3sJQGTkeV8tobmlqygA6+f/sf+mbPAfi2
1DDGPoFJ0aXfSbvyIvLJLyHhNaY0fT5pBh1o5iwPYicYot8wv/BQByUwLv2hgf63cX8PIJCP7Tkh
69xoViM9ttql+NxXqk3FRB1f/YVuzthbZBbKvSotH53NmpmdtIR1Xh5SICTfqpaEZdgZ+Gqa61+H
2eWtZi52QEU5hMCzKh7HUsoMBqO+euSL8a1NYWGP5P0R/NXlENeUytZMZxTc0g+XbAoW5SahB+Lr
0Hg7H/oNAFKLmnQe93zV0f9/ZYwjLY+eQreXiFb0FfMYWcOw/NTdJomw8cVSPu3LuToRIRvwxocN
y4d02Ttk98lkqvujoQYL4qPv/Zp9bXNuM62WHy+U8UxjBRhwauhTCN4VRcjmOSiAw16j5IXcQ1xN
d3MiI/zlGnIWtgTZFEH+g8wAgN/8EmuuyjzbO9uBs3Re6nuZyO8fir34tAvkbYZcDlO3lxvEWFmG
BwZMCiD7yrNvoDtO3J18Kr0HMNl4PXCBmugJkq8i3t5zK3HSDG9xIwnXGPw+bfLLsiCG2QrpxAro
lzNYeVy7cF+x4sE4UWgdP5YESV563wUTZlkbeTgLDG25v7x1nHnrra8bE4ucES+szdo9ESYMw2JL
OF362i6Dew4rXG5fuqQqDJ1R3Aap4CHRh/dEhoZ91qrSDpgpUA1Gf31RtmZweto1oUAVEEP4C+y/
0uatpPktOPduoEop8HbelaEB5MjhOBRKxKdWVX7R3vNVjf98CmdUNxkI70wuXSOJfB8bdMSfofkX
DQKmO+gI/aT1l3WQ9/VJWfj9+7Yq3A/j6GyNvgwUuwTaRlyaVkyssETMIrV4c+Y9KVO3nwAC3lIu
VzQjkaf0eIsiniBfoadbF+zr6tFPSMSTJc1wjkCrng2vmUT4Roc9+n7zdj4tczSjuOLLI6VbNxhd
4iletcgODK4J3sG/ZR9GAG/1gShYW4QW2Y0foRG33mgXMvsJnuPNLRaDp9596QKX5jRyGneNnQBl
qGou0pzgiSxQMJN4uXd1Tzi+AgrQaK5KV9HOynjeYFaP+Hf/ZGlvyprxSQ2joIxv4bLgis641lSe
99hopAbKpqkLygBe674lCNvW3cS5Ch2yfNdMNjxQGr9Hg7dhp/5SAGCD19xs4kQ3yxAPvO8WzPoj
5ERN99XIKvqFUkOyndETiuSrpjATibJLePB7k5Pt+k5lkCCYLGVE0wyjUsXbUVvTjE/SDTKxYQRk
WqPAf0KEvIJ2rY8u6dNy+thQP8BaUZTMnKiOE7I5sRdKHF5CfS5wmG8DmRoG/I/P/qp8hbUkugIF
+KJq4CSaGgcpMnOSHZoZobPmyjDUP0v2nJosPoE6KaSKw/909AMv6P2qRSkmT3jHkss9JN+opwNF
QJpqLW8h7SknmkW11TyKbSSWofDvER7hOq/BbeYe393d6QH7k+LDS/2urOvKFxVZAc0wuxR6l36r
NlT9RSmLU0jja93w6TdnEYME5ZMFJH+rEuWmeqUlEQ2c/x45kF3xX+EZh/W4ytz4II9LrAR3LQ01
eGUeJp8d38D34POs2+QLwxUFEmwGC3EZEmm5tGhuOgvu2AqZsgkIIece+OWFYcO8CbADrBSy7rXx
ToxzFMTF8WXuu1JFEQXgDbusnyRjAGs/Dr9kgnPQEizEOZJaQ6LfBL7TyzC9ESaDXoRr4ccNW6FB
IzZjvodc7u6N1pww+m/6Q/wVuvoLqUlYzY22H7r+jDiNELJdxP4XUlP2eAnnTG4HUHKUod5APkok
1Nl4zwIFoRwmoZujH5P4oW/mvdVYgsdw4RK7c3xtmqNLYJlM5j0MEE0Lsmr68S1Oebd8YC57RvYm
+0b6X08oCDF3kHYBN4XQVbM2UXDlgqZShUoP8UtzGMFLe8z/Z2cupAmc7RAP04Or04OUB1aHGAkS
KAhXklOXRpQT0TXmxO3kClb2SHtsgoxq8WayNi0p3YnNHdzpKt2SEpxvfy/a+C5KCYSo8hkB/vAl
3k97gshD3T+hqAJ+rSmvLPr1v05JxtZn8qyAtkOq+gsk07NfvNsEmpGErF02ayz7gdmjwYtvNK/9
Ly2jmKSMbxNn27AVK/CGj9jqAyxvshAgeYgNHghXXybU5/P94VScynPzCnuY3tJSNzkEC7xWl+G3
RpIo4D9xpyQmo11CSO6009eVokUeRY1BJ6sjiqyKOC2MS5r2ePDrtdu4KjC+mqCr5vmnb+V3Zf9n
KwOq9rVDJ6TmDrL+gBAX0RXpIYi0/cVNSpfODb4zsAA3AAeDS2ZXSfSXNbHFXkVnAzeJSi7rpeJf
MxZ7HxrAjufHrnT5jMTSu8/xJR/ZhGKwC0Q1s3jGmO+liD8UjMj3JOfqRrIBT+EOmVH9c6QU2uEE
yY9jarLJQ26eKOwZ05TcFm9Nvgv6MmzpCgQWb0p6t3aSwEt5pq15+wZ7GLyCiNLt4ZuxBivVvrkb
Bvc5wCIOIhMKEOR/E7o12E3hBnDQ/Y+uLw7B9araYsD3nkLkXyKsjcKmWetbywMC+s98Gubg7cXa
wIrdXdqa0g6EBJwbgN4yxXACIyBSQ930fx3F9s0XuQehnoLVc7mgF/QWKApk0kpoT510RlYm1aBt
Ewc46J2ni85c0fcgWUL60yuDlsRlPyubsdaEcp//4T6zo4KQOb3tjf0B0Euk9j7GWHmp2MzF9IZO
LCjEW/0MBU3YPctU1xUmf1Y1AvFeOcSlLYkYk+aSyCWiiZBqHUGti1YUQVkoyOPF6GpuZ2okRZW3
DQLiXxIuzQgMgLwpoVtmqn7/9ZIuJRZAYveUmlJLwIBYdEJQ1Ql3tgiOiiDavRniEaoO4/P3apGP
orf5lSKotOhkFnDZDG0HnACX4DPj9HtOOUvWTFTqQWPIC3nweU2fVEsRIwrydIpd77Ci0p37iN2G
CCV5UHRCAU3uX/N69l040kfRN0vdCE0kNOS/qWKPQIWVVyMzLiRogXEuIbI5oUv8tXNroAvhk0Ff
UNhaRr0M/akMFfWiH8g1e34u1eNgeCDVR/jMqHrdotu2VDx0FFgHDx9orBxpP1WWPY2Qgwmvh+RK
IzhywxB4n989iQRuCDCisWhRjvful+QEWCG1GDy5VjX6rYUD8xJjcmj3iWcGXhE70OMC6pZdqwKX
S7cmcTFXtp9N7myMx/TqavdBvmMZLVNUtiC+z1Y0E/qSp6lqxA3W8l9areFyhzC4+z7iOY7XGgsV
Gy87+XJLcf90WFUFFJ7T78ssQZJh6UpFGJ0k0ZYLBXD+MmVz53k5cGNyb9cmg4v4U4BtE5XeU+aq
QP+UtI+XL5fCF/ocgns4FlvxjopuwBw+pJT4iBdZazG2k5SAgrga5r6OJZuogdcYQg3nnVuvrnV7
uj5w9hhbgtHbmbqC9lGmnrCMt0y4ORBvB83H0HoEYcT4ayDeKZP1uvC+ynEdqA1N1eFTYU661fal
b4DrWKqjmZMD/e2Fss4TalkLUyuEe0YHufG3kKjdWvdV5ZxjR/2xPXNAbItJmyIvfGgQxJtlcGH5
YgEMCKebSZG+7dYJryuqI2fbp7bqVhkB91NyUjnzLhhgv/k2DHmyPy6efFmrJv2EmpRRGuJOLosA
9dHgFit+yFwolxjUlOnK2ybhAHbr/JtBx/Ae8GIW9LDPbYF4djs2J4CDO9O6szGCGkDcYxpVMcFp
Nix/TJvRVkCXVy4wBaiZ9cnGi+UoytkMzw3cFFrVyKpp5phnwpaImGb7ffzYmaNKIs7CzzJWdd58
NLQEgApOMKi4DNNV+5BJi2lcG6Xly3+QP1WIAMqGwxIa9EbQlsnzjq4db2yySNDtLuAd7vgNlOqH
2It5hFm2MfI2QJhXIci/pQmp6OQW0k+Tr7FGZGp3f8KzF4rIuSj3blDeP+yOtwYb6+ETVf0Xhq74
jLNA4BxZftOpfMOAJeOfmTPFSiRQGG3yeAeWhm+Hs9cIbxHzjsQAN0CgppqV4I8r1TvGn6hlx2e0
wOGoHkxaLuyKDAeZYXpew9S0FEeJBs6P1tMRpjSDwiBdJ6XaYd7/FyMiZ/mxcbzQJsq1rr97it0t
7aTBN9fqkYZF4OkdXryM9xgAUmysVeYdZsM835XGSqI8oaGffFi//HmtUduSWRfarJL5Djt7fiCN
icm/DltXXg1UYdwivmUFgHJYdmMEzKx2Qi1d0fL2ctmYE4oP6RplpmVyI3+dvpw9l50CJo2NY8Jp
vN+XZDxScZJrSUaruwcCFLEwZC8xslrvydRo1E20T7uukyt5Gqq/ZAmqqxqHKPAEpwK+DB6o04Bp
Nf++2/xCLAuvjajGw7DzCYOo2s5Bw4etUwomgZVU4ImZR3m+slSOOiTgG5Vp1O1GhrexszrTTUOZ
W8zRcrniWR9N5tA+7jn1oSMllgXrZgmG6wrq+K0mzn8aR0gla8ZzM+twD9aQ1yGDcRoNHe05XvMb
+NWBMUSX9pa3x4F9Fp6opxeahhr1ZlXT484/vv6sJP35Q6HYs9WzjW+fsTcMy+bEghjjMJj2WxqI
d2GbV+fikNpmkqkNnsFjvvSAYuAbyt7i5zPn4mAAwI0vzr/KI7vzxf8BHp7KZf/jZFHs2Zq1jnUs
evIuYvU5bH0Jb3raaRxQC7gCaz6fyc6ja9cJ9WBNOFTZYz6QKLTQs7BjubI73Zf79WHhhx0gC36s
Ybo7pEtvF0H7ZnuZPpeM9v1KiI0f3iMPVffyHetgwyHzesMCF8stl9+PGNaBG+8HCEGTY5l8m774
5l3zfXFWvp+SFK6S6wHQibmiyk8b1p4cKtGnncF/eWmSYE6ueDhT1F8bhRSPVZZ6dp6Sq/vNLfM/
MloFMT/gyY6tdUxk8lMG2I0jyBDTo57mSDAIOqM1w6rmPi4gqQem3Jb4mXnucfZG0YHUkXdFco9G
ZJxe09M+BszQxA8wshR11NED08jMu8EuktGIiBqjRoFbSfREdwisqmDEDTg59xYrKxjSn3hnpUff
bMWk0G6iwjuhJJPj/dRfWW4pybxbDH/wfTynHpr2Gp5mVDTqdYec3Un7jryFWyNNH/7Sn4lagSbq
/GI4nAKpgpQknwxrhS4HHwFipqT9Js17HEjykglBcWkzEonlNq48XHbeEjycGuZ/SAiTrAPCGebX
u/RqzkmEH7/0KkKAsLdDGWC2qHhMNbtLtxKcWhhxooVzyGPZlla0nMCcSK+aTvH2wCYB/XtFCVuu
z5UE+kBDM46k8G+/gBLbSDCVXI7uwLYs+fcEhWzfEEpVZG8D/Q7swX1i9DwH3T1xa1QtP0ipa+6Z
a6vdTgYggova8n+V5vTlynkJ5LmtoMx95uYJ9MQzb83O22TWEpmYWXIgnLIroe0n1JPtLr0Pdbqq
SobGRc8QGQCCaRLc0JGv80dtBuS59gb7wcGK/kRB/PTh/8Ak+tFkkE/XSQa/KHaClaW+THDJaPnw
3RFueuQ3IMlKRNKsh69IHVQQyw0/iejLJGohrJvXnmlCz3JTIy6L1rKKDCTpU1/l5FpRUQlioLDv
Z6VCCi0meN/72NwZuPPbulmfb/WSQAvdpoZVDGHccg+FRUc5vzRq5PLOmVCNQnt9el6ejekTMmwT
hwz1NfHLON2UhtRMnJPg0GDudQ8DqJYoi72iTENJ9QW2I9x6hdrWV0vZJyqICTxos27R9c5U90B+
mUrfZQCposkjmqjoBv5rWMW9A3q6DVXDMB5Rx19lEdyOcsePPREVMt+U2+lk4EhVFolRjyDaoRQB
/LpRUQUtZcY0/Jqy/cjgivyhDXF8Thcsc4S8fdgOPNEawZJQpjPFEyw41WwfNPz2BVHZxAM1frqA
z+3tZtlAztzts3vzClAq8tvBkg6g38nGBYxfBWQfOvt3+ir1y6P9jAp+jdTIeBr1u4YdtM7ovZYv
3ib6SlxJnRHHMLQvaNVpY9Oex7XWhA6rBDxK9uFnl3JDZuir/qunP9XCMU0d4DPNzi/HFOJBX/y/
m4aqLu6hNsZcQxjKGrJNktxLe2RsEIlPLWgHUkiMYOTj7ifLR7wxQQ+feRkG24lB3K50jzak+PPp
as4hTrjXF1nqEFmopCVrefz1LtTFUY/5to55disfEwEYYHcZvRATCzVLmzem3JDbbWaLBYZlbZY2
RUKpzY61/Pa6W/IZ0vu1/OhmrRJuMNnxnN7d+SD2y1wUZ91WSAjC9E46wfulgWcIHM8JDzs2nGJl
tIsuuJ4SEEj9gWQhQpo64t9ynmlrp4C8pewkSWEMfNWCSXTJaVsaTy/Gy/k4HsjO+2+6eozzCbOw
875wjEBFInsolsBeejEh3ZjOhtmSHMACqLjJKOMI11uC9c8XxWpI9NWFpYYTKdsIW7B3DzeHRB55
33HtCSBycemzFdf7DtVK2aNc8XzFXQ0s7Ohmm0rgxO9YOBMlBcgibkucnj5lYtbpF0jjBk785bEH
RlvtuayP/BfhyyQcOaNP/ggJqoyViB3TRx5Nspd5KnWCt2iaW6bdAE4m2UqZBK41/WSN3z7Vlqds
z767ZR5PFxt5RzZvWsyUL2g6oMQLguRh3J17blfShRq9LBISm5BUP2lT5XkwUArwO7HFYNksuNof
+w04302vvQgqufQ1ujBv2L+SCl7p4kVrv7iJs/6LmlrYLWIx6q6uqUTb18VesspN7xdlV8IZ+dPl
WuPXtkb6Vo7w+XQq7X+a9qQWOnq1s6++3lmaydfAXz8uxrBe8vysQbunyjGIeoyOWkeLben16Uxz
0ZIficVddDehICXiMk0iseRXPLMAlTlHCIFhinzfvztpbTi9nXcKUsYb2fTB5cax+FPnYtlR8XCK
ZvzxL7Zu/285nDwyj6r3ieZ3bEcK0pK5wyo9jJ14qYf34Ksi45hBQtcsD4bOY/y2rKKjTXxGzLtZ
qMe+XTLDYz7cDxApKJmRh/O9jaz/KNxvdo9tFUDVddLrO+F+gFfPMTnx6XVX+HcYeA4RQKxP2mD7
7a7F6lF59pQ2PeNwnICZS418SdkIHSokcmTkQvPf4yzmzr7+h/1rSbes1xM3GdUdIfoa2L+6sbDe
rIqSjz1LCBy9BrwhMBER4ma2AHVy7gUuF2Hj3r1aoauzIK6EYhMJXnLFLz8zBcuxnHSqH+Vb4mRZ
wwqCMTTWSW5AaQPaAxt3v6fSmkd8vOhvCAHYRnQYBq7AlZD8S+saUk2YEs1E2QLV/U2M8bi3hjYK
yVOWsV05MWNxmlJxFGLZmn/ar3mEWb2xK4wL2PX0AxK0vSLMnd3c3AUQHKZ/r4Wi79ViFcXfJWG/
QkZU42/2joC3G+X2zjzkn9z1+RR8qJ9epY2ea/N+G6yp9iNNMrNQWHoxnCwP4proEt0ZckaFmBnt
tU17+TwKvhWPDeJIA9ReeaJftgCu31QabEDR/VWKZFDvpCkqAB2vd7d7JwC4h7/28El12jRfBtSq
l4a1MHCTBff3ODmpRiIvWO4vUI4Df5kvkR5DtpNP48TSZxwcq7YBtgIb+aWij3xUqTi6KZUOWJVq
SRRcwTWOAAQkPF6dsSmKBzVTK0hBQ6r17LGVH8CQ+QyFjWyD91UsF119M5Sw9W98eyhI/oLsywu3
9DX2K0dnE2h/f7+YLAfGM5pE4Ga3BxM7hbcSP+2y54hAaaexbanXqPLP1nQgeccZJhU5xIqDFhTu
Im0khxKUy9ixcwdVbS58OhPNZwCM27rNhtM+hDy4slJ5Pb2EUEl7rQTCIJXNb58b5eUBCaMv+SVe
CvTHb+H8OHISl7TwO/fKAt+TMMWQItV5y6jaraERwzE4FYEC6SlVUqvttDHZmQP1MzcaF9dabV1A
B6GEBxtbOwjo50pbnWMVNtjcuOjasF73NA4MyVXlU94gTS+BxF+qKIHGpXyZhd3idyKqAkGMk9XV
RHkf9nc57x4QrGVEDGxal9vYEeWI8SX+tBChngW32Y/pUV5HhvZH4U10xzwaHcBhioXhGT5a4F0k
Un0IY/ONI+c3oFAo0QZvpvIvMlNdaQ62boJsmrYOqN0G1UVZ45a0MQLqyLX0U2WvbbvhkbXMMbSZ
hAYiuBXdjeLcLUqgumE2C1PywEeLcHOkTi+fa4tjoVlja//fL+yNYjjKU/oSAydcZaQjM+GLbuqt
JUdgLU2EBok0M+WyXGrsFOAx9iS+EmeAMhqv+Cz3elzD7iKs1nscfh3WdiFRwinoYoWn2frkUbVT
e01ENn+YU9M+NxVhYBiD47SxbwszfdsIHvDndo9bo3IEra4F9mPBJ86pOl7UyoNQJNXqmiKgkM/V
g3WzUKOa7/FMrktCXeoWgBUSAvN6qP2w2X7tODAZblSUV9mIlv/0gwdM8Q6n9nykpA+OVU/wMjT9
v5sC4+wNzuILTRjDKnUxxB8sa7waCSY3q7YR7hCEjHOYzr34A72MTFFx+p9ZmBunwEdYoYzV4tTl
/8OrHkjYlrQEIfddhY+3D5v7J3Rcib5zl8KRtxyK7HgLoauwfOswQNGR8Bbciw6KeNcrhbfPIDvU
1TjQJvMr6N3akXwSTnSXIaGnytqD/QOr9XdRUbvNsdsvCKIjEz/3tLlwtX1m3qMN0o/t4s/2BotZ
9UhNGDmxuDy84lm9HEGP6Q94b0zEGGt+98ZuTbLLFTSre+a6Gr2UdJfLd93cEMrdU3PwjREckEo7
dxbcQ5am+2XpllteF3nC1XMrN3PuGKZ2IrtiHXSvN9nE0/GEOVd6YWYXVM0ckv/Q6SPTc8eljOeT
S83x5vm3Ly81S27vxNgD3Br38/7hmO1v74nYX3SzRsOHEY7R/Xty5I8XIwldh8ckAHeLA4FKS4i9
m9EUW+G31RG1oEPI39+3Yj3fYpJMFGeOB3/rj+jiLsVkxLEe2KKB1czZCxrnCAo6MO/GnR7hD5Ru
4lctHQdeqAUO8uuziD9zgwd+wp9xNFakbb81b8uwBUmOgehxEGgiIz7o2yhI/0YI7gI2uwpdKvj+
/4c2I8+CUEaisaQTegsjrQr4TLqM4spmpH6jsKMsyyB14mG3vTCyCsCUaM2h6WAsLjy8cHt2rH1E
i52DYm+lbb7Ujc3Zxe6WeF0IWwE90EKbn6n4McmddICXawhrFQ9OwPFLAKZ7FY48pomtEifC5Nwq
pLNauN8Y/Qhm9ULpRTdYCXWs/wd+vhWWZYHGXwMoFsvX5kG7nD2dvkr4czqzcqprNGU/+ZdXze9d
hU91RZqnTwdYYZAweqDCeYdnQwYE7JRz9JqAEzWdHGKayhD4wqr+RiJ5z25eDHoQ6BiWOZ5k4gJ8
ScnXNMZNVdAG0GSRgzB6kHo+wdkTS9DH5rcjH/Ljl90LldxbAUiYwv7/2SrgFrQyjdPA7lsOWcb4
N+G8wFPLEOIR/9IBorTSlNRbQCnfF3baVuVxhQl/5hQxMYlGENnnXVB41p+5CPudeVd27IQF+9QD
wBebSItWWt/YKNHcd0WZksYNYiFTA/6vOdow2Uuu+VTs6+XQjkBFg9aFl9TMqs0UfGFjz60M7hOR
pi9WNHJZslOVh6Ym6J1XXpE+ZnD3sd1x+Vx4bPmu6Jq1LvAmZCLwMMWp4GDcha+xfr+/GWUeC0Xl
ZTBVay5fUJtfBK460jEvKE4ij/eg760ECTjOde0NY855une7gLK0ojUn+TJp9u5/zTlwrBqd9KMG
JX1bPWo35ld6YKlqKCPuRAUwdNhv7JLSJ+A4CH5iV/6dftl2625WyiyvFQkPvmrUHifEEmkR+IQm
XqnnR6UO2Oo9kj8aPOEU5aox5ZJX5/Yw16cDiPwuIU6mwAbvDz9B1zFwvcPqrWKIDn/Ef16yZkZL
ub9KquOK3l2OMhNa7mlQp5woGoTDAv/WSvewny854BjD5Lwy9Xj+B6dRSaVeFWvcWxMiW4x+eunN
sQL1Hf8vKGArQen9/giPGlFYSyEny/9i8u57+4QcBCj5/5yFAFeNy6LuqkTQL28VFN1w3wDdG7lK
r9+cmsueuTNxuOJfKIJZnJTNTdOR3yUv5f9jHslVCkLXOrcF+qnr9puk7+8m69jdXY5aHOPk1OLC
jfUxC6clDrEiu+gSunwrt2QodmEvOZ/Os5Hh0LFZF5v8wh7igmro7VtcnDLzDpeVy9BJ0gl2KvTb
T50oNbSuSNN1WyO+5xlrz8mtMJNzHNVLb07Ip9LVvb/nJkX6lj+hPP4kzihYnHjlTCpDVvzU409U
+eF0mvj6OlXiMb9Qe8rWdKrOY9EbmC/W8oIREiFGur/fWrzJOV1wc/036DhVshpTRf4JSorR3H02
jm8+0Sk4RvGc6AcIXZgHrYmJ+401O/DwiJxmQs+N6CTxljLBFyTVHqG8EGv7IMkn6nLfnvqFbhxq
fyx11qlje9seHHOsMsFGXaGKNuJmkhiJMjHXIFUYWXL/08Zlfk9gF6l9jX4Giy+st4vviz/ZOuAt
GWsiKRIHFzsR49VGCJp73RL3fS3Rr4/vlMgYUO3pS8H4sqKcMoip6TQEU2UpeKoO6B+KsNimXxcO
qIHMCjsJBVy77djo/1y4I4TUjHecS9UFBPblgj9KY9kVGTKhNGSjgk3X+MNql07s6JXzOzhUaCvx
VWG/0nQVsi6ifMqlWoj+sYzDYd8vwrzu3CrqGHePOv7359/tceeMuRylqFXdPFXWSuHOwC5KZ2kP
TnsQP+w8MN0/vT220DXn+Uyz9H1gvrkvotgD2evdLyXdnqCQdumUCvS78FvJv44DlTvg0C/tdkOU
bDY2BpQnFZEr2+tXWtcbhd6L5I9Dx5yBGxptzMZv2+3JbyF4O9T61sK5ncxragM/g9VFcrk77CrC
TnehQg95AgSVGjEZTcWkMw0BGLWJwRLzdRZJbejGZ87NvE2bP0nlstrtQhiO2AUaFAffLj/rBaJ2
NSsmB8kSEc7qaztvO00BM7uMMtTwu+WMQm48XVeyYzqZgn2PJ6FGQ4cC7HyMxNa1zYuyC8Jr6NfI
HjAnWvSCHwE7rkHCee1iIkt5s8N3oKwPOQj72tOcgPRbv+suJCY9aGAPZBeZ+w85qu1PFzi7ZoYp
k1RlyIak8pDR5HSHLKcC+H0DajMVlU2poCDgK+NrG/fgagmB4f1cQkV7QeJFeL9mtWddwApeROO9
O12ydDmaoCbLVUqpBPFX0DZyeTz9+DHBOxw8z9cgHVXwCzvF+S4Znon2GknhjdY0aUzNPx4ZhqJH
7rLl3+W9juDgQCkUerzn7qW3bnFfHBS6MX/dk/vfxC5wXmNKGs5/Fdphv2v1JvyiGVgyzGPYgV9o
OJJTC57XFHhDPBtw6vcUCiumZ0TPsLOW/sE4yKyjdSOEJF/K/ogZtNTjaYugX5y3cLOO/LSg876U
lzgy3Gczr4kxLG9WLi02cf1igDov0GTmG8w/zqBE5+ngBwtTv6jkvAuZJ+R7CC5zQU1FlLyjdDhW
pNOVFyL8rDAaAROPlPw8qIXewvwFpcq+LRPe88UuVFBT8WUXGfq8eMPu6R9Fb6bDZ5uNKYoKJLLN
zCGs7DuW5OWLUJ5Q1lB53sSPl3zrpYrsm/UtbQR+nJgS2rw+nx8SadLWC8IAHHlF1B3e6nbJSaPQ
ZqEtlwH+cXxOaFo9JKIFMYntRE9JBRM6B+IgYIXLPr8bjAWqcXNyvsopO+6NJwtEPKc56mIssEPE
ARvsOk4uzfCDjGLTSOuWUOeCVXFwCtYHBXGbtBc89gXFYM4pb70C6Ldblbc7yloWSppttNK7OV2A
9koSDUF24r2c5pPypmZ3xVUNr336ohwbAmShhdYhLUfxcpnu+QIVRLaX6DE0eWWgGIEzVmIHN0P1
QsiQ6hD9jneoS2VhNMp7NGBIDWy7La8dLsPvPPZ6Uy1DwQUEII9kCGnmRBKxB5XepOm/s4kNh0Yl
nCxrM8XUikoyMo8TRRwyy6fRHpfODdWP29QHN/P8t44lLJybhqs2gmh+yVTJ7KxmZb2QbrtuRmEr
XQjXS4DcemCd9lTyVikr5HGwVReQJgxU244d4BTT1JqW1zgiRUdFa06EchuytCoF0CEHxi5mmjqK
9cFGC13F4f6dL48vyvA06I6oSSeUg62nEqK9zf2QevGT6pYElrk9Eu0m7XOvcdHJGGcDPRo9q73c
nzsmLyzOAmfNja9SSYFe/7HslDF1mRcdXsAGjSdPniF/G9dj5auqANBCfv/dcRVQzNbgrVaK1YU/
EP1bluZXLW1yQJm82DknuwHEPANKZXXFOv79FwAerx4DO4hgQnjK8JAT8Z+PSigLEvTgAg8PQ7DF
OuP6gqBp24CcKEODmJ73ERo+oLqRoS0+NGRoK4FmustBQmmmkgYPz2kgqNrL/09Wlw+UHEsfXRmR
KlPSusczF9rvu+BrcVb9Ck8a1cp+94NaE9V+SQynU7ya4u61Iskbq3ROBwflMqyGe8t+hXUHb9jn
il3X+BgEhtlBwfXfBNS9CJKQcUBuEc0cCCHmkkRPQXI90mlETRcMddJ77O7/vjmD2zrU68xmIemz
KCDCiDSSH6nwW5EIedHxvX9myGuAAa7HrJFO/j0aiVZin+yQsXQ66bzcr5sfGtSCLHXPKMBt9Fdq
HwmqEbASzhfnVNgBPu2EjkeO5wVrcLj7IBZ8Ew6nuyyJghkFjmoM7fx9Yg6vEAfa9pVQP/xhFsbV
nEwBkUiurAErrqVEyIOhzZxcB69ZAD2xjDnm2o+O+C/bgTO4UkqVlW7toOTv+MzO3gtWRazO6Kl1
zft7qbDIipHtSvap+4/SYKijq5o4GqOPsu0Y6kRGlp1L94n+/IdcW/f8xhNu7nbBwALHMqOZkP4X
bZl/HUj1c34XjXKYcB39SRGnVdfD0RgQhqJx7VoNXf4GeCCQPeLm4eSWIr5TBs0dJmj+ke85uFuV
kG+xVnjijbIn1nt+2UPThZIQpoEAbNfzKvDUA73rrHFs20Hkc0uypHnySxXzWK5AXb7XkbGsaiJU
0g5JLOHDEX8qJfG6CQHOntXlKRoKV6uTufh3QlnNaCvWKFQGTUHMF77ahE4f1Me5DfvYAg0hzF4n
tUUNHSZNJ+wZY470trAxvS5wsT0WvzSo2dE/RiKX+3sWoHFld57Z62d/82N4i7oW3jqmCeudeTSC
bsnaZj+E1hqm/j09104LOe45M3EswYhXS8JpVDRQ+KAThGy7W9u5AhPPjDKvkolBZR4RX6AdAF6U
8Nz6zJZlFfZfGW6ue/DomKa3vVUP/B/38l/kDQnM4YMGHBuTdapgKuxaMQSs1yp0QsxV4tD7tUft
PuL/dH3wIuoJRMchceFFqIx8wGtHOEpWBBUtAMruJS6sIfTKcZYnE4ofvP3FNdPf5eTPDHCk1peg
rnudz3pJxrqeYKtI9JX4BVu2zJ6xq/9+PWcdAbjEH0uiitjQrl6Cu1F8cW7UiHUz+MKM6SJZzHJ2
UiT3OKHogRP6ePQHUFre0iWLWDEXdH3+cdTe1s4+oUW6AStyVZOdDvKfTyZXEGkc7+vt84ZLQ2//
VijujiP7iYbZJQ6PfbhyytCRRynP/XL2r81kz0RgF//g+ngTTEsGMtjkQDWuwKHG1aqbh7Apmqxt
aJW1wJq/H0aHQdXvqF876zlvE3ZtAhH9iLDaugh1bX6oQ9eLm8k362Ez4tXjrhfHTjUbyIA2v+EW
TaZnS+WuLqKA8iESvrHxdGmJNwQxrQEq/5YMAZCyV+Pp4seARiOtwFNo0HYne9TDdSNh+RJhfKCl
OfgcKuWtsdfTdGgObOexVBrZl4WG4zofb0Jz2MhXzMjrP56IBSjw/t+ipuHOat5zTh8tQRnKTVI2
JDlnC6w6cYEyt5VluKb66rAEF2yp3h61womHujd5mbTfHopBffM1JXC13epplQltyDLpLJm+SEpd
uO2Vu5F5TpiPBGaTXybM4Xbue+PVsXT/w9aDCf+5a+2wT+pyUeWqwWrjWWjv0W8uYqMkhrJTXuwD
ZLzw9Ptsv4o/7uXwhZrg/WeGzvAdrm/ETfZWS+xRaQYvcqr/242zH8ZzCh59RtqG3HidZKaRjxa/
Wp1W7JGrIft4wKnDddvANsqhCBln3SsykeEFQt54ot1dACZihZeKVjLGv612OI2US8arORxHY/Ic
Jo25rTO9UOjdXMGg9YCU1mWVyIsQglDuOkwZKm+TCjCTqtN4GhPcgt9lp2wrniFKLt+W5FY1xF4+
JWJN8u3nmIdJFzCs8BMwQABQYtP57zxsOon0rnHR12jgZaKEso/MvyTES/sKNo3+KwplFj8ec120
HXLtdzihzThBETBLqI7K3g5a1oHyRLWo1pcQQq5i4IDkhqJDlS05aFQzpUkO9h1ToWyrJ5QQC8s6
FQM4tZxUsznzZoVm5EnrI+jcMKHbIrt7+2Qcj2+Ukh1AJTvUMvXk04xnxHwQ5JvEGqLgAvopb5Ks
5XuzeP/GqhZXjIo+Kcp/mKfS7/1zsM8HlHi3OUWQ5PlM+ywytF4Jm716NK16PmBKlVoZOX6ivsia
Cgy2/GQXyT32cJc87B/MTEmS0YI8Gp3ccPPTJDYiVciaW/BZKar7YJk2/WH9un5eo7kGXnDbnpz+
qCTD61T7niIOsKB25W+KzY1ScTO2j3R+tQmzQ1mqdA9jUJoJ9lexCoYMVyI6mJer4yVctflaCQdn
edvg8YVCCT+kRUOXXpFez5vqGeQrNdwNZQipuGwnGZfX8L/tuwV/i72W2KFc0GtQ0aFllJcmjquR
VA1CXZHNU42Yua6bqrloM4UMlRKtZyrlKDJ3NaScHY1WZQ1OsvFt7gEB13S2NvWWt1l7c9Hnn5R4
hVEGbfnWBkOmAtDwkvCg/yeS1YVMCTXKIcikSATn0TOSW22CIV4NbK9pBXqS3zUPG156xTdclBC0
z3EPlOgs/yCCfJ57UqkhzLiRMpekvKz7vUX/xe6luhMDuExJjpsUkdFlICJ7uFDoZ55gcjx+kVUt
4ZC4bCz9bWk2uLEZoU6wfsiBFDvVb+YZyUUeJKmWW3XNWZpq2MMh9a61d3yMlmnUStYbVa3i84c0
DSwwg6szkeGzevQzit7IQaIBNH7MeN2W+mfVqXUpWugnApzCjt3kZ8SIMh5B8t86emE0efXSCKAK
KTZzyzPqwdH/7U3mIakV1MQmccGiRd6Nf0FCdX2Mdor99z++bp6b1IHEFL8ivrLOYrA5wXDeaD2W
13qmikQBQWKztZg75uga2cVarB6M5GqlpBioIsmANWBxieAdaQX7vk14G4BgtjJH+Oq05BTqW386
KsQtpXPdOREMeBZBOhzz7zv0mvWzo02WLpspqykvgVqc8Q8ixTAZaBz0XKMOpIN+lXsPw1P5hx1C
AZtgHFBUBdIvl20qmwPoVJM4q+KdTjcmQqZ40pXAnDtNqG9N4Sbadtp88XR4pHo+YQkQPNARWR7v
2SMY0ybi4RKxZX8ae0C8j8YYrPrvWTDqWQymQL0GFVq7rNofNqXlYq6EZQ3E4VqrxIYvcff5HLR+
n+O+C+75A3C3826Mt8GpvqG8z/af7vSNlOOcZuMp8xrX+3r7wIJtrV+3bQB3lOIJwIkvIN3Fg9/X
dqDGICgfIdrdscr/wEh9U9P/d4gOFL03KZFFy8qkxkOnsJlULSriyYsI/uyoxOYjH1M4IwusKkCE
J0EVrltQ2vAvI2vYIvTz9Rn0J0XU3KkB9bnDmOzRuQQm1iMdv4DjPmhBWga8bUsGA/JEDj1q8TSP
nXCr0+eeRhUj2tSvkSHPFA6UcYLyUOFHKgovaumYJa26ad2d0LcaCDTavU2NeJ7UTCPSzn80l+vP
HUwSX07DvWe+7449TNaoAAAPTocMthWqIPNdTOa/PFXXE/uQ1eSMwRmr1GqGXtdrMGXRb7T6YzoT
T63B99UMmIzQ/KY0k5XlxNuZgpSeUs0JFj6zeT1j6WRLSwlUPE2iEjeAJfQw0ytO3LTkAwD9NdQr
1YLT6iSuJ8lp8Uq0Sb5TbciwXb1WXOETi7ix9uqfFvDB52XmLvCb3ynKVKQypeHJQsHCPdw7gxcr
DoFCUxXQQ/2ckBvAKYvXMHSKrqdC11pExlbuDw5begFh0WEeZd0nFIMh15etWZvysZ1dTKWCOrQp
izcuTiUQFVHrsSYeARQmmFLNsozyKZ18fASg/2AsiW0LD2qShJLbuGvInG38MmlTXbD1jCrggTu7
mTd0wxJQ7j7ezC9Ha9gag839oelj6ebIxv/qtdqNB5bl34AI9PsaNOHJYc3SHDT1gagCvibBVh7I
XkG514blwAXerzd/MjnrhsLUjhDD6CHsVqWOOdnVX0JKIWqNExRm45J3a9wJNhP3Pytq2UBpRuhi
/uxLJNA72BFUAzff+L6aEudEcKKRn3P51ALSie6iS0HEDKlRZf9Jc/09rjuzAe+tL4qD+yPSjZuP
ErEWA0GqTT8bcQQcKkX1GOXwavCvkGoV6UqcBg9xkTZVI1HugEZvBT+T2A8b3AuiPaj3hux3blN0
qq3Clgfphly30uD3OZstfBwGoSd4ptEnllADgdMe913VGCATNcPYheg8/p+fwQlWRmGIEjGRO/75
LeTPlYdPTF1Jn2SzwCKas5T+mQxaI1YyEnFLT4B3C2YsX0Jrr4QaJs4uASqnTwu7XjY9eDYyEpi8
S8Og3iMvuTRycqEbqNgURF7MJdLAKXGnJ6CQyNUZzRwZ+x+liR7D3ArLs8Q/Vwmw286cHG5jjKfR
DohB24fHat1j7Sbl4XUJxYUYpAjXj8ROA3Oq3pAvRjzsJcDMxqjXkdFPgDW8rkDKPu68C9/ZqrRB
HU2r0s3in/6WOqZysbzZ15tWb5+u39mbct6NK7XYGQDQytqbeipOlbrcxo/Xa028tB72i6Q6cCBU
oRyFGFw88DhhpAP/TuHtCSj7RPe9lrrluf6PDmQ0aD/wUgOE71cf19y5cXWQIcCdtdGLDtkS9knx
RmREx2/dfgxvFgCFqpPgaC40zga0mCBg/DbQPM5VMEVRrlmRnk7kIEFP1mQQYYAdvKMnFbolGff6
rBRpCDD1VfVRN/1C8OZOroUmEf5JKlKdp1fK2iBx27qSCkGVow58vkXF7YywmuAnHVizNFdqeqG1
5kJRqT4ZcsgoK15yH0N8Fa4Poeq6C7bhd7HAiYlg3YtpdrikzVNq1qUSvee01XS+lLWUgkTTLhAr
chQGYbwLXtr0KDEZ4FgiYaX2MSFhP6pOpAVz/YRbYajRmrE0dj/r36B0IVI6Qua/+LEeRuBxBVZW
ZwuEjSIs3Xw0BTDvMzQ6mpQGmko+B+V7bXIr/fRdX/3w9tNnzYhHnhNX+YPWHQG87jvZf+3V0WYd
Z1p0L/xmz3lBVYms2DGdpRVTNzEvc3lQqw0fuceImBtgrL22AGYlx3pry6CDXNl2g9LEyrPFaXb0
xvF3NBXJYXbZaUH2Cv+J5OJXuwTBxboaFo09J5DjnVnQg/3uRnOBBHgA5K2OZ96KPU+bbesVWLLI
GKWRaSdb/CVyvcYrdmN8lSMoZ/kI19hAA11v20rowrRT3MoyjKbMT+2N9AuoARFhy5NfiVtZ//Cs
7Xpywdy4gUM8PcetZGUJ5alvXbsIOLKogHRjAujemtBj9zjIDDJlUbe+9p+GZYyw15C61b2tsEk6
np1w8iW5UZHCdSka1d7l1VAZ0Sqfvx5cC5SrOK+XxU4t6XY627RJXDCR1RegOyZrPFoJiNak5ga7
JnxOROjEPXB9LRGEUvn0+j8wH5EIfD1T7+IN1Y/85wYJgeYzejMyq1FtZCzYcH9oQ6la+nn92Fhx
nyT86Xlxo17a0A+Nu5FLpANsXTKz3z+k/qAAZP2WwAS1Fi/jbDKX4Ja9Dp6v8DULUUnkj5498mQL
MfgNwkd2E0+ckeXzOwuhR2UyHx1O24eAasOGrOQwJfflXxEuQQr7po9zczsXoxHxa9UXBUaLvjy7
drGUOh5bD849f845Hd93ck1FWawdK9yGnt7E+uIkmfbF6Wdad0aTbfJzXWVXRInHyDDRlu9VyLeL
eorfvhxmi1QTQ5jFvuw1Isn71bYbGEAud+LpV9pAVImtun8XSM2PAylJAKNnC96kryLSg8EZbVJA
cYn6Lo1899bIZyft7g9EiqZ/Xjm39WTo3zzUbZEOHf8LOFBOi4mfqd+0bFASxAhj7xhkFrzImL6I
EeIl7fKOH9z3UWYBdRy7kaQEYE0aEqdhe5gmLEmYtDZLw72UGjbWJ3o5KB6IPtaVRMYjjfXUWxv1
Jgu3AkwZnzVmKs7mDMJ76LOyEnmXi3bq1MLxUGWwT6rm3F/HuVgXysDkiuonZfGX/K0JwEFCrftT
a0g3fEPlR0vcOvW/Zr10laJqhk3uhQ06g7o3AbjzFtTXYRuWNNcUaEGTZ5bWLWHFtRWpmEYueFTj
xxdAilg9b7j7tr0lJaXlxftPwOpxQq58l35CIe9Zx/mBaZ5R5f2llwzUuGvt8FmtF9vElaRTQOw0
VTPP5I8VpG1A5p/ZzqMp+bcitXd6suSy5lp1XWixODRpdVRo783xAVhPRg2oE9ae6Qn0MMwZqfYZ
qDkcBD6Xif3UTGvYNdqRZVPPiGvQjtKzqET7vvPHuF1hA330PfydSC2LNj9SPNbW7edmKkmjaUfv
aNKzakoWxxzExz5yn4awcRCCMPkDnzmW8439DdinR1i8rjyCot2i88s/4DZnNpINs6TEzfD7+cuu
hOCGZ5jTkUUTj2IIqvdukt53v3IHWWe+oI9s/NQXjTkAAEUJQ+4kPYSxVbXcNqY9KjAYV3ASs/3Q
knkdx0vi3XZLglijDmC1AZae6Ku/Xkq6fPTKM4C1GeF4Bf532H7TsnFa3qS06GphTMh8qpYHdgAf
zAaF91Uqs6CqSHLxXgsA/phghlVSe5g0N+xeguXQXWi0dWbfpv+/FI+8i8oX+o0shoPS6XneJfnb
9o2iALx5A5lQbg/mcrGOzdqIth+M5FLqrydVWvAMPpTmTtPMiQlpdZORTuFZgei3keiLfeL3BpWV
ibp0GBvgFTQhIkhch+r7oX6h0HweTD6mNNCnNBLZwi6X5OY7fDd7JmmfWvQaI6sunFaTaQfhyzUa
nukLWm9zIQhXVlp5tpMWa4SX5Awm2l1IpZ4ehwdvIsM1M9Q8LLEb1zEOZxId89i3D9rmuMRRGhN1
xl8FvIXiRJ5hlP+OP1fZ5wCAD1tFKZTwPxI2JJKkVUhU3leqlWWpCj0eQmT7rV/ZaSRYUj8ilkWR
RXp88KGfPW3AuAUA6mz+N7XINDSOjTKkkYjKFoXdDqSQx3vzCpI4cSXiXJGqwvJaJ5qRPOi17KqX
CnRxjGgr2SoJDOfUTQBfR0EFw599hp75l3QEL3Bsu4TPwOyFcjcIEyYS0dWfTW4FO6l4N052Lewg
ETlRNgfIjxHTPUbxLdhcEYyNDwK8hW/LATn/He7U72FLYBnmUB1Eq5CIi5Ku/dclQaCbVZvYGDSh
ib6wWDo01ULlhkfQ8VKNtMcSzIT2Khef6Ns2qQd3vs+gAIH3FUb3OPTfFMmLPkq5CA4NYCPh3nLl
Yq+tg1JaEIezMv0/Dvps8vyuQjkWB5WPi8X8NARRZUX7LO8LiYoT+NH2WNqc2NacjGWad9B7BMlX
uzzFYJrgkN6+vf339nc/2S7oBSMm5J/SOXaX+8yNTsKSqLkmvy7dxJSDfWFR0umtvbtsSGeV4Hgw
mZumzFYoGtieJGYkV3mE3JufmpBtzhP9NVSJiFqXxn8uiBpG3EEZaDWr2HzS5yaSnB/JfvfGl/53
E4HEaJi7FY5S9JwGYCRaIwEo5MGPN4qutHP/YfWFrml/X3/KuEtx8ocDs802oh5GZvADrj9lZnlH
msqGYNOuOLzlb56axbkuxIaCSmx7sfKleqGkskCp+Qz9DYJ2OZJcG0G02tH62rpKg+++88fEAjhi
U9MiMt/ln2VHhLtWDhucZCvW9RnKFGKAwWF+R7M29KGNe2PaYsL70ctZA7bu1YCeCIEp/9tbUCQ7
Is6UjkQdrVH6/tTNNd4v1hL4swqjTMhxGW1DPPAg6banaK0V0n+MyKqUuNKfME61FBgYVgEGDrUb
i9IA+wSa4w+kNjiHdY4iOK0iREviphCpcd7EM4OQWUkSdkzKUG9wXEduGbb8IRE9LiJ/tcvNg6Nr
ykqmtovv6w/2IQgkGIrJwKNaIf6vqYhhP9FjQLGH2BOJog3HBYW9+U4hhKhaq5vr/kKHbwWbA5RB
6h4UvXUsgyjWvECALfHoio3rxQ1sSE/jCae56Noby3Ofr2rC3iyj9/j4lgpKVOaGVWmGJsweTbdg
WcgT8jn5MFzfFVW1VErkhjSpqEPo/OLKC0THk094RiBgRYEvyfropFsxsXMuDRtXHZUTivFlO6Pc
AO3plsVlhhUWqSTCKuuvvQx5utcPwXpMGRkP9iostIOg5gdJUkkD3KqkWyBrQIXxpnbersxYyVg/
miD7182aTH90XClt1QyIfL/zQV5t9/vsMPODBiytmSZ6e4nIDEySQ/JDEZESJky97BIMcJbhmLOo
qsEr8vJ1jPJBkQYoya2su2dl32uVPk5B0ecyBLignUlJAx3RSqsHh3Ln7dS1nGKrqM+S71tK3mJ3
S4N3jortOruAZ7o6PnWK6AdHLy/Q7dkiiDRn9kX6VVZGBAjt+F/a61jxJaH9Wl1erFL97gvw0dCh
X84vU3ilf7nGu21uoaBhku1DDvDa8X+M8RijhNiumMihuNG6XM50g5x8g1sbBpEmmLNzGDYC2pxH
Q43jASpawIAcfrMzNKFcVODVDshcSgLEQ+mdqMD4SsdxIUiu0O6nrkaQ+vRpJ5h8fwFT8x0YDnhA
Snirc7Lpa9BIVGiNE5n9eQch8dpiEYuLwSCCooCYXXcll4tPYmnMLMJ9IC7hzbnjEJLxbIqRSD9h
JDR6eun5ZwQij7HAqxN+Kla8fpMS4pCtMOSWNK0MCoZ8pLm9WHuXzwA/8ZwXIjRVYxLogZpI9H4U
vE0uX/nFvM3A7IBUU8wjghKf1DafBNZmj8y47rZXbbUgo2/5GrrKkjphITJVdLU6/NID5HTiEXMA
L9bkovNwVB/re/1ZuoBNKRnb2Yfnd+kSmOWRIZNLg8COWt5WPdt/VoXrwU8OOlz23j/BxQGR+Zyn
mHRDd0Aub3ovCZ3lDHzfMU8hlzsBHXbIRKGCW2Zy+kZG2p9I1VWsg7k3LYJbQXaiZIT0/MO/LBrX
BuFa+4ELhy/fNyWfHx0gVTayl+LWNOQe8CujvPFqzm8v2KrBDtIEgW4Gv2BWeEVpjBCFB2iKdyae
w9wBfULpEPrzteprrqXIXu4IfFMGlPuvTSJ2ysRSE/5X2npM5iW4hGAs/N+O/3d3opz9gZee78x7
AWttxOSwrTuNrnkupSSMPwc9VnU3p1ubAFnfpKb1PEGgRpyc0e6qlvL6GDARnwbUtTKBQOqsqk8W
07lXB43aNk6lxZEx9Vox9ip1jaJ6kboopCphqiIj8wUlB4DQoCeLJ1xcRQuQgAV089BVnuiGWoR0
TgBmoXhwCMtPicQRySCbM+lkvzyDmVUl7CbbDGFUuC//Hy6RLDbTSr13Zu+oretHAiI1xR06Rw3a
t2N1DkOTld5XDALo6DMVc09PGjbdGDhXfDLq8K7aI3EqcmZd8Sk2S/gKpyChVr2uZdLOymeDsSIr
obytUTjaOZdPf9bOVFVGKvgt50JwE81Ry1tuz3F6SgvvfWCUQ/D/bzkmos3J+zFddTzBhaTqlIbJ
0LrB4V07jJ8GKLNr0Rt6Eb7vHsAkeSgtGeLn5HHe6Th6wmnK61yWG8Xsm1inECnJaY2MJ/LHbpCn
wBr09O6+7+C9T+9S4H21FkzUjivIHBmQvdsm3zwGIrUpjLZVhJ6Y2poMKgzHmxI6QFbzfHk7bF1g
XStvsRWD4+9LYBYW/73GrI721OiqM+r8TwP76NJosGuJPvvvpef6zDf8uN+GqKct6o4tqrU0PSXg
ocizvVDC1FrB2gDlOsvUgURtv6XAHa6aBswVY/ckcPclYjn20tPR7m/7Gfcl4MtApbKLgEOwiQWS
aR/LPsnzOvRkuBt99yEL3vwLXTh14gHb9cmTo+/wySreP+KYkeRCpWotc16E+BxnXeoYNlum+S7J
dt2khWh0I75jK7KiRzmeSbz5gU1jxHVYeKAz9VsnbBbtYSywIoozqiq3kFrOY9TaMwE1RXM9SjQD
79ftkV6KUlXOskiIti8+U3aXYfuaVFqZ/hV0EPA7yRYeEHW9vdZiAVR+IzlZzyNTXOXvVXdn6TR7
Q/enqAq4JkfojgZnK2LWvHzpR5UZ6gszIkdm0yL/u45KTxFhCgpcWVZxW34KdvzLahIGBbpvOojN
Rt/dw8gjo/QEFdH+SbmfnaC+DsCIlTN5F1wdqV6fqXenZR7uiXscMtdVj3D2q/TBcIJgfEAx6EYA
NFCd1RePIuaB4gUG9QC/2wBmbB5nEwHPdPMUy6+hFZgjpOk5iK4k7mpQv75N9N7LJYpW6kn9W2/k
/mlh+axXO+yEJVB0cRYwzO0mxqDMlTjUO9WFkUfdN6CtP4qMJJbXekNgtyNfVksJbUqMz0UYnm0n
rdyxn8dSyssH3wlRgTLHumrgmM1wrUnr2gX1Oc4zrzp+FFoLD8OqifV67zaY0bS5J20zIg5LQ1ob
Gj5EhZDG0OEMLl+BmR9I1F+pWrlxc1qtazebUQ4C+LxHuTDWYmtdRt821UgwjpbPAqBupcuTHcPI
ESn07miLzXJbPw0JvbDKOa0LY39HcV+R/tA+rdRUfLe/4I72h520r4y74gCKJ/eHfeeiV+vKEFUf
ClUrdAYzaumEkdhmJiL5Z11SeAOzakfOf/DsuBA0LtfhQTtLEot0kHGFaVY9bV21XPPL0Nxg2HB8
a3n9VtwlUzNLW9S7nm5PVe9cdXti8yh82M/7o4ZUCDbq9L7EHG1n4OBspi5sdbuEXZwaKBGaMjQ4
hURHy2mh/diOm+vIKu/uVyUbKXYa6SgLyMeEPjmVjnONExghkT7GJu928DiVajFxneiK6P2w7cYO
2SK33EwU27bA9y1EMarmtG6awzOPbpE2zuGbF0+9BEWfzmqGMlCe/mg9/8LrD7YUaDmCr0JFUdrq
h+XOn26IiOH1ZZt2BQ90tXU0nkTed7n1ktpaAsTmGWNWwVq1L7ZnYrNW5xc6JdLovtYAA3DwUyhY
ERW5yaT1HJcH0hooQF4NKZLpx/OSH0zhZi3MDNT3bRq9ISMMS17IpinLZ8Fb4hWlJ7cN9cwCPRpq
hiGKnlsZw6A9yLW49c8YNjI7vPD9qxnpk+VsCV4ZZFsU4KSINOuoorXQ0lQzvkKPUWhaHsYZdEF/
HKdO5ha68NVydP76KO+QNk/rsFvFrrUHTidcC/SgmH0YhyIYyN7jwIWWjXqMbWvrAiHTX45Q5QUJ
ua62P9o60L63LA5FuxrUXK3sB3wNdoysIinUnnxmv2XjRttrH0MHTjC8Nch2vjzqtnrdx6dZMdWR
3OdVPc5BsoKKNEnYJaRKSekO94f++zvQa0J1silHAO5k1QSYvpZsUEqZktEG0I9XtwNBNrEHiqMD
Rsfu/mAl2aOkMvg3Ow4wxk3bOaroKWvutUnSe2UW20099qjdWvsGpwQhH22HUklHVpk+f7fE/ovy
eTB3BbgtQDeIWNInEIXG+xLMoSzfFGZCCsc36wVq4LkIXU1LLhYUBnGIa68YIrxKEqFaM46eBdNH
DA3j+lCQzG6cfWnKAyUSEZ2kCosSfdkHvLtATJ6JBoLKBqFZqOb8UJ3budiuYXYa21R0sDczJQcH
dkaUAVixhBJEu+KVro4GWhJtJhZw5S355P9/D+PZcbWNEbU5wKsHxxvb6X5Fd9LYl/qdt4IQ7IeA
tx+mRdghHdbe5LtFljx5FhSGqAhXfOY0n2IUOL+3DDM5ihO5xjlZPlF9f5mtyOvGNtNcnd8WHj5v
oS9KPrRcZ7wFkJ5SDxVcMeMCZszV88wr+iTm7SuDF7EaET2KOCpIp4oalxmNjQlkoreLNrKcpBxn
CyD2i/iF7pdvo9Js0L+LfY08bhu63dVGhJq4P+nQ4eAMgs3HpmJU5pUdSHFfCX5Oh5nXT+yb3rv8
BkR8hWrt1BNAlDKkY33rXi9ACN/5AlBpvLiSkpDvi0yfTGe+APkeMvP5bxlKqAVg+2NRAatAIJNB
I869aT0R0XRphxH51EWDToCNQ6gGC3kCZ/EOWk+gCYx0HBlsvrSD4+8yhyxMTCCi8JMywrOBNGiu
+fOaxGCeSo0EhNKiRIWhc5aipfUY+YEDHHBwGSEy14utTCYJKrpOesVnC1+nNdYo418qlbrSnBop
jrDdPFbshhifMsqrOG3P/sFlttHg8uRQK3RvX95PBp2q5ZpSMXAcc8qz3zTjfOUc6EE2cpkCHOnB
iMQBMTHtpEj/JRmwZAI+/3wQycjtVS3jvDmp7tN11cag5iymLGqOMgNQ744smAbbucdmgwtHFPV5
9XUJYna3A4EKlDzj8BeT8UE4HPLeyFrDodmuIAhEzFs+J69mKLSywIGLn0n9fIbeIe3fvZ9PjRZ/
LhxWlTxV9QjkgXzKo8IjgbrsoYw65o+aEY/h1t6F9j1VEDb0gEkSqy/UVcxo0Aa5aYH+dydL5gBk
DwQaFtdepw4LPOBCgbr0sygq7UQNwiwfeqMqNG5rb4prbeAtT1xUwpS19N90NCeHotrDWW+VIIZp
Epzu8chMG7h1CpLRripGAHB8UTMVLjCKyMD6ZBvTsf0yyZ9kUtyfLIffwRzhyB1dV00fCikotC3u
gZpZkzd2KWLXSVeSHlbP3qLQzZCawlQYEaPrNk7V117MpkaQyAnHaPFoeoEGl5vGtDnhLcD/57dK
WiP82PSWNbs2J3yqEmNxu2rWcheBgaeVYTJDuEsCLACshyUkQrfIbo6w5g6gKf18uRf+TTuflA8V
biPmuunwS2iA+uiri0w/Xq6gNZc1I/LYJZIYw6TZiVtyS2hvhM/eXlXXWaHoOkBXlGMxqRSOOCQN
YAk8t7u982p7pn2lz+qQOjaCTFvjfuXY/+Hqjhmdt793KNxcrIkRqX+TtY+5+A6alQaNgZG69Igv
no0K7gfvZMnWdgCxSdh7oMMlzjH6DjumBSTNtvjF1pVAt358loRxQdI7a3C7Mf1LJxYkmOREqqMU
8AoYXBBKj1UHiaVHMVUiN1yE00j92QF90S6mW9zRMLBK4emnbEqMZ+vsDLYdLjgt8jN5C6bqenMv
4HaN9lygC0gEekeF82UbhP1iYW7L3/XopW7LlYbXYsmjszJTklVZdY+YR0aEhiRWDgTvVeLHw6et
lpBGJ5+5+p+EJVWfmzERkuvRjd051yZvifX4wxg5oCNqLDhkFQkkn0Gn9FZ/3BPTF4kgomgX5cC/
lLQAEOQOeF1qxqGu/3lesYYeqvKYmuEF8yIzY5BZ+VZ2omoVjUdLZU131FPyAWQDb7z3NscaWIt6
c7NyB+SDfsZCpnhpSrNtMjMhu4XH62D0RqpaQkzrY+50eYDtjZD+JcLj1VDoNROkTv3Dme9bZTTT
DrGCl1qHCFcNJHHNVk3vPPQwmeysCOmn3pLDtj04LrSAFO5kCYVWGO/m6VLAX9Pim5DRv7GlgmAU
T9XJGnV3eyH6izydcqVuxqGV6VZETcmKHXh5HAR8ETFF53RMCZ0SuHrZq09VD/gmqG/W0yphzAhX
9r+YcGJ4iINno+tILMVHlEeFp+ced/PLVyTBfoTjsLItZi+79GjiXklAWpBADpzXMaXPSExCBbCJ
LHWB7s29kZls9ad4nMjtYJKp2zpU+v/0h41HRox84SVx+GxSs8cBd6tvONKkmAq0raDW9R0TpNa4
Kt0r9kDxw0hMr/9nen0/CLdV+XtSdbahlcundqSOU0TO8c+6DLWEibLP3+VcGkii1jsvoaySJ4so
kxDane+g8hyKyE03OohV6sBs4zMbI2/WYSF6/zm61Jm6Tb7qLXANQ2Y+AoZikt5cJ3PEM9Eqsv0r
5Pa8hxzlLL9PfhvXPqwtZ55gp1T0kxbQ3Vj66b7VMkk+0aPolFtKytbUe69ncGh97ToS3SWikGce
DFXiVEAgCcSSTbPj7AIGGvJ2TG8yLFlyAcDRxZRB9cL8dsoGqqIRERA1VHqA48JAPPoqPrlm3fto
r18x1j2JUT7ch7awufoO0devIeLZE1BcxJKLbqZ+TpP+sgU2/Yvjn5tFUWwl7pBO0hpCncrxuaW2
9CyhbhnjFe0GAMmB4HMNTd+dF+PkXqkcTyWXAJ8fH7o5RjKiihJJXz4JWxZ9yFHNxX1hGJqjVvVg
u/v8jqYJeOGFymv0aVJ3sI8ncVqMZzi6SqWGlkcV2U7l5pBTi27oLgaWeaX9JucJZDTtIbwvePE2
XnHesub477bFUfbRW+YepSD4VjikWpq0EdofK5v7ipgzrcWXiOlisXNENSAQZNk5L6N5rDt0ZhVo
GgGwzA5N083iEhbi6tBRRHh+xaC9RQCgE0B9wFx8zOxJrxi2MetHitm4y0lWH2E/JpP8R5rIU95N
liWjeRjviElzRTsLFXmeQz3qIGGz7O8islokctllOEMvZH0vudrVksNUDcCrc58W0xtB/IPoDj1w
KZunx5RW/Co+bypFnj9P3gP5/drD0Fz0prLTDQrfBhsWUsuHsTe6IBdLtqU2Hm14bErx0KdG/jTJ
kxx4nDfjJouczZry/Rp0aaZHwoJY3xvw2CKpcSr9VJ2bzmHiUApHmYWoo34C0wLWT9ygs7HXPw4h
/yM1GEkwfh9D6WgueFXOel1TxKB2BfYAUkmGw9l9oef4Wd+k88OFIUE6IQl2qkDmUoaFwaf58tg+
nconzM33f/2UAELctoanMKJ3KpN7SFzJKpaRLKRvTOUllw6vmpq9GgDU2sJjNXNCXxBKWz3wp52T
+ryVS7EEyS897OwBmjtQBYDn6aJS19K3MEkkeAm33B494IU6rtWwMX3H3FPc/+EJXDvr8YmU21cV
1ipYO8GHAyv/CZi729mrscJg26apQ8j0aYfms6H0ynRUydRvi33oTpZQiyfFuIMYBdoAl9PlNVXS
wc+zvDax0C7Q9v2d4gkVZ40LZqGvl9xF9rlobfjknB5BS469OsfX+cI56gR9Otjp7ESlB6uNV7GV
ml9hdN5URXNA33546pkiBwZKOdEEGvCb9BpqbHh38/I98Fr2j4WyUNgjCycVbbvY4Jx/y8eum37j
PSuF+ucLVzXmnN9GJxeU7s1EhijXbxvqwzdnYnPQVDoZ5BUbcNS6Yb5uWSeFbzX3MTKBCkeOxxKc
b88NY5+Y/4+QfZg+YVKVRQBfU/okcAyI80N6G7+CdT/oQMNWXZi1Y1Bs893eDinkfC/0iSeb3E9V
E2OgUGjmB3pazA84WHkx6ghV7/wFRYOn6lLvcMjPGucVgXHa+pbUz3ZxVHHXfBq/3jHiiuPg3IQc
K5gfHEKNiuHZixSi8vgsxuzE7Nt9YY1YKkvB4ltdiDIeFbtWcvzlR0dYJCW9ExlzuqmKt9lapXSF
JPDITDBsrApvo7dIDZPUyITPiatz39EsaF2E/Qdl6Tta6P+d9ZE1bczkKN1zZSMl10VmrV5RlH0X
oQm2gu9EO3gdX9eLxnoWgBtihgygu3l7InV6njsk/J6tXyB2Kfn6oWvZvlHKwiHXwBmkY1BwP9lp
TyAmhb6XsLZW20ufxP10vim3cJg3CPfL75qNoBDSiI0fMm2HTr1Uyywpohq/BNvC2mVxQfJslLSe
6a/4F5wlTGU1TLG8RdO53sIwu38I+p30c2Iz3IxzLSJv+sdyQWAqb/cKAQVsjg8eSmE5XFiKBgi+
aS1wPvqx6GQ4wdeDH2oxvw8zvJYOesfo0JfmVWQNQMimgakFS8ZS7yrCoedTVShtJgo4OMNTvCGA
9G1vFdA3WbNUF1z2wuhYcPF/iB3nztzIFBuT7H2tG65y7kb3SYwYD5Ovg5WCpeAFg9g3D4FEmZOi
LzQZ8Nf/IjU0Oz5sp4K6Do3psUf87gWO+zjyEn91gKAodJFZSq2Zv0D+wQEuskqdRAou8VoC2A0K
6PgnnFon9Y52uF+aPf0bX2gJOa6OkGJ/4/J9DDrSk1UuqpN+qlQKJiAxDefN6pZxHOvlHZqCzuQo
tcpxDCWTgDNecq2aTRBmo3/cvqeh7ZjVzoV3gmtW1T7PNOv+N/MbaaUDm/Y2fw2+pTRlBIofX6YD
OBbEKn3nC9E0nhyARK6ylfGt8rSE/y7Bc3XIyOTyEyBhK+99KGT/15iQzJu+zc+n/kEio8Uu8O4L
E8xnqKz40ahSoph+osoXcLnr07KOIs/OWU9AQ2AWubNi3X6ZyUi66MJlXVTYBWbEyF7VWGIGuWf9
N94lFuTSFEnkI315ZJ/R3NVWn1ddSo/WTdxlbhj3231IzgCHfUMHkfukZjYVjQv9MXNi3dC7eyH2
eTurtIfIbycyh+ufBb85YnNGgH3oYmKY/5Xib3yNkroSEE3lALc7hkENCxzqPj8uL3Kv439UBLLE
2R+u3j6+HRmh5FH/qfjMYmUG37U3iqGchd2zHBHFlYahgRg6aHgXD53L92g0Hd24F0cAPzC2BbzR
BFvXIRrg9gHgzxTqSerXTkop6ZUSfChO2aleJ3ru0YYLCqhzCuFO7iZ9TqcH49aYiSOtMzlwDw4C
XQkToE2jMiQYNHBtXIaGX46/6OZ4SwVn6igsTCkzeA62A99kat9olniG3IWzbXAY6ltiVbVl8CIe
QCw4ICcVP99AwZKioRB0bQDBHgdZZYAR4CnR3HAXxUPAxrMckTof1cAw/8kyCIk1rPCoOHeVtwtg
tCBUMWra7LVBZqCjFi8VkHUUYuvO4FWSFm4zkLQHC55i7CnD7RFeYJAXect8EFCJ2NZexUIgRgBg
J75iZ//uclYQH4xkGsKf5ZPJ2YP5k/mq17oGQhwMIbsinUTR7wd1uW0zvoBhjX9y2KuPumq4ZTTG
+2nDeGKk0BFSdPTeC/mqoHu1Ts/ApYcFJV+bYjJ0f9UNe0aRtwCcZmCGRTPcyy7jP1oeB0S3Qe9I
LQhr3pellStMeUHqRrZo9hB4x6lJIqvC9J+CQuN/qaeUwq05npV5j+q6bqaXFBzh3ytTdVA1GooS
WSpI4NF99s1GQeNs6DoUmy442DXxp1LIB6vlrCzufKb47hxeD7T37CvJFR+QygWxh8c3vHwR9Nj9
OvvOmBXF6KemSU+UTl7EIls7WO25x9PtDzEBWkbqRKoGoueWdnIYXcCYjD0XrgnkLKNiokiYf8vv
wfXa4RY9E1/IDJ288F5SesNrY9jVSsZc0vxd7WlTUci4cX14c7G42ScT7vhymApuudKotoKCf/gy
gvEiPGYvDr202qQvN3PaZw0q9lQpa+keyXrCd5DZx267eEDu2WoLHFFmtF2HEhq9mVx4P7LTZ+Sp
2Vx64xFCBNbckrHA9CRDt3YgZjSvFOZ/TYvgGSWr1NcxaJwa19N4ZMF503RCG8G+TUW+ns37mpyC
fWBvptG39883c80XRQWEZ3eNVrZNqAIPn5VqwW+7bWn5TWupEoAF6Y9O5Q6KIs2Uo9tHVu2lyBVd
rp4aBgezTmilvKpjbAM61KCDWdMa5zXh7a8ZT8K/vKE6RYWGIptsgEwKGfDFNqh7GiHyGT5b1T6x
BSUlv04df11h6PLW9w94Qcm4AGuQE8AH9kH1dIVjUdyWKDdDo3Qa1krzjNOmv9/IOwASZxc2VXir
l9rSoITjz9IUWag1hvyAqNxTTe0phkld9hovH3rAvlIDfJetJ5uBdmN+z3HIqC/KXQpPgKxgrXsO
eg2PcSDQTTIn+hIT4nZQKhvWLjs2oUQSRyX83+5lAMqQuLmdWsfNnljSIH81N/m1hoW+GhCzBdrI
1E47hxiSpma6FOhUjgTcAyvCbXX2/Q69nqZ+ZBkn6TcfMmJNnXYgfB9204FySt9FA7LnAja5D6p3
OmmFG+P37S4dSXPEBWzIic9TE0JoIRRG+R7IUbcF3ZZz99YzjwxhDwOWfZYYV9grzW8sY7UNJ3da
aNIrr6Mf5k2dt55TfgSZ2cQX7oz0ALJQOcodjcN2e4JXx7Ak2qSju7/g61XFekEEQFpY8Cx+IP4H
mnTZs4bYi+IA7fMXU0RsjwFDGbr8WMmfUhv1AyprPZnghuZpCsPE97m54LhfewKLpMN84xRP/LS2
O1NYdnXQr0YZh3TnHU5hzRRPjfUPzD25FSGTmkYrZN/wqgQF1I7AdtScDtwVY1QqYOZakXOK27TO
T5p5SJTpKdULdCiRqEXAZSOU/pJ5aOa4+PLStaWt5dCPpWtOWUS5UAasCe6ykeuk2SQRkQNAO0rl
Fya7XmiA6rCFMKa9RwHEa0NeDMontY5vfr4929hiBvzAxrl1WzfxbM9M93780gam/5IoP1sk2ujB
asxZXrVCjrIWC6w3KJ2JmZgvaFyYMsQfrZjlatNLfzIUUEXrQjuhV4OEXYq1zouSCYrQKrW00kR/
cAarC1Wvsit5GTaili+sEJMBoNfUsnrc1lLH5/OKgQjIToI3Dkq5zFznuFeWsQDdCLo8JGn7ogtg
gjHuihM96H86HQMC6oLJRBxK+OSZGO6lLp+hYp9KxA5JQ5aZb19f/fMKCV/DUiSbmTvJQ37MjHsm
ocly1UFmjDnfOzbvZAbf6HbgnwzMvvaySNqXrm74IAzqx08HSSGRXyPP6EyVz4FJTRGALAoHsXGX
faeFLv3O5v2YyFOMqdhQtIedx1EbZ3STtCi3XngD6WTscZD0Q93f87NtFrAn0YOkezEpK9UCx5S8
YhbMYipYvykBESbYDpOH4OCL3eob7A0PVTIOxu1b3xIYVBfeRTxuOJDW0kVrgYsGkc7WnyDPv8EV
2cMXRUy2+x8bRpwVu7wzkbhwhzx5ZTQMUJGu5du3JKztrGsSgszeBwIkCNcAWL5C5GDT19uF07hD
NsR9Kfx+44nf1gvGBzaE6jDQatSFicSkTEPfPeb9pFStpdX+DXpm8ylv5h2t/pl2YgEEZg4kYZBC
/WssCmqyCz52A3UienOx/jB3zIvMZdOVng8N1SHvpq6oel3u8xWZu906/FhFaZYOvk6xsSHz7/f0
XGboTFpAUCcMhqyEx7xJrIUubwFV9HHx5EFwgUQfKhyiFlOnMjMXq58ja10soknzoKy3sGK1rdJh
27q8qBukWeYDXGpFlwLhVOyWVos13gXJRMF2WTCODzLoeQfB+gRSK5UFO0ZusL53J0M3SPa918kQ
s7oEFNIEHznInLCUEmq0csY4ItEE0j/3Z5qSZ8CsgLwg7YqtL+XxPvWVFdv2ruKiA03K/KaicQEZ
yM1z4+uU2LSDw694qcH8bz7mhHhASJ8vw8VHeUcA8OpT61Ov+wPZtSiyRDoriK9BBXxbNuBhAkDH
pzBQTN/KdFUb9Rm38lTicouMuXxVl06qkPuhPST0uD+jkUkn8HkJCQkgsRFBx++ki3nnyeqc0hzB
QVWyo98udPrZeKmjOVl5Ez0QZ/9oiW8n9XNZoX2bEWgCi9F6seRt/7NVbFrEaiFXlPkxaRmV7+vc
yosTqwf89l+oaeZFZkvcX/1oxYOdo4L9OGMMxQB03iUPF9fOopEEcru4OSkN9aOU0dudhXFr360r
HPLDxiNsP/AcCcYSpS6GIhCtnJXcKGnea6fE/mPVcG60AqFTwZkCASCGxhmX2ZpEpJ3uZLAwzK53
z+mLtNQRI5c9vWdjdhfya/7KRBm0k/ZmT1zwEvIEJw8n+OfzLk94M9Ww6WRZBFw2qGK5ax9Ffn3h
E7kUIXBHUjBo4sHa8Un+CgOom0Uigg56gQmqjnMVpY6x3XtnOizQLCNYHXMWFYF2rG5ydvOyLIae
jXVPNzOjKULRnjsBOSeJiClxPnnteLcuUftuQs9Pb7jMBQeja9eSqvNZM0/K5f6cQF70YrqmtQ3T
7HxQACu1EuimIhL+Fe/5Ufi1NFuTZx96ITekYKfkYFQRo1p5AXRPNbXazD5X61MMBK+YHNdFWP84
5IbnM3kTkWWFUNpFyL9hAJoaH90v/6mYa5Euu/fn4dJLKFxSIGryEJrJe/FQK1xXoiINyXC30AUV
yGC7BPzy/eTAzJRLM++celz2OebBIUuvDN1ovBnzH3/x/p8yt4ADVnNuuFta7fbKHv+LUBRUi3Z3
0qy8b3IiNmZLC68vu33575DoDinkCkGDHpLc39jUVyAWm99+2PED/4dDjVwEm1gb2rtu5f06RH7p
wupklrRqreIf5UYGAjwUzlxbNWK/MSwYWJH8ZEt56kosUWwSLeSwRGinI8uhqIUOSg2wiWNt9G3N
bvfOJt+C+ELO2Nyj6VZ7wyO3CiriPzPgnZFhe08Tp09LzO7U03jemkfFF/LOwEfXY5cn6DGpig3F
itExnLa3zvizc67Dz1/jroXsnkKt3PNHNbeliuT5YbDbJfiq1s7/rbF1CYlBz+3T309N4OHg89de
qCNTv2Wcgi2Mq9f+A8mOt+MBpNBMB74rSY/gPmk3NErwF6023mrFIapTmoK/QstSLLHNyZp/WeiX
YeSW3My/7LCruAMm5nrFS52nh854QejE+I9BfrL9OR7Lcz8KFsD8nwvs/c3BCRmJ5VChDGmv8hd1
8jcJ7DuZNItw/HYLGDlLnUf8SvB3PkgeO1tWFR3r/HKBA/sm7gcUbqQHgkMYt5XmonmXxTlJQX9J
80YZth1+NlFYeLyPBNNsqV6VnSxaBbbdFm9ZNiDseTqoLSHgbLteplLG82bFcYb5UTzj1Iw2TClD
XeXQ+Hr9ewvwS6QaQyurYvkBGqUBp1dj6GemK2wP5/EYHCaigXg5a7Rkh0OdgM9F61zVO7zb5Kzt
e7svqgpiSvAZAH/q7VyFJ2eXDiICfV0otFcdC6PEPXeq1lfU24WlpJpJTsHMMvXn4H61l4UcAjWl
IA8XQh4BLj127R/w/jvyBUP1anb8N1zK3nTukq+AVkFtf8dK2v0CH3pclGnSXe/z+XskglhvlWfJ
dV0iE1MgtHvsvmvftzvVvY5lXG8XPY2JM1WvCr7xM/B954HxNgiCpwcX1xNGcWqiAsmolBJtyckk
hzTqF2RBZyBNNnSkD9t4aK5U9pV+9KhAy/WoauVb597t2BE26DV4VfiyP28DdWEk2rvXPREJegaT
DT2V5TaIiMWs0UrQOx2YNUJPiHyhBQsUcw/bcOtnMZDtmc0qC9eM2RTX9/LFLJBbwjrvH8avVUsD
3I+gIXjds/oo8c29uzKclyQeey9xketxGozLXMO2Xsi3i34i1cKMAyZ14IUKAucXgpQBWbGVtNmO
Fe6IkxDukORnrXuJPAbblt2iRiVjUM7rODWOwl8A4COucOLI2G+xyvzZB/gDXor7KWV2VR4wRuVE
4GxPHYdtsfTGOOUay52lz72g2NAGplpxvVH2twIAvNxpp6HgBfpVtVWUKe0R3fSV2IYRBISFYS0y
z+SYMY00Se5agt8MCW+WBTMJiUJhH8VWHJ6sUOSNfAPQfxaqB6PU8l6sfp2JyVDvrOOQwypsBxTI
e6Vudq8PpNWu3x0t0SyAP5bBWp1QqZ7EY50sMSHuzw9IDTALkjX30egC3dwaaaF5S3yaoqm49D7U
cUOv5eijjYib7x12geUw23IOClDruybanM2qnRKYGTq/CArgWgNN4zooha1y1+Jhw1fTlXp9klLO
nVpKotP8t7sZ0V3N2rmRoH6wHtfNA8vVXnxxMsGUl/yYRMi1a6f1nDm0tuMDcbibDQqbhNzdhuML
RMs0BXDAhyNMlWG0A9JOjWbbopEZFROT3jEDV9WLpFMna+pRl5coOiGbSXe+560ynvCTl2zdps8t
5V7aWl3OATX9ptIKyDyrzkFAvP3qRNEUs983sY5aZE1nwb10yGuQCpVZumWOHYZu78X5Vde9vqKY
7tH5PaCt84BGP60dJr5C4amnXzStMxgQUtPSoL116T6pssX6r8PHQOUMDc2JnfG7qqp9Vsh7nQGb
0f4mTo4nzon98pn7F2T3VOPXzG+Vgtn/1qbvvGO2msknhP90hta87OMVsgi8eTBQh6/YuIWfkQ6S
W6JJy7tRJMb01e9D8cLHLQd7CpReVyvbHy8nnLsIfbFLGMAfacXb++WwFK7K/VLdDb9c7NfPHyZK
bFZibs94mL3bQ/OpB/cpkn3WBzsQoJldG3WYrkh8pJIe/259+jObgwk7g3aqCV2sZFp3WHiXsZ5g
RPOuJEw7/UTWOubgaJDERsspzX3mGwrBI2APbuvjgXPkrEi8+ObVjhaA/MhmgrMEv6zB4LM3FCH4
gVZ95Et7l15scweRRzz4NXT/Y64nzeejaFlT95BTNhF/ay+zxj6UkxXq2b1L3bG5TO7huBENcHzO
TmXxVzFa8V7SuLPC/SYnLiFPETzWSBNV6J/rdHztY+YaWNpXTKquJ3BpFn5PwDb8+U3HlqC563FH
5Ai1HWUz7X9vngTCIWT9Hjjo5yWmqnFZneguGR+gKOEggkC+yPaanFZ2nIM2cK0sZADIc3U6Xm1U
UDERRUWYacsJVh85xVAU8EJp2mNZDtb1BTAvEf0KtZghOzO0VAEdEsJuvWXwbm3/tkwV3RJWq9i9
LALWiBrUPbv+okpm6zt7DH7YeNIynvB+H/Z+qK4pim8SkQU2KHZwaCiBFOpLlGfasFfvVDkH2PN8
MXfCoWRnqpOIIHdsO75+LnX2HVpVhnibyzsmfcv8bc6qqqFKnkFIh0TSmk7dcelTdy/lpKBctgql
DRj1pbiE6h2SZ2xy5Oqiex7UgryoQWu0GfuSB3OxTjMpRYimpt8UqTXbwjFGIgdTkGYQ6mf8IlPP
Y7DS1Iwg5xZH00K7Mzh2N8a4Uy2C2Y5ucfUyERMaMTU9OgSwR/JebbuUrvfKlJIc0d0Swp0KSjxl
BJ7QNeEi8aHEsBKmMZVD1v90L0VOFTpWsUaHdWh043NkhlQ+bndyIoWYm3F6eJj4a0q8qfNZA6tn
oX3V3qJ2sDvIylvB89D5/BO8nJKrOxMfrcgqf3WftM6lXcZNdb0eeW8GgLc093f6vIs73Gf6QDyR
VWRoiYrEIwyKqXShUopsTlIA9Ywwo2gcECiosMexDWkRPhcRvpYC9RM8OHwy+/vn8DOJqFPAs7Av
28o3irA1vtGPZZwFfSOym/MfKUNOEt9yCigQ8WetoawgH2aNRsTEWL/tVgXE7Rh18Pwi59GcMxAD
fQWzcMn3q2/kAgfgEqS9yuBgkC4cXtBt2Ql0MtZ39mpQs5pB8LCNMguJ0e8hdeL7hhyDbUCAdXQw
p6aQ6To7kve6a0JontujGATiXVa+LQ0BT7mOYap8x5CnjCHNwI+5tuAkcEMcQVwiPmbiiT69R3PJ
llG0WP5fGLEmBz7/JiKFuJkfkd+LMdHX2+EtZOAgO9/SlDtZCggvYyD6nj6VNFEvMe+x/4yeDS2y
wBfGfDa0YFGIzKVtGBGsizeWwMxpLeJWqTGKfjjP/N5asSUKlbO1lBQWvvuWHiyJgi6b7wTVFmQf
VGV/KDMr+FMmG4Rbjk10fsQRVk8QurgM4k+P3R7IiRlVjYBR6qbxw2Ywmx2wJaIggJGPwi4w6wz9
jUBl/baWudkY2EevJemSZ3TB1N1rgRsSp6/d5MYiiWtjHgF/6/uQBfVvYjIVENdvv4vHYLuNIW9m
U8CozsSmhQLEQ0S1c50MLNwH3YR3IYgD1LqfKg2RWRyZmDKXjC62Pd4pmuMSwtkZLC/Sn/aOHXJ2
pIKHn7i2s5PpOScXvkgpb8HKQnNKGrBjygu7Bnx2OwjLtzerkKcPoiXKzv6uHkY1LK1tu4yudcKK
AmleQ7iOZwGhY5mSyHbIR60ag5gH0LkIwJkeIUhDIwhBYMMECKxkZPC/53as2AkyI4a33sJGuqqa
4B4SCuqxeBFt2w4k9vwhw29vzuDEp9ORyyoTnJQ6YgPcChoHB8u/S5gggBkedJBC3/u9GD7ocD3n
mUV9+LJA5hGoImysNzQp4de4kNpTRrSuG/2TC9vXVseURouQuxJiN5BY3QpRVfch48z5UyKMPvVj
spvgw1El+LUDjvxxQQJuseI2/WELZW8xeq1Y0QgdyUKXleKeXS9sfaIuJDHCDH2yF+zC99js6ip8
x2nrCDzkFaD3o/aIlv3LCzLsoj8Eo8Um/8uC8ORL5/RP/gC2I3FtCMX2liN2G21o4tL1qy508RBm
evUB7FZ05M+KAO+c6OQuSw544RWgR3Uu2EJNKPAD9zawMKrseMTBRzadCOBT6NJkQTeKOZ9Qams0
LCtZi9yr5aqYaPq3WxNRcKilyaDyl8wPLJGqgppqS/6z4ve/RwmujOvIqc654JcPaLhK75AJzvXO
Jouxe1bxgiEbp9kQZUfcihC2C7FLj0MwmycuKypEpBbou3A5PLOmKHUqJwmsYGJxwdAAe+v4fUPV
13O8QpLPLF2MCpevM/1bkTyrlLdWrw48WM/WpDgtLzzjv9KKBndXcCxO8CqS1au4wY9V//63vK2b
+4908MIjSObDl8zsiZa/JgnUjgbebuE5c7oRa32UGC43EUp+Qyj/8oYFzmoUcmmzfD9TZ3b2t9qR
5OmOpTIomCksqzXakn8vmheRxyVj4tNZFHbiK5bs04Li8gWjtWVfQyMrfQKPg7mrShIdxKwJtpTf
wDRg3AICCLLd0hPFykt7920R8dbS3fT0aTr9KtehigbJsKQMacyvpaYGWDSkeg7J7qKRteJ4iWIv
mf4I7AGtRsMF4xhHjHO9qX5FERtiwmerJHPqTy/Pf1aEGucQU0ifpSIpMhnJ2Pen8wDwyx9phFZs
kaTWAyXNBsp1VJQ6ZHcb4puzkROWRhoP49K1CRhDDTOedG6qkrAZbFhKYxsqvbsM8k+MF8E/tX2u
l5mTRv8kRA3lRpL347WrlF4OVREdjVc99Ur2U4Qi8OHVhYQ+QQPdHWxyQA6aBEgw7Hwf/KT5hZUC
uJHLUI6iqsBgEnv1Sl1g8alefq4T5Ic0VLsS6uQPNWeq3f/aYSlk0oA4D3QDagnzbCOe8+pTqg25
hM8Y5WOpsYsyio50xXxMBseDGt3hwv5KyovUP4/QurKQiaxnGJtA5ugOm8WhMQCH5qafKGXQnEcj
/GSnJzIRnqAAZjtlnr1royfNNZDD6GAyWC1RDmyaL38W2dg4yBq+jDyBmEsD1AkwGtcuUkuNtU8n
xNKp+AzwSt0HQe/cuQ1iqO6VmkNMsdppykxa8lIVUWCx4mTiVTro7Rj2pIX7weVGcwehb653RaDi
T4wFUPFv2xhBeBm0pFbqwHvBLfeU3eoh4/JQnMT+BDF3W5au/WSCINGrVVmWGVkaqCoy0fTQEi6j
4Z/9vFAO1TTeee8byba6Y+9jCks8avrLNBTNLPH35WUvoLotx3+cdZJQ5wVZmPFfZlnJ+MjtyCal
UDB1MzD/JAb30tfZXNnkMqlXJd2tx0TRQFLThq00yeUrxqrVnTCx/jPnqhqQk021IrueMPKsH+iJ
nj1JE3XANyrDUUrHd5qcNtke5Cxmk0OCvXTaTNuIDtCV2FXUbSVwh8qXQ2FZX87N0Yjk2h7v5k3z
EPIvxA7eXHm7kOXuHur8jvJ0xcVVSqs9xS8HNEd5JIj/IEqhHr1Zk2BpKsXVDFfCq9Kf8ej3oMRj
LttezquEsaYNR6wv8CJf7XeoShGP2zVdugLASIbszVdIO+1cckwyxs/DTa8vh4z+9qLpnSZ5KI3x
ydBwUd8b2SYHruUQWE7tSYisRbiSnz6zV/p1QwM7iuydmpsaHjStMs1pdz4/OoZmV8B1WITdQWyQ
oS6XysnpNUeEfSWi5/Zeo29+1KzaQFaxCP2cIOW9a9zGMgDD49uVrTsO0CysaxkhT6rWK11U+NgV
QVZV/VpLT54QTpM9iZlyanBfkOgrokBTGSYpeeoEGpZqvVSDymA2bD821Jbpqt4jhQuOMuB1TH0s
MjWB5KfvIdTmQt4j46rLENpKhEka7rZFP69g9e/qU2Ri/kl/ekOcfJaruH/ZjTX2DqxB9wvkzToq
R+P4Ddk0WqJBLw6ZE5llLHrZnNh7M6goJaVoAPU/3NeBfiX/339KetlfXjm7V+0do4TzOxs1EnRP
+LbqTPr91LgrZzueawISjypZ7h7/E6hYA17bMJG4Wf75QIvQT62SOXWEggt6ErdBc+laxRGVkjOv
bENe+KTTCy+y9roV690AY9XUvKXF/18h7PpT0Dg46nBwCBP0x2mbwbp6PnIN6/Z70/yc1+wYf3V6
TgcYio/jgHwqEQOHc/gX9KRoFTnt+iuQb56M2eHSe2e7ZBm9yBpQRs7kd1h/s1gK73VIazqrQo8C
wI168mp+AilwCSJHZldEKVsmiRMiiMI4veaikokojAwb8pRjRJ4wCvJXqNDrJOgU1OG7ZrGFpZ5v
kucsOqx3ny/990GRHmP90d8zKCzuz0GCKeXyDWxq4HPjZ4CgbIbhkF6L76U2OzhMCfcM6UjPL2Ht
vVIV8+8mmsHp10MZ/or4ReCGTRbmtIe/wGT2MzFNqu2mUjbjCKGMoJ0jCz/hAL0XzhUA3NdwTV4r
Xo8X93eEiYRbptx4/9JB97WAuU+kCtaYKb+wa4/j3bqOrYj7lnZpzHbLLXuK4ieTbeQfcZEUfgN3
6H8rldk8Q+Z96V2Aev5CIDOpKkIp3OAte6udcnN3q/HCxUP2WFnWVznHb6eNj46Yz+g020xw75W/
9vi9ALUhjZ+GL908VvWTMAjtI+ztYZbm4RWkIFVcx1nZSOHEyfYKsr+amOcnjwVloB9o0VM7+s7n
pA/5+KgXQFWFHsMoHA6axDl914PzLgnTO72GH6BpqBpEQdhSL44T1qqpR1uDZgkNXwLc3e3LEzTE
98/bvClVYEyV7lM2irRrvf1E5a+U/qg2oQKiwHmkjyNHrzXNGt4oRIkpRwYmPB/0CtSM1xwEAojb
mzR+3cs1X7P8Z94k/Ip8pBffEieM4CrfpEJpEwuIpQ+Ocx8ZDmtehevcYdrXR5ARzHjfWITI8iZj
AietiSlGtd8SkyFyC54UbZDyQSMpGswC33qcAXf5FVMBOCngcfPeywHvKyWvMMyAkMcIbyL+wXaT
N8Sk8TWCnq1mFKEwBVLb9eGCxQQbD27pTxXChOHCvy98gEDRcgKt9IeKWxfHmShmQSVmvjtcqlcM
o7grLdiWU37oAebmP2yiv7f4fO5JAhyTSlKjQqWYuwfc0Odd4ziIggYbI/7mbyKrGOPbFoePTE5B
w4zwaZ87GpCmVDPAoFfivfx6J7UIg9iU7nnyuClJ/lmvOYJwhZQPY1ZJp752Xuy1yNRo0tTzW9fy
9xdcE2bLmYY3cZiVSrgGOlqDe32IdtN4p/jvoTKbTXya8R0F3O4WNFOI66Ejx60OXTaU72hmFE0Z
BdtgtxZoSO1BtnlnCBFEeGAnz5lFgPkCPKaB9IS/5fs7DPPDV7amQSWvY3bia5nIxsvVkVfdInnt
r60DPr84eQWj986KiJoNREqtGD4K/7+YGcugDDbnR/Q+ni1DGQ2a4xIve24BB/+CTEHN9f72nQt3
LkhRguUhm0uZg2OEbYjauPvaHERVKMGBkQk5Qw5po79qLO9A8toetFy8NCDjdHfXfHF1F8TZi6nB
AvAlzdMsnB3DvO9QpD9G2UGvY8JViIXjyunixWeqUCoU9CZBzNWfn1qNqmX88rzb3E5bXEV+OaAn
p1ri3wPHD3yjlLuwvASwv0mT10xlYy4T8hb2qZVfDgiOqkFfClV7t478H7RMI2sLmXRngk61Ks1J
FbQUOOYG6rVt/7RMfMukCEHU9uFRIPOFfTxkoiOSI+5n3ojqgubNcq2jXOD0tNIdijzEhdu4dduI
C5Lqb+5WEbHm66+suaonYVsrqAaiebd1Yx7wohYmV0flJJpnc/IgyABBtIfKPhFH4sZ/Y80pNtdN
F8tziO3Fe4Ju+xTpxxI3xVb5WYnQYOJu06R0ajMOxe3QVv01shE1Rx2psxFMMCXt3iyOQgcidTay
qtmLuw7RCPdHbCNVtc3LeXHgCL5O0+2YCVLs6X6QxLXYz8WZxngBdOE1qa8KYBNSAP43p9/oC699
cPGop3GtG5SCvejRAvHZduWP7UZsvtzOg2vlwQ2eKdfXE7CLWPoCJxy0G1kYknxsRp0DLEL5BGTp
HAldQd1ajpst5K0XH37LgiKBQlbvYCFJGE0DvSeLMcW8ZTSigPP6u3DPgP6SIT7O8O/vwLgmGwXT
1HxYlEqjpCbjTLOZ7SXqnj8waoDFH3F9tX4KrbfOHbG6I27SAxdjHa4pyjL49oVRi/Rb0+EuIWmP
C/VHqTWM1c8q0T7V2B+RzY3J4rL5tuzfIPqqy/x+xIqiecJ9qqwRRByJNdGZo6aAvXQXLgQBmN7n
X7kaWd1l6TLsOPybORzYWoJycgtKl2UwjQ/ydAt9y0Ts12nz5JEs2dUbJuzMMst2q6WY58NT/8VM
4nAYBMJw6EDQIdfwGYObdDgxKybXIZ8zKwQ5CB9KvNw2bNl/zCNIB5udx9kkgvZFuOrXUfTs3M4o
hcpL3/zn5DgutVtz2RiHM3oNrNxrMSHR0A2DMeRq5M/hSW8lmghw065Cse0ojtK7ERGo93sxK4AM
rYhEm4PtxFEV/ubFrQpLJHnNueYpRIs2Xqv6ZBc6KeKyqnLKplZwIhIJVbc29Z2YTLi3f/dth5bn
zW+cXx7K0CXffVf8k6ChbAcNB6O3FSXuF54oXnCs6orXrJ8jxIOb4onpcR251qbF3hat5R8LP6Pz
mf+YXruOI3vDR9A3H68kQ7Ad54FtSO+gXVgHOJX/EFHX/d06d0TwhGqxfGMKE257jx/lTLhpnOzx
mMcCuTP4sYL5aEr3OXU3R4F8LVutrimzNMtxIau2rewmas8kOblrkLHOrl4nOOFmorFCwfXGcPmy
uJ/TqOHDmJ9fp5i/uI3F56fg63uHaJDTR+FSGKPp43b52RzMKTV0CGypIuYKhzTJ77C6Vo7bfg+w
eZMnZr/RT5W+vYNIiWMW4WKimlDY7pGvqbkYFtG46hzgXVIFOYCU7X7O5ZoTxBnnTlIROLI0l/bw
Ix8SFIF2x3CyFzE1hF8TG7/d09RhmF/syoC+Nnit3kNcSmhCFb9TvWGMT9e+0GalupNJsYK45XPV
+aOmqFSt3t0r7xx6tHg4JLcajKPg/5kOpKov65EFBnmo3MNRT3mvFx6i96fPQlnSA/cFO+SvziPG
StvcO7RnTtBFhl668drkqRGwzTQdKrWkuic64Ok3h5g2QSg2P6KH/deh6xd6BVk41uIcsfwPvO2K
fljL7LAbx3wkotF11a7rKZAtP3+bR/G9NtuBPI2z4U1H0Fb26Zy8OY34vrxGlwpmZZIucl/KEYGE
zXslH2MjUD1Z+i22+/Nm4eQVJLS6YkSzDj+WmfhRL25JU2CB7P2wEcELHfwmDVPtu6y8mCouhfef
e6yJGW5AAOPOJGDyHZqAutHV8H7I30pEC8mSXjtJkhl10kio8eZAPlsQe27yTbhApC6Cd8lYfGuq
DE/l3poQrAXG2oGMy9Z5pXMupmD8nSTmHfDqis91qSZwdrv6Pa7jDCk3KHqwZyZWEYo5QbtaN7AX
a0UsJVMpvNqBYG8KtsE6q8rhmXHgdTXknqpik+lauSl6/eLpUOzNkGIu8+LjBPeDW7gOEjt7e1ER
dD81fevRtqJ8I7lMArXeGxo71+Hqt5HFeJHffjsZ2QtVQgXjdgc2+4s8ulJAyQRW3zBGP2BR60b1
erLTS8WC3/JedUjPSubzt48MrJFErdSxeMdR8N1Lis61Hfnf2X9bqBtnIti8xoZ0vclJawKbXqp7
L7/SCne1zJiNotGiYZyisCBTW1dnA63MFEu1uKvYPVRuSReykpuEhctoxEk5NA9YX3oMBghHtHi3
kG4aP5hHdqj1W8u4txUXuxQysnjlFlo/lhMfvQ/gZApDzeFitHS96TYYbOMUtnWyEzleUIGyQOdg
Pw88C3jgS74IXgzuoDBVhtOftzm0nMDEDshg+SSE8TuudrfcNBk6zuD1pT7tXsmB9naUDIaqMadK
i0Ftkm2aygxd2t7MMS1HLekBPs8rJj2bLGwAfpETLCAK+pD8JsCqhzoD+2L6jyF7yWtn0GUa+mHi
Fe2B88ayBWI7mutZLPChRRvHhVyn/n4KaOjnYOQnPuWfIgzDxEzjgd96wkWe8txMGEs06TvCYiU+
NHAVhwC3MZL1EHiLqm6u9sRIQOz7NdFyyUPfX7gHj36bsGaWuLaSNfRQ7MFSaIbXSHiEudDecrQc
io+8IqoHNY+hDt8ZxkrC6ToMveZ+BsmkLao0rOBry37eoIKVDQpGead3yWfkoVZL12hbR1IVtwqD
2BKvU/HarNoNdNkCfnQsxE3g2UfTJtOSZFRc+zV1l+yS+Kyoeb42lLTM1MUZqM7VN5O18F6FCcR2
gm9KYNnWfm6BOwEIzO4EFkCgAArwVNyZKTTgQ0rORnWE5RQaioKSJtq1A1AfeM5OI3P7+Kif+Xql
e10zGQDDnKTtPWcszFa8TJRoZvFDaL3gGagxHsQS29fzX/6tnQRlBieSMdf7XNe/Hr+UWhHybSad
ZOD29Fnq+Y0vo5/dHLJ4BF6uG9/xp3W71LA5POP53gQmdpW4ZeaNoOjElBuc8bNBO0kD3QvPEAQe
ZZ95S9pbu47BM2hL5HEEGWYFdx2VTPB5rUW9FZU4yTRQzpCTEKEE7S7Dl2i9tEmzw5NhOz5BuGfZ
G1BzmDZC9cYFHpH0QFqu7MuACPexZAETgTrd7D02LktheMzGln1yoZXQJg8TMdL1w70cCMBaG79D
661mfwdK045a2XVv5At5gw2MNpqIHH26K7jvJTr8Pu86kOmib8dFTNBxPRLEBd2yedzYmmAS9N1X
/uLI5qHdkiez9Yl7D/C9i5RoUoTsUo5zhWu4H6dnttQiKwEOjadvNBI96h6aYEncS3htZ6WAxp29
7Nt9nXodg8zCo7x286CW+OWjv9sajhHCOD7LJKqVP+PauJiiXOOj/dG4oGwkZW5BvYZavKDmWxll
OUjZ+7DdELs+Xs0HIfZZeSUdcX3TB7ioAKUuf0hgzfeU+CvnWFGDFW7MiBOOKHcKhStkCWzUCY5j
P5/S/rPxyn4szwFVfHAcSNS4hIlxFmstxwFTnvHw+nL8Sw3yEWTPQmIGBtkxa5Die5WimtAIAxpX
TuJklYAJLrelzUGyL9SyWy6o2XlUog9DYliYci87Id2PqVOZmIBnuQnObHBy0p5nWMtzNZVAKcLY
PNtDQweM3eL9t72b5ZbGKweTY8uvcs63GsAdqQQR6FGHd5c0Ro5sKyTzYjhXdmsA1v/PLq8BR5Zs
h+tBDNztkodzLNej6wFwt38NnwFY+LGufcZyabo5mCgvMhdj7hPKJgiFvS74wwxZViADbZqJLLhY
ygq5dbKPAPlblkrxOAnTQ0tbgigGz9Lhvl/Cmf/7dOP+PM4nvH2iZ/F23gZORC41EfWyQocbdXnh
C35mk3q0cPBBUycgP2rP1urCaMYUbxpJSf8jh+rCGybxn2xRGNns+Kd4SUsM+iwh1e3tKKzUWBkT
oLP03kDdOuJO214TPWYnYlByl6Fl5vvNwboNO3SdHCMREx8pCRQm3SOMkZjFoVte1/Tra7k/mKJW
GOhxnAMliwpJ7SlakFAK0Q32xmMvBvKEoFeKiJrmBF9NSKr6MZi8Z0IlsikMK6ibVaaOmMq5O23I
SwoLZ+jeA0T4pxDsj/vOi6HZk5cda6GD0CxVZLvnsuCl8p6HyPSZ0XIM6GZDd+TezQWpluUzURoy
+iKoDIP8Tfs5TohWX8web6SrGnJSH+WyEhF6SuPXcJr4T6wdeiRROVq+TjB+Eu4RSGT5Ja3zd8OL
uEa6rHauJoPcU8/Axw7cVApEILYp/OEaj0yC/vOJvy5320LtW2hvtzQx96c8Qecq6/m9VOzDbqHb
pkw9ehK1adortpYRhrof7eThN7A1QBIBofsJ0p2kLtp+ERZWWgT8QpeXQk+zjsYzYJDOckAx5CEH
x/2O6CDoWRt7PiEXuZuJuekqUreDx1a6eoH2Rx0E25W86kCr1GVzbE3CVx1tBAcj/xG2m67Oe/Mq
vW5o70zUvSYsY6PoCkDhINmlV40iEbQ/XIDbA9ScmwTmoj77lBK7gQwKJ+W243uFRTZvWIsf/fy/
o9nBWqeyW/hXMtd0yyNH6hsUIQDDTTGvmKtDlB/ZkOkuEt7mbEbmEqOzlVavaZZrDFhgehImb4HH
2EJrdOgcwZzV0ci0HIZWSLCtp8DaQJ3Cv/qwvfYVO4MA7XEnXapPCnaCjosd2PUfl0U7d8PLs6Wz
GUT6re+2vd3M6VtC75R4mkSEtSzCyy0w/PW9LzJsj4u+Q8JizYSo3McgnxKofhfeC/AafLmxJmhu
OKhdZ9LMrl5aRAVdJyXod+B3j/plUfh0NeJz+2Vt8kPcjDQ5RwgVdayRsrX/1Kc+0WyNYGqNc5Fr
59Y+GoDwHzY1ck5YXWUFlmMG06RC+ayUQufyaahnxW2aJd1/r8xxsmTHik9KG6noU6CdMBYfE7CJ
+TA1qCN/4H7j0H10a2fX/KKCX/jFWJFiggdCh1JYFL9JppmSu2Ub69kA5ZGcy+XjwIYtLcR4PqlX
McA8nMgXqbNhpxuWvRQ7TYrCaCGnXi6jIWkNmSBumVeXA2WJXPNkM7Cptq9YBWDWLuWPpUjs4Fnj
egUwqRfjw8jAvf7cKxmNoIlag1p6pVnGQ/S0hCghtnPMzckUC8NKIo4siuxQbWsIqbMS2+lKqLYQ
XrM0Qir5FCJqYVgHkVYU+QZA4YS5pfh8hk5ypYXxGOlhAzCK7cYgUX41whUy1u/4BMJrw0g6H0wH
rCrja14pSm/RtQMQmMoveMJ4ucaPWZOgrMup+Agg6ejWRLA0hsv2tO3EAPmOyVs/SWSrcUpWPS9N
jOlNDPT4k8cqNrbsGS1OI4NqO/hfa5/xEo2WuQagTJYwLC4XAP/3YTqRbOwzwvk0C2bF6hV6FurA
8ZpxkQzSn+Hq834xlvNl7MABC4QF9BHPpeAeCf3Vnajz4+7tU/2f1VNUV67otczg/A+rzYphfRzZ
LgVhgVorLSDc8Z3m1a7Lv4SF8PU8YzmJhGZSX2L6BFexs0Jqg/LgpxWj9nehEHJBjxLgqQw+l7+d
wKWck83ihhkKZtpTd0lGDXGQce4ZoOJNtsdHjlOkP78860+KYzyoZkHnT8h2yjCI7Bquc5EVn/1a
6LQBz+wCcMPSbho9xMdX0UlkcekI3IyrAxqsabStW/nbVbttW+rdOxCBRRhUeSDSOl1+tV2HR5ko
d8/KHu+ttQgIEH/AOuwYJTnWdryczEZvtx9IeAami7aHPkPxQrpfpqR2D5iiwF1cxbnMQiKTpsHb
QSJy9jZMsZpp7rijOwZAmGQMmZKzPe54ZrhfG9T9rMtM9b2ufnBfbWNtpGXMsZCWtZdPHkMj/7Fx
u0tIGXAGl73t/bf5kz5I9Jc02P2fBs8iTGT2ItSMoVkdft+vFx2j03Eb+wthB7fXQ2t0XBtDACxZ
pDrGrUsg9X82UFm3mg7TQqkpjT6OPcCik36Ccoa3zf+MruGl5xjCWF6BQuSNn3DWHwFwCcENbOmn
vK4BypO0LKKhmNbT6u8rrFA96iyIRIvKrdCmn7juAHnzn06JsyDdrACpjotnba/vd2Hm290Mphw5
9qIki27A7ZiEiK8nazLw9kvduwmNFXFfnfp1kquXtn97s6Z+g0zWY57YZu5tR8kbZ1ve7ZXntN+t
q4xB6Uk8KDAyiDve0OtrTHZ8KKZlg0v82IlYLc/TCTnwjqidyxLL+gnwKdW4m1ZySZiifI84cO+7
s4gYtmE4tyHbwwXnTx1ZF65J0bArBHnAOpTBYpw6OKNjyt9cr2ftmDUABP3Xa8rzT4DmqNOnWjHP
+ocxQNzxRNuSyTydAPPK+xwjkIaa3ewce+QA1ecQSvzF1Nli0t1QXdtD1C5bTvB9p34gfyYEpl0F
0coacf6VOWNbbkaW3URjklWWB+Ea7s9qcZq3kgMaqXP2p36U2iV237Rz3qf0I4NcSwoQXzhfWce4
xwCPZdkI7dqK6hwarMBHTBLjHz2xejJuz1qixzK1ck0bfTM/r1u+EMsmeZRciZsuAOkiuOFrQ4ZX
xnrybRfw4Lk2jT82tUA8QIL/tC/6qJpNsv/GkU0oE0ycUcoD7TMXvbCk+y/Pe+0gyEMHEdrp1gbg
PXhnj8kNqO+HMkeqRCmF9WftKGy26S+THqBn8+LAx7itnzFXo8RD5ZVCC7sP5RJ93qE0u1WGxS1q
alCTY2mEqPAh8Rp4fW7ZR9B9MXeROv3eK0IFqucl4b4TfgBb/8ryrOiVEkdLUzuekZSHmpIq0qiZ
zzpbCVKW3vyOpUGH+G+EkoTPPQUpOIZ1JPkDDYA3a+KETbk1Wd+epzMRxXK7KUPfPYJO3QPNusAy
w98C4GOMt4AkoKmeTHqxsl7hpDZBFBXRMdekii2SfSbtA9dhrjogieEBT/sD2qbT6+M6cB34H4nr
Ur+6Y5JM3/bmbUsjuPxGbLYSVoRNn9bhBswIqevcH1Vdw/3nzGIihiL22wQ4QpQU8+t+stGC9AgC
xuCc+61UDfBUcDSK8kBaBaWsRnJz5XmmHt1HVu8+4XlDH1ZUCeokTCWv+euThZOlBFcasLwYfPCO
7gQjjj+anoHvkVb/y/hLNOECsnWKL2ZsfteTImGmWCiLa9khObimv5aOfEoXMzEHMy2IJtMdbwWS
wHQp/j+2YqvqIMfPGHe5h9q391JYNvQKGZ1icOKccG9uyN94istjEFwn5OMPJVHaylJGXnW+oRQZ
pjMIISOpEdt1ZcHzj5cPjdCTN4HG9SYG3ptg7aZBUqW0M/8M+/u4FibrobsN2n4VEfOXLPVuucCs
r9p460YyBkuza5+xAwJaQeaUXf8tbRat+YkAtIUGm5iNurJgVBo+ZY21NHfwjVKPOFM9lDiG5x3p
K7TM0vHzyFPeFrYv1cKJSNzMgpkVx8ySSH/rE3I2NKsMb1C+fG44EbRpBJ7uCmVkqkkY70uoJPu3
1HdXnivYjZ/rOrQ/jf1iP7vmAHE2HfyBLeJovc0zcvLzvsX/C3OOSd+kSAhyQ4quEaaitDsz5tNq
2KgwyQBPI1VAFDd1131Wo5BhsRSgWqtYfpBd8sq33husQCcgRZ5O+mndhe0yHTy1RM08rPWrvjJg
Ktmio0vcjCinQu4/50JMV84dcXXNtL87A9r6Xl04wsKS7cX4H+qx3BvtAVhOM/7saaCBFHwgmjb9
u9wTR6BnXTDWv4WESADA0IRMI+kXLtms7LAUYvX3Oych68GiiRkf2W7bJmEG6oPAxmvTU0hdu4gL
sdyQCCXnKLYAubVh6zxZTvn6cTZxMajLHq0KcBrMvFiofgj5oNENNSkkQvBURlx1k0ZYwwCFpQtU
bcdMhC6isUZtcWBntzHrNIgi1tGDxrDI2buCXNz5wFTLVJ0GdACyVtyuY6pmPjDr5RudiTC402PV
PJFefZmpJ1J6yEzArtOPRjQaqkDvmGdhCF7xkORqru56tpw7FoDO9C6b8zNkwqnrIfkYJkYUIdGp
kminNz8xErZb1AY8XgBodvTovPVNdeeEbFTni0PdBp6SqorfgqRZN80KRghEd+VdtCttf9Ah2zC/
fgEJm2RaL2PpR2mIkbKt2ObJmGnDhyzrogw5VCkVolzMMkj31+WEqV30X7RG5vUEHbzoQcS7RfnN
79o5DUyonKsfR7b9kquT1YueJKZyjQmgjv8NlWVbp6+hd+rjuOfB/k5nOOPi959DOvq78Iq2gI7M
/Iq+N7KcU8r9QY41cufsnVtLNzZmJnDQwhQoDtcZat4C+VDdneBX3lMPhjRbyqFPAAeOIbUM9bxj
Izp6Qj81T+fwapniqRymesgngioFTDMNtsMvQihwx2ObF8vtUGVber5UfQ8v+gMXOeSJo7VPEGOO
9WEX6rMOd3IA43Lq53TqNFeqc3wv0mcU8Goo6opXoXVRjjhysgq630C7Z3M66i9fUMXq2vYEx3M4
9BmnIG4n5AYX5liVBLHGz/4rK7tQdpl7obX03VkdopOx4VV2SHkgYK+bQK85Hu6M3WL2A6ClxmBQ
JxnoLfgxKf64LgTjLwgk8C5+c540riskH/+6D1Sq4lPmp7hSc53LRPN3u4OR5odhhh96g6QGCSSd
3Qu6iu1C+wFawKBRD2f2f06jw9OLpjTEq2pKVSkMQKzXnL25frbtJ9j7qYtk370UqETwTgiZD09n
t+gPyGitKMbWGAtkOeKuY2h4RRWVZZLlJ253gqQhEaHC3FmDwIoY52WYeqLoQU8NR40MuirU0gE4
3QNL0FnNyPfW0s0iGA+nUPQ8wqtAdxMY/AfGxoi13zOGxrnQ3Uh8xUp7cxzOFoyCza+IaaQA6Sib
j18KNaMRv4vGe3C7f5flaQVopSY1A/DHrEVGNH/bc+6P+HoEvyxYY3pwF2+73upi/uY26pm9B0ci
FuxCLhUI4G1FiaJx0TBLiYW2dShYrvLWMVqJuqzhkK7jime8pfmMZqOi89Y52cXu1S8Yop6NKcnl
ZlU0zN+ArRcHyMP1U/EW9sixKMEGTmm0O+PCMSZzkuAiJLvnVRX9ujoYAAtyX5AR+C27TpB6cEUf
6bMCW5AGdDG2a0yJVcGq0ZW3GCs64Er5l5Y3cYlLtKMW+m2V2cxmhGNJwWLYSI44lUpYiaOu6DYH
vr9Rv2S20Jgz8qu9D6ri33rIWcwgInB/uNyzF2y7KM6C03Lb3lcl93/C0lKNR40Yn7E7QdDMwkWA
TajS6f+IMtu6esAi67zBmmdQklW54jRP7iVMc+a+6iYNg4v4wZlf2gZM/v15aPKKbmW/LRDtHdaM
VXK0QhsDHMbTwGmoeM96myQLSneaph4nhNr41acP5l1JYwnZDpX8O4GQtgrtiGBiaKT64BqIjgGr
+yV0hXiLkdYdfA/J63CQ7LGthRfbG2wvpLsekNoNMk6slVdGFcVlH1KtDjaHLHr+yVfIM1yX65Nm
dKq3MVGo+1odqhQkcnCVnFQcQjxZuvu5toc4pArUBiULaigyvEDbO9aUUyGS41F21FRPsBEIGxLc
nJjZqUGRCeOQZc0jCPQ/vodA9YuSS86qw2XU2cpfhFRauiFzLXbO2U7O6sijnw1CXLwVen0WcxVA
jjCaY/i24pJsuG+yU0PhYlzikHnNpDOJn4s6H3hvh5VYQfJzRPeFFMFJEjr6ARt5RQfn+MhZ5TKI
+TuLMA0nLjwXMYigr9l5U983r1dEgY/MEtT9dT9n+1DjHgAhBNUtWSrQJ4JQUdxQRwCJtLmLcKk6
NHqDuyA3a1bC99YAnlDKJ1rIB8XUWjKGX5SiGc3y05Hkp1Ix5C9Cz2r8o8dR9d/2S0Ki/hatjDlf
O5xonC0eJ3hLVXBtYMd5sfcr/HILvO2hMcYd7+WcjVS5V93YV3BQfHquG4ylg/is6mMJtmzG7nnO
Mko6r2PNwkMsexAfpMCNz/41yEzwF/M1Klo/iS9meINgY426REhCC0Kq2WZuJQQtn0c8y+qq75us
LINFCW4ObjprrzuR/KlBe1rpZ3CC9shgs6K5XTRc1+0thO6T1Th4+U8ftyzkdZg8MVSIHPUGYLBH
SBD70YU3pYbO3GSP/zL0f0rtdt9uZfdPX58c5bIyWGEtyLoJ1LzKNWG9GyOWw7XCTgBoGSNCDH0i
4HEJ6ChGMCeb7A4nMdt6Akg5rP0epUmFGec5+lLUiMJrjOw3ERtnher9FPRJwNlmuXkwtrJoZSd7
c1BLN1OD0kRDCJRMl+Uo5RmDP+CCpxihPL87XVaOntOCVX/JfRHhrdLQBOZCL8VsfNOmTLS3KX+S
yLom3BeEXbftvKOvTqL1s+D7as4/5GHfjwF617PPMdHF91G6vFVuFG4sPtA1MZeu3fgl6xdtSwjO
qfsQqpDN2nu0aI2cC9iKDUarPrDHEF2hULVWFtfiHqEciwILpQU0MUhz3czbnAkI7tVljjccD31J
jpL0fjc4mS5NnDiVWGru9r9fkPQoYpr/eHaXNFi8iA/H9I31SM1l5j1bdrnCe4TVR17MrFT6obLI
2V/vc/nVq/TG1nIvL9j2eIH2WFh88U6rhjO5ngAibmc2YJvDIIe6iJP75/ZMYZ8b5E3GcNioudKi
CKmdYpa5hyWH5UAzQdpR+P65p+qKxpeD27Gj7a/MvIkBSsQMWoPkdoupctTb+g955wB5Lkxjxx5t
sG+Hqo3Y8bhS5LwUe8aLgeE3uxaP2tr3X61guYOi03jzpwni9HVrb5/G6CKsEwJFXvEkXMYppbsX
z6bCny2tBtxxvupxTam3CYuPvLuf7xBtUqLgEpzzCczHQ/ZLLgjAVVrF9LJun1HbedGOFts8nS3b
Oj4EqsdLnAtLiMp9lhG7+2ttITJeg6Tz+mniiVAviLBR0xSg0C5T1G7hA5ABHbt1AelufHdS9iF7
jbJNV09+R58PNwq926KSR6moRS0vqQKb52AX4pkeeZ/4NpFzFBvkl2dugHf8u2iBj1eLGeG6p36B
JiGwxYTdklFfrWrD6RQTMLOXHsatHMzm8uD0FH0yNeyEk/rJ5fFJp0glsxfKFRL3qB5rThXxox1N
AjuKJlXwdIgrjw3vJgTj3X2ucHDEcZ5560rmItPbS8Urqfzho9yvtS09eGUhlOjuw7aKKUZgFPMw
gcjPjgOObmjgDRsWGYgb3MbxETZS+ULRpZOw5MJKCMQexy5HLCd/LVwf6OzRtajynsOyY7hF1XAu
gfkws1cNpmuFvGxgWuXvKx2wMQiky4tKymi9S61SQkF9wN4/ZnEF4KxPsd3izW/w/3BAK6h98CRQ
VvKamXfWA8JzFL35xu/GKopECd4iHS15jBuWZrEZYuKk0rpry1BnAlQyu0h50t2ZYCmOYr3dHYFE
jmrVtC6B2Tgb4FXVJnlMxc0mvDCD8TrYiYjC800oqiOYWj58duwYqgznv1xD7mkV79ktj5k213Ff
99Mk3KJs9BR2ff2kq0zmEjiuPHh4PBCH/8tB1pYR6dVUS1j9jWtfNqkmCEXPpY6X00dond51P2dN
74OhhRq/0O3etn0FiRT99fk6MCrY/YQSSheUbBIGGaoJo3VK9tSE7EXTYZb0LE0mfjH8+253g/qi
qm4mCm2JY9e+f9EuWG6SfDV/vSuYMGC02fwNiXkJKI/936Tkcwa17lUOpmy0BaefOgMZPlPCCZXO
8EgQR4ftMA7bs/rVnkiSuk61zOuNt3agPaQ+pBN2+T7loVJSjZryYnZhwEh0raEHkCxxrCVCI03m
o4jtLSlccBlShSeDWXyGjjgVvGjL8Ic5P2X6gNfgK/8oQam0phfGM04ZM/pny+VRjqTB1v0bznmy
dvw7f/4QJ1MwK5mDfQEptEWmD0pX4uIeRJ9JlfFrLGTl95RdcsW4p5sagOzJ6wmWaHf7hBVIQ9c4
g18qtSB313U5ESXUavHkpR1nguZANYPlqbHmS43fKw83goYo/krdFvKRxhD6dNftk+GN8dgrrIMa
vzhJonS682qajbAsC/OjGvvlL2nG5zEk38kI6UQc/kf7/LmO8HJjvphZRbPSjCjiBLV+3vyXqaJU
nsR54zpDc+CvIZKPS5uIM9q9k8+tAFnlBhDSJGzOeR44Q5OXqncu/Xo++STxEfxPc1vYrr/mFhL8
oQGZCxoNEamK5TN21IBEpdMyO5pAv7OULLq0C6V66PZ4lbWDhSgB5fm8FX0ZaIiOIPem4uwu5/4C
lxGWqKx9s5kpIpuvzhXWJv+NjrNTFY9/YqE+vRMoGOD9S+Rxgocn2bA5J8vzp2KigADKu5WpnA76
xh7VkUGxnaSds+joXeVzX0gExei9dXXycN6YxLslIqdrYo+31c3Jf8WrrZkuW4GrIfwJtAiv/tRX
SZE/XvWCRYy5su/LQ1al6ENjq7VBSV6SKdIz5Faszzey/i6tLdc4npIevjR8sysverOYXsmZqTbF
4OA747TQ8AeagYoUe0klXXDfi7p9YHMxYVy0aoV4Fkharzy6FJMzfsG0p/JqV//givi2Zx+Lbhyl
65XQQHI+j36jBIPlDoi73uRPnzbrVGV/sImqGhJm9pgDZp6w8Ve+o6Yyo0R0cWDRzgfoczkMDYK7
dBOU8vPkgoN+yXppSdJn+BsBXSaUszbE8+88IU5nnlvaS5hcJl4YPsec7blWrY93yVhYzXVHCpWa
907fIdXBqDRnJdRyhuCQAx2F37nC/95CVDbRdhfHR8nynJnZM9TEdzfnLk9X6SgYI5IAXPqxSSeD
c6bKJLjSs71C5DOGBcGpkgfQNWD9Zakn4VM09JU9pKU6eUAuhyaVolOw35Z4VGUCQOc5bdn99JL8
Vpl7KUojFDXPJHerCBiXNP8PvwjQVOv9BHeyAwenqqJgD2T/+JnguX9KtukORRxaBl6U8nZM0PkU
I2ZDRFSzG9bvlXidCSytvW4kV82fks8ykl5TvLw4fVvHUHAIpwagUcj0as9fatQMhuVe1wHtFlnR
S70duNwpgYpbnhPqLfxKg2k6XV20qDNT+smTk+LWglVch6cC5THofiXr3O7484HG7dYlsH6gdU0Q
ue++Oyqb0UzAjt91zvffBNXxz0E7j+Oyb+aD/Vmf89tMQAp46Z51OX/GfPUWKUFTzI4Jve4NgVnG
+8WfERYrwzImW8NgdXMZnVDe58kXI3cmzO7dFKGhp2Q37MpHmTA3XpZ1RSkKqRzxHx5SkWTVLK/F
O4Uk9kJI+l7iKHgucquf18r1rQRapiSap8h9j8KfEYJYrCOcz/v9uE/+c5Ydtq7snmYS6vVrWVR5
JqwPs0x0K3q9mlqW44ZnSSGjZR8fa5IIFfNShRn0I/uOfoCnFsCR3Ub/J2sPCKZPAq+kO/xSs3ky
XZ3GQ1VYlXksFKXEPELLY0MDa5l55I8qDpy7lwxC4IDmExYWdlsQvMTi/SRJc6PQZjSPiu1z7wNe
yptpsZD2bb6JcADtdmisuBOI4JkwjRtUs7W7GLZBExyrJRWiBz6QKg1AmAc1Bu8tO8EJUhbBtxJw
YibHJIDrSRwQ7brfq7PKgCTkVqL6E8JqNGaNvfBX6gsz5uiibi9wxkLEszpUI9oTbCDbOa1koLBj
N8QCJDfVPVMwDgdm0Gf4/1+QrH19FuFlUkazvOqPApHEW92lin9+kevfztj0liyyq+i8aQvX87PL
LZNPgQTrXEzCgC0Wrrf4b47PTHKOQlmIq7MwC/IGAi0uM3Hb7/Y0BoaM1OtZNHYKo8wl90/U6VHY
0JWXvNr/ByevceHw2eNtUJZN45ISodR74RgPlF1w1eVFufetV8IpQBVRpXkdToAgO9O9CO8zBhGr
UV+LwFiF/28w50BGb3ZwDVNoOIB6Glqi6peXg+mlvL0VmiJp0lsQAG6Qak79WeYM0fw/PxQR477G
cTJkW+oTd2e6BlUBlAF6f+cpeCu2PbnqBe78m6DRx/m5YJXscAcI03jqq4hU4jli6bT6ga4Bboly
gLAEB4g4WLCHsNfFv1LdhhI2dWbMXlmc7/6zuBdcDp3M83gu1Qu4QTTVULzwfMvJiwO5lIcARXxR
ZfAEHI7UNx6ExztFzvoFewDex2a1HkenO9idP0cWRBKhTBEeURHtxM0Derh77/EuqT0TMBTqzzwm
esuwttDgHvNE1wTyPFg2rLVYJfvph9fGxLoAcydHur8BANnWqOjh3NIY0Bz6YJNrB2ZHydyXSj12
OrTrjUGrhJCCvYbM4fShT0vQ3FzHfUT4cA17Xa/jVO5KECZ1N+BOk/5zenlDmydLGn/bqtDU5Mqm
zJYHaAT1XgX+ee0vzqaxgtrvmuQir3B2970vpw5AX5bRt5ul+yI0AOBQ5OUPnWCk+wYJz56Ybrrx
g5syNwOlhv7g5AEhmN4SoP8B3RT0CUTP1gzpSAJAGqFJI+1qDqOshvKQCwgq7tNfNFyD+vQkrVXL
uDrcFM/nJO8QO1UR5QiDrcwqOCF2kzyANiA9IRNIiXNMCVRnCqnzLIT5OWLQeT+fOcGa5BM+1ffw
Os9mcFH8fzH8pCdTcuwfWYWQ/Ge9UsxWB6kMP7DXoDgOBpgvpk4REO++SaQaj6G6wTQTwInP1zAF
FQur661L/+G4K1O/Uat84z2DtGaKeBnvBWStJLUm2LPtiGT3DA9CMY9UdEwwtapgZMfru6N21E+Q
lJmzYRVqCsl6RG8mcH76XPereRaThtjbyQN1knX3jtLiLE7700BhVfOFdZPuGSv1hC+m32Kayvy9
t35UoNz/24n2aFG2KA1N55kyAx7JvWWMZ3R9jpMk54dMEly5RTIfA7FX9l9mxf/LHkcp9Xj5Aaqh
2MVVsVG/3+pIDQ8d/9HLVBNORIc1eCZLiDHLyHcL6N6VM/syBCLXbccO59jMNl7q/MZLtxY3bdT3
cKf88iAO+Z6zJuUE4cyr+3rpuPjqmnBHxYkBIJ5KTndSf2R5i6kkEIcY408QTf/qA3HeQNEVTLgY
2suKKczWA13hq4VI7j2hFqQPcDLsYmD7AwESAGpUURC/wcNIPrUGqqCjpMyPFVkOmGYhzcFNLyAM
7MJWE/jKrtLD75ePsGVgia0j6e3dXFq0nCqjK7xqTsqi3+jSdofB90VY3auPIqAvXG5tS5pEl5b1
F31nzZ5P+Cu40N+EBjYGJQVQFMlzCyVDwF7rCIsxq04J70Uc7HxcCvq+xy7QoGOdLApoPI9Y8f8S
tO916oquppTsE2niaP+EMovTbyLKMNibctHZjR+COTSaIgPUXKPRiUt3o0ASNhTcIuvbHidGVpxG
f7TCBUZF3l7FtRwAP4C6oQDAeIdgYAYxeOACh7+sTZZffHgQeMVzdeD58V2wg86IN45gTh4pF25S
61YrGvgVj75qscugARJXr14XonCqN7cDEFvThKtJ/Any48rSEvS975btC6d1lBv+WLkkyoRo20rJ
LOMjA+QqlYVPGW+eHlRW73N1GyoK0x8G+74ZpTOoC0frEQQozC72m13EQnjycFRufN70aiaEUJ8J
yvo642V06D72srlwMGf540xUpCDCeNZIWtqgVNmkRylm8gEV/BZ9wJOVp9Vh0fygr/nd6RLzYRhR
PrG3J2tL2usG/41uzfls1e5dBixNhU7IA7TEPjUZUkJO0dOzktFytU0VwOVQSp2w6etmzzVWo4c4
4Dwp6YfB1CCFzN/B1cnqDZw46sDppq4qODoj5fBDKShAEyLo+x8LUSrMjUetyT/fS11FtfBmx5Rn
dix/TcYjM5BJw1UZ4Bzbs6KXjkzqh8/c6Be1FBpRnyuFC3uOgESknbtiuFIsqk6eg2571b4CLsLL
LOLtDhzY09wsXI0fJ0idpkKKtJdDHr1b+xocjoQNhle3g8OZhRC3OEBsfwXBHpQBeuF/jEEWfqNw
SJej3V5ShWe5DIhMr4q7kagIv3O86vXU4Ly6HEWt3YwdzVGX6qMIKFSVFDtZoSm7e7v4dh7RS2BE
rc2UCnaA6Oryt9Tv9SQJC6S2exFUk6OV0HXYy+L39GpnJmRPyANDU7qfpRR8wz4XTcF1vsAFk7Vq
C9Q6VslEoIIF5jMUzxKckYLPwP0gxJtZIfewho5S/fMhQ7nkdT2fsTiIkUWyD2Kv1g6aUPhpdcv0
bmbRi5c+JhKofymXEASlZzBVmEZg6ykBYO9TK1BCMVwZBRrmTRDq1Rvdl8nrtWStCVYVdq7N5it1
LzQWmW66KT6yz0wf7XVBpgoXW9tlXQ0oP1mhftbpiQe9HH269MkQ5CooeeHX120j51RvOkdOQTBb
h3xykLny0W9rlZAjpIoVLuyimmwRKArikFttEL6zBHUOuhFlh5ytN+Y4XDVwbsS+pFU/tMEKSbqz
zNLFyVlRB2eR251+TVvs8ZvdlDk7BGhZRrR9TzsuzYVhjR4Zdqj/kR0UJbKp6iNWL9TCi97J/OTl
zaIoWOGh6WvIDqUy7PDC0c4SWXLFy1ZzSNhn9iqUdZocmgylaEjKfW83I6D6QSpvcyJJ6a/+eqHa
eolSlDgiY8A40c2w4rw+ZAq8nvhhshKQdJaDx5nhWuqSpN69jWHRYNXMS5ZUBMA+HCsM0EUtmBx5
wkU8KmiJj0znMY3OJqshluAqqLAzJ3TJF+K0TsnOMLARI9/PbP3ZqM7wzNdrS012+L8pJUlXXUJP
Fd/YdYVUH1kVlwTzUUTVVGl79eGeobXPBhn+MTctpN4zZ/0IMF162/BgNu3jyf5HUNxsEFBKXvNv
o2crQdxEx5AAq+xBdFfp7zpNyEjIQ4hz/eXA/PbWfFvVyp+IYSRaOaxm4g+3HFw8axsZLI5Y3oLR
WuXbic1SIJZvpFqI0JpoTg62s+3SEz1fwUkNn7volFA272caD43TQuwikCpYpL9um+Lz+L9RaecI
+hiudN56gQFJ7I59+6tY8PlTTR9ejgGGS4M6TP7oCmZ3+jsUfjD8Al8fff2rXp802LD8VYEo28b0
GDnH/fncxgz4sr6qzWtFDlFR7LsLwKCXtEHpS0PV7F5hBwFtz1rXfRuTh4TzJqGmN59ssRHzl46R
fEj8RUQBPiIV8corq8Q+YhGa4C21dBlc5JoH+2Z2S1ZqqWyDBjhnBiuK6A73bB3OieZ/otkA5g9j
TO2bxVcLnDRTPsckMHEvJlS8Denxztgu1fa3VsXcFXpBMKLV22rzhu4EDkT7kyR8gRCRKSXLFmp3
uQvdycsEWVe69TCL+vpYncObGGGIDG1KCtdBlOsar0IZx5CERpzbIW0J+XY4DbXsT+FXzKS8RVPa
rxH/iyxjMVW5JESQpY74Z8FLJF6+88LXhJI7h05CnI99K80w7GPhb+uYuY/23w7tr6kiQldeFxmP
OwRDvKk59QiNNJp/RTnjG6a6k07cCvlEp0VxA9xIlQelCtrIUVKImIvj/2nk70rD50PEiLqQQh4C
NHozpbCt5dv+BwcfHn1U8LJqUJgOkyMxaQGTmHyqpNyqVaPtw4D8qAn/WHj0rXn1Z8dRvt0mw9az
Ohjzwlvv4On8gWhJyUPopGwIQLcuyJySvbKy8cIcFSAf7oSYQ5W0uK9mXyhb0F47CTS/p/JhqZhT
hL6PmOUEyOcYTsA5nwgKu1lmW6PZCELacHAWQ6YnCS46PNtjTWZOU8E4urj1NTbSRtkl8hvDmzds
P3bON055e/HAxnfQeQ14rAshylDWf5SUNasgl0DN1TapM+A1c+CIj7zBIhOUpOeb5gxve79QSCXY
SEEgGB2W90xM/obtIWmumtPgVQ4gqfdvuDnX0YfLt+FlkMbReeJE7l6ic372XRtWIbk/xd2vyT2I
BfaFMt+m59o5HP5svlPSN3UcN/4enJ3G93+7ERNIey9Pwi8RLocJfuRLQDym0xy3mdQFNFZxFbai
QkuKL+W+3J5dt/rJUFpF2vilXcC7X/myLEOYNtcKssXNX2Iqxy5DVTgRdCKVfo7tWhZzsJi2Fhoa
A30ND5d8nZ9scx5W4GyJB0L1ZXRWrPo2Dtf+CcGDbX/gfkYpTo2OZDSWwgJl6ixX8QjBCbJpswvK
lnW6M8h9y/ovsG0ITsiryBSzEhnItTshwHZMI+RE78mka0+FcmUUVwE+gfkFnXr1+N3lcZKrOaRI
yr9wogqr3qNF1PBvVtLhbRGyS/vZcG4PY7g8RO+AJj7Kx07rD1C5hqqB+67W63C/EGhXTTIHhrnS
tb88dQ0XVQNqBftnRLOFtYrv1xM11Dj/Kei7gW0JFElfnzfFCC15yBnJCCrvUrUozxLmFiY06qOo
7K3pPtAVSbqpjXZwoLGK0/ze5RJp6Isq2SB33a8t2I1ArbJYdqF9ZrrebRxUkXfKXZ5pxZoqn3M0
xfSc9ANekWHbk4fhn7boSmgVRTlYwA+WfJQvOy/DpbXrMpUy7h3qpgYtgXCAsmXLe11lHIEYQi+0
XMBYCfiIOmRwis+YJ7t/tCAhZoC12ckhNS0lDKxEGlfPj/5vscqe5/LiN7XACmmBVn5dZHAUzXr1
BmaYjfc0sOrirlSlfNxbPIW9D47uTxPNp4g/GQlC5odim5ZEBWHMdAwgpNUG+0UhOlg7kJI3djAH
kDw8l5bjrw3fDs5L9RdsxKb10dppKW2n3rJQHenpwT1B50br4yf4qjo7AipTnj4LZ69Fi7YBCvIf
SKAwmTYHmEmh8+zeRDDPAckEB/UmZvRy7oqmj9FC7AabuTcyVfkvZVOC5mZUlfiCJdnjM/e/mpVn
hRkekeSsXOoxJ4qaRSl6RQohzx2WuHjnZiAQxwmMRONbrTaDlQLMyF7VUZIv74eGdllprtqJRYt6
pdvWBA8r8gXf0Ve1iH8CauMlUXNJc1+TQbIAPtKwPT9f8wiDUkLNN8II0Q+5ibqSGspUzEGXHz5W
hGco3e+QMJvgQ80auDdQEKXXyWbv7pOIwQCPatP0btUPLL8VgeSYVKCbyVjfxTf3JEivyLNZSHd3
SzGoaAQd+ncVIn0JfXyKz5rcWVtggoIYq/30a7Febu7RyS6w19pH7Y76eOg6s1QCPr8JQP75kXxH
sncIs4mP2f7AgZ/t7m6WUAqT+AIDHxQq3SS9MUpOz7cJgZI5UsCIhf7Rm7HmAA9WAWim7LFkvMrr
cKMFOkvnbeycnMkN2gNButuH2ssMbyLCYXJ0qEy5wbpvl+KalwL1tFLWDm1l6DsAmPCAqq5qwz+m
oGSzY4bFQ1ehcNswXSuNR8+jtGIwr3QZouuPd5NvoRp5mPmj8PtujWvGggiq9yEJN18Za5zsqU7k
CK7TsI5pQ7icz8B6RpBXHtqT61yyBY0/kQmw0RDzXs40gWJPzAaMtTI02jNnRy3VKoUY9kZFJ5d4
YliPcaGV+ay4Gwi9OETKvzNNd2agUPxP4wRaEFf8n/Mf+RNMWJGOV0xxEdbEiz4gq8W1aTAza66o
T+mOvxEyDh7UxaiFjQAClAJuCcLkaoTzmJ6PxZrdiG6cQTREegaJOGfVaj+nmQSSEJzeoVZW6mi3
m8dP2bF6hjy6i5qKVgoLGMQKqP0qf8wakMCuz4ky/szWKmNrzCYI/TOZNnR9CRhQB1jKfKMsqvKN
RYxASZOPQHzwli9YKgxq5LUA4It6xeLDc5k24HLOLOGm4tqxGC9SHSsDphte1qzBZI3BKvoEtC+o
zshei4dcE8UR5spismCb2uPUQlU6sHfq6piFKBwcHT1FY4iDCg/SDB7/lXUieVpXnpMhnxepI40b
plc5fSu7Yxg2B+c2mgdVPh/bVbdkBlCN6UITnASAHQmKajNIdaIy4yxAacXSzOU4dfX79TdU0V3q
qg9n3f1gwTklB681sjpCAIpx5V8QCqfiSe0gAjX6OWJNlNLDSI32CS4oSsOF/aI6SryIpUK6quFg
W89nTA6gEkIkuaiU2ge0BsDr4EXmMY4YwsN8rAEApruRKxc9TLjJOhjzj3vuuLd3HBX8C6X02boY
hugo08HCzcihXX5TtDKYF5+QqS2EFKT5vzPXpbUsMcTHd+czKyLzSsBKMUcOy4Zgx4KBayQoHPKM
H0aCJe1rhAD5pIlDSHfGMSOwYNVhOzwgnpn0vEwUA7uHukoOJtGCWpTtDX/EBnJSWPMzbUmwIdXL
dI4ky2GYwW15KN8ZIAAOsW3FTqCrhFqJAWEEqqDps5UHH1LexVE9msG910LYNCkLsn3nrSn5XWbQ
dbZqnY19y8n9dce8tgziTBhg62lNjLYnjTs+g5ImTetPQ055MkUTrcjtoZ0bKHPp8oGPRi4Fv7R1
A9hhi6GUxFp9zPyrJM6cOKhNIT28DJsUEFAEA44qVxNSd28ajqm4SqVGD7Fm1oEDg7UHQkRaqH/w
STX5ZaEsTB/QGR1hjlhLERypUH9w3o5195J18gg92edsxf8TKZA1rCbGeN8JvF1rBih474W4PsFd
drfr5DROAJd4g7dYUlhlfoEqL3FqNLBN3FDuNekeYCutLlWcQpO7C9ll5kKwZPqDGbc0j8DmQs/l
ErT1C+YXSRvSKpuz4IrBwq3pmQ53aLG2RCE5AY03ihfw4JQ7BfTYO/vT4mfTMkXmPBFHmS35Q5rH
5Y4QXVvAzxk1dYMuwcz5fB9XtOe6d6nC4VNKo7uaxfjkIOlhgrJwnvPNw6dEok3n5CGiNBImpu9K
ZnmNM3Qb5BcnG1mYQvZoVtMlZbC4ax+BbEZxwJ8O8B2cG2kCvGGoeXj8JHwGwnhOiFVYaF2Peylx
rbJ8av/HQdw3/jcWM2otteIWuSAV3uC1DzINgbDwlFX+49G7TvUmWqsJMxdPjDzUpezMZZM6EfO0
yUa240sRPDKMepV0Zop8uCEqJNcERs+08hrlfcodYRRMGHGo9KcouNWEwYRzANfWN8TozLM9C1qX
qKqkIdy1gT54xJxltY8L1H4pRGFvB4Zxag34r61FfqpU9A0914kVqd+qVLyAOD7HaXhsfdVpEkDp
kC1ycTMM/BYalNoLwQFQTw/kTwOM5ZizJq2ik/2lD5SV44p9xVaMjPMtOJ3JWitUp7KoM45m6Ppk
nZlMpEq4qkj8CgfpIWbBymMjVntI8B7hBmcatGBOMB3B1sGLF/sSVubJXWrZLXnK3ajDyzhr2yPW
F5F0hAG9ZGng0e4DZzTMR9G4n+AF9lfmMtG0xkky2+Id1rH+8b5Ir+u3VvqDIjhimaxkJpTc+Lsv
GWJsCi7n5qKI7zaOPbJP9LnHmZOad99KtkT9TujrmIoGIuTd4K6+HEh9C7Pz70BQOuPnXhH55wPW
aSMxenzFtOv+Ob7s5Ps3mg7bZ7I7yhdHXah+RXD6zv91oDd2k8QjJNQvSjNQUjNeT/HNKlfZrABD
JsHRWy3ENHC4FMD/jfM3wEn5XWvFMKOiucB2rnuLmlHV1T+EXJ3ill76gNVHpak4B6IQai86YKy2
b5oJjQRvx691nbfEDi7zcl0mq35cl/3GSlEd/Tn0aZXPkJMhs5c9q71603K5WWgxSFEiOLsAD6HH
jlzPaTm7LxdAoiOVn9G5qecUMKSSq4t/XSpP38tlSIYX3vvFJIuQgVwwmSgF7wGgbR8Vfz6nZ/1S
XYIc7ZAzWrv+iwUntjOh1SfSnBFWmj4MWAI+qsI9IHznTvxIccHLywSIoeESXJsGPcWIICmEVupa
45mX3PjH9dXfHLqQAZn/0/ZMPOgiCRwWcL+C6mK012IgPc4FW0+LsQfDpvMiUisV+HHHW//aeBQy
/NlG9JyXJsEUQ+z+B1HB3rLzCx/h6vIJ2B63rgeGFAoenrUwwEbFqx8yOeWAid0c5+6gV1F5U2+L
Y3Zn66q0EdLngP/650Zmdz0bkfhqIiXWH1D3+Y7eFSLiTJkPqW/85HL9HRvK5MptoJmwlqquoFbF
TsXtiHLNAVefnSKRXeXHz/gfNNqJ/bX8NdTcPBnccH8StTzAAwJw87cS44VV8RGMRHRId9L55aT7
7Z3PFFkxGi6ceHm1ypvlsCpO9CPw1K7bap4c7QeAfXXdW0hjFK3+jvI1jQF2suahkiZZNUcuLcHa
cdEQgKX2+q9L4aacoJgsiu4i/7lrM4pgs3tW6L/KRGX9wRBKBxtFCJTme1AgieQoJVeqldLVOPhn
8Gs1VGSH4KtGlFfW2/MfR9exalimysgURe4vjOC1uqyNk4dWW0lC7dQ9+U4pR2yqbtO/bBjhGu/6
dnfGNIb9opR85oFzfxPxnYHf7ixscUr5caSOwyYtpkvTF2n9qn/0cUPCqf7U8+BFqqMpx5QOYE6a
iUvfGlOFOtjYIIAJkcaz4sJFjdRw6+qMr1hfuuPXeHpsyYSVvvwXujx2QsygrWi/BfzxhwPLJVZf
K0i3RlVWAAMyB3PQvs7CTsr9TGk6BodU5BKrpJsM8NxAs2UFs3btm2u6pnS4xKyeXpEUpkFeL17k
SfsmDI2teEhhE0m0XUBoRq1LhNDWYS6CWXNqR+mo8hqIly4vQiSxIRZORgnpEDqT9yKrNxXgcq5Y
KejecFgsA+UCxXL6GUHowaWn/YKokMUkJpjLCvRW2QOwfWBQm3MRqGlJ6RSA7xgHxot4xuK+migX
wE0qXGpPna46yIE4+B5vKQX76MUg9CxAlZgAR68r9t4VVdxAneNzarmacVAgorFMIAE6mGuQmkQn
F5wyhVpIwtUHKck2JbVK5c3zKTULwI7VI6HGvvFfopa/7Cj4RLrWW5gn+WNX+2f1XkZrlrdrqJ44
vjxpi7NHJQTJp6wTlRfQJ4o7IMOehlMvWGQovOapPepq8Qnx8TOElQ+4Igt3mC37EIe1/f9EyY3H
lwlcTmIm1AVo3qbyvjbkDxJD+w5DkHqyrX1vjScx42Vj1Gyfc2LGwu10L95wkvk3cimVI6i2cI5+
3E77juPk3Makh4MUWYgaBg3xKhKuPyxvLcw9ivntrBtzs1cVKp7dPbTu6fwpIGnXDKyKHfkNnRBl
bMmRNk3XmFoDO7EORUBlhVQQa2NaAQEjabuvPBxpBc8chnegpBx8xa9ztL0+FAIZdzHSiZpiVyov
ghv7gHi0BGn84g8wdemj4m1Z4/PaZV+07AATP6j95Urh7BxdGqMR6q7H4sErfdLDskT/P2zzzvjt
9PJyUfrhEmL6iDsNrpgL3x3A/wc6q5jG7lJIsrQjjNSofzOIlp5HBd13SmHVhynacbO5qqaAVKNB
rEPGdtWemAMLUVAzgNxffC9BoPtdvAoLTDIC7DGO2FbTUKClWa6f1nfjvJUdf0oDPBovXMxgl9ML
G5qWPQD+0KgkdJoEtm9QBEgIaUJiq3NTFBTL0PaiXMqLW4ICesd26CRiAz40GMquq6Fi5H5Rovus
boDK9/VmPokRRaDGTV9II4bNeJ+Boix3gYz7Ad6iI03dMgCgn9pvJJzLVnp2xNkghTu2jp26uk53
oUUE9mq583CEpSxwciN0hCGMVBpmYio/Mu8alNTxj00IOLZFqJ5peYZiRY5PPDkbUXTpuofwo4tp
FY3VwGE2ujx4LnZDnOQemWVouAx72igaVPo/FSM3rJukTy0WJZnHlfI0l/xRwSCnNRnSmkahm3PJ
KrSzesIfx48QP/rZcPyAVe9ey+VXSQXCP17g7KS79dbBwesqvgXbPSXgwKiFQpIQyTYcel1HeYHf
77NC/isyHAfz/dB1ijCZJ3lZXlOlLUM2IeCqLjr5IgperjmuIHZUxVLEQkos7gLjYMZigtI5f9r8
4QIatM6s2AYCuxhX/56xZITuVJ+yPKvjLwDH0csFBpq9KahT4gdAe6KLzeppkA0Q6T3VHamPNeME
k8eaOJPvVn6oAJOf8gNhrctWQ5PuI5KVNaIoaZ0XUduAQb0rtyuGjQM5UtIBUtwp6LN07eolHmGi
PyG/zsShwrY0M0s5C6SjFtiEHNenp6j5VrEChJY2Il7YtIXtvwSG69ES+V5uklnNRWzhLA0k9bRb
sNX4FG10UIqjpjtqdLyifXZIuqi6AOQCuFjS8L3qZCmOJeVGSiGSM2U6jFwzspnPJUX3TDFniv82
0OaJiMd0jH7IHnfyg8v/AsQVJcEoiesMq8myLcUm/Z748Fmzg40KUvxTs319uxJrQRFlcu+BQxI5
a3cCdvNhMMOp6LPkhizlKLg6jo5rll0oNaiXt1MgPbiE4BbjvYpXYUWKsNLith1NCBbWmaniDbmt
aEIXLUOsnyG3tZ5eHKYj7FGwEx/fmf+Gf4DG47M1P32XtUaQmpOSw8TjpiOMZUdjYiFkjxHCZ1b6
brBM7IwukJAgesv6FReKm8g+1lX/g3PTObzp1aSGE3K+sLeGRuZE9GLZQotCzNXf68aAmLjlSpp3
eAjxB5NnV6UZMc3Al8muRGu0KPBls/A7AAv8A7nVuQjTFdTNm7ppZr6Yfj88JUS8BPcQARJI3gp7
2Pv6bI69hdg6okcZKq+tSVu9zOsIxY41OFayNrMIOz+LV0m4rY4B21UYGytxz5nqybInZG4Tlrm+
I1d+W6XSA/M15H1hdDEuxPftq+e1VwmMNwWbgr59wHZSZT910gkN73KAAE8nWVALFtxdQWHdfSy1
khXcjOYMScfA0Th7YSV1x9dg434450pLeMOmQ+uolMZIqaW3Gx2LUtEL/lfs3aZpF6J/4JzugoLO
mn5ClPcg1Hbidk4/fh3F5uXXcdVnOcYogOwxEtzHFdwPX92FjO2U03uTZteMx4gyKEgj0c7JXOaF
Pwng/T95TRsgmMHWqqAEO5IFIYzqV/a97rqCVdzIx4h0Jf0zPzqfi9eYT96Dmqi67NSfvFL/flHw
DGkRH3kyQxGiOIgmW5IsNcpU0PdGjQUERL+9bbc0o+JoTy5H0H0TzSJD9e31Ujn3k7u5NloZAf3E
2wmit+526Uf2gdhDrvme062Tgs01KeryPjwT7SEsV/SepAW//OAs42ZAbAdnNLJLX1iecmFkLMGa
CVzVc59FJxxV9gEN+73Q6wbSDg66TNL85LYtdRG9CtX7TVRNy+4qQ1QXmHhiXcIcoOwXgwOZ1kE/
eOUW3nVCbdkkEXhqH1R04xrWCf/914I4cedW79KkgXXIKUSjvi24POWRHUZkf21Jv4c90sIS2iPs
OOuoTASV+eHaKYm8hFCA9eyF//L37px1iS3B7GmGr2TP4Uxtnm0f2eQaYonkwdUgd/5tem21kq2A
w1c8g79p5jgSc2tCXfpD8Q+lLUq8L6yyli85RiD1XytEGBMu40lcrvzj4NqZT3GaKj96eQNOpdLI
f+AaB6Sd5lPbCNMdLA7b7FHBWRGrVmkcBpvptpPNcjE6BtxFAWDKcJMRIZ2f7GSOpbiy1jtxjB8g
PYTHi5MyXYHD1qaLQHSllp4O8Y9PM7remftIYkMF2P0lRjAW3p7cZEU+TvS3oWeSVHxqlU8VKkdT
YGknnLIiq3uzjMwM7t+jDOi//luTY7oyhWuUP2bxKPp+8I2mc4b+apBxkcq36KYGWsh9f4An+4gz
RVunDnMtrPM6YIYMBqFsdFLVyhLJdZVX9/ijXl825r8CSsbQJF7mXm6V9tqfhGxqdLtlS8W/0Lbd
Wt6kNAD171W/r1tC8Sc0BvX/mEP36vz47wwQyxNN/DjK4pWjezbwffORu59Gtvddb+YrDvJPvfUz
0czf4ZFzcDxNW/jpWn2IHLyUwZ01TT6r2faQtbAGhPqlMGUO0anJ5PcaHa7b+W6ZSEoIRS3DtgT+
OxPrU/TnvxCiAceHZvdJSzrDHC5/aAdDXKKZ9HpnWFUb3Qca/C3+nSe6VfLWz9r6pi/SxWZ/+RkK
ncCB+hByV802HfSWRnN+A4en5BvYPz0ln9BccJbCGGv4S4SVhcGlHwZM4yt57U/XiHa29QxkBysv
h1hwO7M+3JhdEXaK9uLCx0sIJ97WSRuguZwmBPhJaL7hGltvgYQKudmYKttPKmFbCkH+R3u/Klwv
L+EIhxVO/m8SnGWf5OQzEh4fC0bc063CU66Py+UM5O4WrroPhQ8NKMVX7DwEzYyofR9Ribo8Bk4f
Cxx5NybftW/kEOcylIMo1jHks1+OMoA7TIqJB9kWR179Qjpj3fCxomx/EzlEp+WqosxLmdSoXb+c
BmXXhXXLnjFU15bQ3+qQpVisLVhyc9RlQBEatlD1ZmdXa/aixpNAoyntS7FIXX8jeOK30EanS535
umrVbQiKytMwUmZjpph8IJn8LGL4IXSQLP3PUwfE9Cxmdf64/ogpbCAvmwek/6dXH5xNNFQXvDMk
cwYhAlekwdhTvXc0Dlg8+WL2kBFYFGzGO9Jero+NP6hC+/yGa8bstMQkf+lY2ASVIak378E9gbh1
JVOerDuiB+6xNjVha3JTp/R/UyXj3HlwHhBosvJsrxFriewGxqCiXjrKp1q6unlaksHJqfo3nv+g
7EWnkrvPoNYC4T7ZEnBFXR5P7czvYpBWfJAO+l+NKubp4zgWpk5hO9d4K7MC8EK6vgzpdcDCguHR
iObF3tAWXfBWKIVq2QGlpPwN4iOQb0mjE93AHaGQf5DkOYy3AOyQkHKmMmz7gMgLdtfW+9B7Y+EG
D9q0KtZ2+dc+CDdyepnTF8bjEY4d2zlAaUXKJ9OZM5amDtj7sRMPUibKpon0nSsy5ztGZ3EZePuB
HQBpQc/Ogx3X99V36XvOd2nBcdDD3DTNqs+Frzxoua7Md0kQO0iQO5Se7hUHcsxjKlfyKHrdozVb
oHgjPd8gWOZ3YzK8uZeQRYVZQhoNFtLmnzgg0vRmSlwoLT44nHd1WfDiYhCRVCF/MBueP3fyHqoW
AZlm06PVv2eYEmAMdVrZoT5ZtMZpqTVm0SamnDn2sEctWjZOivNQGhIUDaNjM9oiFKFrs4SKASmN
iI3gzgjd4RxKIJKdIiCys8PRsPESle4HkiVkYbUyMzxBs6LjO6SUXQAXlXUVYDJzl2TNVD5Dw9tT
Odg+csFcwbEaGw692VfyNmXP+iUWx6GmiG4njCJ9ND5YkwpcruqmwTiUO3q4+Ry4n+nEXcmazRcU
S0yCYfgwuSklf33YIh5zwRW9DCBDy7Eu7JIAGKKZxoAW3Dhcu0IEyhYhvhARDd4fmLR3tDWe0Qfh
mN+rxrx7Fu9Zl0iTi3M16UhDuxsZKM0JqpsnQ1jC7gthdD4xgerOwnTEBc6RtM+2703CWh1MWuh9
91htsjiNe0V7dVHMymdRga+yGYTUs09gxFpHG/B96d6UGIMDmzSEu9rX+HXGoEAVwE8/hVc5Tm94
RA+5i3FTzKEPbiMRHZSzcWZ0LRlv9l/uFBdAuODQKWodEJhQBXMn9eSuE1NUxyw160yt5C7Vfwsc
DAZ6Uaw0W3UC8W7X/qCXVRLXHO9YwPk17fcdwJouuCIewMGOwhdHyXbYuNExW5ERCwtiWndMqJ8T
PRnFWnPEbEWgvMLwl+LD+kEnPvhvn5gwd7qYOm3W2SH6gKELc2Mc1Ei2i/vpUeKAURREVswRCEV8
dJn6YiT+9tw9pTf5/2EdCCbgampg3Db1Kxb2tz6EYQFkoRGOr4u6kRPERusFHp4nnCu+TK1dZVA0
Q5mUHzYLW1G5wSaUj0If8M94p2COfsJZwBTwvOyo6rk+n79hC6dTHkJTAv8IahAthNUXTkldWo8V
9gB8qfX7Pdvy1MZaS/5BlAq2Lcr7fkUv4jPKrnTrr9BI3LupvVQXx1Z1/RTkDHrQ5FqpZOItM/WP
ew8yZ/M7L8zMB6H1HzsykUFMTr8vdjJ4+vjXVeXemGuLT+z6YgSDS+J9pQC+w++mKfoOsKoBrVWB
f+WR9xP1a0brxAXs07JvUdLzD6Gz3TuqTQ4tm7+695U+LuIgjem+9uMiInec9TD/rvzU7Uw6hgLf
1ns43rb0mZJYfr92mQask6iHMWiaPaM1GBQ0Wg6DzvHEybd0KRtQ5QFqMAps0lBSrKhrUen5olpH
W4DDDAIwHUaTn/uxkEGsPlogaJ3IPwFVVmAdGo+Qp10geHhQRAhH2fYpb23CnH8/6BCietc5SsQl
JFH6eBX16UqiB8+z6qO9ol/eZQPxUBufg/81ONCmCwsXgkkZ3QHnixteBfP016C1D89pmUldeJVG
xyrPvlWSNB1YQ6HKnCDoqmexehYEIKoByJvic3c5322aJPfbAo6SyUnPDp7dJeQlujxonM8uvjbK
Yh2BLEqO3usk+Cdt6q7yKXXxuGStH4MgdJO1BiQq7++hFnzmZUnaqeui6HAbFCbQMJB+sF26aKsW
/tkFlU6FMCzLpAX6vhS9x7ZBqghnmT0IAvS8JAnEfZgRzfpPBekuyx8UvXFktqFKAT0va7DQBx4c
sgUIJz4uwbdTgV4UjPQ8lKGVYW/oO35Aw5rXt675g/YA9C+4Ik1WJecSuc9ILoQd0QyMLIPPrWWp
pNkkHbcKuavzErLlqd8r4nyTQLxyIBzSIavJh7d83naPnsI/dSmMxtDxy2hz44JP9Q2M+6AKwKw0
4fu1nGRjq5mI6kCde73DDasgtvulT2K6CwlpkogJhTo3kWwFzE+xCR8CQLzUsa2BGPQl5YbpYS5i
OzWfig2zhgFAGgG/DFMcKYhDgLqxens1Wiv2gx4lusy6owqN4uKCoRUuTYkWi1DTjroyXPqD515x
4hFwuubJte0qRBrlwZm04NPSc4zZC+m0b8tLunK6chOTbpC3DVa9m6/yPYP5gXSmGkqJXo4i/eNO
j90F4YWnLiCedm0806wj1+eR2vZrWnbpIfs8pWWAhSkLFlfkca2OhDR3CxdNiRW/dPe/6oIzYn32
7dCiaRHyvHT9Iti/k8EqXlgQ+AjRNneHwryBu7q8lNrJ6fDBRo8TTT6FnIwcDRtkpspMFvImGhyR
ksThXv5ss+AW8h1Bm3/ZPi5q1s6tcjMO7rglt75/3VGL91NvMZCiSCLqSt35fn3RGrVlLb4M4WaF
CpmkZdh9fJ3GuVwl3oMNqWtIGQQHwtjVna1E133EYyY7uWmZtWvBPVkEG9Jm0YnYjMsAqg10t6Aw
LPWU53ZH7NYaZWebgj5lweiSDGvVPRTm1L2ndj2ffFL9Oe+PvEYtLACX6tHQoBFFY/1MRASnZLzV
gOs3igKPSBnBv+7GhTOfr+QAAISG6LwzIRxEnwRZIVVJQOzBZwpdDe1nlgwpvkUngtFpPQESizQu
f1iew80k+tqKfhbcX0Y5hnfUwYpMQWoNpMtu7O3iHGOA2WUTvQOFmZFYxpQAlGHva5X5C8sGTODV
blyeb82tKYMH9X2cTqbD1ykJaY5EDFzkbPLzSCfsvUkAeGX3DSYYvLktLHMwzHV3NBuyGp+3B9Qj
S+QYLN0BLEo3QTVdyCJjc1g0LHFQzgHpE19uFbnsme4tRBFRB0ycpdfz6KpXbsUfx6JVXiqy+NA6
1Q6J/PTBlAk0I6x7e0ARg66rXTZph8Ml9VDvdFlQLgtXKm9nZzab0FyPmxBz/KGSZjYZebWo+qmC
x/rzi8NkcuDC3zvN5bs03uEV0V973FzoBcn/XwfRPWzY6nMSXv8NUfJ2+HXGKEiCW17R00XRuuGf
S26T5HkoBPoLbmicMudPrsu2y1N3EDDfjaIdhD8lOQYWWlCungfnptHWHPUapO11+8n/8IScFGdS
Bw7KPNjerHgXDy4cZ0Fgub7zYCJMRsbKnc3zhHWv7RmQKfw8mRSq/AXpczLmO/bwF8OIPyny2Xf8
NASyo1Fwhf2ZdMq/Ty/fljSxd5p9/1lTkIvOg1SeJTipfvbVNUzRROMK+lYgtYEFOavwLaO3JkLj
652Px6Kl2h64zwy1jthfUcAo+K03RO/TFb5RgbZLmXRS6XEKXDXSMJf1YBDpu/QN9qKfb3fTw5sf
wqLYWsHGSA3dJTcrl2gGboKGddXNF+4rWQ1tuuQYiLQ14M/A8f0e7voeaJJ974pGDJPCGk8u1P4a
H0Karsviyve4IvPWOPq11hsm0geJBzbuCmhDZMpBV6qAA8Jf3Rb+ZOfh/eb8E9KoPraxyQuG9fjq
KehKdqKDabCRq/JvzlIe02/0P/gUNBjwBG4U1ns69xRFG3Y7yQE3lC2I3nRQ0GNfZKc4tGSH6eld
xT81Kk+vsPwHCQ1KllCsqYy5+VpCN/BZr20RdUc3fo7ZL+xl7n1mGkhgle6J0YyJn3VvILtRoQ7k
b2SKYJ3X1xbmqMRg4h3t9M8OZ3wV+KQNI+FhnRClUHK7mStjaBESKFVnQRyKNgl/oXn6oBO0e+CT
M1eew9nUhLqBLElptZBfgkf64zP5Nk36R8HXEE/RYllDfc8MJuroBEI1CiHpGphhy5FuImcVS/7n
J1EqHLdCJ+bZ3Mb+geh1Kyr9Iqrw7h26eb109Jk1GGeF8HFPzMnz/IETS/3JYiEEswcC7Ia1xKYW
guM5pcXyZFShfFioO/82lyo7rNoXWlND7OsSovgbKm7qRzLyaoMPyAOYbaZA2raqxTuF/y7cUTos
QYamTPyQB7J4FU9G9RrhAqNnbwVHroq6BdUlxXGjbP1+HRSTAFgjOerpwDTe3oi/aPGyfitZF/V+
bRc7mQDOGeI6UaF1W+gzcBiLS+PbEBP4xRnv31lCivLfx/bUsd+80zBd1xeUaQ4Tv08fyXizp0Ue
ymYJh8rPzQtzVh36uSJy6hehJSJTh7kzGW+j/PXQhE40qmGq+a6LLsK1DaLGlMPDu6qlr18f2w3U
okcbo2l/dkZj56mU8X5hAWKfpzGMTZDbUTFtnrD1Grxd8IX1zgQdEjBGUz9fVz17IYY5vNgvNldj
vwJYv4X3JoPzJRpmptMjc6Ma8UJSdZHJOcOlMAmtvUgzu4UM67+HUtrHwpGm/fkQWzHUCULEvw4C
DDqVKewpcrzdJC6qUfYFRyg2D/wvNBgTOnQ9XFtiEZEu482ALltyfARHK4HcUWaBksPyOl7s/7uC
80FiBp2nny05aOSTdtpj4+BtppN+qtXhjPi8CBUwZv3v7AsAUPrjdq2i0ie70Cc7Eahrs7a+JcEd
M8RWRj89puOX7/B+hkMnh5+miMp/TmbHB4gsl+Iih0/+i2lHtyADLdzxQE0+mwvZSikLbjbXUAtQ
OCkEU//1zpG2xDmuiJjWfPiWCa8x3/jGsehRFkBjNB3Hi7PBT78wAqVR72x0EmyseSVR+BGBP43P
RoDzpJ5yANRZubrExZfWIazQwKrCEpcdZtfoDrtLTRC3NIp5j023JWYzyTgc4H/RyFrLEeBKzDGt
rZjbaeBeeIeVX3LwcwBnT9H0jFXsJrNmQWnoVvQA4E+zdkiEFGEmj0TxNzh2GwRq4ze5jY33FpEX
E9UVJfRmfJCdMU4qQq8K3PdvcG0gfPXxIgx7nsTLnKhPBwmJnaT33So78Jl1FAnMa2Mk/YkO9181
K1ERLnUNm3tdTVEzyEVTgcqfGt+AM0sOwbf/6A9S6CMUO011azKNxt2uXSXQuZtfgTdZuhBuxS3n
GVWM++qrNVyNnWRpx3139iEDo33ERK6xtFHRUnk3UVl7cQqspFmJDIumfosY/0euWDhtTj5tYDFE
x9CoO+Y5eYa8aVxJ8eU9Jz6kGGcwGxT0Uv/yL1G7ST5xbQ86T3g3gb1rH+8bhb+pzo1m7pk19gA0
CUHbD4R4aZK+FeqhVmu6Doc7RTDkdKWyI+zVBvsump5T0wL2kGL5LN9kKbw3Ke5QN0lv+aOyLkVs
swyKcWnFYfS3eRIpr6xPMhTkmhqUZ8dnt4RhqppFIVIKaVadFFXkA6R+6mBFDGl9GO2eGEw+aDjC
T3czzfVIO/0NVmMYpLONxaei1BLSzIgi+1I00WJTwySUtuo/CwDN+fKNpT8oO0NJadDXevUuawXX
G/WTcYpKdRQx7CSjU4VO6Z3shCtW7laFT6S/mjnsTT+gk6Tk0PHYKypHklXVcHcD/cQk5VwtKHru
v6/BUqmvJ5SfWkO6yMWFAJPHBgUk4OVJRqrxDZbP84YrwIVzC0fe73mh808gCsDo9mgNJ5RcDCKp
vwjg/B+etVuNPo11msGrKjsH5bl2SFFA50I19DoLjbTAbnqUFbBXa9b399nlrIDnEeZlSoJXe2Ve
UD77Fw0+DSLS9l/sQTZWyU8l1ozsMnqciK0wIo/NcpunVfny9/E26RCB3L+r9jXnxfeW3jlU+dZ/
zfsn4WWIbn3BaoO/fyHkKWULsaLQpDgyadAqBWjiu1SryyTmadz5eZwww82IPr6Q73ZLzT+h3Z2x
8wos6aZlVUZ9AuHJRvACT6klyB6KxDhy7plbk7qhuGpSA66QPVVuvclU8Lyn5tlwkv+FBKWpV+5h
mPigBtrSE+bnFwLQ1Ot0xqoZv+kY/yoVUmp0IKFOUyycOBx8kwnVBi+0NaCq81o6l4dL7UvgHw5Y
03trVdVCC08A8pdDTFoXu5vEhB/6OC+GHdl4+okv+LIkrotRmbKIDXwLNLi7ReDoWVMK+8XRNYfk
sCYrE9uLchcx/pIalOFHBDmwL0m/DwaQ7XSO2PmfaGbRu4ebM7Xw3BzHRYqwtFKe/ZWVMV5iDKkz
FPvGX/oxeX4x85anoDYo53hjQilZqazcrCt70i0c8y4SRBTyOUnGvfLbrmCfHULWc2osmXRdeDRw
ucH22PBdDP0i6gNPALsI2XM/VDV0h8k3cchZLoupIRoeGmRtxNJq9tIG3xm410wPsQyyc4wsAmuz
A9YcCjk3sN8CFQdFWFGgcj7UW9256Vkz9tmX8C9Qhzjj4RI1tfsAxScMgzLW5qAEaek0RkURW78Z
F1Lfq6/UsUFQrhlDHWaXL0hpdiD63JbL+P+AAvqVuEkmWap3TtF406Lw9AjkPM80Hwvs8Jjr3A/z
H3/JURU/Bt6LAdRSYW86sCa8LVecwj2DCDwok8oGjT0z3i86jAdzqQZ7lozRRnDRLnG7KJe/QNR4
23R5aJqxUMuOrAODALiqZi/IU5PGQzgS7+fAQysbtgrurBewuFOq4pRtsyC7Pe2eYdHRfc1UV3d5
aah9wOhhU2Xubct8JNnut00Zsnc+x9RTIU082pv85mwegdRB/xIvZPOKlqhp6OofTJvv+ozdCJ83
x4xunpj3PPcoAQ3g2a7VdkkMG6JsyvWwP98IQeTQDxWUmg06AJN9mdn3mRZUwsiSH4AKpTWgsY5/
6yavzHBUCBowYbf7474lOVsa8eJFMPRQfy+Wso8Q0ozgJhTtiDW3q1VI2Rzr0/CXeG79OcVWlnks
BxCFqNwcSebmmUZxme7L59AFx3PuG2/FsJ4stFfMM9cYenW6ZLtVerqtb5R3ydn15hJZ+Ox2elMP
xsTYk9hjulVEhO4a9FA1MMNjPd9xVpz4fOeqS06/TnykYf034DgZHCdtTivEEKhj6sv1PwzhWu1U
gtnKpWy9N3fMYHnLkk3XqmURGX536/9gati7lKt271X2mwD+TPNjmCnp+hIWvkiP/Jtg3Y3yCl3v
4KlTBZkeKy1Qxv1l9tOu7h++aYIPAJgtqVXuyGwCcbi4+P8+w3LxzM+h4h809ED+VaYvg5BuQjyX
RwyVixODwrc+qwQ7q8Vu/4UMZjboFwzl8J6brxkElqZDOCD9xK3saHmJyBCYhlMKwvUCINTgZfer
iDelTV02FelMCN/ytXhgoBqw6k5HtH/YbGhKh2hZ5NeQfGJ24+NvjCYnsxw5Ard6TlGUqObodI07
QfqfRg6HtDVXFGXeKSuhgBfFTi+n/8suKY2zd5SmqRIh2bs2b6k2ZqZ1OuuZk0czsfkWaCbxkO3D
E/TPfT71ZA9xanOfs7jIJmbql0WczgVTbHY+tddilZxNtq6D/L76ByCnhxJVIUqg8fEdbELosN0m
Z2HiSIvEAk6iUkNuwHESvLaBWSDu+WSjYf18ZrAzeBJ9aXJ0w05dwjtVN0aA7vMVvNdUmzw0KJyG
EfRjV5Z+4vxbfmu8c9R148e8HD0tXvZNoRadeYsknxT9Y5oKVsWL8TVFJAmCQeQQN5URYlueBwT+
szeCFL8bdKRqkdNOKKaTquGTs6NnXM/VpG2P6uCST5JMJeoPrlbPxT8VnqunXfON2vHDaMwdwvVk
W5lClU8HaADmhQd7eIgSNVP7BcfqJRh0Guu48OyU1Fe1aANPOntjjlFHAPg2FNJNH8cv9VkQgWhO
JXv307vETAXew/q4mG0GHl5lxhkg/wPjPr5p2LIYuqAmBgVi908AL2gFXh1/nZI1CCyGqKT+9O0D
Mg9sMc1E6qFYCPxmvUGLMbd7OjaUjJxxo1AMi6fIe9R93B/LBfV81r3vgTJapfX6AYyLd/5a8xk5
R5V0F9aOcka0OB2KFQOp5FrYxLyA78UwCliUk/RYSF1URhEpHCZKvRk4SOIwOqVm6sg4xeXps5b8
hlJ7Ee6DB9dQ88Z3fV4XXHOh3TrJgzKiYSwVrKoQEXRivDG2HNe4bIuG3o4fzYFanKiU6ERQFvB2
aEP01yUUd/zYJZ94hOaJOnQ1zTRMwTktLih9B4knfXnC05B90ixp3syvPbn0/F4NLZGT8ywzUS9N
dynvMIwjjemzRVdsg5piurYGE3c+s/hBSYLuKF6ZEFTqpo7kyeM64Agxb6c8lEVQSMo3HNYplHxv
tjRU6qXNRm7tEa1Vw/QrrLAnviomdh8j3zicgLWyjQAO3+THZhbQ/iHPPgD2bkz5rAFrAzG+hCv8
6VWWff4E7ni5kVw/JBAikhqNXEfGZF8RdavvntIjLh0hqqvQwLQbR8woKwkO1UvVhtoeKVpxC07P
xs23oJ1atrnuO6WpsvsZ7BRGXoa2dwdZI0toWleBfr+lEG8Ps/iGbBF1KKaw1NsRxBhnIBQF8off
MMzSQBxSZl1o1urMEWmkqvn9zcVNGdEaJGfgbDLZaIlFdVE88sQ9kN9WHbkc+vbPGKWduzoNhRMe
gduLhLdJR5xUQzfSYkFEvgsSRk4O08IrghLW9+7OufiXNuW7h2/s0zS6uBBUII1vQdUTnjDx88fz
fY5tQ3ihEX9/3TDuOodfGx13EvB9Y9bhS2MezgD+LDnfndFpC/5cpkUsHV3fdhNQcQUHw7PyP3SO
NRG4/+NLk0+6RlUjM+z3CdAhb+ga8AJq0d01YZxbJITyaaGmRG4HH3vO9DGAP8thZMxFJnfMpLWV
9kjsxZ37okOPXsekAACfD0Zdk2IZMLiqvGwxdr6P81Z0uQwFBJlyKxeLzmxtyJVYgFrLoizOmqFi
jMGLlgdrtmmUIJxwp8ZETNF0bK8w8lSDRxVYhUZb9tm2nuy9ZJKGvfp1LJm+vh6R3jNVTpZqMbDW
H9xvQRPK4P5EI34wZNnDhKLiPNSdlZb8mI4dvZImLbCuwMXxy4vvNoJxVioqCyqne/oythFC/BW4
L5ViWJcqPnGoIFvHvB75/DYZ1NcdSV1HO+SQQ5IbWeXBq3bInNR8ixArJ9vjso6/aQIE4koZn/Ok
cq3ydFXprlMFz2kOQlhfdb6V0qD+NjI+fmKwM3JuJb8RsTpp9GTC6yiIMxYhK+yZG8fnZgwoxQcM
mBA2ODeKN+mbmbtryKdpdyFtpTj14P/wfB//syucK66bQ7ovaKoTNzK99j+SIQsQs+vOPzWJUMpQ
L7ODwMHMe1bKfcps9SY/u8jK46H97X6Tx9Ps+yjtqET9OtiGfgi177nB9Uc7mcrYxBPHLnDNM8T0
Wlu2Qc/5Qum3Hc4evqKCy+NmzRg/5Z7jeQXSDXLYaRtLcId+56pk3GCNeY5UD8MLwfHGmJO7BuEg
HK6yfvvxSH2jd+/v80jHcv9wrOVwQpMEX/nFVImjuj9dIUB+Lt4gIjgIwQDW5fOSKKXGwsQOiZLu
RNkfKTbDwKceE+pVf+YRX9y1CSy9PYNSZvmNSH8k6g9MzrdGxCmB94PabBs7qjM7IV03hdEduUB1
4xF+XdXaUeTSLLrKX39CFiDycmpHFjhspPNgnRUpG8OzpFGx2YCkAEZw+LkQdK3AvlhDWUyhorpH
yi5sdWVcg/X9Uev7DP3eppXIZ6hpplLKCgap5FD8Fhi4wIgqdtBO5xOZO+GJ7aA/mGOZzX3NQZR9
rdMBexxBDJgXVCg+0eoiNsBE0bBiVGmq9Anoe+jJc+6hcTvkleb//SEbtx8lQQFd98Zk+rrYbr2q
B8dElqZPBlGHUGalL+QIcrwuhslIaKggOZTlHk8xPpOfMhOjqVnGzXce7kSh2ft9/xV532aCKSyY
lcmSG25vGRbDmVfQNv20YCIaUklk4dm7Gg0Xs5VTQk5d3kzxSm6fXs2rd2or8fDjttd8Ric/VQN0
EgOv8+CxDjxbTrO+YiC70qkGIeWBXu6pBVRYS7Otr4mW1Cvaror25o1LTXHL8HGVTqwzUhzfkhOU
wQ6qqcmp2O1kZ9AApTExNnKXM8hxbg8JNZEQvV7PtzJR+aX1iYSTdDE1ujc8++i5OXkdS7ZsiX2c
NkSeu5tf8sE79ydI3qBYr6jhUPTZc85vj6HMHdaoAvdx1ntnSn4TCFxfQNN/2mCYUj5Pny39SzcI
8aqL2EIHN6pOpftetvKGcaxNaczz2ImjN7hZkjImPerjzfFcaUIwr27ivqOCQflTOP9zP2gd7YIR
S7mQ3FtwJYvJy1EpuMgRhbSE8604d2UjAAxWv8d547OyDC1+CEdLzIZNMAtc7f7ob+3FQ5I+FTdn
t+/Vvbb+y6udyrzMB4CgnrskRpP7F32SUC60dJeVnIci7xGmXglM9+DJ47Sn04iSXEJdL/tO5/eP
qPNdAeNteK0H6arqgNkzlvp21OPhhnx4w9m5mAtbwZJ/hHmqxQP9mfr1xRnPznyiqLFw6fN1oDa/
68TXENPYQZAEuXbdm165gxaWKjT2DywaeIU/dbZyMhpIeuimPnAd1aGSeOnQpGjHFp9UhDYlocX/
faqDlYokqvj4k/Gg3eSERjWjgsS2mRBably8GnZ7Cs2w6GIUm4FO6FH3GvO0RKwt4VCW2U1qfuYF
gLANeplq0Qof6UTGxxePUwnO5KtZx2KbQ7xgNoEnmcwxWwKLpRbaBeZfwurkcsabjZoAQTLMSKFM
eyM8tbPU7x1rkAFnSOCbK2AmGqCNW5GhvW2JVmYDPhpNdw8ZBgIy37YugoxE1lAShp23TZ2EmJNo
MO38e4UEVrkxU6x71o+J1OI3UFvP53f5bajIBp6m9giOvGKeIf+ETwUfjeHQdwfBdlNQSdhaHT++
e/tS1Fxy4OlDucUwxT/Z1AVpZ2oDZq11ID+ugQdTIESsgiN+sbDl6Dnb+O9oK+dqOJJ7IvbrGUZz
q0rnn+mvifxQZOIRl1oGPcorL4qPYS+1/DuPDmgL9SEOpODq0ZN3nIMWJANYVy6837kvUFcYzZ4i
jCkkSU8tCtaXbNlPNdgXPPve+6eUMCCf0Ey5Mo4BUzaqAOTD8QV/oYvr1xy53+UGkH+JZa9UkiGR
xXYVXSRblVr6LMJYdnSdsYCdQ+uUV7PdqI5xNCpJNWH6eyUNwx7HPPfipSJ3Pl9oC5bypiDKCvQ0
qBYOhlI4jBqaGyO9B367ughC18HShdDQY04wla72pPYzfnzrYlwiJ5qTIy/YxO/nGE0Zj2Zp8ycJ
lE5ZtRQHaAGEfOLCwuWsYskSw9gDc04iuth4+m//JcfGd2ZgalgXLjhfV7q0fZpy0PT/Hes4vCQf
QQtrZZbYYU1zV2yPgLQJ+YEA9IEi/nst2zzia3y4qxJe3IU/y91JhB1yMYMnzELDo86G1FqhkH7w
GUUg94hoNOo2Tm5kEDvQeoJcPvfaQ/uVXTg2dBEr1spyRPW8O7T/wknbRURPRTS+y8sU56ppf1VH
6b35ad8ppcDEuQCbbnv0fpP/Z4i7pPQ1kNy6FL0yIESeutRSTvk3HTcO244HJ5BdYQ9OvSE80gQa
vnsSNK0a01EXafiF7CfCPeoK7nqIQ1uQwXvUwiXZjE+HClCGdGL/7+uiCF5YP36CdcV4wmp+jkZs
UmAA9CazjkWTb5DyHYCP5ZGWMeQA8iV9pn8WvhKlqyhjJTcS91OYpRhWO6C76kggSZRpJmV1UVcF
WQxLLznCU3B7MVMdAwQrnj48sVmGgmX9ZgZF7Sl3Q+gSlGPsuWBZD06qvcFKcf3+YA8iB17zxOeo
vEWcAj/f2Ygz3w8WwGQny1orWNHZnfnxxhFDT3DtTwAkpg94rnTZDIBNE6kTU/5dVnxVvsAqJ3nM
3s3xtnk+Gky3KByIKp/2gS9+InC2aNKIrouXb6Lqx36u9IgT7DU03XAAeZqApXpO9a0LWCdKtxbl
wP3j2hPe4F4vkaX6V8LM4ewdCWvj1MEWpSt0d+AdxyYoOgJNAKbaal4hZOgPzfD5U2rj29Q8mPyQ
mlGE0Blh35bOwrGOnO4LSWYlgPNZbTTgD+k5q3GZ2H+jKpvQ2crzIQYNHgWsqYZ6Jap1TmjvS6/I
hLuKA2Q0hpK20PTAZUASfLiuWLoRWTxeIe3bRKwDoHu4feD3mywIyqzOxpeYKxZwDoEB3/T9beK/
l956MbPFlxXq1EY3IAa3h1iuiZmfK7xOwgIuCGkKkM5+EH6/Kl2veaifQMh9ZlJ44CsyYNrqbx/T
NTDB5dyVoeSW8sLx2GyuzJOLDgzwZznC6IZ8huZZF+WSZ7//GGxKJsTtX2mPTOuo2CtLVLjq2Wue
1ZTI/iVOny9VQVOl7Buz042Lq7JQxcGDLq6I612F1rdiTlbJRPcu/Dto0Kxq4K5tEEvuJss6cRPG
Xy011li5CKL3nSXAFiUlf1SLW/pATcc+v2Yuc0xLwW0OF2uSH4KkKdhWeR4kTy/3K/EZyQ3JPTDX
TE5Qd+yUdk1V+6wEaJgshHYjc6nMe0Ia9QtHzrkdkN+nxz5fCsgYCwVsYayV613ESL+SqElxPs+T
/vMHqh7VaqPdNen/fshznjY0rSTz7+542QGn/7duQZ3GnZZRQXwO5GsxnGv0ctTt+3CSAbvadJCY
wQwOqfWnT7pxe08wIG/jJGkN2CRDLFZtUJWXSicLKHXWAMwYo0S8PeB8dN3xDfSpquXN6S7JFu9S
2OPJEAB7H9WIRjMLQ2CACheSGFPwvoEAtfaMX213MyYDgnK4BKsIdh6IitlWYesBwxVyucjHqjK7
h28ywx2/APnuCF3M7jsIO+fg+a/RjN/0Ge2qtYCGe11iEWdYGHYkJFed6UCT3NvxXhT62+sGOmmg
EP2mDTAFWod4DQnTqNZ5NXHSYJ1dxpDmI0ebbK9lRvbNARsv1nodMEAkRLXEqLNjaeSNmAoIgrZd
xhIE4GYnMSCNcVdezM0gSkBOBKmA6P4KaNATB/vWYRABsWmWzp0wIbCdetEgiVRMsQeyAguxLfsg
wMx04nKKa5yGpylLCn7FqycUCxncmvl1A71U5OxqPiXkQoVcbi0JMmzidZI/uo1iTMRyr6Zn5CfU
lwB+rCxMI3jQkz9edQz2HUYyhOwRq9VzXKiB0wOfOCAxvPBBdS/jChMccvfbXCYk/MOcFFteosf7
dNUokrdo9cSeOXwvvufLfMaeOBJFwJMPDDyhjl+0k4FMz1GofSTAeC7DINp8XS0YDYz4/aK/26Z8
YmGa5tWIid8/D9Iv4feC+j8zHdTLdcjvblqVoNZ2e3WU/S6eQnRe95q7c+a+qwPEZY3Cyz9OPfIe
JAh2Y2GO17wtiX2KFSQWLqWQjNCqIgpRYDXSWN4rSHaw2HK6e05WsxN/3k1/xUOvYNiT3cYUDjrf
/u7Ycf1TGW+8RJHC1NK6P1WAKq+hX8EPahCmwbQkVIEvGMfigrdcjvLYiAvlEF0yujFoq74sWick
GHC03M/zt4E2Ss8xGRUGEluzCnQV5AFMa9KG9Jx8xMqc1kbRl6R2KJf936SQDr/2F7l65eoAiWcJ
s4tLanXLq2cs62IrU3vxwQThCWN8Owi9+7rsLUaqOdaE7L6b18tCUW/Wv2yDkRCCtZM8/pAv2WCh
ZQ6xoc77sSbKDvg+3LArmsg48mTOCwJ7nCTx7M8hRDe4irft3MUkB3j+Nn4Es9CB0GQVdPC3tfWN
fVBhGiJQ688Vb/TVdxqSTULyniIzYNf13dRTWgJWvgztlFY9zs73wzhlC0JGMJCc1UTIIfLnc6wT
GNwrvMMZbBpR+iYduhJfuhwei/hjIvI3k2N8bKG5fL/xqP6RhV6PSdsRb2P6LSd2bRWrzOG5OXo2
DJA8cPhVbWLTBjcwbiL/eMXm5HOcNbuepHJZCmHwJuO/ju1hgebe9MWnGDtYV1lXmT/YwMOepBrB
EezoG0CJR3hCQqe8AqCHTYkmC8CDFjUx1sg+XwZ81YqwzMpcyq/eOuPUjWDRZqHhSgOzIE5EWhOs
6inCyOMSnHYrTZIRJ6f4mn1ZIfGx+gKSCXVpt8PmQsShJSnaoBs1lhy5cGZkD6g/6nSmymSP4wS1
gkXEWb8YBrjU8b859386rHO550MvYr/kLLhDwyR/+HLy6FQOx9pLlpu8A/TGmUOfrLHiBcuqH/8B
xpp6+cMJiFGgrTnQYNANTGgjDkPxLxkoSqW4DFwpRmUZjrZSmav3bZQC08QtFMmCJeiqcjm1yl5a
5ulfuS+J6nXEbC8+yNfJyryNayBew2GRXjU1zw6Z4G0a58c4mS07Jm/GC44D1p6hYZ2dka+Rd8Vw
K42DLd6CU6i6AvqDLCxJ9fW2RKfHJDgMGiAUQhYOjKHdwoT5LDONpucJPxtJ3PJlsp7RmMUXiLfq
uhUD0sPl4bOYFLOBpPiyUej5AqBjtCYInB+4D280Vvje8gQF4ueWe9Vgi5sveMDm3XdJB07+qe+/
npk4Y2BBt+FRO5DP4oQfEYjyDvFzHLhvZE3ixIRP5yvaRNKoVVxCtaLEPzYIxEJB/Ns/K3lSUWkL
6h+Wz9C70mW4NCHH2nPHhtvMguHINfj+WNeLo4XR+frsEyJaiKUSRsFbQqJT3uKLXVfyYmaexmTX
Z+jxx5Y/i9khK6+Jm+9Itc118HFT/mknTkA5k4UD6o3sFJ42BjuxuoCp196OtBfqEUP69P44Sr4y
/Qan61h1KLZxlp9aeK75uT3LxurrSM0uQqnAXUiapEjvYjUEGCQttqsfMZ1gRH4YsgPoxKIcsFph
tetibWlf2jU2PY+FEMK+2IDEh6Gq+02vqexVgRq9BED4P515jGolgEH10MyQ6Q7EAsYXKd9OB3GC
kUvv181Nx2K6GgnIFbbAbStIWyCg49RF9zKZGxqCiBVvPFHrGonxM3EgTEZ+0xoFbQ8p9ofc6ZGQ
b1BVSzGX8vrlAMGulWBf0NQ24tmkG9YoT76Fjz0Nu4Nh5HtafmfBhgtAE72PNXJ2GvW4X4ywpTRW
K2PKAFYWd15OEsHSUpng+NSAOrJ6dr990ORzsQ/z8KOKEnpCkrcoPjK8z37f50/w//ShTbhLmlkt
JPHbPHi/8kgwEIRy+WKJyjYDYuvl+sMwvEqlKNlDKdTOJwDPLW3ov8UA/3M7dph68NZGoxwFI35Q
BliwMRk9H41ZXWDsNh4i+ftyczGtuel0kurj6HYh4vx3kxYqkI3DNmTGzbA9Nut1HBusUmYNQ7l8
0+92188GBz0a0XqBwqH6F6rBpX0R9FAZIGN11Z4LMvwmPMOgqdf4z+VxPlkctnzWP7IZTBsgDsBd
vwjKnaKnjs4Q2aeU7quS0RdLsVrZP6y+JqM1p2PWBNIaZ1m7Ws16UVLc/5cqT+QqsJJwN/1tXJaR
e3bYTsPW9iC/tv3IUIJ0oAQENzoMDoJAesecmlNE16iCas0yF6FSokowd5U3B9NklkrrKe18v2Ux
NvRoO/Q+abnxUIpVx30d27v4TI0PXWrXbr+30XLxGBOqKzB6BVTG1JcXK3PxY3ut9FGGsM6h6fAT
bAp6Fnw+bmgpBR7zfVZh4jbVNaCGR6mm82Tr+rzAAHPsr9ZqPzJvMeVRdXv3mKKGizx7NhTnOZv8
4ZY5bvdozUaypnnZjt7xKE7i6IMQCvVBp6e4+SYSrfbqIDnBmfpF/GgaxNb57bZswGI39ZySDC2v
ytOBqLJAMzpG4HjGcEVn8F0zppCMeiFDiXOSAlzRKQPC9IWRqCfY3orAz2QYvL5cxhSN7+YqCB6y
2oZ5tl/jL/9boN+6r5Vq6mBC2G3whprrmimdETkyTqd+Cn1MA8WmpKczsy91EOFwu5C261QnVqWC
ZheI072uukxQfggFRcEEMuEVT3Ec4ArQ/v6qgDwXcGl11j+CAXrJEoV9KiMjw2QBT3KSZHIv0YB5
4ADdNmnHCu3HrfgCFKuXtlbd+2o94vjjsLAGDEDGcVgJyJgdAHBm77+8xsWmvBt7PG41LGNhEtEw
yc1hzmU/fxmetB1zpqdi5WqDp++x+ovvQV3Ce7GCWDlclR24jLZY7MGzFpa36srMRR4rwGrEF4xL
3hnPDTbdShRlDXPS6Phh16oPiaBNZTJxXyJR6wwD/AMN20Ks07doRz2vmd4WnKrTJ7CFBNhxTM1v
AlYxP2ZrH1jPFEOv0KkR6AgBEOmfOiw+6llX7aLlLJ4kvIsqZU+PYs8ZwxZ1c5lPQQfDdOGGghEd
ReVudk5R+DzaPS2Sau32Hd3fjOikc27/jrxW7jxZVoEs6OcWY8MBmK9biCa0eKDgPCo2byreAduQ
MP1BCyzwMy6buX06X0fnGE3UsH7WmiwIJT0O/tTigUmErig1SOiWPyXtnFs7ePikfA2oB2y/ah9/
hKzI2xaZpxaU9S1xh1lEqX+MPS9RUW+zOPLc5A6SEx6+liToLl8J2m+cznYUQBAteQSs7h5+73om
6Qn/fSvze7Od/J9tkz1Mgl3MrNy5UtuMMcaizLgTACr1Rhx6r7gnNOjy1FOGc0RDOD3UE2DDu7e3
bplZew7Axrq1wqQgfrn/Zq9TCmzsEAc6s/k6B32M56MJnIzm66FKx6dT7ue/BoKNNRBVTyuySKUT
m8nhDF1OYJk5HTfoj6Z5gqesIgBuEtNA7PZAPYmXGmu/xy8YT/A9GkFqQ3f6BsGaLYTAN3AZwmKy
7QVNHhjXcJP3fC/ZrNheEuPQL10ZAfxvE2aIeUDt38jtsLPgouaUUmJ0jy+kOBJQlAkfjB2X9r/L
K3MuuKrIiDQiNSkm71W7ynTldSEHIFfWQRZifpnH9amEI5JO9pcTUQrJXRZqsPYLdt/4eMKz/pm0
mc+zkWUlU/XdXZm3HZlrFWOM1QIohn9wfC7Fvm9pTrkuxvrDevOVQ73XoDE4lXML0vE6ZwUXm/zZ
/uElUeu5XKF6ckMpaiv+mnZvdUvaWH2MBkWhS22k3wdxUs1ELbdYAiuImqVBoEVaQbROMsZ0kLPV
c/zjuH6ur2DR/1ybf01/I1Istx2nRbAX4lu9ZV2zuz3K8fn2pfq+l4mwhNjhC9Mf4HXZE2zId2mZ
rSpA0ZWzfCNV1qzAzDERNqPhYoRxR9fhslCsStwptVPPfdQoRHkjP+zKJRUIzxL+UmXjhfNNbifg
THOALZEReDLCNsXYsgzVIDKcOsLLTZkdchzuZKoJ/jHMITQofYoS6Ad/H65fT7szk7NuRCo3uI+o
PuCzFOlcJOk7A001qf3Sz+M8s3juZiXik62lfKdqJJ6+Pva8VNI5CenlV6I1/66JTTxDenVplOm5
0TFhYRJ3tEwpJ3aUK5qgWWBIUCTspTog6ttsua9eE0prqQ+ijodWk31PRpmSsr1KjCtjh10HuYzR
Rx9D1sni4juV/svhy18wlKJ1W7y7sCfL9h94P6cBYrHz0iyIfVdkwd9sotOEoQkM+W5U6buQa43Z
IUMzX+SJfeDeerOa9W4woIZMSd9Hfe+3b4SGRxrkP/Oxu5JC4yxKpD5NnXPEIwE8tLygWWbhG+YA
teNqp2ZFiGQ4Yw2sce7iubX/yFKES2W003VwkmAuvGPYfZ7N3pG5bA7QGEieDKcVZGLNXILyqpYN
HrKfu/iidwsIypgtH5X4eQu6HR5BhgWXnWVGEqmf8VG73VnythOoEiFE1l4nQKOwRIM/gDhhYLxv
kpp1q/BMniLA7SA1zJpZLB8kLhg5ZtlECbkJmRQq5zDWo4xLdZHQekIs4HUJGg1OnQV9te1mKFiR
BAhL4zjFs0pZ09P6Ydi3wAq2KvdVgsV6u/258VX4wMZSo8djSCtbNuhgeTx+k6/krgpLJpSP3aKP
qTfPUo9shbF7QYIHydsYJO081GflWCoTEuJSLbcTwcImGfmimiaV5rzMT/vsNH/eIFirFq5bpZO2
OLZe7pMzkZTawGDjBnBDbHj8UUfHsv8a8MMRb5YPvOFdX7pTMoPFjcS3VOac2G/0CrH0Sr4Hqq1a
hmuIlQKNPgO+Fk8IIEHE98U+v85JjjhUqed8pnLlxdEGwXA+kruFG0cbjm2OMmhlzhPkyqnBP0Zi
52j8fWYc/j7mHJfRPubDIRBZZz5pwM14MJLAHR3fVV8WtF187QyFEH6g0fAvr2pRGI0R/soYyD21
PG/FXOIMHP82pCT3weXpKDK5Uyw9xobH9BreXnQF0tdnyb2h/FfGmzCZy/9EwIQCEp5z3eXv0fvL
kPfAwMAdzTnvU27DU2U7es1V6sZur/IieS8qlNhllIlwVb4op+yf/HfyiKhnpG3Zmg8iAFzqaYCt
EYELS/yCvFKGq1WHwbhw1wIjB14ALGXmEZZ4HGKaLAHRoVZ25tRAUnUHgNRgoYyCv3WSXYKZyYJc
stLcSRqfVbYnLkBXrZiriagalE8/0D+x4s453xoGgd+Zn5vysdU4IIo2UQiOrWRIlr1Y8nlFUker
m9vVyMYl5H1+RAtGhRl4jLIvuRiEAD/wTAKev3Ehr3cr/GYrFb+Ien0Ntk+rAYX63Ro7Ro6Bx8yf
ptPCzd8khF8yQsUX7e+K5sG0Ns4ne6Cni+XNXyFEIxZkh9K//tO2ThIz7lLlBss+Vo742OXcnk/z
dvmxVbWkcPDAk6g+v68FJIgfkxq5FUerKaa3WQyQWJHx85Mo5qGrpmOQlyyXh4cxgG8jUyRiEnj1
CwEWAVe4p98+fZITNwx0mrMGCjgD2OXWBMhwoHDUhdftuyAgTsmnTQEmwgpEc9JsZgbSw29tCeNK
FlKNGAM49q9w1tNRz6YwVweuza24EwtgWCbUwFb5ohAogD8RseCm+xIm4YnKmlSjedgh8jmEev5y
eQ3pT7AR9lsxUvvuoUAGUye1SvHgwHi45hmT4+6IFG3lxLt+dO7qeMWAfb2WGtkpzCtGoNAd2eYt
Hy1JFrvWTqrPb7LfnR0KDYd8VcffdGTa8nRTHJ6dw64x94fL7dFtYqLldwurHpdjJ7n80MgG7/fE
5UG0iNQe1ncyNM0bFDnO2bqVlSNrNCUkJZmPAsZFAqZu2lTDEuZzjHd994xvY9a4X3W2BGkGcrc5
fvAPU/weu+jqkRpZ65tN31RWpDafeFgP6cDr6ykjJXqUNOQ5mQNZUxMY2DMPO8oLZdkd4AP7Z//7
tO/ZCIWs5E8egI289pVgjZ/AlAdct4zdHoe1Wm0eQIH9Rt3aRlKOH55qTrk5H4U02mfDJstaUtEt
M5fmdlHlrKb0XSjllvL7wobaP9yKxY+xQhQO+u9VF8oI0Hh7wOjWwCad/dIEu4D7qZZOvgOB0CoI
T2HySGOxjMhZSkd84lF+ocg3rvLpqvSOjas6whNcdUlnXghEFVPRzMNDpV+75ZcYfgLbsW37S2Pu
bVPr0HE9U8hQmygONCgFREtcHAIbPhC8Ocw8I/fJlcOtYjaaTx1Fzm9yIkhla5EBCOy4hEfzP+c1
HoBFsiTT4LyLAqdO47zHMNLz6CcElAz5Td1SgFlnoYThn6lJrcNiBmb0nyFi55VXb+6JfBtYE+eq
kvxEJivdchaT+hRT7gERbfWMxO8+RfJjUS8v0HkJUKDofWYeuH+E4IwehlWyw5hYWDfD/mDSKA+0
W7uNtFQq8R5iaQImHeYGcT1oSKpAHQsrK2RH5hYnSy7BSN7k5UNMZ+UcKU849QspDmVliG+p1kJx
Q4pCAIvcwiO4L50UAwpbMCXpS2G21I0GdGOTQENuqvfkEfrCczteydHAe3P3koJ1iU+wb661XQXp
jc/HfHdffnwKJuz6yaRxGlo7iArPFixKLF6GSmzOltp/siNDsygnYu1eFevQwoU+lBw+7Q6DHXKe
UVaJYxZB6Qj3NevuY7erhQpBWrxecM8HC+SdInSt3VMXh4jZQ61nJ5i8KKh/L4l4WbC7ztjrFCqa
E0phNhEZ/4Ghu5TInwgn0yoC/7kmBFQg9vkjXjOKwV6QjGWhUYwmC6LlcvYS3Vb20sGnplxS4jve
L5ruYiLMFTpuxDznzDnIL57BqZHxkSx6Pyyk2AgErn8h5d3YsDjVSSEb4hlpVExrcxSSPaKSTv2/
y8U522HmND+5+t/JjRYIMGuJXE1wcNVl+2eQyKD11ar40vdGaMsyljXQL1K9RlLcG8MtH5OfRF5x
lgAt2CEWCLu9JwIaAzGD+2E9OdjglL/3KDaUJlrmg69WlI1wfuXiMfl66TD6aDZozgIk1LyLWhcx
6yc1e1hstxpnO76lSO6ZrxmUiQ8xv1OoB5skJVSzSEv2yalXn17tmOFUoyCCiuEmXWSW93CDmLyA
lBjbxOHKKeYrJPABDYPSyqLKwjjsSUobo05AsX1lSWQ5z2i8A73owC1Et7h0FGrykAnns1Jz8cB5
8mFdhkEGRY+mOWeTv22Zk0Ose+UsNCbhhxNhHrawbvrbhrR8XcxtSfmy2Bf9VWNZx+pbC17fRzme
npNb1QB8wcxXc5i3XMEXK6R3tEV9M94wwS8ss/HUjccHgfl2ZVQbl2TBbah6iCsRKnFMjjSmx+vY
N+DYKnbOwCPexBNU4NYTR/CAcAd/cVQ+CIu5m/R/1sBBiCMh6QZ6aO7G7x/LHn3/B9pJdDPcEucU
Hg9Ibl07ovOdnBWcz/mEYEa2RZNKRsnr65cfSoTdT9nBZeU9u28Eo+o9+PXcQu8gCSApnWTFAcHF
T7zMkZn3r2dISbLwr4UhWW9Vvx9Vl6/GqzKBBQQm8KuBedZcU+72UYyTTJZSikPnXh6d9IVfI4wq
uJKG93im9sfVZzotl5a0i6JGxrMdxqo+YOUoTiHKHViJ/xVGdEItBLQ/cGLvkPniQlJ79lW/Q0iH
FD44vjmxjF7QhNaLO/O63T2cunGyY1tl5uCvbaPY2cP78LFQH15lkfYJivwnvjC3qR6qm1QErLIZ
sUpgxgwMPmtZVmmftF8OOVzE2w7bhcAGSNfp5VsqOvymMjR5aCGJOYMRJBsHw9WbrQXweAlp7h7m
dMo3JD5IpDdcD+eaJ/oZZt5ROlJ8naXUcNH2jxOCfmAF0GSgihG9QZajuJuJJcjUBrQY8tWEVpSv
iyCHXBItIYe11ltmMIDXNZnd4zIdLd7yWUHHsNr28eGx9Jsi/JGFSRRXBrYYvan/j3W0BC5DeYxS
UpQic62IG/PB82qWtC+1x5e5XF5MOHDYEYjutPLGCE9682GytyYAvixZi/5lSaJco/bNBS4kCsu/
fZ8Zv9X1/MJUrlLnoVQvK7JPN1DPUjb3NSCn9QQvnn2Q9EJQaFbCy0+W1/X0GTByaaBZoYanbqHy
jfcUJvv36HQOnxvYNGdQ9qqCKpmZCRSh7e4vgWGlhQgngczqrwOmbLJSHrF47YA+wJ9yN1abj/G8
pTHyFjlNz70mW0ZQtXDwGmZO2MVBav/NV7nYlrO6p9zrRRfbcdG31sR8evkUGhmmd2oepInJykZt
HLVVSdMeZjDisHi/mcfBh9Ws/7TMMBJQBdwM+KerNHcfoSCfIADfROCdnvRWbQzKV6yyTanKiqeA
Vm3KgQaDv+uUOGwTJi2YPp+GUyQrRLXbveoeHLZ6Ki5racdWmJqS7zUnptoHzZ1bPmfq+P2NAIPe
d7u8qg7+4DfZa090PmD/hEv8drmRuytcZg6kIuyPsSY35xiEDHWSymDVjwVgfN2Y4LK8eRGmdVlx
SvabFdhaVSbB8e4qzhk0/NMVHpvIVIGR0BzlTwBOFtJqxK17/bHVQViWuvI8qXsBS2WG/w2ho3r8
TqlO83K/k9N4tRlz838KyiMU/ItPRpbWERK4gBj0L3bef25ReeGk6fLu2fax/doj5eDkxowTq6QR
ai3ZfIpW2OYayffoczt819ZxYYuEZoD1bBH/EagaQHa3o4+bJJveE39mwg5e3wpAh9LxUuRyc5Kn
5HWee5sVAjzOXwrTsISbus8VrH4dJ22ygNAKAww6n6Nya9cwIUFBFhmSAMksOMGcHb3f+LyHfU/D
VDYe0Kv8vcBxQrbxVX5D1WKeW3whYtcl6BMvKXscfjssY10R3WKlINIfqQ7CxxvlMQbWSDQk1+MG
TZLexyXYRyKLQS6xUElRjUJRwFQCaWkRX3m+r8JV/NKvsbzJguy9TSxjQfw/SF8Ur5B5CDad6paQ
dfEoHJWiRV84PhSuuiMueb05Fsrd5zswxvW29iiX58HH+8wYja8wYWhLGdRHF03jbLUrqX1035mC
yGRuQ0g3gPo+PBikpz+SPN6bE+3RzfXKUCxdal8qUgshRdZDxwbnVrdn5wIV0u8Fn8MNb2pu+HAA
80XCv/gseCW3qHbPrCn6U5IZvbNYNLfsEuKIvpNLNNv5Ai8iMqZa51foUKrvL7LVof53LUIcSITq
P8Y/ZzoWe9cnErqak8m8JCneiZ9P/LGCVXjOvP2gq7qra3MvFaLD/rWrhdzp6nFfKUR5Z+NbuRuX
wmLbV6fhZZJIxp3UqBYMUbZuDnvvMW035j8T0xlyKEci9lcOpdl8ooKcKmXdlr7IO9uBijuQV5sT
RCSDK54CZEHVNYh0byZJYITO0LO1r8eSPvA7fFyLy/byVOyHIoltwzKOJ6SJd3a4pZFwo1AllEzG
65CwuJod8n5UZj/J1HY1nal5OSlBg2qpeRKurze43sSfrvnB+iOGwSLNiIr4YpP7+HlNLOmrxvXW
YWj+rc/3yn1KR1bNFxDdofkGqx85AL60xFMJ1Xm4nUgfqx7AnGHzUPQSdishWfLfLMoZU2mKh1cj
hyDVCnEW6sa8bq7jX1jjkiI0v46Mg7/RfwCB8hJAUP1FEgCvBbzybeXKCGnUSTqGomhSl1dSZuKq
l68wMuSFipiWewP0mwLKWMifC5USBsPemg9A9rm8/nlfNLXDJ+WpEuWq2hudRR9s4gtUz4+9P42L
2LhRF2XXyluI9fUqZ4xXnitUxEkk6ILYuD1WJKCjiMYs3K72nRbMGyvQ5nNB7JxXd8cRWWYnxQzl
wIsaF7Aaa7D7QAR6JqcjyPAz4nRtzaIhN72PgrN7PwsnaSPGVwvi9wiH0uREc0Ed6k4EDWhAApTY
AX8Qoxh5WlrNWb3LjGUQDpv7xv85b6D1hyN82EmaV8V/3tlXeOHXDg09LPRZVXoAqtXWhexebN9/
9ni+TEz9kz0lFLvUGXtSI2SyAOmL3dcMT0P2FLPE/WUzYEKHcMuBjynxLo2AKEIu+MfhObDFadKM
p0vxUnG98SvlTIbWE9ezUAekpWukdExRNWnICShtnn0IpCKkOlZYGFQylEHT0UtM6f/v9/udwapj
4uFdjHaPHEoSfDw+xSdNEusT5+hcGc2VO+z4t7gSxPv+kmHZ/NxPEvzgLlS6b7eC4m4cyw3U0uru
tdr779wf05pAXpNGG8o/c3qT/eoeTqP3ZoUAbsvrvFzt7Px0hz7BUU0iZub7oH0D6qPjmhI8I7GU
rQauvsAgoFdkhTdODDoz9nG4Ju8GIj0k8mOclEWj4ZRgy+1eYKXKEWMOPJdbmg837TucCRevccRR
NQ3DRNxmDxxg0OiaBPJcyf2ujpPgU4cHmIaIlZqx4LpOvn5W948cumMfDMeE+4QAEFnINpc4KBGA
qyA9HRtxJBVBokrXxFTjpkPR6HJ8sJZW9lIXxcbXV/9ckZiYIf45FIPTo0De5xve7Y9QaKLqi6wA
T2L3EvRiScq0k2yrTWadwob4GoxSZHgJnkoqrm3ZOcM6oxIOfKOObmREhh2tYa4PF5JkPVuM/GEq
WZ1CsMOI3wiWiLRqhOr0qYgyk7DyRSVlG1hqi5+4V8aX0DHSpd8FNq3dTAsVG4LI/Zp1qYbdIYoR
r4vdiQ9ieM4dxPGWqNb/3y9A+G1BLBhzow/UC1sE1A1VuWpYhwF+YFXIHRaJ2uOifaePjeuj7ch4
LKRWeom15N0DF7h85exGhLS+kEtjZSNGadID8jO9w0KYV+XZpyTdjlVdOaVveP2fRI6N/eCu5HlF
pNHr9TUg7SSOGYNaAUAforIHIyDz4k7z1JnW5Er/0SS1svPFdHUIjjayvCSXT2yZD0a8LTd8ITH/
lGgCY/TgOvOlFSyDds/+58kj9u1Bu0/sWzSVT2hYet5g7KhhV/LZw6PFzIK6cr3Ak9+V3aOyuyg+
M9LcDneHGWL5wOkKOLeRYGF60to5uTKB/KvVSfKw5TtX1AGw1VuZh4tM2MfqCPR9mj8Aiyy/sIAs
H9xoDC7DJBYRDFu1h7USbB7qcnMNbEXE7c3I1W/8CsqHkkJCDq/14y4P7NeVNHoyCY4SeJvh6xnm
fpPmOPeBWFc6zHMdhvSc0zMEGMOlROWcXRRuvuoDXoVNntuaJOhYymwxv1k2v+zBveMOoi3sHhZk
+yF/8ZIiMeZPTQnwcBGxAy1NQofbxn99YTmEvZ7wjtHh4W+QLbqAqH6gxKs0wGovujB9tTEXmG3E
QkbUgp7XHHGRKZB2Jwp81p99sIUF2JUsUiKff9PQY9EUaRk5tY6m5rWrcWo71a3OsN2LCetv87fg
//uez03O4JpD/EScVAUE5BVMCLa0tQzKOahcHLepm0HehKChe/BSEzZOZRlFrH+PaTGLwgoNhfSQ
Dqh00Iw+nRBDwMltR9WLjoLZyHph5ovgjVDFeLmxAaBmIJvr30Qgn2kXWS4d8ZQtqNP9L7s6rxbH
VtJjaMLEpg+iIlBTU6fGAaRU5r0bDQDz08Xf/y/5VE69NQp3Ccs0CETwmozRr6gDdrKMUGq/nwPe
YcB9lRE6b4NDstVJd+DUkp8UkPDWTmUQp0ku9/If/GlFJ0tqvYNrQvdimCiTI/PnDmnsI93p+P1o
nlWWYfnGcEbkbbc/nE9hEwKSL39vKGNWEjkH3Vzn3FSBrsF7lQfaleTPJDlRYETvZee291UKrxIT
+GPPmCHAugkR3CYkCTzH3yKpo+0lVlBY76Y+vRn8wptxQTXmtP8NCDsDKAshNZNEKlJFa5zHDfkC
rN07krJ1OpFst9qCaiqeD41ik7RR6KKPzaVKgK2Oatpu3MJUrkMXHsAn2cAeHfwYFmIXIapITM28
/+DUjTH8/PAGIUpuUGg7NbPK80ACEGpeZNP/1r66wKJfvbjfsqyMWKtR7qHQ5UfGox0OwUS7axyh
1wxTRfFsC+Lf7gln5o/m/dU2uoinEywHmLl2yYl4VzJ3dRV9iN6vDg1cNj7o8NW6OgdiTZOiVhAQ
9tHD8sLm4EdiX/x2VLUooWnL4tlMbszj+FUu/RakZ5a2oZTjPK0mUNb/Um0e8pRhsXrqERE+iLzG
8kJoT4WJm44GOUo0F6Myy1q34d+n9yfWdWT4zCccOQMtIYEnI0ldm+72XyAdWsy83DUDs9zMAVmE
0Q/dwucbUlNtIEhOsHMEzH5jGBhu74nk+W2bhAhUpZMmBVm7PRJc5qJiJReHGYycleqkpUOndLbj
NB7o+lh0Bht76xFsxzFSqP5DUnIfep24cdVgN2fyf6uoofd4XemcfNlzUoSgiFvTNM5Fq1T/gngk
L8MqC4QiKkZeaTgBia7lZGaxVB6iJyqR5HD6ykOzu7EoTnwGsSzQ+T2IkfvKL4rkRcKtJzjVScgD
KYOkvT6RM3s3nT5nvw8I8nZQgX9486R1RcGpgy8uN4zdNNK95mutfll4vA8Vq6jZfT2LHbG8D7Jj
RFlOS5u9PzGn+1NPpH6QLWi+f6/Jr0poHjhy8EhUiOaY8hZ0Hzo8j0/zEpAvG/lyIeP84hQgwa7f
wWV3IWSLvEFcolU3dmQqhCKbeZSUghgkPcfJ9tVS66JtkV6cheOCF32DO8Abc71hI68llNsoTE7M
1ZxiMOKlXj5Binhyiwo7WI4Yp0hbcSUuCvqwSb+KI0sgPtz0/wT4E2Z70mLZgixF7xGPWDXzCs4V
p34E0q9/Ke2lP007H6MrlmUscaefTN20FDDOMxedq58n1Fp/+80HjeNrE9kW42bNX55RPZP3J2wG
eqSaxcJinybk9vkuLKw4Cu3PiTp1ki0JPosweGNXlZOHAtBtzWAgdY8/YBa0OixfqTEGj7wE4FTe
gKDV0/dTYK3OFDhbwh2mGGhYSGoFu4uhVik+TPuL3nH3b+42XZL48XU2Fn9urY4sU7Hz+8EVr2Oo
sKBgOrAuYT4QyiBVWdFGvgW54DBGzL213NgZaP8KqQGAGcg1vbQ1WcD+p4V5LCrTOyh6WnHRD8nC
XtlZ9jRvoJQSKU+kfjDMlBgoc/uu0Ek9W1N27rVPFa7QuEhWnyA/kV+SF1A8Vjish8FIDfu2mHxS
4XV+3zzVpUYx/H0u3eeFU9xf2swFB0HygMuDxa4zBMm7AFkLz0GZCxBpvVWPFgMAL/dpAMEXUTsi
Dr7Pew0S9XmMLX5QWRaFCtSAPyxqas++GrlDHb8JaiNgzfennoU1gOdHtNTAVNa1HibjZyH7msTl
ugQF7BfkDrgERUc4Ejl75DEJAH7lIrhfE5VQEHSKGGAwped0GIAJfft0id9Hm8Tua6DsVHtHqLdq
zMqBXJv00shdWYLFgMUC6HdKyfTSgha/JdC1RFzuzprXijLh+U3pKTocsY91T0/cgXrY+IOADgV3
fMHnKmNxh76UzgEO3Cexp2C+fO9FTjuybVPRxdnRAs7KGiuj2llYOJ/dPGVOjyceBQBA2cWBQZOY
+Iq2luyEKEUDq5tRPUuMTc5dchzy6F3913yLl35uppScNLGkUmEuWIQvKTvZa5CzOEOiZ4ZSky9+
wfs4j3rqed38fuHyrye7ANCv6B3K6lduiAwCbiUT0fmH01+cdXVQKsGHx3zB3i4h5LyMEHVkdUUW
NeOwEPakd2kg+pWkVZKjKwZ3E9xQhD2YsImxBx4UdnVp7kG4zVtI+gXiY04P8ixEgUDJkM1NtWtR
CsX0JDHORrm/VxaBtkyjTYf/oXC81G0dJmeUk9BCxnHkBY1ubq0+tBuITtHVEYZURpA5EGxh8wna
tY1E1Kgvj3dHy85lDXE/iiWKw64vGpGvNPi1CKvxR0DNscxmgAPx/V838t1p2ed3XvAO02QGdaA6
tbY0tj5APAxBN4yzmbTSKngFQ4iZYqx+H+QBlulDEAcX13kqBi8U5oZ/ciBEFHAqS++1iiTJRvVO
JpcV6QufpqevO6SCQ9VQ69G8TTZI4iW/fhlX7Cn3WM5lk/6cNT5VEakeXu2jXFj2ycyjNHUfquzs
yakfSarcX8oYTukcV91a+QMow2NVuVaak1ZVBSTo79q3Tka/lPJnaH7bfSTm3wgxet2QU30xmupW
K4Ywfob1zw4O5Ms8gVDuTfz9BWWFeW03pBBPgeYdibRnGeoBYfnwQQS+ocPXaz51yTHkWIGVi0hy
FOSgcgSOhZlo6wv54w0H8sEjCho6tdq6Qm6g7zJ0sUpB9wHvVkYAMoaVU3N5hQi9XkkkuVLG8Qpr
r5DW9lgY4X5gIRni5rU9GmkgB3hm3rJbySvPqVii8uTObhiMHiVQd9BzVtCnA5SbjcreLSac4ZXE
90CJmIy8hbVvhugMEfdyJiSsQhRxIS9HpTR11GgbevwsZ7FnR/MMHHjr00OY63fvh9bpeLFu8ciW
/XNbpfD1BIaHJ/99rBP8zLHoDzQbhnEpwqxDAeTXTxSOkX+WsdP4wmeQvOCqPQlL/iQQKFxKGrTN
GxQ9kQBNUtBQd8QQjEq6Jre0W/FNR35Rm4Y3B2DIHfKQp/ZxhH7QkmljMGngCFutCBvijBjR3Dbx
WPkSBFm/0l9VtUsff5UIbXu/uMqOzOc2OvbfzppwnnZdhphsuoZCG+iegbmmdY51c67xdVY4pj9a
rtrDmwQuzImPuyw/hIPQOIuS4sNuleRWipty+hN7hOfWM6iRjum+spjqoJgvSRc5dTiryM9ga7Z6
8NmEDMigFv/HCW3ReXjP9b3HY8EHDcYpOWZE/znlHiIB27jg2nm3CC1jE+2Klj12SZVXcWaXbsMu
vIhTfw6G9HWUF1iBcbx1q8I7RcQGXJZZnHFUD17vB40yvDhTbn9KvCz42M6rr5i9nRxS4+0qnsQw
5ta2u9gLEkeBxCNqerVoeINoWv+zrJhcKafH/kYdGdB5wgODfR41ySHuVDD0YTWspfbd7mabBOv/
u7KeWUk6NeK3nws8Hln/jXjcL3JbDUVNJYgK1kr7FW/g+MMKmsEAJUv+J7cdKiyZ/Np1yK1/f7Dy
1Ba2EPLCCYwz9HtBrrsgaKGAD/fEG2vMuX3qk5rE6JRqP0QDWGw3ER+vQkFecuDoB8ekae1gQStp
qx9/d6OwVTyVJQTcde1dGivDhMpMeQaG3zVf7Sn1qm/xxa3l3+Pg9P9VfdHLI2LUnsaM6iaULvPt
MUUGYXjwtA523ml/JRe0/Pj/qygPYIfpNAKE4iRwn9p9y6DTJMdA11iBy0uWJWL3vMlrv2AdcQT5
tMrRCJDuNnVIjG7uuh+OnHM3zKMNEZ9TjRXXbiwqK2KKYL9trNHzYuoqUHWRNMG5ClphraR/ebDv
2Wu1fiUkhkJjpzLwwF2gwzO9l+PGp6G+o+tNimnjXy2Z6WokqKROAkTeJMHpmjdDexWpU2y9oS6X
HulS9WXUk8X90yoge/5y8l5l/xnpLGCpbJkacCsHesgB7rUK9n4IfXgkg0w/UGd3cm4ylGht+JRt
AMB08QHH5+WJwPe7jq21wxKqIBX9FA7HAbHpTT/culpTWJwjNYolAbCj/K+hY/Mu5E2SfDH8ovVS
C84sTsUDj+ZaqLjRH6Y2wokHXtdDVvcjfhZnAA/E7r9pWCSfUw/lUxugFl292UGooCyakW/uobkA
sEI0062EwOLvjUC2HDe0S4tUPkc3Gxqrt+zCBazzOhX7/MJ82kR6SQrEBaq5oHijRTLuy9OGRstv
YB1tKx/vxaWIzvx1JfpfHLQQtTyrB5E55ozlzSWvtaZJXuYtXTEGOTt0bGQz9guLuDjlyTMfhwA/
FBosVw0fqZuQg0waQ/rlYW7+hpnnYIX5voWeV+xXd0so1v5xqplNIb14iCRYRyo+zsQ7ZOGIabro
SXjQN9WM+I4/HqS9QH5EbNZdtE69Q6/ByPCsVAMtMx8D5YCPbkfLpLwwYf+GlJGmxddLKlAmmLMO
DR9bLr4dZq9JgWe1cgjul3CXVKEWt7Q2bev4uYZ+Ng8u4pWC7kGnStXZszstJWKXZRCo5got7V8S
0YTcceuaVZuyNJRpmyHH4zzKzKcsayW6Nf3BmzRSzlm1eXWidMA966/z1s9JGtLBIeD+5d5Q5fnn
uqMKbKg8G7wdOHCBWQWy7YiJzMolObvTQz+NJbu4tcPwIu//IC7/7AkRnasiSEAbYvJ8qxacuh3H
j+1Nmcm8P1D8A6kBDvp2KzSpV3M2lMS0TDQJ3T51uKnwoOdAOTs9zT3qAL3KvJMUslbgAgY7gy1d
vn1/hxL+GM+9azOlOpW0uBDLyv1ncGgSMXGDqhVxxIP1STs4fe6zhC15t8z5mrr+e8sGvR3IKVkG
yZSjHqKvFi9U+oJkXEfH1VILbW/YvmGD/2U9l/+WiuwSpsK0V0qmEp4vygDeQl2fa+/buRTBSbxv
X0RhGT+x3jc2hPCQjg5D+/SKrDw/FpZUJ40gT6JcJToUvklB176TGsQfIrLXhBQdGCVjnhmLe6Yo
obwBq/yCb7hgg++yMtjgiLP521HGBvMGSDqo85YgbXiCwUT+JkmozdI2GFcOcg4s88xMZyLG5o/I
5kFgEkknyLv4jBY1SHCKMFq0nCum/VmOH3KmGHyMqV+s/DMH+o721UaDvVGmu0ymVkw2HD4TFJCg
Bm25KE+vl+X/mVr1CejNpCq/tgPnMse08f11oKANdTI5Sf/yQOD5XNtnyW4PX7636n35oaOE62gP
skjIgZMZdSK+KfZaVg6HgOoAnQnyYD1AWDx3Pe7K2FIggf/XOXD0e69DJF+Vf/YgQmKqrcx8G3It
HPmBadXPo0kG0N4O6qwKHfGC3u0wTwGbY0C+1iDVBNiyL2xmMYKSVIW7uzfugmHkmXhEA5YvcqD3
8IL/f1MHrxAr0PqYuqLD8aaTtVCAl6erV1HNP3ZE4FRU60CoEI35gIKnHhTGU3TFi+HFC0O4hvqu
xRpWMdz5wRNGBx69aI1fylx38BX2oxVMu6mMZW987sFqrigBSwIxJ7O0X41yF6x7rf40lEb8JT5G
OKSVrnEO8648okxFWiIo+85bUAyGqtAqB1FqMjzT4Oz6rVgcwX0rynSRr9CcI00+lvY+lFIQNd2P
I3HBJ+8PRY84jLM4eR3JVCdP2SilyM9hRVWc8f84vPx5B+AwoXmi3YAuspdyi26ShPCwbyUL/k5O
G0DUdKIgs34hov5ztyifF64gIg584PO+B5zh4BwJP7MqsGEY8l3pC9mUxFor2315tkOWAcqtFyKe
Vpv2FeVoEUd7OPtVorzF2/7qcA/HkJZ8QBX38BXQ4q4Xz3lXZy13Ib4LjZApmC+COguA5P7beWtY
o31m5aCPepiOYS1038/1derE7cLEQBUjDv2dyJ2gI+MFFcdu+mkVHg3vpDZg0Bgov1yfx3Y3HT7Z
/4mLGa8Z24uLqTIQwlC+q2gUPxn8u4olIDGjFodht4fP5c1itWwljLASQSk4FK8qwqwl0ADKj0YU
UMv+lFLOkqjzEEBJ2vzs+hoRy7KNcLG0btN8MFUuhBWLGvEeFMahRpBRrOU4zLNIqU53SJH5pljH
2MyKswJr7GW9Lhjz/3gsQOMn12LCUY886CDQqZFvOeiFur37+zbuXOUxv96cqEADJAC+iM8iDdEW
JL8Ih3ZAazT5X8j1GCIm/+wDZF95+VI3uAiBCrfwaRnAI2A9uHtIs2nfjHut4XspQuh0krYJh9bC
aJ0WNpKTDPVqyFyoqpDGxG3Q8TbAwTyzjWidLm/Gsl21CurMrD0nDEk6/T8e6NlY6e0HbAdhx8oB
HW/2XrleqVmsWddl+ohpHkcQ2aAx/htJLTGZX3RJa26GDoIrRFBxA4NchBwoFm26B9KMqqcYVg4p
9PEseUqdmwJ0/GvzEmSAzvh9JXd0wWNb+B+ezgiy5YId02eYZYrILqrvHBRuTvvEmwnH/N9jEM9P
Hqoc8pt5aUqrsmSgBPTsF4nQAtFgms1VV2lu6yFc97BCDPqRndsY9MCAbenohnfzeS4mOZTQg24D
Q5/kxHrspMnQ6SVkAKDWdRWVN3XuPIkCIht41hLoDapZjkIRqyH3yGfKgrjQOUDbn3X1UMmRbnof
bvJd2Av4UgpkZzQcSsTXvkV0fgoOA5imHYt5MXG2rdvb92adiQQrX1/o036NqiXWON+1npDekuoH
ZOniXfYOpVzOCebvoVTdzDDMh7m8SOfK21xrrk7S6peV3JY5L8Yl+WyOHA5FIPwg2+O231Yo5eUq
zarebxLOkMwj27NtlWuV2LkQw5gpD1iIAKdoMAhDjnVry76qygV1Fl1M2djho/XxkKrcasK9nhGA
6gSWJ4bKUcLzKOn97Wy/G34C5nC8FfxOCyFoPM15eYW40kyvyiNxnofN8dKufPCisUzSPFYUx74y
NsWDCW/9PZqprkr6SmzE4j9aPPIAwjWjIJyoXj67QRPUVYg94caos2XSEbHOEwhCR5jYrVKvked4
ibM9mSnju5FgF+TWfYZ6uPakFsJKGthIQfkkzWkTFhrPoh+dj+dAWYa9di9fWnqODJHdD991t55A
nYDVDbGE4CnV47s+QczEHK/E+UBNcwFEz3Pp2h9mnYO4ZUDHc8QoXbF+8A9ped3kXmOM6fsA3uFe
jQT/HCk6/JETyrKzoRzaCyCnblJPaz8+j+fAzL3a/gvfR3NibDSxjsPTHtnjfcy2+QXVx+uxK42m
12Afo1eqKB2XNcJYF41Fvl9WjKnBm626cfkVwShH7hFJunvW69tobWd+i8UObBAqaUuhFFAisqI9
xULEQpAKB7j6EdkaAEJ4Kj/2favvm+cImaa0GRtNehyNGD7klj15MR/Dfk1SMnjuDCMObXDz3lK6
2+qtpqLQUF4bSoLJ/Fl9qCxWm6PVOAxaV8/pEh00mX2xTDLKMazHBacW9vZgcWKWtP6ChRNCwKow
nWBxZI42HUqcCW88Xu9Cr+YnXgy/+sISndKRdZRyMF+OSY1DrLEUaFGQXVQiyNZlFPds798G1KQT
9a8GbmmlhWwW0Q/wX7dHep048BIR10/P4PgkRn/a5z24IOy3CjHCcxGt5oR4GOsjD8LDUaDXnZMM
9UK3GeEZDHXjcnuxawH3W2TqaWxFrLhthjqkKePftdOfFkzslYg06O/YhZWSdZydwBNdl/aDwS1/
UvDTXb3HQ0OS7sC9A7xmwNolVFeKAR0hIPI+OOdrrgW9ZAmrPYgAInEydPWkCBYSKLqAUJthbrrb
7jcvVrmoGpS4KpDOKOzdncZrkRfkgGBn0Ah0+SArFe9Hk9wY0PFYYx77QfkuIr6jVfdXbGcnbhBP
3a8Cm/ZrqmX1oXQ8kfKU9I0KtO8xaUCx/JN7PXlzBmjbI/xLTTube0/Ten+otrCIyjP9pNY2Esx8
GukF6OA7TLh+k2sLiCa+BFwX6QriIRdt8Cn/4gADjZ4vxpGslgsvpclHKoV9/Pi3nr934vDHFDkH
DsRnOC2lDmq96+m8lpfXxf9rlyv+odYSO4ifn51WaWV7YiV8ZKTAzu0kTuCCw8JE/eGwhif10CRk
CEMMcZyeSzZeIloMHZbZTPJwSjU0b/M4ZgNflH/QR2sg5WVl4ECLiSCtpUXVnS1R8FMeclKQ7nhH
ihprHvJEwtQb6WYACjhHTp2FtKmPzVej+WbJ/BjzqPpihLfphv9dIpT5JTEdBiUfRN7IY9IfGazu
qNt78kmPqZ7gPrjNb/4MvmIv4liChszNnbN1pEJdBOi0ouTB3WYI9qNhAlK3PCCKJDN0hmLtCv79
1ype3MG0GBnUZfG14BVfKTtzF8ZNDwxtYCBEj8xSsw31RGeLuA6HEtDRawfCZqbqrQC3Btc4CiyD
rKpUpDQ35UUAJZ53GdHbyBxjuSZxO1UGkSyNrPo/oNX2pBdouj07oJP5SJcUNFVfU7t1aZOEfbrf
4iHwLSl3G0/hhETC8T9mJuWZrjzQW+tpy9lAWwbB7IECnZBCLRQoGchk30zB0YXhZ9w+UbYe7Ds5
fKhflxnbkFemVUVhppoCpnoS1ij+45rimA+83hdbo7L19QeWs5n4E+kst7Sqw6H1T6SqK9nil329
y4mGyKoBoJkYqrS/oyPConM975EiE0gPSyWNbYt1KJkcqzeWZIiLnJdWByu7827VnG8/me9wrzxx
vEhaMQM64TK3X7Dq+GGgzh6p1XSQdFRNriJ3vVikUMX8zFroDOEVJSBDgqGOJadXwIxgLKgb939X
tndiWyqmCuGTsA6nG0ggUyPFJGObVJW5oTFDwNc82HQnUKGnI9dckJY4INEfcZDMq+0Hmf05QVmx
aULp4S+G9ZiT+pxHHiGWPPMDdX8GcjEofnUwNqSmj070Y3wsguU+A6NoPKdfrD1HjORjylpbT6ln
ZiAXUzkSaxw02zq2TyBBTHp6DdTfyYvRXcY1kqa6zPmY7HuVJzU3lAax/5SKYAZ71IV8DeJjOO1/
quD+g7USyel//WbbgeR5Je3JLYDk3+2Z+j4+7A0hVSMEwE0QqB0IIbiB9x4P4ZkVUmbINICuC4T5
C0z6qNowolCO+ofEVQiTI4/giyDVqblyhWJUf7H0tcMwlQWsEJn7SXZnnPo0tg+yeDAn9sbl2/y9
spjTG9//IFZ5i+GIaCah57DD+YiABqxGUtjP/KdLHj+WtakWoB5G3dLkEr7+/7a+nJVhPmgLQNaP
YKiT77mW0y5XCGpQGdwv28+FO/ZJ8Ja4wcH0yWK+i4DGZZFtJcwnnb0s9ybhGI0trmvOjdfmabLs
XS/AbdMpuIKSn++K0vtDBam5fIPp4ohR14A5Sgl5AK0R6AcHWROpQc7gBqoHQVSIfg1BotWTOCon
xsfDXfhgFsZa5xRow6Etqug2hY8xUdqoaSKRdbNx19OIFT8gEFkq+wz+vChOkMYFIxpIHudihwbY
8+GjI0yCEvpOKcd2/sgd13PYZlhzSIatsaLWG9KbrMwu2QX3pQxtZgQy59z39f8fuI74LN+kpJ19
oOjgJlrRXBLBEt7AofVtmffWZqaVdcm3aNkRdvhsCtk2jxjuHRygKzZgZDP4uAjIOyBETNNZVyBo
/zX64Ze8W9DxvFSimwtiQ80RQXrGt2YDu9mPhPiUB1YUEYd8b5RReLOugueA01SUOZyVGxGFVw9A
dWxmY67gzxmYaDAtYeWYQxyF2aBBJGuSt2D6d+fxRsaG51AawBNz5IFXoUanMGu/J3GQdac4KJZx
cq1z19nn+KRMHqckO49Azr5dV4QqVEcP3tX5MViqSXSPL9/34enQYjFiHcKQIfKsHkg8N5VHL962
QLHp46Wp2mbzS77OwbqBqoqajJSeDksbx/6p99QKRJ28r3s+BVTxeNzd2nrda+OvyZemM7dKZBZm
MzkS3IjYvutPcV4rm0OZrfgS/9v7/SDbx8iTWM86HO84YR2crDIgNYGr073mh6IpGRudbYK/hc9x
mnF+35DckEaXjrIIlJ/qONzm8uqIHIV5PAQYH/dneyMGIi/bO628FbUXrGQIvRQELEa8vl3mbe09
SQQPkb6HSP8vtr5x/DTgOQLpKCj2lSrq32reUn06kKSW4BBbXON9un1yg5sOuVFvg4duSfy/+WJN
H21dybqzbrIcHQ2YurNPUgQOyGJhtxdCHRNTD/Jr/bUUPHx4xU2Vw1SWovfnfjiS6DwfT0nINTR2
GHEy76jm0ek2N4mPlNmcBDFaTR0SdqkU+7xPnQDurCSP7NUcMVsUw3k1bi8GcC57LISVea3sOUEx
flbpDH/xEBTJ7NvD8qjSbsGtJ9Ryys97jjRecgZfnuXFGTJpU3MW/va7vOzDA1jrpPLWxrUnaLL3
d9aXbBDjSCRol3em/bxId4CUgSutOzdqfIPXvzCBi3/ROQnZQCDHCu3RCecd5c+C5tPcD/K71rJN
VQuO3u8WoNC9YHKW4EmyPeEKhFFkO51lcaWeXIuJbtL09sN+kbBx3RUmZBHYNPeIxYqZ4ei2CbZm
cmVIAgnSCURGvXqgwkFwr1Ytp2JPQFIEvAut28YEhdZaY2V/+1AIcK0IvkqDE3kRx7z/1lOv+/aX
P7rsqLAY2If8V7zaqu2lTRbo9Dg1Dsb0iwJ33oKc5VG/Ksb69wLVYL92KmNiuYJR4dz+Bknh7Tmj
2KnZynJLY7ZHBGwdad2FmpRN6My88ajH+pO7qEt81HH59WWCR6ZX8KY2LK7rFFbfV/amPI/vNlkF
pHxLrTmEw0whGBOQDPeRqS8UxNLkTGLveWh+BolJuRIK/iF8zttWnHNQG/OKB2hkel+FEpvNIltU
5PEFqFxpGfqWYWwbv5T4fMpUVdN3z178ty9GhzAC0IY8jL+LAcgY2u1gteZVOBs1Fr2+JRESzONW
g5tjseeAs9xrFN6xlHSH4tCYouke4XasSAPCR7W33I1fP+SS4OGTPswj2y1Bnte8O7AxLrTlUMMJ
tHehFaUFDS/1dsHK//JuyXKchgb25iEnatqNGRPaXQYiBvQVtDH4SdQ9Vq75DG5ThnSQ8ajYDBqA
fWTVK3sQL8M/2CRhWm+iU9TO1WgQN4yp4fNUhg5xeSfjLLyWVek/mPEvc3wk8Qh/pK3UH4nrYhVr
dp1RQKVAlgXz1Ug+Ww/KQtZ6pGWYRBt06WwaaH9JnHVkPtYG83Dtt2pVptO9iYFyAXWk0l4PjLrD
3kV7ueH3ZiGJhA5errMWHC1NrwM0l/0yuT9ZIp3ZlqsPZJrmKcT2+9QBLxROnjm3qDaUQF9gP2Uo
uTwmGurKbxJQ0MzG05dCwuLd37yCTjdp88y7MdjHrGTLqxn+cuKUULiyNcrwPVmB4P+o3uO9SU5/
Bxl/5TuxXR+yXpcUpdTiQaHcp8hktjdAjaou958SPVE3noLzqqsadvmLAPJq69scmnJVOlz7q8o0
0vXBk2oV4p19hyPEqAp5csEiv/lCbOJBBP/5o79IJ5ddEsLHYE1X96SDl+bgMeVjLyD2SZN2iGHK
mjjKW1ORiw70+3U0r/rADQsb36PeME6HwQg9Wxtnw50l/99XDqPV+ED4dKAM4QM2BvsIbc1SnIMU
dQolep+VKCXDZhCc7Unno6XGbqbXbsDzjmZ3OFFsjVZN4k3hwMJ3G+eB8MgJIlbTWV+yP3f6/Yfl
q9hddLMH5bScbH7jAjlNsf4CLujmSGoFFgDrIsPC7DcdQGOVLLujdU9WkAdybHQV9YkBycziV5X/
4C8PEScHFXafDOPCoWO4WmTxfMXwJlc7iJnF+jUJQF9fDeuxwhqTrfr9CNOSWUCTcHDZA5oa9qNy
rLL6f6r7HlFLLN18l86E4xYNWuDd2tHuQR+IzwQOQiPVr7XUU1Frf9vsowfG03hdgYuIH4bT8rHN
Jhp9UWccOSjM5pqh4XJ30D0z71ni7dXF4lUTwUZ7Eieaf4LTIU8etlPsEFuoUtHeDlYGzCJHych+
iFoTFbz94+DWi2d+Moum7cdsB6gUzB8ElYA9yHPhebfmsEkGLKBQ+VwiuxMa4AhJ8ngVxMhVr9+Q
zBXueiv823FojymWH1AkSO6BZ9R54HsOjEiEReqwfYY1fZ5g8eSTcXfUbYBxW4iiCF8em8ZXVPqT
6fvRFAawLxvM4gTw2vQEExHRcgO9FShbrpKBuTMz78LPBIvBKrpdq8vUOtqWw2K1yWYkTK9ryIa/
AjMm6/d0+nNcVkJ7udOQk7/2qviueKPCuOEFsnwHDWFQKrM8jSqVjecqPNnxUulL6+l/VSUsSNTk
kklBLov3KJLvuhTPuhs8tbvWpetRtMcwLTeXbhVmfty9ZnJfIi+GkMB1Xthdh2Kgpux+m2VdfQux
chiW9KLqCLeTELuTWzd4egYPMssaVgZoP5Cm04AmoMrVS6cqmoC7TqItjEc/8ZCwCrRvtcxwfqJj
qTYAfjKQCviHOiy+fOhRRho570ffMHUAMUKiO6rNtPo/eX5+wP410UvmjqzutIC/p0tAqOQ8LRD1
dMS/JYpleSLfgXUq6yEmwAUHs7i1siV5ZUi07cJ8zELnMdk/raA93aezC5axP6ircWUdrNzHCc8k
ecUwCZakPPJTxbRDr9YrXBhsNxgURLAXIaEgiLl0KdEvCVP4Tm4d52+KKcw3WKtwF0w5uk9X4bf8
qblsGwktfn4ezsckYD0MnADc2Ww1CYq4OHzNhN+vTp22S2WagFwQ1U+DAd3mItWXN2OMMJX4ML10
CXvOXlGmv9JNCMqTF13CmQUVpa+WAa8QLNq86gmsOMIxhZJkpeX8bZurf6/yf/wzq+Fn5BrZJdYU
Cafo4prbekdeAtSAjKmf7ruNbH6biTJsvl8JufhxnH8vRWYQJIx9kaXTyQSGDk7SEJY5WqGNi/y4
Iamwbu/tUOdn0zVV0iyRvdGjICbmAjet8+8qG5cVYvGNdmS2FarmEsulZo5t6A7xUludahOVn4RH
MfE16TdnELsGzVME0Z2GpG4xRbl259yTwGNFeRbDJ9+Ytwj07WaihMz4PgiHADiEoTrEry9/5tEm
rkR30qhQCkIZgclTtPG0Z5oHbtrmhdHft/8HGdQvn60j0V4QWC4okTQiWnBSHk05ad2BE022eoyy
DSxWNNergSL7EuI2HAYLVzIuLpkCMLbFV3YKCN4JDTl2wLpwCpqAyXDIpz2GS8gPtsIPBzcwYYBr
vgK+XJ9rXETfIVXVCeh/T20ANYoYBzYqg7jlLL0ZWPCbfrncvsj1qWsZNF0ovv85bjSy8CNv+NNd
QI9CjI1FJnwQkjsSKEdC/UytxyKJt2PZCSw5ibYEjTBszn0sEw1mRQC68bOaEaCD+WdVTvLvXLFH
naaS3NttIge3SK0vMBK5zzE/ihYnE0JuCryK2BRRTdiwcOgF/8rzBTyKu5/0BeMs7rI9nvGByyO0
uQRsLetyeWBSc+qAhHnpFDyYgsIuyhX0bfxn+flXD+1TZnG6GJDz6JWM3/jaDDUCgaKWGg/J11YK
Rnoz81HPpY1qO2yP0TxqV9vtPYDpqPVPAqJZElE4F1XjWs5nmdpB0z8osxB2Oy8OBv6WToNmFdyF
dmgbP5GO4KXkQrzZewXM/O4U5G82Lru7dhbFnIKPyAr9VDB+C+T22velkRJ/erBxBqAeCYrOATo0
0y/UXoCDVdZpTxpSpqnB9TcE9CxMUcgyhh8A0dE7xB8ypvj39FmKZvSGX0z+qb/GeQy9SF/wycG6
2Jqh4rDG6JTmQZ8XAV0N9coYaWz6QKB0povRzWiJpwgp0iC5m97xOfQ4AVGSR5jbIjt0hDq/dlqs
O4nqHVw1xwXAUHTMXFwvqVDEzqpS23uyQpFA7h6P+egSASEy+VjUGmRNY4ISGZqttXckCcPhyuGy
cgDjHQETjtPflAz8mGWFV4lVBEgQ3Bh37n+4bIH2MqFGnMbI1C26hsUxPWFXr+xnVijoV91xmIoa
1IEC/LBhIBin1NKXwXSkLR6xtdRTGiQD7calg6mL+YibY6kMpqmo5gbUHvZV8gdEInTqOmw6NlM3
bb/fr3vCBcl3Acypjj7fQjZkAlu1nN0pSSS5zL69YR39alZ5tyV8MeKpTii4g9686I4cwie+umPc
j+mvC8zuS7tVuyJdXuNI5KRjaU74S17IbLPbFcI1riGIbQwL9UMvmF722kLVMBhhHQ/i6WjSOjyQ
cXxVmdVuLFjU0dByfcsScTWyRnU1UI4bhbTeDyOQCEHks1JLoSupskTuEUFkoU7AcBAJtLSNhQD1
xo7HdMEd1vGE1QFaveRmR3o7/m2u5+eeUchcGoaRuW+eXcSlTHCPTosFkHlkZdJteIqMnJGXUK8u
lKlSfEVLn4Wy0gNAg1n1DBODep4BWFwqtr3xLdeZTU2mDF8yH88BKZDDg70JLwljcgG44wGHw8Ip
pB1U8/dzrG+zqXi21iMmyeey1o6jH1ehFY2m5Oc2zuXbHZzL1XGCakxKbzSSQibLwjCi/H0Z8fnk
Mm4Bjej3scEnRPWklR7CT20vx3kf5m+0dxurkXSclHocMwjcSVBanM1LodSC6Nho9vwRLAWtJGqE
JSRYZWzZ2JwqjQDSiuV20Hwj33hGLKqhpZtTVYreCzRA0hHretuQRw1GxhzRNmtADhPdiW8pZenE
vg1xdfusQCKl77HbMmA85LE9Zm2JZZOnOKggLhEGJs0FCQAIAJEreQi920PnXehm8uRHHiQQIiIm
uEqCutOjjnE7tR9c0VOMSe0I5hrn7nJGeJjkC0bMvz/gKvcI+z/A4hkWPpznfUBZz4E0OBbSIivd
4vH4Jpt6QQZVSt/0GLQrYwXdPSv2tvgpJOtJxKMHjk3HuXzGfLfJQ6LK0eHX3edPeQ/kjG7Pbm2V
tUnG0KRzLio1bGUH8SqKrG3HykbZ/9mgKFabJoh8P6ztfRK+QrTdIbAsP7GZcU1h+QehOFLqnY3k
ahs4j7WkaWDjZYvbfvHcMebD9YmoZykCSnLBj+VIyAj5wv9Ta1CZR11/xL8WwvxSYRBB+aMR8m5j
C2sPGfsd2uboLI6tLCTTqEVKmhiA7JwFr5MILVwMFru0fe1q4lTYepkw7wp1rxmhh6Wyerq/mgc/
QjblWKYmKlkPISQQfU4SrifOXh3FHqO9ApbDg7CxsVtkughN7UsqRuDt51llfQ+ClN/BtW/EzKJ7
FSsIB+pgqMWnxJFUJHFrIrCpHzv3NKq0hdwULZKCxECOeobl/Rx/a5KLGNFD7sOhzAwbpxa/rc2d
QaPkCuCwVUlPb6yQR9ZU93uHUm5ab29mC+IKMd/J36GVK03ssxUJ5IwYhgzrtZQzGXsOZnbBjgrf
MqcFNquSBIe9N5jrG3LZ6PwJxtle4CyLGm7EP7IjgDRWfiwYSlgdrGMKBJqXN6N755Px7WswMJHb
BXjcE18nc91My5nQXW6Y/R5BEI5GrfXj34wi62JtVz+rOLgRriw2KJs02iJy8/5UMd8evgKR43WU
e5YzJA5whmbqw57LbF8TnedCfjD89/Bh7kwXnSHjM5NneBbnzHVInKEpGZgRaGeHR2KcaUO4giKQ
SVq8sQ1Xobw95ztsJzxRXSyPQXbXPzoI7yrL+LJSa9S+l+TyxepFqhU2fXUpb6QhzNVZjUey56LX
h2RHh1XbwlNLmH+s5Tj8mdDCJ55fPuDNFgRW0Qr2+abXodQd8e77pmCnEsWqV2U2xknSfKcOpFaD
KJCWH7fowAN19LRTYzmb3EowO3mINbHS5FoesBugtOp0PoU7YYrHYEbnDVntj/88/8y1aDI5+KBL
rbxYcUcUWTAKxnwOZdUJk8T0k52WgJ9HaV79bFaceHwiwgkfoGcBI26mhnI+lekHwpuqc73PpfOW
oxVmtoi5BY4GwScIoeGxMArn7Cmq3TuLvWakY/3VvKKPC0cBMgDPuDKSAWn+rGqw/OQa4pKPh+ko
KL7Q9nLNJk4DFwezKKjZdlOo4tRcQ54LiYXU2ynVE3hLT4KGDgPEBkL6w0NSlc30AiGYfGSw3PJ3
B+pNTVvf9rhPAnelzQ6TtMuSVr+9BxGvxUAJ63UG/oClxl8DkiaCOBy0NQCnuJ4AC2haahap/OCv
WN6UOC8Mn0qHYxtla6qzWJ31zM61KxF3qkMVC9ECS35htdP28aa1Q4KSbtq3fATINVxtEOmvBTP8
A4RRGVg3cL32JCKQc83XNPYn3WIWyTB8iNwF7vGLHx0a9eWBrX5O+nyi4Btrc8bNUXXeoh9XWNyX
NX0ykiRNcEmPJHKPURDd0tIwnR13FSQStAz6DKlP42P53NYKGBbHTMXJhDJftroPLmqWt6nDXZnQ
IKJIXCGlxGE2InWkuZPXH0jgkBJNwSMylUpvtq6BxF+WnPVAB9lXb+Xg2wDKTl4bUb4UaJU4ujq3
97Nn90kJdwDDlHpCWnPVMCu5ltnsSNa5/5rly1Zj3mGhncwUBtvSzBAoclziapbo/dmgHUE4jdQD
5fYA+LPciPpCX3zLYcXvPXMV+MMKfJSAN3QigNu26/rEZQ6merSkCTa85aEBy1kxdSYtEeRoiLGc
EzCqHKAP3Qemuuk47K3HWjOGu1DPD8xOl9CEHLXOPZftpy0HJF/A9Zy1Y2uyfOEPnNLsXPH7Ubwq
Vqg/5w+7bNb6qEYu/L/2fJTUO561uRQxt20T8t/ggl71Gdmbi55GWxH4RkbYv/LgnJCHKcfKh+Q5
aFCwSSq9HAiuSuoPNNJrJK8vNJM6peg6Or5Th8jxBR/z/r0Htjb+qsAKmF587E5aqCxohjoyp/6x
dHHEr+UQ09ZSZYWvW5FWSENFZGVo8IecXaBOkhHUBHtyMQy6mPB9CJA3KRg542u//AMp7OpV54mK
BP1XFzvrtszB58L1RJkTRRPn2VyY2AOH0NyAmxkpVyp8FH8a0wSVTwC1P+agSu3i1+iYh7Toje1S
uKeyr7r96WxKylqAdlLRE7y5Zzj3Dl9XeZHa8zi6wkugwNn1CYR35vMNqJata02eLcfGiepkImDh
iq3SivAfpe8NTqgbX6DvRBrlBypXvMHN5gtr7f0zTPL1Uw8oEkXcdq9BMzLQKP5sbPWLqgtPxZv3
XnGEObRRBjjhkv6kUUEC99RfpgbHXCWES+e4EJc3KHjyOvvygO2eTtNAnFmRlnahFlOUbJ9lo68C
5gz4kOphwgRmdktkhJ0vEwcY0tjcXNQ76Dg87+iVlQ6spqtqu4jQ07OUCefA0G/DV6S9SnOkDi7+
00417P1g0u1s7VCwkw8uDYsAvg8NuMDaRBEZKEWp60iIbTCjR26IyWRKZ9K2WnSkY4TqyxgVXrXX
Ru+vrQ9LuGXd9axtX3Utsnbo8bFFvms2nzU4GLn668KY1UPmHaDk3KVOhd1ClpeHvvsscHdkjCBw
9BsF7+lsHhnSmZIgGrFfbDz2lMznjk1Eem9sHDlw7JesN/KK5yTy/TnBFY/k47gy+S5fOkPAq6aL
BSoIz0xzk6urznI8HGxEwcZ29Myp/Hd7DkZX6q5TZWSFalkqI7rTvO4v9VTcGjZVMjIbEG0Zer6Z
AyaNHgsnNAw1F6sz+nCwt1/1jYmNAgFvn7vCorxaz2a9Ovx8y/MlZGxd0qiK9lZdvgoUHrhEnMj0
jsFTdvO4h4CpAD3zPsVzqJgaRWs2XAye3ZgJaGuTpQix6MqvhHct8EQgnQyKgQBEjsQ3lZ/jB1HQ
1463+Bum4Y438GjDJ6Pei+Qb0NDyFxpIWejr+bw79LZoPmObxWWODez3xGkIwdJYYWtNHa9+K6jU
G/EdHNviUxgKA7cl2BnTzjMRI0a4bQdO1uDP634g8RO8YYgTAxI0AUyAOc1wxUe0KlcmUBKp6DYA
xPBhxUYSzU2bZxbDOzYmG63uus6mLdEqJjFNCnuj1V6mEFRjhg6VAe72Vs+72HsB9M3HlN48qS1M
JMMPD+oilAdrRTDCr7b6kAUaJFrav1ZWsdyCoU4nq2UA7R1LSDTHd+gUYSKkRfoNVM8bZP28uTZy
dqRqwMVUcUCs7j3KjwwwnVw7yLBE7/Zx4izQ3GmIPHYAQ+pW0FuOPpA4qOUMU14bkv4XF0LaRzAN
6j8l46r/bCy7FoJ9kHGAaG5oAwLniWe0GmI3nkDfnzPmtzOnxeCoMUlOorw7ugQbI/p7sWw2GIQ4
YiT6F4cZgL+lRX04N+teMV8IsBISdxzjhBe7s6h4e0oxiBJO0nzOM1SKtMNPbD8m/J6Iqtb946mB
2s3qSrVp+dNlL042mM/dyvYjEWerTOdYYK+U2oGmTs06Wb0KrixZ5K9u8R+tFHt0FL3X74AV3dX/
v++tOfhcZ5qit9CD27nOGWOOULyM7cVO6KyNtgmcaEhCyC3YoLFf5GPol6kCzVq+1SLRRscyZf8a
Z+Dt/DV7EohVAnR2R29sBWifORdjKZeF9q/k4lywZBKqspcRxsk+h8N+KCnrDHwrpEWt4IyHo+Q4
PwTtXZInwbQzo9svNfq6KEfzQ+9GClvBuEkx9RYTN0GDP9QC9kvV81encC8HbaCxxkpWIohdlKyU
XqtHn824TY8Hw3Exk+RWGu9MtdinoMI6tbtL9VOtL2IaktXHkOHfLBQL1RE9WmLiHt4p9n0/cOJg
RGjm3Dk/5z2HywvcpB0fU1MNkCP5myEUzneg8t0900Yhk68yZFwTF7Am5U+6zD8G7KY25PEQnB44
u7QDrGznZDC5HnlF4GVbFvKPxHbGA/xWOJjBPaIUjs/SG1q3lcX+WoHv3RHEulBaN4ZS49e/7ny1
+Y1dzc/3awkDvpGOcaIlIwKZnnCszwKQz3g2aq3zb5HMdPXLKX6M0umpAVdHfFfzOySLi4qKcN+0
LmBv9pAwApViIM/arAXSqVot3DsWwuvywvy+E9smKGPH8t5u2qgz60oc1ryQlnb4uHWpaVro0JSq
uwf+kmMLmUtkyyK+2CnzkjJUPfEH30pDgqY0M3G086ypJGM44aE5mtdfh7IRC3XP6tDCa8tjMUiv
6ThnZp/FAObSV3hG9Ct+X4EIPavHnGAS7GV8WNHmxN9dYV95LDhSXFRFKIpKuIy8arF2mP7o/YcW
SDM4UVoESPjZW057hCx4rvui0845Rj8rWfXYlUuZF1hls1HP9fWX/uNvK7qcbxADLlPVnaTWGhKA
uctLyggOw5HZYNsR3XOyX4BGQn66TX+b1K4wV8N+eH3t/o1MYG1zo83acXsUdVOXbhSzdfppxfI+
HM3RlrFTXXFl8zsOIQy3gCjFUYP1D5ncA2uN3NNqGHi48dmF3feDpQfCFUzgdH1x/E+3IP+cil6r
SYsNBK7MZ7Bzgizx+7VA0B2l2PfKNs+L28vKlkzHHNyKh5U08e8kjfEomOQmEbuLxfziV+NXSh6H
VsbGB4Kv8e40UyfSmRL/KHWxLigO8a/KtKLAk+GNGuU/VFfQrfI2ougdBProDwfOy2QO16kloKaO
Ome8CqHz0phrWt1i7VUc1HFTeETYS7/f6APPb9jyvHvglaHmFhBAf6H4ewC8m5pIuFWHFB8+ORpB
B9fiieobOxIsCIwNHVbw/trmk9WW+JKhb0ebN1xTq7ReANaeZNWDR4Gk4rhFK3ph4212XVAnGjru
lxl46gPoSWXGWznB8RqsgI28WP6FfH2JVlKVMQ/xLxLKp2nsQGyfqIkPb1Cy+vbVwBM1ffHG3MLs
oHC4tVigeIkZHpLsVhb0eib8G1dqVnujEaXznGqS8cRcZrunS4gn/WnfJx2jN47j3i15O3/c7T9U
fw+Z4DpyBHSu4RD0yICrKAl2hNNWN4/HgqWxnV0T3chdAbB42lkqFiYJKsXlXFstZcbVkJyYHVj6
tu1IlbyW0/yPrJcyCuAkBJZeE981z4e/nkpBUKYZM68llesort0aXP6mOiPz2eiJe/QMM52hnXAQ
eTZfaKzTu2mTem7pa6MWj2UjTp2PU3MBDS6Eded5PPflqPDtfu4wWEcSndiFcI+HGFO8L8ELwuK4
R+/dcmno7ro0/6Vav/k+pOBUPl0JOQs9qiFMo41hciOKCiXvg3ec2RML+TwNhS25rPCMkmVPzt2n
0IYXAZChmjlMdoW7VMSq2Umj//kkrMyfoVRnW7oks1p6W5/d7N3i4fE3It3mFeOHXfnYuveJWjns
MRPTFYIoFwj6PHLWlhPlC5vSH+KR7yWLE8eK9vSTKx0f/Pq7oLEjKnD4gwK7Fshn8vmnP5trr2zR
sbGNjoNSum2+dqAFw68+5DcIUl8Binre33HXJcGAHjwMOb04d4EcSBL8C3bryLwP47xVrGaAoAtW
MWe4HyJqvTJ6cwTlXjrRqHzXTC/8sM8lRJ07HSmwpmUxfoXYzw/N4Y8GEqcjDfzFwmOzdnnsPQCL
dXy2ZxlH0wduWEeSP/roWCqRCMd+hmMR+pmdeePwpGzAdWoPuU5uz9/osuAMoz1zmw4aVn8QY3Ld
JCFKG+H/ClDeh+GMKM9SUJ/uYRskq++1GtK3pf4zJARu4ePKb1jBYyJbH0C04ZWZfSmuTfRqyo/9
R6MG3l7jwRIyvXqQxcc/7jzetbH6hWrHE5Mic8ae2Poim/734u/68Jac7LmwT2511gSueRwKhCVE
B3SHzp8pKbNHknd9cuv4zxMM8W5ruPYDdSRoksbVVeiG3HDuPeZ7LQXk5914IzxPyysTPNjpGDgt
RYM1XjMxaj9xOxRiVRTFTfpNaa8ktoIpdwJsq/UvIvy7qvMAU7YLq0WH7f2NL+fZ0Mo6F8A1UVWU
g0wy+VHphQgoB2xQBHn1IElesochcHvYJvl9aPIi448N31J5oHkvW4yhjiRr/r7myTO0lsB6NC/X
NPm2xR5psjW7twT1kODQ5lVyIFp4JCkCqAPVG4tP06oYHALhMuHSIrwATRjf1pFD/rbFUuB3Fqqi
yPZo5wUGIosAn+5nlchxD5C9XUfHO1la0ODcFJzny/sAfb/ACf5mPgHTGm0fq9iRXoUhz9zq3ODM
M2UMCJW6MgYZJhy5cDMHgba3JYzUokpcRS9m7BcFfeFOWIgfUuVKV7kKdsUCsr8FfGMBxB+Ni79X
9+ElRXErgYl2UnG9OZemhujKjUbpbW5ODdF9OUWESOPTFvOsSiDQMRNnVrn9HXW6KkzKz5r5bS1Q
1DqMnwkkDnGfgj/mVUNqzg9zPIbjFab1a0lO5+S75YHl7OkyFlyRN83yguR92ZYSSb/IQBMRIEgA
FTc2byJWJRwogjUdIiaT335Fn32bhxJ2TkTVvQN3idmxOUBxCiLXWYVBOv3A8SYFNPcwQJgQW69p
1c3SZJvSCOws+HQ7fA7JJvLW2uzF1TzUVNnijoIYeD6fRuEwZzEgFklHZ2DL1x4vLp2xP9pV0Ol2
PExQSVRXDxCVcBBAIaKJg4eycv/OZ686DN0myFnitXXQgXCsZ8gADX5S3HTLCMtMT3HdorM++Ld9
i3EH4PB+Eg17rW0nosrXCqxtLshApS0NAc1Gz7QF1iTnRLhppwy1HZHdviFCaW2php58YLlL/kbe
cL+qij4Ssur9Lkskd7O5mYbj0AxNtoYK+jWgkzk0ItQruBbck5FbgrriCY/eMYxLNXOseNnr6qwN
WgxILYy42rs+4kMIqrjhmAciZ30dB7qsNYLgTGGR+5oCrF118jntgI/r+lWsEcjvPjmeUBJlRUez
zgG44cM1yEzhOFm0ev3vy4krXrjCA2TQYxleuryA04T8L8tfYk+WECYNGo3MGxEYVh6aTYDvPPSh
Mj+DnMGPyY6yHsLXAwddnFUeI6txRg8cBGOOxgUjzefBwZNzpE1HvYplNRp8hG8hKBN+MAnecvTB
Qk7WdjNJqFFwByScRhFY7dHZkPqMjtHLOOn8MXwBiHJs6siJxLYsGJ49jknb+3bJD9mmRhXsIRWO
Q0K4hTt9A9KXeGxLubUPK2X4UOpAHInYHKtzbUvkOIkqXpqvQSng90rsVw628paxLXLaoHWMnGQe
YlGs9S7tlpBAcoe2PYnelUxmv4a2UU0JjjVOabQXH4e0JFTbkIpCcGETsEJGLbeoG04N112Eo2+I
dJ/5qu4FId7DDAGtsKFH6cMCCdiQLZ6Yzg2ve5TEqlOprNMdNFIX15AktC5iGu0XYgzd/SQTYIps
zyWqoLCy8hOLqC5Fb4T7Pok8T5uYUMETe1OWR10dp2u85w8AA3EEQLbwgTLJgF/r4nRNv3xGgNHI
eB7apJyaeLmc47kpm7zgEZTuj5c7mLIUNeOmwktwLc9/myi9fWQ/F8LLbnoJCKsT7ngQcujUuWdq
22ewaeA2Ea7V2DqssA13O6qE/hMFd1Il+DFAglWV+hWDPvSE0L65xEejg8owSMasrxlWnP8U9GB3
yCh4g99HUFOo9nNxmD5y2LxfHXfELE2OcV5Ga2YtM/1hMLWthB/gJTu1UxZ3VZf+BQjN23V+hF+V
sftru71ia4UyIclmSdQh/L+2lPhd/RvKdfnu700WswQXX4I7uo40GB8fBfbKHEQoF2do33qnEoV6
UYGJcMdSQCKkTZEVtPYXmoJH1SWq5OMsC1fl6+KqkSlsyf5lPm7yBJk8CSj6pQu9yFqpQ3ha2M7B
AZDTJMNUO09tr+pTcGnJdh19RaKIAEJDT5Zm9ktM8W+AIku86GTuc7m1MebFXrr/LoPDe1szLgcr
Us/y5TgJuFyTBlf2mTIkFbGxEf4ZTZEJzfWkKZecxykXi8JyUm1YDk3aVQ2eZDrToY9SJis3SgGV
tAq84UL4HtvpPYiNfolMuyXW31wFNeQBLHysV24cr5ciTwqmVAIydcX7+f/bVAMYlrsEN/E+1D9W
H1NVAiAcTepCMOYXxQb9caC/4MPBLQrGd5MxRmBrjv2Dz28IgZY7r6iVYNAlhObBmPHOYmqLukAS
J3JBnXYGfDYeBnvEMTkoPrS7w6XvZVjdSgknDrkPFf/5ow1M9TSwxwBytaQ3ZXZZ7VokyIygLDCS
fw4mIsuYKpZoxlVrJ5ui9zU7303m/+fsBbklAiyGIy2nFWrEX6y9BQxSMF2PjHY+R2C1ux4WBqWh
d71Uz346yH5dBP4daaQ1UlyUJ/ZGXY7wkZzil2YWj1G7z0jq4VPnjZYPiWDcO4iQEfi9PP/SYUz5
bnz8TnvFGcNkOAb7Wlor7rzlwp196wX3joaACNVBYNSmH6cckexaizOxAe4vyUIryNRTHqc6pOKZ
zYJKAaiAKQwEqw+Od0Fla3IWiNw1xAASmW6mTO9z9Ql/HbTKVJhCsnBLy+HsLllJorGmRDUeVPR4
ZLxITiJqBiB9Ll4GrHFHPDkEs3ZW54ywKDBiaVyt0QRnFCrZdjTYyMkiS+rgf/7PjBd0VrPjijPO
AbULAmmpu4pvNv4IduPAXNTV0rsmRIjcPL91CXLbaMASE9kZl5oCUIdjRiPn/RFVdmQ2nmDipa9k
D8e4TIOMQfkvGQGe8lFrarBYdmOL3gPVcZEJvyUy8X2Pv54PSKDyZ/ZjJPzkURkInemXRSZ/GpSG
M9B+VCW0T89QSVv0fte69z7ZEnsDF8H/5Dt9D9lyTEsmv98Tz7GuF2PanscJ7CshdTCjdg9XYcGX
IhCIzLhE/5Kb5aYtEa8Lcq5Fk0hoB/FHfXzhh9gmWKWiJfyVdRQ+GqoCmSpM4e47A7KQIqrD1prj
KJZvb2Ar0v8InhHtqnsVKvDKD21RWoDepUYNGWFBn7d+y8C6wAagoGbsQ1KfThBm5ZD/Za8ekitG
R4iy/ATeXB4vFbq5t4QsFpT2Z2SAQjcG3sGBLiii6njAGLCA01GRZ9+MQgUonic4qYuQe+sx13nu
7uC6WNAtNsAUDe5PME7WtLvnJVGK8hqCeqqn9oUXwkk/uvIAst7mo/NhomSF+TIaB7gp60zKinKT
Wb2+3lBA6ohyptQV0ICXAPLZT2eXS+970R5xQHTjCPP+tSB6n/m00rtn5vfjJVk4LeYCbtqpXg0X
kTqOhCWzg9w7XIbM34s++QEVY8iKzCcuwKFB8KaiY9vPc3qHR43+s3fo4aMyiZduO3D+WtS6TphN
toG3GrMMa7vck3W1W/R0omMVlbq1+vr8CmyZ+JSEpiCAbfoXljtRET+HcEtfW8AAVGhfPzpXnCGd
UWQJr4lIQBVga1ucTlaRDf7HUWzXOeloCQnQmxgI0qIfTZCWfIBkBZ1DR4hYq4gmRbWMI3KMOLih
WV7hpFGr9Aj+32gIH0Amto5eD1jm4dLMhxFg5r0RT4Tjiu/8eT0xT/Incyl1/cFSpeUQT0IUbSY1
uxGSXHsbUYCwUV9bRElQaPF0AmBzYdnjjBSsgpjro7T9lu++seAeoSWy2aGRVoELFTm+4DjwQmzz
GasRAugsWa6ks7krtDrreClFQqdI3sEMi3iQW8VAotl8BX5aOed7ZGR+38qegvbm8Q5okbou7rR4
vpAutYHVDnMwpRdywHnU7lLEOqOm5pkhNwRamZO9FSMagQURPWzc51c597XO4LCrMO4YDUijL27N
Cz46wBhtgTukaIqQujzR6/64PdVRqA/ZcYevXPjub1PNb7ll+/TqCJCTAM9hbbk4xVovaH0glKMp
CvbhG4HnK8v4lJSoR9FCH+I9QDJyAjs+jdHa2ka6JjhK919EYs9JMCol3UPbviA/N+mmMRmSWrng
QqcXZVMznE3BbJGY8vFoGbkifr5BRs/pJSI6965D1CzbXacubnGb3ZZZLAUkhlkOufYzt0ZOrntF
YT5Qwps65krpFIDMcayQtHqdVZZ/i95/1b/9yKplR8tfrHZNJdxP9YRaxkubLpY0XuYvkuy8al60
bm9zQijoF7SN92qW7OB4940dpFd+MXFOlpDDVYH/lVRitsSid0xCR//7nPHeTnixYnRyn/C1BJRx
6wJddeOte7fdyeehaRKrnwtxiT9nayOKenxMHyQydEvFwRb2VkloyapW+jD5BKxhZrvaMZot9ixz
YG0Af9Yl42QAGxmWnz+Bo/fjG/zTxipPKdRW2dEJf0xE8JPs8QvHd6p/hx8Uilf8ccbfM/pSgtph
cJOy0ogzq9T0L+3OCqIRLQAIEbVXZSzXt1abTcOnDJ5RYVmbrytO9QQlJNg+lZ0WW8boEBYFd386
JCYGgcrzohmsX86f7GI0wcmk/kCGNI5DDdXwzhj2HuNtzyDOqrDBVOKbhREGbHkAYWUSbscSDdbY
Xi+KN1nI/m7Hw3NUaKxUyczOHIM+PVUC3cBIdeoHpinJU7bAP/LOwrgPgnx3F+lAr9vkjnUGbiEl
lEywTl6UWTuP0w04zNbNHqHXdZoogWPjcTw8vlIK0HnmnAqeYSheXsxF8HJE0Q2p4lTMbpOiojUS
dISI6w5J3emwHbiLxsqt4W7UnrlqN785effpaNuPDdGfXN9iOl5TR6h4p59XH5NiYIinlJyzh/fi
2J1M53S6ZuzlqaorV+tfozQJuYhtIkzGhPX8tVtkGSLcbTYA4l6REZYPwF87UVfSyz7uBoLk8zLF
Jw0Yq4voTu9/THACYyShttVCyS8TJzrV2bGfv0JHkhWjNm53BZHCqoCJcmJr/MVwS1wVL8tDV5Y4
HAsE1+QTZMnY18KhwXWjyk1cXDaewCI+ijZIemb0hNGQ/hEdQvu0TjRsJj6u9Bx8eQAd4MLdKbTp
LuviB1gwXoHXiWge3a/GugE7Diq6A3RuqVjcAk65qSdSyWfFra4CbuviWdPYPJzb2tPnsnca7yDa
CRvIhfBJKvX6O/1a1Xs95K7gh3ayRSPKXrGNRTqOvTn+YoB5nb+31ZMi86ZswP2Dnm+ahFcOx/i0
TlD0hco4lZQf/dnI31YoCD0lOLbsjKzpy53b+x4PMtGPXWJWsG4LyFPNY0yYEy5Jm6sq7QeBTV8J
Ho8fhi5bMq131aD8rEaJVKhFfHrNu2pcFDlmaE7JBmfjuarhtWRXohUDGkSrej6YHrynbloAr5OD
NqDID7ka0sNvQZwwRGvnWTiITT0hN8Abbw5RrKv/L8YtIkJhuYkyyrI83bFd7IZzIUjCib9mGHq0
a29A+klYbrasJ31uPep5ToMuUJZs7guiMmAA10lk/4ozW0UmOprjFFm/dFfvuCpeWqV9JTLxGCXc
wXxnS//efzupgdN/jK50Rc2zGSU9bamvdFbl1FMAslmEzpmWin8F09e1j5edNvCdZywNKbXDI7G8
7ySPHXOtrctnu8IzysiEiICw9ukztK5oKnv15u2S0diD4dxxNvB8MaQqez6dmh7NWLzlNf9VLi8i
QFguKeMXMYyDZC+CYFshJ2TBxkZwLIUR3scLsEdaBD3oCvSxflDRLhFWBCDy2RkXyANoasv5wt2y
j+WJMxZ7uoBDUkYImjv0x54NU6SSMSJRyHt4JCfzYxeDlx8kHoutnGqZr82wEomrMADll5VQIiCf
C7pmokCs33Mblc8inhmUZG27zEEFbEfRwpRnMTqe03BQHRJp6WCwsJU8Y0xyVjgwnhDUQ3gf83xm
xX7w5ojNa7FhJQaK72eCqOB+sejA2RGNGaweCL6aEpqCCOKAhDX76rNsU5Wty4/O0XGH8lV4rqxb
t8G2NGHGrhh94hA419DmRkzAfiA48HZsC4A0uHmLcy+sEmcGp9BGOrq5CBVGkYCX75LgwrpiUZJF
ng2ZA+OzVsjGjLI6xuK5QryLAxbiGND7dagi/geUab3yqjEzaZsPGNcosY4RTuG5cjV+r71eHPwB
8Of9qmdnHFzNQKkLWCvKdFYg6sE+o/Myzw5tFsPh9bjtx5tlpFQ73IxE3Wmh1FMWGSPeXd/r4qmT
pIb/gjr4mwZn4XUdhjpzNoT4b1aq5tfCgOVoL/CdfVtoBuuOuJ8NV0A+ASaiPRv6Rbox1sCklQHr
o7o/D/MC/6NDpdd5rkRn9SJr5gljJfRiGopJOCLQLcnVDE2T5WRK1iU5frgfkOoRaUD6+gyZ4pmk
gn/Voxq4BYpDIL/sCDyqkkzRNFCraKA9l072FZ2JU7Xv7Te0rrFn5ZfbFxeMGrf2Iv/WRjQtRZON
wTdll1illHjSaOIp7uCerBNMMbrLZ2CA+1ZMT8uS5F9sFebXFwGIr+XuLsoAjtPhYpzK/6WEalrs
3lYj1gzDVCKjdZK1PsdH4r1JNXcVuSTcrOPLQcw3UyXS5LEmnls6aMNlq8iy4Tk2uDELC/Cdj7Sc
EVA328YAvulAy3AK3bEHNrkUdAY+NZ+5/Roxj0gUXmgoRh6ZBiGh2ZjYXym1bxUFSb35GNGmnNHW
Kf59iLcvexouMyxusBcVLLQus0wHssuMrHv2Buck+niHJj4+aCBdNTaN3YwxvO84JuWPeXi6wY0X
D1YO08AZx8oZs/iAt6oou68cqx5MgYz6A362cSODaCoG0cM1CEBlQ+both8UwK89PX3uHPFi+raN
Ra2BY71MImqxk9QXhXFJfPwO1gp0yTuuMCoZxmRXHRcRp8yFTa3DokGSJFcKP/UcLZOh/w3rUSrH
I8gKG8cGJhVfQHIVnX5Xp0GKgZsZmREr7Y42YJU/8rhqAnYoBcwEsh58a04GJ7ooWclAVYVlVCMx
M/MdblEbYsOGNwaUc6eP6vXZOANGWHWfvDH0RqBy/RxgYDNHE4MEl+7hjQn3XDLVEcPOyfW2t9r+
Iq8znU0aYa/qpQCMysRJesMhXGdxNZk8NCLUbLmSX/nkkYpYJjiZIj0+jwksspVpLo6S/g5Fotmh
xgQ5YX5yDOFzizfz0HsOaY3+xd6NUW8lLOGvkROKguYEloRtBfE9DpVdM5NrKkOzLR78oBxOp2E8
Zb7Mom4RnvvpTQhwaXKL7aUDXt6SubTifVL2BU1vhna9c9wdcIu3S6Z7Y+SioipKaL3jua4JVdkE
YHfS2pWfyX/koYRx46q2JRESkiML6JE5cby5ynA1OXDmms2UHIXS7Yn0NxrDyeGEuUdRPeXHmFeB
x2iEqkgBfA7Ca3Jnc5RKfLeYSlt0oqrTczs2GRLxpAAQ2dOmH6s3CqH6eiQ5zeNJ7nDMsah7yabq
vaFknUaFy83eb6Tqk+0jQBngQwnRXubjr4P/yom2py3QAR7YEZt8WXmcZvuUUKrhmqqrwxVnMAUr
YHC8+kHyiYJ39GPM8zV6FV/QUNZDTkf2kaJ9DQFLyhAVEvF22kRZ7SuMBNlQODMzxUwi9AqyZpcY
DwUBkqIeaRpd3qbDUU0V9AXO1d6a5ParBRMsVSgYyvenJbxiyIDqW8eK9nSJWrdqc4edASNtOh18
2p50YEnknLkkiRHn6E86j8iDTTThBRN3mzSkxGZRM3D1FCIeBbAToS5cO4bcpC6Pn666u5rs9y5J
5gu+T8bmGvxaYXiDirP75OjRsCRzHXXTAlzH7zaPMPxaBNJ8JUgGJPT0xKQdkPJDQp1nb1T5CLyB
t3J7Jaw53DVE3io6ogJ5YZ8szhRlBKtcCCgJnE32qBJHGRaC/k+wW72w8rkTxg4y4YIB32baFYlS
wvthZDGGpfCy5TNLy2fk+iJQFrt5kp80QX1kcBjE8JwlFWiXUVkXTb84wxDvgGaeUvaYSyL5DB3E
IM4OImYVqMt7WE9lvALGU86ANiFZ6SigBXEs2OfeSEpuVKDh+5S58idYNhjlLgjRxMym0pnLi6bj
Iai5fh8OGLM14H93fpOCO8fNy/+PxnpKoE5qw5UZ2xzUx9ix+Mz+FbGQxJ/y3392TnvX6Trc8Zay
H/QVehg7BfPPlooGcWJnX4/yQR7qYOUrqHy4XOGgBYk6nIXGGeZSZ07fM8rnzd4PsOU7Uvh/FWKb
5AlVmIkG2swTyNeg4UuSFbWLoF5cQywyAT5Sa1eRoKrT9Lt4+4FBi9H/ydsdh1z5JxO1TyZt4mb4
zPNtMQGYirf0KAElug7/07Z3wQej95Na/iTA2BpgfQyPGUFQtC3wr3LnlAzihuU7xzaRoIK8zL/O
gaXVKvUWwptzyrlcb4mWoljlqSrEH9UwMezc5mHMLE/OL4HwOr6tNJO6ipY11M5GM7TJGhxhIQum
HS/ljqTuapW0C95E97By8jW93l82qiFmhh4sxvIDu1aUvsSk7fAVw2pmB0Cezfh8sTm89mzz5fMK
e8C9wzK4qpk+uOrXup2NAAk4Alqk0R7uYWshUknndqNm/ZHUfKhZ36A8s4DhVo2EfpnN4Nh4C+Wu
EC++5O3rZm5R92UBZ/3Jt5BQoUHkK5DlhV28rm3Cmn+VW0bZTVWvJ88FOs35r5l91oZv1BFboY2H
vnsIJ0dVv64L4dG6wI1FpGf82tsJH1Ymdgyvw6/JxIcWcpNUWRB8zgHnLSkk0BRU4ehyOnvkFFc1
ONS5vS1G+rmcCbPeJFxOvfjPtlZSBeisKxiD2qZfLb60RPtY3nFbchUzCg1Nhg4WYUkEUMT7B/dk
MyfKDiZ/udAhsFuI3P8ut9j0Fy0vhk3SZ4bZsgQeX4tkD5ILpQoydgeIup2nAKfYMlEKjWCJNoWz
sJWodehqTj1BimMK850c4/1NS1sYUuXcFbxvNuLF9SkzcRDkx7ISqhFq+WKDMPHixpFuLg6RgxjS
zHgrxIhx/Ak0SQOCK64+p4BvfmjWhhPv2OZk5xCRrICY5pWnzv5KEBdiusoEjfol7AZk6bC9UfuL
axLXmB+NkdRomN3Q2l09l6CO9BfqwbAhPcjGx2ImYYZ5LzjA2ZuSFguBqfHkPsNonvR/fUHwgjlA
vrI7QpZMGqrpWGRM9c+1kaCWy3bWNZXAJpWQBSdAhCWoVuf1YELE1To6tIvy7+iOYn2gN3e5rHI1
goznhbKeMxWIYJftfPjQlwLQa4x+VB9xJSyDde3aBRD0TTE1JtQNoJ3PKMH/JcOaXOozzQAhNW2R
HGIEHxBS3iPNxACIc7vxYAvhmG21PXISv1Auq0Li1oZXvxKOG5zznJgZ1I79qBhGogmieBFgEz7F
ByUOHvxFnahRNtTGb6MHs1GyK90GdRHsysiDi6Rqj1lkwY+ooAH1HxoXnLd3xEbZyoiRl89TVB76
MkPYeJt/gZ8aThU8BJoI7nLvAEnhrd2QSgcCCgv28TBl3cp3wpFjuV/Njk1Alpc9zNCyVGgjJ28w
V7KvxdJTXwZQLn4Dp9TMPMRoXOg6S+W3jv+B5JAn4AH8zqhE62ZzZ82AsuXINt9TZ+x9cXzA2QIO
wQEp6EPJ2XtQXn62UfEzXjmu68xXz5tH8+NCeNHklNweB8bg/T8vrHhjvu5S0GbsWvW2X7MQmvxY
2cBsnXVq/LLR8+QvQ99rK9qCrp2a17SrE7aVWUjZrL8vyR+FpDW7ILKwM6lfDMGXlwqsoP3gCUd4
mVmH5gkPRQ234NLOMtEsbuiT0HjZnr0beC+Exi1zivYo2XqhxWW6uCgzIsK/iqgs61VvWojb/Pb6
lz1oA8H8iL0mAM4HbSdIxYXtRba6HAVc1kNk8YTX+KHM5gih6y5RfWjJr4+eXv6qbt2WiEpRVqRW
hsn8PqZAn1XM7BTCvFbz3yB0kzkFDkCThJmm48z/QywyZ2gcm2cDxfLuQcmrWwA4RbVAaz2/JFlS
2ycqUIyMimDo6QSYVQ/DjJHLi2jEKbW+KicwRXqBdpMonZX0BLt+bVLM1nTHdeV/TZ8VjIiudVni
G+ktzsbYrOqanr3j3zEfGsG26pRcWcokvPVgWeeA5c9rfl6dQyrKLnfQFMUEUKJvfut2S7Lo4/hY
wf072jh4bksnyUd7ENIA8DBY8MLCyqe+dvW9i6DuiLwHHRY5jm9KHTzdGutIQrrE3CI2jWRx14Nr
U0i71rATTnlzcJAl31XWYE5B7FzxJ7SINbxFAmqRTmkEvGcYYKTe/+GHeiVM7WHys3mRt958q0Au
o0E0WXVnuULhCCtRLZ8EngKdUIoXnGpiyMpF0xEFWT4B6Y28TVTrUmOMLWGAi02gwAfVW+fbVgoo
FxMAsgTeEbny61vQcVxXaZDY9eE539rSpjJG1Iyhl33ZZQtIhhXlG14zDzzSMsp90xUyNW5pDlBo
WslTV0aTZo1y6dA3GIFK3FkXqGoMlSnZ1FmwBZGPjF34E1tIsr+vB3cuiNoT8yF3umqpI4QPvUJO
MNP0d45pOjW3C84BGkcW2NrUr0agUkEGZVmoC0/txKPUyBVoryoq/MHq72cdmDOwB3lYyCvgq9mX
u2X0HWDbD+F3kEKZn23rQiOaCzAIeNfv6xpbIrcnGUY+tXYVJVlNYXxKCDov4HTLV8/UCQdPV4Cs
IIe94cBVJS6x+ozd/9b615o4fSjL8jPU8rIYDOrxZ0fI5D+MtY8ysp7vMRNigS+w6rYItJVEstWu
/Z06K+ycRhYR+Riz3Yyhjtdab4+hshUMCIQ7LuMJRsQpd865svqfBGXzZNAgl9t3NxLPnU9YDAIm
ArKDvuhdVQMr7Iq0XCpXfdWsRKKbQlTnHDHMbpx/h+U67iUdMoWxpjCo/LUiRyHn/1qLOkV3yGXT
KuET814u66Mb+CwsVCTg5pFgvj8uXDOzMU63arBsq48oC6ENEKdfQOkSPaodAQ0PEo27dNiB1Iz1
yx3vhzxi0isg1HR8b2RcbU8YE+SqiBQ2uuapbzk5BJzOuE0GyECWYnUV1B6AnCsu7RX0kySgTful
rU/5YYY1uDYN+63rGYvz/ATBJU1ze/0WHB9Te+3AchT5/4AIOiUnLRIHWcxiU2h0UAdkayUf8UKI
dAKvVfkhuN5fzbE92VV6EsDQW33Il/ciObvDzUX3+2BiHnxOqqqlkDUQ2VIxG30RZcNXnxtxeb7n
6fPIPQqcJOwnEFeOCYVYiniia3RYWp2j6HDaSXm2aJ3RGqN9wCNboK7YUsomsiCeZWzwnz0UiZP8
sH1bJY5rTSWYlONTXXIratpJipYRRnbQJYNEY13eNxCGebHWFx/dgZGEbCaGV+nc30FoFY9yMhg2
h0wPmwm4KIMzIxT5pMqti2uiCqo9vYife4kbBXoXUb5NMBvVqsbAXISuOtnN26Fo8cAt74rLiyjN
+oHcM8LBkBWvv4PjtE7/dfizQcbbGv7T0M6WLiNPAABNO3vRqjFsaTmKUqad+jqYbT01jhHI4J4Q
pycyfks63ul2FBNj97MI0/P0W3nKHze4EY6H57PbLjB3wnmw7yExjs/KbccLy8HZ9XsWEaAnUGCg
AsYexjspNdAXglj8l+55y/qQbAugiMwJBg8jgLfhxa2bTI2CoKb6X4F4Qe5vnQP1h2lc6+GQK62p
+Gks0yNb7MU6k2C9VTjh/1MwXRKS70e/Ft5Bcf4yNpiTNX+00JereE9qUMAjDS6rPgutTZHQUkNi
BRw6fff3P8kPjiHQrceq0hhvgnxv0JRdZrnABz/CaIhlwl2lzmRO53MLAmocTjglhbQJV6a7yiz/
TFv3UwEE/hQyPrgi4umcRwLHYvubugr7eSi9iItHfKtN/p4zWqP3R4Ajz+v3gwNr21al7APf699T
RziALtD68TgZ3jZqZHvnmy62GzM+3mHisWLXlDkbmXOdY2oyBCZ6QTPKEzVFR386BHPaLwYlUH4i
OjHjulkdo0IZyb0QLkK1eEIdk+k6Z7TXT13CA8LikS4QVnGQEhYfjuBqkB55Jr2VppcEpxvDbmZd
WsBH2TUZDri/+JqGDMl/kXrYX+KqJFLWZOd3rt/mXoYewcujLVMZlXRe918evqEXFdEpyLM98yAp
439kpB66K1ndzwNSKuLHBlOITWVgXLdY1hp0O3UQksLI44AIg5BgzURJd1SDimONK38Mqh5jBw9V
9An77LlQOOILfvUuvhw693DofdVkiwD4NbBV7bWP1LBBLGA5x8e4uxld3yzhNDwwBydSlEX6Wk1T
ak1KM8SkOQ2NbMHO3uawnwTriZIfkbBh426rr09HHlnR8IwWZQDahpO1Yc8sgehpUkMLVBBRQskK
wsl+Exjw6x2fbK8KZZoo8VIVVFLt505cFT7oL+m50HRv/kg2YZ2DIQBTFbGzccGA7g8POQI9mtLH
TDInrwnQuVBGogPK40A2rUK23M4LBZCuPX4eUHMT8XL3Cfj8pi59WjZMXxQA/ES3MROU2yQzrLiK
6ZeC5o4PjGaxCVx0V0J6exRwF/CZkxjo4LXOATGRdug3pqE1v0lMbuhcCPI1Lvyb1pPMBS4+YHzP
Ck+Cd/xEBN9qiTar8w0o4RqKLj02HuNWwWGDHDuRb+hP953m2xAt7FEz/a4aL2IeohO1GFAidljQ
H/FRVwUKm06Tkci8Ye/GboHNeke2luiXDevYEXCasVNWXvyGGFo9h0KBmPly8/nA0Pe/NxWoTjbw
fQ0eILV1ilL0ZoHvVlW3hh/jIeHsctGNw9Y7GHqFB3ct0/S4T69OMoVartXEEueEWv6sV4CizFzo
r0FcCSYltP9WwNoo8/9VCvEhoevJ0dw0uzEczjnw6BvgEWhjMKn0JY+dD3i4fedHLSky3yKmUAzp
I0Zd3Pbb//yeQyOI/AxkVhVLe8CDxVpW3qce2wvey4/gwXzjwfZaMR86kG5emEM13RSfg7I2H5Mr
kukv2Xyoh6umC3Vup0I2jeRH0mvXVlAnqWKfdCSIqkb2Q1CxrQMRLFgNYFSKCqhHBQ3E46ZCQfyk
wWlnwSdtveOVeHJKyinScijylmZrxuxK5rZW5TW5H+W3kVbsvcGTQRgCvMPHi8DTKCJbgKGnwETL
5fMrGH0KYcv5XllAe+UWNOY+j25HD2Xk9RmSxhFzGsNYaYVxSreYpjyYSVU6aMf7o0jsv8Vvmkih
HiKJ7okDQDhhweDq6Rj0febmoFDrOSoO60A0/Zrm9ILY9EIl2uf5zF98Yc5TYljlqUM0uhfyOZE4
8cx3WxBxewdIztqRyXGgWlqXZ7CxX4Z6lNKYSgQiMNSpjrERKxExcMIiGM5Ug4v5oWrZCFFegCIC
zLT9Myus06wPgK9syMPZ0URW/effJWMSakmDjHh7V7NK5J+snlPKjCwwUj+Pn2iwuF51ZKh8DkhA
T0cIpKOsDRkh0GYQnE/C4WrJi8/X6dodPiaVO0abEhaewrWUk/nY+pQ/OTmX4VoukLnisZuQ9KN/
u71rFeVcMK782S3gIfRIh6Nl3EgnUYCDykBPygjBKEOhgNaC5o7XOJlxU6HK/cMuygFkcJDJL0to
wzUgv3BOHfW2JMBh010xPvQ4gLBp6nmvaj9vT5yPNhodMHhRxHgXmMAWBGBL0nyHkMs0loHwaIYN
8sVV2AhtbIfWOD0e6erF2oMliWgUfUg1gx9OAuCvKdG0O2nkOgkpNfWIQoVix+alop2lvhpO5PNR
87lWi1S7fk2E1L7gFxeadkx+aRsAcRjzUYYgevI7I4nodSv5TTWHjJwamo3WL9nl5sKxTQXQhAB4
XaPys6MmEcK49dn54TbQng4cZ+v5uUsYENsw7nj88sydHRsrRAxTslGjBxW3FL+5INci529LyMP2
t9/d65FqrsAe4dMpCMg9JyG65FiI4omBQq/TvEAKQN63nDQ5rXVrVAlmCf/mvTgivwVt+F0W34XC
Od0eQd9hwB8GVwVeYLoxLr3rCe0FDUZujbS18m2McUL2uJTGyAcFb/e62AaMdm8az7RZAtMUso33
/oTqUi4G+P6mLk+UifebB9H2FiIBwUiQlIcWOFZa8mkQkM5WQAH51FPU8C0Yia1zVvAmyWNZcSEd
VPC2BgUDgdvIsgLLJoy9vvrz/+E6Mah2kbDyr6oIzEAEUJRW/aOpGMmgTM3Ul7ntBghhWG69fnM1
siXFWy+dVpPQpytXjOmaC5NDD3ecESJFTaUPDdL7HkOBnX0I4MrSzNXT/ahuZFnzVATmj/8ICRC6
rHsJX8r7/vdsOQa6HqoFam8xZphwy6130e6rJN7/7VRtywPd5SHEMMd4o5tHbUTJwKPuCcg6OZIk
4l6DT7ZKY5XO9KQAVA2hGWS6ddMaGjfeedVSgI6DkRA9QiFij0GUeZOZz+prlSdBwhlToC2zyOUI
xbjmdbqiMjkk4JMcLACVPKZNOVNQ5Uk2QYB8Xas8Qw/t9zRivTjjCrTDMQYXjSaSuYh7aEFag5MI
otswQG52lYWhJb0LuAnPN6py9QNb192lJ04/jXJYR1JspWFtDBzpseKQhzvrsd2xo3GCT8m5XyPR
XMTXYJYGYvBRvaDAWiIuA53QzIEaKqBBNUKgX7CmOy40BBpWu0K/87ijef8P+Av/R5M0NWHzERoq
YPwCeCRs06uNk8aQv92TIn+lkkLpGuwOciXCm1YgZ7mflmgTvkZgY2kcw0oZeKefXTp1t5oj3WxJ
UlkGq6M4hdntzG8CFoDIXHCFyKaoLbXgCtKvhCvfmhIeAICO9wlx7BF3v8NQbdzyoJP9zx0jLnrW
9bPWtqqYqc75UpsVeMQwEBy1cS9RS9mm36iHBkIeqjcSObCLeJnFElhzN4pRkp7qMwQMFEKLx8ru
3VeGBK9/KzcyvOdBspPl073jvDe2YecNb96tGJoVyg1E96mKZe50JbADr72HM8MkkCubJOMxQkfd
i+lBfAkYLE3TxEkZrJ/5pIAaxuSahujyajhw1k+oVf9jL6ZwubSkvASWCKi2DmMgZIZ1OGkV6dCd
o3+fIGTMwccd6UMKjNGCfFxI0JtAHp5/uVEODcFyUMgBXoFQf4j0tgZl7BB4eMRyA0QjtPh8ZekP
CRw4grcQdFyzV+AHwCDZphSQju8xMVcRXNMXV0swcgxs4E/wqtutz3qNiCp4GW4QCv2DEQ1VnrPI
wORGsrYntrEUrPZ31StQZBJlZkpoJk27l1Uroga3Q0PftRjuY6kS9sdxvAsV+Pr6ZeuDrdjoOobp
ipeCxN8YwFaIxeSRgxI4kedw1pLp/LbAItJJ87UTHX7fqQTzmhK4bEs9UiOJ5GKdN2c39iKkipCm
g+nmhBcevLzka/bKv41MZPuuG/C0d0cZLNjYmio5vXs4b6A4GHs9ZDLsbumNjtiMtq2v2bqqZC/L
IYEf6dfKw69Foc3Ro+otJFM2wZGcI0r534rCDTMnd7GN+m8TWV+PSdyl5Cfq+KqgQFGtpGbHaZrA
7VDxeNrJu24cqMxXs6I6obWfKECXY7qkmQIvkAvnvi6tenUerJA8hf3tavnn2k6yl6ZGlu5St+Z6
daARy7fTum5h7wNwJSYDlqGLiCsWdoS1EsPQ2YQlaHoRDHxJJZUFrpu5LoiXSx0BT3baNNAxQUwK
oDOtYpt/TxM8z0otVKXRjwQe9MPBYq5r+6vsl/nR9K5vel7YvdA2JbNAPArVxqyuwbuWT89ddTg+
x6HywhvI/870Wr2oMoDnXqHb6NM/RfIBale6qNK0zKjkaNvMNTtt+InLNcpgi9IptGyEKeGatNRy
Uff/mzfH3xzXnejeeHpfyQEyDS9ZmWzrsbvv2mUmBe/5TbKzbtARgm2nH3rvHBAsjLVtpdPRcurj
tean0/TiAmQFqML7WnKpEZtodcV4P8Ga8rOFh+9rXh6yuzdqa0I0txabhSixwmJWPj/r5lk8LlML
Ry5N+nDg4Lj95VtkuI0MNWhzZDXGAigcsvHAw00UjCb+aD7bGVvZWXia+hZI9oY520X68D5qmJIB
ivkcYXhHYhuNkuU62VuNUk6wt3nRdUXUlpiVAvM9sgm6sXm098pHZICfJIocebtfs1Vf7rzQwN3s
UMh0HrGS9GOpoxPYOvR/z5rCrpJX93e7wEiYtDflAPUAPuIMkmsMgRGVJHyrcxw1pJgrZBvH25zY
1VFEHhiELfadIOFwAgBIrxOobkkLiiQblY4Jhehot0CAysj9lCdckBVb8NyGE8K3N7JpInSn0HQP
sKSlVQeqFr/0J84yfcU65PF0IGo/um7xs1/1JnRHupthLWWYAaoLmuLc+vpyij9KfO7ebeBf8OvO
wW6Mcv9U1VQUpSRmoMVqd3403/3IQbvo9OsWVlW1XRkisx3o38VANMsoLPyUq4+ioYheC7b1EEFU
bQfLylvmKHW1llSa2n/0mzNqk1kSlLODT7IdBtkl3WuyPuZDz2/wpc0iYIRwzJH54y0S3gOEckoS
KETPXm0uPui2CzBw5nlGGUPKkYDg59CsgAPgFfR0x71TredBiyqBmLApaJYcALAO2sQTeUUZQTmq
xDjtK2ZgmWMbW10uwVNq4fQikfIR2yWW7qbdLTqizyKwYvzstcWd9V2D0gdonsDby9VA2hWqkIea
yU4pAgTYV+dEM3UNI5YMqpMyUDVfe9VV1/k4d4XQBNv3pApuCfs8tMtVAJ6d0gjyNBT+4LsTBjwY
ibK0QEMyIAvFLph7J2qqZxiBtkMZ9nEdOZjhaKwxHblYXFdvCRf0QBCBYROEdSSn8f7bMPuvWPHY
YsT3Uk19vKUmttQz41ududxz0C3MyL1NJD18eaC7qBsjwp5aR4FNdy1Ci1lvm7Gn3ZUprdSZ0EuX
1wf4PZBPkjRhUZt+HR7ZKWMDPk7nPuyM4PR7+S3pD7Syv6hLozT68zdrDvlf4mfBE0ooIyFDItOI
etM/gP8M5AYtxzxJpg/SeWz3KErHAo7vV2BJeKQiLp6YHLOj5VmW/vZbU+AIvMosbmEB3qSys89X
3V4zK5XTZDfqXRsCKEHSUEwEWJra/uyPIRhaEffZ/DLOdOdqd9/WFi1eSgrqzVFCdQ1LYVybli7t
vkNZEkBF9U4a3zbGEbAt22Rv+s0PnDjLdB2PbjmTPWlSBKrbj6N/c4+45v82ZNL8U8kzMCTuufP3
bMooxK4Q2xD+tPnlek+zbRcB2F7OTUjmNUewGEGxgD4ofq6dFQkgKxINdihTQ8+E7xtZX4yUS13r
zuqntbOjwiROHaeeXlPM0JF8ZpVZ0MdVCjY9C6zLQwLkSdxzivtjwYGh24/ezv2IkpDNA6nCROrb
4BGEX6Q8YFAaezioiYBBI6+sbmlEFzuxhkNB3Oiv3RsYMOwz8XITvIJZ6Y8sH4VX9sW0UGUmvtvv
A8BRuWpX8BPUpoPz0C/BWzLShXNm9UJehAUHyjc+gUjtm5ILEzmJkHpsj2f9nhfVZFvlqQ+hH0Q4
jefLjN6+uzCbHSdI7KMwcOVsHHg60fJJc/uC9JpqH1sxszWUG6VKKFQ11+5i/WbZ4J0sXx738bCh
sLG2lds6wGvVc1SerbbEjUByty7UuQzzvUeisB51Q3lmkMaEHzvozyuWgp4O43EK1WzAaUwMZqSL
y+7B/wbUzvqsd84sqgN3pLI5fwSNLQbNwuFfDc6vr7XBPpPNGhDGLGJOEn8dKFP7inXeNdZammY6
OKraL3VM2rwUTEuh4AY1cELouuUUjxOqilTEzv2AvK0USWZWZiaTYJHDCAX1IAeqQv9bjYXwFQO6
VkqAkiIj8p4SG706z+/VuIp22EAev1NZGAl0+9ip3rKZQzFFEU4piHNL60k1GM7Kex/cSOeq/MAe
qta1Y/dAAViOUcMDLfjmFUyM5wHWQI9nyVW3WjXchlemmaeoHqJfrUBANRLol9FMPbbICW4C1eAM
fw98n0amHnLlGpoGPeK/tbDaBQk8uoJqNTdCZBs8uiEBILgbvv58sIcnAGLKbvVPSmIDTvj2gHY5
MnfTBWFyvb8EitpfKaCdK+8BrvKMDBR5q0AoQR6Gg91t/51j2WM8/9hfPGeZS8EdFDgdBShVaUwh
tm7Py1i3sBA+MvPpkYP2fYQWcaY28JXukeDvCwcS+kSxyMB7is+Vzo8PocMh/BeHBIrdGZrQtRtm
g8kJjUG0J0d/+h7VeCLUhZQ/PIQ7k1CiNf4nUsL/5VIMe1s7MmeA2KxcxZNVWlIZ/DHqL/scNJwE
Eix2+HKKNaRgsqbRlglpUB9PAoBke37z5QYvgBhnWucXnbev9tvRgUqLsFI18NtqBko/5XBHxh3O
xck43rzdKPQOmeR7kjvizEB5hzPhH3fwStC8MuQPioux5uShlmUze4Q/ERBvuP5pmgT1hDwymXc5
vps2ykHymZ8gh68HsMCut4/VL6axOmyxfDyDB7zD4GvU0PL6GDpJ8sEioD5KyIBgzYVEemCyEmHb
iP0r9sM12WBCWQ6JESyr4NuZJ2OWYEhtxtbvfpRig5qaHvqifw0jri9ua4DC3h5e3khRypf5q3nK
9EXbTpktkmDHOksTWApC7kkrV/2yFUvQ2LfhK95s7/ekrFwvupfEwPFo0dlLHA43GLApdD0fguzb
C3wveqBrfd1a947YtJE0IT9tYSIqgQYGI3cC2hkWgHqKgzLLNfd50wPmA7U0BRngZS1mLFJe4Ole
koieccJygopTfjuzevyuZjKWS5J21keuJCx/5Qp8sU7HooC2cfoGM0jv2TOMaifHZFKyxjuKdnnN
lo0JA9Zwg21dEnUb7C9sVo3pzPofkSJVE5BPZF0RvtDH5UfjurkMjPyHmTLoJwbITCRB1ff9nzjd
kTfo7pQv28pPEdh61oy+qFxDZOhKXsqSh/YjQkW2sg+lHSsoS/IqQ4cI9tSbTHR7r7T0+x/csZWh
eSWl0+xf9PLYidDvqThmXgr8p3ljvAtMdBxtOy4Oj8K5LEyTLQFMT5Ng2dT3bNZq/4SlKA1TnnS8
svEBq1vswkxg+R0aG+/k7R1KfI6wAd1a7kM88u4LJEgXwfKrZFGzeUfMl40RLZXyE2ymrQwcogHw
ZHPn73j+4PdBtB2rUubdmAnZQztIhMxpQdpx2I2wIaRYZ2Tul3uKjMCV3IhCRfNDSUhyM0IuBZ1w
KsA9iFWkmlTnnr0se817OoSBet+8XqV6Nu93ntvTg96S0dMNeOWFHjPA+ejxdjpwCofmzIa1ypS8
Ld77yV58PCz/oYXqTrWrLG87pVHbhKlzbafGaVhsjbIjAohKYhXtypccNxvOTrZQGSpi+kHgJR2X
C61g0lnMn2m9A3D31TLyCKBxgmSkQk+9xGN9zQheuec5zZ0N9VMUUyzI8/RSaqkWt9/Fz7hid1aI
8NpZXLciA5Ggb2SVLeq4UUpbjzmEXA/i40Z2SV7rnD9RFFpx4qrJcNWo9+JpWhoVq0qUoTB/A5ch
eN7Phz/h5k7Ph3PFNN3rdIg6TM8HA6pRgS0yFvEYm8KDgsTY3/M3p1dsNk/WCkrjmRs3pw2AXADV
P2+GUMj8BntXT5z8pqE8KKyGLZuA8G9wXy6kuQODEJcbob64oLPU5nv0a0ffeT0XhEv7aSOjYlOt
Uavkmw2+APjPV6QX4Mt8c6GF9GwJ/clTSvgtrNnokB123+51wg79Qfuoc6VPm4mMx/kel9y9+urZ
1a774FmaZmAkbM/Pqw3rafjGcBHtDDbGKJ7BgNtxt5toXsNkimHmhj9Aq815vRjIhSxGzR3cvbSn
kPfr2rXg4wYhnFn50OogRViGbwCTI/haNwV2cRaJLmEBQYJTyu6MFNp6oAiAEcqLFlJe2sommkxj
Z/HpxtmxT0PfLuu4x/9Ue/Bo1GxNFUh0DjV/muLA2tMSdcm8Z9PynhVoA9YNQo5jm411fiFIFBl+
saSmTTtZhGUlCtj46Ncl54smjD6w4anxdMVEgFChjNZyPKvSZckkwlpyfNrO5k+ZOOxfRcNHzSSk
IznithVvYv6uhT6sy8VPYc0F9NtoC5dJAmy17R/9Ttbos51D75+0Ivq4AzIt//fE/hpXDQnC0+ik
S1L95eNUfR8r2dtDYR1VpNNc82e7Pj8K9a4T7SKQnpBif9Q/IuAyjqLdksANyM7ekNi9weBbh+L8
jvP+ZsQYlzRck9oCSchI5NqGYNxg0utaLLsUaCGRwYfYc/lfoaPG4dOtWn4MQoSlxpjtkiGDOHg8
nghr2c0dZ9RvE1C9YIfefkHSAaFpPzOZ1Vuu/1ID6MyaGqsBuJfneKQeDhkUjssQ8PZ9TODgl1qo
TVj4ZEPQ9CImpM9j3PfG53KEL+xFv7rWSSU6PpXtRWAttywtPRHTerovMM2JMMLWrFz2oWqkEq43
H8L8yPaWEaTxntB+CY2wFqBSOMeCOgAxjCcrRIUbc5RPRqHXT8ZXO5Us6bwcTk4jKQGi/k1qPVHT
orW/ML9VY9VaN6nXMLLWiHfn0fIMa3bmHpEOLTSfabYDiZv5Gni5R1trIZDv+lr2gg4c9BA7ySk7
48dowKMc8T8FvHGCjjCIJIorHVpmOboylxhWxJ+SVM7FRDkIeaIU/sXPgI1vdH6i8QYtAO+z6bvC
P4eHPaW9Yp0Xaftr8ZfFxu8KUxSfOl0VRh1H3iWq5vWwdLscMyeyH0C4TxJVQAYhsYvXw4b3YpvH
wJPCF6LUn3fxGrJNYP/v/9rNlcda+lJOjbDQn/OJ49thBE73xf/2Haz5lzbmzzzD/6uxJ+Yksx/2
ZWxQZuhWgRhoIDe6bM6WjhH7AVDD9/7M+Z6vzcPf/r3EvvSfymJ7NRg5Vlug2FjXnBpUktffUR4l
5r7t7Eb+QVO53za4nO+rTJytrWBoECiYQWo784MtHPUs+/67YZp3QB1tCx4LavGqlAKX2eAcoBwW
I8+QxttvMC/GbMw/bFmoYK/1Z5cQHmIoZSRAtxNRLAjiLnzKu3v/hwW553ZniJDUqcBcGtPL5Gon
xNZnAzQejQ5oiCYx+2TV019YCARxtp3BH6G1JYlhLTEPRu5LXIADFWRnqOYOTxxcAPw/zOnFedQN
j3OoYNRljmKJ+ISjxsp/yVUWS4yPgMVzJzIxwARcpI+lVtJzI04Ho1nkFr/LgmPbAPdM1JnGUddh
tfXIlkjDBuiRb1u7/nISc6uH/l8hpSBvskn1QebgYegROakz6RzLxTQkxNWrmneh5P4eATfLcw/p
YeBCuC+HQ9GBWpXSN8DUmJLvvr+j4ss8eaWz+fwn2haEUmpwvFAZkUstBrbcqwoyWUecgr0/JSlO
/SHAOiT1v75868thp0GK35ZVQuE7MjahItKnkO4LO91LydvE0TYp3dyJoV8LSW2QUAGdu0Cheu3m
Q4yONTC0P1ZSAfoWxHILGfzqDd4dhc7uU5Ypa5mEppc1LHDn5kKENs/x6mzxpr06bs4B1/JgjstN
DyEhUB8tK8fVokBzjfqIu2CdsB13b4cSONSoVWVHqckhtwmqbwAKXL15e95DsP7OnFF8rtRno9vB
B6ifctZuqtofzkH09KbbNik/VNgp9hSY4nvAedGMsjv+Zcrfq6ADEZSfdJo2+EV6sIruHZxPd9aF
zcBqc2326Mwllr1SdLH58+swAv+6c8LZBh2aTVrLqtiFM6KNm9V69JidZxXKuCQA2CdFFknq0RxK
nGblZh8UH/YRsB7kzmlVqX6a6apAwUoz0ONJranEFmmBG9jmDaBAfLbjyMrfyh4Pgjoul6nLUNOF
kNNMElOlu0Q0mND3S9VgGtoZPaMU8Hi8mK5fc26Ff36MQpJksE+V6Tz1Q9Vdq/gPPKYOnIdoXzEu
3im2SeC+p6AIVtNbDRHtAh95zVO0r1Sm+MnypHU60CKbD7xwJD8/HxcxS4kv0GOU7AxsP7ZMOy2A
rQmjGt1b0N2tPEDC/VOIrZUjuJR1ATtvHLUoeXeEIcqywHOT6OtLBIxSNNvCYdJHMVhcqkIuiOPl
aYlaZ+4/XRMWlRx8LjXASAmxpJs3aUHpjuRk7ix+8pTxJL9h6qmWrGd+11i7nVtp7ym0cx47QbHz
v5E18cSHDgPOekOA+XnvkDBXj0QUFFX7wET3MzbirNkwT6kvMZZ85mpVo/TLuhZG9GHn9/0qkDvQ
P7iXF6NL6exWskodhs/4+/0IjToUZe505a+6ApBRE1tzZ1RhNVj7ei0WzRQ/zMlr8iigDM2DvIAq
IWhWPs3nsEPlRLWbUmb3fONDcpFt8L84NZLD8xV+YepJtFZauxNLjfvePaKysLs6f04tGoXVBouB
c9ajyNqh7MY7s9N2IbuC7+Y1kM/gSJW9hUPJeZgEQRHwdPyAP3vaLqfQwmLkTLHFKQgL685Rr8Ij
NzlSiDdkta/awfnVu7Khkwd0J2+iHqujrwRl5+gEnj3w2lHi4NywOMZo8UTEwDIExfuhpB37Oaiz
He53cuAY5poIAqBbXFKyDJRuiE9ycOu2qZ0hQ8vivM6GUIl7Q3PwZY+AOXSDDgmhnGXTEhfabVz5
QMcBp5JgNCofrFghm+yZcenDa6DvdYaWEh2c2AtByd0sXTEKMn4lt5sJTUmWltNRbQ2sqydc1QYh
oxEaD2JBqcHXd1STZ9PiH+WKu/AeFTSw9Zq3Tg9deSiozX1FXFBk87piBGerBVktkpWDIWtkfrMm
u9FKYYN0i1WjazLc0FaPgG8mnM1YOhB9iIbIJj/43gSaIcqqfCFMfdIVBzXgC+L+qWjKaUcK/oK1
o0JQAaIdHoFZP5Iad685TO6Edycc3whL5eGJJLWCgqDhxkQ3F7c9Eghae+IXD4bGTX1z0NxdYMAC
ZFidFCMLQn4infjN4Bv9apP3OPs//K34ZiJmqQ0e9Vi/e6lrbQMUR1fakXIsH/oKfLTQh0kUJ2na
YAut7XhufXr0qR+Y4f7yGAO3lTnkNEdBijkzVcljzt29pqmD6jhJSCMQDRd8zd1UTydDfoR6d6sT
Ts3jzDEbuXGTl4evoi3q88FyQmPjyFU1drQ/K/e/740epmo2PlYGoKCIO3j7neaCFLAGnKB7XTxt
4Uv/WejjuPpHwGlhL0Z9CW/kxebU3jWASbCUtj7psf33oTX7OEYx1fYhDuAIr88NPiGuAEgzdkII
Nvh6R0l3wXMSIWiI8w8uO28yJyPKzJzFMkLzagH58EFPbIGcVfxzN7QHMoIPD8XporECIXP1siNL
amDKcUNd3tTDyknd7fDMgov7FdQ4Y4fxY/z4cgT8d/fGlCZu9P8bblnsJX9+CWXI7vVryqjG5b78
IooEr0LPMwuoOprV7730+acBatHYIPF+sG7Cz34ZtRLRC+V9f3GgOcFP0BSj9Gyer+sgbm+VpJB9
kZlfdFWYNUFIRxnRKk5bsw5S3XMplafnP2LZIWGGFDLJea5TusJIZ87UITFdSsBW6OPOY038QOKa
0rv1O+gzdlsGaheySr6keQCBTLFck1xBlDZP+nzrSOi81lfr44R7zcyr5QKTUEM9blj6bJAXe5r8
hzFt5XXBONz/cGfG1shP85ZDaoHkL5DQ/wDcVmsf74dqBlqJhTR7zODR7nuHbnznS1wol/r+1Lbg
ivoDUVkhg8l6u9RrThJEXef4Ujtw4Sy0tCDU9Czim12rO2ltSxTkXe3cxBM+9/JLqq1nxkj4Y3uT
I2Emh46ZbtUbcxvX4XcCtuDP0Hv64uJSp0ME/+7gz1C+WqmCKuclLovB2T+YwldKPmIm7B7cCTLe
FteNBlUcaipAy84sQu2EEy9ofOKPEYrhcEKQGJi4M4EdlRgc3n9CU54IMR69P25b1b6BDXuaev8f
mS0IcICh5PPMQwzmPHpaN4Yrw13v4/RqJn82OY6DTdI+mmMLcZP0yoFBoOlUPRNfC4egsSKncPrJ
pXoumHv1MWizpzNons0HgP7yXLzAVeZ0j72ilJxnP9Z7r7Jo7tBbm+GWAipKz55Yx2upawBT4tD9
MQtjnUUl4KvdIdijuuGouLvjXFNrO48MCYzfEiP9QTeODfK2TpmWGSfC2vtUxtTq9/yCvgjwiu7l
wtYLQsSQvuGDzW9mBnaq+UbiCr5Iu1HZnFTCQMghElElY7Uvv8FO6Uihyr5ajheYs9IQWKNiN3TS
KfsGZFla76m7ZsyK0sH69tPCg3aExKq4UyLQ7aPGUFZ+dp1ZFtXPWheOxu8jL/ZdCza1jKuO+ypC
HHfdtCE96F2R5dnIWFIHCtF/RY96GAxeKnI6o5bnFYXlK6ERUGHdsH5HbeVf1qd0QaIRxZpu4OA+
7srGQfVh/fFroGdg/2OktjAqMF8oIosRcEC6znVLkIagikFSYKumNTu2SVS1lBpZTaLao9wyH1HF
Dsvu7ope0tUqmK3CAKgjGxp7SpaMJYJj+W3aF3kR8yUz8dAH6cIjuGKK6c4RgZhKr6iHclM+u8jt
WslngV7wn5Yc3P1lyKixMCkxvWYkdGUbI2BltDEJrTHRv64bEG71DC0ptzd5xMFACOMzH3GRl/gY
D/wHedS4zCIaeo1BLlK2A0NQmYdDZlJ+h99kAWZIo8YciE8WusYNBZXyfuc6Ktb3GBQAaXcys7an
OVcYG8nL5TfPU/unXeyYWH9QQz+hmoInItzfr83RRB5KvTO5UrjcAxa4P3AFHZSmfFH/bKaXfqCc
3zITRFZwMmXenIXs+wqCU1UeG5KpBhamY/77TUcF59vGDPRgQB2kBCyVsB1VNr8Wbad/pehogSyZ
zoiIl2duMaVL37hMHaRCV3Gcn57t8PkNVsgytD5XdZmrZl7tsL6g1mbS+0SlZvjxpAUoNZqZU2Cw
3915Km2UBsxG0rnokIaXxAU1znAHJZ3CHMdeKkK7k6i/qYlqa+hPlNEZjyB7Z9qKrGfa4q1hWmry
Oa8h7SdGI2tGm27Nr2T1xDoS555e3B8G1ggn7MQ4NaaFd7gviG0Rv7whuQ/TEr9QX+k2EY3aQrx8
gGKD/Ywwh6YUkqgXg8cytrALUoRvnRbGDWq1NhrQnPzwAqb2dOgktMhQakH1HXQB/2pPeS0OUXvM
LioiwHMRuvRiHpRplaT+Uv5WzHGdBiNWCN65L7t4TXL05CWXEH+z92lYCs7CRfiWSiFUoDOxUpBt
y6xJZGx+JufnFCfL7DtkFB9RM5m0+jiNfoe2dczfL0bhe+NUp/lX65OCfadjKxSxlF2onOs0tp4K
lG3tny568V22CD6euWkAZgQazQ9O0bMhSdXvLmZo8bsY7s+UtiRq8eOfmNBNs1HhbOu/9DJjNYnm
Hxt88UhVssgQNaCpalGs0/ni+Ouz3P1j2r4wSC0FQ/uAlI2BCcTcJTklEHZOt1z8WFCFQJsaMC0M
vl/n/UnOPg4FyFRat/r4FpglDirZSXezlKi6VVN36cV+Z0Jm5w4N89pfkXwrovQv+JBjmfBx+OfG
dlqdeyxLjVJAuAlzZmrDcFarPt9EgA0NcS6Hv0Usgh0QYmIjNm/p+F4borRcwF4XnfIgV5oen80/
jrbfmKdNiScuYCdCuAegAILvpaVlAIRuCUszY9mhHSVJU+/mr7AZR9bsTzAzRk50DxWFySway/0d
jnWonJn7OfEDHqXV45EdCh2jqHAzFB23/BjkDOkclNNGs4Iu1d8g9y6mtj3G0tURcHxLFpqVX8tu
uZ3MHZyY29qhvywWFi0Nq7L9IJpY2fUj+lb3owY4pIdgwxJ6P8gUdNwqzSt0yR6NGAsaLV2wW8ul
JRjQoGJuVlJr2tRshLm0nlf/glttweMPhYuvfYbT10Hl7jqEbB9+Tog0qQiiHlZYVHfzbGGrHUiK
It4eFqfcsT6mXYzcbeIrTAhqX1//aW+ZzybdRgcOFch+apCGEd/+tIjCl3YqQF9TiMsyCIMLhKJ/
1/CI26p/vHbQTpcfqe36S7NHKeod/4McsoHojPoIm79XhLSOssjhgN2oECJgUF2Lzqa8GLqzmg//
rpBJOUjZ60cAvDONcbgZB0LzLxOaFT+LjfGRYoajzVXxvZmcWrzoaZdfnQu2AU2iO0+tCaerycn+
6ocG76UCsDjYGHmBrYTWWGqjwreDPJ2A8RnirICgQag+QHXkvERVm8Nyf6IyDurpkrh535r9aNl3
rsGLrObkgDsL0D4mqiDgHummvcfJxgWs4cP6wXtEGMstnJ7pKw4DW4FA6V+kjvqRLo2yyx60bls1
LNBlA1NkoeduvLC7qfNmax6NDdOgG3aW2NUkHz48xxU+0toA/u+rcKLn/q1+7prOQLB8X/jofFsu
shfgEJTiRx/GIHviOIJYXyGIKTOGh+psLhJpgCXVMR38548qvXRqI3YGnR1Y1AfjF+L8gy+U2Yox
9fa7v4ZS57/ySw/mAOwYv0qcItfbvAK9cG7e3LSn09Jphlci4IswbqsuruleBiR+Hj4niWWkvveQ
97GqvEUA+5t1Pp4c1ran/he7IH332JF2cdtn1mSidkprD1Y9AAufYR2hnNIXNO+J5y37Hf3Gh6PX
VoK70Oj7S10E460Pc8H0n8dr99zoYKIOCIbqI3SR9VEAfjjNi6OWTKBdyXX5Ut6uzlU7CUiIVGAe
Cbi87gqPScnRTWPJspbO+TZ3ny5LHjALPmJ67D/Xva5ZjlLT0HwO8W1n2MnKSJYgUQYVbBeGLiW2
ZimGYPb9tUklK9Lrgf+12R9x3Ah/cyggFC8ZYpB3fiRdF+YMgRuqibRhJxRHRv8Ns13PdYM9vAde
51zYD3EtZa6v0h5RLUSlhZ63MxmJ/TfaUB9AbBCvZA3BQw2chwfY0QrLc9zM43+r8YCHzaqM/3fr
UPVIlmeZqlmwpgfimI2EAg291MbHe6rgQVj4YJ/OkAakCcAkwyYR5NQbVFPefAd9QGlQxwTWatjX
rgEHYH971oNjMDbQnfbCJo2XMefzTkmGZGYPqR7uHOVA6RNm8b7k9MsDOCadihoJwJxoMHclJ0Q4
8leZvRL3LQdSp6utH664Cp6j2IVy9i62DziYVL05B/bCpAZbSzsSpuN6Qyp5lQECkE6RSYNGr0hU
x8AwW4mSkWOihx5QfdpqpSUj/DRLKr3kWflJpvZHxgCfsdeexEuKuJ19RNqWYf0K6LkNJzRJtU7D
ayz5K6EPoe4Wh02gfSpaIA3y7220z3Yf8IFvuaCcWKxD2u7w5VVm6CBcgd0Ze1h6ihIRVJl+Eh07
mYw64y9SynWXUCC2OKn2ym8qtCeIj+k0zr/vPsFPGJyx7LRAcvqKaxGuzBAC7HURw4VmRvlQh2vU
G/czSS2A1QtY5JmOXd/RQaQzVFVlq0Mr/biNTITTWLdngX61hqPUKgHt8uR8Cy+ZZBCvBHkzsJkR
gEgJgpFsCnpEz/RaXi5pSQ04rwnkCgHcGOJ3bhM7Tbd8W34FXfR0LGSLEG6fvQCeXbnD0FFu0OCw
fOnIwW2dOeW50YAKQx/30tvpUS39VIrkwKXgjwK8onSy9+8NmFZaC7x444WAkZI3z/U+ZKBjvzOk
ss61RR+iGCphU44MdruB+E0SBIMlH13pSjcqW9u7+A1D5fuC/8Bml7LQ86/n9leetcw87cHMucOi
twjWBScA89aZB+exruEiAwjhS6BwLXxreiHdpEofIIhfPoaOUE50xxz9RI38mskxvb4D3PE2Zjtp
VvuB9wfOK7tILjJ/pAjBYxLkBVOLJgug/SoWGi3RYK2zNJA3j2+aUTQYNvE6QPq5rGyBF9r3YzD6
m02TVGBlIK5wINlfjbaQAdjljHQKVLQnn1qJLJz/2Pvl1N/9uZxUvhcL6xY5giz1SnsKtEWhfOrl
pfJfbYS+lM73fbbaEtkLnS3od+bOq/HeAhaeVwmsTCvkkyxtohW1ZoVUopEywgmaUpL16rNUChXu
NgMGowJ9Yvke12EdPlXuVIi+Tr2/5q3QeQpgmNwOUrFHLLKtnxDZiY/iVsJblyd6N5lS/hTioYGy
S3dYXujiBPS6O2FCOKJ/qxGlrke3rrGd+iUIEW6UR2/oggabHnY3wTkYSTsqOskO/re+8j2FAkOK
xv3IeRlPaYIBA9+WtB0J6sFXaljg8MdDoj6svkS82ueVevTAeUwiCV6Stf1r1OpBCXu6jzwCjrxi
wwyRoRfhyzZKgQFFNT7gLW+pRgAHSfkwqfb5y57jzQHAn38wi4Sh1UW+uSnvE+PnOPy6tBO2Fvkg
toPu+l7AatCmyVGcsTIQId7FB5Ep4/Uqsp7HxsLaVRrja+FfmN29tl5RG6OGZ3V6+K3OluoNevTv
z2E1K1XHqxXHUyo345zKJCZvMZaGHHPyDxIubuc2eRMzPYQ6kyGCOWvhFB5dF881S2wY8zMuGZT6
YTfwpeKHRxQOWwPtR/tl1TQlfrVUJuoq83SPUWVVCqYg5F3akZnOQMesu+5v+au5jX6NQkxxig2z
OfAqwNl1I144g5VnzqiBKVsa8RGYMXHY0ksPYsOaPpGm9zbv8kYJ7KR8v4TTssbKvSUWfJsXXjS6
lU1MyMy9Xk/YSF1YuMiTvzXK8QqvZDdFXryY3uh49/zonuv411ljk6lw7t9qgw53B8f0OQStg+Vv
kYQY9JGuRtPQx4LdHv5tJu3WEzzn0voa0+OlfBhfR0CG5hSFst9twLvk4AS06TqV6RZMNsesrRGE
HyaordtckySv7h5a8rMGaFT+JNa/x5kFyDMYrXKcBBU4IAch3XA73vpqn8enEdLGc5AJY1IlSMf4
rNNw0/D5tV3RR8BUw5x1e+k3c1f18fx55w0YmYhuYys5E88B4acCD7oQfT9c/mCRqPex9UKIignO
9oAIZF3zJWCWwwRB0GA23xJ+b9xw7y0+99UgRaVIPZ9Ynu1/86f6Qwc8myjyPawHlONw3sJCFRu/
/Y2bwsCwc7QNdh1HeRcifIIZsUbC2oK4mfsLSmzXs7k3jfQFOzehxyVaaN6r3mGwBp6HtnKcdDEZ
vvpz0SxaGZMdjQqtScyor7EY1rHcRZeTmNj/QYPn+Ejl6uKcbp45+ir/a7dKqXlNhAYr8B5ewVoN
1l7YQKXnH75vLqvUUqlNlHcpvnXvX2HSVYly+HzdBacFhz47Jl9nvLmLbLbDQc0dewR1bIZDxjVh
sh1YTs4qqiS1Ox/Vm3SlmhqZXqWDt1W5eIGOh2lbyGmmbjhke+R8BvQSuPKxF0YHMAgrQqgKSxBY
OjgJSAsCrvziAAPWP2noKdJYwc8u6vem9IyDqzJdM85IM4zEder+KkZKnFNh0blxpZuJ2ilQM//N
EmmXKEStpIwdA7TkFG2HvT9ZGI9lnLdZhsLmp4L07aaagGCtU1OB5JAMszQGHcjTqTt+YbodBar1
tMWI3JB4zsQtUs2E2QCyA51683G2/a0N8NuTtaEEgSEC0E2+/vcw7RgjtSd3xGpZQnnVvavUs91P
NH5A+MD+8ComMMwHgE/IfibJZVLRsFI1eHqHPv7jnvuiuiatHZUWNNUhr4w9iyakiEFPyXxlh6Y3
YZIkOGw8HgzC7HNdtjEdWwfWslPanLc6bIuqcuNIK3DNn5DI0hfnKa+XZKC7GIJXs6WkfYPE58qJ
nG/OWw3ndv/ocIe+tFBL0/XGR6gPCqs7ZxjuDpw2Zpp0jtxT6h1PgNoo3VkvlTN4uqAZ3R/M+Xdl
fZiNQ8Z+1IhDsA7aJFEsup/yig1kllfQHj4AOMOq/1XagjR0hTjqmfeSgbu137nvrppaZGNRdFuH
hokaClwYeDEHN+BXj1VAxFKfGcaP1vE5SbU5KM1kTgVB2VbUfHzbZqTcKukAl+4SckbSjbvhXNi1
wh2+CbS5peBW3J8gbvW0BHkUm2OwjottPi2UFvFD/Gp8tqSkgTHErgOEjIT9VLQNvybfCmAzz+Fl
Wj/MPLuqqQAhX/dkNQ40CZYlkn3Meu+5DegCx7XsHakY1KIdl0OfjLessXXZS3jo5yNME+Jei092
gGMVUOr3mGCvdnhkV5UeQRGDhOOs3+rAkpFy1c7cOGOQ4I27YlQ1HOIcHdp9wcLWLAVbaOItFqhP
Dwtoye6SpLrO3kusH61n6p82QaI/LsoHsBeTKBmG0hbb+le1PSzIWlAUjdAoSPYLqnWZJociyYcS
Ic6A15QigiQ7izGdrGb+nImIHnIRNx5gXtH6FbinQBFt09YXQ5afU772oAf9kW3/v2oFNx2lpJA4
LsPnGGaga+F0S4FG0IFyX5UkunzqwnDAgDm9wri0QxDRydnjJFexhvpV6iCoafpKbRWTgrRUDJi4
SakgoIBWBmcl8nPG01OvQIm4DOym40hoDPUN+WyKF+NKBLpT6tZWW82MuW7teilZHboAWPCpb+TP
VjXTluavHcccC+UWdRaZ+6QD5WXgURH+4WACGoKV4j+cQBkwC1u3Ogv2iuN568LwcAN7AXz6FSUG
iVR6IvDlfgQOLQ4qK0YoU4hCNsCHKOu9l59NMchq2+vkaOPVfg2wFBt3s+jcj5YAFVPH29tqP/9V
I2Pdkt0hl3B18f9ghvUqXejt+jac2j7KwY7tnPzqlPYyCGFFddwlD364QJEv8QCs7TdPreKzkAxq
0Vu3vV/JCrHswnRKsobbHHSHuGeu/KPgO8O6bc80LbjgtjSjwJfPk+TXZIPd+l0eNINOi249hvhH
Xomm2mDBKof97rcyR3Cx3EPpSJrukDXpmAnfcdHzy7CnZDnbXHVYyvEi0jfBoZDEhnsco4ymYPnP
SfChscFKKIYrW59gHJwNnE0+K1JCRfMGfOOutDtPoMk0lv5tbSE5t/fMj3zBdYdNceyctjlvXOPf
yv4TbjksSpQC0rhIhy2hwrC10iT8mQ/VJ+GMZe2VyJFxBw28d/gTnYPfUSvqstYpQVY4XXyEgn/S
6/3H7YrEGLfwc/EYXQAyHU53QUT3YBMZMnE6O5HAjy4VAODUs+F22hBPsUsOIPbox3dBCuZt/xrv
nTzP/JesngX31YqecfRYY967QL3lOyYZosZoPJwZ1xpB6fAcUKj76Id02i3n/OzdqHTDBUflrdF6
gf3twWPSayViFrv8hZfqDU2ZRAcr59oV+WuUVsjpQsms4KSXXV83h/cN71ysXpHdjeh6Of6IN9bW
QDP+uBs4zL2xVzUK2wtr6QxhEWNqgHm0zcrv8L+BpZjlOX87jCg5DgbFrkIX5o2U5GAQ6w4IyZpE
OahTcUNS6L2sogsEL82VVy0F4M2lNo1Ze1ODayVMBmDE1Ohn4Wfj474Y4UeRUqtwbuL0/uhfxpeT
8DWiOqVAyal5Cp1wNnQblXxUER5CztL+CWkXcxD8Mfj6MWG+k7hhM3o2xjq4Uh3Q6w3M619KGd5L
Ih8OAysm/UtG/6MdlOULYptNRIJISDGRWszbj0+Lvr3R96mKTBUoo+J3Rwao13J7tTQONu+ZF/HK
vFs1Oqj9kSgjXQb0R+ydO+jqhhTo931Zc+1qioCJugfBID0ijpMDswN1NfTH68c2gAQFc4fpGbPJ
o+CRQZ8dNvctcTLxYMHrX2vHTJZTpav54bnHPVcH1o1E/4/WGtKH2/0EzSkPe8l/xGoeGy4g8CZQ
md1ub3Wpa5bZECA+is8LJ2bxTUqRw2G2J0zs0WorsXSVfn9c7fKjz9PWhlqEkMdOmTCZoTtnQT93
/MC3/QZPzGAfioNnBzBk2ZXJsXC5x4X8sZNOOClXAZKIM5FTJjqiVhetk6XniMyO3YjVE1pmcfhq
XR7zgyalSy6GWcBjO6DLzZRr9oZGcv9K8A2hxny+TbK7JZsA04GTUua+Gb+lasUyoSifiDycO5/+
JO7FWQQsfeBDvVG+Y/wBuuaWQ7Fg4Wt44iqpDIzBK8d2t1DHWt3qjKytiPqSRg7D/PpS8bnDTr5a
uV79ZrhiiferlWZAJqjkshiLwvAg56dRuc0dVtCE2zn6l0oKDn+v/4UB33QN6EOO5rEFKzsEfFdL
8XMfqVK8Ne+ZgJoQ8IQAOf1JzmHJe6FlFVztG0QENhImbKP1axg2x+j20HeCqr7HSz2LiFmzmQHX
Pf0LkT7hlh878wtumkEiGKRXqBNWWzOLb9YnXqi+EvS//hICpBx2GxTU+KsWE+MOBAll4tRv5SHO
UZPGcn0y8sCuxHv46KbQ3UoxHtSysLMCHxCE3NcbVEMoTDETtI2ekcERbKt4H3ejWfMRflZhKqkU
d3RoEkQsgyo5dv4okV80mxh6BOjJBt5/AInAGBr59FQxHvy8w1z7l4gCxIbIwA8aWFyFmc039PFb
ptIvZOKVSvIxpeOhWgCYge2IUDHAwqjZP9kPwWOt40D4HN9AzwsRdKsjpSR3LBF1Zir0czYzI8S/
4kKianVFMC/i3dmc2qAboS3WHvaRD0Hwa0RhSdJ4+c4xvuCh1zIZ3Z1ISqKq5unGnLbK8x2OhHQ2
ohENN3ufcR4hcQSbDwK4EdwwfEu9iai4KrxW59lMRF8RSwXILx4XfTx4gl5XOBzgFL/b+zMkN4Hb
YnpUObZ4ujeLgUBT8UDdH21oLpVJ0ZnIVdkS0XvuD/+ABGoeKOJdIFS3QxsWsJfSInTSm4+M8yeq
iVXh36CX96p6ezzKAm9ALUWqR8Ww7FnEgzZF98vSVcj1eifjUZ9VNk+e8mk0SaZkghARTMNSb9jY
UwvUfYa0aaCn7Ciu73tXhVtukKxnPcP4CwcQhBmslDVbxwLduHs2bKAq3kuM2rrtr3CJon4Uwtv7
0R5y47NNZfFUDJtBOkcZBqOgrBSb0ie1debw5WQRFFzXIHm6yDqKPzMmuZybhrK088OVNF2rtbBf
7ExKMBAwLkEId7E2Msz4mRqEMlTpuGggXNtAfO5P7YfDd7LDCt2FAmqy3XjXJPf+o5uz9rWvntUD
L/BrC8/aG4tGuACXabS+9/4ZIX2pcFZt99m4KOuMbPw8sWhPAs8npXxwNxU2pm8MReX54BMoGfYk
4ivFON7xkqEZayo/GHnSYSi5czyuu66tmICmtIL0jf/xbHrhRXvP9+kml2A+ox/z5G03icjNG2Va
6zvKg7iooX80w0CdxthTQ4cvmjtygxBwFtPJicxQymVNLfAm6S/jeE80dSacRyT/9s/1t1ifpktl
L3QwKYB5Zu4WgxwivvpAxIklELTWdCyoPGe/3ySsdbfA29RmL2YV1+FyQk6oZKbXuT4Gz/m6UWJx
4DCbpEtplG6xBeiu8xiT260NJjz2Xorqg5K77ewzooxIvBOjF40p+Y4LhZChAKdyf09GM14ZPqZz
5Bac/QmVOzj/Ze+FKQSJ7KCvsYKEetbwUFsYUzfTUORgEtUy66JHYOBVFoXtO3o29TLzIsbGsXUc
YB+x/E2O+4O5NjOFP6QwVL2DQRQYfrczGtuulF46GEmiWHyoNQ1RR5+k00oy0IZWNsqwruqaJO9f
hCdjJeAEwZZu5V1QD5KVIt17rF3qrd9Sdns/jhMjElHRaGlqYgKIeGrD0pzENQHZLDCeMZNKDgZP
6aRE14h6qKOSwmWA82V9noV0ND4Eh0QLo0ivCEEJKNLZIkePbIEffktZOaO5OQ2zcVj9EAuOd/5u
uCsmnkV2ZSSTj5TT1yDYQwiLEd6uCWs86xyU72KY1O98IDPl45se/HAErC9xrpBkAHo5Xr7HheX0
YcOVcTFpbyQ/yyt0x5j7p6ideNhlbMmL5wbshZqnEpWTy6NmLJkDG5jn1No+3EXvvIKYu+pZmzy3
la7cZWS7aujuntHD6WzGe0jrMgWVsZekpCTx4sF7gecy82Ekkd/VXZv56GTrj2UfdXPvCUhCbNEO
cODd1GzsreILC0n8VfuKvfJ8xcFYUS9ff8WdQCA3ao945V75skaqJAMUCX5SMWnfuGQoh6rup8Av
BhJmTudntxqeJ4DKMtsza2aNQ97/RI7vpK/7jGOcfJ4atbbJXJoumXk3rxeRc78n6avYU1KeD4s+
rEExJxptoEAlWNrC+ig17v3zmi5n4EQIJXD7hyCN/d0BDp3XE1TgsN8io0Io7Bb85ITPl5wXibfp
gES5akaGypuVx0Uu08m5FeK7rNJqfCNQmg7vdHZR9OxuZWjd/tM/6fADzYwAArAq7bas3PdMXWpy
fQ0njwve/mC73mGgnWhesEgkOZR1R6yjUeLGHju3Ls4CE6yPiCWhBOBpqrANK7g7n7PXDRdLsF+v
3yoKLBB0z6vF8NX2pbO6zef2eT1ik/7/tp7Bkpxn5KxKAXSMNZ6YI5TpVmTj0WTrlAbnbLTlu5T0
OMpN81TU45KUaqQSXZkKwyS7xDApl7XJar3ByTG2QRyTG4CR7sWX3VauZ8er6NntLLIrsUa1v2a3
wDEEv4eMKqTsD/r/70jS/OAYkxCYCo9NjfaSag2Lq4XcVrP46Up8zVZ+kecj2d24f9T4ZfjQWO3P
PrUAM1L7LKsbpx6Qu5cwyMDRCgw59a51m4J1S7BWVNdBC5bBMVr1NRqTr33BZFruD7+YtVmNl0QN
1S7uXvNuvdmNUQeivFUuTmysngqTn2Vz4B3b+RwNFn3tNF/9eY68fbYvvAk467uhEpHEDnRwVS1V
XxojJAGIgCajAl6T1QudDLyA8i/9qcdlwiJdLwWmstfS87tUAuJBCzxVepilFpktPpJNSFo+DV8I
WN6vd05rte4JzUNG7xgYd/xXOr4FI5MIFcwbDWs2F8h6KOQ8EGcDyI+Tfo6dCMQtugARXY9I+tsQ
EEvPjACbkuff4vfEJLpFrY+H5qTN7RiFQdC53Acj2I5wXGsXYm5Nd3dl5ct5yAnF7XIOAoeP788a
5FCjyMUh5Jd4/iZZkGHeuoFkzgZB7eH23BNaqiVsA3qAZ6mfzWGTrDVlyFIcVrBK6R/x8jwt6z86
oZeoy4YPMWx23Blbtykt5aniSrLpOKxLkNZLYO8yiohpRhbiwDE+wSTOim7a6gCpShCGWyVMwVLN
UbtX73R5Ym/NjJ4tJbglv2wiMZyEB4yb84380QnlfDT16hiW3/eN3brWt3aa6IQmDOMa9ifMcFGU
zU8K034wze9FLv2rNZKl2RlsyOSSR/cCfCWhP/IfQ4S/OcC7eBWcuVhQC8vxJ+TQfSPg/q3XcNRD
j0r5uvnTB+79aRn3BsQX1NazifwbzZPDNo6z+vwA5sktsyzYfaCouXYN5CNNzW1mrbmu2aKv8gf+
ivPAOO01HERwru8iiNTzzYBZeNeqeqmtkeAKxy6lu5IGyrdq3SruWSzOQnEzZKzDpHlG5nO8+409
q1unRWKHLgz6M78B6i7bfxqdwMMqwMKiOMo4NpciMR63gMb1ZR5aM/8s1dgaZR5bGPy64iRvE7GI
HaEHJPoLHc7LWxKKn+Cl1d2SQO3/Ma/7KhAFy1sKqZVnBZ34kMl9CMoA2Phw/mC/3XehLQ+0wHLI
85PIEJGuqDavQbkrUZ8FSzUvCfQ3zabmMzjN7ZUImG9ZlDncjTYwNiElmwH5NLshVP6HIzjSaUQj
YNlWfUfPsucvOb+foh3Sbhmo7qSWKcT/eTMunbaf5BvN0l464Wd72L3Pcvp5PUDGziIKWmDcXVb3
kbOPsRcP6ipr9cBLRd4vQm0qwplDhhFY8YRQuvrxzfXWrYkY2FC9UccswyjGJKNvYmRu5naYrbOn
1882DjKdC2jQIYAk1VAcVs1O6sOg6HBScYNFcfkDuE8IXHfgzY7byLapwyhmi14jO9zKiHmtiaU6
CnxtQ8Q7yQVUo/D3Gzzw+ztbHrREXGiLocXLZVLVQ0m9ZdP/b2IdoANIU12vrMzlHyT5u/jc/hd/
crRaDtzV5Y/o79tz9ZHfocNRMUPZIM16ZMzgFInpTaAj2CEX9uufxS6kkCAYUyn1CaUlALoCjP5y
gf10LqKIoA0YBcT+N/LhBe57iYk0NnhIni+fXjGO+nkFpfyOKpBCMAyPe9LM2gZXUZDliOT1WdFp
T1W5rLrh7440Ta2VCDj/60KIl1bfBPcPgcuu3ySASIWevKFwvi4EctKaWVQyOcF3fzYtp0/WUSXU
NANrnjonNxkzUCiVIyRdmN/LD3Q1M0cA4pdVm+bcnN5dycHq01tT0UfBn8QqimAi1gMKmkN/VMYr
A8bNNZ+gdXZckEEtnQGfJFZH58UVhm3/AdHmm2mtfcdKPVJacPwG72nD5TelC4teyq0NZiH2+Vem
iOJUB3gaZabdMJG+8ElXoOzQ9N8TD3VBrJtSDblmuzSNhiFYmWIe4rH2tmmOk3B9V0GuNxPMDTat
VZTBAM4rtuH0/IqqCWzhJE+BVzpNjQMoxU/h1zBskjSqGY2Huhaxde1baNHi/xDEOEreBGhTxWN9
u/TZl9OkxXFxt9acJ6IS60n5tMpGt8nN15aBLYOPE3x+cMh2rMyLnkZeeJw0uiXXK1De+RmRK/Ff
Wb4d6Lv1qQ/DERJigHn0prU00Zr5vPjuEaAe4NkzdNxe5XD9+o9QtA23z7Wbswua0sSVQMGSBRKB
RPra+K+fladCFpMYay3KIJTnu9VCQj0vmXWbMbMhvbpAgcdjmE0UecrqFImmAkPqGcsWnIA/TjyX
2fjFYuHy0aeJ/VyU/rJw55CuKAumhHCbx3nkWwqZHsBPeOK2KlxYPUbJFxqX0dmTtUYghVnO8i2j
Baxs7gYnZ8A/1YAnLeErpQwVUfq7aGFqZAbkzxuUMNA+mJvyK3oyZOMsM8RUDlrz+qUXiBIVPHau
C5KINFTHAzu3aYpEw/Tio/T2NaXdLn7OziufBfX2JPKaOhydd3NspsmeM8tWCVehFj6lE3oW3zMv
Q09Kwb8wE8bf/KKNhzRKxYvej3e9fBkFvEJNkjpTjJk4t/oAqV9ZnTeS9ALwjk+LRhZwgNqWA+sa
6DuxkBm5E57glJvR1H1avvxBlJaULLVgk7qnu944n7Lr5rG9M0HQBgXJaZW441N8FH0qpK1eBTNe
euAlPv2Y9xiDKFJu0qKD/P1QEoaZ7oqMjRU9g4aGrGn9X4F77lzyhQNbiXcV+zxPm/Zl+RKB2bPl
EijPKemiSlRKI0GLwg99ACBTM4mD00fAHyfJ12FuVPdD10Sk344Uv6H1RleYW7EfNhE00qeAi880
9B8DMLHhbAV07NQNnfBF65z6JggwO9L7n7yPcLq+whO/pAsN+VR8hNKLRiQH0yJe+Xf5mEgMeOPp
AgEDlQqgleW/Bqn5qpPRs5xyeBGE6tKZf3vKvv9Y9608KaMj4QmNBgtS2AiZGGd5IzVOYPsjLQqs
w3vBP23CobQa4VgfmwLnaHByjEgzE/yySkeIX5lVSMJdT5QUV/tI6LpeieOrZMSNFxtmyZY1O6LK
zgFUSziwx+caVk93lcx59ld7Rrhb5sc0BjD5zfs8CNhDdOUNNid6nV8VrdLSjC1yuW2udOkJ4U8i
bgVVKIimMeSCpgWI1pEDLvdpDUpe7xpWAIdeAB/3HwtCi5ASOb5VWr1BQBEpoLriy/UgGydGrGow
4FjFWhTk9FoDxOV5v9NbRUnCNN0ejXDnA/BA2XsVwpqiQyM7wfeZzFE5wLsZA6o4O/2Laa8Pqtci
tRTcA729Ob1FAPFjAnas5EtfIy4JuZHH4togmmZn1i1WDUOnsIIz8LHlFd2cALZyQwSe1aLhAKwm
fBDmFAWDFPvg7DUuO9o9tCkj9uwOYSaV6eKEaw3a/rs7c3bXQ13wqlYeFBcON28+q00H+IPKWIAB
4Y/prf+sPMwYfPIaMlhfXscdhzpTGquU8KkU5vdncC9XoJTiscv42A6Beu2Af7FQ/9/K6Ly9Kxvx
Icj8nAKfOt2PpsrvBLU+sL3k01jVYe24Jp/aYvoVD5gA2+mC2BTh0pfcd+ZKKmjCTqiLZ6vEJPiZ
gGlDtGPnzegwIZF0IY25JXBR9sr5hYbWXqbMe+FeMssSlz5q+ERMA4JLG4TKObMWQ+BSm3yjmwyu
5okJY9T0SmbC+0q2tFhUXkRhIJF12BZUJ+FjfkZ2gbzQpdqy+4r2wLRWbtdxe2CHlOGRWUn1XVwh
ImUxKPMJ+kZW22WN7rI1lF4tN44Rk4YwEQw65Cd440JC3gt85Zffrje5XkHsSLFsbBdQZbFDMi5Q
rGMLIDwLPg+GtxOZRSJb5wF5Xe9FMkw/o0AIvv169aDsndzAzEJtU2A26Iv65/Mqf7zuhBu7O59I
Yo8bbKzjePrEu3XwOFW77guI1M79nMXaHztj0ZOrGt0XUGqssj1r+kOwoOih9GlynjoU9HAxaHoa
3U7CEIqWQKouoI/IDi1/Ulg1/9JGCg3qZhME8hGDzn/qIRfvfw6mZjHtXqu/xA8b8bb7AUNYNSpl
pYoZuMOo8nczFMIEv3B8rSd3OpkU6ucxO7OYkLhugLxUbJQwpj5pQgNxLDkLAui6o69k0497MVQm
mfJTh6ZKn1VoVUDwVa2qSVCXMdoGGrPQk4FzkKuX1zLJiVSgbGzdzBTixkrXWoep5F9GxR2SV2Mt
p6LGTjulh26c2AK9JYasusmCuSoqAGKi2EGhcydKQkJinR6T8IBn+oNACDv22LAZ90W9A/UVlRUD
8Q4da3FkqkpBno31x8E7gQCNlz6vfEK9LCo9Kkzkqo06OjUiCIvxcxpkzogVNQhmp5pjjRLd/I7G
FiFdSKO9kh7J2jaZM3ORkUPD8qnKAuejrc2PorlNSuBGxodOkxyp1gSogr+wpL88W2AJ+lqFU8Ol
u3uAfLYVEY9fQuNEEYOBcBszDfuD8zecst4zQOkwdBOsuS6CH9YoMHnMYsccCMvFi2LP2Mfif4Uh
ngwVzOh85vG33SBp2dc/uSC8283pJT1clraFfp+/Hbyq8SGYo15DgA6rHB7g5TttX6i8reWKIVzY
aE7hIYe7EoasP3+ajO/QSV+818Og7GigC/49oN1nnDPzyFH+FeyeXXf3k2rPnDakEI9jFaK5txra
gSONAXtpPS06tP/M9n9K8M5Z5v1eY+hgvsV7pUBDRKG4tuXNrxw5m7SJRGEs6s5dAOExbw8Zp3Lk
z79IubQENx85MnEy8YUgj7+perpvY1a3K2zm/CGh1+n38mcLFmeVQSDGcJ2IMhcBoFjKH54j1/3h
WMN5qkWOsNucVI++ywbfFJoLcff324CKLJ4IiQXL7PCwb6Kq20kj52uZnauYlggZPs6UAlmN4lpq
g78cI+fm+nqDEw2dIp4zjTJ25GguO2h1iiR2g2B5kEBRiCEs59ZsUH5x5UtYpPw+YkRXAUy5s27H
Ja6Bn48cE1ykp/gdiMTVC5NUPLr7clPDdlol52zQsvjeGAhZgpytz4HOFTNBlruGAL6o0VSSZ+8q
Kezk17UMSL5oFwESa6gOEmiaXLMX39BMfLs6h75nm9/9SnNvWA/5baFLGSr6W7xB3/CYPv/zDMlS
CRR0RP67jDZFtwHozEnHSqrxyNW2Aw3jEZE53SIY7lMjPEjeg+zuT6L/PVqKrRdVCi90ckUoc77l
TdQumbTjqAF2DNk+tt4k/RHFxF7d0WbMyTwiqHrTjk/SwsQnDSPKH2fUNWS+0a52M2Cq1l3QBsXM
FaEh2vsRzni52opv1gh09YkuVgLOOBIzkOCV2wQIX6KLbIpLRqNdXarIedrqKAfmP+9Nhwut5vRo
Aerbht/NPtcLYEVyGQIEqa/LnvWxflvyYmkBKu1wl6nGKxpUtO1FiMT4cwoD1znAyjHFhbYRA1CP
Zd77qdVm992h6dYOdLQp9FXQ87WvYT6L4x5ZWoYwZQ1Jg0ZX3HVXD23iDGTGwL9zKmV64smMMiYo
DyVDOSB4fBUyhUS34qi8wRTYe8oo1PKV18a/2c36Ka7VCvrigx1e2zbIOlelzpHAOKALUqSyVlR6
DaTeWrFpYUXU8IcMGSfp8tXTmT3Qp969SnZzN3cteLib1WrRGWAN7lIDobpTKfzCZXHP1g+z4wvp
4TdAT4RHgENCEWk4j8Hnzsrb1Aiofctobmi1lh0wsnqsuHxhfPiyG6fWf5NZ19rIU+zahEScWqNz
tjwCsVKnKnzSlwJ6x6t+0AQjr+RBGVGba6Pksu8BptHaM/8Abs4gq1eEsR50Hx4FrCW6Ud6jYm8n
fDv9VoKFfCbUpDMR/Nt+ziGkAFREJpMAMjMp0/+kQUl07t48sQg5PxMygHUS9Q0I+XHCXm3uGGRV
BtHYp+okZucGFV+eRASOyzzgWQ56nyTJ+rfzQuCLvf0pVjRPJRT5OJ3kLns8InQ0NZufJnDxEkKu
CfsnoVlCy+w1ehogTcGfWRcYxj8xI/++HbRIcG8g5abhS+yxEJ0mSfTdMc8yFY+8XKvtAt5xyObf
Se7XHfe7fFuHVqJnjcXo16F4WI3u+doZkX8tUypduLSFhBWWxezkofBpAtRZTAwLt50nJOB659XM
2E6SUdNGDDh52W6MVlkBeFrzGvdMIp5EqsfKpL48+BPvADw9Ehe7ynyMTU3roi5sXTNEvhKtnXFP
FULfAHnL7m4au8JEliaZxv0gksNqen7czZbjN/Pr4lRFc5aHTQEH7ksfydER7blEucZwNUZgpBzc
j7P7Q7jJPUUEGpUJ7mgS6a8A5VOqjzpzqNBSxFLZjHlW9WPQ5iwuyOLZ4r7SiPbCmtSroJO0D6zS
svlrVkuFu2IdlOy/X3HaHTs6y1r3u0oyn6mFNo16zkIC+oNahpLtxwEQg8nJpja36bamM+JKezPl
qYM8YrGOm0sEZD5gmcNhKfZ4WH82F0UzyZLKoUqguS8uPhS/yUrgm7/bI6l/PxzFIg9hMOKnzZZS
cIy+p+3LAqTGLv2GlbQr4/+fIa/7gYt1BdStMXwsjq/hEPSm/6TEU3Gje0u0kPDUq/IRAu/9ox9o
jO4QwbrINHjILV7NhQKbR8aCO9gPG8O6lp0b5LFlEm0PNEcHqMp3somWLoUX3EXb+108arLh6sXC
wW0+EomgyVCFV7MA3b1C2FTuYWjvKr3gXcBq3km+ekPgYXGlg4bfEhyM0RqLtzYkLZ557tS24Kfq
Um4Z929BLAUVUH6EzwBaQq+YBcrFYnmwdg8vs8yLpM2NjE3VG0QB6G8Q1kCDmkGhWRBe1E1vtwl/
MJ0x8glm2uIOGPOAjps1jg/etUe87DFJwQRvLwQ2P/XTCMnrm9UVFLOkzkluieF13mASsvh/bDWI
bkfgDqMmyo6yvJah5omvAlRRtOumFIbOKX9Zp+0rfsD10VorfdFqEx3/0DhFeV+MEHhcLIyzAcOC
l8f5UMPBkmXdhU3TFxGBgOiiGPtFndT5mA1TkX9R3r/I0zZeb1aycxg3Ot8uwVo2PhBr/gnj4u9q
fedDen6ICdjpCxfVfBEACpTf7HTMcVx+gZhyWPBZyTS7nB5G5y8NIVxwCQlqe9rgX1PS62qfbL9a
SQJ+gU4FBJzXSEmt+DIxzP3knOFWttaPzyHZmroO7uvZbtppIaNI4bP5oa01NSfx9agcIjIDp0jw
GLcfXDeMRO7UDGfpu0/oh//snwcN6sDA0aIw5EDlWqNJgrethF2Gz2YSROy+9U7pOvQSCZgG7tvC
OQW1gPvBbcgCf4IP4YYBnznup8jk+2xfiAD9uTt/N3z/o+hn/eegoEGvQe8Lrue1QD0zxljeElMn
yncuNHkwXwg/mRsxcI43KlNMDedu5rTtu6d6Tb9GEXSahGIP+S7Gm+ZizEucX9t28IVmDiZ2KVkF
OBwO5NN/3Ys907zYQ4G6BXIlkWbSz3nEU9nvOXUHbL0r496SfzwROu+SmQdvm/JzhpTe9BucHG6k
6Wm5fUh62PHhQwynE3bkdUFJRjwr8UjhMupSeLA6vjtx5pswsJyMJFBDCvVA+ayWv+FA4JSLuUtt
IqTiRtIFFLyTqhqZ8kOtRQ8GsoGGGLMO/c5BStBLUarZcBOKTYjdu8vORYypV4XCfHKulJIR+RXW
fDyh+DrdP/dM+f+ivPJgPB7A2mlSEB5wSLfNoEdut1i3QfpuXAYBwxMbY1CxwQM415MBfHgYgZEM
YOiDoqGTRRDmKm1h7TiF8DqftkNjQjkyCP5lv6u/+e74wIWJsLyZT7MgS3MVM2QVwh59dfakdz66
edvklHgF7nsCohJAVzN8f+xXrMUB7PSP1tk9bcwzMUNVcmpP64JJqBQ/t2HaXGb61N7FLNqr9O1B
Ml9eM6QwxjP/NOgiWTbrrjKZhdps6GrbaGK07Z/7mtyzZ83lQ9qNaVjBa1RFzXrejHVfTiFv9LUH
NVQrZt2+p22UDcg4HRzBRFY+XZsURzugTynOEoZQYInxGmBu72D9rgS6+Ltr0w7rJwjWMUwlgy/8
2m8ufM7olT5znf1Dvdbm9yCPa38NE4xgCOp9D5djalvR/M6DzYIL6xHBHjV9xKSX60Yh8mgIYmTg
0T9y7xNYZj1BN+oGF+gAH3HjblU7gaLtSK5TfMKxJi/jjKHKNOMBBx6YSC2ITTNyMTg1hvOPIUad
7gPj8QHR1wJ3Ugw0tICTQLFEUvDPnGSD6ZzLTfITqOha6mI2cCrpvKi7OiDpyjOPkGQ80pgDZ7gp
6AYqIVB7F6Skk0Bs/pz2QeI58pCWrjB2uF2qF+eQkc8CxTNfhzWjv9LV0JYd3AxfVbtG0QEpR9kT
kJvuJXrHyzhmReFm5xC9qYCrrXbDyz9xXjSVlSyFhZ4RqoxBEjaW8Olx08pdQhJ5PHj5tDizwLhd
2h9hNSwgPJqr8I8TxQQAf06ekaPROXfjJtDXzVlC9u2BkvfPloKHjn+Zuwjz0Vjlbg/bh0xbZwPL
7OlWKGAKWNc3FfpxWl1Wo4JY1MxGAfRkb56yMDQ2IWNn/jvM3miKAaFkz4c9UBu8NfE6UKb8UTJu
l/tTJGDfpHjzSGHMTMQ0fO8mVp894Szji9gR/zJFhhsjeF0pwwvGepuZEBPm60w13mcZWL6+p08o
esUPdLwPPQNdW/ml1TRTmJwvznNYM47mE2QKRVI14WQ4sRxCJnbOGA7BNAX3GsmRsDds7UTNxP5k
GqCgKiCRIW1GtSSMHVd5pvFF2hZBkfFtWACHf8AtW/v52oj1c6HsD64xWYEUGDI9p43JwXBS9Lfx
Ihx1JgJdHluuGuzTky349XGuw8C1h7GhaB7udcxfekqtBj5rfMv7of5bfNtlEw3RpulBWjKZuliZ
uTf9ePCFOmELovrlwDmUGzN4vY8vJMuH/xuLpQYEUTff6a4zaOQzuS7lGseRsBp9zSaO80M6+SZp
+zdZJG0f03U5lzHQln4cpeGPGzIQHcoqX6DnMoTh3267s2wjkEp6QfEwAlDf1++i4WAzHWcXWc2n
6SRrur8Ma1jp6kr6zqG7Knclr5NQ35Cld7USCFMA9rJcyIhvAYvSwiYBhseLUb7Z2/AsGg3KRuhQ
SbdM+ZwiMXf1cAoP3w3SEqIxkYTJSAfM8O9IlaET+IWbEbIrFcdCMQGfuUIVkPt0vOrayWT2IBnY
+w7UUV7F6C2HK2PrwcOvqNwb8mYwaYYtlctCZ3QdE+YgoPSvdqRjKdq+qkkonJ94t8RXgu910/SB
aIzbDlqxZPOvld8//3erwogZuEg4jayyBbxoOMhmhjk4paPqr/cn5r6/W04YMtdTpdQ02KnIKPNQ
Kc1uhamO8nWvxR0XWo2cWUY4PPrV5RavKieTB4X7GWGj65l8N717ats7mwu6OfGLGHioANZKqv0Y
xuYhH/VIyVkz9SAR7UPkrQjMoConkOWQAKznVV74Kuwg2/00MvF9j9R764PcQFc1N+GrFQl4rakr
Fg2kAQyGxPol9P0JJsuzTOahP3zRmJ39l4Rd2CcG66YOFg4JIZBlJG9JTuI4k08eQXI3+R5Ez8Io
zNELoJZINTypIJdM0QOJylHqJK1HUhn7ERLXh0naIcnXQUpF4/Dj/AtxuXip3wNq4Ml9AvKDq2wU
jFGWqYrMN3cBxqMFWVg7/Kv4zYsEajhE5aPTzZbsZ4EhUGRN4UmEYKMtXXe8yMSrM+iHA7lb2mEM
ZAyajsS95/4OZLV6qjBbIyl9izChYgc1Qg/LdjEBU1fWuvgv+DYWwnygT8aP4KwbuEsGPQjBGNT+
VrBsuDo7ena8dyZ4HcG2aa+WaMY/qkgdUlyateQieS29lcngEmNQwlkeYTNg6VjhAzEXcpAwYzBM
/PTkfYKVvZCQuZZeizY/Rez6VLMcZwK46pjTduv+MfEmvGhKBHQKKKYC6K792evmVNgNq70b3ghx
Oaf5uucus5GfTh4GLLsin4xgAOuGGvl1b6FAwhFvrMVJ+mlJ51Lli3fY5WHi8kBgQuEHV2RKjpNz
YRHWYmm2/mAPRjRGWfhB7bhaUfJ1dPDvpORZskjDKOXxulp10zNE1wkYTGvEDMjUBLjRQrtO5mB9
rrbIJwNFMxrqjUZJJggh4Z78ffaEVOXc7qnKjXqZgrGN1/iOOhbxNr6ZOYAdpaX4PLTv/oOVLSFA
OZoCWJ9UTXVu0BWvbsly/6CCMsh/naVuXAhqfBlXnHO/O2tkYokb2cc+XGbbXOtZdoz+1EoclxLg
TZ0O9vfXrEE3ii45JF64ndH6wZ3xtgIQz8R7Ha7y1nz9ekfBHAWxH3uDm0EGAuD57eSqXfEctQRf
Icd89jBgwnWX0hYhCgiSLMYOCwIK7VjzgV0AScgps1wy5apDUnbW7zc33EywxIssdYC16JaN6YuX
fC7a2gYcJ77OOgtYMR9Bw7OvvhHOlC5FojQVRgyikvwkQwWi21q27qBmadwAGAv4aneHij0hs16w
FnxY2Px2n+bANzpoacv3fVviPgew4s75dtVUJuWTmF5pS1jQbJEksGlYkfduLaAaQ2ISOkSfPaGU
i9XHq/qOvk1NN1s+hWO/UvvF3txxafMn6WTkEiF4Guwy+ECewI/8HbdSULdm7YQReuHWC2uz7QAU
yDVCEgOfgPvKfNWIwUI+ELL+uiFwfxGL+av8pNcYFTVWI7oUfIewm9IBq/1yjwq2mmGcz89dSHls
AygiIzdZL7ZDRZpvXnONOM6guKoTVFeRzLFsK3LunwEg0XfpWJsyLwF3iHMUaPMPVGZazwCCKv8y
KySh6ritzvTqFlAOURkCaDmQgKB8KuCb/xXgzu3DZ2ldwdZ2CFS6gNCaqC2EmyAmi/GSEp32LJx9
cYJa6M1oKuuRd/BhLa8Uf07vK7PVo3L0f/jE2Vs3X3jr2waLgo5FFiLv79oBVvRhgS5YtGBXgL3P
2ZnC9gsKSriLt7dn5d63rhyPjpHlET5TqRucJiMobK9i0rLVvUh6Iyv7QItofd5RC/8UgLPBigXB
tRJBvP5dYm9k2DrZO61IAFRo5IBzYkd5fo49KCZP6ii6tbiOmiv15PBN4REq2lZWqvfOPMaHHHH1
9rUY4MdZ8lMes+ttuTj5Ki4y07xkMTgokVCsGmH7cjfZXJmYUtCBznoNjR4BPGdWYD7ux2dP0ypa
WZ1aCF+py2GU/IE2WsUmjCvzj1JcbaojFX1DtZqRh4lv9ob+DMZbWjugrBOo0ybzwTGs3YIqg85U
6bfFgGeIRF3+j45uPD9rRXAjm6IDHUE2C+2Ph+OwuLOMIwVemVkJbK8hcJTjKSrRFvD3V9Rj9UES
vt/jMUzGJZl33GMC1puSUvcS13IZ3nHb7ZM6MQ7E3EF+jeq2vGfHU0UkR92DkMSUbvFrscgwgpx3
2Nza4iIXSplwJpII+Dub46oXwCKJkxhsHrRx1EMcPdvehczXYsw6Tb+Ixxc93gCUj2YgW02vgbGF
xBoN+nTs7Km99+coT+PyE5sih2T/2zAID4w5hmn/qxWa8ByPNhHdh5zJhhh87TFmg4ecLER0ewC4
pQG2vEpiLN/A+ZQU/XwKPdNxMXsLyPxo4lUw4FGRyCvZNuoxYQNgH8Vl3S9LeK0ZSqSbo+BQ7+V9
gmVnDev1BapNmN9SYgMbvmQBrRZFJQfowrrIl8+cJx42zMfniOu9VejtSFYxsaOirALFz+AVM+wp
1VQGniD+az8777eOwY3FOcE4rLd3d0dhhz+W/IYyplzIzBnp/m/lZTFN8NvNx/dUb6Eal+r8dIRy
w/WaciqIl2stSuBr9mbxQQF8YizmXEaxfxknoU+PA5WkOpx2XPJagzZRxc6dq0AAmw9lNUeylARV
SyXBAH2l/shuT4ntA81NcelySeArGyLAradd26LWiv00UDiDVl0uykVB0tfYKPB06652IVw0H2i8
dLfQYlx9b5tmqj21Nco/mjhHPtF+7l7sI2qSsk+kf+GLdKj3iDdXQNdfILlhOQ4YWmSo90x8/UmL
CJ9A6qqrwK8/0Ap7/pq0J0ludT3Icr90lIhNqMGrfCw3ThCXiQnJQwbhOUoF6SOKmphrDiHe1Id0
GyzmkPfUfqoyWgglOD48x1u0TCPvL6l0mb6xu20/K+P0pHYi8Md+w+K03d0k/eaRQiAoEL2fNYns
58xYJYTpz4jdMA5p6oFEGIo7F+21fWl6gCzAg13bpwbntCXrKP8kPaFkzJagOZl3NK8BLoa3G23q
6P1eL/yMbneczzIhDMEzRvrzKIBr5e/LsdOPjbI+bBQN8RE1jF8JSVv5LXI7orH5w4K+fZUlrnY0
qL4xOnwyLCf6z1EdGxbuPrGooAJRf78770GmPhBVwBlX2WcLVRFcJ6VODLalF71xfxc+ZM8jbt2s
hkUpmI+zu7gWv+nff+pWZHgCTNWkELrgfJ8DRr0DR3MD7vo3EF1n6r9TeuGFmC83lNWwFiwGonKv
skKl10HyPGSIZVhjAGdvPc4TlR7PS8pZjNGbocv1acNFAaKHEeCzfWLgp8xSK2XGeD34/Uk2jiTR
mIFFUhMG5G6sN8zcGRbbz/xK3z3UK5W2oNxDgP4LolEFhUEmb2dA2/HX5naMJhmfQu7nSUBDqHoX
nEibz51TwlZEBR6g43p897wmHPvbmuqADDUvVnAsQor8PitcriTj6z8uzHcAqlG0HmqLrLEPblqs
f8mVjKlFCFHpHiOBi1oyPgZWV9QMY83HY6w/OsbBLAgdZ/BA/dh412DEEq5EJGcmr8VdNefEKEH7
lute7dHB89SviutxGSifWHIMt24HLzFHpMCaupDwvLN0HfyrDPVPUmu6OBAPpqeaPvQGWRKaMZ4F
mBlErn3J0CuNgcueZ5FSrN+2tgu0Eoy49X0W4bbh++FVecAGFuWJ+VxvXoEhaulAe/+UYy+aP7R2
i4JR/0FwYjeVx9ivBnAMYpx0j78KUHKlmu6ZWpFQ05k4Vp+fNe+7aSNkiwA6MOqz1Ki5MriZ1RRU
2rGz+jJeRg/cln7VdzDPWEEOHpTva6oTqu0///S0fo8IXvxBJrHOf+2gOHq1THCo7AigzICYBgmW
57T/GfLjTs0aTe6WdIEkPs/mzkRcptBVdsoRWztztCAjKM3yvqthUWdm3sEvQCvwHiMvcD3D0uGa
qCnyuSha6gPh7u1yBJncRTJr84tI5MYV+5C8KR171JQGbR3dz4CmCpsi5TAXCIGwtLoUyXaRJSCC
QMcOSys3nas3dmeuTAjdfGZ5h5Ni25r4Zx3tJ4S9i6jgutVWFFNZR0q/1ng2CfeUecNJE7ztZxy+
zPayFgc/3e29T1Ij+aGE9eHLoBxqC8jUpfXpK8yeA3+lQzaptCSFEW1ElxD6vLuku6S9ZVtFPNk9
pH/5Q408/n36LV/E2Jh8zzVcutVLiV3VymLbOYyfpdtq+rxVauooL6Zq/J6Ti1ck3QS3IS2LR/vY
sahabxa7LCC3pznQ8xapepjg15T19B6xqP1f+KStm2sXquuox608Uxmt7gXLHPJ1Fsyc/LsCGHvv
O3szlGmCMWl2GIPnf1dNGVJuQAvjFpsmf+0x45UICN+UCTgMZaeSTZiimzrkq0GQy5x0X7Hn/EdV
cEfxr23agviLL6imLFbX3tqz96hH1DAXPzWyu/29Y19xGKc5zdys1pUf4iJwPhEchDDMwvulcFPd
qJeBB0Vh/NsI31dDsjzSqEI03K8VBeevtKpqu6xgnQb/GsGTCjVuFNTf4k8TlhkSJ5IX49DZhDj+
+kh/3kNoz4q8dVwgJDcuM9HnwPXWlIf1FM1Frfm0AVcFD+ibZ5nalmbrCsuhRBknHwImxUL9lBSS
7AcrlEDzId/+86IQrqX4b5Deg4p5TopRynZIk+idRaky3Jm2OHFgo3gS6tcOGQuHrxMgeJ61oP3+
+XiUUbdNQYvN4eySKpTE4gHkPvrdXVUVRWkZACVTsGnVmFxikVQRtA3LecPEZFBBvx7OolYCmRpz
O0ynfpGgbVYyekwLY+p6b7gzRqAE3hwYxQ4T/58NB7uEvymrnvrm13Eb+wkUHeZ07fosmrFqr0Q6
jVHFz9MmCBgYWm561Uw0rvhxA6TlX3bHzkPxJQtrdBZxv7tMffH9kT9lxk3vLpHFbcB2V4NKr4DO
+Bv+CtTGP1Kj7Jmji0djl1ulU59ec1YAVwuvpf4CxfP2gqc4CdZ/+KS8CkgURSoq9IvdAL3XJsro
LvPgWr9V6GnFb5g6RK5u8GXVWijljbftZtmqmOWMrmIX4MFomjs1bCq2IojwpDXHz4+SitOrkTrs
ZVjbcVQytS0CpqmFZGP4OanMTXI8/FhHeoBq1fAFgnN3FuXDPmnKGtORTVvCYK2X7oePzUvWroNt
7k0y/nTGEDxV0+32FW+tGGd2kLCi2o0P5Ea6gCOo+y7uMcyGVVUsj4S7PtJHCs/o9XkHnjkIKsaj
YkqDQQ9YUuHXudTiHSW9aEBXBqOqp6z/fEtDhasy4mEVrVH49SPV8WnlYABCuDZxRvq2tJMN0wqs
VcfkzpU9lihZwqxc9aaI3/otICWx6bX3zzTAhNSKu58O48Fe13sxD3NLetOD8ZIhC1pW1jUdrBHb
xfMWyQTBhvHmYU6GE4YVfQxIUVlBU4V24SCK3Kdyldnv0G8YpKIPrk9bkODOOcnh1vBr177AIAn+
RVWg7XVgKrFEiwW5hJsn99kalZE2F8OPvRHPzCnxkK5jinXotTfGcAKlldl0BrbeXcjFXJ0epwo0
MWiSKlj5MPLDfQxuAReQE6px2WC7vOz/QK1AtP6lu3jRL4i4//flzi89CBbxMht7MXyIoG0a2mvT
i7gmcZgD+l9KHAIuvOGq1bcYqB42bCNl7LOFSvho6USq2uISka+htfK0t49gyPYlrI5lWUPS55/F
KW6SlaxN0dfaDGXcYrBf1s+/W72/nv+DoTGCXUOaf4vkXAM6/PuC+56LD4DCMCOVtFiWr6zA3h9n
ow0IG6fIB5Y7AVDCuhl7SfIO+pXRuA5FbD4DFJ1MHB8Slo7cOwXruZBzXKytWd11UBJDJSLQhALg
wsS3Uj71eBAkDTlj7e4bGV/EPx64FSj3gmgiNe3mNoAdneIZuK80MZu7X/q2gA3HpCFCGP6nHeir
tFps52/Ft3rGNtEnOhXejpEpSNTVMLBGHRSZvIRtKhL2NdCuThvBDcGpy+FLA/+iv80zrgRzNiEL
Vv62Yt8WXHtHS4OcXe/9PG4C9A72asL5Kio2InsFZyvutVdUiy+FcQBzdtrT8kp8db3SY0qdqaQb
vPAcskvK9uWXdhnWGwTgjJPcGwnUjqoSFcuKzgngSI6tXmLUfTcZvnS+lzTkAxDXHZqOX7i0LQoO
fTmPlsGRQ06ej1emoNsGMF0s8dOiEtH+fSD8tMbZv2g/aIEYPuyD4tPp9zAJVzO/K0HQiBspnENc
wLJSi+n0vf6l/dT4rRFwk7rFoDvh1DMmpC8DdCOKd4yQT7jTv9J20Gg45lKL0zepu92PpUbbRaLX
ryall/O3frXDkNyK0kS7C0nA0ZfpGCGvWshnKQFP0AdbV/Z5GDJnG5X4eD09+8hIZhzO2abLUXf4
byeNkaIfML7hxdG/eXoEN6KnylIWey45/xKDRsaf5sjH5V9/GDLxb3Y41NSaErUxjarn3eic+M/S
WPsCoBxLQIE87Pk/YEnbkDJlxi0anTAZAbmuKueCx0M4nVUQa3yzdUEdTfPXOkCmnnqPQRaaFiAX
9/cFl7vCTAMDNsgg78sQ/51Z2EHksB3hbjCIeajpBAtw+PcXeDky8Teyd/maOrXiSEeV4+GZF6OH
dXQ/X6OzA+lysiYoXNAssTjkaLRleHFvA8twTV7OIFryIU0dh+gy7dSAiuQmrXE35WSc/UIaK5fk
cqqW/JLbHuOEV9HTFfkf+95gApBioG6yBAkYUnmzIFM8wJAwIAd5nZzwXBg+ajcLdB8+GmlKNHqk
Ev+fRsewrWxPK+z7/OKxJLlR9lvBpXV2iiP/cX4StmTf55ItfJavJybboVOeuno4MuxKvLutuOix
qngIB5BiO+Nf8Yqk+5xzpUsfXqEdNuYMeDcV38aHPIrsEYTdTYF4i7tBs0Z4+Yw6tfQo9GCJDPXi
yun6AOCmNULDFroJ5WgQ26rbb48/Y5V99p0JvFL+PKR5+jq8aT3oV+n1RTM3Gf3p3FyN2VJvTYQ2
aJXzQNKV0tkfz8V5xjdvfJJeDGIn+JESGXqCtJf32j4rhck3ELTuf0xSzwOpJU7UsljBwXAeXJ17
hF2fo0+9fvQ7Ce7REhzoMvWiLa0HCnjIwbd8Q663H1srkd+sS8g3HV/TBRsVDobI0Vz1dn7FZpZF
ZQJSWJowaIOQMB/+lKixAREalkRUnM9g6y45wXFvP7mfxIws9orpvImK89O9tJ32O3lE62AFQ2Od
HBqGan1gmEvFjX5vDx0x6JNWIU+xCe9YEjn55kMG+H5zPb4PqfCBWhm+b1Kt2DakjUB9vq3nxhpA
3xASoLtOvacVVXLaJehi8muhrfnAYaaq5VzfnAuRj6bZDKaxESLkMBUAvt2Y399Si7ozifrjZYuK
05guHABpxuv7ceqGTArJ4zlFh7WPeMfznZwc5Erzt2sqDRXPDA+k5JAE0xKGWWgwaab6BQN94E2b
HAJOwqe7wYXTu8rieVs5js/eYX7R1gt2R4WKQ4CkMn89niiJvyPCPDKHQrQ7Ek+/O5FyRSVSnyw2
d0M/XZS5vg88VLvTQ7+i5LVpQbbfdP4uLpupoj28CrML5Ri5mLYcfDzRgBG9K4+MtzgkbOO38ywq
T5cQv+TVT9N7EDvyq4E7L6rPFurcKdbO229jl3URljXZDcDlKlDAQMjSputTrymJub2pzOR15ju+
Myu24TuQO6WJZ58DIP6XJUzfZLC2TMYWaEPEKAYpDq+iujGumeOFEA2nRbJ02dWrtylfnh70kM8W
bcuPZmAgwgeOZJwo4N14lHcO5BE72GDTPA62jEtIuOqZeROjCX/Zo2KgqbIqdLMEVW1AXLqT6f1E
BoHTYe4IXxwTMHmpOJ2SDEt2JT/+dCpucLTsoKUh5Nh1ulyBSfEX7u3iI0uzPDjF6hs1kD4YdWJX
nVV12m9yDGLN27N3qgmipeCV9ZaoqsKtbQau1CaOwnywv6PrsTlnYO1+bB8WZ699s935M3G5kcub
V6fNPFOvUkRCdSNNdfS5Q/4FdAEe/Vwou/PxSkDm+Q4IeklAS1ePd7wkvdUHImAzfzN1X4KXDJtQ
f2es/XK7T97Yh35Jb9UuADXLi5T4xsyRGMXUOaQbbCugxrKFpdPfxBkGpBH2Jz3yrbwcbdQ+xYeD
R8wDxFbDHqONKv6J2zNlT/2lNHusKOiHiieuwwAmNfCSfUUSon2cuVxPXfY6rP3hHOZsaW0X3Edx
w/OPMre9W/7kqwDHB4arLAciSYzM0XfAGzPYDqkSnwRPIFSyQHKyLpUgQmclRaNNWyOeLwpw810g
HNHgutSxRFN/ecv03tCWEteEA3HpTmmkP04fyrff9pWGJSoRQJSOnSUNZFCkdDlGcVPYG0QUPPxI
1JmcM9LmYKpmiu+2XN8Ak60MZN6+GCteIrvIUKh8HMFB1icQXDZl5OGcSuDUxrhqx68u+eSOjgT6
WLeaKFwBJNZIps8CBGxz4PlsI2YC+MJ/hb32uCPu0XCWYIbr+MAQdifxuvg8tILI6eFUKE6AQCh2
bTnQ0F80ju/EkjyHHze5ekEITkiTAd0udfePIO+17DlmzORVOAEQsr2rxmALGSkHzQ8KjndYOGwR
bAzGxzXlE9ZgN/ZIstMiiEzVbqpugOzaIX6vbEHCETU5+cstASZAmSGp7pKcP95NT5TCCxBNjmND
X+82FdeXSPQcbBiJzxJfUEG9CZRz/9L9/qoa5vxjmgyWrDjkwaNJ64J6RCyqAqNuhyZUcCgSI7vK
iSqvX1aXjGy7kwhr477NdxJ8EZmcCC7Orl3Iucny1xSejRjy33G2kvqdSKRs3Y828FM5WsbcX6Xu
joPIJQgV0W180Bf88nVeXE9kkUk1WMoJmuGMoNw1Yn8gcLyOjBtDhzOiPFE5PkHu/LLZtIYw+L5P
k0zc6J6udiUIinS3ARNsfwJoj5GTALif1/Daoqsdl632ntk8inO9arBkEbvmlW1i7YqAs03GgjrL
G7l5h/YQR0Hl0wApuHhg4iIFmhKGU3uxuhl2sZblvRjyJHv6npMWOxFfYrNf3f82XFQ+fJYBZX4L
EXn/sSJxdbpQwwCHn29soLuuJXpJ+wZ/oBvLyveG5NF3rk/48zwKcFHZrATQ/n15o0iqGyp+LiOr
9bRUEVXrF/Vn/dONDp3Jad8pU4tAxCjJyyJyrjia7PiWLBqTIyGshl5yOVwaX1c1GFXguqsXsWA8
jrV9smsF+vm97RIDR4SbR/eW2Y6MHvAOFnxfp1DPm8TKfToQk9CViU+N0DlWABZNVwDLJY3Rmaxz
z2OIcT5HGM+aSh7ljt7XXvZEV0Nta9UTt4fMZAjzcG5zkCMqNe+0r+aNiEhCdcR1t9yakUMxHcVi
FKPPT4RabeyL3Zkf0/W3EbxqpAJpkq/nyLcagfxwWFb3ep4JIxSkVpP5yIikC/lQYAvR6lo62+yd
+J4i3lVO4MarIKRRk3gHG23K/0zUPyR+IO9KxxqkES5OYCRKFfycL/19rXULaiG5bT5TY0Gnqd9c
A7+T2selVqr7jHT56htOvWJXPUjRyRtJeY4QiG8kJ53OEa35jy0sadK2oogn/BsJL7+vX8B1d/Lz
lWuZfKyJ1VPl0FPTKqc1kSaWX9B0cUqH5/aF6Ec/7vLZNgFANAWm0T/TmhzeJ9k2gXGwIdDJQ4vo
nxGvLGmo2BRBbVQrJe5Tn1LlyGq7lHjJgqjby8MAw63gm+Kxuycv+lHLoTwv+jjMksyIdgg5Z8Nd
7Yzj0hg1xAZr5JktDmivTqP6q7XaXIpEftCugtEy77BkWym6FTZrKSJQ7FbZSNfE5gCO7Wqa9Ucl
KOmXJvCGABrrNkt9ZPtrNLUXp2S5zj/+7KTVbheziqsd6dBbxgLzP6naIjxeCgxJDQikAnnNhD6N
v5zRs6qqIC59OLPbHLUgul1ITB9882kd3iHRy3AYDQfg2X7Iz2lWRwSgMLGHxXwB5jpMueBVI1k9
52ATh5rU/JBrPZQsmmFr0g1evWHvGi2ygaEfBcHQMet+G2vG252CMuLWSA+Y0VubCNDiJI7GfKzk
pfeaZ51W0VgrbOBOhE+SBgGhi9/ZjLykkpZ4s6aQ5u4dvyDEMG9cjMLsBbz6ykj+hQdP97omkjwG
cf+rllF8mf+yrJ09gpbPQ/EMjNfhZNXdOe2x4ad39t3KquJkjJWiOxN0a+2WRg0F8HRdhoPQyI5U
nOtsW/nnPX5rZ9/f6gSgq4btlAjbpVAu1cE4lOMWtIH9Mk1Bb8BmyHboslv+ZDQJkiV6jGMwjdkE
96s9DiaNKQwJkdKzaIhms5OnuXqYZFG07EgI9y58YYVj2vOWrpp9G0Ocns929lBF6XmT5yq/mXbm
8/it47oW0O5639zetaR5H8aeit8KEUfPQ5oRu3IzqYInYRlbaUacHh37uHpJDE/+TMsNbN4iZSBu
/vqN4OxWbsp2U/0UdBvvcAdaviI6B3VzpjuF1d4xHt6HcEPxy0tFIMWN4uJ0K1y29o1+cdxH4UsY
7hbKtVMp6ZAiI1gH0ucqLsjh0Qtf79A+vGxEVszJxGeCzG6b6EkGKUiYnBowFUG1FQ8N9FFFYldf
KzUbRwRKiv2fBtJeigAi02Q9dbYb5IxSmjV0a6sPwornk2DkhTPNnH7rgYNxqUb+ZDIlB5HJu9/a
MIy9wUwDqGxt9+BlFa6TSBCtybNYrMEzzzr3TsWn8naGGPVIVeF074h2dt5hY3YdkngmRmpGj8/x
O7wz2Acr443lM4L68TatuAIKh/wprgXIDWG4X/x8roh8mE5FnbDfcODB7sS8z5yd78vQYQ/hDl+m
yY+wGcjZ9QbV9oowLBc8mgRWThbwICszMTOPqfxSTxNMNDEO5CAdMRlPkdv0rRvRPoemxWGhmPT1
efoO7dOs8tQE/MGoW6Gxn3uXxzTlkm4bvXTcKXiocLzFGOio2lP3MkImWI0RNBU0dCbtVVFUoiQX
TfOoREFNo0Jr3x3kHAT4TXv+Ank3WZp4qEBR2alSxqMB28eTqF3hQrhSHTmKxC0RgDIhvbatiJ1R
lMf2idci00BPBVHcBwBxNXTgC18+j+AiSP+T/K2pNTCqdQUoMrc2ljqdw07OeM/wnvOjH9Qe0cMX
rKoKOltc5oiOcrZz39+WjRfwmbD7PSOWQIBxlEPbFbg3JJJDImjPuFPLkRrbViwudY1A6OHtdYmk
fAaXeAUEXbmzyN5zrorqyQYvNIxfPMYadP0aEdqmcZu/TATa/kANNBTHs8eBlNwrUnNT8OKyloo9
8qmzlOaHZHky8KBCV0fIm3OVhw6pREWVzg6zNIKBuhpN+ly06oEnt6eWLV+CbDLr5bZNWtQm5+07
GCHJKCpBwS7ekIbSpC35OUajCSwtEdwdUn9HMOvFAaJi3J6rpPfEkRz0+9q04MotxmCEIBQaeAfg
bRsG9P4oHam6fzDOswffv/yze6LEuh54bBXvWCq1mwkzijrMMGfxyI6TYcVA1Jchk7RKTILNv79g
EsIHzjJ1UA2FRckNtlzJdE72N/P68N6OKG6H+mOmpmCEDaFpf3PDd+F4EmrbdF1qrOmd9l/txTEa
ByEqm8aieQDd4pLnkjbtPaYt54JhGQ0zOcX4iabp2WCabU/serze6QQVQS7EU6QZsj1o6LyFsg/M
+28pxR/CrRGv3G8IIuJwg6+5mdbMHqsG0RYmAQF4mvbyL63oMDh00tCMsO+uqnTIuTPsOGTfs06A
53tyfG1SFcpF0fUkHU8dLG/ut5VeYTskJJhgyNhh997VnWgHIt2hIfZbl0SEofCTz04wzeg5Kj8s
xZMZQiLSxwqISyGjKon8xMo3+Er0Hkin3SECY4TLl87XwiLXs5w7/6YT+1O/+3GgJ9xQyxqQ+D5w
VLphzRD5ENxjXcJhx+3wmZxi2KEe/7bgB4gXc6/k3bpkILIftewB5T1bRjuvpX3gTa6JO8awviLV
6gMpRgRZhb66ioUM5XbtlbJidf5S3IUbAAmD6REBc2JIZuRyMxWOv4KRlF5FQddWHs6voUYkGWjO
Z6f/JdFwauPCvgbM8PLR7kqvjVpbFfbxCsSL2R+Yc4Mtm3W4r3kpYvoycEgkarT4mbaH5L04h2s5
g2+tu9vjpMjzaEd+Osbjuo/wjOhTvFJcGTdjgHv9dANYJjmvGrJb9M9S4VrgX6i6wZDV33G7UNcL
XoPT62fTICX2VJc83Q4pvc8k5JWL4jvR4GBDtvB5czUiNuDwg7wUQqr0+yqZqo1Zdvc9QZJy3oFm
JIkv5rOcMuYN83cZAJti3yBHN8BNbrSO+yE96gphREesI7RsLGVt7oIELEmw7n/aMCXEEZADG3LA
wqzb014yipePux+X/kKFaZ4B+YihBlrR1Fk6TF/MY7EKTfn+p5F/UwLESasUvIVLAhsN7XQt/egL
YeVyfe0vP8OWAVYqCIkcYCUzAWxDUYAXH0LLDNEmTvwgK9Kq+AChMObMZ1asBJTcN3LZ8stZVcXU
bGOoXatFw5mlAuIGCaAm5xZh+eQXaFz/4vm6akTOMlqQuyQR27L0VnYshWx4a6/5NdkUToVXc6Tt
/qsbOaHeU+XVYa9J8mYZQ/2ylgS0p5pSebq4unnPCEZv/REIHQSK6QJQ5UjIYuLpKTiMWNCPQUHL
QRYLvWS9SJZlxg4XOL+i2wL7ecVs+Qz7F2SJkS77ame194Gyic1+X4aRknVNSPzFA7U2y558zuCK
SIQ2/O9/p7q16ZU/ApWxMjirNIEN8YStLCC2TSsyMoZ/qnv4Ttc3c0M9ArF4P7Khzk/ypEWaHVvH
FYTwxLrl3gKgek9s4rbtILtd2kFtEzRCaqf+wK/m07OLAKP8HdXGtgFjDOWa/WBv508nssWmzmJS
CLv9gAgVG65OWvzh1edJpmreNFlaLhzBY4uzX4jITPMW6fPhOr+PhILMd6h9PuwoyQjiamyMpH0p
jAemvdz0pG8gqGxcf6bKhOjOpZ07rUEfAgH4izMrQ5UPIVSb8/+x2aaJgHOeFsjngxrZnHTmyiyB
EnWMHHWwVbq3MnZDOnRsNfSA3TdB21EaOnb78DOn1X4+wS1wf2aFdAx3G81eHTTcHa5FCRQnMYLe
jhMmZEEglsGHPIG4Q4I0ODm1y9My2GAvYK40KqAkKhK7lvE5pWEZR+c/18iHQ/B5ZPVj31dcFlcE
HkTqAwKtjnWsNZfRd1r6LNWg0TqOczXD8amzz8ghscG/1OZORAhrpNEAXGrQisz+/eYRZBYyEPHr
9I4fZUL+CtpJa/0/G8KmKacB+foG8abMx9nZovMV5mHgOBZ0u4fRVHB4HMXz5Mcg/dzkMmVZAAm+
vsZXPTH3wZfDPi0LjtAsHpmZZgXVQKa8qjhbffbuM8SZzCv8HPs0CW2nxdh5gGr9y8jsZo9ViVHf
pUdKpagbpbym1UkvEZveBE58jrZROdE4Kf/jElKQm+VPj+I923qNP8iWMahLez1k6wk1gwEgpsR9
VM59d+duXhCjD8tYo8E5nGCDYFkcO6/saOurwMn9LGW37GslOVfqAqFLuhscwMyExDeuA/szTdCX
64g8HtJ+YnjkKt9EU/4AEBJMkmQ/YnVM7E8hkFqXYkLvvLnVFo9BY2/K6utaQtZb4hF7dMJ1jrGi
E/SST/T7b1Af3jAaeGlpuYZN+iO/KuQxP8VRbP/uWy+SwaMuP7vXwMdctd8QyWS7JbzvOuK3t4m0
3VqEXLsjQVPQtEJXEU5D30nsaNTHJDIPBjM9GFUZ9TxnME2087J01VrhW0eTC3TP/TeoTKjstlcW
VCrZ6RZMCgfBGBqdPPKWfElHauPTVXAMS3Sx6DpDO1dRYH0yEkeIUWguUc26MHgW/o4bF2KANzec
KWGxVJFIqS81MdR1o2uFXFId1zc91guH6e2xLf7HIpIOpngccABkk7XWK9cc7/8o3bQ+cBd6w4FN
MdeljScg+HiGjjU/IArIds7Lea5z54zEQOFwlefLCwQrtXp3Gr2thgY4DWoE13m0VtURFda0UMMI
ujl5qqcoAx8YeZze0nd72uTB/0+v5vB87L4pzH/rVJptoVTla/lA4Etz8gi6lMMj/9P1gYAm+7++
wpU5m+tbXWA/ILmdkNriJWLp2FzIYa9AJZfg/QK3HS+RPysmygcNZK6VBErmov6tsxAbcnbtreRu
tQQLXjYKSz5DMnRLOHrt0pxNXbium6aMknSmv7ETEuHT8XJMbL4yzvtQe1/4Ag1uSgWe2Wy6QKhV
8ifpmxjLXtLLOGmNW3zKcg2CzvV9ChSwSeeoRTIhCnFURbXUPSYtGQ5VKtiqAK4pwCaOqviENuX2
q+zFJnmrnW/i2y43wRqj5Bdj690xd5G6f3/6tGzJWwnUYbwOL97L5RIlOr51/M0b2G24BFplwo2h
tXL2usB6q+JfJD9ttQU3rmSKfaTBZEOFKsdm+AbBKNzJhchNEFsTWReFOh5dOlGipxTHofNs6mX7
OJ4NF3+Xewqk0YPddLTXz4NZjhHqebuOjvatIqjpNM9GUVaIAe2+wtH8Kc4z0RAbEEGOs4mxhvR7
E6lQcyVwX0CJDVJn81FF+Q0fkYXgtOLtG3MgzXXiqu+EuH8PSOlECJ87gWRRqK13/iEAGFhgBOl3
mpenh7tLIMJ8JWDfWWSfwu/b099wLUrxKxmDk7n+zyellRdTXU8RsUHX9bq1sZV+dS0XaN256VK4
hV+awAYVhoafaNFJNJWMYRxhGwmZh+irHcl3xWWTNBOuqHhxRy3vZZ1IWwgwfExizNp5dJ/+ROr0
SYoFOmqr642Hvg75oa/4mCqkR0l6/6heauCX7Q1fZ2rJlAaofXNccRUoKn3kwnKY67B5tFj3M8xm
KHnv8pTtXq7pq7XIypunSsSDlFUcCJFSnMncLmNCf52j1F4ulHCGLfRiYj96DglAuQxbCAoZ/ToA
3Ty9ejRcAok2I92K987mRF61T9KVt3gIQorxzOTUywJdi3jMHKKiF92dP+L7swDexbf2lE+rb6fO
FxBdqQKwBldAMdiESvj/4pobcrAIu5cOJSoCydSW+r2Nf7Np0yLJYBcscgNq2KWxCqhgFAzjrSNN
jYwaNedUvyoog+E8rvSmumz0XGE3mSyVOztm+yfLNLfn2mjPTa/q6zUP/FiwCqlfvn6/VUdTzsiV
Tw6KQD1DB5fbOHNpiTtGvBiXFJJh0GARBb/Mfa2d169mAeNAyjmUUy/pEUfvIJ++69gK2abVv7xb
Xmn6lbtNv2u9DZ4DCfvavXV3dvICzhLbDDz8DCLPflsgrPJOFugZOfFFPEnSSgjuzzDbWF/iRsPU
pN4BrxRRdk3nOBigNSaM+gmO5HWmwUSUA64UhDvzdVTcAEojRXP2JS8yKXkUAczHilN7Rl9Y5lFF
uXvC+7Eua1KRcTP16sUKvBBh+9kxNzVEuGX7zAc//qLbsW8G1Xr84w7zcR334c7OcWEhbzu7eZJl
mHZNc99Zzd1SvFCRGqn2Gv81t8n8bJ+7ecGevhNDrEI/H3bvAvQTr8wD1V7ROIdiSx1mJ2a7jj2+
Z/1EY16TMp+aNDSG3BqR0oIHJDAz56c9QmheWC5Ggnb82z/vNcxQJhhOsyRj0In5WIn/jFD6r299
6u6mClJpnyssVVs3o7j2XEWdL/XihwH4HZHEvKc4aFPLK1HmggeMY1OjienK7n+T+PElmDhnMShI
wLy5M+QDd3jjQlmphmiR5XSKzcNO9S+0eMfKS3PcoIwgP/giHWbcgVZ3hoV9MsJ3DRotwZTZHeEi
ccevupBz6zYNOeiBdyxJWJPLTeX9BEJ9y/TiYf0iff9f6EFq8xA8NiP9GcZEXsXNjQLAkHeW048C
v8iyiaQPaSsYkrV6kj4wMs5eP4JJQHW9lvZbTFwikB0E/j14AOaQrmx+yMpSWjWjb8c59wEBadvz
zJvwthhsn0Vsg72fa7vvvm2T8hFN+m8WgSwwsNSqXyI/F4Lh0qHKJ91ghWWI0AR5usdzGj5pusSe
H1aWzVU2KA4mX5OZ14B5Jj13Y6c3EuHm3LVIc7i9Jk6Rk9g2SOfPO7mi2ROwEnh13oMISdjF4Thp
+5dTElTLVtSltV857OS5mCg70oe9AdXUKx7GuH3S39VkckBP+Lid6ATNXre/C9qbbtjVizxAwz2Y
FChlR5f4NJjQtQCFjzZggrWkh9BZLTjqSNGfx5ySndGxDvD6xvlcsbom2M2MXB6byTtkGMJi7E5/
WAC1uBG8z7BQ47KnzswuYY7ZcQY4hwirMVl6q41wetZSkvIOWPpiGfCUScrGODXbzI7tWQ7L7CHW
7xRuCx9WBXrqOzUsMiE6204j7eizrstQPCwHPqdkeDVZlMPSbpEGw0GZc9aBm3U2PMhxSH797QW7
LfPy4biR0q+gi8iVJtOlVRZo1Tj4qreONz0qaw6OzswkZCKMMeR8Zuqe9vD1D3/MkI12VTCfHzNN
t9sx6wL88bTmtvh3ipvfTO8amFbOUTLId7mHaeCOFHOURKGzxp0eRF4CDycX0sxmL/uf1QvWK+Il
h8+K0qceI3ayW7Mc5UPvglB8yo4SwOgSgqUFa+wAethVlTocq1ipDCUxg/ZD3fhREaNjR7lVUsTC
EN/fjqbeUWnLlM3KhxNi08ZX1vwZAX6nqoXbbwUcGcgdolC7LpMg8Nl8nKTBs899NT2NGJT3lFp9
cAeYUevJNfFAuHUPeYni7H9oiNC5f950BXR5i5NHkIICqZlb8g88iudPVMP6FtyuRYlzM+WJPz5F
VxOmKHUu2B9qbXV4KmVtKQVCl2HrxhWlIgsRwah8hFCHjJyMFnVTIZKAfpisPVwE0/0M55P6k6wS
fxd45OHAB3S3E/jTwmUXijC3fwOkECMs1Ry9E996LzCP0988nDkevEDOJqB33wN+Yh3NuK0YSUbd
u/6IQRWgg7DsOi6yUVI0Ax+mPJnFWfcn0GRVo+JyYOYh3SktVMOxYaUpR0liaea2oE9O0HS+N9o8
qnMnqrEy9TzsDRp9meL4VMnfB5Nui5Y8maVduSQJryQ7L29pQi5nPBr8x3QQbwor/6jzvaWjnUat
W0SwE7mSfzbb1PJk/aNtRInzKUo4dWNgoSW6XVPGqy7g4CZyx7Cu0sdv6TS4hpH/ajyUip4CnCws
QruCssoeIjDMRz01IiUOWz/THUo7Z09Wh7k+qj5VvhX4qbAn5Roa3YKE4No+yqY1Q2tnuT59JlG9
i60B/AfsqE9z436j9qUqZ4BwtTVv8pOAwmtWSGb3EreCzdsA645AsNyTESa107xkqK01jK1GsPr4
GGx/tLzMqZ9MfH6BI9MA+dhrBTAdMCKJXOme0Bz0MRVZyN21Mm60ZajK1BNcVRLLHZjAQwzyT97X
I3MpLilrD0d6PY5LPJttVeGVBLGGrBkgOG0TgDGOvtLRME8grhljonp39Wcu1om+F76yjtaOFmpG
ixBd16AsQ8ENgq8/H5qVfN1Z1ftZ5FxuCjeUR8E6r9aPXXPKkz2JwDdnVp3CgMP2eB1XQykadWEB
iBez3hodMuwRJGzfTDGqZFSR/LV2f2nHlR2a6k20ZQCOWvpv5gjQbq2C3u9VJWKzV+WaR1mHcY1d
Y0mP0/45KbXxsMYmkKVd6hPsJ3IlXx4g3ukO4QJ+QGtqHLkbHNuSlS+YmfipNi45QOcHZSRf3oZl
JMyuyqfRsuVxUZVqZrp6FJx0PMSj89etdY3mzk7mWfyLMkfQRbLY1l0ztqODUaF4MBBWsEj5cG91
ypx7E31UVc9v1hPQq4uYFhD1lG/efAVKUb/kNVuG4u0pUgm5AXOcBZDzS4V04XkNPDNj4Qf3jJEi
cbeqNDdlHpTxyvvnGh04bDIJP+1FFCQ45K0IJ1WowYYz9LK6qPDPYWOYZPHyu1PZmpbCvH/Zb+tm
LTpUto2tjzwbqWWX67xPsYNbz9i64+hWIN1wBdXVrFzTvViHEdryYWjKVKO7IBMYFU2TMfPhxz1q
WzohRcRqpONObrrlNZP1/ZA+XQf3n2osSJ44z5W7FLSpLcNFSW5wKPrTxWTtQ5YJ1xlfHTKY23FC
cjCqYtRGtrUyzE4sGIXtfFpd7j9+wq5kpUh6UJ2ShlrgzHZuJ9xHPjsEdHWgYTW1SGBfh00zLhBN
r+S5OehpLoFYCMO0TINSET0UY6TbhrQ2n8kGPEFbE7P1b7GhYfDwzGFwWLluMCFiGZ6lTbuz/K2w
XUk7DSmnb3uYZHydSUwadfcre7r9vpmqDLk6SwV7h5l14NbUzAHOVyUOv1Be0HdwF4/aklI3lHPF
tnhB7tx370j7K6x0UAVF2obgPQQjUC4Pitb9RpBOBlDodP+g9uTpUqNbYYj9V347OdaHYkAPC005
2tzwRbMEE9IBXexpE/tDIqLE+YrsjXvVEbDu39q3d/xHb1mWfUV2n+kekp8373LszFcllInppa3Y
Olorxi09CIzqcqe56udSSrhSdLJVdUT/7UX5z3Sc159wNq4hBkYcR6ZTed5i59eDG3LHs/nEaDa3
oW0a1Aq98VuyFjmVzqIfZ2xTZrpP4o2lMNz16nBw6XHFK6oBlFZUhREKVEKT8tLrnVaPnmNI8NA2
QZsrnrxhrE0VYHoo98n9bAgic5gzDxIaXaI30iK8WjFa1Fn8Qm6rk9bXjRi3uLnGsWkN4JK0NtgD
YVeCLCFk8TzeHZOQ64MgN3+6AkVZQnICiebde+yUrRYZwhmTAN5Ovi2IVnUowuqWCqYzivWAacOo
9yYFZNLWgRB0na9GyX/Kpl86GR+VSDYCNOY8NH3wOSRZViXNLpD4g0cO4Lkno6UzgpItnSjRQ5Go
ByR8Os3KbCntyE35+r96YkSWrb38Lrze1OfRXw5EynMGNqH7ezYgOCKWgEf6+FSmq3oagd96SEN6
JokiltwHD7zcdxdDIkt8jmWmMLsEWy0XQrvY0EnNwH8dfERoyZNBbredeNYn5Fcakf1kcoGZWcrX
KMUW1APoi1gqvKcSoBUZR7F8qqmwhhGMSaMtPr9uafxkgCV5g22XxVoOo+Ujuo8TIFCZdi7ViKTK
LQ39uJzMI6e12inAqn2nPQRFNzFILbqYy+r77X50AB1GXboz/VyNiml6atOI6jzYMIc8nrfhVxxC
+fYFrVvy/BqrNgyILrt21yz8JDO+DMnn0y38uUfRzav02QwL/u9hJfl1ATxZqHZUZBpCJ/B7zlTB
NFQFpK3wdY2rI3rEV+tBF08UuXRE6HIE6LmoMWxQS8j0A6+vUkzkNMDGs8Ib2kTsMCfuJYaVaL7U
twC65bjMKWs0tvkbLndnZzR7+TBVhC2KPTkl+M0alXLLe+215X1jIoREkLQeFIUlbusXz8kczBlW
/K0XbqZiMZXhk15Idzqd3nQLmqyV18LG+IYJMhtLmYECVLp2xW26/h9uOUDyqGiZQHC+EmvXIhfK
uG3frPZ+jEUNnv/8D6pEXk5tfXaDEiRBJpoyGptoiOlhkrIpCZdbVpEfGqgTNAZzjGcEWMNOgxn9
wTa7X53aN3iAn9kRKSemobjfajkI3TbdiFqS/Ri6XI0vypjReBS1tAv33Xd8N6ilYuSSAvj+qN0S
7rrfuXMoRwgFAZOD1D0G0ZLQo97maWoNK1W8vqxgP7Yg79JseI5ZYWX9C2AtmzoVl18P4OW3QSBo
OnfAGU3y+mibfIt3S5FJZ/eL9IpC6NDi1tbtrTQiLNuKmZ+CozEaom9n67fLo4I4ycq/y18396p3
PlCGrjkDmR+xvEok1m5qq72YSNlmAzJk6sTEpl6aakoDTItbXJAs4HcXXmRFF+OazQbuxP9Apxcm
kLHnSuN615Ju9GHJF7J1gIwkygDaOql7RsEHPH9o0uz+KApv4hW9iRot87c/yxvBe+wqNqxlNSNm
z+4sDoEc8BUsGtXa/k+5utZMKRCOafKcWHgumTQEYOz9mLVOMcVtRxDAx+VVyqN5Q+BRPFvMisdl
ylD795FCZdqfh4E98TOPQXA7kdgisl3dvKE377fxgnV5u1GTiJ3WBXt9EZCCJA52+ckXImtrGdzW
NAjf6NuJmu9qQjXuhwEzYXPL5rSw9T51yCvzHYiSuip/jxJl6p+o8T1IuFt18x06U6Jn43k6svkA
TVNpNh2jOWB8HnzkqNCZBN4gNdKdEG6FoHTUDJdQGTaYOK9tvzfW1vVEn+Ks/EQ3YjarEj7S7Ju9
N9Yewp7CbGT/rjRdS3eU5yybd+4+fn60Iab3+SLSuJKeYi7LmbkSL35nvocbDhCeX87hOUROGt6v
C+CHctnmz+QKvVvlJWmbMs+qvFVBbA+FKH5tCa4cXvO+u/8GQRGKt8UI99ubqbQE5BPgOKdIj0Dy
MvJrw/N7TSaoM0udV3xSuitecO1dDEL5WushGFOhkUshHHk4wdeJf1wRkAdyBazw3rqeuKfwOnjU
BT0ghDYIwBPbGb9Difl4nvzIj70F08mKZDOA3yxVYilt1rOqzA2uSAsvWO6gnAT8LiE8ecnh3j4z
8anPXKqRq5hnj/3A0H6AIHNY+IpOOzIzcnypSSJuC028nqnzgsamdakp+jsx6yNilMTF358QhUFf
Q22Y2gVBHus7lMb3FtcYL64uIa3sejTSQCsUYsgfeJCQrwE2siovl0RqAb9aLYBmo1wZhO1A3yFT
raCFwssfI3Wq9dZKh81E8vRwkKDZlINhQpTsDbsfMaEXim+Vy2TvV/MciQHsUKdYrLte7wFZql8p
3DiKxOnVbM91kN08nKTlf4ZET7w6zRI3rBr74S1cZCF8SvNpYHpM0CUCUitcXmo6mI9U0APAjuKE
jbaZf2WT5c30ZYzCvyI8945/OE8E9auK+jd8Y0weqSwR+Kh07q2FzA+TJ9vRmgtxYo5I5rK2kOgf
QCUmQSgB5rACJwreD5PY+Xg2nIABUIuKWkx2g0qgXx2ANQQVIdLXqFzedia+fVcWp9YRxhyLCBzc
GAc7l5VRtEed6tV/8XlKlK4gs0nO8iERqXW1ITxcCUHwaeVdBZfr6ElL+4RwCJ34patxOilYDSlf
0+5oRNo8QPhcNz6B89zOlTCv1fke+j5lS7U0UPNz1wlJSNAM3OGtMmGoPIXaSz61Fl8X3iIb5MiE
J9Y6XJzV+3dYkFFA1Hf9aikLkICPeAz5KhaJTPP0hnKSUY/AqRcjZyr9/A+hVOpxJPp5CySF5uEI
Yb9yGUugELdikEjMFzsct0eoSa+qwBXdkSiRJGfoWc0LySHCO+kl7m5nVftvGsAqywvCCyEZz89w
RbbANLtFUzrzgPOpNhHxcPju8W2eUKyEHwW9kXXwjH3DxkT228pmaIbbG390XsWSCWh2C2iJ1jtm
8ebUTzzMCKVSz7pQBXan35+5wXjdZivtmSMxJJbpGFRIkNw9aE02pWMmQTxIAnx65jkADmdxZeOd
lV1bOlNXlenufl1h4Kw3Z3HDOVkwLT2QgPKOKOJwTi0+o4QjyZiO66N/7L7p0vNQJQuxcdY6i1U1
yult8/ycs06nlo7HiXp5uOl48z0BFJFWRTdFWNQUbtghdwe8ZrPy2GBdnz/SFcGranosf2UL5c11
wPYWBMvvyHGtr7sEw9GXYOvaSONQexv/l7UcHmph0ujHl5x52KChCMZQJoh8ls4ZSvs7VnUu8tuU
KEFYFIQ0iul0Jjwz3w3kTFP651IGgic5KpHkYBksA9fGetgIpY0BBb223gIbhIzvr+xw3VybpaQ0
wS3kPQSe5tD8n1X/Tu7zR79IVDHL7imW4p4WaqrxsLC8PQAq3QU9iC1tVUkhaWZJwOaaYpYTYCbc
ij3RJGwKVkTwffekKL2lYp+MfDzgSrhA0Y9nseQpOJMpgy8oDaUANVLNlzTZ4EOUEPOaVR/M0GgJ
u3XSUIa9JxvQ0S8hMBZgmPu0f6+aB79v8NGPfplWIh/eXw/LGwXB70DprIUcHk5Lle0BdASfoJra
wsjwi8DKLDSrF9ajo/goHaS4OK4Hb4HzevBPH+ySVO7nyshi4SBWApj4z+sslpS0beTTjm2s2ykV
ejo6FHyDpBKATaVhVEFkmekEfaJJZRnFtOoi6bLRg50nynrdjLIX8GRplEP0OTnsHGFoxWxfrpu2
aQ2z8kGY5+CFoL3BrV/IF+3+NjCZFnaCzxBR8LhlPSNVPHW3mJBNjVPgAjhfbNheVh0VPC3fB4rk
k9AGmfW2kvJEItnrxSFM+9w8MQ24VF8xXUeBOzQJq1CWLRnbZUZ2xoY/FKEU5ZM0jmL808UMWFMv
HyJt+tqY/VWoRrsY2dLivozfJZLEwGEwbUnaFmtSm7n4tDyGltkTOAtubqkUxSAWlMxaZXMiWIhO
T1/W44dAKUCLZFW6OsKp9eQfp2DZFYx/7Yb1sMaBfP1vnSpXfJu+nb1pyoLGT8OPbwt+jipoS28v
5eb6I8dE+bdFY/g85fpj870JgjnNx9tZcBOawdfPmJSeJRd6W5vQX26tBqCxhYXTvTgcaoVQtnun
9RCKA5cSrBuutoPz2H6qs+fC/6beseB7nmJRwc98qBcyQIynFChGYCl/mdNSkhLzPoXDo6Y6iBLx
eTVRFNhbwSBHLJj6DCcuGia4DFkKQtqfICPpbFiIg6jS4JLairLc4SHBEv8fWjQFITzX0c+9XfoY
XqRmhvWSmXBaCakbd3DnNAxFA7zrZr/HSidsq1TUcq0xWE6N/LZj1TWGyi7SF1fySglGheGqrxkV
d3FJLoQu+w+d18Brkc0SKDpAhRlsBS+KIsnozoT1WLy/blZHfQqPiX0rpgmjSEUxWiOJypFwIQf+
hj9qQll2WTY/8gN9N0r5gVaoXZHseKPUablu0lqQb/zdZHdy+w9GU0fQha0bPxZTxy6ymPisZCX4
VMMVaRm5WPZ3z3UBeeYl0pARltRBVFRWqYRTLxSat0zOFq3oZyZIJQfKLTKAXreQv4tJvtUL/HFg
0poN674yRjMdU+XmBokYpESC1fPje3QYrr3T7os2aH8XMnt+Zs5Wgw+EUoI6iwO5jlfbilnN2isb
yCihFSc43mdGTgLGY5dZEFIo3YCj2XM8LzmGdCB6e/bftEWuYAE1p9D5YU1vWF7to1Wh8o+c5Kh7
AOqYBYrugrB39D9pai+Tcr5Q7DBeeDJEcJTM98aiqYpR83LzMDgiDYc8Cq7/0/+HRvqUMDTQeAVF
D34pL1pL0c9nZCjRBeeYIJW9Xd+/GNN610GLcBDLgEHYMNH4rmtqzmBMy6lo2v+YTriDjwie1/kh
YfvgosUtzcOQICl38IU5qAk+a5q8fkg/HAQnkwFgX4UgU5fEYkibbP6/lbL/ZMjKWRSGGxf+Owak
0uGJO6gZnAhJS3MwtDAYsLWncTV5gKJRT3Es7Qwt1KsgRVc1EW+1ayximji/eBlej1nIY/3tMcNo
A6dJxrOzDwf2GhClNkt5ZjVYeCgnGamyvD+0Cw/tro1pzqX3+gTxGGow5Lx/psovEFow2TMIJauS
/TE231aA1RRCqKgoYOevrm1alXYAfHer01LUL6itgzefXev+vy2Oa1Y1Cmum6fMA/GN76K93z0zu
udehHZQplFVjBcQbTVk/YMc9GVs8gkHvjvBIk7ClXB5pS++Jhlf8V2lRfll08fQRinaKd4EPjHIB
jV8G6xI4keDQ4QLdO5ZniJ31k5ubdwQtTXit1070QTRxrhjTF+sz1uUVugQPXOrj2de7kmzaWh0R
ZOFqgqVmmQWxXvVH6VkQgNWom5873tF8nYy6o/Yp1BhhrmFc1H3oncbJk+yZ9aHFNBajsnmHTByD
hmAysofiU1DU2I4ncNaUxDYGNI/E61iOJIc0zssF6Pzc3lgrxAvO5X1l0Ax+QNqXIrwrycyrSzNI
CCW/xnRmQ8cXnpFFGpGjW4kXVUreadintEIpDL9kbtCUlLp6GJvM6jolmOGZwJipmoCAX0fEozJJ
z3kbETUHWJz93XZbCoHN70Bn3UgoKanLnou3WNEHKN/yusKicisL1iPw9Ckd6YAZPhGDLlGy/UaV
omU1D8v5s6vnNQnxw92swBCP60dQ2MOdd5NsGfo3rYVGALAZzRovWXkuFH/7wc8eIaT5NZ7+QwWX
HWJK+zahgGKcuPC5DafmGwkDiEfIr0rZC5QRQBli0KO7qyexjWfoqpXoCvrcEWMUlRZjjbd+IlVY
MW60sm5zciLhXTHDZLr7nim62rYSvq3x4t48++Gfybuwr8HZAu3TPXkwkEhKyUxnNXJp29BUqVk1
5OXX9l24DsLynGBm/iA6wq9a6I0HE40greur0UmCi2xMgevPxy4z0cbC0HMbuCXs8ymFP23sv7Xo
8TLRID3RY5qrKcXzH+0TctiinaschsSYjoVOC1ixhV2wgOvgVxfyzuZZOQT0p6v+8q1pgPInSOUK
DJZpkSs5Jnpg9pTBlJyrNTubJboxF1nOJEV5xYwpd15oaqkDu1hwMpFaFtnBLS5pZ/bHawdyA6KP
hxeUBFJx+WL2o716rFy4v3N1kv4HZ5CPSiTFNj+G2XtWQ1wsr4KdtDEMBu16vE181jIec0vB1GRp
4hvY3tl5qY0BuwYNgGKy/K7WpwNyt5KPioGnMFltyb10YuY0Efi10t4IiX+DGwmfC02QMR8d31ey
FA1/v28OrvmYFxGTzCZa1RNml3w4taZDy6s4W6evkp6JZCxarvwi5/msRhPRbI+2TA2lKChZCFBa
fZILNyJdOgwMv52B/FE50OY9fh1Iv/8TDycN1bIH7dJoCU5D6sEUD7C3UtR0YtvwwmAVpoSbMNGG
eOId7mO3y0htBm66Gjq9I7CPg7aQJfuCrGG5r0T+VDF4kKLAbt4mmAfXHTWcZHOmUZukE2i487bu
BzlcPh8joXOxldCClPHch0AQygIr/fnhJO5kmQBWYtHn1aFVLsQjNU5sGW9Zx7o/QvtlhZ2XRw65
4rWvTifkWNwSH/CTbMiyWfYJ7p1lyX/7Ty2WwuAb/42e1PGkMrrJUVVKbDojEQfaBkgz/e/x/wiZ
YCw8tJFnW2K7+QDilg6iZmmcgrHeA8ZepCorrPyo+d+P+mE/h6suyl1jmz/cqncOFMxptMBeSOPn
hXqS/Znyekg64D3eraTYOM3l4Xtgor9EdK8A0T2m9iWZonpEp/487vhTANiS4zCt+2Y/47FAcljy
NckX89R1jEUteBfiHwmTW0NMwGq4y+KcEKWYAYH5htnJFydyzK2QKI8xU6SlGt8LUPANbhJMu7aH
5mr60HLEWmu4Nwzo3g3VCa31kyI+lCicAx77LIiHB2uw6tATFVwzldpSnTm6BqAYotFy/pTIBRJy
q25s9vvaJnOPs/pY+EUqxHtq4nGEKbWHqLlz88SE6LNTysYoiRCBXUl0y21dhxTv8jSRK8N7qQZU
uxvGWjKAzjAfbericdceoieSYb+SOcDjwn8E4SJ0RbaO1/iAvxnupynEEIlBZkF4XLWxuP0AoAxH
1wL0YDd6Ns7Hf/5fllTvOSb79y4Fm3maZchSSLVOvlq6O56EAr19R/+m8ji0foq9FeX39va9T/G5
IPYIrtuNOAcjGqfkerBFTbi1zRbFPIdH3ONeRvcTMMKPZ5CXwOWepzLifrt5Boari9Ed5SsZRxfb
go/DRENWoKfJY1+R/vqWViPY+vGodxNptVeulIRAOOKm4T/sGewNnyUjPW7WnAsxTy0GchVpGkZy
PYNWaHjPdiEQ9oI0+LB/7AdL2RRbjD1SLr/qYvBdZfiMIgw66Vr0shS5sIMLWmQ2AKEPvwYwwRQU
dKqrZgfXTnigiusqEDjtePkkBjrrSmb3DBfqCK1Q5E08vwjwFfTXX06vq6ctFiv9FmilnVJ85Fx2
FlwQx+DAitH0v6tBOREMTw6WMa8jQlpB/ZZlc4BKu26KgtLpNsG0sv17Zua3mRJqA6CIgt9W/pwr
GeqKFaqisu0ZoDVUsChkZhf6NbEWpXOh9s5q/H8DjCe+5fUJl4ywwZiSW3OR/Lm5SdKVY/JsRTPC
U1EjL7CRtbN1ZkE2jMjAKbrNfid2qa0kHCL9nPgw/JFXoybomfNyCq9yC+EPxt33XhIQg2ZCPqch
FwPGXge6gG0o+WZ8zNXZHLDdFTQJndzxcDQQnc9Hrnm9A2DZi6+v57wvu9inWL3aCa2EHAJyqBFC
Qvi/M/HUP5XUIzV/TQsDAEe72zpWEWyPfd78w2JurDdnvUSjlzwgrr1pTK4re4SptjlF6AxDZREG
rFXUWkBrmaL88Bh02AhcFi38V9DoCrjFkwreQGTDmiDAuXfrbCIU0H+RDNhvvHJHMpM+OWvnsH+Z
TA5sFoOo7oJn9jSEibrQfzvOo4uUo94i49S2ZXCBNMle+pfXBSb0WE5d2L/DC57X0vNScX0kyhPc
2OVR4p/xWuijzPV4bZkDKHbTiy1yCz/QyhLkHfGBniQYQ/Bnr7RFW2iykpJM4kDnYuQNWM1e6NwR
zd00Fct43agWoZ/WZyLvlqEJil1UUMYSV8AlrltNUCOVICok54A4BubFAuPvzcnkeAz+wqPoi7M5
XHqm3hnrjKLGYhRH+6Wx9InmU7DFZ/VfryiiewHesphU3cxMW7Q7ENYWUngySNQxWzE3LCOkiq5m
xN7aB+EvylwboFPq9BxqW6zwAp3024Kq64Qv7hzY7fM0R/PDhlKobfLCqcZKkjVri2uZKKjlFlRo
5Vj93jbNNKL5k80YsjUnAn4+9i7ohgwb8oC7jfUMJbfcr2ZEJLB/dtGafWF4EvWmCK9N/MVVFdDa
OnZCoYtUBRpwnvK/3lo3r3/XHnA8Ysf+gp/M2ki0Y4Y+QY+o1w1rNr3HqTMlcPT7745Fe9rK6PN5
iwKbeFlB5+kqG473O7IRYftTbGCY6exlpURDSU5XoWEZZ40X8fzMLVm+vOOB+zCik4WNsbBO9HPw
qTOI3Wn/cdWwDIyGT8To8Guxq3uvO2X9xPxeWM29T9Us2UR4K8mNrMTy4wOdYz/1zyhn3QBbKX+r
Ex7xVaF8J1fe92fAlY+GYSah8ifVgc3pZPhkzV8xSQx/jfvcBL/R/bsQhybG0/PCtb/weOoBy4uu
MziMC3OzxwByYvCjDoiPE207DAQ1pTrwpH+Ydi1OZhA71KKzvc5HnHWMARClwZeH/X0QFfDkOB5p
/ws1zqzxLlDYd0zprAn6ukIH35cHcjMRsSuSGM4u7j9cHB8raEq9dzXL4SU34dfqjeqrPpNGlCfO
hLW+ZfuXEXsO9LTSYJIPbXdNYxiGPxSnDMDp8KbS58xEZvr/ZOLT5bdNdHlq0bkLuXgRxfIUVUve
OCoc1dUPwh4IVT1dlv0JfHRVpWxpVDlVtuBoVCoTTjJ2OEa3g2qEQffNos/R4fdcAVnlFZyx02Di
Q78LjaL+YrbHxZGVOtejBw07/9ePWAEEorWDg3OGSGjsU8rrjd2zkGuIGJ8OcGwvwoq/3UKZKG45
B+5ixUVhsy6i237suanSTDHcxwGQrZtE3HONEG5nNcr+lBg4CQCWK8Mq1ve97soBuvZ1yl9m2hRp
H1cOo1bQz3Qab7XS0ljzj4dPBphlcN4dCONDX+PU9Wpl48SnUt5Syc681sRxzueynOcF5ZH5KAYw
+hWmESDwlvIBeK2EMQ7+CUjwGiW74PDzRWtYUdxvaLsQoB6QJ8HI1wIEoNQ6qc3ouc+Sa/XA1ijI
QjAAANQ6vTUJ+FsSt0bgcqYaJvLVxkEX7PyxrqNPlCIoahMrNxdCdK/3N2vLTE+4jPka0Ok5Yug7
Rhymb72ctZzYEMpvzn7zHzpCy8OZQhhZ1Tj/dOVLkp0HMVbLkYBZ78q/FBV2VvAfxhscsLeiF4Ki
nNHgqEj0cJ+uL+v+iOat7YS4vfUuEEZMj0w9ySwX5FLCiscnZwGN0R8thKSiQx8zAMkBt4tZfj9f
npt+qGGBpnnyO/p/FT8XYZA88vM7psy2WwHU5ST+x7d8+4bnISNfFe1qfruR7RVtKYXuqI4Be4y9
YN5pBXU/j6cWxt34aDaf1z8cSAV355b77YMGR+pyTCRpumxmn5TNgGbeRwkb8HaNRn0QDlU2iObI
8Nqepa7HpPdtr8tmoYSApBvvlRu3km9HSWAoYjS/wCd+cC5iiZnUFIohuApMyYEAfNMS082EfK12
TqmxsXg3JAs/2gdywwLO21rEYp5NblKWvuQp7dFF4a1BUBk6a5kIbP8URIzMefUL0+l1n/COOdzv
W6BBKbWJS7JM+o3PzjQxRLEuWY4g9RiLchiGgwgS2hC6DMgMWdASwGlco6QADf0wnBQ3sgL8MHX7
JS83qjx6AzEIFfRXu5vhq7juTWHRBFb0ewKn1Q4IdnveKYE5+FlfpbM0a5XHuHuGeSuCV0VM2O8K
yAIdwGcl3+wIA378Vw+KS0nTzjk1rPor/FnBCt13XnRh3wpRTknf93IMXWldzcv2rwLH860rHgCa
+8mtE+ThlTmUA5ySQmYwWd0M03suP7U2h5YEaTK3NmEM7yjG+Bje+IvC4DcUz5G7PQAHzZ5mzCbW
+Wu4VESVcDBV4viirC42YrNSbk5Z66XheENwicn8EYWu8k2TaUYFx5ivxOHUQowBjwzTa3G7qqgM
UP/IbPFofpuC9gHUkxiCiMC3HwI2GoWon7Xp5qx9++Rhg6AJoK0pjuQu/lIfB4qt/U59dyTpdrqg
mG2zHDnmgtWOOcjM8gUF4K/R9KY/X18cFPYzry7YvkEaDjmqpkzardARkc/K6/gNqJokCLGC5YTM
X31YNfrKYIqBSbRGWWD/KPuRWWa1yRanCleQsSu+L+RO+zjO1QtrjgXUh2ip7AUsJP+BFICq+NMQ
EcIQAwqnfp+2KAQbuxay3Z8Ap4M0XC3FkM9e8MJgwwxMhDTr4G9d160LnNSnrtRVD9hjFibRxum8
Hat8bsU3Y6anJLXFIW4dYM4Bjd/OLVMLcCRhq53gvej4J6Yb8LINb7jRVVbrF7iibiDb4h7Jclte
Lc9XyeB7ZNkISDG6tEaTbSzQB8mU3ChHdpC6dB95sdnFzijjMxWC7MtO4zgTjHEyt2qI5T0VBDo2
lcyPh/acgA0FmoV+2qEsqrmO6eww5QbqUNC2gBGmvK43uu23PetW2iC8vJJs/7dVYhhHWAqXhVeg
scab2NYguTNCtwsCZ/Q3/PKhk4EAXU13C0mf/mqeEI1zafluRLMryhVCa9U89l/Gp0aEddX5+Xbc
1djatf01cGXMk48dOfwNmkjbm2SDoAbMn78FMutlgGLZhhY44zHc13T9TT0eCFgJ+ZJ6Z3x6JLDj
lTwf29P9T7mRTdtRTZwOdvT+EYNnt9MzVUMrCPyg7FAGeLMjmAfyYasEs1ouNDWX8NQPtfk6hD5m
ECIuJhcXwBp7GHcWG36MByuhbDdVaGUk7W9aTBO3Zr6DiXNhzzkJVnsK8j+biRXadngrmkIrUrvI
Q5UBY2Vpr/BT/bjo676JazFgBROnWz/qhFnanOJlRgh23xfdejGbKYrq4Dh/kARMS08bXRkjjnZQ
fMHLxITY3eWfiABDW2KR5dEz1LId91AWwEgJ0KZXkJLPRcuebM01mGuycUIkDmDDbv0kn39BHUfl
Tp9A8c2jl3KASN8J8UJHHeB5RKkD22/GTLDL0ZkqmYPKzE7rZNZHvZrDY1tjHM2PUA+Eu2rM+saw
ZzOEPOG66/rQ4tLjk+FsjpUgT8FUhf5kG3JCxV5Xz6krp5qPzKSdECAqipDVrNMoYd+9WBR7v3ku
aar0mBcf4rl1vY8Kb7qfPFIYlI7NZ91kEKZMOZ5hQVOLvy3ORSw9snyu0549HfsYIhxbrvPYzlNQ
BRHQ1kUZCySwKzEDepVbqyI4lWv+k1H3M7Aqdx7Teix4f99Mq9Ub5KgBWwMDySRKnmn8trLPIIM+
6gi0qVd+oNJra/hhNaTba7HRwNX4IyAZnJBAuzCAXNsaIgLp1h/byNrEt1WUqatDS1Bxm2JRqw+5
+O/Fbk2fY+IVN5O8wt8xD/RWeGtQDx7QuxmZzHfuCy5rq6n1RqjdFcyOHRpypPZYa0Bk7P2aKz0W
/QBeNrW94GqTWuS0A8jhSVO710tutl6fJoyyJKXNEPNrHbcZOkLXelOP6H6GimVuhhiTn7Ete3EP
1x6OJ1sDoNfGp0s9+h+CtL7GvSWTSaGhgbaUggiOZy9Pr3HQLSg1Ndnu5JpWKUFYCZKd3FRdoTv6
Uaq0o2Y88PUzFa9So2aXD0usQr1suqdNNDKb5lBBNTsTw0iuFjitH6aSMtm5xGAPw2kGO6FHmZH4
2msgMI6Gtv7kwS6bw0bEl13h1ySNA/rd3fv8vRxmjaBFTCDP+2DuJQ/0z4MxbsHdkInDS6pGLahB
SwrfP05lnAKd3AB7cRgy9VSEL6spJ00szwrSZZKwd3Dbjs9FyN26Zuu/OrTjsWpwNX5GFeBE3nOF
HKy7eig/VKiVXgGlrOicCCV3KZ34Q3HieYYSceRGOPv/3rVXiNtledY5ZINjS8MKbanzqMsiFHYU
xN+mNZd0bCQOmotU97x+VP2QkNtxtqPgnSre6ZYzcOGx3X83ImNQY25WVzWtVoASFwzZzMthLgXl
PwhFxZlibqNYCKDvpbkXNEuJbGYc3yh6MIfEvN1JzfDtPpJJFHmH5Z1tNfhQucpfQSkKQSnKHV17
1JSyyhlvxk2qjGsaMQ6Ls6MOO/zbQBXdZTDYmuOIHH1Uq2BcclNwPjrBf62CUD6EVgplUxEh5fWy
9Sw8k8eCN01Dsdp7Fk4hC/2zTAASR9kkJ3h26UHpw+Zq4sIC0MxykgecCvOG2als2DqV5AOJH5F0
FIcps3tnn5T3iG6VkBVUiQJUw+NvIHneRoQgXAv+XLmkxeDceH/SkEKw0ouSfMCQCv7o4ZQUb2KJ
U7QRKkUYNjisD/Am3vNCJADbzTKI+hTwtq2Vz35ra43UBHR4np6elCvycoD1p1hdUuxeHQCDyong
bBxKJWgHhKK/necKL/nLoC2V0LYXGNVYg7iGNAuo3VTOSRw66DB9O26VFcveVVxc7jcoQ0wIcE5z
HyVBL7sFwFUNvebmvi6MuZNKA7FJsBN9nqUHsxWMBE4FH750pO0/cDwWmEQMYOvUrnobM1lq8why
wrubehXXRTjLc+GIPMppL6Fycp2bui7ij4BSdIpOlXjSpkRI2Ppieiid2oAu2UbV8zFgKMQiFww3
zwvdxdAHRlfdftJ/cbJtFVJbgIco4QrG0jUEGNqPMqtyOXIa+m1JT2A8ZlMhgKQRsISjeoot1Qyf
gF2rb+sXzLTUU5N5kMTVAf54xajGj1HL4M0Ri554GUsBkxJhCJMGbhrFKkLl3op9BdSELN2R6QXf
nRldVJi5bjTPrLvKzGY1uVjrj86XoXQAdrYA7qEDC88z/nK1oIRoxxGgJSIQelUQ2TTTKd7mEU4F
jVsewIppzp/RFh1n/m/csg+hM4tPYapkd2HRsyaCAp/0UqXHZ2weMReBd84U1Ds5jq45CtFoFYjq
DG/SbNmY8lI4Ej/iKFMUpUWfaYpJ6sxtlP7Qz1liEYlUgTR8bccRzDPyVf5vtuRMEqzCszGz5fdE
G9UMyN4NFw1PuxR+ZUWCmAPrWlhU1VjN2FsrtArpt4+fc/kMLfi4rRCH8ypouKgeQCi+mH3kNzFV
m9q79ZChZa0RKNtjq/O3HF0MHjX+CbcsgAINuLW8+iz9kHkmjwveraj3XwNCSSdpbQPABI7f8b/J
qNqWJq1dBDKnfOKrXFvC1jGpur6AT9p1dgJOZ33mYu5VyvYsL/LQsSkGFKCemm7Cc/j97f5erz47
oK0Pk1NrMEqi0yMU9R1KPRyhXEGOUmqFBoCCgBRkuVkGvrR1Ikwg1Ol6Cq0X9K48Tb99Z81uriiY
hjWaLbisxCNKbSMwtU1L6gld0cMi/hnIgL1IP+l6su0OIP+tIaWq6ZI5zFYUZD/rupGhs/8+EEnh
FSU+ZsVvFXhMz5Pk1SNSDixlcd684s2oOt1sywXzI6QedZgpngVuRdt7s3kPkjvrbxey6WPI6N1V
cpQA84ffXIK9h/z6JyEw3MvezPnsT/gvFvruknEMG5DFFaYhyxhctQsl39Uyx0nMcgpoJkpZyBfI
HhITBbDFboEfzkukfchO6CXoPwYUAChvZu4CIHqCc9iUEW6VlsnBARJ++QjIulrgF416V30MiNIQ
s21O6D72XZ5jR4Dr8dN1oyLqxvMf0UN/n7YUsf/o2VGf7xWFKZdxWy9LtMkDGNYouyT6COfCK+tf
9/VvnR657+m3g6qwl2TfFTafsu1ZEEs57WtQACxrS7Vde0pTZYNdspSepg1Ok5XPQohjdoWIkkNC
QerS/iV8QAD6GpDuDWXsmJwqD/uTquOwuGTma8PM3F5sAqxYG9Op9k8N27DCxFflFZOGR/opJHXM
dkOXShtM8/lT9wAJK3BPy8v16RhEUlWyNR1qG2bgzVhC+MuviUhryVM6nD8gOOUWD5Xk8+QsKPdK
LQS/Cy+0LjlTTEtloXvXA2Wcb7JMCMOMuIHPYbB4YPGH9RNTcEjLFjadAt+NEp2GV8hxt5wSAvrg
WUKvYxdLmyTfFja/x0qE0jAmFnJeMDgu0yGa7/TkWaGBXs7HmdlqZJxHggpDNMQBc6oP/ZNliEbt
6JQQhjiCfetmu1qAf0a2636dkYnRUx2sQ4apLcg5EnxALtAzkyeWSWzklLFfZHoSLnzRjsSodduE
BiNIe+yGqrkWTxaC/sdzXMVSElR2qZXNCRFmEJ25lCxf6yKQvOl92VzR6goWMc2YrD+1zOYKnC/d
sEY1YnwrZpT/fHIzvc2GFH8WEisvRVW1RAEFxKDU6MfPBdPS++belo41fCyxk5+ctDF9oP8wh/AI
cSlQpckCrLtlZ4r6+0ZUxzi79ApPrJG1t+0VuIdbvhk80tbmqm9ISds8IRisb9QdV5kFwu2/nTrh
VbI49FxDY5kF/66CwPtSPKuiwiLvsdJec6ad6A9ZiR6spOzvn6/O7urrOrGyLopP3wNTxB9/uKkQ
GBZnANNx57oicZJ7ArsOvnv1JwdY9+bR3e2TkEMfr1cXdWXwk2W8bDYQYDQIMEMep3uDw6B9HM/V
wQdAhiRgQcQDqjahfoj9hjhBA2dIwEUBker27cohJ3qhRaOdQKEVFS1xvYAqSho9JjFF8xkK38IE
GG9mE05NWtNxfIyf5tTNPOpKM+wB7ejfJtIxVqmdqkOW/k+Bn4cBfrkbODhtCZvmwy2BzNXwsjSV
iZUhl4OFu372dM4co/41fK0RJ85gKKdQbMmnHnQeJMngJr14ZhpGYwIKp05J+AM9Huyyotb9JyK8
iL8+ftHFq2mdt/sb2Od774ZXxgXjnkUzmbABUfb923o7s+oZastUf1ja+cnxa8MQiF7UMDh7y8V9
2ThyZ3EDvDMUWCQTPDFfFsp4uKL6hPNSEYJhM5eAm7tUhxuZ/quIE2Etzb/yyKsTuvo6NmILs2HR
qWDZYd4nisj9XBvXEORDOENuMOy6PRvK9LhdNSEYTlPXMKBSZjGu28BzFTcuNo4vWkXJjJ+6gYuB
qL8XVpeFb3BME78o2gzSsPab1z5eTp8QN/ltkdcEPgs3iMjbNMgijWhrnPpgU4cbgNTrH4T/fjB8
9DWHZ49WlLELNPLNF95556zo52x1hc7IuuriLPZP920YlvFOvQTWUSYfrHCpD8TryM9JMqdaVwax
Px0XGUtZrfDq/3HGV+l3fl7Za1odnvbJ0BeP8/VncmAWRT+h9mwbE7+gsJEzKGqYTXjU0ueBkmGs
5YTu/6HINRDIDy9eghCxYwuBQViAj/l7iOzvC5OkAdtZ+pAZVwaV4RUUa6wOCEM/H2iZ2GyDa46+
3NgOUegTEnPk0TuVRFZg4gQESyuP/j/ZyvkoTcAoNRxkz689FhvC6z8IUHRQLKaAOAsgU+8tDaXk
gCSkthZjIMqjpxEQFLoDw1TktilqjLEFZz+JUC/z7g5Rqh3plfaGp8UBy46+XyjRCbQNypxrrj5h
yTVAiA/RnjLYiZSWvdpAnOIV1KTFgIK4uaO3hpTjKM3h6sO5KeiDo1TUydGeBX9uOuF//CvFqp8g
8/tGlkMX2Qr0p91cWqC1qDWxdKqR8qcB3PLlMNq05D2IoJI/g+WY6EpABt7VWCDhwK0eiZdqlAqy
/V7ty2D85mw7AggZtW3ZGORPsckrVWPggl5QaFMLBocXjZNczCRf7jQZ7UyPFQojofiFp8KUYYsB
Cwt/kSGCVT7RWgv9oKLOWnKT8mhsPx6L/pe+VSFNEL6gsUJmqVjYjuaVLOa8bjB/DTuD+9t5xhAa
AlDTAldEw9UKOOIv4LIVhxQLYiuj9TVp03D0ef7TzsrX2oZc0bb1MTJq94QGh5Yhxbodlb0zSnEV
0BdEsvd4SuHu8VdbCvOgtMKq+nBPD+rnkrqKdTc5alX91APKmOT2S5nfXAJ9Lb5+xu1Z5DPPufoA
DDQpn8kfzgpogtL109m6o9pBs/ieDKht4xwNpDvWxdR507dYMlzPhIce2/u+ONAVnzMHizwU5awU
amKIXevUQYZtUzhJOh3vUEZs6MmpC1f9B/ekzuc/oovJ1V0xhvFZdZhSNurYlWZORopWLwl3WEYm
Bo3xfZcVs5OsmHd37DVlSZK3TCaSXdHxa83zkIENzvA9YMjrgorW3ZOnaiAPC9tvjDgDZBQDdZ7j
hk2AaA1DqBx0WtSs9uzMCGsE9Qcz5b4I3DSFRNIcSadxcPFc33fOR13V8A8b6rX+OPgn36t9RdFI
yao1nxxipv10rMFdNnt2oohXw0outW6Sn2A8Jrm4AkX5hA+/2/NF7UXb7gz5Q5+vN/mLWF8IQkAf
KD/IFCUr8ubJewPiy8yaw1JDKtv2LlfAV2JmmMz/6PMUyd2H+HEt/ps/PknoEe7dpx3hC5CHJ/+Z
0upKdbrpMgor0PqE0sHCz542cSHL5AbrN0G8gdA4fIXUGn/7XtM/F8udW0ylUOyDlEwVCooCW4Q8
/VDERkyypBRVfYfKrHg59VT90h+6pa6koGnzo8z00s0stcjtvhSuNJvzbMM5F3u3GSEpyJn7RmpR
ms1f67LfQ9fsYjrlGD0OiIaKryxwgFrn+9IQEpbUkO6Q/DoyxQKNXB8OrftTbxG6gp+zI4SB8iiX
+eTVxVPyFI0OhW+k9Ig4s6M/w7PkAjKPR9wBXmYr5CBwjpJcH/j/iubXZeHlDchDJNIUkMVMYoiQ
2OV+3Qn4F2QZewQc+oQdG5UdQcfq1qBuligHBhFUg+u6miOPaYjpTx5w+uKoY+MxzrnaR5/rdSJX
Wzdqj6rrN5TBd2Z+jwdpAmk4G2/98be4ArYncunTTqTG9lpDsddDNySLSpC2M26wiVV1rCgyCJZv
i9mAneTSSDaN/LMHVpIEoYK9C5nPpj7484YeNBoYLizdPsr70cDRJkE3fAcfyKBEcgVxafAgGgLc
61VCqJznRDKFSxtijk5ZVB+nJPueTlUhCaEG7Zvy54eb1zq6RlR7BU7jTl7j27wntkgvNgoEV4xC
ZFZJ0vU79fUUWG/cKD39zdbYUVPrbvEpI0xtB/GEbJYeidSSak/dA5MpFJ24ZN9cVgVxRRFHYd7+
DKgEhwESeXwsCKPlgm7eKnZTEW8W0mVJ2ouewaLpqJsUNx0mtmCsIHfvQJ5TxzA2XsV1x3cIWksp
NRVfqdK+j7iQAH3f31pqfv3fDCnOfCf/lR3sZHDvE+11/uFQYDFseUK2MPAb0olsPvHV2tsvvSij
O0SP0WqwvI5rtJ/NZof/X+Ld82Ll5mSg81lW6UW0M5oIOcSiL5+RvBHE14i1Hi/gOMx/q9xOaJDn
LpGPbzeKdl/Lxr3CaZHZ70glEwU2OICx7cZJo7lyvllSNHij3c1RZWp2s6aA3jMyvGKf8jlpCt4a
xS8iaVNU0km7et1ksQ913wp+seBt+X7Okq58JiYl6/dlZHFv2qExwpLFFY0MlCEV9F/UcjmktcFA
6AITdretJojwR5JWpCZmZPfFSI+vkO+jWD67q4u4+BYwToCCaJYxSvEBAS2337tQCsbR0+LzwfWg
UDedCdwo7xwJ8EbYdZOn9tW1XZrnWj5nIEg+Uwnlr3eUBQmWvdV25X7zOLxvqurm8rPuZbfCPs+/
BCnkM8cvfepHtTFCHM4/y1/YvmRF4TOCX0zd2+JCK9s79gUCfr1YnCchkVpszsTXYtSDrOOGKmhh
e6dwP9MH6gz4NBe9pMFHl6LBxVXbQgYWcxn7osKlaQvD9w+GoZ7Jp93EYpkTAnm8Y0gn6HEQUT3m
A/X4c/6qzjOs1IwbTPPFRbX+Ew48gaU8K7P65sjw91sSAh3cuFIpZcodzowtlFAD8090aAzY4tgg
V96zwwklX/8rMg0ykJPZgn+9jXfIHY3cmrvxcVOW5ZIq/xEITGK2cTlI3DjwAJDp5uAXQYfQ5ter
CdOdDF3l/GjFVXsjbhlL2apT1Ok4W3s6IaRJ/42R3yTnEHMKVq2fDGpqdn16w1vRt5IPqeFQvPzF
mIbSgRIvjIFwd8m3LsiGa1f4ACrqg9Qw5AXEWmZobzWeWr/iUrVidFuREY1fQoU90gnFd+NtDjz0
SublZ4OxWPCe9MjBwfetQinHwAL2cXvpldIdqt+TwGayoLMEwG3QwKlKaLdC9yWQFTMda4BNgTvg
9GQRYZWnSJTLk27JVFqG7UCpYBgo2A2O3uPFW7FW3Ck+OG8SGPjlcUKUeqDk1TlG/YnCLYJDnalc
ZirO64EuOq+mUKLNEfW8gH+14D0NAvhMZqrMLFkUB2tXk2YxSwczimxI53oHZNil2k0YMqUIes4R
kR0hXKU512yF1EZggwPIXJQFcolcoPep/o3QepkGOuMG9gnxo0BavrfLpgBw7KWr86KigBz6zRp4
+O9NkgGAgcD7f/9qBomI5WA8gAN6de3HeB2f1bJ6rqP9wLkGSbWSTd0kh6/58pjrSXU4h9/0YXFE
t+Ad9xOrPQdfG2mCtnkXI5t62Ge4KS1gptYz5VFpWNbLHr+98DcR9XCkuyBic2PTYmWupvl1xuK0
eIzRHf08ZG618usjVv8ab6ewADdQ5P+tZM7qMzinZ78Q6TwgFY7SEumNfDzaSMygsl2lDDGQ5XSN
xhd7AgwHgIXyrtpjdBU8rWgt3hhlRg17HAmxh3OXe0yQNu8w1KsdAC52FWsVC09jCbnvMWNyu/05
wxTsppULjpwzKcBQf8an9tRJ/AvW2bg5XbqJs6k5J4qgVXphOWkh5KEdIqtIDihAHiICtGfN9YdM
yJf4G1n/0Prc7lZH7Dng7JIgcVk20kJW4ziC3d2QVz+A2LgM4KCSg/KioI+/cuIfVkfs2QVycNW5
0IWBxVyVolqW5h+uapdoQoYTcym3kKOrbG2zGR1nhjUfVeAbPRfdVDLQ/ifT7968NO1Bvw+RvQ5z
1pmJ1nH290Dn85JkBb4q6COxOoMBgNgSk/tQQpO8XRXGxI5HoP763IyDYEP2KYwQBnhFAp8a5T5R
BCv6K/CtcJuRFFRBUWp8AgBy+F+NBH9s0T6wkBzbyiYeCImRhGHFsNtUFVRgpW7cIUWW4+CYyvpq
dfjjqzcOCubm5NhN8YzFpKm8P+6UuNw7dQWzZrDvGdDF/Dqj8ge2AdbnUHhWuY+snVMyJA5SSWeW
tR/vnN/ApWF6qxTLcDkyW3pli93fSiRbwF52mA7t1vWJ7yCcUvsgn7aBWaYDb9FdZ7Nu9NpqamFE
cuYdKab7bBeWVWw9UsJwoqrSgYOXORxeB4oeIbT3B1pf9TmCg2HyD8vv/vuGBrb2HWZPwBy0R2++
IjGgXlSwEKe7KTaAJhZPcrqbguziAVIznLqBuPVSCsPl1JlfIzH5AqXxQ73RgOZCkdMHqjhJelGS
ke4jjahDa/C52pgSbbdz0GOqp7PkFsi51bk3wSz8WqTpzIthxcpx2CeM/4L18md2Cpl+sYjgPCvF
CI7kMH6+xIaviUw2VLcppL7dTKDBTqhObG4479DPP8+fKyyyRf5NgsdQolOosURJNwHqCjT5W/gM
G1eJHWKOacjUu/slY4UCNw/hggw3AoW4zRgpMIKbnodUYZiWe2OXXN+nEJ8w3uYJomuu/URoliKf
HlcYSbJarmKSfqAuapOTcD8g/4ErNGHDcuDr916iCJBnES795VW9KgT+BYVIPB8j2Qo0s3L/klTs
EcpXWf2hln0nHBh36ipNK7VuKiq4uOMGjZ0RyzkxUyAsqUtJ+6MnRcDRbA7xFzhzf35Fsg+Tqb8R
Iuk4fZs1Fc+f91JVrtDHG84VRmCHfGrhCzGaKkxSJHgj4ooxfAAoGZPNy+bUy609PinUQGRcihEM
tTruTtd9Kewso5YhrXgqB9UZ+cztJo1WUBhjd20Ny82R2+E6xW/uDuyZF+YnEWpVsm6cumozZPnz
lvPz6NcTRFmI4DmsqdRILk7glkrob6bAxhmjCWV2Vj/A/7cB9z4EY/O9jCbYXO4z1ijs2dJl7wWX
+DGvG7b+ajC+4HzNezdnzTK7GD6zr9C0tDbWYpS+tfLxXweEEPy9uH3My6JcllMJ8jYfd9qQX9Pq
3CAMBiBjDpKRbv6Ixpr7oRSI4SPouBlG92CL7gkJwmnrYTngaNhtTFYwxdjwpObgiqpHXU/r6G92
AUmeBC1MWmT+/abLpPFTOhT9L4Opk2Dm+FwRzZhR5P0LMRsRXr947b+1p94ymgDKyIaa7aVSWAbx
3T22hho8B3fb6umu4Ztqo5WPHl3bvstmvRwHLzB0MKZ7v9Q2RFNPy6snlE/NiU5MptVF8nNQGVsQ
vQu7xc4LWt0nl2NEKrhy3kvSIPLxrlgWmzsJ57jEt9Aa8bULQHTfrCTFni05uWO2dLVcTA4hlLf/
TYtALIQuNgBR6PVjzhwQD8dx3e86Gg/CpfYyZOhGobvUIrq0bdnYmKvk/fVPxWM+DoxjScaWL1Pa
r3/7phdbQ7aUiXpgFD1/KW2IqmlT0fcMyKIiou9eRm/0VF/8doqgalLp5+Jez7fCG6JnfU8QkHBk
F9Y9AyLak2wYcRc2Mw4a3aydWKPgBG6eX21zDVbla1sAaMsKdkNOCdUuB+na6ZvD6HaKsiabicAe
AgjXWSKJ2olBozEJH2GHgKiZaoVFaS9ZuMmkzvCk3QlmQpwJKSVuBXqbGe2fzkpdG8jT9LcPhEY8
TP8kJxR05GN/izuUx1+UL7JkiLSiJO2VMbppchkcUUir3lEiLUnmSRjATIIZFiHQzPv6hP74x17w
iinj9mmYnjwmSAMaGOeEC2oQgFbENghNxVcPkerZsgsDKpZnCjbJPWMFYqVIHRL8dGNJIrBmawGg
F6Fmk8hEslrU8i6IIR96j0EXpY1SmBhR/boDXgl3tt9Atv8lw5tkXz+6eU/1oD751fMvQ/i+yuh2
ODxtFl+0M5gBDsJEUfh60jrW3aUZYBHAo5ju8z5CkA7GEjMlS6xS2/Tjxqg8tI5hlIIGU2VrlOYL
dNO6GtjInBOEGKJuSvVdD0doCU7Fmoqm/iVc3Y+JvUAlqn4F3WVkU9kOuKIEvvWILhUKwYL9tVMu
mMsFh7C1VuNoGDMBppVTidI2VXLy4Voe2298t49A8leGdc/WcJf4/h5khGDjEs3arGbh81mZQj3R
dJoRKQJM+KVUyYrfGf8GgUFmoXUnutYYBcVjiiQnp3gmr9Xp8amTRoW79+OeB8QLMX7hW44bYMKU
KqXL8iPMfuen60Vhkf8ymieWDCgG3KMFksU1vyTuXQJO8TylSgeldtCvTFxSQ+hV77E95fOBmk7r
zrO9SSm7Ih6C7hEAdkLG5F0sg1+kdQLGhqFxjZHTDYtJ35Sn6OoOBhgcR/3jv0x5We9OEnUkyRXA
KlBylcjh2MWW0KF19JaRFUlquM2abvWls0LXLXyUhEPSfS/mZtyv3+XMmqmtMX+pipLZEqp1QwWO
YQPgWp5ze395oPcf4rT+tAU9qRdffx3UuauXtlefmPBghcbDoY7/zTQGHHIVF05e/Rsh7IA85HBI
NHX5gAoC+BEfMj8d72+mlZ4b5l8JhB0obw4cR17J/aLKLNRshkZ2qM4umMaaMY/YpeknqXptB+3Z
0pdjuKgOP9N6KA9qdd9u9xBwMbB4fZiJLuYgYy7wvkVSWaMvbamWrFjCeaivL4aspVnAhutTNocY
tXeidbSVQJDj4gD0IOgb27d8WBNyJSsRA1Kc8PGHBQpEXDsZM4XjObJNMyI1F2ko/q5r5QtuwZ3x
JeycCdivDGT/vrDjbQ7YJE/XGANVpNBAnQFK7T5AoVLDpQeOX+58pDYgH8A4GqTW3VGliwS0st1i
Qn1b31DoXDENwyfOdEe28gBQ2A024xIeXO74sJ58oKK8lStGdtf2N2wdDhaXUJJ2Wd3AjG9/frX3
1pAgV9oUFQHlEiF4jFAyI5PaPem/YlIjFJTC9P25syii19NWBMzP9PRAbfIqU/ysfca70Lk0DhIh
Go7tTBbaitmrBXljq0nL43GVXqcS3LnOBBS4K2g9/MR025tsPa/F5Wtb8Ri4vNUzQHUn32DrJRRB
L1gj0S3RXkRhK0YtLpOk6nS9Zi6nha7BZ8mTLIUjUJwXLP65jfv6q5N+BDkGcWLhKSCsStBnEvk5
vgiO4G464UKdwcSnqPBDxJgQXyF0aqcruZix/SNq4pCJfHeAciNjKbi5rU3wwdADSMdv1MfXiT83
xsQS6ISTLDoa+6RU+DTeb19qwHqgwph1utdAgPlfUFywLmEw4dfxwv3lyhRqlj8kSs3mMJ3XaevS
nZGYbJWlAiFfybW5cTXyajGi3daEktnKGvnb3HVUu7NE3F0Ynv4mdd8WvX6fFwrpBdgtCWpXLo7F
LuAPIQfa5YKISgP3lb7GHqlEgQq6X8NwsMNefNrNFH55/f0pr/5Lxc+VlgBbyPQSbOJn7A25b3XW
2txbFWiXR7q9JSWuU6Cup/ImFiAw/Ol63NZLr17k1Dew20OnyCrS6/5byqrkohxmPWxFFZFxdQBZ
26hWW4hyQJ8Of9UJlwk3Ed2qCN1j/XWwsELG8A2tBIZz9pvVsRKINnrTUf9Fzy1Ns5SX1ZYFz5U3
5li4cuaB7R5UYL3pXuA7K4qU54D/ZaX5MO4oYhKir+QRb8zHNWnisWhLvjrEqpOUpPTNEA4Nm4eR
hEs+yXeC5van1WSY+e0VJs4D4OJod7kuVcGry5GXNXxt7VQmFLyD3Amc86TgAG3CvaLyV0UUoWKT
P6ZgFC2RD0ZPJgRNyzmQqt54fJNA84gGrDa9xJAR0wNLdban5/tfsUj96TXy5piAhLCLIJyNXx17
U6qpMOYFySAFowKxl5hwycWLafcrThrg9Rqh5XF1StLe3gvUL407cunWRi9TrDZgCLBPG0gj/lO6
02ck9a/0Rp1nBxtidiIa/fVOi/mLfY67wZOUWXs2MqrzCdOVCiqsUp6fIyJJ1UfGJWp8+jPyul6I
X3w5Rs4KrN9XqdeYR/uLvU/s0XYdkDUMFyTxTywcJYk1xxEd1Jz68SwaAfHfzS18iA7DQV4a0kHz
jopwZaZllBYVO+ZxaL69cE7ab7AlYx2GTHG97XRijUFRtEw1REeEXLsWR3fg7E6pvsAqxKFIwbdn
e8TOPWv6A1dLa1G+UV0bIzcjOT2do8rBXjwKPkrs6QGRvyD+Jvr08OcMcIkri4Aj5ersx9cgj8Ef
/4FCBKYdM3nvyuHZtDzJYgBFlVwyU2KSnkXxZhrDMED/z8V+67JJJnboz9N66CFNJ9O3cnP9NzHw
0UoJJQx1RMUs68Ug1I9KEkV4XfCt0d4Ws2TmCtLwKTfk4nsWVNTDWViIG/IEwQtP43PiCOjHyxsb
mjKgMJOFjoX7u0jHnhbnkCM2RpZT/qh4TG4jyCtVGxDKNrBPHF91ekydtJYwRkMT/PCc3G193d5L
Us+muKzLlZmxXL6X5f6ix0ELKoHK3L3kvpXtjNXBfgarkQ2euNS318rOojSFoa9KKHhWK7ed6Njh
u5Cy+mSKUM8PL0jszf6j07qk32efVLMQwITanVKC6IJKPTzIwUoprQC3bew/n6ce48/nytQpdZGt
W8BIQ45VPzRMzg6lkuc7YtGeIJ65y7recdk2pRgQAJ6KRGWxaBYpj8ipH1qRDIVOkCYhqmQ23exn
mNY/6ipOoE0UbjGAltnaVTrj2KOplaYUnInbeKnGH0RpZ89XSbp79Fh+zjeKrAyUkEcg8LyTXUaB
VJrFWFD1eZmzap3/LYt5CiDwtG883h/aM2+ypMdmioGNra1HalSecTj/yeaC/1MZiVV8BhHD4Go5
iWy4rPdE/LuDPxEbc3PFMmDmi0yOwnsdCrPmn5Z+mb12tO2S0F5GlttyvojnE18ygiX4Vb71q9mw
QNrn9yn7GiEynQbBfNg7WWk56g/uHLhttIKTfclo8JWnqpQtOvt9g0PKq5SKjSdsNhFxMYdnl+Rt
xrjH56Drd/0iMavNxajjZ2G+PLTlFTe6OccKUx74L1KTPq4otz9AkG+LiUlXY9+ql9bti78Y8TZ6
vfxQtYuDOTBOvA7BHN+N1oxDQy/IilUL5vTS+IIgUAevo4+FSvN9+uKdyYZUogLB1Rs3SsX00Tc+
+5s5lL6KUF7unyXqedXIiG2qDC9VdWANf3o/NNDxFCcNJjkFYqrXzRV6yjyv5R22YaL2gTlhfCkl
vJop/KJFKP5cvORjvbalvs3PK9wdo6/mknbkxxqwrRqBoHIm/wtTzeOQ8kfful8h1GA/9PTK3mVp
el7uY5arLKmLGuMwOGuEyNNgcG78LmsZrYHWSUlcsAWoNgkk54xfmjpfvOGpI6E6nsRnZCGEwFWo
rJa5fVWGHt7VyD+/M7NWJn/8A3RBFYe/9eHwRSTFHJrcxY9E5zS8yoHc8j3Y9cAv2+e11Rq7T8J0
HiUyODegq1ByMsDAJHOodIn3ff7/O3Dtm/O6cD6EVqaBCrgoBjUP8owr3F/BsY6pvhwQ2g8FLDpE
XohQJ7FwiIIpwUuV/is5AW+Esl15H8qJJ2XlSdSBzHXL/GqafwG8K8AdmnVUHHMupcHdOmo0dLEg
/aEhFEKth8L+3W14MXV/R6gy4b8/iW6dYMxdpYKTzF4h8CasIcgCj9TEqDxYEGuxA2fKJEXXL++A
69Cj2mzou5jIe7jVrkwcTxkt3OHeqJSwrru1P451yIMrL+SS5e2V79Pc1He/Q1ru1KzGbSXUK8FM
+c+YD2d5jjGSC6HK2k54DrX+bz6nwaaG8iSa/wGEU/6FmmeV6pL62fUOMkswlUwc0hldvIe+Zxl7
z/84MDAISTuKoMZfI3x0Sr3la6H1Gz2H9maY/mEL6VQaP/pZMLvnv3lcR7IWQt+da9NVig/Lv+cl
MMCpNxTBjMbTsctUY0XhclhGmu8L+hAywKvDe2KtZY+3OKoL9cnRzsTAP602bVVV4voLObC67eHO
nfz7DAJak9vwW0c3HPoCvSWY7oVGP6hg2VIlokcc7I9hjYKjkpbxNPjPLM6rmvZvo9PqtBXNbeT+
Smw6+c5GbL8ELKpGzUvstn6h6RDWE9aQYr+8NrF1vYv9t600mTnbdLrP1k/hGx4eQb1Q6PV7ABKv
ojIkivb8z71gUsdEDpL21aHs8KCaCbwxMW6nvWGHsk7qojA84G409MeItDb3k1E804bsFX4oPo6y
haflshdHbt30unp7Wr5+XsHEYM/Fa2bqFYuto2avEfLVjHG/0Pnyezam4Lohd8YqxgdQXJEWPF6f
Sh9WIQFAMSIYcx86/vWb0DexS4w53Ao4RlKZBDPBJrw8eWlhmyVu+tReWLXAwf5BlMXpt9IhFVtP
INUWs7ZwEAVVZCEHtpVlOc/cUYCNWqYKOeauJLdhQ+SdmikiQQR3gDbEMVIbj4mMg1qsYAJK07fl
0Z/8C8YDvpcKg4H+tW/9Tq8pJTq4JP4Nt2ifdGEDIYVOO6eRiIVZvly/7oPbwhrkTIVN++X2COP8
6o3hDQQY9cxlhDerfFX9qxsFQUMa6NiF2Xs6fRu9BCDqetQSEuEuG6ZJVkjhLWb++NS99C2PiMBh
7ckXY66Xv5lWe+lKvdCnnTlMXIBdn89wrDZxOU6sMXeJVgoIKWZv4VeC5hUXnU/LaBiHtscpm1es
wqQS5hDcPKh9FLmMqzrBhZmaBwKDzJXcMSLwHcz6zElV/EgUqJpyoRU0gb/8LXX2cctZQP+AQHNH
u4bE8srN2pj62u4bTDvqw1HObHHlIei896ItJMJCdgTsFpM7ns2ZgeePsY1sXEdAMpkngJyVsvBB
ResuCoVN73/WChla3+E7ZVWlPhuyzUi5C03SpIvGYH3sCcDPy5Q0Bd6vbvAzEPveR1g7Y9GJxiLD
UcnkEvKpPMj+uLBISZ1JFB8CUJ9J00WWxG+drA5KBvlTmnb09FDjVN3w6zY/f06Z6GhtEStY2s02
gM2ly9TKNa9S7Ceb2Q5QtXAT5PXGNPhOLyToCVIqAEuZAP28iVcTrBdoO8PXRTpXzgxxkmlH637i
hyyRn5J1ACck+GbeaZTA3ygV2xm4LRrIMioDxQQm8xAIsMH4Yg3UE64U+6fOyXogZxsyr+HCEwSu
B8TUdlTWaw7PrWZJrkRgEN66BzyTaK9ShiUZKZph57vfWNNbWF1Ze/rK5NU/K4XLLJi9cCJnSS4e
tGcOGDSMp4bl/VcxjBY0tmZ7sIYkcErHyMjNN8PGr234gy+VimjB+Xar1hHISvGKV0rjOcAkYyci
Jo/tM0Xs682iBLYsl+l4SfWqB780odiulh+WvQxskR8oRswsM7IXSUP6H0yuxnpuSc5+jMX65/oT
QWFuC4nf9zSkjIioLJ5D2fDGef6uzN1tyhHT67Nbq3bYVwR5noMas82qjsukG6xtSMCIwMslnPcZ
rR17mbktKBbs4TDGwaZZsEJ5WaABDwNQThxzzAj7AH/iHMGFp22GRG0nWXyDjEPaKGIOyyjsl4LI
CpzJbr6H9mVn3acC43Qz7sF1Yoc0ro+4E3RxPp3Hve/sWlBSvVDGt2tmP+8Rh7DYmmkOX9GDeZqR
ZNrYkiose9H4H+1DeEhiozllMDPgsjWLKA7LCTh1ME13rn5G00OhcVuQEdEyIVcB6QO35YaAb5i8
nNb396Hny51McrKakviKsp1CMJo3FZzwDTAqPudzvE6wBxXG8VGZp0xn1+ErQo/zS7UQnvAMq5S+
QVzPFYO4ftEx2ZOXwrtzjJ/t1XU/hvdO7QDNNVricc0+cdhlsbdn87yul2zt1njHyWV4VKIYm23f
dRA7bhjFAIw1QbiFrWtr5XGVaiGc8f/C2godbYd8yo8t8cktSXXsswVJFyrL4t8hQmXZW6X8UvRz
mGN3G4pI3nwa87kcY+tsuOAOIzdD/wzgRZ8jbmGBF0e8/+7rrk/hM5xYF2+fjwS8WByutv/DDGyE
6JKxREu/HZjHSvY2RGprvjVoHg6/GObDn5odzIrGEyNkF1kpnxPTaUcCfqwKwMZ7h2rZb4xAsQep
UT/zJLhGrTApZ8nct+1binYFpyJO3zs0mpCFMtc8Rccvz7lw0Lv3GKoN12NfXNKz5UeUkf5ayNCP
omqipIhcNwKb9mJD144OO0YaO/Ikh3GMuh5bC/OVLfkLkew7TJh+dxMtscMFS6vdxe1hGkybe6f7
IQW5sCM7BFQJXaQxzOwd6Plrcm74z83dKttC5hII2/uj0EnZ4wZxPqjYT1EPb5bUiJLrFySa7D6W
AelMbSF6Nx/FSS+azp3GXYIdwSKu//cGMVKUr/hqe0296MMgSSaGmzaBZ86N7UAuYG949epbcktJ
4xM8eYnrDWhfX6TUe4MeDDudCOiz3PBt5vlbrhZmJvm5QYt5YpR3JnUFCvzrnY2ubqnkRie7OnWx
zIASsGe9XhZRQJaC8kuzNMrZZ6bccENKLywUMNQXDD99DFoC83Qfytosc3lg12czARFyZtgFMZxj
QNJ+pp4RsV7tsCNC2CeZEoVvQ2nLngT2nnMT6UO6EHIM64okF1mXwOPEtzo4Irps9fv3JZfApkWc
mSZ2Z6CDsro1MEowd6ac+DCwbM6SwU3y0dr2yuRWIki1xGS6vYBPlRlN5pJ2QAhl3RRYymZ3BPkI
XRCw0Yl89ShR0EOEI6o/QdrndNEqEsmt4exAZ/3SBMdGZNp6rqAXopKk+W+jlr6UiGYppjU52YcC
M029EO1VA2LDvv+FaIV4mFZFEorFr0vuiLhz6HPn3OirMEyY/IrcBuO3d/2PThkhbJoTVlu7UEha
dRh2XpXf3u3XUrDecziHkuARvMCndUX8RbckpZAP6oS5xQL8edepyDlx8b0XmsFSSCMQA2LncrD2
zLQxB8DhRDkS/ZDHMB/alLejNLA+oXIwUQV4p8PBBnchETI6P4+E7SXmFGl5C6pFo8GVrrp/Qiw3
vnPRpXpuXWv2e+SLrw/wIUUcWYcMO3fCJ1cgIBf2Gx8IUKzWVvNVXo3y+kzZtlawxeGQHzLN2yIZ
f5/7fjta+HSNkrkyUAbnBGoDJRaOTASQEHduy/iIJIN6k2xkSE0UO1tuZRJiO+2X4kVY9TWdZL5w
34qh9vGEV+91KUNS0YY4ufs4fhMfcYpy0K0ZqwazclNVum3ajGbGsUCYiZkw4qFSUMoxao9g7Fom
yFZc/RUjL0Cp0BtIt0CX59BamitlTeyyjy/ia2vNeMgdZ9kulPoyOEbdgy5rJdOYmYdeuo5wDtt9
qsA0/dFaWnRUuBG/jlb7zaqqjdLG3XVTrSRxvsIf1klRqdip8d6Vir66HYHLAQCHwnhSeHFa1Ktx
TylkATdEptz5VNVXtnr/JM0NOBlo0IDqJxFw/bwKJUHN/TmNXn8bdSEfjB0GcI9Ow2RtG+12a80E
bW4rEt4qJHtY6n92nmzlQ7rclZmgNvlcCSjoXq6PwRETTkvzaLfBajBOuHyJjMl/C/9VVzJAv0rR
2c2m/ZAiKL/7Ct1BfdYhHDB8jPdZmGf9lBTzWt+Yp2s04sxuHMZpRnapWKRlF0OzpVQf8f+26IAe
DOJl7MKMb0elr+LtRvQ3c9uFBn3GoCkqYNcemdh0rvV8oM6lP1w+ULNV1CtKUvplk29k1PrS8uAx
ak1fpYDPTkq3JK00J28L97JRXzUx0nloxtaHffGyQKGWyMjhVNjiVTl8hib0flhRmZxRCLqmZR3V
UWEmP6/b2ELaFg2yoSHXgcUspTo4cTDCQ1Z/1lVddhfUDKiwNkN5iaeh70BZx1q6uFKWFRvzPpJ6
Wvoonwir7Cw/VQ5zQM1fOAivbJpZFxr6UTWni4Q2IQbvsPwHJym0jm2HcDOk7b57ZFVpFW8NQL5p
p+23yj/tN83U00PWKTyoVIXM1+Z5Gh1HzaG7OrXQz/RZUaJBP5MHChedx7j7ZJOEXkTC+VhpB3UD
Sr1H2H3ERjIFwaFEv3qADyJUjHQDgEDTRZ5OyRlwFAr2AiMc+cJX3EDiLA2HegEfa3VkXoEuYg90
c4Lt/x0n54+7K2yQYPA/6M3S6fhtA+nL4ZRag1dj+dZ/qk7hvdWh7ei+MRCQkYK6JsPuS/NGNEIq
O/OYWm58FWe4l8nVpW2XMAyRTmDJWmp4fzztgyHRs6J3RHJZWPhQmwkWwPIDV6X+E7Cz6jheqoZQ
un25/d/jqeYGRKpI7e242ciaLKWh1zoJViN8gfVkdz2Z2zwZMypWedWh7RE1lw+xyUVB9ftza4Pn
o/QzOilCrYcFb4Im4DoqLPUIx26B+FWvaQ8vVBoy2Pbb5TYoHV0UII1MYpma5vDrQ7/iQy9VdXlz
s+WFlO5/zb9Fsga93SmkCZyxwVZe+tLoDRPRRUe+VBvd1gkUX/4HMdiILOknDwg7IMQwhhhU8+4D
Mt9TnC/jqTX/xkoyWmKUmkhMPPgjcfeHD1uxRyb5H0kpvWNt46wnLQfMuGRqXp1aLmepS9ufe/nO
QLWvp7BZaAgxiRSK4Z2TIgHC7LvYRg6/uT0uzgF5Qk9MWuMBgGYK9OrbCjM3KvpsteTZ8+Khg7cD
GevRi+ecLDncLvdgG85E9kF0oQEoi6IuHdiWe3d99Vg/mL3siN2AgHOgIEO7FAHfVEHtjoDupygB
TmYZAwMCk5wrt9yIJgmyzNP+jVYyV4zpGBkhPmrFOhLGoATUh5WX4DLk9lQBjQmNqnE6nY5cpc3n
aOtI9cYEKOUogmDfjK/EJl6n+uRBxcCRSroThn/eY5pV/dWcucgXy0x3IW07C78r740Gs0gOTjYA
LcqnhOF+DLwpwXQpTt3nlMlCINn4HyCPxMj2qPiOiw7vRnNzvDO3xL4IXp4AZguRLHGC+QatxDSh
XJKaENY8nmW487RX0JoDwyTvHE5t5gKGTuUtPDWErwSSDnWDc/1bQcs7pyhPKwZnr7D4XMsvxySQ
anpEOjZJpfSG3BzgykODFEr/Bpalu/Xe8YF/SnFuVOwc0kVO8aOQqbU1NxGzOtC+7jSPMm8muYhp
17TCWv2Ueyx3/f4yQD51hSriIBhnscpNYSQFZYrBoTGdchb0WkGsVoL6tYwXcPBolRULEFL8Rp4p
qtDFe2F/uqAUoHAgtJIyZvSFi50zQEaDwAYmIFJ+eJE/CZ/Q5ix8vpN3P5zangxntZAAMfreSFol
8vZU8XpjmO8OiLfODdo/acglt1WCW04JBNPv3AdVAljDfroFRuqTXnpS810Z0oR6nPR4Oyivj21/
sL1Up+Hex7obua7onJJ7fA183DRRVWWNdXK5SaZK+TwBwJFQIQy5FJn+pYn6xA2CA96enDSLgqaP
MuZzqL6rjKoDhjzi+2enLiCDB8c4Ip/dF9EecjsmoUIH0Yz4G1ZaK6v5N0//2BlnmluWWBOOCS2W
KstRJRgr2P4yLW8p2gf/5RuVReRZFHG9tVfy1EXD7Ne512nFCfOaZEvRADMP6IelxVT9Rb8FoMKd
rx/2aITB668+ty0kL3HRq2ro+xJboWQ8lHKm+f7I8nHbF0P+KFro45MRQW1i+4/jwTnn4QOeRajS
tzSj50ZF72H+aqHtEr45iewCOmo10kTpTfo1GZJ3S3Kdh7W0Vo6wqP+YbvUvxnF2S3EFocO8YRkp
UKiOPE2SUlFyvwDUBBDDHEZb08pROCfXTYOeFf5BB7z5Nbty2ekrUknq/eofIvcZ12DqIhfrg3Kp
NvtK+PX5UvZZVjUIkTP9SRw0iznGbkR8MIASqoWaHNagFSI0tLzWKRwWRBagyiuTirxUM2gN+sNr
23MSpKDgKqNILLHrgT8A4kc8VgfFa/IkKu9glt9PTCxIXJuEDsj+4cQfwZ4CJoMuwSc0ZiArExX0
5b3nX6nBSjMrMCVHD6rLI09Yjyd+x4cIZ1HNSpK9tufTLRV9ndehyrcqLLSIH78sSjNMAXQUCU/b
ivaNcHof+Y1M9Hl20zLwV5q9k4FmmnMIK+GJscfd7ZbZzrpzGHEEw/+DdmwqtHMxtOP5gpm/BHm9
Z7VmVcvZ00+bk5IEDs+RxgRNJo6a13vMa4MEm6+9HZ9m1VvVQwFR+4Dw1Bwp61BW5hlqQyGxiEwq
CPwwYLyY2lkqVXFzDAGXtsk9Oq+pmaALN/LI7pcXlrDiOiflrV1uwowUy+XHbgWvbWPLGtvtlgwU
szlKJiekSU/v3wVAIK2iUWZxNMrdOO6Ww8Rf6D31CVGjHWlceiob2SepL3ZkTGRMzkXmzIldL82P
TI86eAP15hKsBzT0+X3wafbAf39PHWxUEHtqxHKM5zXCrHbC77GyVH4iFZBZVDfFExdW1hBFoopW
v+JP1hXXTdiiosEfmxEg/2rSSZgtq6CxY8QS7qPKFuVhHIwUHgDEBf/7OX0N2GR0/2d+TD3GL1KR
SFsB2wBCnk192Lkz9nw/Z9Z6FZo0xjXain/Hbu6d0XdMpsfXyhOcSFQas6Owy1Q9jW4FT6bkZnsn
qR0V3DGxxCufJ2txcSzc/mWGPUb3WXt+PhUO10hF6A9QUvQtte1+vn8i4XyHr8QpJ5bU9AHujH2I
MfhsFHzhM6whhX8qIoXTJQsF/MC0fVWBTG7EgaQdMWMUjVrPEUdqqi+evC2DbJDHb09+bQJ8k5h6
vPXG6TLnlW1rGSOBAaZpExCqL2LvIvQRHu1rkkDLhPUk8ZkcHF5XTUcsTY9KjGgXj9221z8DFXzJ
WatG4zHBm6UR3Lb9ev77kIxRwND0zhm+NF21hxDTrCLPYxSjc6OfQkjQuuj0++KSGMOHaHGfgwbb
MZLZ7SughQA+LQfJLbGB5Ordec+AVwVdRHy9eouvf5yQsE5xQtgAb+r1UQohr7HmaLN/KciOcgqC
5dMPbaDTxZzXtP0lFlwhauflGlVpPn3eJdfMDdSm2KBE2QcAhugeCL6pGMuL6eGHWInuUR1BDDhv
AePFrfeB3Y/fs1OqbaurTt3Q7DVBp67rAqhc4LfnY+bnbctODRG1OXmYXTmKGAuFRflS0v6myELB
/C8SPS5yiinxf//vJ8ZDZObzE+YgKN54hWwOw4oD7lW5oaOd0l7KdjGb9AELH4wUD/Vl8IJolahE
xuPrOcfr+GJhbfSR+TocfNNM3bVOBMHGWIZ/LEqTwYPmhnjQqBmyFGM9StcD+vl4MtPbozks7/zd
favz5lhdVWpHZTnWlx/esgisWOUsUqak4NIiIbdXvoOlqwJN+eCry32vk+mNm/HZbPb+UKuFPpsY
lv7dGpU/VhMm/eutdCnqEZudv4JkF5X7SLZ6xwncxKmAA1RnWr+ZrsbCWcxAcyBykWZ9yqHg73OI
Sb8dJHxeYBieMYR6YSYmiVOV402rNoiEtlKQlWxCS6MRpWGMXWfSseIx3j5qi+E8UDYq5Y49keS2
KSOCo4abUxYOSeRNCiA64xU+AXB87cptWnAj/Mn2PGpf/HHRFhz5uHfvV5ziR4fw2Izc+cGPC0+o
MJlo0s4QUB7Rt9hsRr6cewlGBYB3+DD8d6YkGhFuCJLwJVSywlvT7OdUGHAfbQyPm53fCozveI3Y
nS3CHwDR3qSLcMHR5SStBoxCTpGNEOVYmaLp5r1kicvJ3VkEteQef1h3x8BsBBMREtxgg8cz6JOx
t7tyzwLiBvQSEZ/2yjx0bUSWUwn1BF2l32BfHjxQ9uXB1lVf5D6RCNY7sti3Ze0m52r0H5BcjXzH
1OApkNuI/9N3POKnGQblc7bHYUoKuM0XCUfI2s9v8rXNcKPX2+CuEODYwZqAhlGGvHXer4wwhIVS
RDpFYaoX2Cwvb5dURHqjRLiBvLaQgK6rgb9jLrT5XidGocOfHUNR6dtKOzRfzNGNhz3bDHQn25Ca
aNVVe6vcvqtC0/siDDkn/WBRkvl51da6l5ob4SwzWStTIqQ4c8XB4zV1t3fNSNILar3htYGJa+qP
h0rxmtMdGAPRGH6qhBBxaIz///zFwVaOzgjczRFoMbCuKA1eoSTNZI7802uLfR0TQdyg8YOB2utq
+u6luBXq6Olq26jq6GyXzawEv8eQF9CkbCJdGGFaoMQBNjJJy81z23qxvZgQJcUx/noEiTIjQcrt
aosYZ6baLnLU6heb0RjYT2MjHBgcvszBwNq4itKudqqtNehVoQuxd7a50jiBdHjB9dG6Mkrgf+4N
9pSk+yfv+HSiKPyhdMrnNlDEj44910R+aBknPWbz8qbNv1yv+F9xjH2IX8D3gW1SjXCHSwah3p2m
TgYlRwgjlZtIuZqu2GcEQ4Y8cLZKYbWtbVOePdEF6mKp8QXEyKOVuX7utTYBLuA7MpaOK2/XUBKl
osAGoB38KDqa6welll4tdKno0KRqhBkvXtRmcffaPGUvdPhOJjluVpBAUbsOzeTr67xkRjS9S1bh
OPW5KaSygzTyeB5vTxw92Cy5QQXsakAsCcBMu0gtsV3BCn3y6IbyaBMnw8DSoG04tHhbdpMungsG
1FkSRtuL6NBrSL0E2Pu1vGQFFcknft58eazrf18kVkqDpxi8mUG6Hp2jwV/nHhOzsenlxPcj3UBs
OslRQiQ74wvEP0EM4qv/ahWrh6itMu5YK2bkDKtRBCz/GSMdp83Sr8qxeoJJM0WEwXZ8enai2099
F47Wo63M3t59Ff92dD2tCJof21EOxj/lMbTfn9t7dD19nRH4ctc6x36fqzPGUEMqPVKfPjuyFFsP
IjdRVof+K9MvFSTbQWOpI2Ft4H3AVM20j+eWEqEYyST2RPw1JgM9rZP7g0qTjORrBRgRaogrqTrV
EU3z4cBnZOe0tRjxWfMCRtKsIF7VH8bjlvbpM38OzxBCH4ApGIJFymNgyB/eVRapKyM8iJidxUHY
eF9Hkhi8X5Hvb7r0Buu4Wd8bX6jMrAgopBFt+3399l7+/KCJPEDR2ZRxSzvfzn/Kue3fnRTQ4OAp
T0UzIM8Zjrd8XnP8g0+CQAOfXAcTMxhRm35jjyzSJocVwOJ0YCuW/zU5xI5mPkshaF/0Vwi2fll/
Pwr9DKB3QzgpMy/GirS3MXqFL7Y7X2li3f/b2ZAuhErn+1zl3xFt/qL6KBqLxBoQOH9DW/dJFiWr
OXPdR/rGaPg8K8zG/z7kdplOUHVf9MCIPGZG1wMtVjsFxCD+R0oHXHnyaIbKax1hFDnZRk483rvG
EYOaqOxtlYhSKdN9yLwlMbljAa9QdjozaLELlx79Pm2NrDLMFW0LQyyMJAVREMRFIUmSb8dS+X/o
OGoXFY6QqZHzFm897PkPHSQZO/4Dwjaj2M2hv12emgwY70s8g4DLDnmTDFudVrJnFAImlKdA7XfM
43mcUphXbMQCtTcUXhEJJPQc2WZj9iSDAz6dSj6cYeo4lGNopUjnloYq8jHPdXs/ARZkx2rDCzsv
0kLpdkWTiSVHf4qUWYuDoTbw4JuD7pR0EdOVS0/3K/amArQB73wDw5I54PCRfeHKeMGmA+ClS7G/
z861F4q4jFrD1eoclcU/hcFKc3aTv/0zijoyXtDSWRHCSoJnayeFWfdN5RFx6FwaN2B+vkoPr3fq
9OyzzNFw0Cwtai9UQrg2vbyksUU3VXR0veZpX/uQmegyOocU1aXjQMroPU02VQPlkd6NMeIYLih1
DPEYl55vK7iJK9xq0sugIiH1GJp0NoQH4wIH0LHbthvLGIRGU1PIoFFfeg1KGAZ+URZMOv0xisFP
NQpNzsv83L8ly2YKGhSyTViRWiXD+/wNDG/lurKiZsGT7+Xq69WnCHJjDbN0/upBJC9FgDHhSKnh
Jf7iQiSPCKjGgwmyj/RiJTyBVC0UiX86Ucb2rswsDPITOMTGo60eivNfdpP/8+nriKF1LTF2+ZP3
msW7mjLjjfmxCJkKjFbu5snHXtb1MeX2JavEdbgNe3jXgV3RhqaqrQ0QU3+YZJp+zMmeOthX0qOH
EX/gAwrHpWNFnJsHBY4npaR5klD/PaLp/0nXw5gdJkjKyvOUVxdLfLznSBgcCiQpb31Zz7grT0um
UxDxBuRRQFIO1+9yIvLhuKl9d47iLK8BURNE1JbZlw1AYszZ+/0qvgJgL1Iy3El8KgENme4CSsgN
BzbrUibZ8l8K6NznJDSKJdHhp4Hmez10cm9sh8fcu18ZJU1wFu4Dhv59m/PIUDbilwqz7l1a3GK6
XZuburgsTCDnv7rhV2t58IXFyfJpBxP97ETTaeckAeJ4VqDrSpkyima3alTf1wbF8MW7teJaJgr5
bcqpeefn50RLkaDLhAttlbdLJBN5zI9d9M5HmP9BTn/bm4wfX3i6dq5hjqfrPLPFmgHZBLOg8bBd
/XUDwJw5pbFzUBPsRByUCmRqogSINV1oHj1yjiurLmPcd8vMwiTllb0dlgrT7xNkS+jc33WfrvmI
CgbvaMKCxJkuKGL714NDG4WgAn6jCZewu6GwrFp4a9lLIQtUWKNkdlpRX6uNYXJzXHiCKeWQsd4o
f4nxNZ5qJPOMuXychNbnvAs4LovRvZL4BmrutO7PN6FkkF/EjN1leIc4XJuxxq9PY22JZD3lUVCt
WU9MMvdy52FPKCwJR97yG0rJI6D19kpmBQBsLrZU2glC9dr4W20PJIYmDD/d3vEJxhOwoe8Kh3rW
Wczuec2zu+6JM5H3KiMDDu0skd2Ae+HGxBU0qx4WIx18TzV3GOkT2OGTY0MYWnBrlItCq+Eul+k7
u5KPd3pdEZmk8uouNLeej1/q4eIZWV93m1iyI0ugwCxrAVQ/bcm9MCTv3b6A4VxOntu5aBHzDtI9
UXdX6QrY9Sx6Q1hwIMPcjaumVgqvvquIjzQ03XhqGgE5i624E0emya/RXfEoYL9DUH9YSl+z3lu2
iQMUMF8ZGJSLHXMuyEAKOG3Op4SrPmQZYbdXy/c8xWCnsj0X8TKy/0MzE17bHdsJJkWFVSD9u1M3
R+YfJkDjHSSzcexfKBoG00Vum50Bo7K9VQWkM5XpA5gtuzCyQO8c4PslTWkO7Of63MUxPNlvWhZF
rjbhxxnbpDp0D/NiVOCXu/zuuitSWtu1TIChmo9AXg84zYC4qOqAwN8Wi81lgD2JzPYX4dUmrOiT
FwyB9dtPSGw0UYtDV3fPLGVxzlaSrHxQofMNL8ViHFUpLJ9XNDQkKvloRfH+PwFLD9x9Pdt8I4C3
igMvSp6rDyNsjlLX6sg0YOkbGwxTxzMM3PyN74eL8MuPDkuvZULy2r++EXwKjYqeW11ci54D8TPN
wneOE+lfOflphJOea0+iyHUNW3NAHq4+8gppJF70wIgu3q9vo/+nI4iY3JTdQ2nESIzmAvXWIEVv
gsQVAX0CvqZJzMu3qaKztdLilUDObOoivceRgg3iBR5go7DgmeCZ3dJkYCULTjfZpYJ9oNNwuJya
KT+T8iU0jN2icJIWB8gubIMyYZ3vPkt8iNJv/jA6nyFi7mvKqIsN13G9GEM+DO3woNsOyJZ8Fs83
aknpTYDf+EY3VJtKJ1UBGC6eGnwdzxKy0eTAaw5nczlolhu0mfrpPYJjcM+g1thuoCtwBcZbHmmT
rmSzoftKCcm7wl8ygW+dKW2Ycdj5zP/xKvgY0FfM6Tt12mw8iOTRCx5tLzL2gG+z/9Td4TO9elJO
dcELBiEaj+fyylrXZL3VHF/dCvk9iw8Z7iIKmZ42ERoRnGiGZ/nDF0dvM2ZL0gzNZKVsCf1fUgsD
e/Wc6K/vvRnbyFjbIECslR1wg50a8Xs9hUp8rlLd2IdocBVsB9ZvbMxFbN/NXEjoETgE15NW3SA1
/USQDuBLJMSuYv7GbDnLXtIjBXY6XY+rJd2bviy4ugtN30hON99B5tTxe64Nf/daycUP72j2OGaT
QEXXw72QAInT6Bby/0N7FSFBumTOLlKrc/Zz6ZFik3JyFw3MovI1DOkXX4ztUSGA34R763+nKToE
OVetwRDDMT6zQdC7MDTn4eAQ8J7k7iTl52aVMaGUH06QEetO/gknTrDUdcV1Rd12UqzDIF2Kf2+F
Q+XpSVBjwTVLG7cWNuTIG+ffYHQDKxFF2G8N8G/kMN8yfl1Wx18g3Vt15kU2dc9/e3JD+Qoh++ag
ovtcFilA6+aSRY5kRnEjD9Xv0UsWuzcnz+kSXBHwSsWUhke36PBSRpaklwuqRGg9DuSsuLJwCHv1
yOffDgmDLQDp8K3kSbZjz7tBWWv0QJsmKJjxs6l+Qi2/K1/ePDndW5tNwssgTLRBcRpujmYH65cA
j9T64IQ5VBtL8dDW2Pt/tUR/yb8fcEZRPsqBJXNnFClEMnxuSJ2Bw/5v7TN0aad3ws88DjP2gHId
H5nPBXiR4A562MGgoirhKkQWFw6QPHqR7iUhJbj7oMK05ld5VFVONequdni3X4yhiUw4FNGVz1Em
cjP8SHhbVlUMIENSxfQCIt7K6y2ajTuZ+OXMnmzb3kz/zM3ClUXSw4laecUtc0Rd5vlLcERg1W9f
6RtHt6BzAGNI5cPTXtHf1TgRdJlUPfrZ/PwB265/LVUUhRjWXdCQpvt+pIy63IDok/4evyUCWujR
JYnzZ/44a4hCIPFKkZ/TwKQAlK1FlBfYXLFJXmmk+0SK6yO3IkH44DB6oD1P7s26xhXtaWYN9ca8
8q854m4d5CpfyQpZ+U0TSzBIUBkLQO9NTH7n32sfL1v/cvlC2+bejHCZg2JPQNCzLVFYMi5v0b7s
58CVx2z3Wsu/dCkFpvWARZKrT07CmGMK0S2j21YTZHpqe2RzqGjg7/+A0U5Njl2Z77QyuhaL4k15
U0pzYccywvaXNc/v5G2k8Iog0nc2UZbJO1VexXRtbFCsCGYcL2cUg9ZHxCKLoy5utc8yxKYiyINU
AbrvgBlhuz6xLqb8d8R/qhVcKo+S3tLhywlo9fmLRhF+0wSjWelbQ7sI+K3GFKzbxIwLfRigOk1A
4HmZF5Wk6wD451DlM79zFWBhY9YoVechlZOfNLITzSzjF8E5lmqdVSD5cpCIotIcgtwVjfVJlJs8
fZeWfl5X7kVxDBt/ZMvCMgwLKZRXyF5R/CcjtXpkpj6om8qOPnY6LvtfTFQNeJi11PygMRo3s0zT
XqvdWPPhFZNC3V4hVO/719aoHg9gRQOAl6IjuoxGaxjYEDu9dHyv7E4Cl6zFBlOHONw3gcqKW58F
nPBjT1wLVHez1SA+IHHiTnU/VVzOnI/tg1RPNtf9r9DUXZKPFEjN/PL59aFdUvo39qDTfu0exAJq
IaXEOn9Kn9GOU7thmI71KiEAFI+AjPYPkyMU36MdwRKVN4Uol3vhZlcvGEE0U64CL7oDoEwHgvO7
37htUQAg1/BDO9vrFixb4rD0sQYha0FOoKwa0cuNImEZB52mubppkG97mfGrDivJoYhIfuR/1Iq4
bwBQYd1sktfNaowGV6dcFCPMrBJtRKg+lGHhW+HfyPM7uSS/X37WkicVqRkEBw9TZk4I3CpAzHmK
tjNxtuBMGunpUoOm2FOt9vcx7Whj9BxIdGKUrpVGl77Knm9/VyvUDYl7YNvwcTD075+1antuz/93
IU109LYW+6FM6Z1wizjahahIWjltlVjX/Ttsz8ANHI7tdIaQeaSc+JU6zWobZkckrPT315T2E0Of
6+PPk9Twb7Enu5CItmmWfiyycEqHulUe5Jk2rIeAfaxBgRna9q9tXgpeyB3xXGRVHOpgwPjp8yRU
M9cTcWsZFCyf/Zqhdbwgjv0MSO7yuctjmuioLEDxW+kGNPN0rOeMnWEyq2zZQyCe9Zdr/1PziC23
x4RZKPd90qhJMdKFt/pikKJApT73dWmGBBFPRBETUV4MFi83ybWvERxohJUgPJaFsEEGxdY7FawH
AbtMr3FcKpnRWTcUvE/rwG8++nHnWM46Zo0wmgLu0GcqJSSqCuRvgBWxBq93gv8wdNBczOCU+Mah
GTBBRBxiXuC6BgeEnOAMEvW6M7hZTc8xCiYKmWGr1FeSWZ2nb1l+ygiWlPNHOaTTdTCgXZv/OQrA
9OAnFHEy6597egwXiG4TxANO3Ckpt7BhXb3JhApMaANC/azjTDl4jDC4c2OECDXjvneCUgYTCbdE
o6OCWni1KT1FyD6Tvuel8njmdZOClj9C/Ec19LDML+e2vQDDsA+QxQVc0tJTrfFGTNjXJa/z02FB
FlFJLfSSscXs0VtlnBT1kdwOFYFvRPGmsvOj972asrBVVTp/wGyieroCLQbfdUJu7rgo9wL92NdH
eKt6+wl1In0fU7q0li5PuKmb2KAfrQ8i4nxrRzNwGf6Yia3fGb1A+KTBkPXB8I8MpNZloioyrrvT
/jOf8l7mcwyEIVcuwa7f+d5BTJU1OBeHMIabaVIAcUb35zytx6c24iyvLboSxxXm1VnrMBenKBd4
aaic8V3kqasYHp2APADa/OKR1i0nwB6WM55E6gBwFsGYmXfwyfM0/ieW5c5vJdM3sPHciEKFbqZv
ee/sF/0WTzKDBE4jOuD6/sb/5MwUaYBjul3XUAuWm6ZIh31aQ9ls6IMTSKZSrklUT8I9fWW/3AZr
YMUmNJcFOJtTg7sKwgKDMvTkRZ+grKJyZdZdL5znh+jiITKyaOvBoDTuUTbJgZaicfYE6BYWwE9R
jo30bmHgavWVLwHMnye/AA+kbC77SrxxWfI+rsWHULjNZAN/zRDYJLzxqfzDXUdl4Yvs94MSjPkB
iQLrzCdQZ9LV3a8y24qyVo3O61kWMB8ES5lRGTv0/aV5SVGhIK4KF33k+IZLY2PDtczSVuEdL6Y6
BppoyffArx/aIJFw97ux1qSM2+BvtKpTI6a2iJB934nq7n0rUyDVkv5dJWYjLLMLWpoLlCSWuqzd
ZKEIEhbrrn70wwjhA+NcYsn8xj4X0DyZx1c9RDui94b1q9Ge0vEry3RrkdvpQz0ADFcmmcmILbuX
GqlyMWF4jBMzoxUqLt89V3+bolLnVYdvHXZOBbjoNURmRotylb2BP/v+Fu0ZdT+1jVV9Gzupn8eG
hdFOPO4lYDuH7fU20wI16psDLOffRkoMliJxXxjoBt7fi7rBPCQ6qfYc8Dm9FnXUTG08SsWO++t9
5IbCExVgcEA0/lu9UWlM3AhPIjVscbDsRTv1/DEs2VVMLYXf9BCKwasvPUNX7tB50n2aOT2Fi0fH
T/srW1OzthqcXTQ0K45oQPuo+Wwnf1ChAnBypgqxR5EZAXtheMtgDyaTtgApcRyQtaLnpKy3Ir3T
1rf8QsqlxIg/rEznivUTtIeqKgfOk7T1XMpC87Ei6Z34IkFjQAHSnik1MboQDUOgZdCwb4D8ERWq
pX4EEMYE1rDxVGqeYmD3GI9y8xDScfZE7IWIgIifAL5e+bo23ahKSAYD+od/Qu7y5P1Ik0YHFY/0
5nIJUS/wadrpFlhGgV+lxEyhqOTeZhxm6R/+RboMSvempgyIOcoPSHd7hHYgihxDkVZHADlOpbNx
BIA+8n/b+rvsXHArDkvPaotaAWaJ9mxNpy8d51wvhn+ESB2SVj3radDx3h7akLPxl9kZapbwmLll
T8xxtOhpxR2t+nnZe9wBnxOrbyUJtGGjbQY0DrMcrGXpF6aN0qcP4UoSW3Aa18ai97RJhHgni3k7
aaO1JYPeViYGsKiAt60jVHE4O/C1SAQEnhRfVLF8digw1drZqNUR5Vmplvzr1t3M1Dn6I0L4p9zg
NLS3+z807lSRzSyPaytDywOUAC/IPThA+6QF/sqlTXoBhjATGemhjdj0inD1fupEN8PeZ8oxcgC6
B1xvLxsQKcLE+/UgxKLJ4dkFroWWha4Wwx4t4sbSb00PcMzk/ZJRArDz73ytjn/lifZpsRQagSm1
bJs0ajJ2GtFwf4qKAYvsjuIJZ4/F4OQjTu4iTMv+elnMvfY4yyKYFGifiTanqkywyf3pMVJ959d4
frmf4PcuGv9uWu3lSJlrrFAYYRX+Pp5hq+D+0rkhTgxnqxxCNg7VB0r6xNBXax7yH7mGcbbNgQQ0
RRiuSm1rgkXEYpKTM9B47RTZ5P6Xv9B5cKiyNUVltfCXBZvv4T+JsD2WD4yj/ukQXKHviiKhZkbl
GJgXpYCOErIfFmWUeiVTiFFeFo5jUSXD/E81GFjjqtOoUYN/niSt5hAZiqLW5sge7Ao6shWGuzbA
QgzWcu6tIkiLCoi0AS+2VbDR+D/g1Xm6ek00hZk+gBFmTYqRtqX+8ucK/SHNcA9MqbIBhKMvbRvJ
tzxGt6CNzeI/HXu2oTu0QdSTUDCz3KAw4puNeCgZx2XaNBl7Zg3BjOerCD4wwBQnyzOK88OKBlCC
7wWJ/kY9pvBnl6f2v1/zmBXIFT7apsuKV4VPFulshjhcpCklpLlF6X2+YGU9bcC9MPslgNsovHLO
d7t9TiTsy5ksB0valBk8LAIPJr2D7ROHbOkxPz4+pqbC5ei/ArYjN13deqnwgDMASSbI99yN7NsB
rNBGrZhLp5NROF6dsNbilzvcdfYq8wuxi0+rZ5iSHBCqR6onShqIKzQ4jhLNUUZLFeQzTbixbfTX
EAmosYXMjv5fheWfi0nkv4ovo1ZS3eKvNtjAnK5oHTMObKfxqGftwt64od1uF2GIvhilhkRW5zuu
WjQYDm/7KO05j7tDdlTx9EsH9vEgK+JsAb4UqpmZbjQKB9qBxDHSCWpYNoT0QI776VgT1HEJDq7i
P6LvZdSoZgXNKgILHcvl7bCd8nrVSzet7HwgAFzb3yclBtbttK/ONC0FynAFB8t84+RvjNTrpGP2
AxGkRaWHo28+ypeQJkAyaqnFaIJ0eBVPgfA+tTZHRzH7L9jpu62OI6LFHqzy3TpJqHYaZ7oG5Xrk
UmSRbx1HEmGvhuje293kmDVNfCR07jp1oapE4SPfDRYPiz/i2qG3RDlCe2YTRAZjlQpA5PIdnmNW
FFH9/IiIfPJgdtjEpCzfgfHjD2u8/Agxk4uBi9vqB2v1kM3dHReI0G+LPIbKHSZcuN1PrTkxmBYu
Yc014PLsAH2ylX2xp892YEi7Vr6a9SugQf9UmuZb+Uh6/AGhQ7qG+Ai0zYtaPOj++wWEQ7C9KtIy
Gbw1UFfXAC2Y3sqiod1yR/9v9wBswZLGpd6Mht5WnPt5G63WnuqZwu/W0gwfpzIpdYFsP7wdg6Tj
pLkxn4x4Nn2xm3mJYhrHo6gfHa2m90Ycb5vUIOmFhc9x5o5FwBTSYe7f9oCkpluG2mWWvsu7h4mI
U2hvVztffsbUPVXi7ih0pjRWbuQ5TGMxkn8siAZIvcn1XN8gSSadYsfO94HUEIZQBwbPNEdOLoDV
Y3YLqn0HOtTQEGN46TsADlZSj/uKRixZhiJzBa2eVryhSCV65jby7y1ejOMtsIy071B/RspAMyJx
JBmYQVBUlKLxTo8oFA6W2F7lLitQLbZJ0kHhQXyd17oVCysYSOSL06iGk/PcLuEWvW5Gei4+qkjM
boq+bp7Tk8ifpwQsRRbi6qQJIMgq2xRPIWPh4BhwPLZsp7Pw76jLdg5IP0xQ/IBA7d+Mpaq/GVU/
GDrVJ+w15b7J1odPx6F0BZzWjJnwGIvQ3u+TdRHK9qHKRVED8lxllyDV/mbDGw2Fcqssv2eUhwfg
qlbLBBuHEYPxuPID4jdOwahgRfY5Y1mTyZJpdT4V43KOCxf4lGirR+tVUIxtqWg1jlZ9IZhEUd3U
ZTdphqQ+8YEkF3xdaGj2Kvvreiw4h3HuZDSPX0/qZfirXfp3Iz8uWIxxW+/4HlMttHjBIo+Ns4gL
HwoW8CJ6ArWa1AayH1yT/edMyCTztHuZ5VYtEEmfk9p5fMSMMClGUKtROxLEZmFUOgDNtJVtqSsg
4x6LryHUP+zRSC+QVySGZPVdXFrd0PE066455ibl1ohYk8D4Vzoet0RdC4rX+/XApX1xv2x+/qNB
5wjqjLeqaZhBvvfJLv5OS8Vg6i0ivtKEuVBF4v9SyYDV0SI93o7JleZwaZUdJVCkNji10/IA1FJ6
bT4QYMUVtuLKZPTcSs38Z+daE93JCGTPLvp65aUhfindPKAcW7S3KgdkjIpSJDRCqXGjjpKCeBsY
eAekQ4ExnLT1ZnrUxkrOL/+seSBO0yyCZZi0bBzO7/nVA9SQkQ7ezBmG5cJooYfPVPojCe4vpUy6
uqGZS45T0do1ZZcDZWKIvWt9qHLerbCEEm9dgK4YytQce/e87myUGWUTgG4CxQBFAbvqlV2RguKZ
yBBNwhxgovcmNXZGhrT5r33hNTAVi2N5owXCFqA2ZsudrSAiECrLHo3SjHRDfLj/ECuNJpPSg0+L
0HXQwZPyXfY30tCYTn/6hrF36fTdgg8XernqXuWChzm7Hhc7K8ckyAI2vu0+APj+JPZ4xRsKEt24
5lZoCcLUq0M16IzacgmnqdZ0uNh7PcZGLP+4uFtSTzvtfKPy9vT3KxbhgTak5z9fMQeymFd/I35S
9EeqjH+iOOhy+kx6e3XNZ/FOYiRk93PvPCFIs8whCeL+gVOpsc671ZtSTD4VkvFYXLrCWDTtrKPa
c9L9kr1UrbQRyPx4gD68fy+/lJxlHqWjSgsJ4E/Mp029zGl/lXp3VB1fd2N9k/diX03Fj9J8j3cX
TdvGHnA+LgPbSbEp4ESptvJVfncd7U1L6EtaOFtvWXt98JydszunXHZEcYMk3Sg2Bx6Tco2VO/AK
3o3ToJhMvEnzfSQU4T0Vd8HY54X2LWm+TKnZybdZgAJUxjhZvVeOJokVfGPcR45IQbhUPLCzJUSG
FDV1c6mtmzW6QMM1IBOfNUHYdgW73PWZ7Rbg/fslg05IwpNx3ZeEnrF5SmQW3RBnwlc1Xd0wtldW
3EygZ6G8QRz7SYxKESAg4shFEPXrjdezbjJPzxyYOhKvndBxCJZ56z/f3b63mNnpWAUgWIOI6ON/
Gt4YdJ2gxX6DERRuAEWYhM9i++ms8ZuDjoLVeucNcwrfEymurOGhdqAlyPKpMNCbqusDcBEAq17q
pqSuTEyXq+UbEeVEGtlwy0e4V8JMXk1iyS2IsuOawDOvfwahsk17G1qwferGlu0K5yzqf8LLqQ5W
EEwq9xqx/2IkOESkyKT+Vjw797573xObhqdJ+ZCYAcX1SpZS4dARxXVzunsUXsHt9J/xT2zZwt0R
8uR1kdKLdlDMYkwSHdw+zKTGWAFoS5VSKFPNOI99pmsifRj7DalSd1prkwdZITj8M4u7GMA4110l
xi/iOsKvV40y+SOqIO/mmZ3SoN9urhf5ocsuz5AWnQxMDSNQcRC+JfyTEpgsfcFNC2m0qouJcLmC
WEnvYXzZ3yfv4iyRWFOoxoyTnw8usIvzkGX0tSL5g7r0Qsq+6JTYTiTkokKXOf6vYOPaQzC4d6hr
B4/3Ux8L011zXrKE67IChzWgOExl7ssZ9O4fYe8CkvYJg9eNP054BfrUAObdYxDlom1ZSKQvaxM8
KHkVDu7z3YLX3EflHwX+Wbx8yVLQj3MlOYiBQMJPBgepOZcVMl3BWy2BblNfeA4befqNqqOTPgCh
IHJRMNpB91+4jkpfeBsbf1L1n2Z80fnGJVLwNnmdBCk4gIsnup45TTsxlFN+bjGkb+T9tlqu0ObR
XNlF5zkZepfOC/HH7kPEKP++gIZblweqyuzTrJU0Lzd13YEd0n3cCRcwQzdCsdYwlW931XdkEWA0
wHJufipWMqNfhbzP6ptpgYUUCN2uR/g197JELgBQlRDKk4RVKFxGnP3GnRsqUOBVeYxZNDYxH5B+
1zIkt3Pg11ZBy2o/Rdx+bk2q31AJhKvUvphAMx7Dn1wIq8ERTtcLd3U29i1zlqBHjE0Tdwq0MJIn
Sgi7r5FaCgYquX1wLMA19nbZGhPL6zlVc3tJcSZVu5MSdWxdO4o8jWeXUj0wzFMImZcrj7Hd+ZuW
Rmo971OnfIPmjLUFbZC4m4lLTNBOteQnRKXnlBHhWrp3FRMiYSRRuNrBNjBt+5ZRw7Js7ujBJXlq
cUTLjdSHLEQNZz95Fs8BMooxSKVoWOHPaiiHHwT9zLSZnSV1eGrPxe79ForZM2uDq6YYv6xP6u1/
3Yssj8xhZEuHfEi84MzcfRGO4Dm3by5GufSJijspoL0nfAV59etEfF00V1iSjEQnPkovsNF/ZGPJ
gwYuc+39tQdyzZeX81k1Gn0yIXhor2FD1mAqGJPSJ7c3xH5zP8qoIuUPfmrfGqMyJWSbuu+DGGWr
55JQt1FFR9WDPXkjqq7l4NqspRW1P/yHVHXyAqdIK28xGOE4wgJjbdnVaGdQrqp1MTZwfBi7CysX
GvMYbjJa1Xv+HzI7BhJ+OKJFcc5XHyn+WSugo0KrvAedwNs+9L7OIYTkhNTuojDxcmirO4575NyC
THKI9IGZMKJX1aZyNtfJCxwnaT1A4MEHXFewUclzjbChqstmtRnMFtiycx2QuN2L4vDLamCfm96w
fro8Bj2oDPRt6Hc3mdxKZRgkuHi9rtFsOmT4m2GJUL/0m6IJtLO4FBIJbvG6xwQivrJL5+vSWE6E
P3JlpmMRmWI4XqcrswnVy548s5cN0ZgE2SdtE1A0/wemP3Co4fmjtp07n3dTKAjE5jbf5ca/0SDG
rTH+6+OuuCWcKjpRX6uabUN6pts7HpDDeJ2/Ikgvcrkm9uUuRaO/q9HVzMq5D4fH4AcGA5XDqqxe
jEPP2sCEVc7Z3foI+gSSGDkIafMdpkuXjjL3h0tEj5p2/xB5OMPKOHGB88dPtunSG8qlYJDGIHcS
hyPkttb8GeOuGzOUpeNFEtkFuMjRJ6Wei1N/7K8fP+6megsmppOMyY2F27sVpO8NwZtLdaeLEAow
naoS+ArJHNcNKBFZcbbqGhMcRK+cZzCaARiBpD0pKIlHQ7moiWqXZs5mqrZ1F5FAsvCJF1oqqSyO
PuVuaBo8lpiDEF7W0qnfbidtGmaJAP2DE9N4mjp/KNptj+LalZ/PCjQlXx2bEV9r8tEpzRvbiWmq
gBc3yl520SUS0MLSsvfJhX4MtdgBLnCzi5o65HtyiGR24Hc757SOW4ISIsLUS/AJ9ztmBeHG3nGR
H8yLj/5k/SULSB77CwrGLn68KvXFKuyGGSZNkvX4/Yb8w+r6kScMNGHUkoiaCc6HQ5Eh+7JI4ZQg
9GiDUIYXc57/HsYWWMSt0pZjUbYJ4RbM1jDjkkRV508P+F2JUoYEgEJgm0zgLbsTk2cQ1ByVDudB
PPz2GuKKmDztKZczLFhF8IG4TPx+zWp7RvWP4ZXtbPK9UVr8dexQ7+clbeTTpAyCcnbfbghOlfd0
uh6a9XXZ1/EcbyC3QXq+nV2CYeUBwFwupsiYKIQH13RBmdUIsqc4ytpnGuWXAEZgsDlEVtuj5x1x
2BpArxUBFoBGu8yAVyP1bcizg/wMFFIRb5heKbps9DCbcAIH3crPWGA0z2bTvGAmv+iyEpxGIxsr
zACt5pfq230MlUzVicU2jQzye88qAs/7irOeHSoGUO9p1h4q5eEKlgo4QI9DW81a4jUNrYrIEf9I
Q09p6QGo7gpt9fsdJQ27ZRemQhNtDh2SXFUpoUgKM1U5DTleyO02NBr0Psq2q7xkh1qFColMa0xa
6l3LSuMpNyhBCApD1one+mkqQyeOyIBMC08PobZ/PQ7jbE8aXiDSIPTzn3JQRRBRI0P05zhPkc+4
ehrsZQGjNEZYxRPkddKPpBXjItCiwAhasmvhxQKTe7BSB12/AbK4nTwhT5fAj3W9OXuA+uaWW53x
6awD08IAZOvZZ4gHJfMnVICd1icAhhLRMkzzye044G5QW9oj3fW1FnPhCsDOQBGpLM4mch2PcNq8
XKSxPXVsJgHzPn/nrgCZMvJwrPLsbTD9hMoiDFFH0giuK0b5ejQlc/aH1llXCUqeMtF0VL7NEwRt
YCEbY2z93TXfnxSnW0HizXPXGc185Itj6H/wshNB0CbEctrDOyZnR+gJ+YyfaU0N51l9FyuMKnHw
YEHVwHOmzaU8zHCnddAO+Lv59b9q8sQUWBeTh0tkZK24ikpMM/vgW9eLcwOQaZjOBb47So6KE154
5QRQx+3vhUAXny1FbiRzFPLEKx248+0AU5x0P2oNcqmLMaf8OwlHlSiLdW0Hr11BcKn2WFD0J/Dp
DB1rmy1H6mtG+U1tgbu3GKKsTTaS+pynpOYchTxo/ywvpiUt71iucTz/zZziD++8OuxSWu2jjN0c
COd7zOP54WpL5KCSLd7QlIanr8g5z8nZTmXdLUwW8C4z3mPNiHwDykhqqoVN1S5/t89AXl4i4I76
7/KGL8HETp4vcmvgwHRk7mkNBFTcpQTE+bKJMxpzc9MXP7VBEnTNbxP7mCAM3iZfpEmGYnYEyDkB
06/z+6u8TWXdIwf2JdHyG70Eby+dI+CAiws/S1Wd4Iszxnzt0qty9g3l8OCalmr24bZormWsxQwz
GMzRdzJH50sodD68wOUXbWw5VcD7JLGzdfwU2+nC++/kHjRQt/Z69gEOODLUfHHlr/SzJcFPP0jK
zYJmvQOUgaJawjbCmgCHcnBCQREn2gvUqi9djsXsP9/cufKYKpbqFXVnAB5f1ZT9vn4zLV4pTNtd
Ymc3DHUH9IG8Y0Dhb4o1MDFi+E37nPpV9ety9KHyHhU3xwynrj/42Q6VQ09NdjECBCoQe2/gtBG7
6UmHXngPkMoFwQVJv8gmYgIezNZULTT3cMoYrJXe/e48XegyeFGGcSys6qyTSMjMOb+yO3DNASri
Scz2spBO8gAVe2T2reiyMTD+xDUSyw2RQkIFBjWbMHORKznj4t6eEcvufycEqeHDWuHqJfMf/EIh
4zvorBLdA0qi/+WUJLQ/STVHeFuykozVFl6PSsANZRzqVVX7i9gG3coZdJMK52MlHqyLQVghv0VZ
hk1Dhehj4sZuUfpN4nNq+6+lyPbRkLLXNaD46sye7cSTWjXTMManajNn/Exp8WFlaZcKdmfGX7zb
2VcANBR+IC9if4qchV34ukrsOiyhx+Tnua+hVYl8/NmGtkH6iX1hcrzHnHvHli+LZ8KVEPC7R6fl
yAit7jNv7YgdbZUWOOTlz2nP83c3U7kSGlvzTRnbIROvoL9K7U9lFrzxN81HsRyCD5GI00emzHfY
WeUWhVltL/fCvNEhe4QBY/BFpPNDqxqkRP3EK9t2mFGQJ8e4UD49SSx32yegeten8ffEUQ9DBDnj
2q2viK+PDGSrSG21Eafj1HXlIqibQJvM6M3RdcN+b1uo8sU4NpA6qzHqDAabFOf33ufLPaE/bVc8
gufdv4kJwYBQYUeAT4emCka4VRq6E1XekXfbVSf9foKm+nmYcOgc/Cj3MVr26TZyDrQEvMkI8Ig7
rs31qv1IXi04DzEqlj5NR3I5xR0RqY/4u4sJG9lktUPJf0MPFStpMktrJO3tckABDte75ui4Adsv
oxFZkcADuhwwBv6CDAI9gNOkra9wRwAGt5X+27eYV+NZG4AhutC6NFPmcVIcPjmiQSDVoOFu97X4
4XFnPWMsIoLQpg2qX4HwklMLdMtV1ZZLXNPmgjZfRne/Gp4aIdgYlXILZmah9DJ9gRQTU8RU2+pC
3LY0vz5cD/xMcY3KbE0pgRT+JajsOsBXeAcfOaBJPvow0Uye2Hu2VXg4bSDGDpNmxKsocFqED2R/
TT4jRbW590c8jbMHTyIvcrFa5LeV0RzW6pSSipmwAJocZ4Yr2owvGFZm1bare6x5cHrN9QxlYjo/
fbbmACs1cXGvkQlxW3bCBBU/83wE5qiiE6bKBzlCF7oy7jVxprVCXB3H44K59dty+MuAzGIA3qHI
/48214aF/I4aPpWTDpr4OxeTXGoK92d0HSkNtspPXOuJfw3zWtVkWGJxGkCkAJl/KhBbvVuRFjkW
Gv09XGQHCylReA94dxOpfqhg0R52Q/4jUysJM59jlCSAIO0WDF932s+n0KP5EAQ4idvmWKGX7Wv0
cR/HcfbLv/X1qN6xN/H4AzGrHCKPffIldSLxG0HnfF245MN0x66a3iRoWiqNk9uC/wK+TrpM6Lnq
Kh6qikjOvbbDcKhR843ZtED3W2HW2hVMUJPFthdetr+lQUfEtPCFUtMaRLmvP8GUdPSlp6D+NRTL
OQgLHBHtB+yPzFWf8cu3lfQmr3S6qS3g75cdPSUOVOFYt8/lM2dV4ZbMYpY11ZF7Tp001N2/qA6d
JmVCx+OMIY7YwsMLfD49/+DxCgv+wBXHlPO8WC48NmdU6DjV6I3JXTBarjv//9WxtDJcWpy9oQfC
+inc+uEz13cDdh7JU4u3lSVzHKHcymorvLvvGKCqqak1IpkDG41iU+7lFa1lN3RiRN7xGcAC5aTY
ACHSCvYW3graZNvDYOQVzLe5HjiYdN/g9IlTWk3qRJ6ithCd7IhEggFTitBbJbBbuwwhQjh/p6aU
dbB8fZBMjXBsDvc2So6ygzfYfBujmFQnu8f00p/kyJMhbJVZqdSjCNEHUc2tivLE/a8WkgWEEsSs
k1qNfmeIqCQi2pt40jI7h49tRvM5gOCRXbfgiXpz70BtW9byQTf0UQF0jwO+JniizKq0lRt3cUdi
jEE96cDief+u6XCf0/twmzxNsHlgGR5K/xu7AvqNJo2+VV68jsEa7CGzQN4dfsGAmxcFQgszEqCW
1GkX1P+aKzxf5nO7fsuClDAik9I+RSmxpNwxmfNT8NIkBWVvGklpNrCgi+7D5ZA4UypZmh0jlS3w
zuRrLUgnGzfe+iM6iXgleNl0PELgOsDg9p7uyjaQgs+u+tKcXuDJcWWEvLbxvsYEhPPx+CsEelFy
N5zbRXHUqcWWSCgNtHxNFo51V/TcQVMSsJ9kwd991J8+DFkpu2FpK3zi39GMB6s54Z5tDzWXH0oa
F97+wXo1Ua4h3od1U/7g/nfZ/pxjqYsTtNwh3OlRG7E/GGxKFyxlLXSpI70eSdPipDLgRJXKUoMp
dN7IbvFLLzXf0hHshN7uKZQ3RxTl4IWGeUmvT9P4po7nY+rkqtuJzjMC5gODRh1hPt0thjckJ2vk
esmhiRti/psywaU/COiPMTY1aqgWQQBKtggyJ65OGDs5EObSArduYo+Vlv3g/P2/CKOulRAlQxFA
fNAJ5vZuj8N6hU/hY0L5I8/okQoGq/W3sBWX5Nc0PrpcB5/Mf9pvOFPjxOwBrN4NEmm+1Yvzpi2R
nBBX7Rm0dyGLUmRD8plKuIBzQvFaE1I0Sp4HrNeUay8nmZTcqoPfQ1vAkShq1HydwXD1YYmaWJrr
mnr1Y1JH/qY34zDUsQz1wDQGyqIQKoooRgrSh9GMPxftSsAUZuq57OsN/WP3MWO8aO4G0gaKbO4O
RuUUAiKCRr1SQoYO3q2HxRyp54+GidMcSOKdp0A/+3SnbDFi3igteZgzVTthbHjm9ZPkEYtV/xmt
D+8+UbqaDBwD3ATyW6mCdi1GOb9Vjg+TAtENvm8AgXiNmI3nEem2l2oTG8ZAgJC5OPdpeYA7O016
fYIbhqj8fXaVBO1G6TAHkT4CHfuHks9BnGGFCvKL8WiYtUdyGat7DxXulfIyXV4wHsyk38qucDNt
eU1ejBBf/AYLiLizgF07y0oFF/IhvU2ZnL1X/u0CwXsPGteZWyebJYLzgpPTyr6hgRoxiRCjFpLY
TEHBg8sjEoBg5oK9C9uuphg/OiXwt0XdKV8dUafvyRfFn+pdGhGGzN5x7v3vTO2pZeTlyVoPVo8D
lzrDtTc3aCeox+g9qdruVktb/kU5g5SamaeMrsDy47ZfZ9gre2nRzUB0UJlFkHfyiw3s+sBqkaWq
9McG7NYaJkP7Tz5tOKXB9+l4yOXabtNOLzVtMaEA4WFXkTfQIxsS6jzwg2BTonj2ONmqO0Wr7uEj
5kL3rdBXTX4IDTj0hWAizUgyj0zUbSjIpHMICcSoXVMp56Xd2m5s4hESmC6aLa57wGNJohXsakE1
f/jf+1EG4weEHZNSAPaApk7ds9OzqLZFSPAyobXa6NF7+28bXmDFVvhskQBLHYpEmffgJC3EWVOq
R+QPNUFN1hJrus8ISRDh28JFaCaAunhC9nG+qMidEjBy9JJVPwrUq84ErWrEG7tM0Nl5Q5zexjwo
MEBAbxRwO5BMvdUzSaMRkKk96UEs+hqC5jhVfSX9SntgG13/vsoUhB0MOtn1C2vzlrDlLtU/MC5/
Wrlkhg0JFwLZYiuhLYGKwruHXJMt1NZpWEDhgIX+qDx+aHa4l6cJuNA0cpYDzTKGnIFqIdvf4TAM
Fxzkt07ynnANQNE2Hs0Z0uDjisBFLUWoeRJXNco8d4XnF4rfPnfmIo0WDDEVdPgMh/Sjr0nZm8U1
bCGoz2aeTBNfi8WZrWn4crL/Dtc1FIc/mh9NHlcHsiv/HiCp4kEARRD12VlBOVoeJCzOL11WRzva
32AAmqsZCXdPW/qLvTFqVJp+4oXA45yC5vZlYu4wEy5YXNNxePV7njzVsn2RdZRIXSEZIgWYsV7a
dkO7F6LaMJ1bHFc3DrOfb6SBsxWps3NxI0+EaCqWewEiNy7RD4MAg4lRnyDW4QQgCNUYeu0olCQO
HdsM3ZpWYASO+Rb+evq+kJPNkMkbgwrKbgMOmGgTdHIza+GoAoCbKr6Qm6diN25cnkta42cQdqbX
Ozeg6ZICLpt9+uj82jiqpTC4dKW+A6pVXqy/5J/VnxoTfELuSBl7yPY37iKPWby1AoQ0cXG6IEqp
6KPyHIFxXrPzBafHacUi8ltOZuO6IJ1OC2RSjCXb/phDHpeqjhRPr1Zk3ir63x3B7HHGJR5GLi+m
fTCqCY6iDp1gUx61pWcCayosiUkNK3RFUmnYA29k8lMPEXu2s2k4Iz7PThYmGh1p3/xiBY5V7GZQ
2yeIWkHx7Q7FMtXizxZ6gIYrb1ophB6OV/jm6cOBAodaAP3sPoKOTiHETo/yDTzhLAyl4YmF38GI
02+CBJ1GlxraKHE3+jnPAwaBgFeZxJ5xP/kczM92nDFWhcIQiDj3VxdXyY3Iy4AaEt1NKZ/hwjSQ
4AeZiNcM9bu+IBeX+tggKu5lKh4AGsnpyDqm/p4wZLYWlei177FpybnSdtkG6WZdA8hmecVAfC/o
qvE99UBRd/1a00XUmex6MHTuLt3xGTM1Z2IeNtfxCEWnyi6vMcnhBa5duM2NiAAbrhKQhSYrn0YL
89f13Xjuz+BB8uG7qJsbYN1Ntmoy9TyxtZ7pKbVMbHlaPCq5kys+eARM3uJrp/Ophw5Pra91Q5mY
prhqk5zsqJgDaALcW3YGcweEYacsKxDq1UE3B6S5tebPgNv18u53m0ulnX6yzUKLGE8F5iLTczx3
OONaC4kRrelojgScYXrxotOWRyae6x8qxb5e3Kn5u5hQX+LuWtF5ixpEFlDXDXbUJTv2wigJod9G
BxrPNcg9ZagYfj940MYWlmpITexuvEM6E0h5uSOGxob/bmgw2Wz2L0mWlNUlbij/kNuA1qtClam7
syjILPzoFsi3YZ+BbE1KXEG5+YvUtEsPbRfMJaA9TPMK/BqUbOHFZh1szNujDjqL6X0bIjQA7PFC
vb5IoFWne6fgbrM2A4w4OTYdbgaIIBdIS/ErtZTJutbR0zonZK4o27kRurQzdNpLYyothPaS/YdF
X2mNfgbJ6IXoeKB7blftpQ9Gyp1KxztGYgnmcWr03LDiIGekAEAW1ztoougGebjVqm4X26DkaxkX
nZKhUeMTIV2JgbE7+AeDWfX+75MEo+hxdTxGj6RFdvxL/IyvxNAylfDW+zQH5hRqXi+T3Uyq/2SJ
18UhSyb++JyKxNJXXyKIpVxwbsjCDo0hRl8XbJLW7tMWcfsLxlLuuaZFeyXrLs2cjDstojWhEvdR
hb2cbZ7vuiQrdz2Tk/o9FpNYNQgFOiyrUlMKu8J9BE2dH1ePsAxRow0MmpA7BCXcL739ZoGjygTP
OKcdcgBifzR7rtogXlrPqZLEaBQXxQ41MHEEF3vfDUyalkLfgsLvUC++sKufSyupodQKtOXaDAvX
a3KY5z98rnR9ygKpON68+9iNbB/6WlqLWrD8YW9xJx7TVKv6u0ojltcQn+7hJy4Xg6QVftlmC6aJ
SS0diQzHPJPEyo1mCRFx8XXoqcTelFymFR1og+baaqvhRXOOyA8wsU3Ijwj4uEXS35qXDqhlFWag
WYjAR69xq4ZPfTfwZqzuqiUqX6nzS8XdOfDb/RbPDTEBnw3b3WHVmdXa2WuD5tbp3DukIYexnHGC
saA3wmDApoJS7DRsh0Pwe8NyCuCrhlfihI2pZtltCrSOK+mq69M720pIwTPiEAIvCJeg2C6oUL7B
Rs9U3oQ5rOgJHM1CixqHTBw/ChbqfOUEDxptfn3UdVSTZX+TlVMyp8WGu4PPNLRVJyOlCeRb0FRQ
qdaESPMRPaJkz0v35zyBIkUM3WTdjQ/z2nsvEo27ifa/3BbW3nstFTDCfAg263ntMe/XqTCtX2Bt
Q0s36aujH/714ZN832g/sAi4jP9wxiApU4IdifmqU0cZXSVtlnZ9BQP/zSJKNxfwRP5V9nhrPSDh
aEgfW85MHwobIdmo0+qCaP3S12Dz82/kMIjiw9RXnU2HzFv/dmAJ9eVLDXq/QiMFrmZgZ28yV30b
T0Q6FGCDKLkKv2SILKaeOzi+5Xl7GoU0KJOxUXsDOEVw9zi7ULdIJ2l3XTP7U/AfT3i2AyQGTCeJ
VSXdI6toSOO07FjcD3Ac51pfAAnaomLLig9DWxzvFewbFsjj+hW9Sec/NpukO/PBU5+ky0mwrwNz
PaLsoIT5Z4O9JqVEQ9i0sqUMwose8f9S9ylygkAHu4X0aA/ZiCghKh8U3J4r4GUYGzcWtMTjedwk
+2WkxfoBnciRdpzoZ8+OVE4VCaYGtZup3RAsZ3iBRjywpw/uAtXE5iSQ/M+FvmcSxQExN6o2upno
+SGh5fZz6qvHmXNvfdoOTu2fc5MPoxkeUaTw1FCblW03FjeEb+yoJRgTkfe0W1RCKZKSryz1HnhQ
Z0fzcAp5c+9Z5qq8tuRaXt9o+JBLZVLSA//qgxTnIuAtjHyqp5DH4GLYFGWjL6cQo30MCyPGMoOS
BpGxofkO1Q0iUBH4dWMlSYCcT8T0sE2l/hC2LFCLV674Z1bt5JyOLZL4N/G+nlS2hIPz3oy3BAod
KqXyjPpmmAjr7hYpFLI8/ddXCWtV7UJkmlav5OQCmUJZNrs2brfG5GsU4TnBTCJ/H+FalWDNWzqk
WhC61of+ouh7vxQtV7TX5f5r1ImOqq8P2emulXChPfDOMQVxM/FbUiNCw0HsrAZS0cGrVm0MICyF
1q4+CqfHSrrQsDj06lEtWuuMXr/CKHKn0uNaXwR39HGMDCMKK247kKhsA+5nILSemvOQllqYgeKp
LllU65PzZhYv6ecnb/eVt56aLNDynAZvCSBp2OmDnZF1N+sh3piVPzlW5VMqYhsRzVHGJpdi1BVo
6IdHRfGMFsL9q2KWGZLesBLZ4a5DLi7rPCW8kKd5wAhFQr5/F07Y/0buX/m6K7tkEQIcw/AsbAGb
jyoLAHWp2m7ab3mFTz16shjtskUKjL6BP7cDl2RMIoMmMdZ3Eg9GglfOnRgJMTCPUYoflHtU3mmf
BIUQNQEpb/8gC7EviqYHsxOqwpnv+25Gz3KXBWNtkQLI4nweo6v7qSmYhpqgd6GYuRestQxMJF/9
VhYCCbd3w9/1My5lri1ySl0BbmqXZOAvv/7akZbrwtpfc8gBZmtEaiF995p7x5c2cITsrFznuE+o
/x6DoVEa2xUUnsT2ZgkRxEQdPHs69lJJXXyxWotMkP2imZVVOWGY/T1mMo6h0EiWFoidhQCw6nYX
OGLJ8WZLJGcionUpLb5QjalTsqOEecvgXa7KmjxNoykNDY2CpECxlNWutYuVY2l4SAldCzo/Gx3e
IFd4MZTF6tZHeVYTCYrEYXL3J4ybDk63dOffJZfTnK6+mttu/PuiI7YwbGBvvVEwNgY/iARsSeMI
Ua8jHhTzHeE7hPPIb9OKfXzoMLMRLOzoTdNBqgKi22aXWOHP1QXLSk8GEcUI0wMGBnCsgE28/HPW
N52skctaFalb+lsWRm5eDHVokXCbk+7upAo4On/ACdILMEGMzclfPixyheO0kf18HGxEfOPdcF7s
CApk42vnjdT7g0bMBlPUt7ZMZqOzTqOo4rph9OOOyIIhCWpJ1vDdGPM0BvHT2ZOIvsiVArf+NMYw
RBkR6PM7+3INvemDoLLWQEAlKGflCSivZNJLKZ+XQ5PtxYSRKY50S6h63er82Bxrs6OOH6MEcKzt
rp32ijZOUGh1B41nJ2u+PyMYKZZQY65+XzQtl/JoJ2Ac2XfrU16cg01QJMNXyZCD/UaBdZxhvNuW
de3EK8KMjEUJvW/ALgNXvc9NUJgcxW+oimgJpHplm1OlN2/Q/3bfPeK60nZTMEz2l1I8XBDF2whG
UcJnHQWsyLPvOLUJZ3485SZKV4hioOW1wi8p2gl12zjsnJB6tj+YU/UAAmUay+dkQ3JhrfRLMoqz
N5guu1gGuKE2hJKSKfszQ319b3A4A9ZmgSCtGEAHBkwNNb6tuKE7+TQs1FYgKJQFdYZhKzRwRCd3
AxogkEifehHDWpSrzJAhxndJdRfyq0mYgg0izlCpjw4dV/ZbSV3a0IOFK00ZxqhL6eH+dsEFR0jY
zn09u4YSUDd8ApufxF7Z3apFOAPu3MhlIJRGMOBNeHrLx8h6IC1ZaEuXZiezwe6hi3woOZxgUcL9
W9iYmMr56tYyXMxjkNL5DuIO3ilcCPyjZYsnX/FH2CQMiNYaz4IogbxdtYFIvSacN0thi0AhGNUL
T3Z8W8H3ZdVxgTmDr+XTMw1+eA0uP1w9zy26relbmW/t++EZauPUQEtd8+1wXcKIcs/ujc0iyq3r
CaDhq86xWsxhWX6y7bJajba44A5Qm27WBLrOervPLNT9ZRBfdg7ibTHfEhxq9DFWwvjFeb9xp+44
71+NnUmHkJ83FoEiuM/5pQAdb1FfAzR0KMY5HQMDhMzE3P+CcjQR4NzipSwaOBXq4D/3nszvad/q
S2CfUjOgmpjJ7QMMAKx+QW/10pipQwyB32Hsyp6OepdVg2INHaImPpbo4FOu2f7GGycImjZLWwKW
6nAVrXBOnaz+zDKuolKVjFQghaGqQZLzRdwWfNdhF8YLD6G+1v0cIKJ6jvg5TCaNUwrDJcKEOfl9
KmEd0DrZNGH3Z1vbqeNZmPGdxduYqNXiy+ZSYOTfGINk2eZRBFj96gKzRVLN8IE1RztbGkOJI0tB
Ty2sbyqjexwWop6moE404Othb4pazZ+85sEaPXxD8ZBC2M9MVbNP+r6qO6g2uCS5WxaTSuz4QHcs
rZ+Ipv1ZTCrlr1S6x9P47AIf3M1lEuFPLYnw294FJv9e8wlOM0YAZ5msmPsM3kaq2KgHsLlOb2M8
ktunr9hnip14e42xOoDXUPlK7/tHB7omKXdIM9+xMh40oUQq51/sFKTK/VWt9An7qSQ3+3BVKaa7
dDn0NPbgLooc97/6ysjjpVEZHedFRZR/QaPALfY+VSFpmZ4rvf7HIqbK1+T6qtSNg31YtHTNqbi4
Vqel0yNUQzZFnQkurXR4r7amZFpVHk/JBcNUx1aYdAOjIaqZ2if66a6F1LLGoeF/Pq5QCJ9oB9j9
qEEQfA7TE2teHa6hYu+Gj3lhqdgEWkUWOShJlsvCLVdxrGgUcQnXouJDqNstqHDL92LAqqniYYax
/tYbmYoMcBH3AWrr08F2ZWj5Bu4YJn38icE+eppIF4E2351Jkltj+wq2C5vVg7hMelLGK6ws4IaG
b8/zegJ7mj8bv1UzV7xsp2bvr6B4+zIp5QCJnT/DbjC2Qj1Rlcp5KF4avnGma3p2vbDBbEwbefwb
LKsMQAvaH+1RBjwW6u6OWfh2bbnmVsU7lKT8gps66X4Fm73A8zrxUu3fjwvUmFK3jaD9I6Ge5+bq
hVY4Xl2Cyw0iJdz7MkMjLVdrjyp6OsGWdojXJUc7Dg1rcELCHu8/3Fub58RhtRkqAVyHbUnstFh3
Gow0d9MIDTADLTzmDBT+rfoB3HuVuigWdwTahdYJGY4wTAtoo+ccVaahQ8oE5OlOpcMtHlbZC1zW
/at0OfdxDSuyqwB0sgi3nok/UPbHvc6ZCW/10kx0BGdgB4zKUDZ4FUThHpym5QxzX61LEAJ8dV0r
E6vzqAYMc3ui3K3+zNbu6o34rRH9iOB+aHibCNYjREfVIw5eyD8myhsYjVHmUxqzE6ayydsI8rCo
vjr3iiBrwfuFbfT2IzOo9ls/aEtvP3wY6eiGyEmPTa2XayENRxjysG663SdODkYOBduNpI4ACKGV
pLVFG+ewRZGTBp14BeYiTnDOwjnmjD1X6u8HuHmmWhehJomck80PCKc76b/1MNsFF8vDywSazbVj
zIoPBxsk1b8NnpiRyMWjaVePkI8jMfrDfeCAWiYBxVHy462t+7ucjs/tvmkFP555ONuR4nqnhgcZ
hVf5aA70dXpeu7MKb0bq3SPIbI2z4QQ16YqVODaYVS0WTWFkV1SWrs1pCFxAL+9w1gSFlwtxpjez
gADYs2HuMmEKKUTn8U7hlG246EISCOndejGcarA8DIjpswV/S3YHjINK2SKz1Ycs0/pRdl9E0rCf
TxqofVFg30/kUqvFDZodMUW0SDyLECjl60kG287nh5kGr3+Su3ixRwprRiAqmbFhr2O57d+PaAqi
JuTJd2fgQiqCA8AkAgJOsDvC5MEjFhfv7o99XsXluEXP6rSBUn6ME4pSFQsgRvjnH4xTR2eBmZy3
dVI7W3p87g9tD4M82zD40HHzgXTT6Wi4sjcxrisJN0GB0Aplpw3YlBSqhSldwiH/N5bPUMOL25Kt
soOpy2PO0kMPBg/EIzwyuaHvHhiatRa/DfRLeE9kEyW6etdbq1hWRXBRSmFhoGJGU1uDFFTQyB6k
knqtAOJ7GvWZlC6TWqFrC5R2e507vsknpkTh5jI4mS02HatPlokIcgfbXvkPNI4rF2N6qVmu6P5v
DKYxcTZMFYsqMBggiGoXdv1y+FQa0wD4v2Skcctox8DMlUAmKE87iKh3qqBpn1DVyz+m8NnFU7lJ
iae9jv/7o0OgweKcvIbh8ZiT/QCvyyovBwtVwuMszalc8cDi24k5LvdBWSi1EwVrxJqX6+YQs5Jn
1+4seYpx96/ZvRxZMT5DzikyBtrmNcoTq2jefjqSZV0F9X6IJtF52EX0X+L9usyIopB9smSmrGV0
xiQr7Tjp4yfq4UyRXmHoh6IPuv7pT5nEz1i2P/hjl3L+Md5OfxmW4rGNGW56P1onINLpsBx8WV4g
L1FpR+NSmMAYFZgV4s5Q1FQjH2uVVJ0PJPVe/a3Pu6xK+/s+vymegOVHBik+nZdgNuS/dY+RfEcI
Way0JTuN1KM/kPpmBSU07RIeqJWTqbdDNYp2+r5YJA4Q3is15bFVbfDRc8mb+g+dl7XqowUR5pUv
zsjTmbzV/Zs3wnAQeBlZSRZWQ8bBCYuY/zqI/fe1SSwnVyMAvPSAnPKgsb4W1s+e8sTf1sCMqdei
/Fm3k/9INH4ZUwTYwRggMb4YVQzSvq6a2t/RHCDfT+AdrDHlS7vbqKp0WWjqwfZw3/A8BA9401zD
M5/ZgsdqEyAvkle5iAN02mje8KvFiAQuDBRExJBxnwZPT60ZxYcPqk5+F5PBTpf0HRCe6/2amOpp
+MFJnTV5KYRg/mW/KdZfFurt63gxQtakXugGIsPQV3Q3eJfvEk8W4cDXuuiS9GEC73fzoivEXz0a
1wUwaTxZTTleUlHWyvYmAm+rm9uStsOTs5QLys0a5PBFHT9bbOiIrjakM9QMrha58phYoCgcS9NG
owE7IrT4xNb6eo+7yzcH+p2sg5MZUPUyTIIyuQTh/7DuvEPDMmXxR2FcnnjB5NX3T+YRUV2vBblb
gTi3i6nn7jn3lWox7EJWWKCIEnEL1qXndySAapUwJ8Ts4Q3H9ab+N5oVBl9+McTYhTC9VNx+FLT6
Xglb1TOqHHpb0f/srA7bmL0gD0SnwDgipE5fQMPCxSnAKCUYM35NoIYOTLPYqe0pkIO7C9rEVtTI
VznenGyG+mDOCYv7+Ncg34xK6hn1Hr+VYkCR2JABF3ZdLVsQd1Jsx6r4vlhUDsL5vD/L4YH16U7+
Fc6jsYxFt9FmXi0yH7l/D6WXq5xTHssdGdBwU/A76o1U3S5u9xNfzADMh4MzJ7rk1xOQSWXF01bv
QZGwzH9H/QF3K0nUJDP08orJbuwXZLM+qbZ7OeyharXgZZA+skDOEFCp7wzgSdBplYAsEAaXjl21
H00HewkgU6NDua8g/ozM+5BhdEFDCMfh5PUNUw5VrnIrXQ0t3aokMrofoA4Bi1+0NRLay0EQbN2a
XV9z63TRc0k27b74nqztLRfCVH/3XxPCDGqd2Amr5WxmlzzfauW3lMik9GEI1pEcwaw7eFCgp6Kp
lLT/8U/SRVtm1n2SKRZZXuRS1eDRBBMhcIvcPNCr2nc2ZfwGiZ3mAYoprEOza2CcNXnUZrpcYnz9
RZSshalfchNf5A7ifoYkI1IIub3WDAAYh2darf2RCFFxH/B/9jyGLHRml/t7hhpX3EG+a5PBF4Sh
ZflGZRdBKGs8Pa7WKXZqgsWXVOqCHdSG7okgMcwR8NtAEQPsq3TU6V815aQtRdVAbpUaueIepXBT
OLnWml1yTAqhtnMOkM0BlqKuo4rc1YCKDliVdHY/ib14iMnVjgYsdfjEdlSPSKsdxs/awGYxnqDQ
gYliIAW+5DZVgPRC8wnvIY9jch5hzumWZQgbOrVGcvEXGzf2Qh85sMgBY8taBKXRh3H7ZkYpR7jC
SDwQM1DtB5ZcMo2phX8VxC4AZnXvfw5EobOThwG/1ULd69J9qsr49IpVSdf5BErH2ayYRnW9jxFM
aGzEU1ZxVxZ+RkswJtCRZH+mTFl1CvOj++qum4jsU/YcnEs8F9b6C114dZiff0cn0DR1QqXyDyHI
52ZYCgrDrUGY4jGNX+sXD0dcfgoLObyckuPDLGsivTB2H9Y+vpSmLQ+JEuON2A1Re2fF6PmOh2YC
OyNN7Rh/5fqy5WgG7ue1FjfNbA+yAXdIff5pRYGCH3R5aV2bVHjzbJ6Jh3RHkKsSS/mVvlL/U8zP
fxAedV3SlBeqINXEEE+oh1wS3oTKyOC1GMLKGuonf+bhxCtEX2YwawUsx1nKOTXi2QV0SR1u98Un
UAgXGnfGNvER+tZJca9RyQfBfX7ytl4w+MCKONnKwMKIIjluM2+41Ux3De9N2UqT0+Iiis5g2NDr
GQEOvJyvfzBGa9UW+mEl29lJFRtqymbClytLdnixwO56Dvv+fAHTLjBU8psEnblM2n4kuY7a4M9O
t9nfQht1S1SlHgOocA3UM/hn7kojRbBBJ6C7Lwgs8RnSxc/DwZ1QUN5kp/7SXTyk4MYrJqLXAHjQ
hzxRc9o3XVRq5ru9kKuUR53Sbw9HIS1KQn4ZmRWbiYy1gmeuxGaGhlJJZ43Suf/vCqkl3FRxyNTB
IyLqxAbAS6nk2+noYP7LySpxN0nwXTRmFkNE8f62mdhL5X7ITYmfBLPyk2CcsXZ58R9SC6l82VM8
kw3sXPTCqTZow3pRX9+MOwzRl1dKPRTT/8ZdGji9Anqr1j9Kpjtsxg4NPnls1NNnoGl0aUI5O56U
xirtR/dzMDefIcjEPAHqPr+z0E4GurUmAG37PoqG/gMtCbWV/9n9x0kNEWjofEdLCarh0aQL2+VJ
/5QwquARp002XoqW5jC4TJXu2alf80BzyJ2rhvGK5XIDBN5Rji9oOY8RkYG7sj2Q4qZpHfGbXePn
6Q8BqwFlHtUSXTU9vl699Z/GeFKqYjN/NrO6YJXNB29dRBg9DxeE2QeIdamQCVdQ5GcKwA2S92go
qiesMIGD0TqQToBjHupDuyzfKMGscJUI9c9ARtRKFA3u+j8BZ4T2ldwFh5jHpk1hq6YNcUJsSnk5
ee67B3Rq9rWTVtM9HUxO3dJZY9M74y6VNLJWh2oSyoWWuBWk0fg89pKzAAPzyqYJlPCVBoGHU+fd
D2LaxFZAJIG33RNrLr15qdSUAXvBWoljh2oSbefNbqzSMGcRsKJWEhr8SzzEOJVP+pXQF+BD2xDb
SzPy5p7sEAq5bxyRUlabxQkSQ+jXp8RyIzfCd3wk3ricgKw3jPlasA6I3xjjM5UDzkcxKfwpw0gT
oigM6Z+p+cS0802ZCECJWLOcxQnaG151tqLTA+lnc18dxXHmEiWyq8Dp4IyqbVGhklxqyeahgwqk
/UzFlUUdCvLwpXbZgifWnDlqhYcd7w87W/o8xP/NwzOl40Rmjsk4j9KPF80qSww8B55HDNl/is/y
j+/SnPetlXVt37/YXTUfjC39fEs1cguijFmD8jNQPc8mQ7+odxrYQFFruB7WKhLZKA+uWcZ5lI57
ap8tGcYsKK3C7OnhLTvUyK6Otq6nABxnGcVy8FshptKGcgWbhq1hRLkDyUanZmeVHoUnd6JORDf+
18HGxy7Lvcm5IsYQxogWR7W8UgcjU7dfiullkbDINZ6ayyrm92h6y0hkp5O8qmnrtwdTfIbXRJX+
rrIKvPrnw7L02r20A/JOwN4Pq5ADZCcGIUq0dker+o1lgGB80uIErEgwZgSAifMbfdQaw/IFHKgI
u8u0BapJq4Bn2Q2UAylxLE8yCHi/sauseDlA/bGe9k9QVCrLAE6oezdgQ22sFIMPJUG3oiXCrtnI
DQWaYZJTM5vTqsTUgK0hvIIKHQiom2oCUjOrDL1+iE5pPshN5ugQHV1+rGX6KJ+IyTeLVrC7xrAL
L6/QnIa17e/VFFmtKEb703iKWX53eq9LmoSzQO7XUy+1OAzS5im+bxdzHG/QuD4uJfUz1NIq6kJ/
mqoiJM3gFj69TfaGMe8l8l3rclHHOPTW5S73HME6EYcxNTdTJamfgDtA4R8QPWMsP7tqMZG3G8q3
YuoffWgQkC3iig6Bawzu4xBRZBKfQ2suHtMge4Rvo23bT+85aw0xyzIFZD2mCtRkbS8ZjMp7w2cf
hLo4GDTPNNU0Trj7MWV3A1STM5gnprBK5bg2AzYNsIbdLuPpsIlJm2yiSxkmv/LgjiBQga/hpJ1b
dODIUtWji0uOlMRB8aSxRY2OOqKIDiFAIlpzFor54yUrsaV1yVafU9mUax5JK9z/457efSidBcWR
A6U22pR1NmcnieDdHMwanPy8JEz+YffB4XkI0ts3IV1J9GOySXEtqLh891cXJInJFqXa7C2P/pK6
f78nr18TT5GPXqvFns+JOeP2pMClQW3PffxOAJ7hVlLxbm8ROQ8qCW5UQCyyBbcbSx1kZmimFMUv
A9gP5ocJ6lzNYxh0nmn3W7j9F7atqhSqc95c7dAYxMo/ONM6Lq1NHdTK/qtDixajB/qWpeUcLZBO
4dpg/ljnHZz2gahg3fB1QM2QfYaV/adEOk8tdO20bCtT+Ctb1Bc3MQODauxbNZxhl86FMbp5SvHw
k2xmxtdmBbct8P+T7d2m5rtdxuj3ogXdClu0V2jUN8jYcrUNjQdrfwQ3NqC7i68s1qa0xe/SOngG
rGqmEZms97C/3UT/em85jQyhEOOZqqwX3rHWEKrG6TciBBUXr3EdYMfO9rVXhMlHTxH1yO1kv+9q
4d1Tn2cJ7L/prDiqnA18R101JAp1KAHYk/BwuUdPgv/1zR6rNEaLGf3TITrh8kt0Yl4IYreFIkAd
wbRD+jJzvCoNz9afn50F22rhD1JZiwUqs8w1lEi3AAzPz5o7aawOFFbs5h3wn5DfzfWgMYshA75C
cbG6tAkQQzi6YAtWgdPcf2jcCIBEtbtdR8Zf8xSVxOnQh+HB7mCQm+el/TD2BNzHfKkBa4LrUNNW
PqFPyDdcmgMho3z/f0/rYjy24vjqVm7fcpDAJg+OKTFkFyfx166GZOZESXOXf91sk8muyw69gvRT
vm/hpsE5RJovdyjiMxStAPcuYTCC6CfBPGyGvTdpgEIUzGy8/r9mCNwRAuYpE3cWUj/wKf35UCbj
MAeNLVHK/Fm8t4SbSCWD+1XplRZc0PfexsNJq5WXLEMm664/hoAQfpsXa8Gd26FKPR44zFKoLgMg
ZZ/3goxXFuVTzIXfDMvZyRytqzGN96/nH6LKsHTaPF+fgmYvwZdwsSXooAIwpfwq9Cg1q6Jz3xlV
YhVL7ZknfP3VUfJt9nJKp+VZitYtqUGfiwd2smxmpw8Fga0MMSwxcqzVT6hL4TOPy9Ynh98XToGs
puZp+bfpHYPwXKWZPWfgPWLK/MuCE5SvmQT0tyAH0KexQgHepoxP5cqYIOsmfVO6c/8XS795GCAT
gGV+xp7IFuSrcpnJM6Kovv1diZcWdKO9OEF9vKABpG0eVYAmHHPK/7SnsNJKj2EOj+yQodurJDzP
QODzNnbQHzMEmOxBEdVmZ0rcDNIN362855a2IZYUAa3R43hahs9AeQ2Ohx5hjAIck6DJs9UaxuEs
B5lm1wqKKEjOEtXnsLDBRzayWYO1luHKVT6XphGllSLNxXlNbw5BO9qV8anW94JNTg+vSpSVZrFF
b8E27kjdsACGZYeetz1ssOpAc0FS0WSDh4T+21kXYVJt+xqpeAIvfYXSA9D2dD4NeJgTEIy0hfvH
828XMFmiFk/th2xhNSma5z73TnWLtUszafQHCSwMoHVWtLUDl5tDR/AuJ32dTQLa8s+rye70OidU
BJHmivLbpaXWdcxIo4X6IUm4Sxn8J6BokbhoijLlMSyofH6k7M3kdHwtynC+RgYr0+kBes0ZSVWj
HXDFE1ASXPg5IhkvI81ViMyJ9ArBuTBF5kILl0djAiZyQGkeAniMAs5an0MAVynk9MxJz8h9nGMw
mbpAibGRa+jJ4BrIdIsLxxgzrNSQUWXK8BedVcUVvO59yoOflA21cundEsZWyS6oe+T/pPztG0U4
gLbKr6u/87KABVe3Dp6LAx0cyfCPWLmQwQfkW3sntR1vU+QBt6odt7lADOb21Id9wCTqkNDDUXJm
HofwtVSX7bCSGyDln2lDKpjDVuzS+KRF9Pm3D3i+z3L+tcDAkGE7mk5ETuQct2HtN+fHiiBRSAW7
fHj1p1H7OkiPYrmo3McQFYtpXTyoX+iwO+KY/4gvUWpRmC/u+5B5hABkm+oKVCykABfh8/g4KBoT
fKfp52cyTtBJIsRl0cDnrh9qrh222kxI1BAXjYEPWGd1tQL9VdLd4Uq/m0OJtoyAW+qk+aeFXsCb
1Vc9Lyv9m9QUuaKcfU5VzQxV7NKd6NurrTl6WlAW1mMh8bD1rbrcQpB+ugSAtUJhEXUpfLT6vB9z
Pw4r0G4eR4wTaW91d5CHSNxw/9Bx7O9ZYodyHakMDXTfkuz1nHfMEWe5euPTFZLY8z//aGo1jWdT
WVUBPaKFlAL1uDEAGLxLv0AIctZwRHF7zykjT/XkbUX6EtEmalKG+AKcBhClZl/pB9GxO0wyRpIc
9y04Ww0XPSIui4CCkYfLXm6dpkrBC0udUcrlizMvuurWn0wuDd8ekTIw4Jt9bigJMCaR32CqFrXD
5RQ59rBh7Z62mVIX2ObTRT8JeQIIUywBBuWSFCgbVx88s6cbtt0NCK+fbQ96NoujlJI64AqoCv2o
nv9UTE31HJLMp4WHoQ1bAnOaCa4BmgII4TALEs50/TAi2bvYuhCNsA5DXzX0k1EbjZjkzNP1MadM
3DntPGXpde+MF+7gJG/yuDGcxUE2GHslG1iZSUdAiBc675eM70yCIRTHx9HuQ1szln98p4H06vlO
E4iyUvyKjy5qIHTMErW5Sg2obiSzB5aTVBT/XR88s5c2RXC8HFGMZ/u3bBjcEZ8VPM7Y+i7zwJ4+
M8OH/QdAHCO0OIMdMGNo+d24c7AHAAoWVU6LUvWKGQjANtge51kd4le1ACkVGU4MbmQlGlyW6jbY
1cHq0aczNL1TMXSVl3fkraxdVHddny7Fw+vPAJbUVc4UnznbbsWL46ZKTleXuLP1jSHEKPJfK7vj
Xkgszyff23McZuJylE99sinF9CYbn+cM1eAluJf4+zq1SuaehfONbLd1h5VoSE6klLyWAa/EkkTS
p9UAMMsjIeJ7RA5+nkFPqLA9j/GdxM5Cpw1GB++tuzT/p2HjhSL8uTi3lFKB2RPkewOCmDmljSQr
JTASTyVgVQ2c9KeZNhwEqqS9trWL/Y+bLyb0ulzBFLXagoTm8EcyeSfzWjrYtFeE6ZbZD3tVNKjU
atpsGRhU0keWeAvrgYr9wl+6XldqPIvOnG+fn6S+Jz9fCMz59CVYjc24+kdnBN6W2J2IeNxftZVM
uldIwVho2yKGlBSdd6QfzDwNjsrE9hSHXkXi6pfOWvjCsKzWosdPpYZfrhG7qffVAoitiMJMeQwI
+cIpoIfr8B8RYg5X2yUOZfO/1BVdQvZRn/l8sChEnCugvgypp44URJ2pS7kYnpDkEdvfMUu8DVvj
WobKWpF6/MJ5AXHrXxnZRQR3ttH6i7CdiHCUp58i4isrfzTjsR5CUOBO7Ued/PNpwlRUdNVgB1L7
OMi4TgM5jqq4vat9/mVNOyP7x/JWTJdw3IaBcIhiOzhCeG3LzvdRIQdJ4pfu/7CRaAZgU8P2wjO5
joA2TNsa+DcJuIgmiudDOwAOLOifWkXx3bc6NDY/u1kp2Vgx/gjWeuszmH8EBq7N8umeqVYbVJN6
yvhAr/+b2Z0kkOX4/6C3HWGbHsel4yZ24Y6LAysAeRx5cfNuqjPfQIlyThnLL+/Xuw55lRnc4x0y
hO0dphRpFjIFNVufu8RizAhVHIPoPvb+r/f2TH9rP1MFLZz7/xeiq69wQQXjXZcvQ1ufzPTlBe55
zwl9nRa9i+0jrxyaXGp2wi37PBZ2WtcMfHhObiXg7xzF8OnH6oaf9d9rN8dffCfY0Sts490AOzXf
DSrhxLSqKOsPA6M9wAM7Rvb3DzqxiEnIiwfMQTTXeX0FmACkUhRyMSuQhLpQgPYXDkIGqPbWGpeJ
7zWM9+DvJh2ZiLrkl3KfKXexulF8akqb4ymMaBkc9cDflEA/TnitVjsY+4GR+Wfdzmn2205uuuLO
4ROzgB3DDShWiTUyypDT9vKtLDQtx1Wte2vR5YEI9zWFqLpZQimJG/x21fh2BNQ6V82DRGSEYgfn
XSvfYGDG9T0MBpYG+ozPaaHFPwcJesbi10dQjC6Z+mISFDEOkiMZwSF60BRpDOJvtkR0LbWqrbgM
WizTErALGFCABG5aL7MTIDbQcAzAyOT4j2+lk7idDNJdHGAx6W3/M/jcoBKRRd5S4ORYmNh5YVNp
kROTPy2dP0n52g2pPQ7cNo8BKuZgWNgqLr43t1XAZZK3kDYyhT+y+fC1CCyG1io3EUypfrZcPHbX
9GnP3QDtt1mrtI742ErBoYaUGvi4+ZjBqppGfQFP1F0LgJzdGIpsUbxXeQoaD/lH1tOyXPptfuIv
Kxwf7YWw6UgOaCJmeSW5r4uYpiPB/+voEOPq7x0nzJHtdjev7NFe9al6nxA9Y+ArlMmD31/Gi0QF
1NQlXkQ5vIF4kg3P4kXVb/JWZyfsJjdCn4jXqzzmzjhx7nAabWbS59MTeVi5/8XLhzkmU0wX/YW2
MUR6leORiyIemHh2vNoZ37pD4abguz2nDisoyhfs0H44wsLDUkecpsFZbbtv/4MvRssLijsLdJe1
jLyrXmavkfX08uKkI1pRxVhn4iG64MsXBKtRUujigI/piDCAcPr85x3VcKErUwzTIQczXc7AxrZB
eJocn/iRGKHvSl8HmYv9HEd59rzZ+HMcnfna4jmmH5AaVniSNhkSSSL4sADTEc0V/faRIoY7ddsx
FNlzU+JD9uL/36X0tEDyRj17+XVJYRJzkf/XLmhTqMbgo7Spd4VA0092M0troAeeKik6x4gTOgOD
VVv3a2d/1JGJlk3r6yqPUKWZPPgm8xvein4Vb9ke17YvxAg1QJlYobjlFZqRQWbknfwYwK7G0g3T
o5d9p9LeU2AWWXNcEcsfcgWT2xf6oftOotPpgG3RHCXTNpuNa74fhgOrpPuDf8Ep/EVVINOE/G9T
NqI7JcLRG1IH84T5k9/sFdOMC30wyk3odCWOywVbb2VNvkz6zwi1fsr5zAXMbiD+P4K/1DJszUKN
M9ffSU7nEwfOglRfbL3cDgQVN5o7PwPsqICKH6FVIGNBkyUa7VaeH5hIPtrEBJWJw4zKHpOfF4Rx
w5u/82Fy21AWJaW3sKpskNhZtHnbEQv8m6JMseteObmcGRSqwtf4StUGk+suRaC8o0KwlNrNFnFo
E/ou80FwnoZ1i4Ct4NQ/BKIF5at9YaHdLXWclP4ZqfQwn1cmHqKVpDYgE0JJKGUnevfx/kyELC6l
FGTY/3RhdLKQ/M40AYNF0FoRbtub/9/t0X6E2XFiPXJkWdhQsRtZLkgKRDRrEiVS0tRiJejedVUC
VHELs/17cSWJXS4Hsa7FMkrshYqM2oAGwOl+hsRgV4C6EPMNIAl0xk2HybN9T3d5iZpTMftc6TDJ
+UhcYJWV7mhgNt7I9XhEqvwgMRDpxiG+OlvyWEvKhvqsbnMniEvzdrebNUWZLdZkJ2WYQZnwKqsF
tsJ4szgv2t8cgS1GQfvcbrnlOI6LtuMo1hhQZGkWZV93AG8vXuxq3WGGKNQkVAwpXvOhGYT23QSj
FzH7IohWLfNiueNL1W3Zfp7IBxBHgKcUOkgRt/GtHrn8Wx4diTokXsDMb1r5G2Ep46nOJoFtFtfc
yonqU5JytP/hI4/GmSrGtDUI64SNCrmWWo7E3QeBAWK9W99B8IvFIKiRrC7ZdZ5Dln0D2NYg24eD
wlQ7saWqfHvF9Vmmtg7bDktYOneTjV1ZiPDhAdN+lLKx08SXjta9oo4wVgv8f9NUiAPYDOZrt4vx
6QkfFHazERYKwmMqTVOEsLtYcnYWGhhlpRn946xHUMou7Xz10hNKWWPnRqZG8XDdFM2amyIGeUnK
ZEyr1mUdIb3aUT+OVGGHaKlEQ+c7sUNR2d49MjgAWn1s8B+S+OIeQI8awegBsMTL8LG3JUAzO02y
D56JyKzOM0RWavvjQ6er3I/tQ/N57wUFGL7tXGHlSVIJSiR3V9Y8ViB0qVQ74jX7WaWXK48QqUAu
akfllEGbs5BfndJOYr+fYCc1kZl61dLPL2+HeDLFyqjFKm6BMNcyutwrPqdH4rz5/5OPvhcRSUqO
LmFNhAEMVSzHCnR08F3l+GmZvdIkXjEhpfgNzK6yplJMlmays5kuV3ufqr3+1vpCQasPz7ami54l
kU6wbUtrMuCPAh6SRokIFhDhyZI9UgPKXUe8jnTJFtoTRFyYOGqC2Zu252Bdfs38gOnbFFFHB1J3
PHBJwjb9lQ8KPM25XAP8oaLO7xcTiqG54jUpw/OsHKKOjlcucTL9hEY9dx8WHaGJM0xW1qOETXhw
Z0uffzZzCLLsY2yL0xibQrfJapC/KcsFzeMLGJQa0BWbKUDXutRnS0mFG4J9oqmE6FPZPuyc813V
hE/afWzM0spJPNmtCUrTLEnud+cy/Wyl6rFgY49SWFW/swXa34n2ybUODjHIwyfw4uatU/tIv0L2
3rKTzIg02Lqb4JWaSC131PAuIJPsYzS2Xg31ApxfD/EXQDPAcndcWEioWG9jvlshNKrqwJGLwfOR
LJONrtwZMxUVGfT0WE9355DsYkwOO3a7ElpmeCJ+cCehTAK7YGzlUl1YlFobqZiQAFuPVpneUXGd
3QKN60NmSrePs9Et+/sfgut9D6f6rDatmVqdOe3NWc4BS6YjmSlH0nMEilhLOeVDyiVJ8cpBB/2k
+3h6vxTgt2YjWa9xVj4zm0Z7/g8LIxpvwe31uXUPQKjxJUfSNI0EnQ3NUPn7oeR4fUhpUh7gmr2N
r4oTdUnz45nmVyD/yBhcF7pK5q5jngIa5HR8x/CPMaU2bSSWZwQ+NCg83dXae7Vxkm5lflmvixor
xPsyfjFhnqP8O8POoE3ZNBXaKQJ6dVbQtGTfrhBoyPdv7r7anntR84bjcJ2nQK6aj3Zvd0j0mll7
asmDosa/ihDVbDlLxYqTxg20DNefn8PWN/3em5QFyV+/wJZuZ0y5fxigihlIE3d6HfMr4+zurVtB
/FmqGvMuwGgvQ+pfHwbipwDk9yPM08DiLwKrp+d6+JAxzFXadkvzwy71lc4MJ+muQW/OWFgdRg+P
G36FzcyCjIIw39oyGRKyQNN9e8cNoswJKKqDBJQfC1iN6f7XG6TLvMqzEviclYa5Mw8BV90eL84I
XtlLu+AuxlfOqaxPEhZsmhequ5cVDY3U3TgfIV66JDZIva9YR7ghTDZVUDU2b1otsVF0WWqAxpV7
Y7bpTrXR69d7NGTzdPNcgqdvurp24KArZxErmAQGb32iQR/J9u67oUXuah3F7QU9fnMtruMByn19
vxRogbD4vmx2WNHIWd2RmoCEB/yHOWq3QG/3nNwyCYVXV7iLqDpfn329yoqEUqqNDtqhffwsvOmD
RPzcBe2xr8G6clXETb3pgyIjV288W/FQiYPQAauDoT+i4yJ6oICN6P6QaMFFpoTTXdiML4t6FS0n
ksX1/CELWZG7Tw8KwebOWYeG5WQM3ohktcWxBbU7nDxes7zNnaO0ldlGus5GUm7Rju5t5wnhbmDi
Ck38RG/uCOuyT7cKMUF33UvqYS9znFQU4KVfhWNXVh9Gay3oaDrMHh+SYuPhrwgXboSQtdF6T2Ew
IZRbnrpq7uc0QlYIPvS+n4ncdZtWKXvpc0YM1PLBqxVfBGjUayGmkuW6V8Dydmmrppblek8R35Jg
W/Y0zM/yWSQL0HsvZ+JxSm39120/LzDfmGXLj8n9u05OMELIRUtk259TrD55pND2Y8DDFdal+L5+
1sW8AUx2cwdAcASQTiRzK5yXqJFURRXn6zBLnkUWa1GXUm7X8DBfiDCVv8oXjyb1Bv8eW1hT6aFa
imMeX/kLE2S2jLolcPpmPQxDedP+ovjYG3Qk73aKrM5Do/XXNiCBc8Nu/odLzEp84mI/DCxJ5XkA
OtrwSEXpl1xo/9hfOMg1G+ek0qT0c+hTE3yp1M+w+vsL2RKKA4r1RVbO56C1XPjNYVNhWN45EChM
lGBgPKCQ3SVR/kxcsDLmop1Rd4Yjv+fQpUZ8MieV/XKV1M/mTIx7LGxCl23L9yLwp3vDvC5D2cK7
sC3B7XTcgN0wrYxrfgyALHIqlC9he+6rcFDzqi1oi35sC/IA3nlBntQD2EUsMrh8jodrkaqNu9aP
Ej0F87ZfMVQIy2Q0pB0BqcgAEEb4DsMN0m6aGtuE/mlDJaHTOqqxEDtcktuLnESmyb4lT06hRqGU
oI6SfZAKl1zh5rlgIrwNl/qkdKbciXkkywNJM9vU73An1tqh/l1P3JqkfTi20tEyADnC1VGM/Bkg
14e6owHiS35iusL6SX/OZAdc/KZxNwdRAopvhr0/vHXsD20cdHGb66215T3cmXYF8W6PmbHdWKv1
2predj9qeyIFBuQXH+fXUCRXBv5gvnar4q7ElXcZUxPUkBwwOOFysZaviqpnYtD57eaLVJzdOHNB
koML1CJUezmqXh2gJqHYNFKxXf1JILb944GxDL2iuI7jbYn7B8HlThXvX2kDAqTUb6OxwHv7dmTt
9/r1lYbAsKpBYmGFNU1z87GBeXKRQmdwptjlIls3ssas7DYuVcTLpSDWnOkSy1Z5v4b3rB8J/aIA
er9yhlwFXeI7PhW763duMRHxkva+ZYNJbhMpNkiQh2z7sOTpg0xdqtAYbDkTzWlJjXW8ZT9/MXEf
d9iEXL7g62SiMnp3RvKynwWDrZMr29DqlMSL6nATyPWg8FrYNrzGW+tNq44GnMVLAPqzXJg4j4SP
1GOwMYA4GW0O6aM4/Z1jP4pxj9fLHSZF6/xaTfmnoCjNtSIGjpy/q3etji4X0CtHK7WJ2dN97u12
0oqJj+0ggdP9J9fR904Wj5zanGREyFbWblmrCufXHjzha+EKkaTzEiSQP3/kjjscUC3WPv3Hs8T3
RgAmr1ylVVLXkA3L/X16Rav8D33TmeqP0FPlpvVrBr9Dux3JhK5kHVNjQFlHGH5dPkp1ssRXNC6U
oSX0qCK6wMBFiMLzcG608YZifMA4a7aMuMahhoAGltPOpAeTEBnz0pBqoh6Jxvr19kg00LewP92D
k/sBgYBDSKMXVPJ8C6+mn+VzH2i0ERDn4qC13t+fCjv9KLqceruvqkfnR5e5WIx9GUJjcpe4bUNy
n7ApRIbS6N6nLtWvHvLmn/4i50xIqbWYp2CHN70b4miS0oOs4zP1lm6Kf6G85i5cghPO1jGbChfm
5vrnTYwNubTxsd+ckdaCeaFgkwDLNIIhn/QF1+OmG30IM7AyxZxJjql1QrifpVno1ZpihYjwK+uw
6Kzig6IpVIpgZH9Ae9kuvMSvmqDj0AsKeCIWxqjikDN2TJpyCt16tyYb6DYv9GobRvUU5oHwtNsF
i6kcSZ37aBWJELUs2OIlRxGHCfS5OpmDXGYfSQKncnLX3+K5B92ayi9quq+p2zRwxzAUV7HTgonb
MxXEsBhqanmHJCs7OOvyuKBQFTKTRQkOJSmrPxPoj/reJK8Hsnu3376FBEt/ez5dmYjcarwVwEPg
EA3yQW3BRoZRG5fMHkco9twAiQLxuMwEhR/NPK/ZzzE/2Q4xBSl2jWCet3MIuJXeNrFaMwF/vUS/
PolhalVhUB0uL2y8XABvf0nKInTTiXjobeujBFJSSxT3bjMP6uIhsNF8rblxLgKnKm5bI4pNxaDX
h2H6HbhbQzxB6L0XZj7bJ2U0coEZNQAkJah7niaba16kkQQLxaEqmaPe15HfO9uX7knstciuhm10
UsG8f3RcsCtW13VkJPXqZc3nls6qucB7kCmlUJRKg9hBc370slOye1N1Zm4jb5jPlwJxJnhy6t3B
ZFA2HSyZ5cTMtYwiriBNfQ0jmW13YzMmVbQEVquzbOP4DjTePP1wgJGivz5Wz4MicXGCpEmJK5om
FnP1tQB2yTkcUzn8jK34Ln88iedCiBcDQD2q0DC0hOHJQ12vUvW+CpT6gus2kEAtLuax0IQuOkDW
g5XFVpohX5Qp446+aNfvdms5csAc1e3D5HlbA2zvu0bwMUYHs7N3fUlWDti2ujHqKu1Wzr9okLcl
2soWg1AQ5C5l+368zh8PPev/CKPn7+1Ny2kB6wJYTs5ah2FAkS7OD+0XuGO8x7jnv4+XbpxClILG
0t4j3+qSzpfpvuV94hie+yfkdyg3P8XBLtUYULUcJ0NhVAEH0c8WCmrzZuoeyCii0lw4yzUn+P3y
eWac3+iwZ1MkFf6PmAooPEApUeKKQc0nqh7czCrX5A8DWcJKn8pX5omL8iTGmg0WPfJV5ldp66WN
8+1vRH9mpZmAd78BQbtcOYXxD3/g0EyMWzD6ldWNSllzyLfHOyzkctBqoeYWW3BW2Va3C04MLguC
e1qpamuDCk4ykUUuZ6sxyD3xmK2glLr5GwqUbRJuW6tClK3Yn1t9h+eKBhc1Ss9sYyaoLpdTXtuz
JVUGUu+8HLAtvFYsXfKuV7OdU0tArhGxzVWohCl0/iItolKKgU9+gWEs/QwGllWJTReulRvEjh59
Fz01bznB0oQ+tfrBr3YhA8axwxjDB+wXoOIbI9z71ExxKce/CscFAPxlkQ+uOMLLVa3bcCJxG9Ow
nRizABjyF35yOVmnTQK2BwEW7hCXy34D6Qs53XzVhUstYQQ5GEbcBzmN5ZUdg17/EQjyzhHjygMe
mLRuRDoRNMDG/xSEiEQ+K9i3IcUpX2oZIEvoEETIwqTzlsFs5lyuLS1fVBdhOE9VN+P7qBykzp2w
ZzFvnlWuoLcp6g6CNU0nP8FnqcauBrsgkSVIQR6QU7eYYC+8m3uHiWxQO9CUZeUSoYszpe8WQ/IT
GyvHkifNsDofrUuvyOhhiLvQKweEOY9LdlCTvYk7RkDawmJnPiKxomLTPGPdo3FClyiXe3wsb9wS
bfTlxtNgJ20X9n7n4bSwblWUSaVhjyGJzSVQQX1UH79M5yoHwEBUDGUIJWGf5hiU5l60XWykpYEv
UqkVGaMkCkKLILRPsv7qs3FYh+GN2bmr0EO7x4yCSWf2ym0bbRvz4ZTxzhnH0uBYJUvUBzKH3Z0s
KfKQzLLRU2fUhwS0KHxpJiVIuSWt991bOt14FoF4+YMU/VSXvctCHAwyeH7krw6AvnqBhZJLsjze
e67bcbsn4bWst1NqZFNJ/kI30pgmAzk73Tj1gpvvKMiXzVsMR1CRY1f/1vIC2MY37eYnSt/MezRH
O7SdLKJryZdw/4kl/TlPoE5YytZCwN6GGnuSwztsyaj9wSdLB5aAEH4UMQP/THAMNqNUhGtBatrm
GZJcfJ1dlz8HwmnZUtE0tzhvaBIlL3Jio+UPHpW9gMxhTkKeuMU4rawWuVcgv8etjN2UPf29BIXZ
lXXYdShdIPftCuhK+iMg5jP1DLXEIacnF6TFuz/yRWv3jljnAxndbZ40Ni47xoXsa9dKER0uv50P
aCWpfXRD06e6iDd6JqXO7XfpE4QJBgxe7ruaF8Ri87FfqE98rm42DTIDIq/tDarq9cE8ZotrT1EV
WMMrcEy/3bSV9DhZ7Ccye5Ki9tmqudgoVbgjFX37wF2yW+h2dBNljo52j1Q0H4Ok58iodQtf3XwP
bp8seKpGEl90dmPRAEah9QYV9sHfIBdMdAOSUIlLAZ4cuN7f8p78mq4s4uzKWmqszvmBRC30ArX0
j9iB46Ujo4X6Y+KzBWFVYV26McSBrb45qdVcBjVCIQHc6/q4H1Bsg6F5SxSRAdvDmLawyPzgfI0w
rGOEzw8MY3P2maX4sMnnMZz7QbpWG8sGhbAFcGIZPBFKg0z0vY30RL58SUdRyBk8q078c/+vJjIN
u3zigopLU5GJ17vQUCeVHGbEYGzWfnR7JuWSPWK7b7NyfOOjhxTDI/tItMF+T38iihkKOYaipCh2
OVqN6z4eLc5x3xfoqZJKeaUfJRYHQVGxqsUeYzQGS6cMF+BcAwLGYBkeNw9ixoPz/NsARMbQ91tr
ecwWzabBwrd1z7Qj3Donczgx1HAfdUMPd20ep4kXoF1T1rmNZR7VOUDEOGBBDW0tNKdJ15WKJp24
twTtVPzSQJ4ifZaWmU9GPt+yTXkGAFN/oOQZFZqaACLpUOugnuzSRu4w336M339ZgrJJe4TnMMGo
NtXSouEJ62JA5bwrVOCOlDc2Nx3TfE+FMBdfelJ6wwgv/Fnot674sN44lh3+xO9dGB4QMJrM7tQQ
wC3dHPb53e1EnHAIFCDrkdsNkKt++6G5dYctTZzdiI2o0+p/zktPKW10Jp2LdQ9pbeRO+5ZV5UCY
ON/xuDLGRgzknbV0AEq7LaiZibVO+byjcjPbVFGh0ts44tUFY7BAo5UBipAQCklk70CWKspOUNW8
860pI/t/uZBTnQncOZt/2ZSWndl18WIU7dlm1HixJXVUNyc9epQYiSB4YK1hOaCzKslaody11MUS
SLFt2YOmoRnJvn6E+FjoiqKIXajPFzX8I6kgPyPUr9bldpUh8S0i3afOrrjQSlSqZtuDXnVEsE9i
/ugizpPWfiA5xrWrvdHcA0/uRD5FvNlqCI48uEW0R57a4OCEPXGtEZWDOjwYJN5gmu9EIrby6gaZ
xzOpWaSJMKl5yyRoulZ+fETrnw2npQqXQmi+st5bYHvGYQ7c2Uh1jUl9wRVp2Z/sS0ZMHMhCTfkV
hiiojOLNgoolBLtDdWbCtMKymQ33qdNANkAmS7HEsdEP1SnPvGkrI2BSA0fO7JBsumMpRtB8Xro/
mX0b6BmzOwta6k6kZO5lQLIy8V/QJFnMvt3KukprxT3x7KDf7i6n5TPAmYDxWiBXWOLEr4JZ0fmV
IH0+uZR4ZBXbynwc3Q241pwJEFyl3gM2yDZaQCKThpfNFwIabj4WTzmGkRRdllCav6pf/vgBCK0M
SnEnBeGcnlIcqZlhRL2I7L8aMRgKWvIztBjXyKEPm5nvmlaJLAtm1uplqUIV/o2DYvaEEyj+VvhB
mBn9azwClmo9/6vtCHtPcndLqHREkZzpjM0lc/Yt7I6cg2EkM4pS/kQi01qoWGENKNDyijYznfC1
2oj61m/vZB+nD6aY27LEm7MCazKHd8LxrTjSd1JlNbmjVKGk1rPUGC5Qt75nQ6egPLDDJG+wCFia
KoM6ULULb2ipIeulJtl/Xw3nkHVdEjeBIg7YVNY8dU/XPkkn2nuipIifhtlBLjm6+C1GDhL0DKuc
CqVx0Wh6iiDQCD7gwLwNt2n1G0jFgvDx3qK+YP+fxqloAQKtqp+UuWNOceULmpBokYJucNYVq2QH
/IUY/00HxeD/ZxdACAEH42g4CBvW+4X9p+Nn5IzeFJlERm9bEOEXyz8DlayqN3242cbHeifskbcU
Gr6JAcNydDEqAJKHuIZ1pvz+Q2c931m5m+ezu3OVbgX41lp6TIKBfR1W2e2OKsnNBFGZ7Y2Vn2gF
fVarb6svEz9HXA1TAfy1lsxsPL4p7lT8x9eG0X9XyqX7AQKjHJm19jiNDmhjxNGwd9K6UArUj0CQ
UtK7TAELB0EMG0JuXpdgqmC+AIT92Sxm+Q+Z4NkFdW7/dZy2Zl//7PokxKZmjOchvbS0SeheUQ2X
ThdozhewQS9hrCawkHkI1n2XY02+CEs5ID92ek9cf++jlkiDMv62WDuaFdp3DVyHQ3sSpt/nQsmj
3QTBndfxUgvG/S89hJ/7Bel0iu2dB7bG1s+6a/HbM97+HhTVjIyakdjgHfu8erJ/6RZu2fychQNb
dLQwLx7btko4jMD9PcLFam5lCnli/XuyRQDtOz3c1gKQ7HkUadVHSlsSheKK77PkMc21On5F1VcW
ty9GPqxmEUjJycf6liQcC5Znp3RSF2QjO1gJNm9ruH+vQ9qCmH7lbdB/mjhWnFQbn+LlY/jn2r1m
1msRXyoKu5j0VbwCfa6lRPIJgYfgA6dTVtlTUksrfeVviiQ89JYW5YRxhzBuP55ujYwIw2Uo0Vns
GUig6fg4kYvWJdRwl/+Gz1qa2xo2UfC/7OoyQtiSYOsxZwBHz1zUcU6aiiVS2MuWzjZI9adJPjvD
CC3HN2RX++OZRGW7J57UF1+iLAJlojiLmAH9r8kqCRMdu6hf1z0H/nAeIE8CmI/zcA7yTi5Wi9EC
icojMYg2qzPzMVFuTLYt6rdmJtJZXrSwZWdp65NZzue0KuZhbHeZjA+QrkhZ3TpRdgURLDenEqLy
IUXHjDBKA6piNY2/dXSsyaUWqFfEziahWuyVN1ECZqN594HlSgovzavC0IOLlf2syuTNmS+D7qs7
ZQcgRgELjEzJErGtCN9P6bSPGdbUqN6a5fDwji0IpAehi5fUWX0w/PKwDlM/FeIXfosREGEU5EuS
Pf0qqRmdPAVlRSEObyBd7/t5MyKUV/zoWg2mRT5os3dntYrJak2avyC0EDGSmDl5N58ly0KuFPs2
0PNbdt/Rc7loQsofCzZcmKUI+m56b9Dxw5JQN/TEQOtKDl8Bsf3v4JKQbRcEc1Tm4FldjfXdbZ/8
z3jN7W02oIuRXGBubwTRJtZolmBHIpSnRi/L8cvCrGp4W7g3EZEp6ZaSX9DnoUolnaMKbMMBMYRe
kmcdUMhwd/hznHpFo7T7SAMZGNTOY+MRhuKuwI8GtGR9lwt1iXGW0b/tksQJOUPfDzwkyjC3Eh41
/4gj6zKHOLvMZ/SnkEEypMQ/dHltqduXsK/ST5SLWBvqGLxnzb+8UWBDduo7zqMPzZk3cDzPSmTb
Epdq2W25T3s9Iz0w3QcGff3r6mdtH6YaWNfupWDs+s5vkI4gFCf7wPD3y5WDbPF7vR/GWc+TXDWU
j+onJlOsAAiEMEIvjexuCksbyx1rCIGKecm0atuqhsRynBppiHgoMyQePHgzBvlgl2szPnoV3dmF
KtQ3MEoniUOtRsg1jlkwFMD1Xdpz98SsyVX0WBDMIGZlt9+1WcEKcpEhQiriik26h7/pLmdXvh3S
223MzMl4/SDDJCIrMb4Z9hPCgt7ZtHgAFx/xq+aIC+zt0MLkTM5iOeScs4NjTS1nZhd2+CwcFlX/
DftWM1QFjuc48l9kJ68BcKT/F7a8sJCTZxmaistnw7h7tjK0dudpjPYkxKgXtIJT4tWpZEUZISnt
DnTfRiKItK68Yba1rupNrzPLRoR7nMEvFVueXO8AfdIMNMDPg+ST7r/V31j3GgHqrroT9BHYwYAC
YG3mtSN4nQUgqtRS0wxhoQWJ6k90/UAK/7Fn9nE93ArVOvXt6FJ20EPdnTuC7NUKqLQu2NomvgAN
Ug71nDfT8GcWXhf+ilB4PjLHZsyikFs0x/fMS6AKRDReuNrZ48jD9gxi1i33gjEjHmGRd9b7K0g5
OfuS9T6kWCzfBa8P4ReCVd2NGnltrMfNvQ9scLaHhNW3TE277qF8qJCVhJOVYkw8hKWMoZCY4HL7
k/Pnv6j/c1rZB3ckLDrnDnSnmErOewe4ErXeoT4gcFH0ntL91DUFE1ACwdRfXGvpsLq2Tk3+CKCb
5wgpVVSIL31N9tMbYzn+SrmsH12VXoYj9H7nlLNnz4C4rd95ZQJn8CZVm6/joUee9kaAGsfCBW3s
Kld7/D1PLi/p1cvclJuJMDeNBfrdkR4MJBesiIo1Tjxbwcpd6fFa/R5w9QMV/aSDZ15akklnMmV4
XVgbXdOzoVmSIedRMOOblJi4W/ZUqGjKpsa871U8sinlg4X6fQJOQmHzybszlTyhyANQjrLFogBt
l2dqL+S6J9tjkVgTvK7o3mcTWUlserWjjUa5tTRUsLpdVWw3B0YtT8xfiUkZCRNScx1otjwisfbH
W6l9D5e/4PqWhqrg8noP03qyJq0r84ymECDgPkqTbCsCzKGyrEOuDqGxdwT081m2ZbL4C/+J2qj2
Rm53YS0w+gwL4tkbOZZePFrUgKZVO3jXTUeQfLtjyTN6xHyZA77uFI8n/dS18y6c+A8031CtFhqv
tmsflQ7SVkgJ3GRDPPQ5t1yO5NaRSPGG3VyyVEFZqyuq9xcuOZKkBAqDANx3qEcdO7H5wIh46KqG
pFzV7bX4P5qHFvF3dOq39U7+L7HLfqavUUhtAP+JJ5F7q61DUch6Mm7O0Kg3aVqBDhbOSEy8PsiY
slDB2J810iYDD1bZR6r9uQ4dO88wcmLymhalDFYU00mLi9EK8dOhkJXJZt9Q3FCdkZqyZdFoI46K
lnAbrybXmZZZ0xzQFwRVIm9p+X1V9uEzTjmjTfnAF7kmx8Q5xXZODoUIfkl14QGPMHLgeetE3DOT
3EO7bF90ND+T7tA4TNv+ZHBTrSU4XE9gQ1TVPQ/EVS0pot5gEqrSSXKyuQLVLI1bvCgfniMdxQQN
Ix6oREvBJS42IH9o6NGFY9eudJ7Z84hflDnXFnTq3Rw4PskFaGvoblN398301wiC4kKr2jV6FnXP
5M7B/xUxUQYKtGdFgpT6mDINxL7zZjvRyc7jtT69L0bTNpH62dQokWj78f5b7oGMPzJBzyUFjN6K
WLSkeBkLyAKIa6M2BmMgtbX7vi1SKcTGHMABec91hq4AT7sCuADHLxVmwnqyEgG9e0jTqFXAUICY
d7raGPg0okZJQqwXVej5E2QZMpFtEtmJyTy02k7GSIA1xOP2w7AXY0OsDXxo6NXyZlUdwFLU7G+N
8OVe+W3k5l5R2R7IuZR6rOxVicqhl5KerFo0cIqiSb6W91hw2da4HJ3wjN1LzC846FqWbrBIFaY8
g4UiLTF77iayvvPxcg+cr21Nf3zhRyaYyShpoDnaYnOg/b0DkqrYbQTK+7/ZMZWY6klMs0rvraSM
JtZuLUFUD2Y5LJLMCM0Ra/xzZwwMTvkN3fMHqQzvW8gKDWBowfrY4QUalGvM3eSWsWCAVhNnFz8c
/mHPy2YjewIamVFDLg5l5kev8fhHTfoJXU4I/uXsZlqpBjcdLTGTify+rNTpE0RxdhZmnkxknBgc
ANKMq6v2sGYurl/FVbqdVmAIG/q1I9KD9YgKy7daoHsmPQCBloiN8M19+z1Cf1ZFEePKbXiQl8Wq
vUerJVpRDEzdhJr+fcpEdZe90cWzjk//wCdU1Elcc/eZoYOYwIuaFonzhBSC8f+W0M5QL2P59GQa
+5oveSPe4RQ2DHrog8D8fNOpqqmQLubU/UwRYkNbY2pIOE5dZ2MAKMcxQ4WE2SWbpTmuVDpIJ4i4
IPC2DDOCrG/h/7PYWDWDA76bmHFfiVdaQBkp51Qx95VWMnvFRLpn0cOdZnx0sTmwDtyWdbzxLEh0
U8+U/H3IuMYbcR3ZXKoNTFiKyH6Ky8gK0r9e4JilX2HjZNdyVIXd2GmS7UEOnGoT8tG2T9t0GS2J
2ze1+e2M/gSDC8pRWUrA9etLEKnwu64zDHEL/6AI2uFXjQoVC2GH7+8TKHWfaFKRwXwNdbguxB8a
66nJUiXYnWjPb3avK1svubXqSXLivlVSbbgivNbAtMP2T38jSJ4+ThQ3R0YU5PtPZNsGY6BHM6Jz
UdVKB5EQbM5ZKPvsXulCbsDzjbwN9cHRewXSMOfinOGPr3oJExb9Xl3I2rmRwRo3bK8IuFpCc0UN
qwGFbh+1ngZZzS4Gy5iFD0sAvB35bIqUFwGq3VWmcx2ggwGT41V380AsXjnktPaHHESng4AlDdHx
krDkmswMpiWWTspwibI5crPAjWo9OIfk4d2U4W0Hf95Q+3Svf8nsntko0wvO1EVGQatQ9alFGkGk
1BcO+hnNPnAGHwINWHetT9x1V9GdAXor4V9PW992VsX5UyJeBmbMaKJ8SLqd5hJCkn66nGw6IAeM
qOTJqJMV72b0rYg599MWPE9e9e4KovQAdxRJxOtepHiGeU6iDZgVOjurr9eMSKLPuV5sDVL79P3w
6A+UrJyuxiygQ5WWpXWU27FJ9AGIZMJmTeUAeAquRnO2/g7VB2IAUnuF5CnpalS/SzyWnK/gsvNG
wzievNr1d4yRdiNikelQBcR8WEmMZymr2zzi1jkdDBLsuPJOReHD6YByc9hx2QrklTLf2K9kByU6
3udKKS/MZRsZaU6vYQYSseXsjrTupPBjkpbeuR3CxitbEBJ2NwE5mqnnuhVUqUpDottWH+RJsREE
ARZg2hkOciQWEun+4a4HSJla1XIc9xa1UNA0esWjIUXs+ALQsiwtQeUKs6Zk+Ie0jFCGMsw6f/o0
ELyKFSxpnr31CdhbMzukca9NAZ20pdCkcDpJMt8J6p2nxPjC9nbCryYu6mOuHJE4KXp0YrCsRA2Y
3N8G1mIm70w7Sb6OcYGWmtvM6kIcztmI8XtNNl6mF2wkf857F5PknTPMzaFFPopHtVJuIylZcUO6
Q314Nnn6Hj4FCzn8EHnh9tPEhM94bHi5V383QO5JKIiwGqUp08CR+TTDR+flPkzq4s8wdg2U41hz
dH2QlTvmEo4iZE5ZUZPlUPMiWPBKUJIWj+OU3fFooK8MDvZ/YpZKp/Bha9KZB4hKZRA5/BVS7gR3
QLboNn0/4eWG8U0FwGAdII8tsHUf4OSvX2FVQ8UFph7DCFwxTKGK4zR+LVz49tE4PcevYgQCYMaQ
8RCRHCRIRyMKag92B8+CtlYZ84/urEPHN9E3UXM/0ycMTlOcYKevWd+Uosh3aRiYni+PZWPPuYnV
lYKJcGcgoC1cXJ7b6uXky9D8kOv4a9XJJlfmMCs1e0IqAU4PLk+lFJrWe1cih+s/KBfbySTTUN14
VdTc2XaSBY6MvIT7ZaXz41pu39IZZZ06zX3h2Z0UTcpwNTB+L1i3GkpPfxSQI3IZCaQaF/ERH9NH
xrhRI3uz7s0CdNmRNvEaPeUQngALZMGTd4ejNSy790MEXyo1GuQZVKSdNQkRR3zFZ2ZSwecx12QR
nguIMbYyKaEZGrJ8MiFEVOTC/DRomkJ0pbLHSsUgBldm1jkhgxljX80eXVU7IQ4B5vbIdYjkEjR7
9Q7/7r7f/frbWJWON8VZCMxxTo3WoItWEvUDIt61uS5RLqD+z5fcj7pZmLigzLAYrzCvhdSj/Va3
mTvGNbwHMNJAPVP41eAy46rNSTZccMmS3VTpvVAuibceCSV2pelCx6sF2ivJa54eUYsMWD0dGxIE
8LfvY/DDhuGHQ+Wb904y4HMcV3b7uOJQRNWL5RMFxzQp/cJvDrt2TGkJzrpjEe9EEtMDxq8dKBBt
OEbHE/JU/JA0R5h6JO19iz6dKR6ISH85mkRPBzWwJPlgKrkFwooZ7jBnQWvjQDSIUWMiFDMcMkPb
82MzjmTkfSImjJfpix72RKUHFxCybsxUj2w8V3PK/SioPCqaWSS0lgbDpZ+ky2mOpf8d1yB6OIPm
a/+EFQNQq/ApfYWcd21jTQfJgfj8OyJYNRjcjbpwM2BVBwtzFnAIuJ6AwOO0/D6YoYpZblHEOp/J
QMUvU4qgzVxImoc/gwayyXNLNsntGk4i8WARycXhsyix4ghHephaOPil4QyAC7hCppnI42EsNNqw
vGXvifDp0uBqmh4hbHnvxUWF2/S1Ox203ikGAZqTZ+dJDKnGXwRhWUsmNDCE+c2xnRkxj5QRH1NN
OxjXvYl2YYRn2s8G1AplihGs6S+AvnxQ7Gs9z0poyB7sGLRLpNKJ09WumowIW6+WKzNpv3xddgLX
ws+Fdl3MtKMAG3M9pvjvJWEkhDI98IOjhzC//koJD5lSYE6U5lahAVQbG5dt9Wl6iuEkH9dHgTlD
4SbEZqYGz2iv2NWzUCb8p7/knnCzOwoOoPqs/vWnmQetbMCGOcJ/lp9RuFA4bSXjBw2IH9tt1mSS
Z0oljjDRlxAAOzs7cBJHpCjPqbZ7/Z6AnbzA/drESHiNoMVvOyWesOo/tIb243Hh8YZhHrv1XNOp
yurUT7spB9DuQiKm6/6vDJN7GSLvV4rzcWiIsbv5Dq1Lwl/ecOw8HeiYStkOpKxmHwUQ1LMbqutA
LTBi9FRCZCpIhiQvfslXyOrUNNSRTJP2k9/KrzySXnILmUXRx6QGAJoy+JTbPysfVp4R6Lb5W1RN
tBSfu42Iekrr7jwQ6H1pN63sIAJ29kSCP+6Nkq/EmZdHIZ37JX88AMw6qKdUoJdM9hIbfm09nLZp
GQT0pOTj5Mj6AQhEYUcY7zim9du/kjqUtgT9cQcFFv0+jvdrzJnPFmNYR/bxLYwknm7zTg6U/K12
mmp+UFaWlLQ0ms6CIlqgWs002GwYQ3m++8KHbp0yz3uotmoN/4idd3LlzW5FibNny8WgvPPmY5OP
WKukmWbNmKrgpL+sNQGdKPMw/l2jSCIGcdPUSVQwHrcOq431WBUEYTrgCxRnspdYzRBnwFvBiFFQ
+JxjJ8gu+4Utce3EfuiuE/0TAP9Lr2mdkgBlNKwEiFU/Z90j4jJKpUiMiEbUExtni4hfjwiCvK4v
au2MZmq2PUcx0w+HLZ0adHnZeALYbA/Uo84cQz2Ilc5KVNdvMssR022XnSgg8GioBPHPxmIREgGJ
hv3b2ymTsIFGXJBg5AbPapDcNHzkawPhKlEH7UIx2jHXA0XfRMXLlu/V082CxbqyM6vyQKEEFg4B
uGjQJzh3RXbE9wR3UuDF94Hg+hlTQ20QyqofpK4GHLbUPVTecMlslYQF/sEYref2pWsG6r++U8Nz
kz5iK3y+iK3Mnglypc4YBRTYZa6Qbk87EUi4IWOstKX3s4/aXKSylupjeWwrRVVfJqUIIsct9uwF
Bke3niqfGl4s/on4KPbrn0vwPDF/1wCviDVxASFwWItEeReRnV9ClVs+O02RD1V8Jxa3l9mTpQYl
6aUyZ8rfa/RKyckqHl52lwKCF1Y/1o5jltenXO6SEGi7WeZdV20q/tJ5PlWVVM7Nn9hxzteGUhzS
RxoTTeuVCnkjMId16UZ9sz+NHwHooofRjcDQpK2ZW/L39Gam8nfGLLjpu80MThHoF0kjqCwlB+Qa
ozZTq4f4yFlAyTwX+2LK3h06lg/l7IhqFSW5Ov8gv0XyKnIQj9iF1rKQBMjrGJn4XrxTyzk5SPV8
rofCP26pC0woQZN0Dbe8oDMC3Yp0BEIWc6t69LUtGX3BVaMicBMGbBC04eFyve43SJRVWaojKdZT
KMQ8tm3oA3xM+yvcqyee94/CTAQizIGO1MonzJlwBXCQP036EeAaoaYea7oY3VPyv4IiUR6QS4bG
ZwFHAMgUjz2zHTD8kt0Pc9wUnbyU8V8/x6UH+qXvDZIwYObB2vDXF0rXvQ2qMdpU0Jhb62ENGc+j
CxNSwPhWKdNy9zNOz/ZP88WsQ+tcLPoSHaQYt9yK1i53CkBf8h5L1mrBjde1NQP41+NdXgnd42rV
t9yPIhTHEfYeltWAKDMvkMU35ygcpBkLeY5qnAxTbxfZm6Lb7eLU6kIZApggNrzbTUFwjs8vR8ho
CbLOJLGUSlVFlRVX6s8gHnyCvO4qZ6QHUwfl4kTBA7Mp7kEEy2sQLMecj0DcbeRGXSjvkr+MGxTb
6BX0bpE/nW7+jNqXhJ2BWI7d/oq+4ZXZN4hiQlUocTzvY7WETq4FQy8ncoXpQJkmYc5zNc4gurw8
smDG6OcdAhnXu7yK1YNpYwWFvqLnAhe/GhWvUyfdVjQPTVtuiRm7AFZkEQKbOuhBBcu+snNVsher
cjshVXEeYYM9mwgMDwhpqS0++lUI9f4Ppki/hdzir6b+Sl6BIQ2/Lgn3mPtY3heoqmvsZ47iVtQ8
8M6Q+jm3oAYD4ttILlDIbcm7HsgIi15bo9/OVASoM4cRCOcmyyrrdrn+gyDx+Thpox1ABooM9/rc
aLdn3r7iiQIrffRIHjGtpw7oVuNYYB5WRqr4FkgsC/nXB2IAXvz2jKekqTWzW2/ngf/lHPuOfU6x
eKh3MzZHD6z5DhmZv+vWRtK+1PHRXP//idVegelowiFlVgD+HoXuRsei6J+AU02LNDxi6snQcJeT
OHjlRcLhwBruMxmlGE0LLIKkWhpDeIyNPVJDIGBZbLNIKTYgMlqvcRXgmarelJKOIigvhM3WcHm3
0qgF7Ah//r7jfvVCn79VSZ3UJgCmKeMTXbXsa9t6X2Bdz/TZk0P2mdlyHn/P7yj5fNBUpWhmy4dF
JOnspusbQ9aMKDseXrx4pvanpMm3KwgP4boQMQ3f5Ha2xH2GXxwiHiHHT2A8ER/JlugSxazUOL8Y
nSl8nu00grSZc9iKiS+4n2amflwDXwWjHjXmyjCmMjWGHp9WgdrsDAHAKlBA6j0UzdlzxyHLOQ0V
+LUOLeCLIaAP0GsJJGHruqu4moexMdpp+em8CvswdxNZUM1xTjgUFDCws7i5OOe9fRolyZqT38y2
HxnsJfgzBSWE2/uJiKDIedYehttskOK0q/8RZCsxI7D0lezB+JufSxexCxaENJCdZbfJu6XEd+2U
Ohc/ePZHppHWq5l8mtrHwYzkuJDbi1564loKmBeXCL3TpOVs5KzrcU/mOiMISHCtMkO52CIcM7EO
Dcplka77d0F83hc6kV+CCFQymXylOjtaopoxWImKNql9gYTl1k5de9KVoKcj27oUYlcKx4Dv0Btm
iAqnvi09dAuReSFFrwCbrWlywIxPrIgg4qw5tKqdiqB8q2c0yRTw98ErwmsVbj7D12F137wJVFjU
2eyWQkNUPJ0S2ISdklTfs9Mt1CLkIGDKanteHvAb7+ZYdDC5OuwVo/WjVNXOtHh0HOtS08OBnxvJ
AiU+Wo7iu6RWWDLXU3gMXav76fdoQbg2Zdb1L6nHUjyx+6D2yTZKZEJ2AO+mT3cYNwGK6tw1BAnJ
jFWsCwVzkq8AINrRQBlBQuIinAklz+EkG+2lia+RCLMC3QKbmryFNtdM6+yZ6jaFyDUPSCAgDoRW
ddL/m0NE0LiHoI/jIyCUvD+Jbxx5tZoI5B7Uas3246bPhAkGaRlsrLcf1BkknlH8l39JxfLKGCQM
r1bdLTPiuYmgfF8kLLfKVf2RbVsbS7AZ6VG+ZEe0B3/VNCt1kV0YGPSu5waG9DD+f/8Ch9IwoAyG
HsMa6nW2pDj8oRBt858sSWcbgQInTq2TeP78q74dMCzlPYbfQmoex3Uz6LvGQ4noPPAhg+wqvft/
sYqYsTRA3Ss18zZZhqNVUFrd+HmTQmzxEq+sjCXxsijyVec9MdbLqFiAQCJRDHaSU0A0V9G4mN80
g4rpOzEKrqihSoV/qWzSP9jHWQQ7a9KwXnglINvej6jLILpzdYOVUvL2HnxUY1wgzk7Xa9pYlR1/
5+tXf0nWsGBf2pac+IT1HMUJy+W+ZhjCRlW4kKWhFu2qTwJnK2gUE9NuNpb4ylowpo8zbj8fANPo
6ZxIv9oHZyILj01sel5NdDM1688sXiIbiPkIoUx3K+O15nFzUWFF32KyqH336jYCk+9BTTY7sUe+
YplGKb3KXaQwQG1AeFxPqCUPoloWClaEolSX+gzQ74fMFedpCKjIopZPY3fmCXiaarRt9J7uskGM
bju0m62Am9TuuoOLPR1n6SgbfXRBVQgn7pgmU24WFjrr3iJAGKM/6Fv+UJmBqFJNvGq0BmtLcJkx
D53EKSDObXmySrCcWBtUNtkLDBZbKbQlHbYGiEm1fdQN1iJxIgki+C1nkRBFLi0aMa+7aOCD2b6k
eJSL7/SWwTuQFWhlp1CFlg3M2s2bpFkziymZ5ul1hUpdkagxeTRA8ffkxGoskkaqelZLpNTqVDKO
L7rgxpbWTYdSYyjs9yzFwy3a0B6j3Gmvp5r+yr+D2ztXTqgoIlGUZbpJIRI+klYjr7LsYJeovwHN
rJy+gDKRJmWPJPGw/Tba1lqkSACY+LMWqSkm6evLn27iapMXcK+xwAqOoWf2pqGIU/OCWoSzCgG3
bCf2RXynumSphINkpvzfQzmm4kmwoiHSiV5QUyObngQaPb2vL1cbXLPW9Axy3vfbvcZsazS405E3
hkXR1xzOWPXEjOIaOd8wzUftxyDjQLt1RegAP217g74UVDNDhd49OcrL4UkANcZFx7H6WyPCbd0V
c2hNGwGgTxyimW+6pZK5CQdK3z23/kgmDIMxE4O+oKQjXyhh8v07sG7/g1GZwzw3Xx+SBC9Xuj33
Kf2vnBwQ+g2ExhmaicnhYsjHmmuejr+GunqMwz8sIYVNhk20K6LNxf+I5MkfXkNcfvWM6/nWgqCf
3Jyz1xLAz/A5vL4MO/cZnlFnVg/mgt46ipXYpb3UnSlrGT5Adr7Od/lMb9GTHopPE9gEoW0s9bG4
IcvhTUlroQc8WgOxBHhL/BpswhsuE0woJM5ytLtoPfXWVCRTnD5oiQHjaWHwVsjQVY93VYsiLrVr
QMHHG/n048StcnD/A0Ha4PzLHijKDtjYBhMNhJIubg/gZUHhGOClp2XtwKcBYMdlaQqTGUPpwrwc
Aw6GVuVjjuAsJeT0ZtB9aC+IVpNsJL8pLYsJvHlm655yVOK2lQNzLCUhgv8uJY1xgIM1YCM5wyg+
X52bFaxjX4ODFOezYzZuEi1MBQiNYUP7NkO+7jduwfHRunQ11LgYMxui9HrJojryLjNsbsFrB61C
aMLaXNrJqCkHRcXyQ8mJazl+X33iUqDzwdCLji8f6Om4iw3tC2fKc1nvpARXS0BGO2KyRcPWZxqU
yb6y9FOAymqTONqqO4rA5eonshThnUviN7gHIzzxZ7MbdWI+dYQC15L9hXPPpMn2hkLRSAL9HV4h
e9ywOJ3I28rS0E/j1EjOWPuFR2tRxsOkYRx06Wg2YZyfgoLntOKt6jDXGDDM1MHMdmOzN4g9alG5
dE9mw3of22XPCNKanpOwF1GyjuEMJpKu/E+Ctlq4B1CpOTRCUEr+s+mSoid2vub4MUevOch3D+Lm
GkufDfRjHUsMEXo62K7Fv5dHef9qmZIS1dHz7H/16Z3X5uWeVj26navKivRCADT1GhL4iGAMGd2O
urn2ANuMO6zosk5byzNkdX+5A/KCdT3xJbn7gsk9+P0qv1lSda16k6Nud1V3rfenZCMqZmUxvTIx
2rUPf0pUxEQ/nNY/6aywq4GmFM7jS725R/60ccRu1NEcGIFfGNpwwNlVttnIkRiSwW1dUnV0m6rc
4ThMXnbEBnHeVRcN5s6nIid9iL4VmrssFdf4K9SNrsBXez1RIQvrUScZV4fO7bx6VI5yjekMX/5n
nnxuY9VjsFmjiug75OhatB7f5VqmhCZrKYSi2LxDaWFYhYIn36uDDrWTCnX5RzOrlc3POQLG6OIj
mquAFNuFXoSAffaHfrkte87uVt2M60wrXJhmV4C/XIR5w9sP5ZYRVT4YdKEha2re4TCqRw0Tps5Q
+LXneIpzttEpE/LXW+qqsERvFhFU1yEp+lpBLtrxzozyYWxWrtCgsodEpE4h04pO+U/KsL+1NLH3
YSufsXcV6xAtYgnVflNvWANsE0VTqLcqnjqO/sLlgTNDUDhaZI5S776AVAqXCApA0Z2RWajY6T1L
1TbyhiV7Q6XfFSrHCxmaxLg3KTzT+2uyaOYbl+k4zb4yHZwhwLD+dzSE/mpmhyWSbY8qvFnDqZAq
ok/tSra5ZKp14HSRXqHvYJuU77OT/PbkTRRCYEoan+zV/MuIErZpKbavt6gVkG3x9p/cjAfXgnQa
unTE8CcwGaHfrfUBtQijunE9wgtzV/KYM79xLA03lqlj2J1aduI4dqNAPL/dK9/4CLj8lfaOvx4U
f4fJB7SGP8NecoamBI47BYWEAqHGnsCmsEgWNVGHZ3+6m7o9XefjBvN8ZLZ1x9cEtzJVjGclLfds
1NbVmE9yiUg7kjHHbaUIgWHd1Gf9EQErYvEliLflUP8LHJpPrRF6bHNKu9omlAPyxN/NahLi2yMS
ebmZP+wP2+a6tkghpAC+ImV01uGJkRfNe13ekmzIvoacI8yYBgTyvWS6ohNuE+soEe3nfjxH+eFX
uHaKjNhqaJIdLK4iKwAXppx7yKuNdfJLdVPR0uLIx/ENoxBwT3xUGiLJCqgi1uegywKm/vxT9IEb
waGA2oFnjQPGYQ7mSzpIeQW6YBLSZxzCS3YXpV/9fwM55y/2H5mEcivjgQ34oXPME1mHy/exPEFh
8ob5aonYhGDwf3HqFM180A6HsnKJy1o9U0hWtuG9+1nEZghFSYN1Ll3ZDrArlaRARYSt11p/3brH
7+QLdvkiiA3UM8oMxDM89DW0TTr70eUHNr9Kr3oSQ4Tu6wwKpt2CkUwAsth+RMgMrcVDXUuP2+n3
syebaK6tU00NwC0xz6wIfMHzUK4CCA9XaaCJNVn89vQIyW3/5jGnWb0K/DKDFZtLZcH8JXTL6U1R
nkv46Z9irJrC7EWMhlT3FqUlXQq27LqnrA7zG4afySt+h+bmZ2ecMjCIFVaQb8u0qBHbn5qcvs39
m42SCc7W7+2rYljTLovibxgkW5AMOKCgg45iZd7UW044Q4OPJYSOmYNGbsNbkZRp+AyfkfJz2hLo
Jcv2od7WnC3l7Jnn8k5bV9FWFRzF4p2HXxWU4SariQX7uiQn3I6a/sPaqmjCzT3fMrTqAhqnq8G8
nSG241IXlfOjznItstLPAgysR2Z0LsTeyc8BvsugGbDjbcgoYNQe2bBApWeHhYaGMEwUEHGD53r5
QFWRPCd+DlOV5pb2Zj8Zb7EJRy+5H8SUIuViNIXh9Y4xXAszkvTLANyhYLUmw6k4IJWFQW3Hrm2l
2nFj+Rpx21Fq9UNAz07gxDw1yTpbbMAjYNSli4vwta98FQPzzdcqNS3s6d4Rm9MjMRadkWKJ1mIv
Pyk2qbRCJ24GeenkuOlprGJdBndaGhEzxFSemJdmYwrFn7tdoaeyImT1h5jD7v/3Hq9BG0ZdrpxR
Ta/3BFbnmSke172FSY+8M3ixpnfLptuU4DO88kg445P2RPwp94VpMheisfoBLjwdNzPczu7T1ppb
DXOY30zhZXZz/0Qndm0OnZy+bEjq3bf5siH56Oj1uJB2g3pUDj7eeLmaZZi+hxJZ/dZqcsR20+gj
KjKmaMwbP11Rur9qhFvB9KNdE6Tv9y8vYK6kt8dpA1gRFs00Pl1XZeHMaV/ONyqNJI8kKDB1ek0F
vXkltBLfCqsfF1E1wFhr/TUbl53yWa7kC9LVzg0DenoXbf3n1Kv67sXH1tB41ZoN8xDzo5bZqR5/
DGvHcqENpC61ALKDaoEIZuHuCV+MSy8SSVShWmF0klMAPGbrfVa0gBslbujvX3RSA9yo7PCCwEsd
t2DQ0EjXw1KjmUTNCRO1O7f0+YZpchYnLGbXJ4rOVvNjB+EGH447NdYhlt5Stk5IbC8tfyvr5W8n
e+2VJUR5hKaImLBQQgBA8ROcEIZZ8VC6WjAjtxvKgT4q/WCGBdrKgcZlE4Duu+UzyaVB1yPwtku+
b81obkj8i49eTL/9doegQ/TZ5x6YgeUGzE7wDGVVtooX3Z6H1uUqA67pByLh+U5PWAG+gWScwdM0
Ra33x7H8Q8i0n9hIrp4D84IU5rDew25sWaOleURAnTqyj4Qipza7c6HnxAt+MvNp/JCQ1YUecE29
CO53jsm3xd3x4QmihW2ujsY8r+V+FTi1/5pe2ps8C7R0kXKayCAUgOn+oAA+xZbFcRGwT6Hz7uHF
4ejg0niRK52t0w1YjjgmD2rkZqRJ29uAlKJ8ZakRmkPFiGzcDFaeBPayUIJIWUZ2x0t8biZ99QAG
R7ix0XyKpE0K9fzZUkv0KUl1RYZ3f3J03FW1sssHgLC0tSQjmdV4MeojaUjOqvVoUO0R034IDteM
XEHTP7ipqGlcLxemwdgtU2wnCXMyrj93wBB71QCtoCoF/6+95edzzUNMo7KWOJ9w5pMsUpT2cPuY
U/QVp2kcHAKWN1iWKxro5qgh8H+8zIs0kzpX90fcPWHxrqC1bmKPrg92dFS/cvCbYrMWktPfj26n
0HF3XSch3m4L5IdBZBsgw9IRU+5gDVpoAZvdjgI9LDWjxw5JrXseQdpeKFwi3ubphOVIQWPwhDMF
LN/zb+DWg0TAAN6OBpjmfejWL2QgPK2ze6oWgBmN+3V/erIqZNKK4IQUltBA228Y55ozsR34QFN1
CzCHarKt05Yb7/cmCy1kXBjdyRoW+jVD2BLjvFqQ4NEBBcW/cGrAIKpHAcKghT0pfiDdKvnymbmq
ZuZInKySMUqrEVdo6iXnhVLhZhjgzmZUYGJFzCo9yuWAcHQdo5jpx5M3qc6AcP2xB60xmUQfhUYo
ro5H2Hi3uGt/fU+zE39fKrFlOvxAzYP7zRjeCGZYOFN+IJLNVoXbwZFaFYaMSe0EkbwtCDXG/x6D
JKsl9nl7PQy/cfs3ieTREG6fTdmRAI31f/awS1KdzDcX26GiupAzJv6TiB9NINF4D5o27w3tc25P
FH9O/gpy5YfMIicWgp2Dbe+pKVHzy7mu7McC0XjTPnQrFJ/Ejq5POlTOr62LU558QTjMpipRiU9h
MfY/wErCrSVsTTwoKN3r0mf8FWhicqhgpKy6H+NuBjysMfn3N4ADTvsTVDXvXw1Kx4Ag5ePRMqVl
S6XnJMM++ngsuQ7VtNUsx+ath/Ah30/KD07maSFgAGp7w/Axv4u/I/fy3G1NlXvhcwsIC+58aPV9
xbUzg/GLcPePTfWfLClPOGzyFJYp2lCjPqf37QJXwk1XiqQX9vT0M1rYNr1xdrECya1DNbTdCdsk
KLXO2scUdl8mNSRRyReceXC81G3xOw7w5beuPbXP4871m5JteUxmwM0HOlYTZWzt+N6HTkVwr2eJ
vQ9+W7NAdB+jTvsQ3BUcum8iwiikVjK+x66X+rgdYSBKKm2ICW0vlEz1mNSkqK3UHbg2lHp8hCl4
3SN3Yo4D5IGW0WqFOS5aW8TAeCyRxkacl+3z3R5MqfMbDo+XjSNOxjXha16iGZYkfo2H+XVOTMiX
kFMfmtPGODcxLeoQhIlTTBnD6MZPeHuNxkfIhhfe7WITzqXU27rjiRdcnG4ZjCW9QIAU3dls++xi
6QxWgTVcQPcWpotnznG3RAKz+t2itZEqfZX1Z8tb137+U88wsHaAAeFKEAEaF8E9IDVS9OQhuaag
XG8l4aA33Jxyc7UUMLK1JpixQwjXjt6/iMuHLAc8uXwxp2q64Py7UthrBYENwLYcx9SEgjUgF5Zr
aJwPqjZemmwkGZvi2loAWMdUQCgw78akoz72s+DBYq/ABYirb5k0p/BW+s/IgncrcrDBTGYKGiNV
/AOr/D4HoBXOmeS55ZviXcoH8VC4VKBuk0HkRAimfc3BLwdbGSBlzIKN+uvxPY2GgHV2uipj3xIQ
ttxS+152E3fMiujytXktrnNgEmOSc+fx2gLwFnOz2gO4z2wrl8WqNQcWlE6cZ56Ba/fg+jdyenbn
CVpP1NWF7fMwX7kBsHuQ918K7SNUS6nNKk88Vw33d093ocUxi5/7cIl9rBkClycQUqn7elD22kdX
jOXhqnJZgefNc0op5uKvZb2LRbgaSKOXdrp0bbc7FsRar04DBmpjLwckTkLtxAAZpLe0d53ByiWP
aqLWaZufHMBwQliW21Zti2SYX46j3D6h6fRvg4vtSqAKDOt7z7Fb+mzo1jYRFu+HpDjOS1VKTD20
+Rp1CRXJcXhpahWhb/fRc9uU38+NeL379hVMGHSfx3PAFdA0QdfT8XWZeP0iTQeiQVVVzX0JZgrX
Qs02NyHrqDJef/3NLUiutuwfjGRXu2IiLdsJifj0d+dWRdTmYNfX/ZO04hlIcoi4WaXH7vxNoDih
iJM/fcI8mj/r07tKlyYOk4TgKlAXFjYp/nTI7I5mPoUS/evBSKFPni497blO84AJ5dRyrx/OjVua
Tt0vBirCj0xUgHo4Ivf0FrITl+Vqwo3ERj3C77Mow9jYcsE0Vbj3hWC4AAOGTuFz3OMDjJ/bivks
G+1eEGUGn0RchUjwsT1JaID23LK1S1DZEvEZVWvwCdbubO7/QpD8t3gpqbmW0tp5FAiHPuNe3WrW
y/e5HcCPbCif5Om3rwD6x6PAIeYWRPNxdTWTBwgQPfK1RSCnXigH586Y7h+dZHwVd4JFXuzzY5P6
h5sPgCBTQoI26EfyPaUUWiRq/E16mYAdWQm8dH4IHuFNDdawKhtwn3PljEwAaPOPmmzhX2JuoQo2
NeX3tpFOr5VUTv76UEQ1zKLpafRdkyi+KajWwF0H/VHpEFGRLGHf6ZqFtEykF6pW/JgrS3ogrDd4
2PIuM1x8ip1zsfEsjM3L3SFZb48JV9pOEXH9T+TaiToDSO2Y148hI1HQD6clSS2R/Oye/IotNB1a
uRMpvrv8YTWwTLtHhyOUbMNvOfyqgtS6azpIw3q/NTUvUSFhY7+uqaSOEp6SCULz21jEND/61SIM
KVAucc6YvyYYxqXYMokXrdqlHB80FLOuYVxmKtJ2OK21edCuKb+hN73P89KGA3wlgwi68HwMLKlo
SSjF1ewXJRWk2FypLjcf4TpAwQBDAz5+0jz7mXa8hDoMTVJ6zcw53xYwtWOflOBPaCWCFKAus2iz
SyB/THjjr3aqXFSPTrzbIo04bf1wReH8DEdlRwPjTKyVi0IPxk3NcOb521y8+zJH2dJQVXJOJ8N0
5Dfeg7iA2kkfZZryVjGi9DNFKHUZjxl0r754ZiQTSFSYKsPK2bctrQ+kXz8p2rKCaMn0pD7WyCYo
h9jQLK+HTveslsw5u4WB79dxcu6hY5JuWN6EHLUO9E3iL4c+tQuu/6ZXnRfFpVdc54RfMw6Hezou
v/P1k5sYVmKUwdLFpglsYGRP4XV5+gIyP51N+Vc7980kfA3qs+qre9+3pjd9CpaWhMjPgmlfsrCc
Sc7VdUwiH3m7PARTQhngNNcW8CGsntKlWUvf78aG3OqMLjoZWErs6ffkrWzImkRSBvf3aXrl9KC4
gKqlZ1NC+1Hxb/q7nA9bbGv5rBRRGa8HuuWCSiqxeCEVKtmI8SGN1CNJygTiFxzBXQvPzUCsgVP6
Iowty+jzRBupGU5S57TygvPZcGP8SIlgTAM2qdhrWgcoTINfdIcqT44aQUrPgioHT5MIBKdwNnv+
AihxH76R68evnWTF2O7Dc7fNGY1WcVSFJ7nj6oT375jLu0HCqPB+OBdwcFggDOjz9wNEqDYDp34Q
5/BgqOTkboSNbca9kzZu0nAAHoXc8x0jyBv77qJgI07B6Bp54lvJGU1ZBqtoQXGCUQ8Eult6R909
sEbuzoKswQKP/VQIbC7DjQTjdx+b2DaspOSrETs+XWt1uc8XSSF8AFensw0VNZ/k18vXFJllqq6H
IB/P0pMqAB03dYDSZnY0Q8gfUQu90mPTk4WVUtlc3gg3Dk1GsDV48IMAStwWIH8S5TsEVr2FnWW8
TtZPQUUfC3yH15ea0xezQ0Go2rUT4ONEdkDjYIgh05ymRDcnNGeErBVvTxT2QJgcBbzoETb4p127
FPzE+cBFjltKA44IAld94zNshxPg2XnACEASKT9BQMquf8x6FxM3fhxpP/7n/8uR1huWq8KSBnMC
38GXdr6A+MrJEELW3lJcqlZzA4zWbGIEVGOf6neobc4D+zYrKbyHCkSemszhrCGf7wTtXJulmjGM
pJjI35EBGEmuYl3He1kXjf5cGtjqh99vdW1bDLbkPB9RMf7Sl9QayBTSCz/ynfSOrWjlaqxjQxE+
78svDiYGUH5iRk8SzffDHL2eldCeEx70OtaX8z6V+Io0xt6WfjLqHlzALdgpFRSaTvVmFpKfUdTD
Kyhd6tia1Py1NXJzd6EVrKUAa3nb+8ZSUd9pS+wsbCoat7qfSihMt+FrtmeLmLdq2M0DuSR5j1BH
lytUgRqa5NIRq1xtyZLJh3swBE9Ak2zozJFHBh7tqYGQKvIGtkDUBrw4xbckoxF2rVCxDWDFOdN/
STAMgMNehJk/ZUpKbcEOSG91XrciqXHnDa1I5hbzPNX/CsUCwIQU6teKpsDvjPQoajFsVww8CFOo
nmZGIPu43aJgAaTvTDKWeeD+vAPdwXAog0XPLIUiBJO1s2Zbd58+D5ubSSY0i8r4717h6C2N7TkM
gZWTOKlgEYipDFSIZg56F+Wy4fG+Z0bqzc/Qbedu5TWgMQD08WkqVAQmOqG6k4A37j4VzBsNh/iK
vZKRTyyN0/JOLEbxNvd8zdTpbsLL/ERZcWuSMIBxyp8QpNOn4cldvuATJl+i8kQ+geeSFCMV8m4E
F4oijwwDCTK4BFIjLUIzhD/m66QbaoXZYQOiMm2awfV8QaphcGU9TQM3KTiDxRZHR2kkr8RdQdAV
g3x0SoDrYd9YF9WlLT/cSJVoln4/rsj/V8aHQq0lAb+nPxp0h+51gGtQ9dRq86oGjB8c5BPsysyT
O9284QI7mD7lkC0lOf5mMSw0PQ/371NvLPB+gztQT6MILs0wqieVaS6LQ6FmIVkCYdp/GwdwF+Dv
ehHeqkFQt7EmFDYmQ7hfsHwo+6ihSH275bjhWrkppkseIYp78ZjilFGqHPCc1y0dndlvsVNZP+Oo
BtE+g46bjaDSn14OlEeHttlGKuZA3UJr/J9mC6cGyWK/Td18l1EetMerKhv3UyNOgJY822fqdhj5
2LEh1/mHeWhnp6+CcstU4ipElBDF0LyToj5f2F3GaQyvt5m8a7bUlYAT7NmifbV110+USWDUqjqV
HSJjv2OkeS2zjpWTiIsd4po1RkxOWgdfL4OIGt9gJ4c9KiaxebEDMoc8PLnLcovUT9YfOcgAqaxP
6VYyHDEAmLSsIedKvBZ4MiYNsxGLc7U8M8PovBu6+75pNwFZoZaujDUp30JHVMPT5s2pmSDPZsx1
jh3vXDmZX5zjr1R55wEgcjmhXandRbVfIbsKMKdffX2Q4lI938bed0LD1B3XCXorZY01gICgmFJa
KBbQoCTF6KKG1gHhqc+ianrZfvyIOtaIjcYyoh4CYSXsECOMSbH8/CzzwraEP7ilYu0euvK3ZpOZ
ErP30nHT4ME9dFzz48PKobsErHNUP1LnnPZt7iLSNpYEnsZFgD3eKwj6mgJRtlsSOt/I7o/ADvUp
Nr2E8QuCXZ3xwbpuanf2kd2yHKrRWJOK7bvidDFo6vP9MyUZxt2tghBcVsBfPgcZiORpmC7VbGA2
FUlxYGqUu18FUYXHvZSgjnWSNoaQWHxhl3I39yPuIlnmtREDrfqJ1X4xYessinIcFzAtL1V/6BN6
OCr3+A9xpxvr56eC4XHE1RdzgXvKy2AIg+xIlKIbaWjsYDvEjGvtCm9K8aOcNqJGANFtj7ZLAmGO
QyZ2wbW4F9i4MB2hVe1if31dPdzW2Wzrz65rEzZxv+eo1f2P/FzMWv8nWLZbqhW4ZdrILDgDZmxJ
0R7gs3w/y0QI8TrK73Yfkt0oexILbtZfwOkDz6f3p1nrs09FbhFu4VPTqtVBbD0x0Fdsn9pt15zz
ep4kRQycci1i2aCe5GR+qDTI7O3ElHboVmvyNimN/4EhxT/LXglae+RQhG8k4hx7i/jpLzG3eJpM
vA2MxK1sXxxwZc9nDmX12n+dnuRHJfNkcDtHmvRbpGK7Zp7C9wLtOYVKspa8HLB2sR0jTa9yauSf
q51bToQQEjJXX6KrooGMpq0fWO/xu4Ovm9j3ffZQ9NmY9pSd6uTFO028mYbAC1NiE7fu4WdY6tcO
Hu/Qql+SCGqjEFgykQktLxqibeKjDWT929jXsOo51GTdam/aiSLWeEDVOGGHr5BTQmnLUzJLlCZQ
tpGKsfTSfxL7AANpkUNAxZau8JbiqACPT7RRe9gCD1Pz+iE7pO3U4y/G6LLANT3xFTFG/xXGF4Ps
2jyoHoYMW7185C/DlpFhS2BwKGAWuQ16m9p6cLr6Uvz9seuQWfjR73y2Yk9xOXEoUdzMpVxPr4UH
R/H+bcHjvjjDTerNGn1Us9Zu9r54OCTXo1/tVTrLGHBU4OhzCjgkZq/Jmq6eNM4rbDXrvzX2HMF8
qVR6khj291EeLr8bdGgUprKCpHTChDO95K5D+EnCivYC5pr6q6lpHsO4WYQUk9hiOneKgRErkJKc
SnqhdJe4UM5u8mTT8zF8+BiPJUJ4Kn9xm59b+eBy5QA8lKCwUV9PtbBBz7l+jbv5e4P5L2EBjtb4
SECWOFEXLnjhkfCVofBUTJa9/KUHtmE8qnr6LmA7ztrmbQWTd2y/2upSZ6iWNNdlGtQtYXa6fo5V
sPOJDLBN7CUUd4SSn3lOdEVjolG6it4KxrHDHtlHO4ATkJECN4Mux6xOhH+IHxjI9dAurt+pIUTd
/cQk+KB3nkVAuWzQ3LAkWaysqdywITzpTYg3nlMTP6iqJDuqUsWxitR00ew1rrOJxI1mhO4rqHdn
ge9txneOovW2IkeoGIrZkqQ5cMI+Fg4A42KeGGhr1YLMs7o1zstpZWXxCuYUvl2qHA7GeqA7OmeV
QstUsL4gwdJ9F5NCtuNWaJ6ZwIBo8rPqxMZZ24OSB35yZcjxrCxQBMRvPEmTU9bLEaIKutTHtp5u
R7S1je5/aV3l3CYgOFYXDveNaGVCWtwCNXHBn98ySzV75nZegy0OZzTc0n48O6CaYxPithGPM43Z
FBSB5D22cTwSqy4y8UyL8mXyzCg3lTmPdQtMbj/hDRXHOm8iTl7llfOu38PHLj1HcLozHfy8A0Ay
vB7TgY/y81oNeyyWphWHDLeMW0h27t444qNu2RJOptq+yvVvbSIpPLS4kfEI2ZkV0hDOiu31xGb/
tFwXDS2wUgOkdWdBPtUrC3eyxB3b850iPdS6pC3J+Jt/iRa1IaON4UsAbSd1ctAbglhrUgPSqRku
pH56QJ6SBr/SoED/6PJS8Ogg0NUId9LWtZcj88qOxrVvuTBdvTiUMjnGM4BDrv2gg93aXMFbZcHl
dhxkz5m0orjx86AuelhSecJh2B6G4MjG1+JqBK1SgSeJ8djNBean5nhJTiUKP4RIuZglrfrc3HMs
Y2YlvgXYIuBYsmcg7fdEQK1dcpItPYC+za163wpzd00RKXwSx9JvsRHdVFN4ursDFqGOY5e5Xzfi
xDnbqdFDUM186S7YvdlgecT2uCgT7v7DQwnTg1nixJA8HACc3sr6Z2pZYfKkiJmx7LdXIXp05Wxj
7cVF6Jl2/NAXpVmvSVG6UFJtKYq8fGlvIVhz8ypnAXd9Mrw6vKO3qaFS07y5Tsnl88S/rnzSmfgd
/7chq+ghOJZen5Y0SrIjXNnRUg26gX0n6ejEuUM2FduxjBTd2Ec4HeVEfwuWHOQiqRqOejLP+oMl
Ro1FoGMi0ZnPUIZz5AF99oPcjGsvb61/dX+g1T8lhF2WJVeT32UWv61rWzkbd5IP/bAl8v6Oem6r
SJ2bMFWxEmHk9NmLzVWAYH9RsUAkY1VUuz51/zLLC3ey/RVLpyRTgSJIWBsEx05XmLgUN7+c4jvD
AuuX81mhEmBj12jzOnvHr3gmvXSekgTlda6yWwEfANaFzc54sIR/QftkIWNA9CpVH80BGVQBCVYK
eeNgHCdzeoy+EuwjinzIstrwMGSE4jJBviA8UaEbvPE7+bCEGOQ9Syd8BtjfnwkNv86dXHwL/rdI
hrKcURjWMiJKEHKndofr81ouHFO7vy5mEhShvm7Afou/bQJ5h+ypo6uHRKUGqWGwMi8dcvxs3Xc2
uMrc0mz2+LZ6rHWG/MvoMX9Tuqmm+OGDijjZpY7tviz7cD6mvxtkS3vS7RTVERHDw9MsW5zxQ583
TBFBHba9kLgmINFPPqWuamZ2p/yna78d4zd16IEs5vGXcAKROq5d+r6e8qPSCuMO0hq9M/iEQdEl
MnFjgNjlhhfmwcaoQefBUQ8ggNd/i/0HVY7c/mTS0sIORjJMAGNrHj8JSErb23aKMShuzr9UxnKp
Sohwq4MEbf6NrzmfUm+hB3zvxq6Bi90Z2eTO1ViDwjYOwco/9gys2bFAIdSgKYRT3Munp7N9K/em
Ay6k4plBwqrCwn96K1Q+Kbpr2fxapV+7mgkSynLsJLpz5rqaH4hsRMA3IrG5jTcLEzQqnYAQWZIl
TvuxkI5/jSn2Vi/HKCxj6VFScBRCqoC4gM7qzWdjRVHMJDALexWgHXr4BYwGWURGxw8dwOJInNrx
jAvUN/nev1ki5XS4oEtsimfrHiRs7k/NM16AoqCHVGnWKq4DaRw2mV9ECKaYxGyj5FEDSJ8lZWp9
46DeyqM975uPGnx0HDyhiql261kh6xCQ7IB9a5tEzBuehzpgiRqgVl4KVT8OVZXivX4wU2av8zkn
F6by5XuGyx0I1pY92HVnFpTfhVAqerLeBUV1dr309TfMWFVo9TlLXcDzOHdmr1qRCMr9qsuM35lJ
I6mwCpbTSa5lQ+FirE5u6z5eR0jyVxt+Pk6dDJgR4YDZc6XDZlfqGUsE/gmDibRsNKw+49EP9opY
8SrZe+n/kPwBtdbvahJIEXwBizpF5QCjYrSH9h38IzC8A0EKZhPeViqceimFftE9IImZclv9BmST
PTsHDKtda2wLeYoICdDW/qlx7yCdmVmON+v8vqsxzWIOzdnNtkwn7FTZ06FiW83duWipm5FjxPgt
wuNd/HVYpdrG6dGjzMwft4AY3cKyHPh1LYYbpFEFkpR1MAc+w0nl7yKIAoLyIO0mnZd0AKyA7dDM
517Hq4GHoQRzeZC6gol88UfcnMi/5ccMNkaXnEFvDeDOEmdtbniPt7rZ1E175++ToYejSc/JPYLq
rUyAe5Wn/lU//Hq1/1qGzftsB1hK/9gaKziqcR2dt/YcNba/xUcVVPV1eUDnKe/5JqT6euUXXv6D
HHAO6cCnzYG1vdAegP33YScblWD8tkBNO+bmzY7hGuPGGmTjtb6TeLkkAkRStkLvRn/4Y5J4fzDU
jgdxdEgYmdeJSxDyPubKIL+aplq7XuYRW+PUnxc6zjU2uHKw3CanCoI6nG7IltLZvu6EhKF3sM3e
hGAb8eu8ksnP2bJdoV5ED7g21HP/JGRVpWQxw0o67y1b4aLXW9W6YCAziVXL6USkgKSQprzEDCAw
KYJ2b3Rz0qj7JLTrM83eotdLXjVlPf2VlsMWzrrgU5kkf0E1kEhKzb11uAVAkhVgSP9iIT0P7Ymj
ohZOcWtlm5ghI/OHtzP2ug5FUYdl4HlATkBgXEY6j29dpN1qqXTtbAfM5nfEhuB3nmwcT/Hm1SvD
RrrSe94d79YOTK5TMs6OE7WZwoVqNLZUf6UioAQiEsfTWKtxlOCu+iAtqTj3Z2mWNni08fvJ6cTK
4EABoDThYK+XGQ0P++Eoa8XJMdV9ctM4bbxqRncNxju9fcMPiSlTsErb8am8lOhxwUDYsXIKhnS5
lpC1jyzf2J7P+oRjCYJ+Dw3EnR+UYo1fNjpGIiDD6rqM121Y2KBAm5ZN4B3R1fmo7gRCCG7GIHhC
6HlxwvgnORGSJJX67f7yZUy2uxQSJihHA7XaRyeUmVAh5k3SgFyzMvsFlVltSr2PMi4TPxu158qf
2qJr5NK/ClCPw5gmUKRlAKGfR7EKSC6uXFmTEAaOmzpU/vV751cuGWZm1yqcpsiW26pXBqkQ6mHP
a5zgJdWu159czxIX6GO5Y9QxngpFbfb/N9kXGodsger/CNsY6SS4sW+GHRcWVjxWH4LE4hfdo9V8
j4OePPo2M61T0ol70VUONabLW1+to3DZnuS9qIzizJot3PFsyLX76t69qRYDcllXco8xEJu97rvl
/FV6aQGxyTNrf399u++H7qV3muGrii2ZYuR8f4Yjn2eKtJFniPClldd8bWJS0FLOlexJgZYLJnSq
s97Cb/vtmlwnsUeN+3W4blpo+RSSOktNkzqKtwdkP3oM7HYKIkrfk9sH4uRTwU8dd1CLn51VjDd+
RFUI5cYaikQ99kj0Au6tdl5yaEcDMn6qS+XwwqWg3h8ATq58o1VPPl63uI6UyiNi9MUOOaiNbnM2
zlVqieVbHYBhPqwxPXFnoz/5UuW+mmQKJ2NQA9JMMtADJLWThggrJH5Hww7sSJ/TlV5D4f+UTikP
S75p1JQuS0rerq2I0GdDJAu1/xZHO7zWlZyHhfCGwepwcudgv1S+Tf2A7jCUtrYAdZ4RHt52Mvft
MM9BHrt+tXUbDDmeB1wB5GVM53x0AfonEHQlG14og5YhaOByMfPUXCSN1Acnu8kxAkAKPCOBuA2I
qDo2iBtN69TPsGtO3+Xftg605hAKECBXG8UljjOvGVbY+0n6J0izB8g2lmEQGaEKBODWlWpvMK5j
Ot3PCdELzrGWGtZG6GeYTF6jfi0gbrO4oaVshYlIBeVBpwjyJ1CUXuQwNbG2XYBFBBv49pIoZhOs
R4btaTRqDnl2UK1rJN/LNbDuZvQukD/PcCArYj+P1ec5G18prQ6Q9SrtCUKKOFSLE2mR72QGO6rq
mbEWtSHzPeYqK3weMM+QNmhTl+NsiZ8S+4U2/g7EJF6wnI1sBxsZQGOCTCT6NoFTEvbfJt91KgkG
LvttozuJnBhGhVTgEkIZ00xavLLvOcki33ZAheSJfM+kVWXQ+U399cQ7GpuGhfL/gvQweoZcaX3B
3qfpu88RBWVXkPsNSbNrArXvUSB3Oo8af8vM4y9b3N0A/HBUQJQyPlwvJ5LXdhhFBbFdWOhAdGVH
rpdJx7SK8/p4EeR9y8FKwj/HDzG0mvzH3bYll0jjjPZBlUWeYQGZhDSDSRPe5Ju1vRGMmWxPPzKq
6LCKyl2VoV3097vcxZg4BvYyWx9dZnLabjcrtKWMyEhNTq+SmlNtf7oQgJQ50d2yzigLyK2D2BDm
oJk1kSvfOK49N9KGiPwWNID4Wiya1ZXHwwHrlKfRdveBkOooocuTfcTlDXQvAhNdN+BH/vAPePz4
kSls0lsAOxQCq6Vt80lXpsDGwLOdXf30fXisn9/j5P/wSDJsX4XSrC+LzuMs2OmEel0JQyf3f7ap
CaI8/ouOkxIB27rHhKBuAOLUu8yTM9OVwCF7HAKqAIcr/5tsY2F+g5qsGWjTMG2NFTbOkx4uZqTe
EGnnlB2IPoo2ddbwEbwrTyWHBDXisHePlVVT0flT0wazLrpDdhcyReumO07bv7YrwD0DqR/M7a/n
KBa4dAL0ZPR2OEiAjiPYSaPA/lZ23bE0MiPusvRG9jGYRAWtJXfI0FRS/VmbUzt/VT4kagH+ye9g
+g6GpluuxEF9+dUqX3CMi7qSDHTCfLXmGYEqP4urakuq2anIx8KQY3zBArt/s28zm+JIl6fMkt+7
MtjZjIDCkyAsiFhQ37tx3icC1cpop8nCHVZSMHglHkYHxEYIhiz8zuAYcVHbNjG64sD6Y/P1/E+D
NxtjGVYcZe2S7Sgl1Q+ppHjKSzn7XbWGaPN5veUEzZQPGfPUBfhb8+x1S0izAUkZNbeH0cFGJQTC
aA/uAov5IUyHIVq3AgP1iXr435d1ZiITzzoClYRNedH737S333REqVtkTi0ctW7PbXGqMUbNZc4+
wwo1FM+Y9mC8JIm0Qh2p0Bc6/DSuZThrKLGRW2MQ7+5OMvUVg53mHb8chhp/ZNapWzLqpFpClDmp
QMpRYbl7W5mEum/2usn5l42zrjNAv/sHCYiTQOB6x0TfEkf2MyJpSBbrcfUkixOijSyVUG3+ok8M
wkaoBOHy6459R2jStTfAtYwYcFUgcG5m0q7Qb7aqS1QE4OLpB5mawAGv9iZpOByuVW0Y3srWRHll
4FFNtmOMtFQuAszkUg6phBEP1QmRZAHCfOav0Q7IOUd8jUYI0kuQJMlWnyrswnuM0H155mTOxJ0Z
pFTjdKWXKK3GpEreXxZQ7FxitC4CESNNt1YFW4KVlFe3vdaaK71iHG6gG4v+G5QfF53JiXWxgUDK
Vv8WaMDqmD9kEwC6qnXIuCe7KvPkS5fNdb2MXxhJa+08b9TgazXgNQxMBoWjg34LolXQJsaLFKNY
woXzVnahyWU6r/Emv2iqRTTMYAVqR5AY1k4IbDU82Ma8f7x8Zp4Y89/IPWD4n8vsSZnISlyeFHKs
HdU8YY3aD3h1MDKTK8VS+dfm02xHAxPK/+i0a7L/tEQItF+dv6A16clzDDcn5KdRJCx5sVOFGVLD
Fgq3E0WR7zOFSzfrYo/3CuHu3vJ73Co623Bl3V3oxN1F4x7axS1OTb8BASmoUCvzotWj6q3iCquG
fanUza/Kpc9tVgCra+5sMHuRzMVRJpp8G699TpU/b3gAwLeOJgRZftfRe94zyIM60VSaSOKfV2mF
uHbG2p/dtntYHH+HVK8N6xkdYMhsF7Mxl1vXJrlgR6dGX8MlFhTegknLBzLLCRFWvvQsjoiuGLx5
h+/ShShjvt991dF2Wc4VbhKXbN9Zw4DBK55FSuPuy/9XPClfNbdoe0DBZR+yrNv0pnscReeOp8s0
hmziCBBOmsneq3M6AuReUAkeTMGRXChccnzTzv809yNUbfT1EiAEyGonYoqJj1nq4uJH72K2pxib
XcIbBRmC97Ma/MKG8qi0JG0STNhJ8uiIMnz1GMRxpmvgpDujnBBTQePdDnd6eCFBak2QPv/mEivD
XfETASz4vbz4vadFFlujvWcE5a/w4JMJ02BfyeGl4jx3jGMCVTCJ5uDb3/NzgDooPzSvjAB5Vn5T
9BoUP2JcPS5kHtO1rMpp0zUBtXLHVZpAkoo9m1mC4q7T9/XuXG80O0ZzwslZxafMeAZj26XjnMXc
MUuqEMjQTihlexraaHWGAtHd4G2/9gwKnekpqNOZ0sxbrTBw79ci5Jjp5U1fFP0yUobqO2m7SnUQ
2laxAUcgvejXw4XsroROlxv3rPZXPElwu31iaKfXdYykxB/i0xeNvR16OA1RUlP7H64Bfcf2csTa
QG2a1jJH/U4hqdTILM/0/a64MKywQrqgXqhOiZPYoR9ficrjbkg2Es9k/5DoielqZhHGfkRTjWFu
J0MMAFduXZrC+AmfG+ZGPJZk7//+YEttjybl/vITLN9ZfUXb7RCAKgP4nj6osW9rP7Bay1ZaIz7g
kThMfcHSQz6sTv1QZH+RssgpXXHeKPzIR1deixq1j9emPdb7In7/jdP8BZ/rFD+LJ+gdEBH4eLRW
oOHKZuF924b2RkJTITw5mthKKqz5uG4BxbWXkJbM8mgvVhTnAHZYffXUVWfrqGS+gOy3bhvpY/ZF
YNJGdPx9Rf+7ro6B5WPBafJmifqPahmgeEPqgS4LxsPQKECKbF69w6vFQbsZSy7QqynUzUBY7Kbu
MB6aRb9CQDnPD0J7WmZqJK7KZbWk45An8+QFeW6fnR5j2HmEQawE8gl76Azc/ZcKk+J1616BqIIR
QhFfevKgy+tjeT2sUSPXByWSjJDxPzSvUaTLyUyHChUuwbTL6CaSOAR4LnrXpDorsBn8GKf18CeV
jHjs+5UvVNbuxVsvn/C5+PSuoFjuJXlKoxZwrLaRrXFzyI2tugb7FQe8TorUf6NIPW8Uq0SEi3w2
uboY5UoTrnOK1nA6fFjaZzSOmwRjpBb9FLBG3U+MNAxs7ftUu2VGeXiPMvfRcfabz3YGeJchDT8v
csVQThY4HkBz4XdTyUrfepoYZAIFLOlCVML3iGATNBkkbZnWGiSH5IVBgkaacvLD3S/CNyvL9DjZ
HrPb789PQuMrWfgMBcCZX8oE0/a1rVoLwJNv2CBKVL9EsE4R7TSk1FsHVnEI1ciHTrEoXSpBkNxy
NEbik24Asyj+e93WwzwvvwZylWCAKYKjxyESxuxPf58LYM30CUuSYuETxxnlUQNm8Mzyanrs9fM7
FV4vxRkVpluDbrpnHkIqfih2vG8r3xmHLaK9DnwZvuVqHinx7nrzy2GAfE+DmGomHVbAcUGerEuC
euSYYXMGcHwIp1najLeXmLmcYxuSV3RJJGv47jJogLtqKLVicsUHRVDivnGUzHyoIRKT35JKGXUe
5KMPlA8FH3LbaZAFMylMtv4DIv7fKpL1mF7InMJXJ+LWb/q3wNGUwr2RxEoM23gHS1o5fPUMUwN5
AUxv/LHUNmKY8Neq0g4toG3A/howxcGoq/M2l1rQcYMsm7jwRloWMoQP3DbT4efjX2T5AHt4VILK
Um/8xqdKk4x6232E7Grb2W6F41XvMCQAfFT9XdylFMSpvMwDkkh+P1YzctxPRRYeMfpeAKMVwhGd
f8B+FvRYjT/MWu7m9jkhyi0VSFCzBKXZXwUg69/EqU7UjOi3zOIjhjZjzwfPYXQfsOaKeOi4arCB
fhHdPchs2tPX3dbcLJFQEuUoJnPDXAXOX72XSet01/Xbz555Ill4UVM3u1SHI97UNev34GvF33CH
iotioh4OZl4iigL0By2nzqXZL/C09boNQ9pOPi5xt4esh1pXkn9N5QMnMo5pVRfNY80adCr0In5D
X6381Nm2/Bl/+CkzXE2/paRB/xf4UJJGtHk5yam+7tpVELY801squ8C9zL7FeRj1NMNXG7ixeCTc
fTtEY9LF40uXUggTwaX6d333AaCl7YPyfDZ9X3Q+nbra9WYz7oX8O3/Q/SMDgldYZ4pMYNZJtrYv
17TRHZXzBj9L4MpS6FRVGXMk6AeKmZgD2ghowgJ7LB6dHMFCkqOfFxMhXDGQ00N+vnBAklyBDqnX
J9gqJKoVuhSQRhJ0FSzQ7MW110m9jfnvqfGQf7HJRWtUYRkk3I4pE/pT3U2vesa5RlmFTyWDOxJt
alZgrIUoA5qwRJG1aUvc/frJZ9NMIM6Kr2LmgvyU7MtdcnVzqV57yS8O1Pf1KomuvB1RckR34c6h
fBq8CGJ79qJwzQDW8vSoUvIYuBq0lolNX01ZyDkU2ewIrQzlINB2wDJgG7i8qtyILVrXrcf7ZyDT
LIybty14NGhA5BMJq+NqDA/GGO9zZXZ9rlBjz9s36d1gbPr7GlaSGJwAPWXWK23pxmLW0J0DEWMW
eFMuBzmc6xSMa8dIA2VV4OSpwgLhtmZhqi+LDCB+Ic/TY47zys3Y29uuLTTfjRxbFuhV4gE/InVi
wFBzNp5cSpEOe01SCmGMdfzzFEch66ZMWphu38WxW4hm+fXres3KEZKQ6DOvBXJKcPm/BSrWjsro
dqSmGGNey//zxGX93/pfsygTAB0xmeQtaPJIz84zulyQgeXECkUrbYMTZPuNghes0GDmMzs0a74n
dJHhCrnu0WVNrlV5YaoJZwgz1BqY7sIm5Ybgqx0e4qVOA3G4EVLhALFHM8eAYNHpuqvXWZgrBdDc
xbv2ebGRVijvt7ojXY9c2Ra5q3YQcWesefnzU09x0LR/KhEK3JgMQQZVgyCecKONTU66+XEQpOCW
jJi4vu9nWPximgxXpRgRA2QSW50detAq1T1lUFZI8ikMeiKexvq3sWWh1LUjnbrWh7r32d8dfDDM
aAee3U14PECUj4i83Ov3EnmDnH0Qq1MQuAwF0avWkIZEnhifMN2JzfwnJvhG16zBhFCEHkOK1qtB
BLAR9iY5kcc+ouFgu+2jtv/oYawiIvXdRgS19FC+OHHBZkIY15LrtyBGcXGgy7YKFfUWZ1DemEtE
MJct31gAYfz+51EkMHSBHLbPKE8vb1zXCiTEoxt1kiYz7wwfLxTjkJq9iGHqMzkZ0pmUeKHB7xD9
xkkrJqAeQiBaz7+zwtqMQclpaLL68cIYnmm5pnUeLGtVU5OXrvqhnqcZc5al0LsxaKK1aMrHIkDM
mh1cW/CymiJVT0rD9EImOsuCVR0uqbjVpywbD9xZxGFmvjX3dMO4PrZv1v5dwn3TXEPommY2Ov6a
k1D6c7YOaGNLgGIpDdtWvCS7BKJaS5+hIUfd0lRcXfnzKgFupJWkNIoZZJDLAOKJ3yIhDA1aGIJt
Bi9yDccMJzttapjSwSyrl+pTpLkGYZOLNPC8K2f7NrnJ6OIA2cPVcqg64rVE9d6wbdw9AtP3wXQx
nTlvSFk+/R8ujRUKJ5j6FlZ6dpGXUUpNLiv8AttFvBZ542ApmCjroFt/srs2klYjy2W6X85HyNNX
N7yUaRpjB4S61nwQBqyCx670xEGyNQrLggStTgoU32IKC85EvXcLbNkJMEViIiLKhQ0RfnvbnfCV
6DlId92hWZ6zsF0yExXeuBjek6FlxnesVGC8QZLw8fg5f0naP0OKQQ+gYitHhWMZEyNiELf8xfO8
cWuF3THj4b2VzxNR9SyDBXp3woCH5nJw/WYjr09enB1BTIYkVi2G/oSnZJ7Yhc6zyZ9ZrCYcRUB3
CtX/iZFuj7LoFrSnBiGOKExzzgSGLJc71agReoAzf8V1Aj+0vMgUf0bzRTSZ2cw7O6jiAsNCbIoq
J4wRXuulVYQ9CTxeHzGgwAbDidiUKhHg7my2QR2fHPdZELCIZR2in7XwrDsfF4j+Z3b6qrShTfk4
EMxfwVdcz5mgX4i54myr8bRkRnFSTOOF885/1qZT/qan/rreFutMCg8C5gzBkGUfvuxdFD968y3T
nG/BMPwn/2o8lM5LztBZTtpxIW3cjitzagGRVenRqXAGoshfw54deBIY2Pc3QGqC6XdGr0aMR//l
zNhfaSB2ZWiSAsVBMNO5SyWpjoHt4OTLsvjPywzRzadVanWCTUQluWAwf8kBObaJplt2IzkrAiou
G/10GlD90/reBUuGDj5Pj8QFywF+d98pCZyg2HHbaIN4h257eeibizxYnsl/rLh3ngYvFEPlqn6A
j8tNE3J9hl0K15t6IsPCLrlwRTh6nWzr9kdhExjiMimi33GkF5/Es8McF2bq77uE64S1laurYcog
agawFn29KmH5ky8qhh2MssrLNrYDZDSD7271pZXr9dNvnit3wRD8TcDvlOFV4xV1Lui4mL1227Lt
QwV78fOPKaMu2fd+FdC+Yy9F/KLRdhTjg0GhgUjTZv3bBYOdF8i+uG7oGSQdvubHWhEcK3onl3oY
gBGeuX/eeqJC8+rHSGtjqpWz7ZwY2VmhYU7AJjnZboz9hduzD5a2sO1Km8rULeClfdEh7snGDSq/
77JdN8eZyzw+JeXX8G6PYRD7yKjMizjyFwu8TQw2o6iVAgIvMgEHViXha3rRvb9GYPAFJUJgZKJB
oC5VidBfG2WoWEtU7sVAy34sHhOxI4jNgLMS3aDwYUZDJ6U7AOt4J/OKP82b2vXJbkkffpMw/D4z
PTNNoxsluM3M75PpZP1GEYtKHMeRlP5sM1Xzeox9YE8XLuVMFAHU2rCR3pQHQW5wXsbD9Pj8wucZ
9sphcUU/yNqv7CMLHP98DLz0xQ1raxv7lOUci4D9YvlqzIdVz1j7JufLi46ZcV2uIQwS8iJ3jItu
hClejgxdOvSltQvlnjMzCfy5yvHbPGdWznfz9TvHv96okrd1ay9RR6uDmy9PRpgq/2SeD6ICKA8I
qqhjvaKhHZg8q5plJVrPsOYcpbhmBqr4A2jZWb1cKAUN+D2JmghSShzdJPRPG9deZBDKudmS/D9M
iGWJjn/53hZBxK6PFB+UYu7HYNOs3IR1A2+1qfJyLNi4YDMMUFJNQ0rC14i/jG5hbn3vx22sezmy
VJwA3CExR1V77QHKR24iwZTCJpUDbjAP9zAGlJsSWgBjDR6sSNk66VcwRV6wypfHQOU52XcpzfoF
Ujc9+IlWvlvF1ZQaA9wJSFCpalDhwNwjx2EntjWBWKX6paA/xo8vorSE8IGY3jxvg5OIlUsewCKG
2WNcGJGh1sxz5A2ZhO7ZEE7M+yTa4+npUHuxOe4f+/XCRqVgyH5vMvLYAsuyhsYGUOuFX6G9PtNg
7MdSwfBX6pZBf5Rnmu8O9Xk1TqE/UNomTsdhnw2YdH7fibSPHQFIutYnsO6+2jKGZvvueQw2cphL
G00w6yPyd9qYWIFZGQC2H1yryclcbG29PHqx+zBHxucVR71ivZGPoqen7QI7MmPgQzJ/yrc0wLLu
2WNyl+XxiU5yT1q02r8Ku3CEaJW+zJr8x4GLlUxZdzLBpX6R2PkAluOoSlAy0zg7Xpw7lNJ7txCF
J2XyhpwvgSDBs8eVHFiY+8Fb5MqVbefObpWLdsAxEm9E0MfmL8o4DjkLoNHknqshpS4h4P8KJSZ2
Rb+cx1SICn3HuCVuQg8YeAadGNsQJ5WkdgHIh/xxH2iblKlqDE5QR52KvG+qSKumVkaLg8hwv2id
TaSrtzZq0cCYRbuG5Og+rQia9GBA+X5ghXOz0XFn77uQ9VSWkFgHKbQu0y6ZeIbYPj8FgeNK2Wx0
oZJrzIDdL0ZgvOSSGknPMMr38yfiGSZlaKsBPvRToaZW1XHAomaLjXwY4hNph8/TcbF5A5EuD9Ss
vKJKHrkcEQOBtExu8ajA2wKBs0jUlHuLfgU2pKqRdu1qlxAByNISI0odxECNlKS+9J+rsgWByyDz
YbU8DOPu3OpnNLnop+IwNLrlg3nItz6vy+HI06T8d2BE4J/JRwExX4xCiHewfhgGawAn1E/ExBGC
zsXzZqEetqLZiGpT/IZDrQb2kFVTdQ8QXitnPP1vF5FirjKcl8pIElzH7ycOBE7nPq0/v/drQh3b
dvdlo4AVnqO+DmXF9c2O0Mf4Etv+hSrqwWm2OTPxvlb28j//76RPmQm77k1kY0zLlDiS8fJG/EjD
Vl3fo3W+wnoIhA1s1zh8OrSqthqbuuMYNG5rps2PL3JbS2IJpaw6kN7SlghVIX59YBzu/toPdqTo
UYdLUG5eLcm4bMcxDlbPcthqe2fJ7SNTQgnZtUe4YvqcwOvJhmtYKR6dbPRETCROHzMQ83nu4am+
lTQEEcAGdH2hZ0N6CCqWRWht60qiNU181S3vbsF+3ux8I+cSAAIpsZKOvWKSwEnCU8uo0wQLp/K7
7jh13PgHDpXYLNpX5gvV4FnFNRtbWEiZP/Pdog84a5hKKoE/C4k36b3yHOIkyEGtbvF48F3kqLht
8Y26SxRu2CA4UbRd9iPZ2+rRvRqhq/TBPSSll/od7zvt+wTcJbjOUVSxBS/E4K3+9u6lUmmeOQ45
gN9AUmuHv4ll51jgK55gvOEsZnpCZb6zHyiQm1Hi1O80asbFOuH9LDXbKcBJV9UKyt1X3QfcFhVI
s9cdfqN8Q0DeixdX1mO0as/+vUoLTN5aZQ6O0cCCZByIhT7o8QduL8x7jVAiqsBHH6mhmjEtG9ug
qB4UXie3vlKkDowEpWS/o0AXn4LnQgrIWk4/3MBtI6ohmDB2Dg//+kWoYQphvMEYadP5Gu1rTf5D
bmuqFQrUbi+TWGWogE0fWonpcaZLmLAAdB9xmOm3PIWyIh48gHD+PV6U1WerRtusRekGrn/E+KTi
ajwaQYr5zfJAhL78kH6Wu946LE74enH2PiyNtb711zVJiLBGFtegaWGYRIuOt3uhAWJpGYSfwQlf
9NLA7a6jQ59+SGwmmrDiaha0/03ZNt/EbRbPDzTts+f6dCLv2vfPBgqZkZ64hZ5MwOWU8mR77kyd
t6YyLh8yKC7YkR+q2jbJYHVE5PpsO6qmEKdL60ccT18y+O+S9nZvxcsGSPtHPifMcqQN7p+6WaI/
AXbhFGWRwVSdIg5fMN6ehMrH20CFlkULSz6ceToDDQ4IOPM5c9dVVngDOVItZ4YpBD9/+tVHfLhV
9NoqdYdluyhf7mbiZhTGEYI1W4mW+jaFydrej58x5qrM1W+iCOx29oGMhRP76GxLklhLEhWj7jtE
rKCa31IjUsdxMSus9eIbafj1BVbLcA+bglPjLb10jNQWebTpPNuD8FLW4invmb1ODyHSJuzCxrvR
4ATMi2qfU6suLLqrVkQ+QRJGsPpkmEbz/OpJNtPl2SAT2UXhcuN5uyccRXJ0MJEX1Eyn4javu88c
iit1WVm/gbALfKaJKYcGo5tAY4dfwhEi/d81qy7YwRY6drl0wduoQNWT0fVLmtmeFHpxmGWw8TtS
o6gRcMThF0B/a1PoIcriV7ft4MgWuW6V6seY0Xo5iOsQ2FIT6zn737HfKCHPLyqtFjgW8aWiuF8d
cOF5omSYX78uwpbwtWfZFtZQC8BanhEf3lA9YRXiz5fd2LCXMkuP+/cpcT2x363Pta6rfU3S1oki
+A19xkhraERX1UKYi4NTlBUolAQYC0DPOzid9RPbNF5FY45ujWIywPRHtjegf8nfpmwqsTS8CY2+
Bljhht3nJNTcaKGhaZYXRjvTzEzSQXsoMlySotGMHli17szYwDUmRgBOO2KNEK1i5BjQdZWHX+u0
iV5b45quw/GRF8ci2Y+btFhQBYvnvdXUQeCzELNdG2kAPtxyvDbW9ETLdItJBZuVzr/1l255Lpit
VpRm0kmcJdYhWJ+cPjZ3wJZhjojWqUl1uW/uFnBJbB5mocRfWRb0GuSSOA5tBmFHhGNUV2zqolcy
KFTntUrEcNDilrvQjWloydlbUs74XH77Ppit1Ueyl0oHCwSEaxPqCrYmkcSdgCgJkff5Xb6rEfT4
GcK9oc1GxbPXQAfoMfy8g4Fl4NihsTpKJZaQ7zmw3/l0pH2ajE8y7cwMtrODkSh64vADmAUHa7G5
zY2Ek2rNHygJHbyAW78LzBp5+UBrIcgU/hTKd1XOvh6WD8jH/86UBNSbp9AveEnQdmL1AdpdoK43
eNrjzTBgcgsYuCgqyKzOwYoi2O/CQk96VcvH8XeFFpPm02px9h05pxfnKdjgHNy3qrujMXhNq178
uSjUjV794i4915vJQI99sD2GjNux2hBUnEkO4mh1m8W25DNeLHwPJ7zjgptM+w2a7ABn2lacX6eS
WVFR/bL4AAstTdg/Awl0WsiJNZ6TLaOJ5aNf814rUhrSU5Ph5C2ll4j7iJ9CQomoL4+cCDTqayOc
YxkBavr1vsyelicLQKfr9q/gP9USIuI/N/MgGiqTNuOMR8zd9Ipab+17iMtmrP4s1SI2QV0P7aMx
nUXuk/qaLtMP2Sveap1bNli0zGB4GN8fNzeW17VU10v/0mwpjqe8+jsdxl3n9rXLXnLjmlIL8pJ1
tzik6UFSxUyxzs4w29RJvzO66pnu+1gVjPfhMBjb4qtXFQhoWJtHSGpOI5SgcL46ld8bCmUmDfKU
1CcfVOZyWo4SWa84i0YyY2PQ9VnVK0BfIJuMoj2SLqtzB37/oscTv3FwmxWHVLl+qCsapX4gSqUk
iY8+0wnFqZXhj5pgCPEpIKxi4C1iDPXEXtxddRWV2PCcBDGBqzqtgrKtbJJXFytdqmdmxGQZf+LG
cBSq0uL3NqFIef19Yfc7eyJSnlJHDcLZ8hj6nRGyPK8VG5J5SreOhgj9ThR6UqIrnqEB074TMgXa
zD3pt4euSifXkXEPXxxgdLEd4vZgzdIpUH0Yi4jQEDObrWWkW8z3GgAXdeib4Mqs5+GStNzUHqTC
P6CgVPx5QLq3J0m0jHyEK53urE7+nqDEdOSJwS4siBUrby6kiJGLKEAzXy2LXzxm59DEY5iVk80J
XCDPcucpBYZ5fJnUWLmrmxwfjTUYV+8s4o2o0gPM35h8T+5A7PYj7uiHNHkJdzXVTyAJeSSkY4GG
jDSRasc1qQdGjiEBDlp9YjTUqvTpmxRUNrotx+zNrZFd/73Qt+h/WHrqen77y3XIJkqX1PmA5yrs
d0763Z/m//OiCO5RDyZ2vxKx/HzztQ8jk/WoTpjYLvRkUBFCo5MBraWCSNpryt4Wcr70yuuPsiAo
vzY2AWAZXKBRXjEA+0cV2l6kXtvAMdeZUPvZuRexJJeaMvuaAXf3zvUsBMO5MpuMFMWWygALDTQr
R/vq4tlzCrXx8DelJqfOHc/gLF8ruyxM59UUQTEeb/ya2LNllk3zOfZ+MwjtKo9z22dZI24LdXFV
FB+qlmfy/B0y33mEmkgZurCfe00Of4U7BDfva3wtMiR0JSVYnj0QYDiL946ASuuFl9q03OErBpVW
xj+WUQj5Z3DPwpCwsTCUu+O5Y62jfztpzfCcxEolSre7uB62oRv5Zna4emiVjLYuxpaYp/ddva0h
EzV41ADNwYW9Z5GHrmpdu6iXA4v08wPSTgv8OTbR9dW3ZN/T9iDfM5k6YLvOww+38Z4mNnHmKuyr
ManUoUwF6bC5T20LhzgPLVVMAnIaxh5tmfT/Wf7raKEkUoWdzzVr4sBC6wVISl8J6SVIz0B5ofwx
kcrV6EUQzs2Qna+b4V+YJkEGpTEA7zN265XDtgXaSyltfV8toJEop8+h0p3sDdFM2THx58CnQlOr
mj//hHzP1DlM8xel/uTRF3yslVWFBA3iTdWplOA3FnaJ88kmvpv8tdN8T68KrAJ3E4tTyPpuuS9z
EiyXhX/nbD43dYpiPk1fY5R0+bifZkBPETiRSrbTpFpo5DdG4hlnX7X4j9i90815eImpfUAW7xqv
83dl6viPjyzZAung/tfVtn9AwBVAPB0X9emYaIYbu6h96tX5QdDkyGw3M+VtC/2sd0lIzf9aSwYn
BPeB3Yhr79bqJypDYLpRIUHDBJpMX6whgwRohVVBfm0BScPzbmpgT8vM0jdsFjcqJT//i+byyUlA
xSRpqr7bbdoiRinvpBGGLzNCdUl5E1bZ2hf1n+W9/IuI9AZNNqS/bR+7qOWdk///Fu3y4sTrAsV4
OmOXhjJ2gJsU5DZPc8icbOl27m2Mde0MDe8VbKwWymfVK6lGKYbpBXQT6bj1s80ULJebXkSYnzKf
P8T7aortHT+nsLQEfCzWKZlBbfHiBB81I8oR35NeGuHprdchiqEiYsNJKT4vjuOi+yK5AaKRpnD3
JmKK3/qzbSDPYIAF72H9XugZUESUbikxkRHTiKlRERWwr21BVxkCNPHUy7COQfeYQymlERBEQZcj
e5E+jQ+zH8RctB4lG9RwpDUBkD8IhmA2SBIWZN7iCVO5Wctxx9MLqdD0ObEIWOY+grQ+QIyRaGUd
6oHq3jnPu6WePBkJeSJfNhtF7LD1W6TsbXnLv9CGjA72oX/P/+lN1BC4K2ifvsoa/jbYkdZKLZFp
Zyffskmi+4xpOjvcDhIdwPNBMMjGrFjysQqjTuYnJ+8bx8WRUG9jTH0UiV26cSB1mnt03UHYbvox
eR1i7QSBBixCl4SDa9WHk3uE4KyCBj2bPYNHQO9mFYDYvUv66s4azEN9bNNgLUtvUlfEJzhhM8NO
IaJosnXdLVFBISYQ0ACVQxNbpiN9NAOunDs6No3YBQhT924x6ovDEenmxse8RlA6RfNwG9o58+Yt
x2XkzPqSy27ODkJEJ5i7pYGSVj7bzdqbDdXH7Z5gOPiwXl5vFeO0Sx/6L9QtvJf6jMnu8Ccfpc5J
t72nSmf4l9o8xyOV9sibcS2WWoKBOKCtSnL+z1HixTEJkqZ5NHgM0VFTzzPNNI+k2XTQRHQRkx/u
H1l5CgHdd0bU9f98uC5pk8HQqMRzU8TcH4ZR+fugfuuZIXqqO7PZGdJHgAkWisg6y8UbwSJLVHv+
Bekq1pD16C0xuQ7EQpQfviCWNTjQsSej6c+7EQWpL6uEWt9b+P5HGQYNzYLaefgLXKc1z/M88g+c
NpUjQRXLo+czB1pvIz8awiBjWpCnPHL7Nvk4oFzrd+SwZlxKU6kQBdU87x/b5u0qhaFbi0fagmAx
rnffrRzeXnMihsbOpbq0oG3OtghVB7x6botBTQ2WnhMxqWuHBFl+FUoMYFfjAwfAMdrGvDebfs3L
26b5EDebiuYQ0f5rqXNKqKVo17Z0alCaedXGRN4QOPyYX60QthYjfHG2DbwK1fCjeBL0qi/BG8c8
IH3vFccx5HuaAoUcXiVyjZ32MsfCUTFAf3uGY0JjbbY+wu+BiVesYbb8GCRc+ajZHNEIpCcypoF5
oKi1IBQM6g8T9yHy0uzQ1sJMajSY8AXNM9+9xx1EDIpTHT8jnyGIMNIXGvUArmQO/5hLEmtm5PW2
acmTnyy8jc1LT6D+Hh4+AB9PSYagUf7IwT3X2xlyX8FmXsyFYbVHDgB0J4lutARHO4EzXmxC4nzz
Nk2XrMq+NI9uHGYFti+YYcE85yroGNy/BQYcFcyHN9MRJHSxCQqphsKg50GDr6YauVghWOqjACMZ
7nL8rOvPfUKww7B5WfVIBDESq9tmqotmy9/jWDj7S9PO5HIYdWosf/9TquLWKkPEoYApuscKalp+
+j12crb3AYY87voAJfRMShWrP+sqX0/zL4k4Vp9edRgteYiJx+Y63OxDbmK5pzCfU4iT6y+AQuOA
QWQ/DjhyoWBJSHJvRLTAW/RxPZMUmiTiT0+mf0V32KnEbEr8jit+rkHNjLm2oeZVdB93no6uWXwn
Nz45x5OnZxXZ7c60QFipb9J/VUW26ip/ZY7TSQel9Gn8QaAHWazJx6Ps/+hQcVmcsV5bSbeJw5Ng
NX6QWbkvw6EONdcP8ObaFmiTq3z47U7VBggyVZYrcRGb5I14e+YNAZhN8Fh88ezy2Tyzx2HiPUjd
BuU/AK28Yn0ucWHPmuuS69zT06dwG9KSzAUzMjq54FIwjTlfQ9p62vqeBFPzbCpF7Yoqfh467Nuk
yEYyidZDKOGvHDJ1CUcrX1fktZvBFodnQK4Udan8TIFwMl6YB8kpkKBJdbaHwEAExyplQry202bK
+kTzYa3YCTEIug7lMJDgV1aB1Hicn0mk6qruXfWQ2lrlSZKZcRkQLGwrInQ6azneF5tNy7oeQZ3w
O861moczsr99dOdp/LqxFAtLoZNzv56Rfxf6H00Bk7euNbaYIzoaaMTMDujPCzfMJjlAgewCPAAg
XGalMBpCVtbiiTD4U2+QvScCNc5tFBu/aCqAZNi1/bLJ/PQoRTBbHQcKaZQQMbkDIX2qOqlOQWWT
6v/2CR/I8ZxyAU4oWaNi9xgTt10XIPNFIrvYpnSu48SLaO41eynMChCLq+CB7VlW4Fd6kYEKr8EJ
Mgc1B3d3qVByoXlWDDBI/wrNl2zu1gd+G3/GqZ/GZfum9NBBMD7OlEIQ/Me+QTqmBhATl6Uebj7P
aUhrSQpr6cGEUvZHB2V14EcIHOeRQHvB0FtgLcRNBMdZFqnv4h4+sMZmVmT94Op1/PbURe9XwW66
R1Q4dY2TbLEfAv6C6NdX0cJ1E4TVhTZVEl4xO7KfoOhLhjeyywiR+EkUKI4ap++iH01UmtOp8yMj
uSDrdJojiSMyWpfrf2nhFmWRE74eqNiGyc9JnS0/0cMAfFNw+AAmn4fX/7P3tPnEvy1+EvXDQdJ3
lLRQxHTfrFZIan1ViD/pqB0ax9zcuUpZmdjrBhhBQwgaXJES8K75tWKAV1lf8NauCmOzGHM9D9Ux
qxiKKE4+KK7vKLC/qvL1O3+f8rZoIv6Nc26ie3d7VP7WtQ+rAj6hIAgfQZRd2M66i7jjmOYOUjEG
eBKSHe4XcyIHQ5ucmK2kiMPYAU/W9mKyZfIuT8c6YAK3FWGI5PtY4UFrgBIOwsOqG+j/E6DxSXSs
LxtgJt4X9YHHG06D/BQl2hhVEzm2EujqWRn+yIs0y3UW3ARXPoUKWNrzy+GKlBUVB4BdTx0gxrtw
ZzrHUEKxdMWX34JRnB3nan4yCi4EIka+olYk9uQgz2rlkJvpUwZI8Q7E5CSvZeZrOVKYkwdWyPwz
qkdL67G9q11WtulB4eraqBbefgYSWy12jGMCqepDkYelHpQMIh1vBeVEPHY50gnGvDL08tai8MyD
K2ronVpEt43R8gdMolNTypM2j9DU6xpupzaUblHOH3qPAu1TiYuYeX7lakR8NK7x4DX6jaO03nea
hExtNiGe9qZSnJN8+HXhQXPUsP8JwdjJDQRxTNXRuuBIkUqiMpt/ERah/9TT6XM8Imb+21JAR3A3
IRqKlgElpadnk6CeSocJGhHmQ2SaY90KzgpLjQG86/j/JChjbB/Xpgnvm10pjeQdkhNxdF7vTxgQ
nOgQ+4oXpxy4IwpjuthikFzBz1eLFYv3IVVYp/dkxlfCN7jtRYkRUnnBFEJkZH84Vr1zd3BxoZNi
p59SMo2h9TH1tlSmJlwTSgQ+4x7/RAvjhKJiIxHym6ZgndDSdjsSzbde99UPgeKk1eo4k8o6olEA
KAlbhoWZeupfMBm9x7qPi1AJla2J2Jzaw/GtbK4hxM1pAWFuDFf31lgKQihz9A2ZXl751/Uk2HA8
i8SRvQHLuDS/4Nv8+Za9OFCprM1kvae7re+42urdMQ9QdLmQlOF5ajc637quIjEVd6UxGuRvf5GS
1jfi8P0x3Mk5vCF6pZ2AF/SHEZ/jTbdYZhX5u0h66NyS9P9i+nOzQFHWwLkso3hVRkDcDyUmMxHW
4FoujQtpJ1UpZ21HozZV7woi8YYOKI0rQunVkanDE6CGxkGLbnnnb9ens/TyKrSv+CG9Dl86jYwI
yIEsc8Lwk2OQLP5zZlG/k48zpAotNVFRtoxMR2GxkNbKp/7hF8Vmgqvvm37vZogifPVn7c79WQtw
vHLq3vCNEzzt56NzwerjxwEWkjXPKWUIoGI4QRW2UtOkDishaA7U+cYdv4aswgmQ1C+plBYo5Hga
Qpv0a5+2kBMM8Ccy0DXtjK1Ra6D40jyeTm64Okd56l/N/sMU52tG3s/VyM5w1tb59QlCFKzHv9G9
E1KTSf8+7SKDtdsZ74zPjbsXgHoIQJiqAYp+a7Bsg1VxPwYH39ROnVsBhs7pCwTbsb6Y/qJyPXJN
KzXi9+zoYAJ31KdkrsW+h4wwAcvlkCzFuIpR6bdP1e4mgh7ywDGyCP3uTwEn3r/xw1KVXHcSraC2
ZdnkjfjVGc/wunLVkTaic0qdvm8X35DTBI+VhXF6oEtyuMf0Nrs1zyKLamneFhl0Zaw28SE0WBrc
V6kpQRl897kVFm7bkfwRhVCXoPzGAjTpGiOGfp3n7waHc6dgBRLBJ+A4ULQCGQS2lKEgE7WQrW58
XEQPikOfhQHTvOiGMnm4NVC9oTnrglZc8qnevJ4obbEAdYS9yxgtq2QWlWPm5lV8d4ORLTUDvrVK
pIQ2/0I4mFKlbp4QdoBSLjFBcg4gUUjh8TVhz5hQylWWpUltTLEqasMEapJRnlLw/Jubv+6PTQrD
6deU84OlyrElD5lyATeFKdveVNdE1VHbNDZSd7DyGMy3AyICk868oVeEj/I4cPOJXkmp24JXRW3f
8l4RGvMFScvHiqEwSkR12paHu2NoS0Qr+EtdSULLP4GI/Azb/G4bhE5A9FoFuszEGyhaFLOezrBT
rCgeozOI++AGMLoMZT2o/xH1ja7clN8nKs1D77XRRujkH4rSs3Zt03rFWarEO62U3aDZ2craXVY6
PcC6ZipHx8bmKoMW0EY3rzn6jN7KMGgYNjSc+rtt6EIIFRsE/3vPTx4wq5xC6k0W4N5Ka8uY+dn2
Gi84XGbHVQCjP65xiYDiRb80PMlemv/zcIfD3XpTxR/jIK0PRRF0OEMhwiAo0TXPGdkr34Bi+AkD
szBHX0ZRjP0d3qoHh65pPvhWQj+KF6qWIIXWXtYeol+tDYe5HGnnV2d6ajAeJNxS798ZkstQVlCg
poqKUiu8BZcFEYCQU8yJqfC0FI3l3xryQbsN2N+MAk//kXJfwHNmZNiom16qe0/YFMozVdQPmXHY
hWhns578ZtyX7dBzHrFcG+yZ8vBTWaicl8dGstVmenE6qvY3Rc14FtaiywFCe72BBm+zcApYaUSq
4esmLVktA2USwskX8FzgcmKsS0uIvP9T/5pb5/jgB1k6NRVKBVzq27CIic43c4FnjWQJRxuHzAZB
i++SfYrZmIqCxliO3txm6X9VfYN/pYawNt+eSsiHSKQvUZws3w34cD6KDbjSoaleawrhV8/JuoIC
OIP8l1ovPrNiy9bUxNiv8kkOxZr4UsZWUqZf7TR5tsw3viXk29626lNpN6cYTou+7x+vzS/GMZj7
puOepGHuSHhD8df+OLpAEkA2uTX6PAsXPnG7DJblE6XXP8H6yo2UxASFR5KSHSW1Y8ScE8jhBrSw
+KQiz9Ug8nVjvFE0u2e1+fcYRTz7vadYiLEX9W8iBaqOeBozCQ2BkDPrX4rrl0vbBPKwKLgeU8Wc
o1BKq35l58tkaKSKZHCNDI8UTssMmZwzFUolRBCr7nT9OkPw+gHWwJkSa7Edy4XFlAI2lvveFAc3
dgDSE7HmcBoVu+9DFf3/wwFar7P6E1TrbnHVQzgMslzEgGFPxHkbNhS8B7Eoi9wZgLnZErSlsXX7
xm4rBBfZ9S9xdqLXdjWqmEufUND3uWj3sihqTKbMIL+71A6KkOcaU3Tg5LETAlv8i0GKiRstNsMX
8LjBHLV7NdxSJyHQlLaKmBPA3q68g6FRmKyAfAzSezRLKJdXcDDS10yZ+kv9UHSbCGIu/yLjVYiB
wDg45aDHSbFCb6qh85JNP9KLd8MtFsns5y0SPBZdOvqGB3jPbBMlhnxnbwGTSQ4fVLUZKZKHP/dN
9801TThuyyxAJkXOLDDdBONKFu0TFnNpFkMcl5MYQ2rsAH7da/mCfXEWXgWzuUWqloLvzQEeoKoR
dz7hcJ6i1SFooPRfFtmZsq5QmN0+jxDCSCk2JPOjQy8Yxp2/sb6OwY08eVXT8qRv4uMe0YircHoT
DZDFtJ77xlGU9PFOXPYsC5S82waLgkemRb13Gi0xAW9i4idfCLjdt6hwtPpzQRRW0BRZEVzJMSIp
3tEcgJN1bRPuqB5WlFXKRRku3y78S4+5kSrMzUPkPhkaiA6ZkqbXmHnQEnmcr/RToWnlbidU4/1F
i/Yx8RPz8zRSlvPmty5HzNhRxY4serI2DY+Y/GTXyJJhIjua8EnOTCcPT6siC8a6Akrj3ZNz22sl
Ijw9/e+w1voLogRM5acSp9014NjKSVKwJB4ra6qtiKETx9s69VMQYjLXibVX4qypYFb1EBCLcefV
UMHwpL/pBp08L/EQ/gQvfjLapCUaTeli3WFkfojR6ZLJXIH5d5EM61by3e55DAS0RRnOYT7/1lal
xhzRbiR8PTYYdU5TURpZECOKar6GZMYWmWTObDE5ifQiiCua0HU2aD62nbRIPlLyG41fJgrA0N5j
69R9vRtdqo6BS7D3lmHME40CrMHHm5k8Pr5ovm18EsIGjT/su4EeiMca8c3dm9Lul3FscA2MDXjF
rbLgiadsiRjPQPlVu7OQiggvRUyQE83TUyqNDX1DP4PRK92KqnbpcRHKW4g6CUPL+lbXT3WGT1xk
z6GdSVw1uqeEqzHuTsWTYhFnWMY9rdVasgSJTCi9GvJf0VeY5LwKKppaM/W07U/R2+Pgusov3VhU
lnolbvh+k7j7FGnaPEf7FS5ENSt5kQsavmFFsSDO+3Mrcdbq7oKH4pwceg3FkNJQzfRj2hApzv7O
b+jhrv2xlK93rAv+SfiQqA/M0DOiF7A4Y4Ia/o7ZUT9vNCOykuD9bqkq0lkVuncenon1AKJaru8K
86OkmXPHNabhhARx5oAa/zEqOs394nYQwrwaM3jo6NkpPU3Oelhe3vKHar1F4pd1jUbf1Q0YT7Xq
blBxdU099v8raGTUPqSFuUWByyTiKRqGVMxAvCbzz/Nv7CnNdnqaslmWEzDm9kjuJYk6/t7d7krK
tZojBEnv9xLQxuEf0ycA+jDy7MaCLf4hzp3Mfss6Z9Bwe2zkT3mAyMWRVa3BASnC6EOYz3Wx8ZOj
YhGa+mkur8fYQwd+aqbC+HJtmZ/t2Y1MOFX23TILNveC1P2fI7LaYC8Qu2uQirQthBrKdFvvMzkX
h5WNH/8Psh+2s2hFNfOdqo0gCOh3NUYN5VeRehiLv/JABKeObTLh4FDLZosZ/BhQR0tu9rZVIpiB
MpH0yJmGNL0LAZF7McHw4n1XbSmnGwR6b5eFVOVITyPoIlA7Gmzx6No0S2TuZJkMqcyHGLoHckUa
Lgd4IVxkscWWsxuKl5H0Ea2LhXCyML7Dkfbcb3HX6/YqZaG1yAmjnfGq790aXz4HlbKR8GP9hapU
BPnnhirx9nrjI3pCe8Ri2ltVGZY+Dqg8+htsaKPYnhg3gVp+F559W6cAmeSBt665PVpiTLpyEOfY
BaKDl7d8i4wIAFBa9Yvl5bJbeNTLDs7SfOX3zB7wT9RYK8NfrvCJz2v7DuSt7yGiondIIBMC6WAW
NDgFFiUOAUKyCmyUVwBIGdEVaY5PxPCpoVD4PMUK/3ieMcNr6CZBcxssY2O1JXcDQeHCaBMl/GbS
gIZYKSZj0MhrPN087SrgNvmXRPBMp/NR/hlSwBxyuXclOH9ocjjSDKFutp3ZUGzGzZMn1abE/jjl
ETqdaM8l+HC45GlKzD3h/gop2TdBPM9JMUuls9FRZZiGOeN2DDcXX6JBmOiZcERg2bnHgDg7ClId
n1fCDLl0vElbmoTtOx3kuR6we9ARP2owQgnDPNPWKgpjEZlEf0nWDkf6FfmRW1sLbwVgfXraUDtS
BLY4fP5UfzbDDwHjxXsbOpUruQyebr+1yTQ5JYR/dPH0xoo9jh7VMgTeGJycgJs1zp5rRq5dhatn
J2jnJp6FQsT9X4o8BqbrLrjERouE7MbAAJW1rE0JPNcsrpqU1vqgPojvb/pfJSAZgD68/PggK93F
sYYavQHiCQvUxAqGAxe9PbYEStUMUluUeT6kz2ArCxyIWYAioi8OEV9uxa5wqMnpeevVjlbn3KFZ
tKgUofAQirs4eiKHIJh9j1h7lbWToyAsp+S1ChVBuUPNk8zulNj70R/6tnw52/CkbEFNjAlB+F21
sbFk0jOksKh9ericAQ72YS4El8JVD7uWeHxgME5lK59/oo1rMUOOUz3HG6uiwUMPoNXMkP9wfObr
XutNBUs6597D9285AtlST6PDSLsjc6fcF/e+PqOfjBKu0weblUXRZ4mb8iHqEFiuPz/cY1WQcLCy
63sjoyDXc+LCUxYcr9qpNZGNm2pJH52IEzADXV856hPbZyzI82RTyC/wKDszrNo9MgS19Xas7t8c
yJU+1x+KTgqw86BOtgx7SN9jgvMkrPbUA6sfgT79sAwZ6UbPDgCE2frrc7qXV4nN2D3HrBN0zd1e
jsuNxjg0L5ltv1npvMoHNSzO7FrXP8eMBTyInEChrRlPmNhwzr8O7tFopl4+tTmq0pXUFMEzSnlm
uUBEnrLHAweEMcLNWc+c1BOMfcMRTSH5nbepZeAf7DNy79cnU6Ad/bC/7vkpFKZBeBjPxs0CEKCN
6bFy599pDkYChWfFrNZs1cIvYefboStiE/kpXI+dzzqpImiXTftb6o5cw/n96It9vzDmOZaCPfE4
zf7KGEXuZ22MlY/LM/ew/Etdm4VPaen67r427dAosbGgsJ6AIK35HjlfPccJGESjA771c+XY4dpX
8k5AfyXjhvrs6idrXoJI2gBHcdPUuayK2VIBVRzBKPPml578tt3RGvSGsRjDf639aTBOY4zN7YEx
EkB/tcZThGCbVCRYkFNDkPuPK81BHN2WWZKH1bA39h+4v619N/7zG8G+OB0k2hIAZOLJVgX9iLg5
oZxQiIkC1Kdxj8JLE+Qrymic5FXdlG+iiUcpWzcSp0goN2ETY8WCrbNJjpKs9AnA++PmLQsMr0mM
KpVprR3g15rfQHUUFuG/j6VNdyubI7TRDviGgWuMLuwTEEwbyW/H0jgGGIlHNWLI1I37oHfGJVEI
bZ9b1mcgZxeQ5m72oU1dWy59t52EKt5yPvJ9qbyUTwp9+XA2d1A/n1q1oP7GA5HIubO+MbBVw8WP
zVF6DkCgeNLvHdlafyZ2lDAycTw7ncLBNt9P3AYkCpscrto+KBRgxMZ4hAwl4zggsQMQZQSP0sx0
4EoMLKCS7G+JgDQGxNEDCbQpHO6iHsytTMq+0IINIvK/ZHxEX79FEkgEuzbiMSB7Z2rInnlGPbbE
tukC72fbmcyqAn/oMunIbEd2ZfB9v3vsFHpQ5JdlxKq5+TxkbRUFX1YB54ggUUnWxRAw68LD8wFu
TcPrIvIXla0WWvGFVoi0R1x6QKbXFgkdxpSNFxSAAn+rIekOI2qU0138S4AQ8Gr51AJI+1tD+qtv
JkWK4uUfAuCTK/u4GTvBt+tusyqB2fiLLYRsljoXjjZGptxJyLUepERqEQZxw3a3pQnZ1rT8EpOq
Wy8tBjfoaSihE7yv08O5+6wi2bY1GywpnZp98nMLA9YYF7G6CRTt2dzaQpwfq62Pn9YWT5FBTg7V
vJPB1RdxHUwr6Gl/XBypFEscAdVp6udjJCm37bt72j6BeqGZ9z04GgFPWJl6HwC1OyTvifL7YbPL
zOjN68AGqJsTGlr0YJ48XcSRh991qOsBVZg4S0z5ZqPnDGxT+aA1NhU6q99MxOKOw+NTNiSjKDzh
1gZgLWErkRfdZA6ViCT53qEc7WVgFHC/9VJq8vKmSeauqALSgUabzPT9YH62pyDX7Gj9YeGRR6a/
WsHqcGhyboJpOCHW3hzqBFqGjmZRsp6Z9mOWEMcUApyaUYdoKyIWlPxIqrhvMyICFB+O0Spi+cKt
W+KLkYNNNUAwfkHwqS+kTVH8X98skBqOXojw2W0/UQJQQOVoIl6uCBz1Mgvt30HQU484HYbSIHUK
Ltg5XN4XtDQOHEVq3KYXOXNbfaOwfQ3cimnskAba5yyVTd7sAuDjF4hzcBDoa+tEnnGkacnz7yzr
IiMwZeHrW3qCcRmxztqXrlD76gYkatQ3CVHTun/9MQArNlc/JfrPnFa3NsViZ1sqTrOB9of8JSFt
HwdBrRlIh6DdKemsnX5pIY8BXtJ5UfzK4xLypXu4VVeHSaVEKeoNbefJ4Z02d0kyrivX3Y+FaNOx
aRc8PfzhCVt7/tdqy04bq3PuKhwROaC1l145KIns9gjP2QKBms9XJkPW7T6BuQJ3MNz1TUy75ToK
XtG1dDLLleh3rCQZnxUYXtqz5hlfUZBGJwZu+5vTrbOcz1f7TVCgQCTZ9Y/dH2peIn+EPUuZkO4h
CrlDgWJ+JXVzV0HL5uq1b+OWBhAs8evdVx9ZH9LwGo9Qy93iuW+Oe02kD0ThRM3sjSAk/T/sbtCb
v6c11KI19FEynPgncetlbgdWpxNGcFYqv1TXVBeFE2h4zvk6792w0rMdqur6tNpjOU4fWOp1gXaH
VBc3tLrBuM/o2Fy4ca3DD1eKhNdg67CNY8Z1O735dQCqdgCEYLFoi0rABookTIR5Bs7ole7Oqi4T
kjJDoQBQyPKIXrJ7ot+RwtcqHH2bm/e2oEN/k6fpNTKqpfxI4wIfqRkENoj52gUy8gluuXkhO9Gj
R5vskKPgPtDKmnlsLFatxuT1m9TS+AMkE1RCxsCjV1V6eawRxJR7oYvXJ7Pj7ld1tPhuVbBIgF2d
HCq8X/B/ifEe5IR85HOgHZetMJPzIsrFpYhZqOBN5jrFczeOIxiEKmEMkA8sBDddkrGoIvfWqQyY
GnH3IapgwJ/dpGkzl3cv18hqVxVXx/POlBK97oJY2AMzpaBBRs3Gt1Z36fJLTPek18fmnk7/jJ0E
YvbAkSiyZTUXJVLoB8qR4uxXEaP34Rdj8GXcYGHJmkEYil01hkM6czPMzbA81Sm1LX1tdozeZqyP
qtk9rgcQ/mAL/yzDN8dtlb6xR+4X28AVcX97gzBN3Xn05xwe8IZx9ir7SQ66n6GxcV/P9e+S54jK
K/FqJptLmzEKIN0GkQcV95mpHz82rEHo5lpzzMUOTkTzzCO+7Q1/LB8qSRFulI6tC9LFpX3CrHDp
Iy3P2ysnbdsyo7dpCiB6kmvZZLlNEeCdob1guwM4bsIFZha9jUNbvS6Joxo0KGCcFKv354jvMZY1
ioNAh6H7AnpH6zbUaxq5v8XpqGgIAYFmNEt0AUkrTKgNwXiHyhWY9XmhoxiFld5y3kzhvCzxg4hi
/4L8AthqGnI0xjab+WrEPn2teNg04q0myTDapsTHtVopBKQPHOCzkk8cZ6RQYCP/45vY0yScsFze
dhHxCaqR+SK/ZcG3IT6Pq/5yKEs1Gtmhe5OL6UGncoIGPNN1p9gTIUxoKo6ZbHjj3alf9reL32Nc
jUVPXyODsFhLV9OIwtKPHUsvg05UX+hfdyqVfoMLiuQL56RXkGyxdctayTnU5yy8nB2V+5vjDL/O
wuDCnR67WzFOzE5Wz+qypnqVvuz0dbQKIlU+WBqFD3NGtlAoFumkUmUOrmaWOXHR/D0F08tp1W3h
lI2dnZMqbeqleT9y1WiW9oM70CDACG1VB7LehmXIWVy9aRSVjZcwLj+wR5DIS6Axi0dTYkeWvums
mXlwJyndUykcK0NuuF+X0f+hmMST2Nqrgf7m+BZqbMvt5LUK1fl69P1zjvKINGVnK3VYJSPwhD8n
olvdzxfOObw2XXtP5ACWmlI9gopXyd2hYh4BVZxdL41LdGRvskqDoJG/wfdQ8DxmrSizjifmUaXz
QzlmEVa1tOkevRL8eUxFTdjz5cnmkZ3ClS0VWxLD7q1/Nm//zFSN8sbLcpPkLzO0QtxOSypDhhOX
GnsySWw6Xp8HBAf7YxsQYGRE+qp8SijWi/Iuu0GPvM6GTeDuaoBVug3JbEeSeDHCNMB6Qgkh8Uoq
iFwkCvQJKnqp4R5NxEQqutQsGWjMz5qKqbRmEz3r3OCLdefu+vEHrv10f7yn4CNlyI7praZu6R0j
mblYEPyYl6ViyFfT+3PGL97B6v9U1GrTd+GwJoNQhsXHJ5wTPyQ0icawTBA+DYhHglulYd11fnfc
DCxJ7njtNSrcDv1phE7WFKUeTI2pySZykaZErixu7pAqqjZ8mYBsH8ZHOentvpbO73nxAaxeo9QF
S7uejoK2mf+Sd90Coshxaa6uS99cHx4/Wspye/YrWyl8V4Fe1grdjHzkGhpj1ZdhYHRLTddQdg+H
hVcXWbtJTdZmorzU3kF+Bc5IbfZKb3tuzfbQzwipi/QlqcRwLKzw4LjMJamMXrRSMXYBLXhpzOEJ
8WijF8522WnRAIgxjt41aJAHPduhhdQY38mL3RwUEvHrbOpqEcc9PMd0I0NIa8b/Nxx7h7UM2tVJ
ey6yfgFt+5foILxZ2Lvs5Uv5tRTMV89UjIk+U3PmQCS531k8QzsfiYzl/paei8+63DuM3QN7CLKl
EL9QjllZDi+G0zOgSxiJFO98iI5TN5Ml1cuan66hZxRqAaAWib3Fo6gjGp+b+Lurl9fSCbWHkdUU
QQdudMNpSAfD0lvdCJu82b7jJOFXLg+FzsiBWcz82ltxiGAl+hg5mvkFVnsyTq+STqugv++U5DGp
ol8KfcyH5zi1XWBRfPoUENTuoumqhdP7QewxZl1lL/KE+8tfWSm9Ivv5rqJBr5T8TC9UdOgMHVTT
VwR0lhOuccEAAlT7op80ciGvfxSOn4ZRmmagXGGuuTgED1jh/b7lxT0G2TSfmBp/eUKbawn7BT0p
HCV5PZ6mISwTS5Q5XYhOC0+6uRdZoKLbWkwtnVlQ8tJ03EAfoU2tTff8Yv9EKDQlwYsKpD+niHf7
qXF6cAko2MZ6g54R8EkRexDbUyiATCuFMl1SU2z8m3ORRdlueo1NzMqdTU2MpTW285rNWKLM2arE
BjM78av6hcRK1X0Lo1wRzTmqalVhcfDHwXtJ1DO/DQTsYrKNNYhRSdd939QJ7nt/GJo2aIdTcdzh
mYyYu+12AdJmAnJNM5AkUY7yAQmvjsGF5HFAg81Ksh+tnoivLlbSe9GqV0l58bK1j7lBfqTptpB7
Ua8LwnK1WeZZeoGXRiErT6GrB9bJsmJDzrmzHaO/sHyzITF6Q7LJrJjjh7BBo8YgNmZXo1g6LKn/
mEGKGpKylM2Tqe4GjhyZuZj6nPta9aIa9rLsaYznc8RTw0BJmQoPAaY5HP2KrnVJ8RpfPzcgWKiQ
84BfBqMvQcCuNp/WcITHU8RXLX+OHkBa/GtiMijkD+Nmpra2aTd53MwDVuZKMfTK+Aymqd9P+kVR
QnxILaJkmUKjl/SYk0TyuWZoJ7D0f5FYXCmSjEznIw4wlaQVH69VQbw2PHpeXPVVZkVrkq74TZPx
pMtn4z1VjZlnbV5W9wksdZxsB6qi8xl0tU1pLUOacrgKUlIVZr9/W+ktVmzfCQdDlchQhxrly9wK
oj1oMnuwuICqALRW2JwGHgCpf+UnNNS2O8zRw+NMa+T0CqRPUV4nkymwb7SllxbyYV0Enu3kHHfH
dAseCy61GtuIzdwxx5iJ9gyLijun35v23kJ3mQ5slTYmBGcSF3XZf7dzKDEBIgd0t6j4vNAN601E
k0mfTPaqrIxDGSSqyvsDLn2Yybnfl1e5m+PU1VcqH5YjKHwwSUpo46KM0Po2WO21ZMeTucIAQB06
fCsD+ZIHUqH5sCEPKBT9ALbbAlUjLxgPXJ/kdE92Hn4Pyny8ijfnifeCMjW/0QZc6x5DZiKdcf8+
uhkMC2VoMBM73XZz+jLvgUK2t9gb9tzY2bjyIk/vuaPqWkEr2zwY0X9Ckva9yKXKGpgeyi5ZZsLy
7WoXXnRSLG95FJ/oenmEM6xuzQa3+Zt3p4NeqiVD1Bu7eZlQ9ZQZk5DAQ5xkov+sl075Feh6uLAF
IwkIcTLdNTWrVklkUktZY0Azu/rNpzwk71kI0DQyanRuuUS4UnCOipmwBwBBZQexQJsiXB5u1FOe
kIiC/B3BslCvn/RamPoYBdEXYBng8w82jYUAq8+2gfaVkjqmzofXOVksPEyX5blbtxZWICU84a/F
rJhC8jHDB+u4HYyPA16dERqc23HPZXaXLKJ1DeEYMiE4/HFQAD2RrbBlBnx+F+TUGj3aSlqJbfRq
52fs1bFDq/9IZG5LNivJ66bvmKYCVTytJTfgHe9mrE9nTblHPfYODZArTqKSl56XBaODMDGTC5Ia
A41mONHf4FHK4bttI0QuzBjN5KORrye57VLO1PexgIwlhaZyhFg75BLrnEL6kqHzMwtm4uw8GN1N
iUk27tmdxZ4etfjWcO2GOUej3/2wsQ0dYBzxsos71iUHqcOvKg5z5GMLMj2rVG2waonHFI7RdHQe
pKyqFSpcLT+SqoDu2RiDVKMzJWGslTYKUo272jeLltdiXgTn38DBF5o6WwdXpW8Ttrqnzk/zKkN8
6C60HO7L73dmpDKbxNlYuvddUGORf+VIUhKHhsPqt+i3AgaG3kcOgSe3WRqLrbaN5iyPC0gcxG6S
EQjGc98RxLw/dD96egsd/9RSCmw6nSAFeA1SGnadvwka51LbrxIEjsy2jOWh71NE2mxGy+NxlwoU
F0ke2thp8Cb7t4GEmmQj/1G35HzePe1fIFRi8wpDzw3nXPsrMzVXYtqitHD8AuOGr/iCsxrR5Th7
MfTrLPl2tKIj9EIxPeKtfYJ0kDe+KI3TrIupcgnyCVYbAQE14dVzlnfT5sBKm7Qbs14ypo1fVT6a
QFa6dBMYzS1c0NDl0r7u0HXsMtC7Nu7Vrdp8EwtCFXW326yOCveexcMWtLcDAJrwU+7YJvR1KA02
kmCJAp4sb0Ra0hhn5bQACDy/9meS/LnhrCVyrKsTASobrR+/1tjqYwlVIGT2in5mLCtuFtkC03Kw
DaYMAryRDGPk9TC8HwyJK/wixsXl4uVMDtVOIMwf5L0Kum5Nb7ZrETdvjULBdhzwRtOsU+npQpnY
fp0zfe+mdov05BL1BJBm6f5ujfU0gE7U5qMY61FU3geHXhom1FwM4cHvSobpJSEwrtzD3BWrJAzA
y2rMNjcNkDanPBreKMG00mlGqDnxKIocdLbHFO9hFC283EinmEmxmhS3DmdJJ5V3Y2pD9cATROZ0
xvcLQzFUoOyoyzh8Q10uJ7uc6/sMDxs2Id/wo/hho2xFKfYyBGowr71CSidWdfa4cchqy6AD5gKZ
2zw6YvPQnTocCO5SU4zgPtR1Mk6SypW89rg15KzfqHZzv61gYxMbls/L2WAnVm6J4Ar9DpoNww3r
8oaIjJuRWUTT/C3z+11kXEAmtrLHqap+3qlS5N9PVm6kiy3+A9n/YuoJwMPzGSQ5UIRuWlILv1tU
gU6t+RTmWPNVhbQbb1csg9MPLEIrNUMKxelkm6s1m9dBoX0bY9gmZVdPACIUbCsM4t+9h+FDOb+s
ppA9O0PaM0Edw3rzG7gI7sB2IMi4s4uNSx0xUi92OXbJIQVy+LZVV8PrDKpi4snN87JJlNr6LZ7T
lnAXVOd7vRMkpd52wz8pZ9QV7cRrX5/JLkXhttEydOqN84waIcotVAqD0GK6cCUx1xh5grmUkOC8
Uf/bpO+mWCPBluLsna9pC8i9/iOQT1xZ8N1sHG2iBdVPQL/lfnoyzfaQZCer+CJGvNGXQNBezFA6
uJB94gxS6BAp3VBHDwHLNMCUohGwkQoYhCUKUda+UeVdf2MepF4qk1yshNEkxlJbQ2IYuwnieE0Q
iiaLA9PGSfAHBi2SUlsWv/8n3ILxT8nWM7StuDvgKynPtytnZI/ZE2GrmFDF8Q/FYqbUrKLQoiF0
0Ez39bc1fbJM+lLSHcNUkFSYUTavnlbFsp80V4mYcQc7M+0JIoxiz6hk+jTcuLTrIJXd8oLwU0ZF
Npw448G5cHMmVWY8TFGdyGCiyXkjOGOqRjGGqGac+t4l5l/CCFbtqIkwTRr7eHAkMOep5vkYd7xH
Fqm5aAUyh/qQQjevk5qhKqSbPYU9Ts/ktbzx9gSNPpchXCROGS5coUU+vO/7khYmspKWmUJWbfM6
SYeZRB5gEeJHLOkow5C/HUK8IOb+JaT+zop6HAxH8ISMbcF9GYnoqMLtj2CfaNSCGOQ2K7YrNAZL
sGpVxwio2IDROri8bhdK1PygBnTp77aQtNcjylLqP7UETWFubp9Zp5OYzihbMzsU3kwqGJltK9Pa
KRZ9xWNlc1abEpTTim2m1yNEmDGs05Vo7DiI40nGl21Y2o/HzS3vHzIJpEqfYgk1q72G/0Uvsvez
20Dwqs0+/3WoqPeLBh436RTNo8X47jiQsRwoA4vmandK76UixtMcVA4Qoi+y5puDd8NRt2aueDAQ
k3KP5c7rZrFeM/ywTFCF4OlbaCYmsctU2NK+Go7JU8BtG/3FUmrP82b61ABbFmwzskPI3XjM0jR/
wpQ3HlNKe9cT/kVhdkV1QqygD3czOyRLcy7aMOBw32o965XLvj9j90Q8miLSUTO551U5KTI3aPdD
ZYpj4rbVMkUO4su6VwaNiIW2wfyboeOexq96hdAo54m/VAgCDpb5VoD8sNmWA6YGzMGsqe39gGyW
gbl4mtTsI8oqAuIMWq76bapHvYhNxohrjaKoEEbvbIF69iXz4E8gdBQV7xcmdpfuoYQX4/+l0UO/
qDsVFQRKxMAlGkEJuVnHartTv8xIx0We0OJdblxbb9Peka7vVoLr2haiqIRwpfhB8LeR4AgQbQ9u
5AYQEdLmqHsbkNkeObJt6n3rMT9lExtsTqupHAzfWctHROIjrU+3ZRWRRUwwzaMZyImVpyOSG6x3
d3WIhYc/8lMJlwyyXpLhXzp2zMpS3k74sELfkzeIGvLkMPrmqJKsYVmR+1qS6v0MmDR7kQYKGCnP
5L0vOaAbinILyB/hRvq2W05uYGasHF2A2bSN5GkQRQH063FqXQQziCtsq4PqPdfLKoUMIWk1kFoX
cgPkiXCRk0fJIxiLwkGRV+g/hPCc3ZfJop2xxAgM4jthkqQAdcZA9q1A4uUH5xkf4o5LN8c76xDm
wdfm0A5bmmb0OxQQAKDaaifAtdmimQTEF23xbaFC8ew97Ckvn/3vKjh6V/JrpqvwXkp1SG/aLpdw
GhhBs1fGMq5xVj6wmNsXNGaSw0vvqJIxIDoJaayT/zO+5qXCt2I/RbzGwyH6YZwomsnsDNgNq9gC
9cxe3Ze0jItkmPAhhcuwlj77+ouc/E342NaokmnOsN3O1iQSay3o6XdkDjbNwiyn8fuhBWFDB9Lp
a2C5Ai1s6jTt66OUXog2EUFF+DIPXYryxku5VzzFUrbe/Hf9IRBvyExiVgG/UgcMtJYitjxB1QQZ
rUlYCt7L4pRDOj4L7k7Ph2285/l+rd4/0KnB9kZbDQICg+1WmyChy9X53f8lnGEHdjQvDk3dshqO
mwxw9hK0nmZqAbNRtjkChqlrvyRvYv4HrtUzh2RWUZf74EfUksX7zfVYscNCjDFfNQshWv9pMn+O
XyvmhnDBPLjycamIC9cij5m4RZZhod+MbXb6HCiQ3wean0jYludZTSdTmW5KPCx4nCkzotkFMUQt
WJpXQQs9Ma0QcJAg97zq48kcWNgz5pGm+UySFBy01OYSa2taRtDfRvwADJlKPaVl3N9Vi3+bfQNb
MYv4X5kVaPMN5ougIy907wIMr1KJvVHqrysYoVdn9XeUgfblWSKSDl/urz1Aoq3xlJQBgcMYffO5
VS4lP5LTshH2L+IwmuENRk5N7r8PkoMR9j0ivqtmW2w/MfICPV09MB1qQhioeJQQdzG27UyRFlHZ
1TeYR9caukoWf+aH2SjM1LnoDgtfAhK1BLEZKTO5Zfg+WEUKiJ7oyeaQduezsofwoNgsZGTDjBc3
FCmQc09G5QAdZCzSr9ryFj/7ArBbxTmpw/SgIQoCedMf6UX3x6ED91ERWF7GHSDw4jAuxEuI1H6U
Q0ghsxjw7B07HzYosqK+pgTcSMv0iC6+v80J6Hyzvf9WOur3QEcnKqO2EsPsqE09071oGGeGwcHb
4AMgbmoQpbj6LQ8fAvpykKpMhfJHV7JdUqxdrNufa3FbgPhhaJ8VkZR5EmYr/DTXvyc9FiUyPt81
TZ7H704vNXwRtnxyEbXew8DD0PQWkQP6UaKorYFj0DNa1Bmf5gWsEDkGdmx1Q/7Z12ubHtTjq8Tf
eeJXKEo1bWK+o5eTdDGTF+NxBazywgFyInSIqrvBS/0ee9mHqDtd0lNAiOM0QDaNa1LL8BNlDrQf
q/C++huKb9NOxyPU4IynCQ8H+SMOpHVruxtRFjwe8GibJ/iADpOVuGCikQWPDfl0jX6L20BxuHSf
4el2UCL42be8/FsI/Mr8dTHhd0jeEmwnufSuZ+vVwXdtOtt7DIEuDMuf/U3ERsYF9Tu1vLlWeCY/
zwVgQNBQbBBVLavY1eZVnhqb+Leno6n0/eEVKr+y6bllucWty0/sGSlDUGNBiCH55E/XmZdC+TBX
5b7LsZIvs5BS2wM1FmKuov6serruj+JcREt9o2pINrfYTGINKolzoTwCJ/HpJY56IUEUARNDjLkL
aG69FBye2oCR59iXN/0seLoOkirM8ozRu5IflIBGiDPxQO9nr1zldeBjIbrG0yN5ju/XIN+AjGJC
nrpJsR0duUkBS4Q98i1FtlTw0j+4GnnENSMYz6aZiEanUrpV2YDwpHE8SAmZTWarjujiNBgTL1a+
G1XLhco4f+WfXs+nkMPmnLpsqoGgfLI9Wf31ZveYuwL2S3VpYvcw0pvbsiGY1Mxp5koKzqRNX+iH
OMNC+YLJsjdJWfLtL8ApyHIu6FcXVV2rA+NvvhF9aMkEOiBfVG57oj8VDLA4UJ5Utrfby/fBIId6
QdVVU5IJ5BQ4a4tNNQxE7cjmtkhQIJjvPJfazL9zXNANISWrpBlgbKN8HTb3ZYJS456RR7h6aYnM
NDUSnmsqZS/RcUB0SY81VeuIh3B1sLmo9AiJdj5f9pBVEIJKkMhptQgtr9f4OBgtiKLDDQOMeOQu
/bBbnCVXUo1qF+qJ9z+lKKtGokjwQEux52O0uHIpsVum628ZlYsG83quzgXAGV1jdAHkYMIvmO72
pEwAs1eN+eTLzk4NExB8gfk9zPnUMolUK8xdXwGChoqKKSRLm6Lk0m9Z+dBwg6nXcL2qWIOTU2Ac
2i0bu0BGKCRxYUKr1WK23tA2hrMc8T1BpfrJLFc2QKb/YI1q1cghrxvtNrQjWMEc7VFF5R/WiBeV
KTN0Pz98cA7DAFrs3w+dHygdcNN/YhvPEBvk7lMbVBD2CwQe2L2RLovtOKLXFZWe1HdA4GaHZS92
y/6R0Ray8Qlw650VBUCrUkjYbDocMe8uy5o/cxYQGQr8ZRgyf/1sBvIlbE4RFvcpgbC31qhH8BR5
S65JN5LPWdVexdR+FwKSJYNznwd0j/bVSLjZQlpGhkqIlDXp/+T+kE/JMfj97csRBauEgGzJldwo
IeMv0QKQpo+eeJ9T271zKuqDqSqEoOp6dT3NedYbR+nHOVLuIZg6KJ3DOEGiDESqPiH6mOsOddnP
6+vX77BVMcxq5XbF1Rv+PTq6CtsElY3AlKnSbksnZ3fgBxYC8ZtfsBiwCRVh1wIQspW/8BtUj+e5
e/luYoMpcCbb6UsSlbWPEKz7gqmNKWNd9jajVHvuun32SxO3/wpt1DALXj6risV0f0mlOUZfkYLY
U7TQauz6pvCvzqEXOjfkXkEhifOdCoRfIlXaqC3VKHPpB9Mz9mv8sKfZM4v5XUkF+OqncTImcbMs
UiRKr46lS+2oB33gq0psrWEvzVZTHkDBbyXycyr+b7yWeU8AEi15to7FmP+h/j2332ZSa6JcY022
3graN6P6i8qNBoaPDqWXWXinPGVjjYYRa3SxAnNtE59bmOs6i5HB3dHYQ0nOPBw25G1OJKNaf/K8
uzN4OoBTbycBF1gU9OtRwQvEGMsxfVb2yI8qDVZD20oR1YxjwbMYwhzNUr8Fo0aanjtIWKxcc5uv
53sny/gNgBWB2t3UWz+V0gEXL/d8SkAJs5Kz4q1FNPuHZApDoOVSNgk8adgkSUFPF+nUI+js0bjx
Hz2D+WQbNBPRZ18GNo3UZS7IAgIN46cbOR9Z7N6TZxAUibd+q7E5c/olC1Z1dh9qsVJfrCbXQMM3
LJHNh551rKiD2r5UrsXKqn1Tw936pLSoki0EgSImOaLyLU/C0NHXiJSUF6Q6JefZ/MLvjAe018J7
NppuHK4Vofrvej0d71eF5syIzD0w7hthw2dlomTYCKTJ2qj+Hz0jXOqE/mLBP+R4xHiFfPcfytq0
8lpTtC37O2D4kddArmIZP2v6zfXoWVdH5sPgbOtS+Buj0eWgvkAPts529EhyxsoyNgRzV3mu0YNT
vR4bo4yJDET47PAQzxpjN9DYvoOGFU65uitnx/SOGVRM2Tm4TCmoY2WR6riorOoyhHCbjuk+z9xO
dEONiojXSNWXxwBxWkENEf6vRCrjgy7opbO5V1lmvylIE3BvtMBHRn/P/3t63kXQrL6RzAcrU4rR
EblqDtE25r4Nj63HWvPxluMLh9uZsSu/M2akJkewoWybopCWnhJSRzZfMZrX17RIGtB7FRD3fGgI
gvY7tCvtpBabRWD7hI0bcFAAajHCb5oxorlNlUa+goFSYaatmrzcKsv1SM5uhJkrcJsnACIvO8us
RVUyd32t9AD58alTeGRrzTC32oQL8fGW5NKUcCFBFgjjOjpqDr/5OcjOIIY/NgTkHUylrDaCkcFK
TKAASAtBt5IJAAwp9AOmU2WLMa8ZRnGXk3JLyWCvyUEX0JUGRdy3diKhqcwIOLOCSH/jzxInkq7u
uWXkhYSNhSa37BUnZvU0kIKpg7berqKT9X9306PYNBNgkczf4PQVjwjglZ30s/xsqaTehaDnmedS
Wg2w4p3zm83kAA8uZCWgynXsMeTQMcOBYxW9apaok1OKUtindBjAXDxc1u+MZmrcF7ZWe8FJmQO9
k3UnschNcdxeth9DuDljowSVfmnHEodyryo6/LDeqX9jef1UoPFbuPY/Em7rZYSc8FkoGC/daOPA
JHHjACXaxnYeCtOLxcxUwcidqJR6pQFSFspxExNxhnTvN061d4MVAWKw6PFN3rJQhypwwV3jTzN7
mmZNPOQrRrf7zIz94iKE10H2rZex9fE8CCkh1EFcy83OzoBR0EGMUeeZa1oYUoMbFf/DQmlkWeIA
puYasuiVnjscP38l5iYGIzttrGOiWTo6F596/JCKRaxjlqTm0eegpCs3TlnrI5N6vbZ/WsjyJR07
gprwgAmxpsFgsscACk+xYz4CbPXTQk5DDmHOSlviGnHZS32EFCfLHsORxYSJAx4FXEX4sbblsHb9
ogqZqzxsgTGW0q5hlQZqANuJgvftGvh2loGdgF6cBD5+R4SGsezcPc6rEaUu2LIqIdT8n0+TpbwE
MofHpXNKP/99GjfRBpOXOWS2s7bHS/uxSUnf3U7VkELdWimcW4C1BR0FKaqqxwO507cfNPtEPPTZ
wP1LNZA1YzoUm3mjrNBnh+X0C7Vg2aEO+y1yxsr/UM3ensL19XpIW1NvfFsvYICkowxnrb/uM6Gr
vUmT7/6cEe3B1K0An+J54jDHHOErI0l45+7hbp5m/xY6DbcoDMFFgl5u7xZIrigpdikj5cfhRe9L
ngvfKcWMSpFMqea6RlQIlQvLElQBDTCjMO64HWwMAtCsGx6efjQVlQiA0Tt3Sok1gP/TZ/LN8lHt
+gh5FeeBuY+5V8HDDt/Xwz8W5Kilpv0c5MEEIZWgEDWeMVBFQi+J6RbcHF+MapVctz0B2UDZcffA
HSVCEu1+CEdXlmMvGiMwQgJuRYf9v9mB1tcPnFXCqX7RsKQfsC0QK0zEJb0VzSp4xZfPpb0FGcRF
oR9jxIjYmJ6w5NTHZYhJGqT10WaPwWcUolndAnIjhM+3A9Xz34lWexh6xLvlQWzOfydhFHNdLJsT
9w2iz77CXbwCC1lmEHXC9dydDnzO41KotnTmqakn+PKjf1UWsCkhdgoai2F7IeHG79aec0dC1BnP
hZe0sg785WzKcZsbk3ZXsNPrLAlTE8cdkxnnPHjcMxvjB5lUgvo3g52+Y16dNO1AhmHVz7F2SVdb
xlrqOJ9qamZB6qBO4vILsQwODIhLvuWW6N8QyTD6zlfRkc4Qt89k6dobWwpaxaz4FznJ+m+so6Ma
wYiO2khZzsUWrO6oWhNYl9ehHxRo6CeBvqy2DihIQbj/vxC6KiipqkVmXLc8ZVbxgKs9UG2MLAwr
9y9AOnxKacFOQrhaOIDJGK7IK1YBQKOy7XsmD5uqXbUlSZ1hJWdYv5ouefDnXJzoaqIoV3C72m45
LGq3/hu9Qt+/5Ja2fJvvN7hc2r2CRlF33qRWdxrDQn5kM2HBWqLY3UO73A32OtGwciocRp4sLWkL
9lt+grSwYpUsUKSSB/o3hsevJx6v/YMArlJW6N5D20qhiLoaPx6ahxThlUA9936A/z/uWdyfwuB1
ojx/Zimfg2x3DGjTzBlBiK5Kg1jX61UAPderxpyOjkn/qUaljH36UiRXGRK/Zv35P9Z7W2w9AblG
tkiVWkDzk3Xyq11LZSNOprAq48nsUMGJEmVofzL4bQJew5MmaZ3FKZFVQ5eEU2pqEVwDRUEoTtsM
+rLBYsypU4ru0lUFxWPXtZLnZ7S6SQSTsLZcFWci6yZ4hULvbH71b7k/+O21w/FLHFaph6o2JgLA
joBYzdzuNL6RCrtEpmLMwZl2LH4HLIDHrGTMLed3dZcv4ywCTSD7ch27u3LwhaNIpuAjaekKhbmG
woCKUpng0hJbXgbPyeQ88F4k7D9Vp+GO4I+gf7tAc3OVLP/fN3FrdPS6zbk6higeMYoOmGz59K8i
ajI4i7EvYzD3S5k1tU3LIrb+HnoGsazWYXjZu7nXso1tnDF3TE2kvkfBlgBtmwvfgqeU0Basm3My
BXwkPY7MgvMtaEnI36itMlQi6fzWjIt2dXi0WrTD4Oi8xrvy6tcq0TdzZM7YbEfzTamFHnoj5uPI
ptddlxf2Pbu3A5wdfYx409+abmqXJ6EoY6cVF9Gv1jK0tvPE80Zzq5LwgeghMatf1NGlzX67PDK2
izWvfoDl44zMv4Ga/FKDdsntGCYp8dlgryI1PwuMvGt9vM+h4f2Td+fcxg4ntPsykvIWlm8a8bO1
2QcsEKjNLvrkII+ltwJy8IPswOA1u+HcRFnvNelfNNBnzmNS6HkKIaVaAoLG5HwgarWma1TQ+iyZ
qUNIiPRUl1Q3RTj6bzqPfpBVmBdC67IGFseJJ1jBg8whth4t5KhSJ9Q2pdoCEp+wY3bz5Ic+l5Qa
WCVWzK/TA/xfd8xwA5nCxWs7QOOAaNDSe38OOQmg9kUhQu15cAwhx5U8u93A4AopAbHPauStJ2/2
rnwhnno5nuvuyR0Txnz8scntY9NITLQWn7d7LKjRm6C5Np/lhVbrKVAQip6cVkDuoON5u01NKmRm
XgQlQsiKsFkY72yw+KxYdVlZbgjvzPkGKLyQp7/m/RveToJvY4ktdd+sXcIns8HUgMUxuXcntS1W
VflfXxDHdKsTmlR91AoErjmci7/PRZpHzWbTj2zC3G4NJwDUPK3GiLiMw8RDirFIAEIGplTIFn2Q
v3+W3ACY00on8zgOtOsn8p+3FXTshx7NhRvXG4KmsgLUx8qy/unobmFpu3r/zukW5SnbipD+NDsc
xDVxbpi/4Bhm+utF1jXIPyWPT+5+ktxowSyHSDQVaqQyW0EaHlibavJ5l+9kjUAozaZsipl+6B1X
Sv10h8gTYDoMhb2azFma6QY3OJzxOoF3fz+AohiZo31U0vdTH3pid8Mviowopz6ewJbxscigwmQb
dj/Oy92kw1PaZIGI1LXV7XoWXHKEIpt4mhRcre2kLTr1pRvBU32b7Ze+LICF8qUkcwxqG1gy/wM+
+7uMF43FTG42U67QIDTqqhnAwt/GUe0SKi5SwOewOq0GF1Rix4aM+9bwPXSu6NVgGCqcCahym9sQ
PDpzFoxUcsxifTAX4v4gXjOJ+IeZS5fEtGY/pfWR80XHSZsL6cew+UXu67l6uSTmKjB1toJzgWdn
NiSyxTwWJsamR/ksajETQWy5cMWRM/F7nSIZD1bv1XD0j+pcQe+aqcxThQmyFr2Skiy3pgft0w0G
4lyJfOdIN2AirWQ1e8gnRKE+Q0Ad/vuezu3rNN+AS+3ZyFPdPv+69JuUENa0J4kNY4L2OX78bvf0
jOjYLcReE+/XqByGDsI3ezcZrSkc0uiUO2At+1gvh6Gxw/FmIVRLenvHoHNUIRIBsXCYBcXig389
ts2dk9xVHOzfWxe87k3qUi1DiqHzaYFIPn6vDR8PVPJ/pye3ssWsyuMDeDwNz5T2oncex4r0PAeu
kVXUREec/Dku6O6/dsM/3fAI5RWdr0Wctsd9sjGdA2LlFLdHcd5WCBgrldtzRw7GneZnDGqakgzX
Kuv5bXkOjHSM8PQCdR9yNlt5Sehxs9bnwuH/JmUJgx7p9Rt0VKlLmwJ2Nyr5YYuGEUYw43JM2re9
zJm9nl/Sh1GFnAMJnn6azm/ZgpAn0SLzYt+KdcHrk4umt4X3u1Elbb3XdsAFsQtYjBchTZHTMh+9
1LfpnnsD0SyPYi1Let226Ag5nMsKxS50atQcywzQL4xvvFL060ua+yQoiolP0QjmDjxCDMI2y9k9
Q4vHpJc5EA+sJQ9Gnfb+RLMw2MERr7BBttHQ14EK0JSCKf1Du86EaYuI0cBmRt5lFI2zC3aa9l8c
cdK+bEosvHBhT1OC85yRd08cSCCg51VaaJIZif5Jd8s0JgZAQzW2v2H0SZ5J4+fM4irGKxX5rbMp
JG5S8Qg1Xi/c1htcWMwkhDcBLP08QCguMZBOR+TkuvzdtXIJQgITZh8hNPKui6G8DrqVhfTRRPrm
nVorhdtWAH435HLcEK+if7haOJayKkwWT06zZAnxECZmRxdzAB+5NcXgCKSHZWf6TE0W8eES2exp
qVKZVUTebDxdU2W88GlHRU8Ebkgmk7gbAr2Bcsn/gKu62Hp6wO5xLA1Hk3PHtI5y39GnHojsslSL
Tky3SepOdSCtasH+46Q/wwUQdXoGTYl9thh5c+FRlVnm7w8VjiVT+9+oz3WusRvKPbEkTL6p2ooY
26YWjXNrSwY4FVqF1/cHmO3zjoWSNAlfbNXPVzpN6LfflHbHapzRNDALUXVRT8LD4/ATXzp3C1Wa
vpibpXSChEaTUgJwxWvoUuIwctkwsZjgfAmzM13rlk0zPHewXDjcOssvTcHPNkpLizb0Cx6FG8an
dFHTcmfIL+D6iI6J7ci+FGfo3BNkgzhZ3xcincIqwBRdcm8dd4Rvfw2VVNa2edMmppvN6+MNGoCK
EzQmasSY51hlzsRY/sQfi3KGByn7qddA1ARf+yKAsgW0+J6sEmT9IjNhq1QhaeF0UmBQLnS5Q26z
pgVSDetRtAPBPCK1qkrZ/vhcccnsAzvLG3M59qL/NE86JAKPf69Gg7p6bbydhXYDHP/mdQfUWBlq
ylZO+hNn2qLiTvOXZbJ3Hwzz3e0aWdR+B4LuYOYAuJc3bXqxkWMRERb9FUiJ2a3uUN6TSFFNMMlX
V8Sumvh7dNhCTb1Bo5B/gkW4H/7U72R3RlfJ13cVKHJFasEEvLe7Jg9+13CgxzBpDtfw0dmajUNe
M/dozj0yHCemvHfDVQ0AgCLLfPGg7AjI7E769TENS5LHl+q0GudiMMAyhKAHOkqj1SVbI4+gBz5v
DeKA4n54H474b+uuFlyRD+hhil4vIYpmGE/lmWpLY6MyhWQsJP5xJaVnw3BveyZHlyxvdDGo/1fU
4Po1Hx0hr9Oxn4Z7u8Oe20mzrfFUiDogQIeUNQxt6ZWZw5IAV8KuhoDgAFGDeoQuD7SQ2/Ax3MJU
qNK1yVx2Hn0jdydTf1pYGhnTggG8RWEhLZvJytaZvPF3xkM9WJWnPZg7uzaf0WqndtSTey+0Hene
XMUNKxDsDcsR0UgYY+kuveLQo/KeVBEHER5YDDTLhSNii2WzOBLGvkM4ij3REYWB8B3VwEkG/Eib
atXbygHBCtMxCUSP3kRaCs2gw6Y3h3Aj9ibknjviQzVFgFQgTRE51XJk7CAAfORi1yt8hz9DgN9d
ZW6zlb7YSkV6OMGpEhOnDr9pjK4GyzNHLlWsiWXtLhCHmLIzPEm4XQMNnzsGJUKaPwbs0dvGiOo0
BkeYlNEc/KIYQp9WLiTMEPGa1EDC2NfRjkHmLqbDVFoe9T/A5kbzztHcE5iTAc3TdzaOSSVmzV4s
dmk/ig2oC5MV0/jqd+9P7DRMSzBh6AdXwS8wia7b2+f2KgU5QoSSV/pwxvfRKlZ26HAMHlMfjpZS
WL42uLXLgI5nyoyqpncy1DJE1nWUfEFXK83N+2xPGesfkWPgFjPkU1MhOjWMVWwhj64PXo59PnLT
I879ZcwhMfoWmu30gHrx+DK2Z6QOLlxqL9Zu5mC9irC+jaaNyrQVvKyAzQgxCB1i1rPlCY1wC4iV
GZ5lEVQuY5qdEE0g7bj/iUggyFfJ15WRW1xA+WxWcnB7OoCfmEd1KL4dNXrjO7ODKCsN4Y+ZSbUG
YI1hccuEfbmzwu0xGrliFkLZqOASRR8kWqeOQSpEAjnmo7ba0hz9+iJ3Smnx+8scEEIsajnG5Z2V
GSIw4AOc+SP2Xxqvu1qlyK2omzMg4EW3pLkQFLKhjgvTZD7idG1GbP0nE20rEcy3NnZ/wnMOgKNT
/UrocC0kAs/nvlH+UWaiI4q+dsdtHh87DPyMHtvaUF6vNxTcplqdtooW0E8VBU1GVtX0YzBRc81L
PVBDRfVq1iKwGiWpR0HG+c++6/TZ7TqD2lwtRtRbeMNLwzZOoFQ03r9WdDhiX9mhoEc0zdcq7o0P
6F1hsW2+d1KO9Rc5y1JNXieshPo9KQ3l+57xDsUf+qJBMAvIQ/AkqBD6a3Nb0ICyRlHa53snQYEP
MG9/OEsP2uEfTT++wiePU1tlEi8eev8OGgZpE0YQ7jF6BwK5dYRzjhxhkYKp2AQ+DHQifuFQopmq
G5SxdFYNFKcl39VH61q+iVYDG2V0ny6zP2nnw1fSwzmESSI1OtCwxY1zGoq132+J7TBjy8Jyh+Pj
gsd2H5Pe+vWogQfgNny6aUlXr3c3wO7izY6HBsvz1lCXQh5bHKymHY+vyYfyEZj4kMAHld5ACpga
9ZoBO9jkEILqfhRWjGgBeiQPb9FB3+JK0YjH60xYBhCEh+HNZ7FUinagtzBY+u/8XP/0lK4O1EXK
be+nfyNRzBCurZZlkej+ndmonBE0SCcscQOOeMtjkl8UcqzVcsRkDkZ/w2DnPCBqwtGJMVUWW43w
gngw28gzU+tHY76u0VD8ydmJxgBzVsl5pLfu7BTEx++hOXmfcYB05nLzEsGwffmU2lRJG8WOzxXZ
ZKgnyQxk0WquKn/yUB1F7mRpxJ+VVZaCCU5FJE8pANLsp4xL+2Xk52G51+66UT/3CsKe8dXU3Uxg
O1sXj+Hj4bNOfihSH5nXolWqNfKMotuVy0pEQfrW4pPDWKvo4aiRE78TsrIcb4VLBhotLY5TeDq7
MmTkfpFBQWEp2qowq3wsGs/6MZjwGlbaHJrGRnD9+DL3M0uStl38imuU+kIQ7Z+EIT+n69d3bQ7u
NK5OwBfe8GFnXF9lgHDgXeaZZFBz6rSp4BkwKJN0IBbpLWEVBGpRA6ZdYAitFvk8RxxHM1cRfKYx
Xcon5sMqXO2rqt2+Mlib+d8NrGi+2tMRd4MDMyMqkB43jinjMOOvQ0+hAzS/hlhxvMrGGuMMUwYi
f6GdSoYj589OHyVF3l7L9Xh9GSTOKMDfnXAclR3QB0nR63rCUK+UsHBRo1V3mTcZ+22GrWhZHu9V
BlujYny8Eqh0eVSUFlZa5qxyc7et6cHBp+SZXR1FUvXvlcmfTfF1rp/xowfoKU4Rrry6lWA4cy6z
Q5fdpIc9GSPNMbOODFvy0TKm9ViFtu5xP0pEiqjDgRZBPNP7T+I0D06iv7BTy0p8M+8khoKLJOG2
7yolMkQU8FKMTT7EUyjUmIkraNTLKo/bzOhZwZLuRVFTK2dC998wytypx821Z4VkBzhk0VcG+Kzg
8FEprCgCr95VcVEDiAmW1+YRJzk6iHHcZ17os8XSBXbx6H8jjnUitZAJnSyEjSCj9H2Ax0H7j20I
O50K0J/G+zVuCpZJZUV75ZuIur4tXdOTWHiffBL0I24dINrWYikifZPfdx8CHJS1UX6733JtNRUc
OHU7Q1cz3yJrMEvPs9Uxgwu0aBNwRm2a+KtyNs6dw6E1bPjidepR2agyILgS7Hgv9qfxhha0NuGC
b0KXU2I9L8cEfYXOmAZ6C3wL/73Wgoaw9g6WvjoxTKWZtgI4P9KZn55giuos1a4danMExmQK6o7d
p2Jyy4P6SOBg9/tvSNUxduNLClhM8bJbvN22XdOZX+70tj5Zx7nvbp5glJrI/MQKvz79tQDJLnqo
DDM1RhCFgmIcr2jdus1CjlAhQsUwFOkmWs0M5ebzin84gbVPyiWzsAgx7RiNo0Znafg1EpHP9Oua
CEMqJwLFFMbPM4If0JSpINN5/ozODfNu6sOqB/GpqHXf4gMSKlQ3ru9k+ajD0a8cnC4Lrgh8M5Bz
ucKYG1292j5n7iwFz31+11cOUsmXMYvgJGCFj5afEi3fYBnesjY1M73IepAU3egLZngsr7/GMNrB
IudkbFZ7/nO0ZieWhNfoh6EhPW2/IMxnyEdCaJfijT2D9C8spQ1+dEnzLkKTw8Vb3IMoO2tbDQWM
NdaUf2oNQjVKl9wE/VnH3yOrtNf/V7GcUF9cK0/GXfAj2y8Ns7K3AHppg9hW2fuk9NzjZZP4W7qJ
Lx9bhx9+Lq449FCnMkUVHpAnVgR1aguljWYBB9Ey4wZOKHHlJYoDU+z7VggUK3F/uMTqT0jaAv0U
MpM3T4ji7K2kknx8Uu45nd93qlAZgD9JtTvaJMNk2n0b1QIUz+tJ4W6N1RoWiX8OjDdnRMvf4+/1
gm60WGgsSsfX8JW7LqoBQatl50nA4VBFKPHbRXSdjswjY4vfT5ewhihhjpSh1m0grJeueOWJqt7x
40DKwf1/D+/H6z4MVger8ICE/WGwcSOxsqZgeGOyc9euUzM3XhMSf+U6x74hwVXwsF+6GMHSWEP2
eALcuI3NcDF0xLjTb3vq1cuGVUzxrvR6A/F61dEL0BnInBWnUMUMFZWgxe9tFEowV9gMkNo1R64W
0lALGI6bewwxhXtb3UQIbmA8s2O7TbnLoaKWpw4XZfT868YuZsb6fbsKoCh+R4C7/gHUGJohZdWo
oBe6A6mYmk9by7UdhULcFeQO41nXyQdldTmoBNcO8n3+4UlkiifwDgoHQxIMlodbpTTeU7ooNwYV
F4GuIzGk2EZz1jWUofGyDUqPwJca3DE1SzR6MFLMNGMI+pgwtyD/w6uoIr16w0M/LluFfEPkBIUe
hlKXwnib+P/n2U3ge3s8I7G0h0F9l3mpNb4hxNCmVjdIX8BZeqb12haqGA9UZI7XRho04JCPkqkY
pMgtPLvtHoC0EuOEu9gqlB7YLI9V12Jwdd7Y7/aUBtBbcm3JiqzYF4uzbdLCC03Szk0ZfYVJSgvs
id0pnoKiSNirx33sLjEKX9FOfCV78NlvJG7eZRiO/D+415jl8xf5aPfiRKbBPtzrDev7zqIWChSg
OVcXJ1HwDQVH+zW6lEOJYMfYA/CHu9MFll8DADsE7YWMHvhJY0IWvcPG8GFpA5+qeRvOPz0Gp7sa
sKa1bqLIM44jIrHIKVwgeNe+xvoBJNNSd5TIUlqKvLiIalCFmhi7SClCmyHn/rPZkBDmNgkdCgGk
qqCm1gKBKRo2ebwe5hySmQvrq3Tg8tLFOdlSqrZ9/uiNKFWjTdtlHerF4MxgNMmdm7gqsHvT5ZqE
U/aZzJSil2dBAnRiHa2Y/NWo20sKAu+gNiYun8biCTLYq5czLEbispgmn1xBd4wwmAico7P2Huxh
dJcMIwAtUYQvNLt81dXvehVhJxCukk5Cz5LTKCF3+peH/H6pUtAue65P23q0RNprTCAu04MzxvNy
hKV7MHIBzsffDOZ+Pedd21+xCK1b2mfRYXgKbu0IZiJ6WSvV90KmHkbS1eYyV0PMYyVEYeT+BSp+
D7FhN4NJ3r09wgfV9/rgTQblpdbd6k7FgcgX/bdTdYs9L7wk4iHtY6aoakcXM8owx8tRmVGvcTa+
1My0y4CEtUnAwQ/DZFS/x4u5+RjA1q4A0eGLx/BULRtC1NO9qoyYeqJNg14ncIj8upZ9X03YPdOu
wRevISeDbGGCi/mSoCMH0q9YNeqzyGZm+f2A7eCCqfis2OzH/Qj7oHohzveWZZwpKeo1Dgtlh/iW
KEPWrbmin/ZNFuiXosYWxRPRC7Y67rOoSnvKfOpO8l4QX1Vs/lCO7m+XgJfEVdaKeFz/Z/hAxXRr
3LvKoMkEYO16boEhNjN3Ug0gty2hbsflL4UHy/UT0p6YN1O1kMese6wAOzmuIeiNVUi/DL4YhC/s
S9w2fwqzJJwugl+hlkao+bIa1DCRvBqod8/Z8z+REHIQsQNq+OXoRzvjuU3g0AD41s40HLjsw69e
Z1gwyDES3A6jy/k+2NfrA0ndnESvPoiFZWIjDncMMqp8/RFGKcJRkKFU60PaUJ8uYPA7d8qKdRLu
bZdNWs9h/JGYk/UKWSlSBlf+JU/Qy1Q4NpSA3zZDZjhMwxlxqTZGzsxLBWpl9DOC88mmYS8h7c1Z
17gg/Q+etwiY1qF3mpXZT1vZYGB3VKQRATQw/kHN86wCqk7ZuuJD6XA1Tl8Wre/Sqixoz9Pg6nWg
DddOWUNd0rOhUNaCOoU9OdIZ12y6AhMBDaAJPPeBnpaQqnM98lYh8kHV4TaLOpQGo7qA8+g8a5zk
1D6TzjZUTJfVdkURRMUr2y3XCrDBeE8QUG/m0mId0azMcuOjLnlH8CBh9+qRCYOmFkoDcmRFNCB/
i8f33zxOT7R2y0Ac0Zf8BGqpWegYXfQBIIr5hV7XfSmRm1yDNcnvZz2G5gfimSzjAER+IFiHYflP
IutDh0sLpACdYJWUJ9B+7YybPqyyFiWVxdglojQJlu51vJRDhHCyr1hzgL6ttvLyBFUDnARegnsd
NzzO2amZJGxmXmFYz8yUNkD+e3J8AB6PtzErHOCpydp6c9PZVnErzUzQmN21ljha8TQ/+5EqQRUN
t87HULz1gNFBRxkXZJW/LCnO2ndop9CcF/NneG0jsW6NB1VxJuRdwNeY3zO9qR0UFY9fXIqfbkla
vXEbyplsJQk0RR0myy+fpEVc/uDxKUviapX2kWIkP3KNbudP5shbZwdwbIETx6M5C4aYZTH1t5MB
vbEIdhKcqSneL2PuG+BF4xN+rNxa2r70ZJYJw7N43Rs8sPciTWgYQdSxm4GGVfYAaXRaScMJNDq1
RE5MG+JAFhqr171bY2fwrfTWi5JPoysSVnbljbeMZ35xM4u5jj54yv+GB7awJPZaOAcdPTNtR80/
u0zOHAk7zpAE/vtpkAANGyV3M3Qm0oXWnAhDiVTe+/iSZ2+Sg4U39crfjMiGNOdH2n7rcVqN7/LW
3SDhWLlcmSIzb5D569TNaLmPpV4xXuQuRdxydsZLt5iceRk4guu6vKYwBJK9L1qRKdWRjKbq7Z/5
kZeBPVFVcIO0BRIcP5DEnW6gtI8TzS9a+loTDkm5HIEW3CZL0wLQeioDl2JnOLHlnE6gGz3aUTmt
nsUAb9bEAY/JBFIj/lvpGAMz5tXYeoLP5PpaTwaAMca0wqOctUunardpERRaud65q0kmKJYbdVA2
sy1Lkgh6JxQ/6jYMfx0pcpC2lGi6x8j5OMy9f+fOtSquH+E9Bf//sHDEuJUNHqfZ+6pq25BCrUaE
CaNT3FKvZ2Q8+28EX/+LNwM5FDvbg/cNtP9WRSHU3Jqx/NQdGa0u7mzzqSaitGciNBsVwDEbbrEw
QSIWLnmJLm8TejpCIrlTXqpv14V04GY1ZJRIG9hpqxVYphxnhMHxXD1r0rx6jaT+oLEHZ3HCpJqH
rLzG25AeMjPBRMcKfxZl5lk4t4duRUw5JoETjRDKQsb86yV90SvYFz5AXF7a2Tkr+2uHzyqCuzrS
joyHSqRblbfHZSb0sirG/dHOwCjX9feFnSUWiIkQKPPzttr0OOGAb7mHCO29dnRxen8oIVr80bep
ZNNQK+7ceS4dqpCJm0ZtWTPsf7ZlvSzXxlZV3Rw7JjAZ62Ei2nSXhQyI5wGF/K8AFKhMOFq6lUOP
gudxUXDvPQP6q8d6DfJhnKWp2YsNY4V8nq/PGGv2Ma+OBmDNK+IWqh9MaizEd35djH2aHQGhWGnz
fcwAjymKkcZ+5WcvUZIx4KPsiBzGEPPJ3yFuWeJRYk9Lutl0Vy8zgh0LWVnA3Oi2KW0c1GLcA3Yy
G+dfGprgvGLC0SoXd9n/DdasHTlxSC7KP69gIRVgyHmWbeySMnU6z8SomHe66cKAk0WxfqJFSwZu
mzAaq8g1E7X1DqLSoepgLMYM2DaBua78yrG6FlOg4qzjeMp5Okmr8w5rYBH4mpvB68sKOgW/wQaC
8fOXssTv+DnWn56juA/Vg6VkSuPx1fNtuGTUP5jB4OB9PdZfVnikMYZKzlndh+sSq9zDZRy+TYf0
CP7XfJb/gQz0Mf80EVnDm+mjtdBDpaKBQE9v9U3agpTgWiAgfaqCc3sLIIZum/LpDgP2Vr816PJt
/5HjkX3U+D/Ltql044h/Esq/sIvbgcAJiRRxe1OtuA8C7RtEmhahkanYemUVmsl/S/1TDPV1mW7c
OaR4DFVPdrwrGcYmz3a+7t88SlljGOrVtZxHdomoTHFt3FstpFrmFOUC6/D0z0MHsO4mDPSClZsT
nbU6mhsuWEvK0pZ3G6IZ8U6VHYzjx5V8spn7/rMtOrCuZ89W4T+Xdufagi+b8h+QgMO89DER+nB4
tZlQAFM8fcMN+bRvwq9aZO8PxRp+CiqbYBVAp0xOeNS0z0zpcNmwCkwFQE+ze7yEAtzoIiv8Ak/o
0e+7G7jlxSuxKPtE+7hxBCznpjsXVhqWbyuljnAmAp67woAylNVUo8WTIifMlDGjtGT8rIZFaLZv
GYzbyVqNXIgmmMIe/l+QRVtmuxnMo5OINWCTAmVDDrGIeE+H964W5zDMtJs+p7OtAWU7q5qM+Qfa
bdkx6oakKjRm/bSzCO2vEADTV+DgFG5P+93XFPxG5z1Q/6iOBUonsxVJ1cgbCtDNgwQoX/B/SFvP
jVkD7teR5TFL8YTyaj7GaDmsdUH6TBv389PiKPubapf/2MdGmzOcEtwnqN+WLmd28opRL8rlvLlU
1RyfXuyDm2EXWV4vSLZhAfxXbXsuuAlG/Mp2SCzeYmJZkXLQSdcjhnK9seh4eYf9iV0L+Hs3jXwk
j1kBW3RkPlneIsTV/eAfSqfCS/jJTp23T1iR5PsiUdZ893FED8kPfOcob6PiXTiVcctE0k8Rrs7s
UY6bXwrV/J59r6V8VqiVnKd3PuSxXllcGegRDWuTKLpOLky+y07x8qFul+mURhG1+P9zaW2uM3+Q
1fFwaq8RL0cpzEvFDJlAauQwasolAAGKXFmgYBAnWsXBqWqRXedAbzfMYlyMcUR8GCRK1WXWGMWm
mYdvN48uhbbjuVTETfKedtJeUHyBSGPjbs1P54nXs8zdLb9Shb2haeete+s8h+5vagWY+tNmbKe9
w+QL6Ks6mVeAui+LprzLxH0Ry1iYt73jsI/0300Jp5fj2gs5AJGZt2kzokNubj3jbynNjdmarf1g
cMCNi2As81nxFy1JbXuvu9D0B96G5ftOjj0ZC5z6mUR3AqjUwD58XGaT7yYMHmPMsJNYNE/kG0t+
RF+ML1DRO/0gNRTGQizPCKH29nzjODNn227cvYl2zbjkq8VQEqdlJgeCAhmLFoVIg82J/fZWFZom
HxtkvEBFJx/J8BBgLZeGwVktIae9MFsCuxODPreOGEAVgIb1MbAclPIKB0Dmm1JOQ5g+UkZEc0Vl
ut9beNvpPNFdV86YGDdEp3RUnS69lauqM/PMGC5amVucoGgOZPkSKv7Pdi1h3zm6ZWQZGrq1kXn7
s75bTZ1FyK/rtwXTtENCU2adWsCIDVqwWbpBSDTWeIMp9RlL6vZOJLxUuMWWFmzWwHjhN5AFsOqx
Cwoz1wM3gmeJsFAGqxs7+2S0M1E32m1jXGq+9yK6uwdexGMvQxJqGxV4d2poCxv3PERkjZ1JnrS+
jVxqFBeDqCmz9Gj8Swc8CnXEzPCqNbF97QuuTN4H1StlybnUpqsSfCu5x53ZOHqwneE0qRT5H8Nj
4p3H/njPC3JnvCmi2R9QOFG5lstrTAsX43YH1AEJz7R7pVLjuKUG0zsSlhPYdGE4K8J1gK1tzft3
zCE2JQ0Bjd0z1El3wBs8elXGmo5kpGm+NNX9YWDV5DS1vNpC2+D3AYSmcSITvj8AoWhv2E9em9YH
qMbnk2oJZPWujwNFNKN4L36VekhQCBtRz2XeWRKUNZ4j8nXvspmKLzTpL44i5UAKFGEh09QIm+g6
ZsRKCRgjSeZF0wILFXqMjnfzyUVr/x3WYERQSGZaexnV0vVj1CxsI9x+B6lm2M0BoY2LR8hKK9rH
V0Im50thnllPAkr6VeN6Sy1M0dqoDfr4cCl2dgyr3Tap2oMQHlu415DDdGplCWQAAjBj9666zFUE
x2yV8FDulU4OQ/o92tFpSiHgOt/0HTmSfV2fSREqOxPi2V1jwwCGGdIUfpbhJR2UF8c/3Hlzs7Wf
xQLrNj2rrjv9HrvEQd0RwQ3rq9ifFwHoehmpLC609qh8KPTfPHFXI/QcrzMp1GTyUKKNbV9+ucWM
oU1s03V0LLFx3v/NxLhUvO6Chd5cnJVKjv5OVyUEp44ECwMJPvYmuXnOEBmhV3PZ5e78HbejtqEH
aN2ge4FjADe1+5141dLUbn97vNT8F/JzMQa6k6Z2QfHep4W/eX/1kw/QoroSm423OjTjD9Ue6bEw
Wczw0TE7YJmV581RUKwWoYF/AlVTM0QcFsYuRsWj7AcCc48pFmX5wzrho8xn0nJRNpqfqLqilnvh
j9nKbFetc57PiTnSRtV+RQtxQ6MbyxW0LVOXyJN+z7wAxykzLJrQIH15Q/ubo0Ojpzf0yRSkA31X
DckNxxT9EuIIDmXnSoqAkwGMVhYNOU1Ztz67uO3feIEEUS7cN1SELXBOAsunqLkwWqYP4V2gY75u
rx1aC3ybOtgycdHCAENngeYWJmyozKnr8Yk2kKkXtudU5catHKMP9Y7bzaHySDfg+ugBCaXtjp3X
qwlLnrDKXlzUr9rclBAH19P/Pi57yjrlooeNyq/C36BGPBZ4vNE+RUV8dn4tYfYq1x2PMVwiKl5C
FCHb8N3CEgXXpPoToLjaKBdrwxIWeJjgJrcgUAxHfpsWEOlOqrjAbgiG6bCF+j5ZzA9wdmGkbBny
GOjY9cExpEfTRmkWe3zKvvz/eKBOMrO1FGIqYycwWwbKsS1c9oL/R24WCio7y7q5eeD4YoX8u4Qr
A9esy/QxF6NCt+zuojyRsPovMZgEdipNUQMnV1sm8HKYeQTO80urZ8aUBtT8PbMhBqP2emZ/Im2A
B1ww3ciiDuoTta1leb10mAw8Q4tOS6EZ8yT4TXIQuFmUqFQ+6gy4mWW3o/uabHYOzL2GKSwYrzAR
3Wr5bJdKDXGD+adTdxRdUQSzfUJgdhtiGFuqjQs6hwPr1zrVqxS3oVGz/RGQj3x31fcWwyc3ekG8
r91sh9y2MRBG7T/VlQwvh80dH+rMb6uX4yLpszoGHxkonQeS4C3uasgf51La3WSCLf4L+I0snD4P
LdGrMa+TFb1s+6c2Rh5VX9p5hYoOkTJZmTLgadtd7ZWjJUiwOtghzjsJzdkhgUCKIc7K3TZot2ja
R6VbRTmv/egCeWYgXqNfqMVoCbQvtLAew9P/fKcoIfWWc/bZtRDP2h+Sk+bm6P/E+9DwoBBUZT01
3BX3UECh0bs3mB7KzgFtibkoFzwgeghzf8ywnQr5pQ1+7Xrz0mH2X5QMuLaJSysbk5L11ukrH7dd
J4kt/J3nXTVBxyQIBj3Y6tuhS0XamJEJv3+zT/4pAEF2UHvUT4xuS503URtjh0HoXy7OOZafeiuU
GNtD8iSjSXFEBkloSvp1I9L5/3JtNiQ5BWJ5Dc7aB43hU83MsrJI4JRRUR1Kiwkxf4yZJ+C6HBb3
vllbBPUdD+4C0u2ZimbSJs1BtibcFvM38LmsBVoPYWzcgmOD+lZ7JQIw2XD2MPivrYfc8zBHZsW2
kP5RMnCOm1iQFZWJijsTJtQEYcfM2cAfmMy8Kg06AZsQpr27i+sW/YuU84tdpueQyRRW8tSb2R8Y
cndbkK+AjwG2prCiKrMQ+mblqs37lB2IgI1wf61Y8z+9OGPfoqzc3xBSDlusT1+yHO+s2MQPZCow
PaLsK7bNgilc2Iafsei+JEXqToRns8iW7wNTij9OoCpoCGg8fC5tMMilS/aQUOvap/1MMGEyCVQB
k8zj5dlu45f5VS1cm5yhBEwPIgraObVU58Dz/LPLU+wTNd/EJYO4kmc3AiKkuDObl6XTkeBGTeV/
bUIyQW1DDKHZcDTwuZkkrRjOARFTBrGlZFIxyvylpzFw272mBF3qdcGiW6236PdG5WKY4ZYO6YIQ
n9pDzr1SQzWdF9RkHkKa+FxnrjYWb1K+P//1ZKXuGVNxEOF8B8sVL9C1BDddThTI81ZxoVHiV0n+
RViGewg16L4b39ARwRynsN8hSV+GAdISbGT5rZ4Fd3rCi3GYqz6vZn5Od85cnmXrJpjFPN0HOnDZ
uO0ImAfFQX4ymYsR7IMDyytITwaWuQdUbxpnTZ1yXoUO5kF00364xU84XBzv8OpeutK6U/napWZ8
xDcRfPcOgqJlBJXBkiqsGLCmHCMrVljIGrUuRq2nEybHub6TDmIb1xQu3Ygo+VCY6k/43+F0k8D2
L0meJ4TANQuGH3i3JR1gtNecb6t0queTaLwkD92nHI88tIEtRqSlNgHp9DwfbuRnLiCR9fvJP7YQ
Vwh+11OWkHtRqF5Z6IPV+OmSLtI2vQaLESInnDH5cLRyl+T3sUikTrP5cL7SlEVLrpZEo1zB8bRU
yylpDhMPE8G4xGe0zjvCCSVZ2rq1xWT657r404BpSbpvKRRxaPyYbgyaZbypwbTVHcBR7ZH/0nGt
U5XUX8NR5sNxI68ZCx/qWBFzwxNObTxsT80e7tODA37GM4xYUy6osHxOY6+Y2P7OqeXPK3xof6ni
Z+RulrSr3fJegPCZop/fIUlLMpcUvv/iXdnjycePPjOBsa1b54wazFsmywEZNNr7Uu4Rry86lnW1
kVDZdh1HmMzAfy1JC1aJ8mE1j5erNo8zF3ik5bepm8cdCn5JE+TOi9/p0FdL9WrmYvyTexPGCyPT
R8pOYJdHKzV+V1Zxyk0iH5eI7nIFK4gHEU95R9m0AdEkaYEzX7lA9qhazjz74EkFzwyoG5TU4PbD
dVAuw8jpbYS1bNGOQ456jRKS0Odchz7wRo2jnYsKRbI0+oX7BIU2/tYWxdgM72t352Fkd6/lkALk
X1LtEIjDSzcxDWyTBNqOgZpdjRBjPSSV8PalgJ6D20eOJICEoZl4Wt2jSiCuwDxRsv2tq18xtqsJ
Y7bUqkJtP4QXMniMIy70yh0IAQCpt3Corn2bSrvri0igpr/XRZHM8xfiCnAGqGghHF4DYQ7L8VZg
j5i/ybFD5E2Fu5MRJlO4iElSDN+DpSbPvSk0FszmxG/9+jKkhV3tny6IFg37X2wDh2rFo5b10gvB
vA1YCC0658GQqlQImWDwqu6sfW5KJ1EofeoDYihncCrpaYj+cPnE8b2xkg0bejL9h1VBsRs0llBI
6eV8xyfNUzh9xneaXtVn/i2aNxE2hIyQfvt1Y5V6mqQtA3k4brR1n72efXwP7ltpXQYajx45NVXl
oT4bxOs5EydpNbpa/b39535+gFqxzk5wfQT52d+XWBUYPQwWYngQ3pqz3ICn7r6FALqtVYX2fz1p
lnj3tFtDEA+FgaCqFrE9jxMxTa6yXuGG5rYK6Zx3/xBzHKiUyzOWFzGVz6KxYVda4wZzsYJAJ6V5
hYTKG/FBDdnaxt5peH1v9602dqCTZQWorOW5o6Bc+SqePTSUPZwIuttIswfw8Xu/kLXUE5v7AjUZ
WoiZ010IqXbSog+82lVuMEs8604pA2S7d/d0WGVFqXl/tON0jQDeGnI+WudcCikTzSXlP8ssNJ2M
LDT0uIg7u5W71+KQqkzEXKpevwQXvogtDoPHKeOHO4v6KQDZ1KomPErvsveutrpx0Hg1+3mFp4Ej
5dscjP1Cj6ZDywUnuDeZlG+AefVEr+g5tNkYQ1rEzxCW6pIJkbvVceTqKWuFHWIrba7bEyxp8R1f
WFdVohdGc+fF98rHNHotlY4IpNQZ4giXHojXyXPRa8JJ+U3quyZ9wePSmXUibiuP8W6z4TwGodim
qoSncUQ5NasoFKv55bXTjH0abLIOBhI/NWxCOXoFXfQ9UbR2N+VZ2jJ2TFXe4y7cpcBXfFOY0YXA
Fsvt8gp1QVUKbUl9srGQIp8GMLxkVxKMA35Ffng4zO1juqAvZQm99d1d9SNALvqd10Ucl2t9SnnL
0BWQiW5nldUc5jnkvfE6L1eCKBzIzKVPb7t5TGqBUrTVKK6y7a5UF6bmhIsCiERdJ1GwJPKq1U9E
X4vcSqJHJBhaKZFDdgulvHCNOvh/+U5PdpsATdL7xH6M/9WcAhhhvQtuTYvPO3cuvRP9F6UZnb0J
JWO3wQ6zyuOp3vO0ZUYeisDLP/ebmyyFq/iV/6FxNojQH088ObpSNTBTS9bGKDBGl4UZB1n+Aow8
A4vJXOgMBJip2cBI5qShIKP9NFUxNOFlYwIpzqAIGUXvq/SadWrwOqJYXHRqLG6anqwMQx0tsklz
j5awb2GV2eyAD3aCoc+froBG/SB6gFRSfX9g4ceb2yZvsurIjzPHgzckoRJBGUoQGJLktWMfmvHk
8uAf4Xz81I1+fnw5KXxUykx/ujIdJDyQRM9z+6rU3NNTN2JEA0+biIKVsgHoSc7tojJJe1vnWkp/
3mK7rXTE6CrZdY5j8okGQBD8oLxxS8Z+BN6Acyha6mvDKUeTxZxxcHuZvMVyey+pS0RRN3c2o5xB
SQIHcmK7YkQj1tRRpTX1G3MhT2Tk1BzjClzI/rAVnoUKcuol3wOM5j+w1CvaJZTQp63t21rG6brX
nLc0SNuFnxqmBxwohrfHjEjhazIU4tXDdd9eylwGeevGH6KQ0xxejQuDmeeM2UV7CVmhy6lG3obf
5oEPvco6kgDM619wdGhbyxxqlXrJLaH7C7eUj9CmXQ1EMJYh4vvXbulEuLPg9d82xzUohkgQoZXi
OagFKYrvDBkJg+GiYsiImvDqB0Ctl+gO5gfWIXp8Dv9a3nRoe31YIh/+TB1FNmP38LfDGPbu70Lv
/D2+OoEQ0xdkW6+A9YviywMI0kxJ6fRtHUwJNbAZKny39JGtYupyijthljEh1gAtYZhSg1NCw7Zj
z/EX/xC6hiMXE+fWFMg9WlTnlttwYHYdS3aB1N1zzRC4nVP8UwVGOCNn1xRJyeWBvDj1MXvrYPPN
KTXJvnHvdTXccMWGIf6hBlx50qRP9MdsMzXsxa+P/H5/LleMIUQZXCWi/sZ3hUh9f4iGkN/cF/OB
j1Vuzt8Gq+Nfw+KshZpmEoxdEW1O+s+qj+fVac8K7wL5jEDs++FrbZm2eDWD7Z+powvy4JCr3YMx
plls7HbvJwXeL54dK0CcbofyMCVv+0gm63U1Y/7xZdsJDsvvwCBm/7HRa4XlLABR2mQ8DB5K/m5N
0liYvgXtS1p6mDTJVmgIcq0eq6DtdlC2iaje4R0ICHRkEZZ3Ou5gumQGJelsd1D4bNKRsQcvZ+VS
JBeVlF1MR0YS22HVuBtTYYIYFa+vdjwxPn8lApcFAOhMVvwx3OjbFqfxCVi+jKFKtKa99sYxFdMJ
qQuicM4yfMzoh0PL3xh1otLQ/ZSfaVrtG0fXBzxb0HQ/9h8SmrcxRt61qx6Sy00wYwPyf6GEjHna
U+xxHW8N9yLTuazzM1T9WaaFZA9AzqJ9G+Z+j8uYPuDq4ce9f+2+pYbxdGyx+EGZdzUtE7i0WJw9
M+8HEo1iEHkZbzS8yGTECa3Bpxfnuwmzs56jg/EBXHsecDqsvY6jnahhibet/PHmdkcT4kx5dvd3
tVDfNVxM6E706ecD6Qii1dvFkTAacmdk1V5nIi9LbcB4TH7eWP0kY6uRnffYfP33Y43LUjnz428v
5kov+LifbfKEbWXxGny9Seu659tzTzYBK7+6WTPqmB0nF2b2qsEu45ReYE3ygaFi2+EkRkFxV0JL
clcGXAk3x+ZnS5v2IsCgFcHp6OqTUQyUP5UJzGAGOBgUGh7NQqlXvfipAUQ3tPpjjKnfXQ7RxDfd
KKg7Ud1mNN0pWBcPkJ1xwTEHR+26qwFdFvsHn8aDHuNnlBcmR0acVwd4LcKf9YJs4jDqxl0IcfuK
3TNmSQ7YzFVegKqlT75Q93iwFaIiHZW43KGTF6vJRMiw3bqIsmCBvzTPltzFCjGLnUaQ8MKoUmze
Zs5hI2E67OnFsvEUFYPshCqVhd5O54tIZpkOdWq9CNfMfrlvy1XSBSeX3xcxVgWyMprsIsDxNH8m
qcpfIkhxpiVBKRAFbS7gnN4d1UYninvIUNWFizH8BI6XP9LdVSSwa5rwdRqWDVfZYmcQKu/Jd6Cq
EthajoTonWxE1M/aFQ6e2HAiryLZ4xTsCo+Ot2vA+n1suyrmI5PmWGR0ggZ2RpIrJiIt87D/nzLn
+JaKWS9OUSdmP3wv5rl2Ah2BAI8WG/RAcrAi3KAjHRkX86PE4IhFizDpnG7/cLB+dtyv3YNq7dY8
j/HTt4EnoF633i4U+vzpdLUCsLntKePqqNIDuqerdzHkpuRDNkVKA+0l+Z6zxl8gfVuPcmEeSFjF
pJ2btWeUAStrCLcDN4d53/N7Yd7Xkb9MUB/Q5L1j8DGxBXBGL1HDHJTe5V4aYrGjagKCxlRm+zeV
/UcPOgw8lbEDvHhBB1AEsTDMWB+GgrU1iZGJsW/jBdP5mYonusS7uyKk6AgjVLqTkG3E5F5uTVvP
g4jPZ9iFAi84NY8K8MXdqvhdokPo4Ydh/vMZ1JZGgMMIz9EQpQBGUO1BlOGnHHJUi0ppzzNdT8jr
qDtbGlnFp1lMTAT7HiVlQ0glY/Dx5Atg1duYrPv8QBUs3eaw88g+hTcNwBwJyU8cFDNqrTZdRa0f
88r6y/CXPu5tAI7BucDkrOWUzt7FEiA+2bS74kuNxffwwYsG8BCEYNjN+XGiiWfIl5GxYekLn/1c
Th3vvNVVmzTiWeIsewfDMwtMMay2CY+DioP8wMfr1HzWK3gmpWnwc+32lZjuy2QkghMuPNxOw5b2
PiJ6r7e+0dKj2wamCldJbMRKRE3vQYsFCIj+84qa/xJvp3TmIescKrowbnDlCqiab7J/VgClUgdf
+qNtDK2uyXIHyzd+1szCDEui26crVWzYWwnur67YAUPUVDl3EpKWyiOLGpZnMHKJ7rweNrpupzlL
v6RtYnLc0BHgV8e+DRpXXo6cnkWyLSEyxrsNl/ZXmxWIrt91/ajxTFSIKVfQjQspm3zMkw1de370
2TPWXFAFRChnKE7nDjIhHhtvGYPJpBxjPTeQzrpenG/0Ama8frY5q1+FDCBoxqtfLOih2sB51zJV
nYzgh2rEjhlJJbTSBOkbCUCsLX9o/l8gUL9hfEivJF4jlHp5ZIAFrDrWDxIxWI6Wn5IXU3W8kmNf
+dzA7RNyQ7+2yziOtPe8mVSPFdds2KrFeChKzCa3eW6DGQWw2IdZbhBkbh2p3UYSMg/teqzUtp8t
F2XoB9l5wU+4VY+ijkJntmOMICvRwxyF8SqeZy2fTR2UAaGcbGJxmwhyfyD+dZ1RchGvPEPfRWNS
a1AU5KUyrWWnu2gMRaEPEt0FgfjUTF/kM50GNCvD8gYWI1jXIVSO9X/g18JEcCJe0sUiqex9/Bkw
bxXjFEiFIEG4TjROSDX7OwbSVhjbN9ID67ZDblIQOaJDkR/zPONHpZzrIlZ5oxVwJ/zG+DJuDqp9
8ys4jlQH935t8yiVHitqS1kp72l2F7h9TvP5f1rDlwsQNWmK4ifonQI3T/wYh5Tt7lgY33DjKTGT
ay0sXRE8yVltPdJ9DmZkWCifEW2yHzB8cErwfbGvPt9jr6AbQpZRRVuXnO4gEh6+0AG9daXFzqXS
5aS/9NTSnwVzLkhmOhyk2pQC/L+j3KpsurP9ix6isnXvnR5l3FfaD9waE8ym4ds10zHPNE8JVuhn
CDdFi22yFYbz178QypcfExW2K2+FI20dT3WQhr5T4wRwycXHKSO4A1dGZRvck/xoCdXSUChp7rzX
+pjOV3trhtncQQSPuIyeYw0W/jz9fx2rsogtiXXrWU9P28t9t5W0vYbp06DPF9HZOo/5QxauugGL
tL+TAj+9d9wnhD3t1SWgrNzJ4t65v0lmC0/EPAhVQ1l4Ai9VpJaSMe/q/0Q2Tbn35hZl9ZEScewT
U1ITV9u8XwK4efNG6DJHi6/FPwFX77oMlb7IWIswPmldRKjI1kWunIP1QTSrDlOJMfJsUlcQA0i1
Ke86NlIPgxPSGacqU/Lq3+rrf9X54r0hJBEGKyy1jbhEFMbDIEwuW+apf060Q6cDeygpRhH+O64j
vtpPtF7LOa4NfqAOrEcpeCL6xanrI0K9By+8nHDStjmUScmpyPP3Lef7VtN1f7N7ZK23wVJwkQiV
T6VOn+X1a30hGi0WGrbgJ99DOK+IuMjyarweYf+MMlINIcUPwT95v704f7UgOmD+a6HJG8daZeg2
xNnzab8skEcMRqDajZI4LnCwjboMzb7ackXkGWzFFCtgDiZSL/qlWjJ1WNm+/ARf5N6FcsQl/56Y
CztCiYdZ5i0vREEoGKFeAzeHz2KMqg7sPE9PzzR1ESf7gZ8K71DXfceB2+MidYd+EWtO4d4r2vu5
6TrYeQL0ZNYOIisOZ2SDP0eJiMgKtHJ9qMq2N1Zw/mCFq3RgURub9dc1wp/gOIX8SFgIoLntT5Vg
fTtwc4TX8i7MKEgwelwsZvUWvxFZ5zZs1tr5hUdGFMnrMvCvWymlzawyTnsdwwxCwU2d2A4I/mxD
g5XlzV7qUDj33X08RK+Jcgj7JPtSBxV9i31vrW8g9JcijdVU3l/6K1ngTRbWl8WfTnCmU8ui3jBZ
07wF9C7tWyjpsKNf94vE5kRan0UZsCBYvLWRpOqC5xR5WKoPT2GjGmL4352SNKgOXJv4D70Jcg1j
8B6zOOdxepWR8hIO8O6DPe/lqyeqCKJtYzlxqRNRGuyPekNIGklcEKSxrdSm6r+zzKgXlKtQL8Vl
g34qML5GMrsAL/upOOGTLZuGdTJ0KX6aFNB0I2lrCu/ntavxNyByqOV4vVNMqwVhqHfq8CVanmHx
P8JJ5/95Xn4+lyT37FRbpery4nCCip8nNAfBXD3Ke40GLAw/X+BKDUuH7+scoXmA26wRuTArKFid
/jgFABGBJF1/kCAM/fHhEyMTqySEgoAxP3Yy/C2rNhtBAggepkqyLTZHR0jCUgvi7cKWSQi+/9Ts
LXVCxEwnu7aqqrHnXbHhyhOrklgjBX9e2rqvSVvnMPe0m72rN485mtWh7bXrS5wBZ+OKwCK6W/HU
WdUq62Fw+IAWIkJc8xLBFNbQMIzzSwvVUgLr/Fbh7j6FBJd4cNZZNAoXYbmbfaYJ9QUrU/+bU2r8
L81WG/pnn1vvPz4e8qexuvdjzCLePTcGjpFAjLR0k271fpx9xP0EuP0IQAHiSyj+vPc1tMEV/pN8
A86M+1ygMQSz3auHsBdAAG9yMCZH2LJ2PfYKO/KF6stAcBtQjsI0A+glk2WaykL9HcmX7I9S6Etu
hVkl8QhnSJhHNsD2T0KiwyULIprCXTZ47EB6kcI39KDZ7sI0/bDCi7hVXq/ycLVtzZsVCfV+KVWt
WBaK9e+06UEqkjSCJkb6sFQEOAD+J2RbBivvT0kiUrNsDlTQWEwryVZZaA5+aJK0xfttAE/Lsw1h
kUL/nfvoAfJuDqZAuLWA/JcO3vHuKtnWs2ExWp5ucHy6i7YNgg3qEc1LiJHZB3vqTVVaJCEZnS/W
BcAq052v3LeBDc78LelfSdW9MvyR9OL4+IPu+7CPpdRXG4Mb8Irabt7Lg1zPt0A4Go1O0CEESj43
qOubIfA4HTtNluHjBngXRH4Jp47JsvzsCtuwJiyuJbYNFNNrFii2GiI7LXp3LgEuESPu0Nkv1acL
K2ijESjQVMFafr8hzA0mxu+rrmRO5YrYUZef97eELcN+LEM2oYOtmSNl/xYVvk6OgVW5r/rlxGzk
lAbrK8DOWEFZ+giRc1gqzWpWQXw5pxkIX5vAx9Agu91gGTSelkq1IrrMoTR7sFbY01HwSCFHBNYt
+x8tXkuqdMAQ40Twxb6uD4SZZUnyDpEx3gYi/DyCDCEA8JkrZsEiW2fVlVwN4g3FokGgpyFi+2lp
K7XFANTaKFIZuADn/S08sVE+0qw9VlVBJzcR6zC3awrjU7qdH8Yzgp5IGJnXHl2yUntL/bd69wJ2
HRpq2FrKAkEcRyRFozif/7HIyOIW+YhH34AHYYwWEQ1G1va6C8xlOQln2QQR8RdyJIP/We2uJv0A
rfh4nJ72jtFks78wez0HTYb5Zqt0xSS6y2KZZLFhHxXYFfnNvoUqh4bLo9jhyyt5Q9brPAeCIAr1
ydsyinYIhcNmJ00GiuSz2ZsvbyJcrhqXlMcCSd8JbPdXM/3M/SNLT2t39U4KY+ze+UHQMJvyZm4Q
1u9+coywEQpbPucsUGIYFKeKl/dj9PBU8ZadE97OK0nGfsQQusfLVFAJHesEyiYIX8J3Pw949Vuq
iH9JVuQ0vm5Pvmx4dzDiTlS4pKfMyGeDfn6jSO905VxKhsb/LT0V4Oy+h2vk3oWrNyL89pGP8D4K
Csb+fMKMfizBzE9lNzjEEHQ6e224tVJsCCY+bCKMcEIIHfJbZrqLJ6/P2/tGieKAl8B+/Jl0kRvP
gUrPEmnH8qU72zCxXvmkDv5xbGAb+Uo+prTyvHVreEctTwlvQ5tuLe7mL7x2HINoV9qZqhJFTMjo
OpzyduGIQRbGFD3SyfLTIj3fZETlHxPWTSMl7MhqC/GapOYFpivIv6zI2S8NrzUbqzwBQR88h7h6
DLHz05+f/QbPv/jaUWb8E3oH0WTKiGplU28PsIUS8YfvwSLukUSShFrsb0Xw41yLqQPvePMIhlBQ
dA1Q1AoU5XDU7zUoLWNkgqGvTsbOkdouYvXa+Jwqu5SBkVLUGec77LSY2blSsHyjS97n134T5WLx
RHIPNfFTeLDk6RDcJ9WqV+MpHZJGlh8lRELOiBefYmBhaoaPRQx8kE+wcApGBI96FBcydfLD0+P4
p8fJix7moYyxTQiOlXQCOBmVOT77U5Ina7Ca9f+ehuWYGY8IiWl+bayfo/t3K6gS/+s+CSmCkml8
Xg707slMOwee2PtEQxPWK9DOBndJQUArI2w+5jRXrR16+z4J/oBjcw187lEmQq42UUW3n4NsEWuM
60mJIjztSszkPxrlHmcFsRhk7EuhU/YLXNmG+FQP2SnF9FfTcYx+kJfOv+ezYply0aSnqDo8m0o4
P+x7YIJKQsHIcYIkt5JT+s/khzlxjb6agOpOEifv6riXRj3TjqAVPyHG/DpHP3wg5iKgfs/2PJgI
9zXUmHxe6LUgz6YddTfE8jpQsJYp+07nwUcT+Vng9KpI2CgwjyJ70yb4FC9VKuze2udq6FzakZge
56LsQ8W6oEt3lsf4ZaYU7/5g64CYymDP0X9K9k7EdsgE/ULv6T/w86HzZUZGtPn6Ao6HytgIRZ4Z
im18DRjuxfMamskfhWcSGLaBSwrkP5tAXs+erYpFyZ7qMfrpVpm91EBals6vNAiVPdKpf3DkAyuf
0tGwsDXZQEVUY0K2gRTQ1EZmY+LVpDs3wBRLaTYwRzYQ18bAdXOND+GWZcyMufzAnmd0LyO+/2Ie
MXKE2IDe9RrzE+Ch/gWZ/Vko03/f+8G6E63BXIkL4FYr2l51s6xHBDt9KGgQGk4bLz6qARAOxAjX
wlaDfz3z72oysOGipiXfAD5uFh0hxO8D1cz0YDh5gUCerYPSkuW1YdY/q0O6CJYmhNEKlb8me0p7
b5q8Mi+5Ysbwh5NqcVcJLjKjL8stI26vUxZabm5/nQv+TxP6ppFtOvmnEm2mDjvFDJOa3u7MG3hD
q2hPvhRjnxHy0Agc24FWe4AE2nv5iv5MbnsOaFl9L8nBRB+O29dMdGvIedNhuMxiLM+4zvwNQGBa
AimGTdH2CvJQAvgHKkHg8fClEDtNh7yvcp+GjuVx4689nyCERH+Jvi/QeFZ2Oj4mhh17zTGxDzRl
rRxciXBhekXwMvJr2Yytkz6dB7VB/PExBP7pAY3re/Rbj8PA4d/pks3bzaz1vL4MAYwEGC+AWoxJ
/PTUhiSX9jZkUHyeB6QN6SEKLCRU1MxIsrJbZIzq7WqWTwWwpnDNYlvL4dmH6I0sDHu+qWizmaGJ
2eKcQ2T48gdCxFzPDOopJlVNBv/VjzMes5WtwjOHSikz0Y26fxnodQY8JKBLbu9tXowV8SiNhtO1
oskg69cPwlmNCmN1cZ6lJdD4UVbb6fkOUKxRRT2ZIngqgHfvqGtpJiv0ffhPWfzhxcKUbDxPbXxT
APvx9rgVN/ThM/FzRKwVE6aPBSzAZBmac29NDcQbjKvG4q62qJsfQAWCi5ybmfTyfHiGawZdZ/aM
Vz8lNJzkHoli9lHNDhwtJUydcSTD13qvwQqHtdSRD6zrQaGP1ZedigSUzZter9lN9kOeeEJk2pqL
ZudCTWiwQIxbKHXsPixB5iRuT3abi/bXDROEsJctrDDN8bCkWgKuR6aQIfkxrkDJ3OdgEpuQxeXd
gPYzCUUnPE5QC8UR0NCHR8JOJ0jurmx3XFoQc1Kj53LctvbWRZgzSAwEcgl4hkNzMyxeplK6+RV1
cnnnNNgGutNNYLXT4CnV5AuYztCQXVgYrNhaYmzPNNSopnMQTAZGQkzUp8ZBwsZrCQ732XS+hFm/
f9G59OmwBF4EKDkYtpff07dGq3XpwDQA2YfJRCsZudLjF4excZKodqW0VeVOd1Asu6Lug3v+N+gC
Byxr2YzRkgP9rIxMz/ku8yhETHtYmgAPkM6qYdpH58FVM4TS5HYhKmP5p7Kt+tU5iQIC998+6Iuh
sNssdm8OC8bbMfTP+XudKdO/8MHkKdhwaxpRfo4BNhoxYNU4UeBr81qJhUU5/+7N5OvGY96Lo9oP
oGGhEroTGNs5bkEkp4MdGh7Jbk1rmV+Ea5WEL9pIkOBIX9kPV7oIOB8zTuxe0oN19Q5B7d/DqVMi
IuEDylqOqZJUkSFHeoLlN8YHfMcJkcEKWeP+UkoHPabnbf6qBm1LRJfN7iEVrV/Utfly9B/I9qec
7S9RPixFdmb1ZtDer7D6dd3h3jlXS+zoF+gKMtMbirxW0txP/ndWPDvwXzBW2Qf20FTrn8XRf3RA
3tTSz13wM1CPO4LptWdkwnYYobVX9BsfL/HRWp2lAxDF07H+T+fFqJjVo3p/c48HACfA7tY0+ji/
5y5cxD3nCJ793j9Lpor1pKHzjSuxnXQdndpDSkXLR0LE/ZNxrQhZwgSVdd51TQfAcvZgXpivOq5W
2SpN65nm1KnwJT37011doU4vN0Q/NFhu/dyRrFy0SD5HAJg3FPrTAsNbeaXvSA40z1vtn//6Lwi4
2MaNGoohnGXQthxhIta0KLsKx0EFj1fG90YGjMNQ9HCg89o2STqVQSf7LsCCbvn7A95T3avV1oCR
1s4HEWIDf3o7dZWKmkYBWLWNJes1ZjkZm0xC/f72WHTECoIl6ZxgYXRasfxo7fjm6x/sAoXBQdAU
Pr8HmaYYLHESVLPHxh7RwB+aoGVcsCyutQLrXKoxLOL7GbDvLk2IjfMdR2oNDg/MxDg1K8AO2y18
hHph6nVwaNCExHecqIo9VmYb2VWZzWSVoo1gA4nTL1s4O6rrEen3jgNiL17fnVdI0J1fntt0MKt9
UF2vSbwIA1jAKd+ycR74scgWYG7YM1+Ix4eQK/udWUbBJ4JetToUt6yRImgx/Rh9YLOkvdW1JnAO
KVsx0PgdRhbR2XCv7WY53PKnfqnDi5uP6BO8wUIx0GR3ihXzoYvJsMYOCtci6JkmjM+LQSJPZwca
fnwrOYIi52+1T4Q+VoXqv5ttQ2JGuo1QuntOPNLpoXx0qZ04Wpo9RNI/jMAEGTqhk8awHPb9yObn
bZGpMQHw92mmERSWyCNfX9429H8WoBgKnNguyTBepUoSB+XK5CdahLjXscKqeLNlpaDOwwEZKl9/
vsrkpTRmaf/jXMD/0cCqo+aRh9l22C0IUnHxeIwU3i8kTh0hlP+uSpccC0tMUd9kprfvx7N/A2Xr
vZG2rFmv8EtwEqAFRTQvCvr3K5YBJmxBrcduahMzW0FXiDnmtitKd1jqpU3QPXuHlEI3gmVF/CqR
ma3ARPwQNXc8lMb1v1c16YyHeuLos2NxhUUZZV+8wza33wvy2a1WfRhzHB/azVnj0YvCOHRfswZh
5Q9eZaLdJ8lk9kSRiuv+cs862XpVka0vBLiW3mH5MXwJG5+TxOCO+KK6FC29X6S4XmVtwZoRtzqv
BFcJw85Y20tZwfpa9yLUdAhgQ607bR2b665fOMCFUQHx+EQ2HGDV4sJz+XPCGisd3MwC3XVQRsUa
zu5FVqIDF3usaFVfXUPr9ke1qmRHYGbu8P/wHa6sBYpjal8KEj8VKSMDbPeuOf+bQArg8xkgEdW0
LcPm/GHSlbUQeSkRslzsPb7XDo+yxTvJF4ejTi6u8QamfkDzz2kFBusp0cxiQz7uyiI5JaLt5kJI
BZQEa/vJG6/MsF6AlnCKFnHJjAv2Zq6tOSUegvmvJKqxH2KaPH2DOxr2+fiWmUCuJuR05w5oSPPu
6lhJM7WZKAvxZ8xZj3wKoY7M355FCViHGzED191x7K+Wq1LP5TIzgknhwL7E1OI7Ytf/yfSZM9Az
IsWt4Ng7vhR8l4KmHnzhZPvV+qL5QgnPVdDd1A040DYXykhktXGuSmVAsr5wqPQz0W4auKkrqI6D
SFWqqCz9JRgFzSLWFj9JPlS2AzIJK4Q4EpWqtgbS4UJPHxw4THvMM9/pTAzQ9hdjnLVlwKIEeAVI
YvsG5rS2x1rGrf2UcMUzPS6RuojeiLD+caLiTJJ8gOJda2vDKcVdrd36dU66gbPRBlVBMln16tDo
AXfA2UXImjcr38DmOyoBAYMUFQPj4+6KfN/c9888E2LvMPOZyTruL0vm2nCwZ/UFofqI67oYA9x/
X0lQGC6gMZwJpAcdHRs8nCikbQtbXsfbt9BONlIsfld4ZpemMttNGRPrf2ogRPIG0DviGMRg4Nyg
nGZ1DSh91fdT3Q45u1zSQLyMcHf2Oms7yFbNpMLP9NOR28QWbk7jQ4mQ4z0dYhJur3RuVFYqu5bW
NPVztsaovucwopIMeUeGtBJ/TAfZf6HHJd0mhXOr1fNyiosq06v+lGyYaxtP5EokMStw3Dmsa+Mg
xssr0Ukwb/kfIEe81uwgnf0fSS6GFTcy8dzXENW7/fLvxqpe5ztF/Vke0RFrWpBPxYg/oNUuwNLA
NIexodL3ldHGbKeQbvqXnZAVpawNxYx/B/73stmhW7xYxOoLqXiaoBwHtn6533TD8/5oIiLZacVb
3D+7G3bl2ZJnnPIkkxh+bP1F6eEYkxnB83m/nQ6MN+5TzDtTeMWRHchEMo52EWpkGl/s/zxl3/4y
K0IfJwgFgbfn4WW4sOCGFEOfCeXuHu7p07WM1Zk9GcFaxnPr9VKf03mO+9F3lG9C/qXn+nzb0EZR
IfFjHvkXSqelWcj+7Xpp8+qnOU6EhUj5sgXUEf5zyy5B95/V5aG9Ug0zI9nKQ2I51yVtiEEkciEU
WymAkXmwuqfmwyV/qh9ESjPQJ+cRSNWir8vFesJuoIEzhJw8uR9w1vHmNoB3Jj6qhEYTPi1JTEQE
lbk3RR70HUZdzRaY2mDCWGSaSG5gAdniQJbYBfaA7DIiR9FXXSXOkzDTsyKZWXoR33EhD/ViH9Ju
NBU1ghpXKfd/a7XqXPFSEXiCf+BiZP6KBozQBD3/TZ0sIMzuUaVZaxnaruH3eiAFJDvQtKqQcjAN
i+i7kVc26jbIf6dw0jGnTg4DbVhcEhlTOSlOhmph+bNbMizclETJxfgPfn4/jk2SFzfXrCchkd9G
qks1hSM6wrGrFQ0TFf+QqiZ7JF4ucMJTb3dHBIxtJDIQ+vWc5qNS+myfBNe6Fz+oWkfhyrjCaiXz
g9o538dR3h1el9Y1hzkxkxOhP3JCjc2RG2S735EYLrPfRbvUpvq+zsTmftqmdXN+jDFKfM4qETOu
NNAztvxUcZaRe5lWsYzbbJgFLTVUW2FumhNWUI7Tdu+cx52ZputykuCFcZQRZXdbGtkZdGND+H+K
Q9JEdX+PYa3fUOb2ww636AgfuxnZSlYBRHmWW3dFX6m6hMCh5Ew9lnVoniekZesaG6SNuaKTsc5A
KCu2zcwqRcGlrroKn4MR/WK9xwfcR+bvQie/At4++P6VVhoFsm31FtjY9hbcmZX4kAT7zh3ohNu9
cd9HuSQ3IFqoQRS1w4CdO7j397qMVIkmzEYAg6/GADd9qtHgbzijzAPPuwlnd045U8qq/ghDX3IT
yijam3ng5xMinYh/CrZbo6Rxf/KGyEhLL1KGEjCjeRhMbyfKH1iA6VDDSp5SfcHlqfHFrzFfcDkN
DNLqR91DNGceS+YiHrTyP2iX5IgeYzMGLlrXaufp7XTfzoDrHm+zxJnAhhKX/YEHQGzNisETH/f8
OFxJvfjkINvjyr3LtkKquBuDuYXqSHAfmHVUtMOytwCximzWEGwWqS6zKAuMcIOF5aNNMDqoxMyi
1yF9I3zJJ8MMgAZ351AECHa+7lzft5NO2A76nA7o4olorXFDJcW4t1ERa7vJ7IstnKkXYUMB8Nsd
dPIDFC72sx3KuzItcVPuVOf1JSe0PIDVqPoHK2C7vpGMhgaTxqcg3hmFZWE4Dz4pNR5VDM/nnlpm
9SrA3pFic7ZdRB1kxfexwIyQ79rcWDIcUY1/Kh2TX/lWqWyR9rQ+McM2wRTyyqCzB94Z7hwdhTDc
7rZ/BmnSYd0BZ4jGl5EK8VpAAN24lr/WBdmAwS4Z+wh52iWOlDpcU6N/kQFB2kigMWldzCfC4SbI
wQZkpOMlEqMXBXW+LDpG+rEGfRZP/x83q8R2CZvbjk3IHFjDEm03gljMwFsByKVWEuj3WaNLaiO1
xXyXazrth/XqBF8SGdf/VPM/7qH3NCfEnK1C2vxYn4Mlmk0cBBdwFk8geUy5CYFGiTbaeH/9TUko
sNfchi6oCTs08wPC9GA62pyGfxtRpw6y8cI4VMiKWA6L2t1h1v3EGyh/OxWU3UD2X0x4PUNs7QUf
AyHGVy9FC2ESAWt9u4EFb43cVc/VDiC8Ws3NaEbRCzQ6NhTc/YpOWzWBeqYQAIER35P3rAHaDUgv
/++bphn2o6Zy5RNAJTfEP/hIdT28muj6k6bj53T1xw2TgzxmWmbs+663ZjE5Ldz9Y7DYma26wz7O
pI72SznLHJkbMg2nQr0aAIuZ+VB3QuBjF6gVZdIKXN0A+oHv/qw0ggXw0JzM84BiFKWiyWpPkO2t
z4kVAS2PLpEPFjka2YBvucm4z5AFaLO7H/MSq7Duzqf1rHHvyBQ4xhYRVAqHARxWCWNaNHSdJqhI
uZnaHusM/rdpYvP3uqOODfIHZZyuZSDiwsKve0LdXofYiLOi+zA9cY7H8ADT6kOIcNj2yHH6iirH
QHgv8LaaKNpJraw+p/jjwU/9h9wuMUl5JRQ7dsA2nD8DorT+ZggDWzqQMzIsVtjuzIt/LzXxeCdI
N9NosxUi8dp4V2mxfas7i05tmGIF63IYvHJtV1w4c3pQ8ty5YuoTo/la3QSjhzl2fwKXn9sm4UN5
ZGI3JojGp8nAdqp3Npw+mAYeuZ1Lr33H9jrF0sz5lGikLlWIiNp+47vQj1NyPUZwfvt7tDL/5Iq6
7CVVIp6y88n2MDPgReF30QNl1eJcCMKxjzB2GwLnq1E1V0jd8ES37sxi7heJn2l7OQTH4afsyRVo
+U26BnI2+4sip1e3pIeZ5VXSfwtUOllCoWF/dEvh/Qs2Wr5i+BByW4irEWWNfqKy8I4BAUcPUhKA
LNxv52VYTjG7q+V/XANdu/KVJ0jAE3ZNXltp5E/Y4Y37GyQ5wbmAG9C7WMBrEjH2YvOUX9xgcHto
7xf4Sbh+s8Vw8deEbI2TMqTEwb6/ZlQk25FZ0BFPgB7xC0J7XeIyxxUofw06jeEJ2FDhlp925qo6
ImJ422IkW2s1GwsKEV40nusn82/1+fQmT0oOYpJpA2TXmPREVWSgyoAM5va4wzy/m8YBwUHXcB6D
s0ptPoPKsCLytH2xjh8vL8Yces79AkTIWosxQX7KPNnll66Ynkt33l8ar0ExwPUr0qq72S7yf7jJ
eou23vImFCRA6PsgxJeJ3cd0R7WdEe1LZDvvyNKq9BBD5M0n8rE+XmFl+mTpmvF25T1w0SiBC5V8
bglhT8dmT+shPeZfnGDKiK/9MsplV+KyL3vCdwYW3IlPq8vnatoYqVbGV6poNoj7lqcoxfCeEuYR
ZAZYuPk7iWFFNH5cPi6WZezSQ726kkmEyxsD8vqIzWeyO8UmU/Ud+MZ27w154OoVCie3X9Q91j4S
AnWX6oBpptJSvVCl34EwLotsHZxExO71VI4ISOKsBHYVcfzYQiJZeRvvN6+Un6hgRhCmxYqj66ad
PvsMh/M2IMdSpHmT+wWl6jwPmUkGPotQE8/9NlJDFY7qGhYB2E+cY9MXcIOEohqNiYgDSZZzoCiy
0LblWABKe6ASen2bUIY7wKco0QTbS10kEVJMP6p9TufVzkoOtcFH+b/3RaH2rL2TOxznXJrFBrvk
56EhhOe0e5GJrrgLVjj9ABKqx0ZuxIbAARZPV3iG1Jo+AIkaOxbgJO1dosUc1HZzmrdvjVJsHX//
S0gEaV2QtnCAGYvjqowSIliGH3I/ruGraW326FdLOyUmiaABimIFVE3xNSf5ZsdcyQGfpqwH/Nd/
3rEKyt5h6uNvkSZEssL2bArvbFirxTq3dI6JmRZzfhpgFMTMwltRe9F0W6qqHG6bkIz16ZPvy7/1
3xAX6Uq8GRxhwZYy4RwcfbaDDvKm2bJZALPieep3jvMR5BTCG6wcszClxPrYCz5CYpbPyz646Gm0
gq4Pmg1DDb0Juzd7pRIJT17L/QOiOkmbzB9JAHImHhfwj1fucy+yIs37+LbG9kLv4gsn8k1M8LdN
bvojHI38AU7IkYAQOkyN34xiA4qIufOVFxtMY7MEvGgAjGnFnzGU2GMUVLyCco49JxJPakY4gpqv
lYEvPWM+bx2TC8kNRNG12qLtB23Yd7MZ+NLnSPO5q86eKvM0ssk97uWLC79GvTOu76sNwSL4y4XT
QKzApNxcruP59AT+5jaLF+ofCmAf5wWNReF88bg13cp81ePlLrDSdYJnPOwvmVPFgy0OQH8Oxdoz
CvkNEN++y31RW2AicDzzbwS+2w35gsmKBxxRLtcknIbCaMmpwH3bP6wUKFHBOODFJlVVbT/mHSIv
wXXtRbLAvl9CwJyHEC6SPW0wZtr0NaHWatMPAOyuuYk4jZv3J3XMCupblwpQG1sUtRnxT1PX3Z4n
rd9RAnDcP547TGChOuvEVp6Lfr4Gmnv9inzaSbUNAhGhO4ZBrA7rVim4innOWZdBH7orUgnL8ubi
TPnVSlEK6EcJlmNwMWE4pU4fp2q3FBg21eDLmbl6XWtJEpDlxMXzxv9IbwfCtixwfdsKhZJwZ1cp
O+nrM8RekJUtniX8vjhGbhqZwRtZ53bd2T9XxVJvebcGdRAc8w/xmrxbYIsrQDf1qjK8qxsi9Ign
NLdoJ5D9luMdBvgpLWNreYrnhUo2OPozYWWD/K3nTSBBP+fJff1l/GMHeQ2cgOIQkvqCP12nGgXu
ROzbAUkYxpNu0OJxkjOsCyLs/5f/UPk9UlMT3Wi0SdKcN+hb/tnej0SVvlsaZ7Eni+KZcTxHOOl6
0EgjcIIATr57fgSnApILvj+jXL9PCyDQurl/wqBy8OCnz8FHZNn5LN79s+B4EweFdQtdkogXD1XZ
BHu2oH5A8vWT9vPB2DyPKFZo2SSyLQ7I0ZC4502vge196PKl5YE2WrTnjXTcMYyL0eWm5cD+ZYZc
RukjmQMokPubQxiwCVI+UdwN8hR1LIEoRMqc6W5CgbnGFnfvTpMGL4qRs3Oy/6ic5x/V/Z8dYMNA
Lx6YrL0gLI0pn0UN85hiWNOHztJauMdNCxjKZyGfiO+vkGda9JoLbBt63SoEiIZWCZOt2tuIkOU6
FXPIIOySuWWWirzxWz367kHP5l8hhb7LHgd01yafJhZxe9QkbN7Ri0lD/tXJpjgS18V6EvbTYBDw
H8ofL0xcvqleySSsXFMM/UWi7B8TwQUuL/B9j+WxdTxreDVlRoHgGcVglkrbdddbkyzQ4roXoRbg
aw7YCdeUBBBloaCFr++iCCjq7QHMuXMRX1LLB4o8Co76w7U0vjT0iAfmn+637J+YboOf/YG3X9AS
/PBbGUSrmRKvpnlTQeyWB2Y/Y5REM9GGwlwxrCAYJcWjeZV3pgF96DkJnBUeNrASFredn88erKjl
HNwt6FSXAcVGRF302YXNANoo1pfI6gUYsg0SbipaDIm3ZbplNgycHUqygy6BqZyBmg7B3fh/orYv
pDSCzc+BSKman+N3Vjt5ao/nO/dgEx1sRmOlcMRqHh19xac2CvSa8nLufLaZWlEjO/59UvoAPZFT
Hw++ssZVcTPgTnk/5xfKrylqgLYBSoH+raJtqjnR1+EmKLuAeLq2/Y9hgYgUBfKZXw+bXh+JZZcj
AJnvkZrdM+mQivOWtoD9+m8kLdq8yyWmTUi0OHFm8EX+ffSVI1M5jGTPWH0W1X2oJW9vketrA4Yd
YFtOy0XLIIXyFZcMfVTPG6mZ84Wm320NZ2PCUzL/WedPx6TL8grzANGWbp4wplYu2xRCR/vOIxgc
FoBvjobhCA0Y/XZ4dgyvye0XwzRhE43cJhbzozyOkePmAeXJWGmgFsE0VgiJy8yVq9AL5sVc+QBq
L2o7x/Tw672OxIdvRG/Mv8oG4apBLgw2uSIMD4luqL2EsG/McetUxOpwHldcuafhZc9/xNDAL0Yr
F4wPAiU/9RQkSIiQVS7wdQRdNIkib9ls1BnZKkT5xulJoAnV37L/WzRXmSrBMY8xbyW0C7Seq5G3
4pgB0Ed/ZuIHvxnc1mQSn4rcjnt5H/SBxNwel+wHY7ODV2gP7fa/PgAhOjP+Gsf5FBjfQqISZhDa
Y+9Vrvu79KNEdu8DBCM3VEmeUfQCqrbZZHPshDD1TB/6iqYDsAiWuGRoPRaisXQwMZQLtZwVrMNJ
ci8G/W5Fdl1tbDPhox/BkJP8q55rkax7YP17s7YQ9zF3LeiCHBjUG2A5f3zvPosNnsd7YjGsTHwu
4O0LTn6e+vKsxddqtpz4ecBwuRanBv6d4BjzxZihuWOBA5lxFfRze1SyjFBjMc+ds4mRKmQwCHxL
a30dNDmgxoRVe1eMHchSXkcYAWVKYotFF/c9dIn4CCY6uMkIqZOLDVHPiAW8jEv7grRzI/kcDIl0
3Q6A7Nk1QS59urWNKUSyzdqOkItM49MN0TnmENfM/AlUuBFjxTShFPiskaRxN//LePap2O08jgBk
D19W0jKo/Xr/izCc7C6KwdK/jVHnxoKQ+Vti/MGg9/BwkL96foJLczE6tfjS13poDRjPYl1i7ZUl
zokLskIG1KQ3yJLgkiuuoqCTxXCnUhOZ0Po0B1Gy4Kuq5KAodg8yTsLpex1LXXSIwNhiPI7XOYg3
JvIZIiuYTT7Yet9seLavKu+D0kSew2e+qSc3WsVWBXZgKKj79KSf7Jce4CFNaATEhhCz6SV/DYrL
O8tQ4S8miN/9W+2zoZ2hixtWi+DuYng7Kg5ZGeLGMJpicHQKTMfZA7u5l7tIEJXyKqddWUkKDmuh
wEJcMxSVWVsUqA3Mi5ONQHm40gguzUbzZS7sq9wvrXT+yKj4qyUxNR1bdXHKhY+Dw2109WrsGN/G
fRg5SBN9lKws2xwSczDlkDoUlNmHWC7l1IHE42zkFokH7Ea5+ADQ9CV28UU/snqy1L34olJe4A3n
IuEDwfWS2LVDmyd6oa8JbdWDPg1+JdAihNUkNV9w2KRZyunhb7Nv96sEcUifatyBJB/wktAttXAa
uXG/DnrY2wecNm7RX9+ktRG4aK4lzBpICPo7c2EMdYUrN4MSEQAr+DIrXFlv/wMFr/YYJJ/zJx3b
Abz8daG2gEMGMWzu4plQrcmKefb1xsl0Ei9sNgTCJriOZ2GvfZL5bfQRUdgnOZESxsiNieFMAEEc
UT8v3yU+RKNSgb0g+b5UNYFATxkeHo3CfRvaaq6PdDA5vtr2qK2EmxnpRtmQcmJ+hePmJWTJtc0v
6oAk65rsTKffIb5nTpX4ViDFN3LDpaZex5eSiqHHzZAffiLHD3rpZ7C01blMEUotyWUTEH1E1Owi
LFxZZuAk9+ergnwf/AVE9yOC1keErp/SCEJAa5VLG2rbSnS6zRvSfIHVadPUNfnI+M0/HARzqgKm
KvZq53d3JWHtlNWsE8soFet37YG7M/vEnFAzqpV5Ak731LloCzbYJ/fUR6wmjACcwISV6qHekCHy
SgSyAYFIoVlZFOfhdTNFKM2c6cjTNxOxJppPr8Wg420SQcHfzu/fDKRFk075o/M3wP19WD7ImsKh
C08ezTdj66kfSKGL2zf/q++un4oIPjKQnbwPBNCVkaZtskO1amX0OL9XrS+DlmAbhOYdJYrTZPdM
c0aoTkjSIY8exUfo24lO/Yioi13yvlp9Bm5+vJxy2zrdzoSDY2KK2gpj+lwtbj+joO0VbjVQTQY0
w8M0hnWgCw2/QY5r/a6iTfmOrv5bgPpVvS7ThK6eekoMoDXIJfGS+rbC4lrWAg5jJ4rmRNObLai5
uHbd7PSEcmUGOthLNlGTYImtwZu3Ax4Ur+8YNlEc2j29fuP9X+o8ig3Cp+4qA9EdfZm18pma0qRm
1LaFcLYMQhzVPryb5nrgb3cBlgUPViKpANQTwnN/iEviVxyE6lXTZ6laxzjSmCZH22IIomOW97Nb
RuABkIM5vOqdrSosX2dKBDneDeoIC6eZSHkY6cyXhMQvJWfrJ2rsAyKA2RCJbHzvXDihYWeyLJfs
4vYzTKkO+1c6ztSeBnWF+yggHey2qK2aRlwoSK22QwstOHpIaALKH+NdqS3iELmqB8/B7sYLbzAL
f9OZ0M+hpOANrWphPphzuLxbMwGzAuYkFzfT+JKGIyzYKCQ1OxRmasVzeUsnl925+kbFy/j33iti
rstYtH/gUkGQixGNcGn2IYvSfwTwZ1XUc4wUhsBp+51SOS2rAkCaheYvH8Z+hamCs+0GMzkm/32N
OsksFVeCWEv33r25t5Xeapgi70YxPM7RUp4UzkxCAG6d0pBztdVyzyJLTlJtIuGfq6F86nDF/yri
JEUGPtnSdRFXwf+gN/j1J1IsuPbGOG92r3cIWuAYnLErviINsWLrvwrbMpXLa/quXTym0FOIJ6bB
+m+v+FIjPxvZZ6rCKjPTE1URs5tOMO7XlG02GXQj9WANHzV/gTLrqMZr66wZ5p1neQt21jWjiVMh
EGAegALgOI+mtneMT/T6rpxITo+sH4UctdTr3jzWn3x6Ad6EujfpsmmA0kjcPMZ/Cwb091P6qcfL
y3sSsJ9/g6PD++05/2QONO2TO2AbHwdSBrQL7uIVW/hUpuDD6h+JrI8mz5rrpEkp6M9VmMYqTz/j
pQhcrSrOXo8QRf3XhZRJO3zcQkxo4oQtSUeF7VeyPNS/cXATMNAHU/CnkVK2HabTAtznRLXwiDcx
B37x16L4pYV4kixgvt5gaHpO62QJ5gO8B3quYvp8yLXsQALAGHSuokRNHaI2HZuNJeMiaqfz2cMp
v2edo3xteqWjoGIc9tvPdQ7zTwqYK7+scDegB5sPey+DgLvO4bBcJAAG++oIO5xvICOEC1FUZePV
Wm9nnYsqnoywhkBe1ZQBLc5toLR1GJm6FB2m4HdYLdNJAKth1anB34ObA7XKl26oHGKiAu7kGN3s
zTQjeCAAXsdztBdLF1qAz+GXImUGJUn5MO6tllOKJVLTB5YeO9x/73T8uGggTzEWmldrRlO8bNpI
+VGH5xWL+D6rs1ZaiXqMx3gnaL9Mh0E+5QOKA6MX1OaUA+/Gs68GXbakdDghPX2p7oq3FrBDLcfC
b9f2+w8wd8VbAIkSAtHWKlA74vNE1grnTzvWyPOp8QB4Ik04zynlWCS95TcZhExfchVMwFzNosnB
x1OanR2NiVxR9Fw3CIeGS/SpF9jFrJYacATyXn5MekW9JwHE4iYTc/QrE2OeLP87eOhL3Z7v1JFj
tXlx9tL3FpY6P9tzywysD5i7+DZmkNCd73T/+8RsATlmqLYXQ/sPRf8FRO0TrPEaP6HxHtFlygIW
xUtYIC3bhYAQ75/wPWIf9leHP5N3o/1fWiPDAeW7uSDXoEu88YS42J32ctmwZTcryXEkXIicH5Ny
wMiAuyALhyqZtTTssOtr+ypZHhiiwAN7yg1QL0z5VKEo/LmLTfqxsXnULLVXgbFKdc4poGzLgMj1
rXuwzlDrFxSq9SFc3UCubS10vpkiGB7U0tEaCXhy7IG2+TwuxO8iDuUCjlmw8TZAv3Q/iAAlb5Nb
/bsQLtehfJ4ifbeoHodgR5MbfbeFcr3tJjtGQj+ejPRxcmGofYdrzSJ0dm1iCJLATAJTQNNVt8xA
dO+HtZ9y29DHij/f4nYXbu0cx544tdCpWzyG2u0mFgtZICkYArqt+vQY8PQfgU3iBU/m5rA0Xffr
zgxgDHfymPDtAVRi+FI/q1m4rm0hDPIRMtePbcPWO4P2uTYbWpUv02UYcwW+NQN0sqLFIFTBqxu5
1PKmElKkNVd/O5hvEVUxFUYSqEK6CJgM4+gQjziB9UZEOMvkamasZ2imWER/3ua5lQQgiC/Ru60K
um1Xm+kzqEV9Wj5lwtCbE8bEUSVNPRh6gD6vgoFtLS79ysspEfdaVMITSfx8qpuWSEV5WKgb7zhc
8C0s8V1mMDNUYNSggM1qIQk2p6yCAFUCb9iUKxcnQZ3O4/0uX2MInf3wXdbIr3rCi6RV9R/2b1oS
O/THTQGJ6tjdQmo6MxP+r16jjhOiRKxQpSi45PzWalgfaXMODDE7/g0guLJ+2B79o2l8EeJ+x3Jt
o0SR6OTxTeZw3UJQi+Ofo3dpVMtBl/7uVpVtroH4Z3H7idYyHOMSX+MGr6sUbhtOrYQ3Bkg1wRs+
TLCN9RPvMDAP8OQtSBQGZp/PvA9MRkLo+Ad72XoXMwlunjxTYYXt/s8vfOaG+Q6haXmNm4X8NDLO
dMFsWlm95VBpMW1U5Xutr85gS5ELPL10F9IikDilrxFhM6sWZDVa3sEmT9rHmhaS4M+zZ0XxuauB
Iu9YoejzmdgidxLr+Vv4/vV/VH4zIO4IHOPbKb1UaAAm9MhQT/kTB5CTnXvJpeYG3dxKc/sgaTnm
s/BG6JMgja62CdLdc3lF5KJz//l2HK/YgHsvrIrdQELtEMbFJUP9kd17p6qF6DiMBfX+pmlOO32c
jYKNWT3eDEohDE6gbeQtAO2zRVZYuB3XNfKX7pJz96FmmWO05OH1/IyIY2BeP0jBS2V9It8mZLSi
9WSU2+P6vj1oxZYfo/3P6+dEq79TPwBqQDuxKoP1lt15OTBB3q5QawUjlRIuFBani50OKDC6EGFH
C2ziGkj10ByK9NxoiWNEo+Xm0o6AUQFwzpdsFgaAsf18QPimjikPuL+ThRPwU2zZ+2xnl+Smqn/W
w/QtcH74bS+RHDr0SY7PMBNndYP99lPbWTY1ULIDA63GKUqrLTZTScWSZT+h5qsRWH9BpMUJKm+a
rppKymIUETZSIGGflcBeGD9NOELx+cLokWVNYhqw/P1sRPNinsNTG+HCxwCR240lyzmw1xolsDnl
LnsFxAbenNSsZPSa3OETs8egYvcU7rsubKmEvVWypNgm2KQgUwf+6mxIPScOQBvLhUfpYFQGf2nk
BHXeWll1NAwfzMG+trpsA6soZYNWsvWzwOSXsGcMduOJJ2qo/rTI8lJBNH+l0bEykKnatqvDHAlD
/nsAZOthmzAFTaheeQrdJVLbzLUc6Dw3lWGEqFQf1IKPth3u5ynwFdxVR3IgDZWAxmve5YZbOLLe
Bl3nb9Z5A6H6x6d0dkTTgx23YiOwJdWkISqu4hU02jgymljGe0w5stsqeDxEUmxC6M14JBoPkZSN
MmbKy71NZsksc/9gXeA9MG1hytkAK2C+XoNOuHIb/M4tdI+iQmvMCpjPw5pZVMLTU5evor6qRlA5
k5Tr8An5ICpxRgds24DL9v6avfT4u3bwc5PXZfoQllIpSVqSIiCtwVuOXlzYzCbKn1wFxdHK3eiq
X6rsKmE4tEcqth7fdy2pOrm2maXKsSmR/M3/jkqO4qFjSUZCnnEEQqatTr2kMOmpUtrgJRzUsvpG
gMWlxa4ptib1G4lqeUgajGk0HbDQyJmpRE54nGVU1eWsD5Uo54Qusd1E85sdYHUJ3qQ8JsYJqjvj
a2aMIm27FfrHRdvC/cNRLBWVBCfiMoN41ngq/TsmjCItYysbTCgJnZ/BZ+Rk/avCYdCGgrW0W44b
Wo483gipdZZshoqCG24A223tlWmx18AmwLrwwht/6o8WcRcRqhXAdcGfb8uMUXqw0j0CSLiuvmYk
c4xxcrJFPoe5LjzbLuWNf2h2TFMvQ5vR+/rvDKOZsG71sa0FvNGVn0lPt7pbIeKnq6E7FQBeC0nL
ii8tPIhduGCdYvLqV4o2LlBJtvoUCte+pbXH13rWYJh4UZP+cD6a0xHh1oEQfTz0KpXNQcKGFTZ5
q5pizGx+rZtxAboW8g1jrSB84S2jug84MEvD7AXT89P1Gst6zXFyNVEKKa41aA+gUMer9HzSSVVZ
XgyLs9xq/qiW6DLEQejzSY1iFZuI2fANGGgvw9Y32gg/8hAyc9igr/vbJqHIFbqDzBBuS/jjlGAP
dFtYqwA7kycz79NRMJ968lgXZSZOn1bt1Y4gT0vI4ksVsuIyLJS07dVlonDTr0hyDHDRpXcA/Kek
CcbwYT7kOL2gWJTsz9OmcAMDCX5kGUcohw2PxBzN54lJJIKqfrWwTbicu34gDTLVP9n4jbIPoyXI
83sCBgYBWSZ4w5lhQkwdgmI/bE4ewBD11kDiuLZSSRzCnJt+c4TcUvAhFrZ2oOFUSCtOj6VSywLH
jyRuVv0lKKgWGHYzDjshhNJVCW0+Dlk68OBVDANiQqh7wXgx5VkMFUosEVyJfm354yAvX1+VCeYM
t27TqhljJDf5affNDUqLT61iJY8l91caAuKt/59Qm3cmJ3i+Mso9W6l9IcXKx4elzokCQx41ieR4
Qvr9SEIY3nfXlya7RDVqHCnAzrVxOOs7S+JNX5WcWgA2amcz96ziuAEYzi1VNjJhOg0GrrGwYqoh
lLoOrB9CKF3KLV5EsCJxI/hd585p2Uw2Awx0t/5CljObAqqOjn02i4SUk1lmxmHRvBrq1ancJi+a
TOWHn6nKjiNmAcrNEarq5XwGUUJ4e9W85IX293dN2GBuFnQ4GGjZRTEBMgf/g6DD12RBNXdZLQgd
+dTSNr6TUXxaSRCdOZAywHZ3UAun7wTy+f5DhWXrhH+Wk1nnFgAvsOCtUGADgIZT97ArUCPUf+Jb
vcDrrqfy2KiZAOLu8HVURYAPuedv0ZQdVJHHofQrvTJmj8Iq8iO0zeNZUE0Nexa7SMBs77fWM1ww
xV5uCHMdP9IzE6/oQvybVtyi26ZNU+RXkJnq0vSL43g2j9YK5S3MgqLq8h4jXGs41Hp8isgKZEXJ
lv76FgQ9LiH7DHkZZQvl5iPFTODfq9hHKJG/jukeppZdqGc4fU8Ec2iqrWR+Jk3jrEPP+c0uvsQK
IK++KGB3E8axmRhPsHp075JCaOuvbdnomHsaClMue+IT26+1+RZGpG4Tz4Qegh6pE7a4qLhrW+HG
cDqulVX1pSfriuDHPfa2hPZajR7vMYpjE0TVAENNiTyPxfFe+GaoGsRwbNRBBRdB3z+Pk/btglfw
cuUGKZsjMF4BJr7ozF6HWYnmuEBau/8Gj09vI1bO4nC2mCav9ovkIeORpZ8VT8pc8L79UP54oOIw
tm3TGCD9zNyg9d3iKeDomUMLQXLo6WAadJNjAlyASmH5cn1hF596u8ppyml1Aa4sbI4Lk74vU8rq
X1S0wHVS9Qi/xzhVMhoEkyZGaBPyZIow8e052xaO6owNKzXLsMsDpHI8bPSUI1TtEGRTlyEQVJTj
iKoh6bOgBYQc5vQO/tqmKV0oIAy1tBDIHhkXzFBUaCMDzkRYbpIJvum3b99FX9sMUFtjaYl96euU
DBbC7A2zXI67CKCDTCvVKOKGiHBwqYBl9El8fRiTk1NIUY3ZOC7Ete2l//PclkASS+QPW3sfZ1Bf
vIF1mAqAWqEnuwiWXf2aOH7ig29H3MZjImtYi9wP/EEtzKormVB/7Gx4S65Bin40ZicDassYMMel
7QFH3afhBLkflk82QEuZbz6FK6QsDDJuxVRdd8ExaVN3bEKiDixNCyOWrLFCQveO1pE/imN3meJt
hyoJ5F7JO2OwKpwPJOcy7kA2FMPzf3xKOonU2HZCNq4fkjX5bk11nyYi3lNB/C6je8z9EDYHIO8I
/c6qQW/B2xiuo9/jW+NlN9/30krNtITxt57Q8iexW5l1+vf11wD7KcVAw7N0KUSsJdMWdpHa4mUd
JJ2CCyGZenkAf3y2vQvTXZJ0kEz6v/iKEAFSQqjadilPSoyJM+jPI25gjWwq9ImrWN8khq10Ked3
v/yhlSteOePlO3j73N0wGtgv7q3DlTnunPmMfryev/TuMNBWXbQD8fTn9aYJw6xhR3VK8q/jo33y
J4FDgHFzgSfXWGjzP6rvVKl3qsBoGROelDKb9Xndcx81hcph9NIwhWUUv0KND+yqnv63acAcKlC/
GPNpPmyNmcTk8bdOC0YLw0P05faPD2F9AkVgfONiEKQOY6p8S4eq+wSSZucBYnVc58JHHKxurIIJ
aiZ6C9deSoi5h8UuebkMdJhi3JEAW0wjNsWwqsKPBYGm+DraT5g+f6yH3ZzgDm6pjXg8hVEf9722
t9A3nGu6/UavhfH5Ztu4R33fqkCTKAHeQm3I7V6tOPEW6vBSZ/xEbP8n1u/wQoVvBVHnldlodiMh
ewj+CJs8IWAKET6qYOhugWzTqtTOcvnykjcvAh2WtHg3a9i3rinv9q4/rHJkBDGq1HLQ3VWPEQ7E
kqJ5VYsrCKJMprYRzrldaw6PN4/nOnWOm1CNB8GDlfWsCJARp5RvqAwDpyzEkMNpGNBoSiLvbu1N
W6VR7Xslszaaq5A9OvhhOfYXnGCiHu2GyMtqZ4VSICxRlLz6hblPQ9WGnryUfyw2ezvZpC2dhDZ/
HflKxp/gIOnt1jdE5UlmU+VhVkQ+BuaPSwuezGDvSk/yfN6Ovfx7/PEP0d5LcCVNkIxUbVNHx+nT
GpxgUsMTbNCdCEN1vEr6VJWdsF6HGb32Hn7J5rSGqPrLvDZ4UR7536BwsUj/CIn0P/I2G6dHXlt9
dA4bR4kfF/lFaDYoqRqdwtUQzIJW77cpFlxxcuOXesk0kS5vjXz5XqFnM3UWzc/4y6Pww77nxo5g
dWB5KBJGWDLhRbcfIO3pvMJ4p3LuXzybO/mU7COT4byzw9QVQ21wgYxENDsWsSHb/ffETKGuGldk
blQC/ALbOE/ImeuabwG8odTxY9gmwpvFfPIrdt7TXc1/Lb326dioSc7KnMppiLJC8kf144IKqhR5
94lFwjSaguXwF7St7LBRAu3PltDMiVgfww4cpyk9EozUyTz1HrB6SMkuw7n/ZfE37Ey9EH0sto9l
fqVP7Tr5ZukOdEpzSGk+5Vz13NBAopwl673woysX6/4q3/J6ecrV5ovc6ynkOTcXe6RibB8Zbi60
QeaVrKv0nEdLPIZ/JG7UYuhh1Ov4pCMn6E+9GPDv+q0lvyECuaHut2W/aBFwbVehYg7EdTHFyJCz
6fmj55LwWWsGcRJWE0h9puTJhtmqFX7J9eMdIsI45UrDx6wkdTJVvH/lNnKlgCC+tsEES1WDxSiD
7LIOs3ObyxzuDXlMiisUUQQBZ0jUPRJWGvrhdsF0kWaD4uaNbpRJRdcED0g3zV4Er25t44yZpQTh
W/pbIT9QCDnJ0ne4qeHkH0cBebmQ6g1xm869u0dmJY0t07A2RNyJfQWfyswyrdQv5HeYyZQIXRgf
Aj/INYZUq0uY7/2LGkYLnPHoBLzyHgwlDGyBSCkUVqcpCc1Vchu0GYx7Hv63Q+6WolAqoa2SlhAO
DKRUZuO3UmDenCK/wV2qs4+kWjyF1PhMd98KIr2vFf9GFYm0cB1zBSXibOKen0flkzT86y0vBSQV
Qv3xoBTTDyJpwlL0WgaHwFYymy9f4TTkaWr6SIDp3tOqUKLIle9d11hWdOhP/GOuwAj/s9jjqqSs
B2lU6fpNf8P7pG9JDXV55L3P/PqztFTu2ydayP+Mv/hAWM9OpVuvKm0nFxms/98ZPRVCIBsT5AAa
6E3q7XqDyNR9Z83704tBjQMbheY6Ey/E/6jvwSD4frXAcj7k11pWERY5JLxVGaZ1np65iccRusas
AeAJO/5wBwcWaMNhuW1oi0bCkg3geXE7wTbIhwmteTjCCvKFBgddFGmLde/vG7zk3hhEvQMHhxMc
iPgO1D7IWBbr1oleLLuIOzX8MCn30p9+qy0ezA8Yyi0q/EKhzsFjSg0e442wzYJsGj3nhYM4E781
Czz2LLcHYBCujl5ie/3We7J2IOcuOT7+uuBmtYK+eYgQv/FARGlEY1SOifnvO0Sdw3iElFI/DgHu
/Pwc+ga9ZJ13Yji6REq5Q9Z9hBzOJep56yXQR7quPwqwWLi3M87pe1wZPBBYAUUcAx8sHaq/1lLR
m7jURfxrj+6RgaezMw3kXIdyIDqO4gqMcRpKyfRnADNtG/8HthdUTi/CiraTffBQqdhIv/EJoNFt
V+M0Ot8mievAhGuzYTHD3ejSDuBy9XbMokaoxA3LxaYOJCqAeYnj87Y2Gxn6Ms5RLg5iyhluKIK/
+xY+QYT3O0xWOxGz0ksz1MfdJpZMlXtZyuDJYTAtA8d2EChTAXWOQ8cZgFaszWYlAR5R5yKvK3La
b0WQW194WZAK243SRdE2HFpwTDiLJr6bl6gviUGcVl0nXDYdWE3twLBmisrzRafs/U3sflI2ijlL
/nBRDXNnXN8+MsNPywP4seh8dB5esQ5NPHFVK/YU4EsAVQKGPFqqwNiWcN15E9EBsiVAQbsWkB05
ylKwamwXYRPAWRSFSJMvxiZAtiRNxDfwd7W4tVERCGRhf0gLSV30750DcuNI8me/IxefXx/w7pjx
LSqbyXiyhYFBJrUGzyL78OFqavvZIS7nLa3FhEHYEJfousa62FP8AMHvoLziD6x5p17vnW/td+cF
QbYpOj0ukjEqwVEOvkKQN7qd5cBGaY8xDncsf/ngZTFG1F6RzEEMpLeplFvRBzTKnprx9YbDS7MJ
45CYd5l+YfjlQ3/HywSjfAl+bB7uxbxKIIbm5eremke3naWTDZOKD/iaDK4OChuqQe4A5tyMmTKw
cqNBtcYl9WS9T3q4J7pAWNxiRbhU9SyxBcnUcqo/NCUBHEnwPFPvM5dRhSca3/jqQbDmSxkjUEcd
WASVtx4tj3Yqrgs18tWkmAR2S6nZo4IxEAn92XuVmK3ZjIOlWjUi6VTTQZduWVvjixLAx60s9a1E
j/6en62Azrfc0UNDKLDzD2a3FzxYf2S+/9BRg/7QxahU0DCt9rK3gbPw+2vD4MolItbMvBQESt+a
0+EXpCOM1lMxxP5QpEnzsv92BbLqK7zsm8HmKpt17V5U+PtKBNRiVtEDVfaJ6EnJwZY917wFkJz0
ceimJGcPcOCLGCxExnmsw0s0mZkXFRzlCHZovCF6cfoVWWKlcxNSNeTlfniHrr3mJgVqnjT8vijy
riD1CGnAbRu1U7NluRp3qw/z3f2qntLtJMwdnteOmlTHL5rVBfLIHsoWVMnVt+SS8X5ue964fiXM
ZlBbR/J9YP+Ok3l6khmnakmLhznmFrpM0e5it9bnXrVZa9NVB3JwP55/mmeMO3Uf/Cbs6T+y+Hws
WUh5BkSgi5Ud5FuoR9cl7e7Xkb5MB4wd0wl2hW6VR9GS4H4yODBaah9zsFOxANmfBv3gwacScL2C
Kqb49lo47xeYgOzHkqsi4gZLu3TN1LmHeIWO5A0H4hme0ejw9tCteiU2VbilXfQoLOUASBwatGAM
5IFmDBCbE5juYIWjV9LjT2QVMjX9mInzzkaA4a5dmtr7KXRYkc1nxg2vRQFTppuUE+PKSTo55NXo
YYfirYGlPSvLSMzYeVU17CS/Whj9CLg8LmN4JYairbKesIGBEe/9vx3MGJA1/A+3/zncyaxDMdpq
JUotLi2+LpJDYa3YahKZ1A01MO4EodERZiAlNRPv8g3W1PzW7wTYLMKsv+lNTWEGdQdUQn4qHxXh
gbd2TBTaHaDBnjn010sVbY4i2J4S+7cD4NXUhdcrvxi5Z5OnwEdyabR7EwBqQ92GH+XG+gECcoXN
I4c/12gRhMbOEuz+uacX1ONLmOxwLu+89flIy2jDw57cDnK3vO1DvfJIBcFy4EjkX9PV6/kfBs5n
wuyOGP7R9cvgSTTPWVkQrfi63Wy2fzKmbRWThASe+KRisNM463wvgcYv0ZlNFpIGGw4Wbff/VS82
ZErzdklRYMhQbeJithxIAd2dEW17F7rYoZ/LaMjAAE015AJ/O3ZYHMm8ehvyuXwzyM+0te7lvqQN
y1lKK7s0ou3qvcs6syVQbp5GCGUC+XgE6TV5aRUNSEHJNty/PKwbUAsF5SWjbMRU+rfZZLQZZKHc
sMR/mkeHo1AVu2PEa6+5sW5z93b1Ozb8WpO3UDXwjWSpKtDteRHym2jgA6g2E6JFeBgYUywShJHg
28yyblh4TrGlCJQe2tmzbhbWAQY0RYm8m1EqPKuar4emtT5oT+6gp0zsd9I9dMI9vlZAKG14Koq5
Q30RppW5PqlQpnD+LipRm48jkkFFhUugKPdojgIV7h32vKhH4XSZTe1hhjrDx3Aw7UiOhSyclNvc
wi/4lnEck+GpetH+egOhtL1P2rWQKHOkjSnrCfjpUcouVcxkH3NXZu0j777tVGFTJ6FpiIk3MJ7G
vKytQYOjnj3HiI7+epDoktOs09YlxZuKIZAIIIG1n1tX14V9QVlo8HW17XONs+ZMfqND+oBwMBAY
x84TExLXe61ZpdVRdYCYPOE7wW1EYgA4CIJKrPYs7yM2ey0CjsmIFlOS7WMDl1SSq2LwgcmuYBHR
rpoWSf9XSLjaV09YYkeyOsWzNz9ZFb63/jzJ3rBdIjNP1O4aUoqp/jzqZl8HRo/l27PdQYFBWfve
ntNPhFlIwZg4tuxCmm7IvzoXiIhZvi1Q3SGILAVESTaHapB2bhMbMFBaYBumTEi//nsrIRGekOqf
P9zuymmI06KMeqNB/cfl84y0iIluWxOBI2DDrimm4GHoq+TXZ9C1EeCI6QZ9iK/dsaZ2E7vHsXB4
rDCHXIGeteOnKRlDcGZ1RnVvxANSAgbaMpH63aHbaT3ZIq0q4YtVVc/BA6CzcUorBvLgmDFpqS9R
MzFeCk9qpMJ/YXyDiCvGHm5mbmrFI2wwWyqeIHsWfqt0fiqUPKYDfJYWYBBKbK/fjMevj9pdjIs6
F+9IElEYE4NSCYBZ+C2EhWy2aPK7fDCbb2DG3MS4oMRzh/Eoy45bHPt/UzEnShaBV/mIl/hg7W1n
SLoWWu0Spp7FggleHy3WpmJ7THNn0HnsSQyPJZWvurUxZjrRjwvspJkIvRFghQh2EWcJcPp+XX6U
xuih9KKcu/iAqlO0CKg40jmJo/wBi/H4ycUAxUcD29ZGVBvIrOOE3rxFCavVbbvgBWo6lLfDTpcM
28GCyYcJAZJT6kxDORii0JUS1rcxeI0c7i1B2+3Vxo4Z7TS+wRz2M9foDxfuQZ+7MCLrPBp0lDQU
aPnuBRXCtQO5LRNiSPoMI6fJojq6iQzBJslKQUKc1nDt3UQvfdQB2cY7sgZen9JMgfd9hCPybHkE
radG/mYyffnlA8lbWGR+43CrdfD+nLUuEaBBK1p7vPbkp8XvzPZQYpDUybdEX2WzEkAePUalLsdE
tuIzUaPc022s9izFML6Rof5UvHtK5HNcgfqo8/YKtCPGjyPMl9jvj8wBEk2HlaC+iHcKQv2RQYiE
j2dNafZWQobM/v1KawFGjEKzf14T5/AsTjbVY/zBtNaz/ZqVC2Wh6hiNJv4vlctAxllJeCOfMpk5
2rvAVIgH1QJ6xnyWzfkNU5uMh7wy2S4v/107JOXTP8Toiq7KgGiu34FP5q7qz3UaqL8ZtXreXizc
ILNHyv9n7OY7cLBxg7CpjI20p303ktf0iu/eBoJgXp28hI1rUys3yDxi9UWsGE/glPNPzShhKuEs
nGwi/hXCTyl+owjXY1cwwgdeO+EjMEexP3bugvaAvUuCpU5r7jlhbIuY8zo5Gifm3oIa0aEtjdPe
lFbYEu/9QTYBZlYcr/JzkgD4BVCTahIb6gDL3fBOlGtUS8oz0NoZzP3DLUdgbTGV78eBAK6famPx
4IXHA0I78ksiEzs7yaTmHziQRDhFyt0QO2otXsS00NSGOHOT6/4Hbxq30iqPycJ/Tn03/nKPisWG
u8++i2VnU0wBg5KDV6PdvNgvmFhS9Ok3Mfv3OZwioGvnt7057lpPHvZyiuOL6EnjYuWB183azsFC
Kql40d37Wti3GXoT+WocVzmuzt5+KhCTflsBChKycwogMep8vD4xJtEwAp9McRyoeyexJumyWya5
xJNabllNFP7CUx0gL7+VyaVdf8wi07XgsKn4Tje+9XYDgVzGQsaZb++/aI9v2doMICB0NBGw9rfw
wH2nJrHAVEXsRg4HKc8YldlXlexS35xMoTuTtgApvMcc/vxLdkvS4baINV1KJPCyalQee5nyq9LW
DiPHnB8Jv1tV2K6zETc9wQKu9v+MG8rVx0ktMN9L4MwMHfcJWIz8ek9wV2rkLtPnemLD13ZSf4Zy
Ca1OqZure7+KpCJZbK81gUm8ujE52Ks5Udsr6tO+FAxKtI21sXIgRrFApk/REjCNs22oSqKPAR2I
MWCKRH2pFho4Hz/Z4r6u2DDPs1fyFQLI0vqF/OGPiJstQXZel2xVcUYpXQG6E6fIOcL+Q+VUP6d9
sYeFrLkAOyQiDAnY9C5XmLp21mlJ+W+byXh31m6YeGUt5lVSU+6EE5/0v9YFTtXRfP1NOEuq4oKi
SzPnhwqP6HGPhyNWnQUsJtwihNfojEvYEnZP5kEzgjyRzxRIuxgC44oGHteY12ifhCnu2DHcEIPS
Y7Tm4FIVBZs/Uj7tGxakgBC1TGIPO7FSpH3R8pe+6CV+drlCEfSod0CK4djHd3VZ6q9usKOt2SkW
bPQ7li85RuoWgRaxXYgCCfFeNARXtb7PV1uOypMjH2RQgz9tySkPF+MwuQ/OK62p2BhFooAT3tBO
1LPZbKafyJAte/BZ84MaSDTGgrstsWxU7tQSlDwP8wKqLjCZhXXsBCH4/MEbYiCsOPUS4WNcoJbz
apDdI1PyVU4Ya4g9JqjIYWf5+mUtCFxbpA2Y23730BqR3xjoNig1K0A8cMTu6SC/F1K7GmawK6/m
APiLyCkqPZUCWnmFpcbWodEkMjwpAl23pVgvOtBCa4UUNBoNld29FBNmpJCoMjCyBpw/CL3ckTUr
mXwuXE5s4IvyGrHGHBWqBc+sP0Z5sT+IBs5ErBZPLDu44bxr33otUFTr4dHUPk96nKgcbB/NmCpm
7w0mLJ+3XQIvTrMnSENhEBp/96POEj3nYm+ekh1zFuxjkXac6aL6//rv9mGIWhGxjxdyO/v7I1CE
Ve19P1LqeP/3ZYMjSxLsulF0OxrSwO67oHnyvzis89UcsRsRESxU8z0DR0gUps509weKjFWBlo1Q
K3SFsTZSJwwMmhaGrRpZ63HKZpfrnIPo56FFa+hmRdwMLtllZkC0TZ5/UYcJFw6SWBz2mDLtedoC
jp/6JEYoAkead3RjbYsjGvqfRydyDWiRWA5krq1hujQs9uL48LLg/dbOqOsGikLuBoS6LXcNHUMs
4Oyl3j++Qf8ycJVykHeTvcx+m+/qbTr/t4Rk3Qj+zk4arb1nl9BTcOfpNwwfmDBNMfKYWUc4topQ
Nz7lfGyD+hF7CQME7nwOCkl+KAyOu9IjIGGf332dNlRJLF+vv79nGdsThUu00ccdK6Sn2I0iDmah
3pWIosykPZ6LvRLoAIrC2Bq+iXGnf7at56ADM7KpmxsLQZ0xbuzrCAxCXshAIqj1GZ188Ru8zXrv
hInegS2SJg7PvUbslz6p/TbIM1hDr+UsoNUmkUm3UhRDHeQBH6gm2z3HAAudkgNE0zKe2+JdLLR9
EtsVB/AqLYlVJuQ9ozIB6076JzpQdYm0fM38GVcGluYO6cwrO1txR24mPh8m78VHA3f49N4k6lvl
O41OepOEcMYRvSa3sV4lcK4JaZCTNv/8YL6AJ/8jol1lK4SbIlfNuZ4mFAPglYszdLbyq81ApPNO
i/iToFe+jrLHkB4W7mQe41KsRigggQyNOt5Ux7rNFovLigTcZNNKAZ7Nsnmh2IRj43HnUntPZD6V
vmV+zVaCM3wjnXaR1Js6RFfbrNvokZJaQ72CMWgXogTQmpQsEl858na9q4+kNdeaX56WLEX1kGMo
YrTfJHz1ucEprGKXV8NZ/8jrjMO4ZeH1ZuaZ6He6N0Os2iQ4upohnq6t8o9N+ABxs9tWl7zuFUcY
ephsHILHUdu8MqwhNhWQi0+LsOoehiECRFPFJ5IxU0vFT4cLGhtMVvStsXNNaT+mIe/jpfrN9eRc
MyrA+wNE0c3FMwDlQrwcNdXYqDyZAJGaT29ZFieby14uq+4JDSUrYID3N/WMkP1ZzhpfwKfm21Rr
B9mW1RUz6+DwnK6Fv7oVlNihlWoUD+ewveSHH2X5paGlG1EUBIEjpmbW4rulmiNWAplVQ8W0zg1k
++PVwEszNwlmVw2/9tJQpnEOWOyXjgV3NQKPXXG5ZBIP868wDV1K00OfADhbdTpr0RSyCpzVnTkU
Ae3EG3VOs8LRuuCqI1feMgW9NdJG85TDdZ/P9QWgRcdO5MLkKUKUe072bxREXV4EIN2kU0aBFMeK
6AQOrAL9BloGvPKa89EZWnawkNvDR08TWJ/lriFYQjVAgaU8KMdKwZNL3q8n3U5SBSkBWbSKddWL
yEk8wICGL09YrD4gPRrVoNRKyqaXPWrLflHPqG+zV206TF4R5YXgAZUAVvalr/LAwvbHZuRyWM4o
vhNqYBWnA+f1V3/Ac/25QdQlYDovj3dtNjC5U+/j1o4fU2VaxKIPRF14+sMjAjeJ/3Ytn6CzLZRm
GQSQDThums77pC6Z2y9FIq9zbJnHssg5rXI2RLmJnvsJqijPcAsU9B15iIWhAMORo2VVD1cOHcWk
7YotOI9Rl3s4SRw0MpgVFE09R+jxsbea86XDKMP1/XW5WPESjF6MD4MUOy0NLnvylRdxoqYzr1qY
DQZAuMqN4I+VkCcA/wJUtDox/tRtmKpgx0edlLypDYevKeMpzZGu3UqLaFHb/H2G193RUkN3t1IF
ddYAKuW0PXoUAXuMGgWnPyLMGlfEEfS3Xa57oyHbIVIvMyLzOHSk3xrt6WWLGaSNUdXQA3UFIN/H
rqz9VrihVSPwtsM1S90ObN3B1U4hswO/gZlSJxy51H+YeMH82S2SAgvagtpz/i3XxjBHch8mutJr
02nSeXqTowiFM6XLPAMBmt7EUU321CWb3+/+dcN5gw3U9CmbhruYPd6oZH9Mw17vkbDX9nbiCzW7
xqSXteFeiTtCEA7jBJ6l3sbobtuh8lzq0DMYD02b8sc9l6/x7YZROQ2IyWwsrRiPJaRw6bfh/eaP
xypT+aIjxFGnc1X84yoo2Qw/gw9VRzPsJM1/q+WPHa8RlcjY2z9ojW2pZi6+dNiwC7080K2ndFSh
3/dPdTansNcMDn3Jn2WlzWYvNUbWGQYBFbXU46YgWx09GFmuJtNtth4rhl5f4EMCiDnNMD1GJYwS
PFqVNtsEHa+MzlTCnf+zorbJQMiGNlIzaIkoROj3dFlLExX9an4ur+LjlDJlsM619oBjAWuafxI5
Am4OXqbrS0g+mTwwvyW+6KUZ0XAJJd6ZPuBGie+Cwj0AH2nlmJZnNJ0Bg8W526EtA1qiJE6usa4j
mLXw9OIlUqiqhWnhMsxmXpbIOJwDf9W3UCocMwlg2HWLttYpxVQV+1D/8DB+jAt6rntLNL93EPuY
pR3CDsb28eAyrp1XtflBtem9gTMJfcxjy5H2HyzGJZaDO79BREEbDN/z9J77vcxvodkPLb6z1HUA
OX66NTKqxSd1rnoVvEbgl4GRJAirMgaFabYs/zdHYQFBc5vhy17WYiYxKZYySSv+YKRwxn7B7Xwk
Umu9q6IWoip832KR2/lsFfjMTxgjl0Wxe8UrTSaUPmLhCFGpgUTET9A1DyZUST8C3LwyKvFzEmLb
iNQd7Vi24IbJtYmwHVonasN+XBKAMu4BesAaOZly8KutH15wZ+CqvL3NO1SS/YgsN91ENgJg37l7
oHxRUIT8C19xrSU/6b+Zq5ZEM/nlX1dKeGsK7bqdq5giqB0h6MQGcYh33YBCyfR7+FKxVziBwled
7EzkRRuKg6ZiwNGeEVe8f+Hw3bujS56ufCFvHEG+ZpW+DHwZP7AwvHtY4PBlh0PMgbial3gkJpHi
Mp9cDlveN671sPEBC7yuPUPF8ll65YsQQidHbSAqKTrIy0EH3OK7GnQbnbf2PuNuQv/8/rv5AdnJ
2pPhOPMHE836QZZcIg7iYq14GNJiRLjMigC1CisD13ZQ4mkIQyheQWM6Oqw49OCKmZfB1s/d1sCX
8bFuiCnaOjxRLQV/gKkzVq446ROe9TqT9RFn0EQ5P0kNYLqQjoptLZir6mxa9PLO8Ygu6V2WY7Ej
bM8WiGw1905MYMoDdeWuny2rgDi98acuRX2bdaKaGiW24NHbbvDkU6EqKSPJUUtq5z6elw+HE8mD
v85YVoEGyOQqJH5VwWwxQZQf8DoqKH44Cfyorh7Xeo1MxqxhAsfjk+gBe5KmzqGI1hWTC0OuiPTW
APmvigvmA87fEPNu5v8eHpahd1nkIzGbsmw6QlKWpG5gRQgJs6Rjv53TQjKcDlKCYO8Xoo1oetId
lXBtHdSEdINDBLh3ivkplxiWz6dbUb0FBWlEyZOiNdY1Gf+ERb3yQG4p2Gu5qlRpFuymISYwGNPm
ECr1rch5L5V4ijJb31UjhVkqO1nvHMHWMx3gyfXwOODBWknTjonBuqzs9xVndRTk3X9SlY+2APsc
Pn7Ssj9Bne5skM4QIec8by/almJQkmPuQtsmE/AaxRIT9Xu7p4l7kro/9BUnzL3fGFMU7lE0Kw98
IEGuzQEICSMs1j6P+tk/yES3ZI3ueQ9Lljtua1NTCPREj6XaQZ0j1/RI91tS3/EeeONrartwiATx
ee4HCmbOl4Uuy4aHlqbSSyirMXalqHJLZn08wjTt35jgmxFgN0adiKL68VpaZ6yAENQcvWNb91MZ
CA222dZU139P5LNL2bWnwwr0+Az1K9aScUFETpnJYYjKAYEbD5x96PIqY770O34xSWGUG1Pgqp78
vY3I/cQCUo18imi2hgHEeRZbWR98zMz6AVaFd7mKXQfs4Jysz5RUpzv9nb+e/dRgb8FQN3Rkm5S2
PunbURNTPVBk/cF38U9SPcXLwy1FZ4w/X3kGTAC11e+1IdiWSakLWUJAuvBdm6RGO+ycpeLsJaAV
SX41fWRu9IsCZDotiSgVYsR59mLSs6LLfUgpglMQdNqAXEgRnSh8x+ah8Q+p2j7nZV6ffViifmWo
3ooyXKtuWobO6bUUar0ev1C17FJAQsy6C/V/A5ej5O0/VkwUE16o49FEn+iRv+UzgoNtlKI2rXjs
S/SdOuI7DTGrlG+xUbzyZxgJaanqeCDyl9ovQI+LbT34a+ZrfqQO3U8Bh/Y5PsUDSBgZifkCjHNa
kTlaRs0udWXq9PNvGlUCcTQg6NetIIZGVE0diPfxuX9jqogSrdZxi0mG5VTVLvus1Uab/gL0j5IA
OotDIYWB8AN72X4dxTNHyQQ2ie1owO2h4H0fjFGEixIn/x3Yy3C7Ho5zySggkqZhUm6A968Nl8f5
hxUM7nQqYHH8KIkUiPGgePqI8C4WB/jXIDlS1LdLsc2FL/Yy/c/IOc+f2cQVj7rTJHDT9B0ZRBXe
GTnw8Hr8Y7rMXuZ73k+tKdzz8WGn74jPom5rtdgX4zNXljbC82vNrpcbNo8MZP93FDcC3rkEv3Zl
/b8DU66mRgNXOL+Bnr5MRO55j0WwJ7ZXFfEk1IUToIiManKIeTWwHy1E1t7/EYVtw+lOmRMfByHY
GlANTjy5HwPEQ8cws7QZfJty3LAKjdWVSDETOY7aDV2FVq1Q1vdG1LG1nR7pPx3xfZ0WHWS01icg
t1P4FJRdsXnyXoIung1uVWrSeD4EDksop6pM7ooF02ER43YL8BaK73LWC9b7hH8ZRW5g1IJO9b3x
95pGgLHouIqOAedX9cxtgSxyOFL3YHqKPFmQobsj5XaAWzns1cvZ+UkMw3MM+cIqtL9VQ/OBZ1j+
L+vXqoXdAyHSkXR5dsmeMhqiH9oSzCctPtsN4f2A3gY2aVs+LDh0cJXBJmA8u7n+y4Bs25oMynlY
QI7tgNsYGpS/ta68xZPeeHqg1ZXz42yOosc0jpdYyasTsy9a1sNjqAG05c0HZgrIkJtzggiwUSPP
Fd80zOoGtw4yESFuPi0T6G8ifvaQfGtIgC+la4R8+9fsOnSgaYxnLdxhoDNctwUST+cQl4P+bWg6
3sZaQ+CtQTPagAMLYIfNuSkCYVANopsmtwXJEh5j61AddvPqVvuWXK6Hte8nbOdlSsKg4bSAT+p3
bGZxvZj5AXY9NiDGcKqjrKzaMQvImLY3GkfFdeWOkF8sQDecyS6T6dAV8AnVM1iVHypsYm0Xgauj
BQCzZOnSUndpVHjD0THQ8QbURKlHInod9eFnytrNeaCklnLK7QDAmBLbRhRWMTifgfWPonSyMXzZ
zSfL2/2U/ITIl9rkUgLETc2xBFT1V5V+BLdi3PMD6MxZqcgfsr5492/5WckebqxqRmMo74I+4wUg
9G0d5kt0U2WhclXw0MabVIN199UkNE3Bl6uotxQNibKv+CDk++zEuzX9mDOk3M1Zhmrobff4GIv8
8xFRKF0+tnFi1rY3dNnKbC8glu8mJyZ4i5Xi0tLP5MX9+ugiMFjeAKXyxFEXGRqYKqVtlKwNMe2e
I44dAFX2nsycWRjXEXtY1waUmjmTQ53MkNV8kDY2ZtW1LjByVvVz1Bip7R5wUBg8X3JN++FdLAeW
9xu3n4sFO/Eyj+OgiKrP3NZgMx26ldnkkqKpVLQZRScsM3y8+al63dojAVhDjxf2LQdqWWltv+j8
MLiZfDZ5FOPmiwFHRUyCPAvRr5UvAoBXYmN6Cn+IFdsjWE0fXh+FswGwGIif20SWyR//e14+0Vqp
9aID0EWGpG70YGWeLwLOT7ZrXp77YlFaEVdY+EJLb0WPL8GAOnrmYp/2lYzpycdsoFdiMseoc2oP
QdyEZg8iwi0WvlpUN5AxnWwodkfl3sIzv9tsq3B8oZpinhEQb0edE5a2UTBphRlozkRDGJQv5ZZD
H2WKxmMFXi0CRdGLHTwIrpLJQa5OfqGWoyiCXGrNqDWshEwzbLKxd1cX5mn82kutp2/gZZ/fK3os
nkQTbvAMbnuRGprNaHkTR48+hFMHHgeSQl9RQcILiP6LX3GWae4f9963WFWdanBgAQgDwWy2Zpwx
2zD/1Z+31+/2iZ75Rt2D4SUZtWKoxsxpNPLnBMhTkX4zsqyLAJwqf44FIJmpXWDnXRYISk1asF5h
RuxGus4s3+1PlqxaNcqzkf3yruHQ+obRISlVHcanlseLFfWRCm5RqvOggJ3xU/5S/EFZB7MJJD4R
npaMyGD355gpl9cXAzZUJLQCIR6B8OGgE9CtqnWaLxiyTByheDyKJRxfQFh6zb54NkCZ66ugdQn3
uTlIOGeWvbpaJpXXw8CBSQ7pzQaCDmt7YhNUA06i+anoKm07sfNzrE3lUFRuldHcHFsl28g3Iwf7
OUJw53KGIrSE2rA16hkLb/Hh36NzspPmxHynA7FI2r1jIN65cOI2T3MpDj48voxXUti6fAmXheiT
jHoU9ysIiOAZUknfwC0Z+905UNx4QYuBPJGU+gx56HzSsbFzDVNgtthv2tgVpMIhneo09u1ag3We
flQAHKVVLXvs5nMhH9X5VPEIpelnJeLMIVbB4rmsSNGK/uDzFOg4zHH5FfQpwh7ORiVf8qWd8PTQ
6RM060/+oNdxit0vhoPHBRZRaoqTfeBS4PGAcOkoYtvOmsvaji+q0ku7AbhIMiqRWVu+c/mW/Nhy
KZmIhkkRHRjn8UkaE9P/HRwaQQUN65AHHVIG86u/Mab5Gjy2QeketE9SP4qoAmUAiJYsEloA1bQ/
D/WPrgGEQ2gwNMMBVvd/yyy2vW1dSMEV8wZDWXgiGta5VNt+A2BDTuHWUvByd48Xa3l+rLMi6rJf
4O0Q9Yqmv8HW0rC1QGVR435b7w7nrVab/5LqUoee81Ndz/wSmAXYifBH/bDvwFn4efZyvmtmUMrv
7iVFM17XgpTYObYduSZmNpKE6QWgg63fFaRc3qQkPrLnP+uzMbzQhRlmnJufzcjNXJl6nT9TZAbf
opMW797FjWP8gGGATVQMGzmFlv7VBso2Q3aWBmXIeHXsilNAAKj8XlME5A9qytSOlD+8LuF4uu+F
g0mXrY/797Xvo3HZmZNVO79dWBY9S8yRUkjlfUt/bE3A/R7qu+xSO3al7w3mP2aGG9uvtXk6OCpR
XTLfLVZqQDMnMDt7URtT1qXYa2d/hitPO2pVKthrAegZXsUiGmvW9F4gEnvcplCBDlVdwM6djss0
CLtdpVP/H8wGflrXQbh5IC+Y8IoaKCdXyT89vxTCLTaIpWF+jXa6dEPMV+NQkOO9tqed+VgNu36+
Jq+SJGMh1YmpA5Rxw56HpbRkXJuuDw2+KI3l3qDDj1imqEw4+O8G/rVFeAb8ZsaN2HunqFPrhafz
uYinl+lSoQMpbkcYzbbSq7sqG0o8FasuvTApW8sIRO9U4I4h8d7LIYvlKWfvUEWViHgogzEO/V8e
ahSjboPa3vSfIIyiU+R5G3zSOkza4vtoTy5QXlrPUVmVeHtds/ADbxQ8w+MfDwVC7S0Y7LmxnX0E
QR21kwKyUowNuldafrZawTTn3px5oVm0d8+rjBfdZYrgOxybrF3fZYOWE/nFrO/QwE3Rl1ZT8Aev
e8nrKRa2sL+yhX4AlmbLDTrmcd+rZYUQeQiMfo0chl2SS0jYYQfpvXV+TY1DMC3BgkhGPDud7JZf
0LiZhjTHkzH3HlK9Cik4nWSFRHjVVOhdVERlawSl1Vugb/ATf3yDFLJ/AX6QsEThkv58hjCMNfPU
kNKDsOBLrkCsb5y/tzh5xAJmXKH3tZCqdkO6GGdkARZ4Jjjj6TTAhq0slIjfYHqF+DSi67J33pLd
2dIsIPodqIHNNv3a3dSHsw/ygZqvObt+IcuSTZ557A+oVa0QEesvF/iUtqieVDtGKxO3wrX1Aga+
FOZXTpGoJCaSnPip4GmIjoE10dNdnmKNkgf+1SfFvTWaZR1jWRCzNF7BOhtPT4/RVJ1Ckp3pZn1B
N5JwqMuGMkEVvyharnGUZHdnZVKa9lYDvKC/62KFc0Gq35JgpmchpNICGs5Vv0u6QqlgPUSigaEB
t0ZA9brGsUvnz4pa6zpbkQqQ6eDmPrhVoJKf0ab6HDSOtHlr8Z9YVB4Wi+cT+xTcHThbH/CoNb3d
HZN2zQcd+5IE+6WFxEZMoRcMTW+TpmrboTBGITKiayKJz30IKPHDEIy425V3JOxmuhMND9OYBOmw
Yn0my15Xlf4g6X6oFs/s9lMh3Sfm62p0Z5kkxkIw5dk29LEe3z48cEwxajynqw4dzt15n/NmqdVz
6PJ9wBvEwRfFHhJbzJ0LBo3QwDW/watPjrOoUHgyRClxBGSL2rfSqiaHCcqE/R0JlwJxlYDONr+9
5fW4lVKtuKp8XCG600iB4SPNLK6aut+gVlxeico7VahmOrn6zpzYPNfh16Dcmyn16TEudR8aersL
JZL2LIo0oZR06BGY3hyN3r+HpqXsEKZrW/rHVtVKVVeRSid2rjpkzaOKKfiVlGyA4UCgORJDtaL2
DyCYC6dB1mmoLCbSrko0xUn5g5hpnlmq8IrlT1tKRfSdH9WYUy7uhVv2M0PP1IiYvENFTVn93PCH
/wc0IhlLoTZf7fu2KJmx81TL1gumS5dJ2pzsh/9eNxpsdmw+q7DP7SLKbyzBWBdxRP1UAGnf0bEW
aBEprC2auXPX6HliEATil2svBQtHoz0v3k5YIgsjTpzWh0tOmmZtZe1b9LWUiy0NFgxVrdWNEusK
0FcekU3z+TkKzoHZsJ0aS3V0T3BbGm+ZzkF3uShBTg3k6BzOZy2caKITZcq02unC7+Avja4EszAr
ZSInhnU0q3yJ97yDOQ4RMn5QnWd0fjpoH851SN1tOoCP8xCT3ZOYqSdMnrAdMgGzPgshwaK0JZu9
U86EvNx+2iwei3iGqJg0LQrqkbZ7ma67523hRThszgWT081YdexM7OWXAMD7RBQzLLYix0G49hh8
CAXjMzw5jx9AvCLfWxVcWTRkeTu2iY9XzI/+WEW8T3qVwhFt++7a+nXalSOfydxaRXw4wc2qS/g4
doe79h02d/ICZKtMsD49dSYl1LW9sg4/ffkTaPIOGSD9iiuBVHQXshUJ2YK/3N4J7VM72egN5yCh
WGUg0hrBil5e7+dKgVr88yxQPVTg63gscBR1PW9vkzsG9XTgXdk/uox0EQ+oRaOEodBe8TKcMD6q
iq4cBN6+1YWOWCHI4lyYdwJA7hBTy8a4dFydwImJLqwpPLg+zxYiUNH9bGXxAgVsKiJthXTS/8q0
N4mrpRpfwGU7tBWjDBdX8wHynfYJmiA+cf37qrMPZLr1+t/GzAvEThR9gVJuRASb29SiVWFrDXnp
6+/43ugaQIYpnssySQ5o7xE+8QImJ4mevo14SwcpIJUBa/cGNigiNp7V2pb90hlntQnVvyF77Nao
UW6f36lF2+lh32u6/ANsEBcTFHr/7weWnCx/XvA+pKenK8Ml2WnNdTi655lAGMjBM67NTZ6Y+b1c
3ZSzc3qCyXMSsf1MeKU02QbQvuqddCVEG6kWRWElu3TFDQM5/1V+T/3iJmNilOT4fgh7Sttt+mrj
+9PlVdI5dMFrLfjoQxva+83WPPd5W4nFYydwVYFMM5mjeJ1fM9sG/TrftlS8Tuxa4D6Q3iQ1OCrk
mVtVzFCaYUeOct7TJr5NwD2hPBYoR+Pka8N9jTb658rjrkFB612A7Ajam4iPdatEWTsgdOfgOa1y
oG9hO0185JCtbwEtnWdIdSw+WprfJ8sJkv5qHGuRkpOXfrsyA3gwZPRb7cXGMtxag+pM3lHnL5H8
zzykDtbjfBaOuyVjTHCfKas4rGNIwqZS3uTx1Wj6kJ29gYk7l9hrFAxDxmdHSOP03ZlYddtamIrM
rkT4GPI89OlvbNHZH0X4a2XUrXhw4HOWidEzWCFRxWFHBEz2NLucSBvgh5RUfxG/RmpdCbRfvGat
AfrycW7Vr3wRSKH8AIlE6Jk4LKNWX3W7EFD1mfpLkrhYDSEYUhHXhTOmfNWLTl7MT16UyRyGI4Fb
seZXbMPDAGn56zqefmsV6+KREb+cvbEGRf2Iwo4wmOqYRWwTfhNlCNbVynXBcAol8laZLTzI0V8+
/q3BQ0LHJ6+grJA0oXbwry7l9XNOwXiPX40HNvIxxJCP0ng4+4lRYLbsVX+fcRLqQBVUaPCebQ8e
fNlissWpkxxsNZs37EcyD3hqarbBevVY3pC3aZ9Q9RCRLWuiDoZjwihLX+yesxTljfcXUcqMNSBx
9q5Tb0o5GaqMqF0OmjEuZt7fkEiRVYH5whhIY3phYuHoiKE38NdKnrn5tIXBFWX0+yl9VOQ6PlqA
6fWbA6UanJ3Q7755obXy6iCQM/PMUdSr6uVoHHeLwTFUz8IKPbfdyiiBpxa1FqGJ1Bx0MZ1GqJAR
FqByd/YeF9VlLTGHEfQ7uJQBPTcrDps1MDs5CFi7BGj1eJ/+SBe099f5ZylOc30SLWi4+UScy35o
x4B485/2vjyBUQGiXGrWErr4QbmHqXTKGHR6agx7/yEtJfaVLbog5bIuYkiXsBGS4EDMLVPXgjY2
NJ1/S7a67DupPHXWmtilr9pY1eUrFrFSTEz3xFfY5dgYrxUIV8+5oSHhukHvdmpRngzgzfGqbx+U
Vu9Y3jTZ5KEyE9MSLEga99evpuJvBd71p+afmnTi89LQ19K2SxmGx70aw6hsYWIkuQVhZLYsJr1A
Q/XbsKa7x3KKOlHKDqwc/jVl1k7NbT4hfis1VoQa+3R6REGvwkJPhz6+BDJU/ftOSClGkGUgkD7U
SmbZ1dcH/1QAdE1hlKGfcrRocZE0oTsM5NiSoDaBK9MkJp4mDeFKqpIJZDhRtGdYTVetw3etJb+p
D2fkQbnOP0nmAVWY0WeHhVlwK+5HWkdDQqpr/AaeL+ncJjPPIJQx2+C/Fp/FM7J9xHQzLEeCx6bx
ifNAHOyWJ3kuLk1kbO08AgFY89886K9ANVDiycFaKMWgTCDyYAFIdhi72kjhPPuhnwSYzvzg7z3u
zLnr3+1DeEeGQlyNG2DUiBEmwuRM3YwgO2xBFsBjgow0bKEjCFMJLkkgHiYWdM03NnmIkQGIVP+Y
WqJZWrH5YOLM2AG3EbpFno1K7qS2c02V/WYMkyGo9jMTt55WqxjcP1qmnXAdotxb890LCMDxV+Dq
MkLK0ONBTB5SeeWodxjVLy0Oe6VFuwP852YAEB2yrzUTnoNNl1Blp+uSReTVHZggtivPAsgG5dl6
5N8nIdvO3gpV/5mkEN6fplaO21iwyPpxaHdreN5QGA8w1Q70wXrAkX6wU+KWe9uaFciZPsq+MjoK
0aex1ButhJRhdXuNQBLZGzggPu4NF5J34qrmRkjylD6dD/eArnWCYx2TIp7BXs5yicFeug+4PngI
DxcZvqzkZOJyz5h7EeXJ9wSsYYqPivlPAzflwMmyqtuODplPA0Po6R/eq8PtqhVE1PPhxFdYIoSa
LZknfnQKL/uKwgr5PPZK92wkqu4mQDuxLFvZEqIFIgwE1YbP5exREWiXx8TwEKMhtQn51FwfEqAN
ky5NC98lTI1MIG0ebNvjyVuerOGgfY5vmoAo3iLivX0kYcNweBhq1GR+8h4V/BoqDwmUOy5isvD/
jszTHbbBm1beLxmM3KbP1Tlo1Q3hcYQS9mU5vtxK9uT1KMAdsqcqFSjBqKFEM8hPDBfaAbwfeahf
BCdaNfQaXgiGNW9tzrkdZbDTaOdIrPK460aYb0sQbMSNk7wqrlX/c5VxyhSx38OrByervQOE7cR+
PxNXPXJ7de5VFaZ2jlVJk1rJ+ZxMr1wgpiWIGN4Zh1sJFLCzGq4RF4KztjWg86Li8PwT6Nzc/z++
0lTy2uAZks1BaYXq+j9wLtp+l9AYRwNgL+cFih5ZKNSxkVBlGjLsec8TZRdsrEvC9BbJdgl/qB5L
rjUT8oiJ7VDSPBo6WjvwfQOwxCwKu3T13qOBdklhjNUadowGqmDGDGhqFKXsGEijOHX75D4tr/PA
CUTtakLnPCjBakmeCc6YXK/g0MkH9wAdo0tcs/L67ZL3q8/InMsmfnQyS0dAy6Vo5wF3+S9bzCu6
YFF0C+m4flwRHYm1/080oMKVRV3WZwo1O07eC3CZN+U5PEaGQ3TyO0OOzTDJnVsp3x78MJi8xVro
ySVydUTH3YsyTsBn/AZgb5kLKopXzBAY4sJwuEz73iSh8BFm7zkDijNnBgytKvZQlt0L599e4L+e
+LEOcTtSEmuVxoS0H97oX3EQbKUrTSOQae9gGVHLbwQCPaYmxBqcmS4wxym8b8CrvzUaxsylQU1P
W0KEneACTVMLFcuolNPGVfjPiCDVGqTHaW4Zr2NAOl/AdkOyJgsO0nR+d5GnSSVAodpSDztalfLx
l7Rb0XKpM/uPUEV+r2rXBjMesZXkJqkjJfmza+FldgcA1n3pBTe9rrUGx/BxTfnMQFHYVE9Vbv15
mraHQnjH8rcptOzlmMVmiLEPls6BQncarJFTHfyIvhs/gt2UNeh5t0V+fOuM85G9Dg3uLjfOES/1
F43KtGpYKq6FlZfkGxfmIXyJ/Z6TITvTi2xD/a2Iyc0vBJswguPaTKZcHU1RrYy3o3sBThJ7VlcP
H8sGNObMkYJgltWMCXQhGxdrwkTVocnUpmY42bCw5WbfMfD5JOnGf7PGYxulB+yFxTOiQ6osb5NF
wi7lDGM7moCt6jgkbKWymn6PdeIxk82RoByMFyOdj/LW9ULZgjHNH2pLWYPVsrvgPzptIIJ50Rlv
QafX6wtN6roVWenWxtxuACnop5KVZNyTy8Ac/JnEjBsu04GaqZz+Q138i8p/5a5xCTRueuZA5WI+
lld61weByjmYG8+jo5Ta/B0m6Uhms90ljrBHtFJ43YmvFjG5PI8uI9PGI+Yi8+kHobF4WHjHowuQ
mBWAYhTqE2MO9wyxj0T5Li7RZBLXa8bkUCmqIshBMMxiBkO5XOFGn+cC+CmSlwrJq98qY31bT1b7
VMVN1M5L3FXfFKUXuPevNHmbzCfL9tjsMuxauhw3Fy72daY5g5vJ3swl9EJhDyjwNJRex57Hf0iH
jEms2OMbGfVettUWk4LfoYs9E14/csZaAhntpaqwzLQVg5fPAVrI7wPyw2RPsRM6Jhonbnt/aVHv
162t2IQMaJYLitw8szY1Dseu33Un8mEVpN9RdLUjbByl5LVzR6k80FDsmd+htObth4UaATvsoXGK
OG8UXNtAxwL4gWBk1p4nZr420oxfo+PmZxa196pUu2O4GVdfG7cuBrz7aTN6XbjmrSlF51rxAbXd
1zeLaomPm2XhlJhEMUcv1XMfWnTYr1EGsroiKdZMKsMIp0nDBToTBWGHWKZAGFy4mrNOKsw5SmOi
Oz4wkpwa7lj4ZrLTQmpxNqRMZvtFes72cIS55epWjNstaCkCOMv3iYOINDfFFSQI0dWoMGUbRHnN
R1Cnaga9h7GvvHGehg0lKOQXH4p/qcD1hzm4hFbLbpTlFVMR3EsSUVFYFJ9HyGFn0xOOhn56RHP3
n7Jb3uw+sVowM9SWXfRw2F+y3ZxYkFz5jDUGUUI880sMbyjI/yB/IraH2LAulwX+g7LjaXcCegiz
RKmqBFNCBpa8Gkf0IG5HMPAacxHJrwXlgwjaH+08v0HeluldT8GNqGouQ+8/6lUsS9y6lTa10CYp
jJ0TkmxydFu6eetMXD+fQ9dgeHR+l4/NPv08zz/lMXacNp5deSfu9JdDi1IsuN4KaGx0wq9b/rcU
CkKlGWjpfB9Woa1tSYaPH3O6jkHgOHd/iSQQjZdfXg6E18hhaI2Dd1mgbn+jGKmh6NQZtFIozDWg
wFQNRDj0N+36NCE1W4CoJvXhiIhiY8jA+rNs+CVM9MyKSufR58sae63jeqo0lRbhwtYhqcnIAMdc
Cnt5HsmHDF4YiXACGeXOQJPY1J//L+NqJse66pSfEitOR6RsrE01oPPGqKg7qe2DwXEVt6ISuaYX
t03iDbBNcX81a+Uc1X+9qoxjpzFPQbgWA0xiNvE9fN7y7nvt+9GkbWZwWaYp/uZOKHcbVn1DGspo
E0mMUyH1V4SSqwGJBBQ4Bd8FokqTsBj1u9nS5xQYYCTeTy+3+AYYk++aJgS+Z6V2yEpAlhObtOsi
ZnTn8/65PKnsGGFGR1TeeMsJ4KM8P6ZuvBLVoombB/GHNbSv6F3fURKEt4yNbyKPU5eDIyk1B4R3
gWgp5VrpGjUXy1EIWni1mV803suH2sloPRcYwf2v2fCMa1Tv9tTGx2Eb/wP2klTAPssB6HwdPmEA
kEir8CEyEau+aPl9JHpdUVhkUpDy+FHsTEHfl6tUtbz2M7CtoqFxXOxWJsNwv1pzp4v89JjLAulu
LzGGVuUnTbf7ntu2F9E6rD0+Qphsw7/sb7DHsh+qi79xkxnu5oY99GoXAgF6v/VwQ8uVxGCenTCG
ul10deqRoBSM0JFQ1E3T7RLCGCXq+uGNoxNi9rx1Rvct5c0K5C0dU3AepXnZMzt+K12eAMytFESp
U6/QpZuugom/1lBdYU0B3Y2wmxn4/ORTCDuXZNOGWtAjArQ8YBn6sQf7X9VlDDIgwyBKybpIQ0Fv
4tG6Uj1PV+7NG4Su9guTmLBHo3qxyGvVxoA6CdCCVZjiD/zCKWJvZefvN1IYcD8JXjnua6FUCMYq
KcfyB9picPyWwyVqNeGT7Q5MN+moQiEdVWL/meh5f3xqAaCaleAlwKoh7ABF5W1WkELL88uCvgd+
tEpSA8jvsPQFCixShEZhFtZPHkMokc7CrKSavXZg4v/azr2RP1e1xYGzo9TTiRTcIKt2+bxGVvBR
FKCNP7iulOxMQzlzpQ/RV21KnzFjgdyZ2nmtXch/Gkb0AkPVAxnQ5U45KCuiEEhfcs3tjfKjk6uY
mIWZGxxvlSHyJqM43JbXzJoAKLo2vAHvxJHIKOKqMTR46DpixiSUbZfyv4wbnjmpoa6D4Yh7oYEs
/wdZdO/z3Q62A0nojAM39TOvNLjHGFu85dcpG0Gt+M2mlJ8UpK1+WZwMBz6J+nnhGhYgxNyYVpXi
Vfxz1OMZ9LrT9Y0gqxJ15611zxV6ssBZNXbxKj+LaGMHImI8OBtbVpUKLnMBu8qGdTK2loJ56aVQ
rmg8dm8I9qNgEMrYjYiH3sb4GupoINoFHD+MoqIlE46tHE5pEJ/OJOSBWvq+esbUjlBLTiSgRXF7
XI4xqg5/7FYpISpfH1VDV48SYjqyOSGsdWu2bP14S0yx81+C1ATrhIZniU7a7lNhVYeyvMKHDkNR
AD/I4WirAorBKFvNDoX3rD6g8ApQWNZy3nne6gjSl03dZZj3Eg1iPkLJ6XBNUK+3TiQTKRvSfKBc
qmt1EKaGpIbLJHPEtfXOR7ydnByuc7vX5yvNmPfyH/SPiXRb3GwYYIOWmJR1He4F42ZMZQA/qCYD
cQqxom8uMwbrnHczBMaAn73o1Mz8jdfXWgNhncivYDXdInJYWZ7LDlTzm+XQs1LTjK1Xmq3C89TC
btmudxhjOAhNvJZsVq1E/HNiFxgeX627qFptymnHjXfyvRoZJYnKWX3BLCF9j/BqNvg24pg0D2mr
XuMUE0JVFLJhzd+ocdf46Wgj65R2Mw4eZDM5MZ8KgM281zZvFAlHPXGsFVbXHopz4Pet2HGVjSdT
wbxsRms9x51zGR/0X3xHARBOKHz4/r82+1VXrUEwEAP68mEaAEL0xHsmuJ5IxHTOBsNZJ4hyIFNj
RwUBi4t4wbOebb50LrJiXihkeU1SPO6p25CdSImGqNJrtRVicESH1drNJOsDayH7hl/MM0RclubY
TyqbLKuBo8c+5UejUhk9hYVvbbrKTqASGvYH53o4pZJjE/q8Jv4l+8RHbMnldRt3RMd8YeNL3Jo9
QN2pjOeXoM6U+mAUXCm6W82V3nEoIOWQ9GDJcxFqibHzpnCurU7qmwTcvhBVnMdnSgtaqoVT5byt
dYFvKFJZECWeZdOiM1xNTYZUqJcdmQtB48YR/uw9FFK9e+MVv+A/VNjX4CxEc2epfe/D0yol0g4V
+85ifVChYwp9Su8BbM/xYgFP4DYFAAzefdkHpIVLNIfhV2u9yU6xicRJCntBwoXDFjyfAPsA3vKe
6xTdZGZiiwgiS2p1KwLKXnSlXQ8SGSCfo8pxWdntoeKI20MMXNwdWUNVlKlfd5Owygx9MEqSMsno
DAuZGr6c2JUDoXG3hfwh2bfIQlgZQcaKpsBlcplYU2To4Ys8ilkobM6eVVeTnw17RKbGh5FETq98
GefC7t51q64uYaraM3g3adhyODZgPrNKx1PnXwaNR+IoBz6FzbqgLyjj8pkqids50J0/r2TGHCxh
TWaCZqZM8vjTUJtXvWjceSkdiWAphjSVgGGfyycrnzxJAkJfTJOkmIaromNABCUCt2rC1ynGhSR8
CR3WaLM1CS+OJ30dNcW/xMS7Hyl8fgqFxvReNRKeUEcnYsjBKzrFrMjSU2nMLRbdjwMnzk8OC3+c
b5x7IXn0jg4NHxzKfNOhKIx5sq5fS1B84cjxulhk1/im08ID3XE9lPNglIWt+UB3fmQwCT2n/BC8
+nFzRJzwfuzRg2gAeYxkbqeBZe1QhZBPucYhSLkpMJbmS/hbEl49AggshsM5Fqp98fivNliitJ0L
7g+H/LV+6vGjsZxIcmWbT5/AKt5FmNgMahIM1FpQXAcUMwH/fOG2G8A3hEh04zkspTZhG4eMkVs6
z7TXAtvnFKaXQDHQXNi70hNzaT9Q86EmDCSytmoR0Yb6r45mceP9VN8eLpcPaFsUd3/75dplxS8e
NEUK9lAr0BUwvOMngKG475st2kCTR1HXNUFITGckpvVPoGvcP/Y5lXCl+vPhcu4T2fGADbk4yIuN
A6CF1lhCiVZJglmRdj+jLFp5/bf35XZzViDdt1PLXBWijGx0mRgRfe36PR/XUoAiyvHwSnFQGWKg
Fp4IkipxaQu2wpr0K7RBV66RE1K3uuuIIthf2jcaQReJu/nJckNED3RiaESgKzumqHcLEOR28pjr
qBPGSl7RlU7i9HlFJ0H2ihbICPQodpQYBNu2iPOddR8jPLO9XgENS96XubejRPMoV0/OwOz7/yBQ
AIsuFB48ctN5R4WCNbPHUr2AOrTZ9L9X3I1qQm+PX8JEFKGIov2kq5ubggwiDnmfLf9V7GfvoiyF
8B6OA800jTTc2G6RwCC/8W3sQcyzXBlj1Q4RZ9MCGJCync2oBgvmJhd2Cyb+fQMkZkpLpy5dCc6R
slgbocvs1uX2k5dVX9sah6S0DrBYN3e+LbipggRtVA87Sy0N7/HKFXCh4eY6tfKirAxv8MLASpyP
IiC+I66qRNbz2gUiVaTXf5WNYX+pvvu1JYP/CqO4LVzzdgynBRjofRAD8TmGF2MFjYKqeU69/fb+
akN9SLn3S/YyazwqMbTLF4FO1ydi1OJTTcldOfnpHbRdFzkuzqG0l5/HuVqWn7YfYlwHm4IJBelE
v5etjnEZzPFNRCgw7SQlzDQQB/0Z7Bue3gFFNJy40DNBTATTDweqPIFXsGzKUWWF2pgAxIFOkPpa
z7GekFyxpfC40adJSm+s30F3B3JvYcF07Yb4QJnb2P+2EEAcFaP+82n3Oj9oU/WrKVHLK/eAtNOz
2D0GZCIAyLGwE/wIwFhZcmKObswMxKTMDOaoHUrW2lHOsy5jWFhp9t/TUfWuRhZswHftC03zgR55
uKqFNSiT8ebM7zeEtYXSZB7weuN4O8+zC9ibX7Qqbi8cYHTz6NhaNO/rNtr8BZxJOQpdaDjoR7VP
m4kPr/be2c/Dttt07ierVYC/BjVw8SpGv4RqrB4Fy0xJ1IdyuSoONXDqeK7lUB79Q86wtLtAFC9k
HZCNtQXhObHEyx81d8d20iiKQP8NiL+uYL1+wdksuv7AirKcihzFr+NwJISgVa2LpUgRTTfKRzrm
DUmqvnQ9jh7eSy3SR1y+2pHkI7s8IdW9wqI08u4ZhfMFLtA95R5MofMWZdP9dDkluGQTyoZje8oO
EcH6H/IrIe2+D+VMS+UdPsm54jCGLq1ZSXOA9Hg4G0V+1E3nBm524VaKsah/1L1TnOufp5l3njiz
3iSjhiVoryTJJxF3NnQSBCmqTLgddJ7qWKj47iaCnrtT0nIGTkj0HUI88OmmCM/YcRIFk5iHDOeC
dfjGx5h34hMvgwaZMVSFlPKemLeBiQvZpyDLEN4mKivcl8BAvF/s5tsFqNojNQFHa7dMMIboE+15
y1vcoQl0J42a3TjfLIDo/vvVl/ia6NSBbCpvJ+cagLW0A18ymco/Mrbhg0Y92L91l+KXLYzYWPvR
NxzzGlkdbdYfsJBspvvKz70zhmlhpoJsqQA8VzNIBl8/KddLW1lh3G92sIlve8tT69Zzp9zZ2/Gr
WxV1F9EBIndQK3l7oizFmfogivqRXeuYslYBcCNGCjVS2z8iM3iDbiUTlxbU2hD/u21bu+E+xfFu
f/oN69ad4aCjnds7u5cqhuCHKj17//uEd/pFagZpa8lfKrjGzo9q1SZmFuaZiYqpraihucBYIZkl
RCvuokkjzA2VjF98sjLdlULurJN7A9EqKuhRcdasPJHQfo0e1fcK/22VNyInBjlvUKH0+LwW/8WB
rTiDKGjQTS6HnXrWnYL1T5ttrEX6UrArROUXrEyw/au3PychjPkguMU8KuWSsvHn6nrPIAu4PoiU
q6N30J8Wuv+ZLRtC86x0qjpqzCaPEI8PEzVS/O5GV5dGJhdUCWkCuaJgP/Ftk6uLzrTloJ9jn0Rg
zfI3P5Re/dnN4RYgpnlWETFFKnpAAzdV+qRjG+ufjuJ8JjSvUagePIcdSiNzgBUDSVY9m5314vrM
so2iLho0AjEu63nkwOZCjzBRo/g+et796zn7NuPsl08WQK6/LLHrO3yBoxyEi++R13qtF9UBHXyX
+/DCRFBiwQFv9KAz9LnXe8qA+/5P+yj0Z5NQwBy9hheLTifbh4gxNUqaZa6Y/XgayWCpUlzuz9DA
44zBhhi1Ne9MkuGQhLYdZoY70gc+rnbzLWyZurhLhyykioLsFVbjzD1YDvE13K7/Fr5NdfZf1sDk
8srFetgyO9q1E018YAFVeLWEGkJM/wgHJSg7dEtMoMhJVXw+nGxBtKDwMJ0B1mrwhMHTtXIH1CBB
64tIBeHg6kRC9Ov+3WNHJFQMdOITM4MEip3Q5ZWgFpwCQs30htR7CItdbT3Kmf6pGGq3JW4XTyZi
MlwUtwylMBbECnBEdSjMyackOnaDzCrFVreTv0NOpJ3k/sw6Gru7ya9qEDAsl28Uccv8I7+kEb0x
Ddb0wz3qPnP6b8sFwAiBtYGxQtb4HUakO6aX+vknu9Jd9td7nNsWxrpPh0a2vveY3wWx1jBgK+HY
c6jDO/X4s5cUMPklXJy/azUUs3u7jhPgDB3q5qawfWtThKi2xIVmQ8v+QxiDmkVgPnQVcIseJyTA
Al3dsMi6H9H/3cGlJ++8WpyhUCa5+J4M+Cg1W5ksBrdBGFyrYnl0RHbdGjc/tQWw3vBtm3YQe2bZ
DfmKO/8aOaXPP+pZKFQzX8W+y1TRCUML+2X6jfwBnGek23ZZrFqQtDqFTWZAnRYRCf3HCqbC5vkK
w+FCVOZCCIto3cTjGFnF56JTpmoyuTsN1B5T88hgPQ3w7mgMPBFkqjtCRa/qxsS1A4yKtMSYHIQV
Hj4aHPEuNLjWdqVqFoO32AfYwdiA+wctUixY9FdgREu7ug/pWZS+fE150ziO+aWEz6OgTq6Inwbw
OG6hNWCl40jmEr1wYbK1HhICkvaCRRiVGL0JosN3SUPvv/eCLYSjmmVWVfDytttT7hPY5yuQAgzg
EEaFF6gTZEKiTSX2oJnXE0v1iK7IxzDyQ50quFHcXSos7mu39Rz3aaKoSgrN5VzQVATzflUF0nKj
ZClxQyAiA7o4I9U8kqsrK/xcJ/hpuTyYSaOz8Sda3ZuSVs4TaXZaPDRce4vIJHH2eLm7l39McDoT
c1HnyFj1FCVQcRtxZ5GuyA+eImpE4aJb+Lpc53WU+u/kA4OGBGrdeUFidJkst4xg+OKwTBIiTLkv
tRl/H0qV818JdwAiveWvZDWbtJdvfzmdgFZpRWK/F1BipGAdTUNzFUfrWAvWMpG2Kf5yav5w0Jlv
ZepgueBDFfR6iJ6QPQ+MpycM7Rz/hcT5Dre4sQdxlNCRYsaTgUw+iKkOQFHSdM28sy/Bw+8bGxhm
U8oAF5+JVBkKvhsMHwkpcaMJZe+bpiBPsf6eXP0rNEHm3RjZobQ+/cy9fq7MBNFc8kUQKuo7MYIs
oVNg5zS1huVsf+1mfXTvrhptKaleSuZqmQ3J1VKJ0Y1VLtTVwhCiq7K3yVmDABVJzSJZA/dD/VjU
RAIwq6OM3rAn4IYuy84VT1DM3C6cwjkPxFTdBmLi2epch9/QaYklxfhGvrWBDbRqjVx5P4g3PwoS
rQ5a3LQM8QF0KfIVSuM06CfshlZ1BGkRbq/N1D5IgYR9xjrlm/hQWiKEI00vLj+f0Guen2p3T7Dn
GpprhkB2QEhGAWMiULUa2Ti0cJfkG2fEgJoNPsLl7ZkDHBsKOkAjyaSuinMtjEzY6hEoFYqKUV34
F1r/g/oMKg2t4He7MZ0zgB3P9DPkzAmD4vmVVdwDgL3JdRZlV2Fn7xx+NbIB68iR7VPBTTtIAhvw
L0PlszpcpayP3vRVU4DjKRYnzbFySnzeBTroipZ8AO1he9AT1JiOe2JGcpkIXeDiCBxz1TCgLZxb
udBEzQHT+k13rP19kCOkcnTF8i+DJPD2tflVdKERnM9HHZmVk4wouGM2VqmRrnybSJ59r9QdlOQ2
aoCZguWpm5WuwJz21CDHDdDdThqiuWtzPWVpklTcdsJfW/LYP4Vqyt/AmJChau8LXjHCMtSjN33J
TeLix9NEaXXvfQ5k7PpRYvnuz1M2ohIcF/1C/UXe7Nz6EpResAHChhvr/j6n5t+LgMF3QKFCeDjc
lLn5hMfjUhzR2q8q7kcpG8rMZUuOR6SRTS2fcAZ1T9bwotPYVFwNllKfRN3iv1EZA8U9QABTJk8m
2ti9DCqjojzxURmaDj0rRm6h7g0t/WIajDworRdCs7LOXDvnq0bywWHvuOXo+TeDiRlR7xmxpdUI
NWsgdFVef6JLj3DwnBz0QXkh6psGNC/8efOQGZF/TUgv0e7XTKeKJJW7n1daEpvrlpu3i7Nc3pou
pgBkpYmKKzKZI4ZGSxDfNXlAs51a7ATHsr7RqyGQh+roeLoycMYRfKbJI+yylk9iFKkIluOGSTqD
akyxemQXwp0QF+pxHvXpOuD3TNEMZC5YauFGw6qwuqll0Z4qAkzFinMG636R95iklfgcnf4WPD5Q
wmunDWHylDJQSFthrwF8225hFWo/2PioSpg6+HStGTh9bz3C9BNQoyr03iL8Y0rAlMOVgicH9Cbq
f0CVa6uVabT6wC3IGjoOMSlXlErcmr6v/9qBa0rNHdMu2pVnpywET5EyygG8w4w2IyOjTTBMIZ5g
Wg2sda5f8EpQW6VpZPGcqtzI/Jl4u5wLtaRz/nX077JmhNEJXZWkXMR+t+1TJt4zyIk1BB5PTX/h
NwNTwv8dOr9cwUIAWjigVYl/muFh+8gSechT2fisJLcDZpgHH3+JvQpm81Civ9zozXF99sfo3wm/
Lywc/QGIs1K2PW72Dc4IwGqB4wAlV7MQgV4p37b2Z6/T8NO0vUezBIVWPGDFkZeJfSTq9dYLg4Wp
ty5SCNyG55tHUrkehw9j3VOeDbPm4foJx5SlAS5NUoohxZ3SPF95NW8rIzp7bJJTxeqcJ3+Tk/Wl
Uh8VFyYObW1iWi5R5M1XHeI8CTFEkeN/RWTPccxrZ00CLPkeZ+Uvg1rBXzM9qRU0NnEe5ceUfjjO
R19RCkgwZ+IM030GPpTeAF+WUqjPlAh/HSw1L6jyzuRjCmRlblyRoU7z6cqp3GyClsaPJzV3CwDq
AwPdk1l7Uqt6ud7sPt7qRKeLFMUO4FMC+tBdhlH/Zpj5oB83sMNmGhO7nVdj8kdJix5E+63QVyJR
eqPQr2loOBtZsA/zsdH1FiZfa/TEfZKlfvmQEvw4PAAozoYKrDgu1/k6GOqEvjfu9Zdxk/FRu2CN
dQmXVQgEZVcBZqGfttfudxLcu4M3tIhNjKTXFmFINX/jOU1/yi3cQjgfWSHOxSInGbLu8higqw3Z
FguTAqVoEKpQHZ/zEm/fkZGcvG4TXM6XHcHUo5anpzr6Nj7z4eZ5aS0ava6TEO53A6ku8fHEK/84
CMN0QHkvCvHu9bQknMXcoB9QWW5NJLVz7cVr8OxmvQ/za8Al+UGoN0+B+zSp2TvZzUwMWAjYvS9b
yko5XEGO8kmK14bttut1e6lhOpL1cyd6HtV/KlVuOyUwGQ/sRN2/6SPrQAxw8jqzliTFJSOQu996
DOAGkS4813g78yKYwgpzswRT+terI3CnRdsgGBwP9DBWD5QA33SZitrRX8CGv8ZVzAN+JiTkp0KD
3uvFScIfD0z9B6rvnUkIXoSQbmVy9L7NlBkfcDIcNTmUNd03g9U52NsOkY65jyj8RXy1TxKiAP8p
ZXgoEgSrkYy7HSt8bjX+gknp8CRgQPYiHo8on6QjSa9TtlnEsOTMOpbvY2gTHcjowpgTT1hqJOqH
mUj3CJd7LQQF1uMNLIEo6wsZh5OtCNJNg4FgLSFRqJ5vW4TgpPn9Ks0iYTCI3CInJ+DTWcUrWGz6
PrNQlReGXvORPpMYV6vKlITg5oYRiGYiARoBbeBTB+CAQGNBoO8RkkGFLWGfORbwy7ATN6sxEMYj
RNHGE3PZwddJVtZUXXAwHeYhGO9QsHwvdaEQJOY57ZhzALBY+ebQ2Uk9w6mkpRlGSuzeCVZUrjtQ
4YDG1nWDhXKhnZf+j57Bp1Nicj//J4ug+hUl0ZFtg9z3gt0y2rSgqyn6avg6uRZnFw1yqh6knjmB
eZqnE4vVf7iqUCDvP+DqKrumzDdZaIakrixYAw+tQXuhWHuorokbNoa7RBvJGm8tFQrtypeDRDWp
4F43W1I5n61lVG1Gtptqpp+L746xieCH3bl342DcyCCHMr+em68zdFb67IOtu3mTfthLUUTIyUDb
ot9YzDQ4dxZJBS+kzKytSmR30U/K4hpfLxH6dPWZxo5CUkpMtwrZDV5rlahvreMW1U4IzQUxps67
wr+I7Sx+PJ3w8qN6wYpkNvl0nfle3G9XJLHE5wSQP9yUMpME30YmrcD1c4VTERHPD5np4r+/V/GE
td2tMNhqa3UT8wAhMDh51TWsG0bmjDkKM9/LGl3UJjp17T1mQj6dJh+kSdkQkGkaohOgwxJtfbuR
hAV+6DzCSjBnMfn/wKXL13XvWN2LznnHuSBaUG3KRbrarFXPm1b84KBTSNXrnWC7MQW8ySzFwX9R
VUejR08XP7R1kPznWpj91NUGgOBv9lNmpP+oS5QgkJOBCczh6kXG/d5siUxeSMURvgn4x+cG6S7R
V0MTuRKn8rnhAw7PMK3FthbfpTFn7thlHV74BAUaNQmPay0P+GWsM3fTvkU4qxy4WM6gJsYXXfEW
biIA5fL8YwO2E2wptJoOZwx5/2RRTUn5DNJj4+vKB9tg2gL94uMFdC3frNVdl9TXU3Lu3MX6+Aem
+J/nuOUsO3uFfWqMK/sHnuV/8/JMJYFkwrWB786FuNW8sx3OMbd18Lt81eoC2Efw9lBQHhqGSn+y
Suu7BbZIHCOL6FF6Mntrip7mxo2hXrdqAdJUce9mV2PszAtHxczPbChGSCt2oWlfgWcIexBcgP5S
5SYsweel+WJnGhrMwGeFSb7np0cnT7SOnqhYHAqyiRxc9agbfiJ8/nyMNqb7S+f3w+wHbCRlTDtc
Uwx87NK6cijLl376KvkJ6dmpA6aE1CkX2weqXvSIG+29RPlSmItNsJ4UcS0WKWjLAGh7AFtV+r1p
drJieRrF0XHyDEb1MwlDjj7HF9ARvFEwrwUbivLvjn+8ss2lmVj9zlHCJw4fZJQC95nIlh6QXe+T
osy6AQwGLnBpSN5NGZ1XNN8SY1JEfR84anpZIH8WvDqqeYEjHG7AAXooM3e8D/o4JQhQdNuUPVPJ
/KUtS2rrx1DfeaNGWJfGG7E1DuQ5LJYLMwYtLNqKun/ZE7NXUD6AikEdYCQdh8J5yMBnql5jsTAH
+FBYchNkaThILwOuhc+a++B2WzJuIQLtNmay3k0Dv7hJPDCKOs7jEJEZlgF7OCT7mFUYn4wCWCXp
IqRGO07rTAfXco+4sKbZkgIBbybT+/E17I2Tpq6b//3vSiCKq3aLN0UJBMZ9RdZpC58xDxMNbhdg
aMtqZ7C6WgtnveOX6HrbYREbr8IJ80zWEyGbqjKgrPsckd1IsRm5b7tjdT8ZRLFTfuxcCQSST1KQ
vxgNXxTcs4vKb+RwPjTgtawJOd6HmEW/owU1Vswnic1mbpCXdT26jQHHi95bYv8u+4i+8Z75M+1/
3gI4DSsIyuEgxDGH5Q34G+TqCt06B9AJ5XgjJl4NO/532C5Z8I5sE65y9Vuq1aEtMKTwqhqjgjzo
okEQ7zsuPOR4RYNQGbBALoLJRQhjZujXxRbT84eecM3mRTg9/kbFAPNI1uqeRQPpyomZGlnf6BgO
jr/o831/PA8FmVAK+B8XdN8nOs2neOstMgnw9x38bo3cwmopyHPE2/98mW+nHD8MFk3KaxGaKMIo
RlQeW7QlIdjvrfE8yzfb+wWIbwEenQBJ+T1l8pCP0nY4/14H73qkGFoU3w2/Icrl6+2AB5m54k5x
TWwUii06U8pXZ9qtTbmNyNK6NiTDHfy9kNL8YJaWiR34ummw879EF3oY9uQv+vz722knx/Z/rL7J
hER8mA2RpGJ7tcuMNolCaluXVLokTBymoVtmRiWvi3MLNKBqs5bY/IH6G5hQJSUJdTeMZpPZqQah
4q1tdb1a13E2I6UoURr1oYPfD53WpQpQsnZGgIY9+DctmHgWftaRy7duuiDl1zK2RG1x2b4QzFQz
b3GILiTC9ItoOx9aWeFgriFwGReNxfpu8Xa7ymfr55StDZEFleJXHvBq9ctOXQuP9OI5zwkEzVPD
XAqGgiPS+BCxlVEnaa88ckW492kI/wwaIk+SbkDNT+Ijk1a8LP6k5HIkyv7Xieheb0TksLcf53Db
EziKXG/z0mqICxj9Rk+5PeWs8Kg9W61dOvCz5LHN/4RqXOIhb8xOgOGHL4f+d/AYLmIVzWL2oVAa
lB5XZFZzr5q8p9KjLW/2lKcGDPntXMo9k+oOv8jujeGiW9v6DD9iZsFfB0a3/5csSvnlv7cVoIeO
7P4rTGrLUh5sUb7Kim9byTxSwWA1j9lNb7/PHIfhh+DobuEhSd/0VkDUrs3J0uPxGk21qNI8G1Qz
4MZQEi2JB/XERUXBxf/GIX18Rqgr+Z+zr4ul7xvIgoVnaEvMCLqxayKOt+GJF4IgO7fY6CBFTnTr
bUyIh6XFoaZq33+UX1kUnClNGXmx7NSVxnX1wf7cQIvxTWD826aS3ZAOf43/VH1r+4KmLo9060HC
f8DltnGf5kTJZ4oAz+y7tX3PC/9ertbvlVigDFwSsgoqDb/OvLY2DBAFs7D4kZOvEzPm5XHzKyw9
pI4olUt8QwHgvr2RZuvJbDynaL3pnTN5keuvpmFZBvdOaM8R14Y8dz7XGHGz4WofXtCFqSkWoJ8G
wYZzZLkM0rgalsYewX+MHWApeU+G6VLXvyQ6TTD8OddwlEdSPxvRtKO/E0y582z6XH38YZzTdg6M
Fp/ngQwB9dAmqPhWMgxLDR7LPTwXpSCOb5FEruHJRMZt9emSfgorzBg7FSNRmjev1FcqlvwjxFUI
crkwGpZdCy5ID4CuZG8jSbCyTDMUZGuUiYa4LIqyvWC/tlXwak4oGG0WEcSKZEjj9sJKI8UaqMk+
bC8BdT52jYw1qpYejzxbNI/vGDorl+Ppz4HrBcewptwvV6M2kOehTTt1CQ8MfOeHS9YnOIG8Gf5I
Nq+q0ay1AhVQSBetYl/JW/DSwCJajVl8o9sdn4+iZcLX362aZyBSZfoZvkZdksGDcDKCI35lutVV
2WEoYxjzeUiyezWt6BihL8c6gi1N9fVnPSpQBNNu2yrbufYFnfF/i+Qwtc1NlYW0XkOWgcxQrwJz
tZGGr61LBYt1hcMpFp9Ps8RHmgemE5+nDCkMiKnA9N20HchQf2UIhmRN2VagZzjqKKa5iFFrrxAx
FhhW60TeQ2v38bkXjXaHvZ8wmwCL2AKUBFkBKM1aMP5FuhxgSZvMbJht3iQmBfB2e491cTts0M8d
Ixbpzy9f8q129hXC1UyY+Lj0FV8feGXHs+P/I2kr77WVIJLjcBGD/PcUi1Y8WHStvx5ZpSF+z4LW
GQM6egvSjSPY4opL60oH8Jss05HfK9vFD9cpmNnslQeXuDsT/S1bu+w5WutLCVuAYf9OwGJwRn0+
P4SleM488zzJp407zVIM+4P1M1G5atVsb+pLp3dMGdhiELY/skiso7VPU2xsJ6cTVNi9kBiyYUry
2S03uo5/L/N4UYp/sqlJaV4w9C6JibIPB9/AChEweQ6TcLu8ZCyxyfQbcWx+Ioc31vUh/MZFSPt/
gnLe+JzNDr/IyObzsyW/JfkVPgisf6AVlhft4v8IRojlX8regolsYCUYps2Lj7G88aPu6wmYB/k6
EedsqCGsyqrjW2RpBewm4/z5YMQYE/m66xu03jjqJJop4NLjxpIFH3hMmBDRWfgByUu2FsQRJsX7
dRj3RlNB0fl0H/U+yx/SUZoO/YIzcbTrVShfgA3p1lLcgsSymjbg7faa92g/09xVJ86/GSQTtVe0
gSwKCfz+xughVgd+x9lO13kVMBWkxXSVBg4S9znT1GfXwlbBlmR75Jdd/2VOsZeu8OYBMflcWrP3
M3IUewYMM5cxjhgalf238QnVrBoRma1XlwJ3RkhIRMbCf4IdjPP+IU2mbsZ7twDkxB4bkZUICrZ2
OErC8KicHLbY5uGpSTAcK9bq0vzpk+DLjg1+E8CruQoTRMmN/Ekm24CKERwDk6PQYQk0T0Tj/x60
Dz1Jj0gWajjuRxeDr8NhYfTqjgRIv4YKCJpwJHHHzbwe4A6tqkS6beEmO6vbXNIXqiEGYWQ8AKYQ
/qbA2aJP6OyM6omVkFlBnhaX+rGTgTc5/sTxFm+rvlpLe5ND+dlY4mZ7LgInSBNtIUTJIsjPCjb8
uZue4BqiahhsWq6alr7ShPlOFf9PhNY4ZOnxxa/5ON2xM4igOt3FgfPxTU4s0uuFZIEnN/fK1lke
MEsFWyVzzpNmCrlQqdv/9vVu5d2uig7DQqpIxomwsroqT1XTtOd6ACkp8lHFYCoZS+o3FdvdJN6z
Hm9FFSrcFTsAnwTntpjm7mXOH4U7Seelw4BEjUheIXcfGL/mPUOey7peA0CW5FHtdN+gxI2S2sjC
zMjomI/wh5t/nEmhhO1rzx9zO6+wXgtlqWo5CfxdQN0ESSdl/0iN7/bK80NbKXUScLg0YMjM3jSz
HYXCGignBYbewd+DUY7HKE/tomXp5Tutjk/cWuYYvotAXagwiIP9gZotq6gUA4h6zsBxD3e8vmf4
3opfX2vaVhHIUOIxLnYWsbQVPYKJf9yyjStMy72ZFFS7heC5tj1Xnuj4OdpFS3uF5JPL+SLgXwlX
cXi9ZynKIr/HhbkzIcLArXcMG37VtxcWcL52jBY119aWVxC5Rcle8agohsF3KkWMy7qvA0Z+f0IC
ADUWLzQhAbIpRBUdPbFShE4xZWIHxuB5l03kBqv+RTrTbYqT6iOKtf8A3l28AyO9E2DEAuiEtm2Z
M/lDP3q1WUef8wYpl4G4a5kRXt+EPEWtQ1q8+9tx1EtgJ/d2VozUV0EGXOr/e7nET7Qw0ZRspRnT
9QkyeWRXn75MH2eydNVMxgQwJdllf1nc8BBLnDf7KMfbe187NhkJ92TEk7VUfkZavJ2BEhez4Aa7
bA/an8a6Tl09hM5SH1M6kRiXG/kDVr89g/tPaigrTnXX7UPTmSPaZsooFoHgXQwSrlupD9yp7YTM
uEltujwY0m7wkgGShjsveagNzXLBsHlHsPfzHUz76QMEawQz/TXxaWSKEAch4yxywRusUVbRsd1g
5OFruMhm0pLcxeriMzTcd03q57kR3FRqyq4K+nomaou2pf6E2/oQyC8bDfiMoVZgJ2MUu4pA0FZ1
DsNC6ucg/4PrVFsalU2Ac42f+D2i3I4bUVLOgmewCMIWkr02ov9ogeZaqhMkSzcbHTkSJCjO5/Sd
xhQhVoMoMxT1IXdYY5gq04RsbPL2ibUHn8RrJZrW2ZJKXL6MGGtA2a4gR+085DypJ3+anM2JWayp
ZkzAYQgWLaISel8GB+CjY1eHcwgQNrxRzRy5XzasEdHC82mFHhpUrUiYVKxS7ROFmE9vByks8ul4
N+C8q3q/xGEPUYMEGOXr/tmHLgRx0Avkfn4EsVM9GVRdh0KYntW20Voin5q5L6Vm6fmbBEHBPLcb
ZCFRV5OfOE6IpPel73eIvwqFXD/HHl7hEuqE7Nzbgx58M2MWlExuK2wXHWOfVk5fqKLWII15QQx1
u3XAfeXackcTL57vMgsFGyzXhHuu5/fjgQLQJFhYkOfn7+zQQJm6xfWI/UFS+Z4PQLZnjCARnDMW
rieECg/jQj4XF4XdvA6dsOjUZ3zbH0OQtc+GUFe5V3TGk6sOYMZGuDaTdrYT9uqRH7reNRqvb69o
y/H+IFJGf8wnYbcfj6NXAoV6o8fQk/brorkZHnuuMmKHkxbaG3n8ccrSyPwDiNLNtD7cwtJGO86o
fjabb9pGpFht0rKLhtA0fsPWlhljC2J2b/CfWGnyfTz1mPFANkjbxvo1SSgzEa2l41UkcZPzvoS2
+qiz7Cy2hCplT1YUZ181RUSEq84AmHYuZIivylnrHDbp2vQpNa4XVpwDOTHjjCCfll/ciRdAc2dR
kfeBAebP4yLSSlToM4blM9IpGxoYqeWj7Q+xvgEi2xTdMJG0jCmPi3dL7mDU8avCiR8hhX22jSBM
0IF5iKAMgcdgi3d+Oq1BEgyQW4rvz5Ug0yUqYnE6rErnTEmEr3wRWJSJxgQHhj66X8cWTl9p4wu7
+si/VbeFHVZmwOrwJ5mM35V9J34Cs3rO9Ur10RYFpA9XgQAF1oztQDPnrjXblZ9b3iYcQ31ceAE0
puiBFbVVZPlYv1UPNyp2jQVuASCm1VA4FjyzaXFb7W1VQbERZkImoP4RYLC4dGPRP3ytcpqQCZ/J
lezC2jOFBZDZWZSezJmyLkkWYdtsawCYZJKN8MQuUxaOr+Ldgcpip83CpA09/pVHuiRRNv5YXG/Y
RbEmdYP0Uxy3EFk7YdkLYOJZq5V4Higbokhr5a6gfaSrS8fIXK8NLjTiXoLTKsyonkYkrlEzieLC
vZh+3f0gJM4dA1s5mmpy91sCa/mZ+qQCuZzNljvnsMs/M+GyCS1wCILCBiYfznnnX8QZ1wO2yVmU
4AC5bssgPwEyDbuzrhew3jDpuVWP3ra7U08o9H1qF9BXoIRrYsC3Ht9nverf6IRej/aUAuYKruWD
RPZWc/dUE8AW2/GA/3KCMSPNlrcWi7P13ANfRZUC1mEPvhibxKyuHCCkwbuJ8WVLG5+O9lrbmgH+
IGCx1/svxP/6vKBw+PFfCbRi3QEzKY3M10Pit+vnqL2s6mKdPL+wbmN4UypH0zLq9oYdy9VhiNtl
okNuIfjakfcfXY6Ln/BVSMS6YhOeODnR6pucEo3VZFjzKl3ZXv2mpMqrj5vGwxsu6/P/1gwTr+LP
IrjIibnLXqaRUmc6QuhYgLO7QnQxgsqXm3+DYnGmhC8XSLdzqxZkMsGeqYWxPPEaLeYmIFnEkPYU
xPeF7FAOGXVziy6f6BPcFc8MOKuWQ8zFeNSS0ZbvZr8wiVtX4uDxX3xSO6aPD7+JLa2svJJ89EqF
Td7xyF7orejfj55walomdK+/iiKxbl631AwOzhGWhALKHHB9OJWKHLKUyMtbXdODaLawj5VqiY5V
HuCrdVXM1Z6l6zQfheBRQajtzlUfFS1ud4cxgq7G4SbH8rTDeW3S7Xg1RP7B1Y1DRIuyVzvlvqJ/
x5mvL3t58VauP/yHZ9wRa3NWftA/cEbAJACPwKvyFiDKRsSG9ikmfIx0l6hIql9nkbD/9hdKq31E
5fVZNdaqCBlGOuSoHWjPTpGP9o8ELJJZ/BB8itk/MNCJi4LA+FL3khHYqsVnWJpW5EUiOYnYHIU3
QkXWXnkT8HW7kr5o4WZzPDGEVuF5dNCwWejSKrwaihBDmzTy8u6yEM9Qmm0vK7xIHUrrSRDLI3V1
fPWP5OqkJn+J6hEDVKKyHmea7vfHcYUtjIsiJ97LzOo/XmcJmJb7VV5TywbRKr+4Y3EwQF3965Rp
kRQmv3MyN6+0ok5rUySM6kOJjbYCizyc8t/t6bfVXV4dpZ2mtemQnXmlrKjylD5lim1szEf1buIT
KB8jR1o1WaE+WWOW6AjSxJfc+BcM65MOScO9pXlWVNuhr66lqGtx6l4nfyFlW5t8tfUH7Vw+mwwK
TtEXupTIM0WOXHhh50FaxB9bAaDOn7Gvs6eUtmjb4zjiyKoKrmfw0jT1NtHwNzkqrKaj26CZmel1
tI3eJ9spdfgtm4Qg7J9RK+M98u4b7YC0KuzqF76iz1+WzDfh8BTWGBs3XVudwytMiXcyvya4qtMs
2/k76CrKvSEflqgiMtPWwCiLiE9FextgQuG1XNiqVViKel2wqDhtJ0KGilSYbDZCfmqbMiGBK776
yw9x4tUerJwT2MFe7J7Ye0FjLQoxCkAhWaALA9/rAO9ZUfKRtwz+MLaq0c9Pwlu6VLSIH2RtT87G
uOrC0wSxqUDE31nBrb5JWIKnVHpyAnEQ9ET3h7zFNvXs+7kWrGP5A9msM+aW8A5d64spyrPM/Yq+
+zajSNHr5i+2H5Sd+DfVjPFXoyLwNe5zDNKFdHNcaYavurEGr8hxiYowTE+aBkttco67UsM2ig/x
6PT+4SFW64y86AMQ/n1i1ICn6+9IVm7kRVELoFs99PHOsf9p44UPZRx+x8q+GzGntrzBxCwu9cib
hkJ4BnCpKLciaWVm/jZ4qMC2Z2DuGoErmtF/Rgyprg4wF+AOWikY3ykWY8qeUs7h6W5BMfGNG+3U
JRlVrjhXbwrxb3Sb0aqM7HfhVpcEHwCxWov9t248YQFVLCAficz4hX0OW+lJlso02qIxpYsh7vu5
RMjvDeBGoSnpTz9Fjubf1P1W9gg62bSY0Auegc1EgTqKIT5W+IP8ULE0wYT4RE7GzqJXwzb1Rx97
/ajjeF+2I/+Yfm/ifegsLDrS0HVA26PKledvyQAM4Gg/8iiQl2WzO/wr/8r3GqXavIi5m3sxPXJ0
zrQrjecbJOOvDoWyuT+GlorRGG7bZ/3G0Ct1K8gjyNGomQZ+XCp8SjMlG3VQhMhm9GrJl/oI/3Y4
9Qx27Ah9mP3iHpfOPLtg0v5GFHI9LVohsILp2rUG1QCw26ojekkO0pBG17F6Cee150KXi5WlYTxh
HVA1VRzmM7gzYN/4tKAe+KC8BCn278En5nMvqKeTyUjAydsCf1XdUazfoz/3s1FYbzEVpxzqu8lg
iNSDzXa5bIzEUeVD48MByrhgveHvcAKM/f7kwvNN50djKaZprHgprKa0u/oYTcyZ0P3Plzoic+dA
jbiNNcH5kZXYNlHhlGedqEhxcsrYG2ueuTOOM/5jJLuBRTRdJcfLHGwg5Xq8D/Vu8PRdvlF43bDJ
dAj5QYjI1uWmvdcvuCNZ3hdf6ELz0vy0t8xMZryq3jnQrtzU2CX2aUrL34TisYRIsrWLGIYE/eUh
+V5PLV6rK7jbRvHhRjRgNtEhvvnPgSh/kVYs9L8wrkRH0UrW12Y9+aibGMW04AW0ZG09EIk0IrA6
6V0ialzXF0GPd9a10V9iMAW9pX9ZCJ+zTiNUClE82AU7CtFQu6sJxP/rwsGXXGkX9UqWk0cJiONt
2cO83bZOYyZ4ss5s1k5pKCL+LUCCOty8WghvBJSAu3BhNRQH/b1T2bfleJwmGyM/wFMpDLKSCvr1
9e9ATKEY+x/YRSgpWX8ZucFuK+mhxQ9297YwCNASBgvvzOAA4CrpWiD+ehk3onAa/LscHIYmsMg4
LQHMqwTkMQzhMAqxHurxqfDLMNQLS+MlIoCSM7FH25U8W1HwUKcFwEvYqPgs2Q0T7YaNWDdMrWaB
vfzZ70RB9bHHJ5EwreQBch8IzSn2QocrVaeVs7Y/YJC20EthDhF6mQ+SE8FXkoC5QyeOj8L0WXzR
29t5lK7PbZH5h0xUXavstb1hioHXu/F5p9T+vDqqEi3ydbqI3OWbuBS9iPUk7DJIvL6/NdYKhJ4t
xtHzuOUF1Da8izBXOYaX2g3nYse1sv0jwallzCRrTraLcW3eYO+ZtypuUOFwIVyKwhBcO/89DOAA
QFWBWjy9F9thPtmbwDGtUANhw1sF6wNm9sJpMyA7Y7NlNxx+W46D7n8PpBRumhzBwprctLwFQjng
nmVmdXp/K8HVHFdfRKi8fTvmWYEG5vuosIywYqWTCG3tTgla3iaJ1m0r9DczwuxrbFrSTAUH07ag
h4buUMpm3EEmb7yXs1fjhqOQN8t7HH3IpkNyiNYYE0O5atODwgKmhPOE0pKRav2Kchj2LDi7Je+G
9Zlt+5hDDZuNch28KZ1ViFhh5ywnJT0lXrfSBW4AiOy/Q14CvNot8ZV9imwB0ZfqAuM49/qQ8d9l
KsIwfXJapak7maOgykOFGV58qNufXkoyy2TLi9tzWv/ffZf8Ne5vt1diPiTSbHOIkq3Km06juzLX
Gx41weMwaubPBcb9PNlJ09CcLElchL3SEOIMupRSVASRxWoqVZ8Zyd6zjoCyRhbQc48PlPA3i9GI
Uj/qFVHV4s8EKQja9vG4kMtFOV1ZyWdJW2fCHyJnlOErTr8UhrDkTRFEpG3vwEhsQYMfdWPd7zPQ
7Ra36ktAWg22iKpgGh20lrObSpyEta+yPyfdYhUdYav5TIUa+TArf3Ncl6TuCCwMy8sYnprZOck4
cBfpovFwFBLKzfiS/0/G0vh8BzsdB7JWtaWKelWbNgSp0X/UBZIn9nWS8ta+cJiQvXzA07b3AT00
XrEAQu8jIWCZRrl6+e6A7uHVlQ0AdwMU9bxPD90dXm0MUjky9RUahEoUwR9rfpEpkINnKX5Q2V+h
psH5Ef2zz1DzdQFtQ6cvfR83LPcY4XAWSVMHGjhw/OBVoiTuCdUZ4Wn5c4gecdlDCy8YXnx78j5n
aygutjhR+Jw9D2Zks9J2wH88sNDQRnLDyM4u4GoHE+70i7MScJgiXcvw75FXKolm4CHNdiU1jcBF
b1YgWH84xBz/I8IF8IJYaUyNhSSOkBXZOWxGDO78meIMuXwn9ldiHIybpQpSk7eBXrnbj8yRdtJX
kIgSOBzQws1f3lu1Os3nlWgpwZfhsKYsXMKfbC1Ev+YyOq9kIvEvVC4anTPVdtYvxX5X83UOxOcm
p+2tDsXbMAGLvkGz1WBqHt+L1K/n/oQjDazzNzR+gpCi8NG7p7MNpn/43G8QbLGTIbV+vmy76Kvv
Gwyli/Ex1iWd0C6O1LD1Og2N9H7s4hmGM01O1V8GozNcG3aJ95Kiclm3JUm2KgvCjdNl/iPNc/S0
b5A2EpkSIsnBsfACkLYbtUrzDs8nf9SNgcYE6jusTXsmRCdebatJ3Y5R4lMp9G5GRWS7Y7OIsRtl
iV67TSiN+Ch55dhl6IFjtJ4exmS2fF9KRJK5aaQ2/BU6P/df1Rb/LsvjNQjB4X3hMuvpLeZVlGaY
nCwgFzdXwQ3l6w4mx5kdUxUY/Fg5IuE2Wt5W9jIwU7QxA5EDJVZcWyWos5Q6n/Kbcfhe+n6Yr9cE
hSl6aLXL8Keva7S4MbGctlf7ZH4sRRhDfcO5TtKeln4MT5F/QugAeZ2OJ2Xjvtp7lKAH3U8FmEgn
AK2rjMX5RYW/B25vcRUy0zloOAUi0kG1i5IqY25FebpmaG4JP/NnAnXgnE6x2WWxeHAnLKXQDu8m
u+eAN/laRwcKr/oelO1NLk+VJc5HdknQZdgMdKAKJrhk4jNjzb8nPWSA3Kg+Xz5T5iXSYlnzjTdE
vM1Zn0LZpHPezh4VYbXDWUpUxYKj1uYKMMCQroZYIs6YNXdraEFpB0xgpRZMYeP3yq5pbcPGNcbi
vpr674KjlHJaRhxEmOEoKJHqJOdFiWaCf+lk4G1BT8rrIWZhtOCjWZPLAm3IWBqzrzD4OMW+9slJ
Q6Bgn3ELQJRMWpd+uVbN5KlZK8G3Xzt2ulkQy0e6NYlvUs6v5emKsqPqfw5DsOEy+ed438rep3sT
7LOoahy3RrGBiFoUaP2B2WceVIhy0u5n5RWxyyybI6X4jfgn+1HC4jvOBSb6GlDaithdRWX/sRrz
dAObW6gwrJyqL+R/bDlL1X6bqQ7meerbf0VYUpZBAdWWhwLn2o64mFPiZY+//ogRv4oCWRWFVtnu
5sJf4MohLHkbG3I66BaqbOA6lsW3ACaiVaqFEU0gomik1Sd1WG2gA4gs67VMQsKghrQqbSEUORM0
LUiNcMyswN9yX6npo6tuvubM8cz9nevf6b+Q8dG+bS4wenf0QUUZPw6tfoWPjYOEHIdrxRJacLq8
mVmsAJrbFIL/O/ScNNJq38IwooiA8i5gYlVvZw69I+1wFNPyo9FYNjTvSRBo+fPPNcJ5X47URh7H
I27AiMjUS4R75pssoMiP3Rtap/rYQykn5bBD+VgYTSwbBOzPWPAYr7eVk1r/wMXGxAMF2XdWCzR2
YwZvjREU8FnEdEapp+FJlPN/epHrDc+okz3FUwPXf48ijKjzdHszYbcN3lLH4Lx+n1x+Y84CZ/JK
Jh+XFuTNStLUMxLaXJ/vzJAFadpI9ecxm5QxRmCkQXFugjKLQ/DI/P6ShWS0d5PR/qpuz7iVKtgW
VKqakTLhatStR7eM/ihGsqqfWbkCbIWYurlEY8gjrhePQS0TRPvhaXs0eslny2fROAdArC+t5lqu
u/R34yS9N5FzjcZ29yeVQNmqhzCTpA4D5mRTDgqsJ3awNXBDlFtQAzF3LQEvJ/TzT1wnbntbstRp
UyTHqOzgpyDVmd2Gv1HMKkRtIjMaFzuVd8LLZ5HMOtbjxyG4FJvux+KuS7pZ/OZWaADhcvClOGnX
R+t+Z8JrFrPVPN0Ztztv6EV3jenkWeVmB92TKAaevcnXvSY+THs1V/q4cM/wA3l0oSEP5OW1CiqM
obtpgibincKSPLYw0JPZJUie8Fr6zh13zz0+U/gY1IcWQvT8fMsgQRQveNHcf+KqzKKEJXun89xQ
7oA0Riua9tMMe8CHSkaRWdGR3jQAfufwDDRmH5iReUV7F2jlyHRjyrkOGD5FAfr00g1SguH6506L
YiS0rDyXSFYwoHtrjjYB4+xuWvkqCXNelJcgtfeAlRJ+44luaa5zhXc4XNz1cnIyeJ2nLvXPka8d
f0yeyvxa6OBFsA7qHFdi2PLLc68k3RNGbcXOShU1DnGP4sjYZFoazg0J29N2sjWX6gV5tQ6bF2+b
H2+0fTtbAQOqyxsYpeWhkGtSQ8qqH/EVaWHRqsoXF1HYZQvRAxTMGt7Vu7GY8QrBkD/rAUUlxCS/
Y7Yt4dfZztcAOV3a0f3O/pX9orm0QEFHabm1a6Wwkt4C4rT3F0Td7WiaAEi4LnORbL86DgDXJB4D
ghXCNXXCehcoVVMx8lqRvHpJaTSA9Fu2Ta71dz83P0AyEGaLn5Shp9W0eJtGwRbMX+nYMpDn2i2X
vBHjNz1G9NNXEFqd0iasAoNOeOnigNyhw27K/T5/mpt3ibyCIpK4lNEVuvgrxv6Z6SmIRCH0oh9t
Js8XuykDGSWibLkLhqC2NVVQoDmQSCTy/9cNcQLLo7/W0TCyrGqPgccPo5iSe9khae8W7aN25/V2
uHrCGF69XHk4EbY8BqKri7bDgPEDeZUAML2VJoiEqUoa4aNz0jIl/lFgekM1jIRua0O54aymRqnI
X/9Nvz3TDk9t3ZYnshhJVAt4o9a+FH2YJRK9xqgYA91tlpX6/vuIgXJOC8cdXqGE9qKkgGYXS1Jw
8XB4Ba7MANMm01DRPXF93qe8h+MMMwhle6oYrX8B6iOjUkn/0ZzwwXtkeGHn1OEG0tMyCNP6vaFM
8hrxoOGgxX6WLOBakmb9lyYH8XESyw2webr93OUMWJgZn4GiEdnqBK3FDqTIh26ONZJvjq7QwOz8
cjwPz/9fPE9Zi14zBdNCAuYF9UAubKIs1ExzqzAkkYQWyoaVPxpblfT883PZDOUD4pSEeLdcQCKf
ls3s4pqP/v03BQ4uPuF7pOem58ah2YAgCTdFXP2qsnpjmQct7QBAzo7rk0Otn+UUV0WrctAUALLB
mpkYeWiu43DU0uL0hZbtmRtHYRE7XjOIl+v+LegTZgEG2m2sf4g0O0oiM4Dnj0+YWmXWEs1yt3yT
6rcNKua5jzMnMfkmRIQ9lDmdIAcMMzo7pQxTYvMS+Z3dQ9xCBQVflfdPg/lHfM0DSeTgquSwrjW6
pU6K6ERlDrn0G7hGsbneFAdbOPk3hYGsxUl9ML4h3Vcicl4RqVz8m+GS3jAK2SDSPVT9Nlw40DwY
RQR8Ms+6l7lPpOS3JJhh26KY3fPSwGD7IlcsRO6oa4Ijtze8BzFg6FAXuXIEvbQqQ+B6dXdmRhq/
B5AjiEGU5koQ9bnu7FLi6ndqFksBApFFihIk4vLnjKq30Kpf80cJcypxU+qtsq/dQu2bG6U/Raht
DZJ1HWk6GCgkjHjgfxHamvBsKpMCX4vZfmPw3BPJ0fkFBzOs/CeLv6f6DztyASVlJlAAh7B/N4Kl
hiqcBgsnrUq4zfIbO/1FQyvtZ7JRayOL7K9sjNvDHGcn2kPBMCLPjoYFlTap+SL9I+CTQQeCYOHQ
Xs+S9+ueJKHTDYpyxhWfV5fveTg0z1KE20usE8H1FdotTmkT2yFn/D9bfm4WGdRCnewF45iSKM6e
SPGL07r9uWG9Tpv8Sn0+qLMqNM3fWdEOOXnVbl04APHXJHc7V30c3rVyJkS6DDvElOPsxh/FOrup
/MI4wyyN/tA950d+Y/zgSTWCh3Y4cywTgGlwEEg+QMnZFmGFcy9wAjVKMkn8LW8ykYx5E/6Pe3nQ
6spuexvReqAPl+qWVgTJs36RlxxTVx4j7xgWxvl6i4h+gzwltWAX6wZe+VwkYjgOP6uq6zNG0PMP
K9DBHgtFi+MW6GXUE6GWjkgjNdu+pnZDDNh/JNAqBLgvQUDAyxsIlJzdWYLcuqa+lbIaUgRRyk8I
9v2D3Wb8wKfKbZalj4ux2IU+Gx5zNPKI1rArOwLXLOZrbd5/IPUu5s24gIxw2pwexe9vbMS7jYPR
A9Kupt8Y7wlDD4w/AekJIwH53wE72hbW95ZBzwW+WoaJMUb9sF8Vj4bjhqYMauct/2gaoTsdDYHp
6KyXUWhvU1mi52KDKCT1z4gd/hXKn8VXdQaLiI7kmy54UNgF85tFvLlbnCJEBNAvEZi7HnzG2cgC
NJtsu+jzaKpK5W5mL0Q0UsOoqqQqLFEMERs2NUzhpOsnJa3K9ERJYbxaX+CpODFF/Jz/iDsqNAR6
0LR8ul/GEcDYu6Tu9LZdGQyxbXLC1llGmqTsGyGhtMnH4zMyQn8UEKwSHyrFR1iu4UkoH8Fj+T+W
mk8Kuo5ZrVUJ1X/1jcs4Fsq6oqSq1jyPJdnJ7daPy79Xug8p4N6KHBPzp1h3bCrGyC5/5naDsZ25
gQ49s/DyfsjQZmQ/WyKQKs31SzJshafeSl/kvjXy1fKZRhlvRWzhwIBcM9jrC7KM4HEJSxrSsR0T
KUqWuP0fQa4Xn5W3q/HHaDtJC+6SHQomuwusV+tO3Y4ov8CaqGoKDqMcJXgOAOYjXtqfdq0ltwij
Y18pTCRdXSqwGaN8L/ovJ0qlBjFhDlvX6+Kd5oOwgyxB3ME9ix/KpRXFOr1pWj2gasm+DKQu+9fQ
MjDx3oswi0CTXxgWHTr7fzEDktBYBfeNv01gDfkGCuoMSVtVGnSJu/xPM5Yyid/10YIh6UqXNuIB
px1wOYDO9VGsWeCA6jpL8Wq/vdh7PaKK+gbniSVVk0yopzI7axcsn2Mkroi/7zTHWpxGuNu1wbzk
S4+OvQ0TrghrFfF8sAZYNO0o8WnkZ3KZlIyR8jux5mBv+cVhyXrOeGS/7xkp02REqcKTdjCDDy1Q
nCW+cJEW7dgwQdc5fB3ZSGZnwBP3yYiax5t3zAY43iGtIFo+090zK+goqKjj+0cUu86ZjP9nj3Q6
aeNcrNZwlOJ4995YhYLf08AD+BfjIDMROHLpZS87ZqnIHzCpNK4v+USYAhxMTiapcXFToRXEohcy
cElRrSd7LblqIwPkUl6ADF9U/0uDIF4gMK05PFjZ4Ib4xHxxKTTDtPmgqN09l5bQUkt0/GzXhiFr
LZEjpO5ZySwieVQr+R4Fho12KQv1f+7JtvC3oBiXW8NvjmilSqxwDsmnlGnnYltFxLRx7mq43lE9
4jjjGoLEtj/VLYbIXVO00lFu7fVU7Ri3R2Aj3IzDUJei4L3I4T5X8pEg3/TacqW2p+eO9U/aZ/NP
AJ0eHOwQCI+rVO5sKbOlfj9uYpspxe/Y2WZg22TrLlW1aQQs4Adwod6irlk2eAEm6tjlfhcH7o1a
kTXqJKP3ZuurBZSyCxQ2AtfxKeWchvKSplvnMye3v++2FGVw4qyR0TfrEmP+UzCGaeh1yFNOJ+Vo
Cnqr7TPstwYh3Kq8RQ8tbTc4y2R68xZ/r153gxP/Ur0GS+XbNDwTVFzTm/mFoX8Yhzngn8bsDL5l
W0ZjFuwPPtyREYw/uohiXBvV1c5WUW/eqZP1/7wxxYRETYk6298L97AYNOsEULODTMK/wLPbylnx
GLJ99XYD8ufr5A3Qb06JD+A0PrTxjfx40VMwxbsKftvlfHHpI/cc7M8xCwxgOV486dQt3RAVhIo4
WeTX0sm05ZaL0j72x2d7f1DPrMjxLzdd6X9JbVw8ATlkgYIns4qJcPZsSJ5vjXFpr1jaaamTI3lo
UXs4whlm1+QV71fQzERZOpcd5VAr2mBU6mSSl2WZFJHxlDAWORcmA5V1fQjm++TvEdRu3CM2MDdq
3NiLpTv9mLAo0xjeUxXwYQaUciIPXpvOtA94n1ad/+E1HaaW9oyZIv7kDL7FeSY08/w1beB9AZ9h
GB8UmIEw+hsxWXF1CnG3fzmRNLU0WS9FbNU4JS9FN4xbt5reMKGyvgzTDq6Fv+hLzLdl1YrcY3VN
XXaET3ky3xC+Y7oQ39HpXdaaadk25TY+CpJq2KjKVr1pPSZoT5UjvR83PuuqwYocaaV4oPJdDZme
Rupgcx57ugybhXnpvOzjWtuPYz9iIxw838w00mdK9x+HptueAxLf1B3Mvp5/bd/RCCX2aPqYoT2H
uj8e8w1X4L4X3SvO9RFRFzUqIVQEGPuARhJKRUy8q3Q2OziUh7XrXPSiTnhxyG6wa9ZajjzvYGXY
lFJ7xEgI697Bb2uePmukijuqFXeQHMmmyRcLvT9FqDkTi/29Qsou1/DmT95brKYYBnKxL/I9Kqdi
Jy6Eo8S7VNOErI5vBC8ksI+QoKVSxrzqwjGF22hoyDKk0d/oNlRiyVVCz+xPdJd1kSs/MLWnCgt3
oR762ptmfHVbqXJAJiGEKHks3k3DSs5svslT5AnVvTvQyv/aHU7vo9nCzKjbbyUmfJHuKMuAkI9f
iNcxffnWPrLM12kNQwheQ9jfrAvAjxrVxSnmOI8QFgQCy5NsScnhL2KTpaybQwMJcBH/PgrnzseF
9QvosC8Ea4N6/bwwQ9YzejHk83tnjknDJijTuEf8T3JwWgEKOhjgsKaCA89Mi/f3debRbyqEJEC8
FypBh0fs6xPERd1HbRqSasAm0EpNpwjv1f1z40iTmPWeX7vDykI7HFjQtJkcvEClTNVXZyq0nQwF
XzohFIa1gYsiyCsb1Kd+U7nqNZMYc5v2yf2P/50hcmCFETzReOcNwJjv319OlvVudQR6/Q9FwSqU
duj1Q6Joe8G11V1WtXqv7rSu/6jnIhwkNggWOTVGqZyWf9QGeETbK7AHDYdxKrozY++1Ame2Q+YO
q0OGNXNZvOkkg2lzLHbdeObbh8tQm/TesHPb9rszSDDR0fu4AMjID7beYBXgfu+0asWGWAkoi5DG
4lwWHXKNonia0zTLGnyGDtyqA6GpVRLfUoBIv/+N/t8YZF5vLIreQpbl2fnlUdPr6Rk9GzAcShl7
gPQsHtnwvlOIde7+If67m/NVNxoOiSttoq9eECWFW3Qqenpgw/T6/27wAINFrjCTMO6Wtyi5IOBC
S1ynPlddA+QYGes21GIsLiODjtrB7qCYPQcpjlyCROXL+OKWvJvzV+ABREL6fZcCr5J2sHuX+rYn
ASpXiJS7OIvYFZN2BDqkrIbV1qAl3ed/XLzCQctLzrkfwmGZbsiPr3PxLyse7S7e0/RhOnVIYCbJ
TmSiRCYJ18u+cC4QGfFmToLqJ/Jmw+S1JrNBUS10aW054Xm+lb45b4VY1/63qjeWURui8jhu0XRS
GS93BJTLauxGMHVSD2kNOL247yvUW3udn76DZxjXxFewpdNKMUXvG1AHrIoS2AQewK5/QrwdLbI9
rnqfp/eQJqyqLPh+dyuyQQ/am+qubTETcEn7m3D2Cj+a8lZI6NIT2uK2FprQ1Z8VMIVJXjJfExS5
0PkWG/DkUCG0OfX0dgP+EMwbBNo3Q4HEcN5434ntqpH+iDeCJj7j9LVefn3LjMuYxEXlElq4WuRW
iTkdiQx4O7FmMmBVTOyxEzbb7cSMDd22aTcSZGkMNxY3sBDkQB7g/9LGb6a062zGFXV20rNoUqU1
D0aQsVOlDyQHtMG+/TOmgZxbfyT4O/wtK16dGmTYlGHMUNkYY9L7xw4zz72Di3wSYB7CbQvDKjll
rM3YErQ3MSTnA4PVlg2XnAUXY8tXGf+JhmkfbI6r39/hTXBbu9lNsbApDIRKFfwiRvOUE0xw0Y95
CqXojO45Enci14zqzfIrzopd6v8q6HPgGbuNsjPqDNvWOC2LNovNPmwmB1fbzMhL66a5C5rh4zqm
JIQ4xDbpLxFwmgRssgrWsVbMOJZZ4hoake9sb8Xp7Z7Faa/vbHhHFMSyAs8SMBPuZlZ5dv+NIlKz
LBFUQCmJ2C9HHl5XpR2Ok/pybaPwLBn+ULv7+ZkUkeHFZkYb46ja0p6lGDiSw6WmbbbtwLrylYg5
O+qZvuMDTzvlBVgVFHna9g1BvaIEwNLx8y8H2DE78syr+1zJaQKFlURRdwfCyisXVgmc97ndi4Lz
U7BIABVsKwUnZMbulpm1r9y5mQt1VrT1BNXOgwlR7C0mkUgNrYQiKQcBqONt/U2aQjyH3qeLs0M9
jZZKUEG5epPC7J4eHjBrZ5VsKqrwTiGYbvriEQjh42FGnP3F65RyNlLSrvfnheg8kyOB5Pyc6Urk
/a7duV8BPRQmh2J0f46ny5wTXEmZ6kCtyH1wB4gUQh0o+QDZ3yUKKUIXC5+gkqgGoPbUSs1ORf8I
LdhsfVMemBkYptCH4xQn4qhFC3qHDn23GXq5tCNuUIqBxwACL9cvgrWsLVwdAJNTsx6c8qVbZKhZ
TMcOQ12BLdw4HN1u/YhuDa7r8x+S9kotYx6dLmNzksjSB7kPLBtjyBVRmsFs1duxVmEee7A+tow/
39fcMeKIa1kn+ruWuWKU4g6L5pfuqKhV/qS4Weih2lfIq1sMWJX/cLkUfPcJaQqBV8yCjX651PwL
sq4TrW2aiboZMj0jlklnAcK5S4ZUULA7p/Lai0H0vkMuM/yQ9ZGp6s9hd9AEWu2bA5cJuFROVKYM
5HrNxVVjBy7lnkkVk9qxESKYqBa/3u3Q8TpVjZt78xeYiw2Ofit4Mu48euVQWq2CDmpy8Q5WjrFn
/0lSetzeBm7mnCLY6jWv/S2yVR2FRWkz471i55/bZ/YKgllGd1DH9Clf/c80no1qqHKhqTWEHEY8
tIyHz1jiEz4SpKRPHNOvo3lNwcgBZERXpag62IFxCrX3zlBSkgiS+FiSmhitLtH98V/fu5Qmncfa
oLno3sPFgOArKuKrjuJhxdLVtaqKhRYSo+mg7PIQCUxKgrws0XiZfWGa/WAiPMENoQxQioOGAJSj
0YxdCoMGWxKLZCE87hM7xyzHoFxt2OeMzzgwCycohhNkGiXwk9raVrDn/Te701TZ6XVOdM2WY38S
x7Jp2NpMbl/3N5lYcZ1/d4MdxXRGqoYef5QmskgEv7kL7atBUTa2wlnKwmSL51lBarq/AMEz9+GW
9W5Ik03carfR0RvQ+HsRNBtryZuItktjD46q9a2bunadjsmkWANKibkOOSPRZ+T3l4PpDx5tRkgz
ucXNW+VbNRa+aVBjYq/dW+2325rO8Aa623Rsej6XmTKYII/hiJT73bj++PIDmigS6aM/O37dd6/f
jaqX9zuSVtyUx7luj3G5xvwKsUXtJnKeWgtbJ5x3IBWNohjhbNSb/TyGA0fK2ejTzjxTC6TAYwuX
9FkVnRIIYLYoBD0rgj1pX3Ah7PB5MHRsu5nGwAD6zjeRG3oQIqsh+E0bEUIyaUIVk1zFqvYIHdls
dTk6tgBSHsGMMfWbQmKkkLm4Jbu+iAUj44ywASkHXN8QIe/+7+681TsAcAJvBHMLSCX/4A3ySk+3
Id/6iOqDLRsCcDC9NdgMHbQ1qqAZyvMm/dwUe4/mNGsRn9yb07aar/WJ8asWy3L52cgyBWPxWtW2
Jnmlh7LIeAvWHxYZIFJCN9jbhzC/RXb9eTMuzS+927FgPm4eQ39QQVSEhCiUB8Ko+gZAh1LA8StJ
lJu46nUTPkCDGj9c1AWa7v86W+DQKD35UXiRF/cy83hD3WsZpBbAlxA0j6xbFifATM0mF8CLHDVF
6O9YKtSIU4TUC48gcoPzQqaZ27wcOhxmdox75gd8hVZy3HQVDq/Ej7F32phsm/YRigaOV9EUmgmx
z/Y8VIQkINAZ5Xu0Qno+fWw0/TsCB91xmJ5YIO1ikswTdlh0SheCG0WJzkSVQnhzo2Q2VzsVHl67
mUu9vbDnISr2Xtml8hYYlm8LxFPGBn5RqGVcbsCbBbEo0Cd6MAbFEgAvbiHGrOacE2lMht+1HGfZ
2x95+umlwNotXIGaF9MzGGMN67TaGadlIrFHKzMWaYmiYB0dSDZVH6QQTu9Kf03WnNskl3cy3x48
VrehmJ4qyiay7EdJpyZJWGWmFm5m5q5ejlb7Sgn4gq4sDU4rcbmEIXdd5X7EfQdqHxpYpwdcukzS
4sNHLrB8u4Ds/1gwu3CfYVNaK3XVOIe2BIHZ0T58r/d+wJv7FL0JU/M3vJ65dlaFwXEo1PmUOB9H
0r1hQmTvsoIoTEzOmmTeu1kfiG4q5cG2K9evB4eRC/Zls6xs65qKMSJaIQ1CrMGpCRwku8a2yY+J
HDl8P4OEHOfXi12Kh2Nuz6zr4ffilWbPXBUJ3R3sQ+GdDZ9LUkSePL+5E3nT5r3tMrJ+20n4fDKt
Gn3ptUucYii9aVnrisUUsWf0W6XLWJDL2xzHevrGjRV9iEuDeg6BKSN8mrOfWPMuAotz/hmpTtNZ
91TBafhBiIpmzo6GryIHs8ggDwf9A5uQFonDA57JqWirLA3KlzOVqM300sEY/hVllleI9GB3PupF
TjdneSvRaLQC6SBkBV0RgCuzUotJZmFzmJRmrX8JPD9v6bfWEA2UUXpDI0tYTEH9tdVMr5x8iRjM
BfIe6ZaFztrEUst5QPndPUnXCFnhIeAjmc1cPtodzXzJDTRjYbVK1eatReZvP3UXXFXnA0iBHN5D
VEKUrMOLk/PiBRf6Fr6apV7jj/9BK8mVFOebqKrd9iMe05bALCEuywjrTt7ZMOY7+WCJ5LqgTJjK
WCxq86MwVlPW8jyYXAPb/lc53pPXDj3PQvt3l+u5BgiN3GHxflLJ70uv3cCmmzmIi7v0L5NMid8p
rvBAtnuAURbg6ak3F0DjZVFdlDA1zZU1oSXwDF7jLWzwdVK+gyBSAq3ZVtUppPlTYzM6h/F2TJ45
Aa+Mn7bcU6sUjKmiU9zC0fgPUtoLq/2jRVRpC0sl6SjU7XT0KOqDWK0X5eVTE+KJ8pMdqmlWPaDv
ob9WVWvAdGrbwk8+tqE7rPfZ4WySDOuC0h6eZVpLzJuZ9YJBW6/tT6T2tawQqJM44Rv2TqxpEsWU
JRtqIbAgaTAWt86IismmmXtNhTDzJRYlaZJlCH5qCuaP+UtAmhwaF2cfme8ggcw3uPp7kWi0+Z9A
SvpQOYUDzia8blZH3H2ol06WBlIianyjwzQwWYZzcyt3Dv2laKDedJcH4/sEACq5iieCKhGLllIo
Bq+Pq2tEi4koHwuQBr2M7cQi+U5gShkRKyhaybhmZ6C7cDX6Fef1KPV+hT/aVqeg/2uSloM/IzzJ
MCM70Ax8uOTDrP5/wyaFfUHZOdCIljh6YUJYOlqcu0zrAT3NIdCy+1ZLrqAN5+iR+Nm7Y7K5PJeb
qxT7o0RJ/HhDe/caKhXobOHVT01lQ8H7VnXSWhnXH+ztdt6SJ33pbFOvzsU9aPAR49UyhVyLUxzP
edIHcV/8iJinh5EFuEU72ua1AlMXlVJjE+FNbHTfAIyt3snt3BLY59q82pcAB4UIYJDXPLZ0Xf1K
dfLD6tVj8vs6wqiT3k3Z8YvSdQZI2t2U82+JvFqWBhUaWk1Uk7raqzu4Fm0HwTkBYvc898lL/dxs
FCLRFUoV8grXZObokreG16hzoVRgtxIZPqlmtFE6D4uy95TWBsYeDvd10eLFaoWiZjWOr83+Svwf
+Ch+LvosTaJI0V2+kwSB9MdYiQahJIEFYqzxX3JKk5HxBDClALc0bfLRWLotoYsJI5QTVf3vS16N
JLJlLzn7ECaLFCiBiYmdIE0oWHzqFBCFySpk3PNE047Hzeac1TA88zDHmXiulJ/K9TxpgKK1Ts2B
TGOxpZFZPXgJR6zivv3gHYLV8VDC7rRdIwXcq+/m1xVAubW0hHsDfiZQnT1CI1poKv7/+qN8hCKR
vC/raBTe2KKMfgSpY4+9mHcQTP5bJ+sWEJcgC29tEe2E4BFjhn6+ZprhZYKfd12E4q4NoGY0P2QT
ujGVh8Q98iuG6E2/Yzzz4EMfeX0q51OKY7r8f6vYw6sfgeKyso5jdFIimV9zxOUV5qzfVSI+pR91
kJb1rJJrDtZEaMhtzN2n1eEfFbKwApBuamXB33+gQNW4fADwK44Nu9GX9IEQUhFXULquH0Eb9IOM
Lq9gD/NfxDPJMny6iOPyt9JPthw6FXB3OUX5SAO5UBCicAfrTRB0rhAsslLI0eojxCUA4yAEYr/M
rMk11fHTcJtpEyN2qWlzqAD6UVUMsY2/x7mJxLvZRPUqUxRrQxZAJLGUOvkujwOOsxjKIW8hZJ9l
YtXnzC/z3SVz5sgAtUkBNEmCp+Iu6lvhWfWVIzjvNOpGDT0yl3Hx+7393BKIkWEMV2OGXc0snEpX
H6Iaq6WAKkqaQoYu4j5Ygb34UciJop4v1emac+XtXzK9HVyVWtnJDp1fSFfJuBcNE8pqrkgcCpbj
MSdNjrGYnOEE8YIn4nsogn+4jVjESwa58BhlQ11kBGPc2VP+2Kq7W4OFXquO+MSu3Tmx3+3nWFql
3wuWP/380QfnrwixEXqycwck1buIxTfnf1GjugcSClCt/11A+OP1k5BWQrTbwoql/qVjT9Aq8K50
gkQyj3m8bqKYR+nSATnZ6hmDw3RJ8MeMKY38tnTdsJDIAkGB/rtuGNDugvqkPfXeyWWdjq5EEOKr
2ku0+mRtVdN8HGXjTqdk9g85pBBOpiHCdWlv1QmtC0YTqeayNnHgqx/zxblv/SFeTJrHr61IgFgf
0FsaKjrrNqN1vxBNuOk0E0DJxjrxx+kAATQcW/ytyfL5WOTfvAX/ohM+t1shtR1R9hN55TyQGG/3
rLuyI1uWcYkSZgJZMscXA+dJCiGUMHPiq/ibpzK+X5rCRIhgSk9rNS19mf6bfAZpbJlLkKU3hLcC
BvpUJRmOSMmi83OHQnjpVj9JTng8VMCBbphqooibFOckPx+ID0FAvK6org36w/VgcPovEOx4PCWh
UxYVNGFl8F2oF8Wi3i7aYmjf80Zp0TYMsXG4g8dbRyctppkMajH/T2TenC9/O7s91VkJ1hn1fPbu
iC+K3vq09CkFfTx0kyg4kmDWPt6b9cmGWLf61WKmwtzVHzqobWNUJzKit76DDFt7ULdQWxeGqtX4
3W1m/V14yawW+/QU6nPKnscK3vFYfwyFReTsleG7peboKaEB+u2jfb6Agl/HWdUUpBqWAez5KDfG
uvjdaRjglh9LfZ4eNA9nrYsdFClk/nwT+AT4nrBkgDprT6x3bsHeV71y4PwADbOBRvGsFQMUsBep
rVP0NSZF74GNRBrz/hFVSdw+LCnlTrjG0NVIeTMlOZx4Bb8Ee2Lr3xApFbeV1ERPlYwF7DIacUOi
c8U9WmYSQk9qXLnj07/FSFbHSn3vRrNJhz+t8zRm90TtFy50aBPcIRpo+/A80O4/DaCezuqp9wKk
uZQcE7s0ccUO+wCUmOGLgKvNUzSKmCCF+TxgAG0SwpqVl8Tw02QkgXsqrOblMXQThR/AZOCiy6yH
5hPsBDXFjIdpnaJ5lNOetX4DQ5F0Ku0HsqrLHy3jWJyp6ZUhnGuE5SrEtoiZ8qJpGAo7og9Tq8Mz
FBgwXj0RJbKdvG1KW/5NMoZgUp0rU4/LZ7h0uh+AV5bjUpmKAyIJK0KH5zsboKdmaXcZMm/6yjf0
qBbvHkgX2WE7ZojD5JLaTiuHxM6lAiz3cmRVveWrBIdXzr4Ra8m/INii9HiOSNXLGpFucMdVEMOW
jN/3MwhDZ3JAv0SVnN5jr/2ojCMqRgbrdzbUXueU7ZWRdhFAQ2NwJqpCvr/KDZoskQ8Idxbc4DUb
UJ0gvcspoRejMuYiPl0pDrT/U/l2vL+GdocuHcWmQNIjcvn6BYcJG5Ypu5J/NAM/XvSwA6v3rMF/
uAJTi9NPw6YeuYIdbyC4nqCNzye3taFocfZeaAhapr+h8oubKxejf6OuiPegHZAm1yvKI/g4aALI
Ft/DlM2oB0fyHVcDp/mvezLTQuvXN/6LqfIjc8gYDwT8sxO6VRLBExngNxnN6tpfm5ctG8Jfjg2N
9+7dtdZ6wRhBCfiUHMISuRPpDoi6HVoEkAdI9Xjoka3zB3GzzQP3mF9GnxCIkUwWZYZH/PpDGuDj
23bJJUaE/h27YdYt5MSsVTq5mwAYuoGD/CuRFT2d/bmn4WOK8+wCwG8OoecxW5bbo/aYElOu6vsf
6WrARtPDyVjb/4lRHTWoqgycSE6qtMrV+toTgpt4qXyV8QvbpX2kcMV6LqZYakP/vFANFlxXWbf9
3I1J50sB5K404e7SMLUl/w2LRbIzpJvGjcZu29vh5ZI5oVFFxm2dNTimuEmAheWmRkOYPsbOk5o+
QvEroxa1EOfRHB0HUhwHV/SrGD56nfXU9ij7qhG0WjnOvPK0yhAIxydr0b4eAUH8G7YOcYn+V/HL
kQPJ5rY/xI0rtO2y9pRPw/cMo+jTc4Pp4nAeGaMBtsaYO7/Gv+06vcZta0t14lmq58zIIR+JHEab
GZapRKry0tHyN3PEZdM/Cknj6YP0wr+9QLTkfP8Qoomp/Cz9hkjXGmIStCs7LaZW2trDSlHa4hdz
MPUehSyzPeDJqzPj9taCh9NZQhxE/219JtPUq0QObrrwVIRohUOQCBdCKpOvqcTK2dV3SndN39yQ
wCbAxYcWjHBjY0qLuJ89geiT9wbdsikpcKSvGx/uEjPb9iR0/uQPj2+Xb7yZJs3KAdIeLu9KZxjQ
eEdV/g5SkkW2Ieu42MkJqVCeWOBLOyRbpxkoWJlU8x3jOIkTFJHn6b3SEau2dx4aXSrjk3ZN45Rd
XGpS/SjPkhxz2JkAVoJclvPSegzk557wPDffU8yh2A63ZnqlsBsJDGG+WYdnUaYdqpQKPEppztVX
dLtDO+dGdxdW/enZXFv3QRacaGCqtU+4bGjZYO33/vHcczsAUBP9uEGNUdPnDVBUZxfNU/ucUvCo
rACIPX/N4TBv2vY2my4d9kDF7P4dGNPnRVTEl7EcUQf99/bAd/9KsDTiYadl9xOm0tbq35zGsCcW
s4m2lGzitstkNL+RE6Kh6DtEbluE7hogDXaClVZoABmC8gj8i10dXsYm/0lT0RUA0ngV+i9PbWOd
CLdYOpW1QMjU6pcBr2gUqFPBWIR/K71pd62qILkD5Lt4jb8UVDwptO1amJkLPCPvbKf01+d3+QM+
AnztWdTKyBIA8opSGQJkicx0ohBUotUjhg/N9Wlu4V8mV+pdweYXR7aYpBzCxa7KFVblzLbRbDaO
eavWM5d9enm9hEp9iBZigO1L7RgZO1GRa/MO09hTo2882Gbgeg8+R7gwKj4FE/nCM16yZJ8MbXa1
kx2ZIvVGfm0clFW8nBubS+HGeDiuJY0Dh75JZVW2KJFcjj60YmKAKNUKpn1SxAftACmcEJU+oATJ
c7GdaXi3f+Kf74oIJvRa7cYuVlEgiMXusTPgIrqKth2qQSIvnkexs2YO2UufF7XZ+fcu6tcEPFg+
ksiO0pJ8AI/EumhutmFhTpM2v5iWZeCafCLYYd4vR8rKQ1R/bcjhXt6AdaqpL17L/c6rlufYaEBD
nwrMlxf3n6XDFFCfe8iI5RFx+uzvq8rOWZuedz6BGIml7+ZpO6+N6FCUZ7UuTqi2cihDCqUY3FER
0b8FjWAD+p2Sxi1wJ6sn/QwDCTQ0h8ZzLDg3n9EsUgTfcw/SKffwVdvtZ92IppcvjhkCPx+rBHtU
0vq8S+sJpn/5JevEAPBeoK/PcKYcaJIw07KvYpmx4fIHC8M5U2VwwruXngbDFX7eUMEv3jM77R57
UchDMddOs8gSIfZcQFLbo+izRlIfLB5RX9YUNKKq0MmBalWL7tu9SlM4+Kxi2GKrH+AlkT/kXeN7
uNXajqMQVCLkactXU2FNfLY0bxLC62KW288utyjRNgi4m8YyRpVu19WnxGQZy2DszO/Jo60BAmfJ
YBVBihZNaSj5EUSDRnrGViNF6bd4mDB5/2dRvJs4wJ5EWaCAjzVVcCxVDQ4KKh6a5uiTu7bLKHHq
NvMdcnLBJac8A4OVGyO0pq6QylKlcxh+Rl79DD01VP2kHPQRkIXsmusZWZqgVUt6mz5zETupqC15
3NgKZphN4nIrxIq7/U9zPnWkK90NYFdmijvsbTSNWnhtOzSjmVnYLODbQ0BwAx5i3mfkIlmYbUET
Cy+WbzdR7EHorfrxhGSHPB9eh0ltovFR3r0WcejNFtuHRZgzlMT4dnJauRHBxeidzrKrs7TB1Ojt
9v3C3R+koMpQPIcypaZAPb73iZ/cKK+/1bj7xuYtcPVHq9ve1no2mg92dt/oujqonS9YITCmcQF4
R0wfDgjObc2ahZ32GpdCX4jjIToHU6twOGPCHA/CLthKjUIURRzca/c0u3sy7vI6OAnGAqYQfezk
RErKB0eNlaOt+E1Csze5SY80+QGHzGPHPAt0IGQnW4fGjicVbVEt9bx/S/c8/N/txD9W+xi11c97
BQ/wydxVA/v4yncR4sRiZlc+Iz3d+sawNMDy0iihW4kXzk/dWdVgOwBmwS29RUBTuLpDqgJat6th
ABYUI0EFAAI3ueNDesAQT37z0LTfF336J6Mv1dvzkW2dl6ubDdann9bP5slmINBsbx6ji8vwX1JU
IWpX7VAp6gXxhI4K6erARWqI6gxP4rOWD+bl2VRcI2oOWrqA101b8VInADgPqB6LLS3xP08Av6WO
k/EQoW3lhovSU9cfam5xsqg9HDxZAqNKypIsGrtViNVYzlTED1aWh/amlVP9AF/A3Zy9R/K8D6IB
HDVzWjoEn/08mFlxCexrcWvqqVYPZyH3OrQTS8za9CM4Sz1vAE02ZOxQnvhMU4mvOpc951kXA3FQ
wI2al9cT4wQcNiCCA82QWIT8FrUER0J2+uMr2SkGRsKySRNer7Tq/KlXaFkqIt1gseH5/vH5mke4
LRk5n3ZzSKKAPG+PnMt+3KsOtz+MAm1qi9CrsQXD4qZIkSffw8e7D69ykJyzf0Y6jikgvr5aT1uy
L9L/2KbOHrRo+f2x/PLGeq/1EeJdKQywhpKLlgh03EWcZIFMq8OjWPKCyIYdNzTohExbA0S31lHb
Bmh9Mb1XlqHIX6O7Xqsw1XRDkW2qw3erMdvipGnTZTJAgIB7Un3aibGbgKjHynFNbQR7KLI9qH5n
iwl5cTtTlSCVGvJX/ZKqhLVjueR1wXNJDVUFz7MquCXAeKXe6dQfpkN5GVdbtZrIv8K6Pern7L9z
En+WUErlqc6ZYPD3seCy9LX+2czDgUeQPJfqIFlJw6BtFQu81fzP6mz7RdUmYkZt/cIWBw+KFFiP
/Pn32fdpydxC/Sa74AWwhB/hiaQfCC2LZ5b5cb85pW+qMBWNFRM7B2bWPfXgmjDLQI+b7imXUN7x
kGboQ9N5aSeUxklsO5HoSKp7cZtJIfk1eAYs84zvoN5EgDWaUL3HrFZZhsJSIez6kJEgpgHKViW9
mwfXmOQYPmjYN8Ps64xsfJQlLxOJmOOuOdwbFf5wUuQtyigp2TALb3+YWadCLVJDsfqRhiWlKX2P
V3pbaLvhTXs656qSbwOpO17iHt/0K3WDRtcJoEsdxgOucHkkrtkukYLbNGUn29FSXwDI8ESGNiYp
f77+EuTxkvVD4h2X/2/vOWJcLhp1dy7GcoInoQkQzjqyvCla2cV51NT2a+bLBW1S3LeKP8zbYIBO
p3GrIU4FzkGKz5dwG0nfUyNYuSqe90ues0o6SBvLSFGBRIlfIQcuZZa1YM0svxA6uqvl3M1E4I3Q
2nmpswDmp6sSLdQrnPnUI3fFlAl90pnDjnOQmdD2x4UEd46n+tjl3T/x+50Gwm+LHrc3VK00Tr6h
rRHQQn0Hz5rN2lq9ymD5p0eUBP6m/xnw3RclPIAK0xAGB7fMcvuDXn4/Augm4mLtq6e+Jg7LObEj
NP5mQjI1Hvzbc82WDM/6o6b8t7zZC1QJ+OGN7E0r99lL6RfixwOgD9KHRO1cXeL0ZPExdoGpGSLX
QVFyKBsIb9RT0T0GChLs5bribx0ZVhWt+jwwGsqXt8j27m/WeYvgpJgiY8sOujMcxl5hc9aU0AIi
Ze3BFYzF0KbEY9Z5+CpBdkWmbYpLHjBO53x+XwYmolxX3OWPTlhcZmdbrl2AMCQt+XzMZ7L08o2y
jDRb9bRA40/t0sUlzo1wpgG6nBGjOQ98jDSh5en6FVfaX9hjhT3k54qe2kfa6KK1UaP5CjmPKVd3
Re9okzq4ualMXyTQj/LwAEHYScJC8cZT9ljuBu+bcnSuygO3toyCbOawtsdBiJekOrftzm7vqx3x
MGY3ANIFaLAOOU0ja/w+BYwpxvZ7qYH3JF5DsnnxCyEObL95q143Sx1qccFEViiMmO59/j00AjLF
uCAhV7MiDFzcBs59codMuwtJUcryEkUO8c5oP3LcC8vcGpQyKU69T3WBqbmiTxmvU9XmS6kSwCte
303txaCMA50JgX/Of/41uoSkj8hxVzWLQHi4WNqONGZ6wXKmwZTC88VxD5rRhyk53SQaO+Wu8/pZ
Tc7rdPd3SEOTgjqUpY1ltR4Lfzg0+tyVths75Qbx0k9xh8X1vK3rlFHrXm0za7afH8+nSeLBCsno
8JXENndbfAQ0i5mv7maZA6C79mwsOJR6XK+DzrMCyO5mhz4A4FD6ewEN0FVnNcUHaQq7vFzzaxci
gJwRs/BU4L6VoMmXks1gnyGzK0Rs+JV3SjZ5yosfOyJSe1O+5OTyj5lAF9P7onGHx/dJvBgFuYX9
lkXeUP9Q3qBRh63A9bmnpVRxuXx5ovbkgsG14c/ApYX/ue2u8ArT1udD/5MD+l2tBZf7yyFTjQlA
sOKDQbqvqWYqbrKKqZd5eHT0L/YkEeDeQQVk8G7Qu1kKbmdy4pxjFLGjXfgAPqz+ys21VKvlyJvo
3OPjGgjqUgkpcvMFxO54phEYaxB9eq9IoGAqRltTwxM+I7B2X0gZFpGmOgpFOBWHjFSl/qXcnENP
evEjblka1rQR0LCTA7fp0wtv7XmeLHdOYeI2EfB98kDJEaINO5UswvYZ8AAz+y8gWdUH5uV6LylU
URfPnRvdpaCsYlEMV304hUNeD3pl0hxdTjyEsehaMQegMrNeRgmN65J5hIy5VHJIXXlY7zgL1KiT
kFyaJ/PIwhOBI2ZWbpxVEDY5KRSOo0wKx4q85UThOF3/LJ+68eG5yoqw5xRjV5vgpu0LBCIji8CV
SmZ+bQLBWoce95s7H/e+CitLuBrMy4Oa4n9tA/xw8XJpnDMJyFCmZX0aWeBcikynlNazDUT+YBXu
DCwVUnpm/SWrlMorB4UBmMm7f/hxB8BYebJ6eSQiWc92LldW0dXXIIDBtz9eNdeevNz+U+fOqd1q
5MUgmNZqkpEqpxSEC5tstTWVcWkKH0Ne14S3gE0Jj50EMwROLqcyzzWZAFGWCb3aMKMfB0dPjT+6
caD067DfKNsqR8Tts8UtEtV/jHlm1PHhqU9MuiVt5Lxc7m6aC38F68Li2FrzZLQUSdweZltaICYY
hx7/WO/1Lze9Eip5iDi6n5oNlYk2Q2giiwoKCvThZGDdVdegUgB+5r6BEL3vGlMxfKHJf5Cxp6SL
q4N4d7EIggIt4KfCyBNTkxRcDBT7HYEdCA5T14vJGZ+hN1OIfhIAQ4bxJrCJIIosBkTk+p3CK0Uu
sRFdH7T9XSdoCh3UJ+svNXfF4kHbMYStunOt8QirYsh6V2EKUCV/LsBZJPx8+EGewLwF6zazfprs
cyoJqG5uSemVAppsoRATp8f1cExvYRJPdlJXMvBTwFa7QRksNGvCM1OZv7tB0AgVnvg3LPqwHxWP
gOKKYEd3Xa5z9NT/hMBT31WVKyoKUbDc02zcxKYuplEpCbHYiDdTcYbb5Pv7J+VWEYRyXDoutKrB
0baKglGTeXlKKySyEB+Di3T7Qrza7HHtAK1b1rkWl58KZ8PAthv9kxxzH5zV9LqV1rsQI1lTcGPZ
NdDcaDdoeUw8/zmkrNZd534pqbbxM2ZebAlLNvzqI/g6QuP2m2iW6DeiJiqn4qEYXS/pqglM5iE6
QNfO4sYc+B3wAf/Mn4vIYhDH7fKM/uR1LCdK/WSC6/ynS6asvA+sDkqw4qwvDl+ib/u6P9KFXhAn
DzWFqMQ2GatricS6O7sFQd1IJfFwGx70kFQV3TiM/2l1DM/w7GnbmOgasR6N+526UUyLkKqSTxz6
HpOUJOpuudikBgUvXQYgvQjJoyAPCBMJdSL70E2fo6ZBWGv/hU0xFli92580QdXx4oM+jtAiAcI1
KL/l3/1MdMqRDUIgx4IjwrTZ4EdD+jlGKBA3dv5yQVg6rt3Rh9lCxIHWmetTcCsELL0Rq500hv2A
c9nw4NbWRnutumARCWckAPrvBZL2v7DsR5h/+qoWj5DzM0d5Uy4rOT1wsgxUUFJ5yDl077TEp9Xi
+uGvlDrmmjPxbbmq2ZzkDpb92QulE6yyq3u92Ig6Rwso57K51fJfNUcyJoYSfPUmiOZxDnMSuU2M
i+9Bpcb7wRgWXeoBuGn3M51Trk418E2pg9PYoin+4axMd6Pljju2St2LlZrRtDns4Y57FTVsqbxp
GFed/cMek5i8zw4eKF+ApELprF26sgkIWKqwFEqC6UmvPyo4t4z6RBTZedk77wYw2Hg/CspVTfl0
9VgOWy3X7bPr9B0XS3zzxiWddtKgnRuV0MmfEAWH//sjjLWWJBvXcw53WAPYPaPs062I9wnplHpw
7xRc2u7R55NOhajlyhrS8LZQNMOPicEwG1Xp0BRPrupWU9iBbeUqEcP9vbbnABBy7i4kjvcnX9Yd
+VESMlCu8xbywM+zkNSIdQnGsqkxN/9aUfG88Ts1eq/6FblbSYE9RUCqt4o8C9wwYcspuNygooDE
hQ16aETItujRIjVoFyaraWEqWYgVjmqogle6X2vzctwCMJVnZV8BHt16WTjAe7Z1p1BCtBo+j03D
yFrUVNXaxoIaOBpAqkjV/ukxbz3trCyjtk63mww8leJsNVt4c7I164AancwdmeONMuD4l9DpDHCL
OoSMALnVfMCAVlA0oFuNHadFVsQV2vAOrlvxtLee5tlWCd9gtL4PAr8XdAHR4rskVU4BGOiaSEoF
Le4zgNza6a7SVRXAr1PToQ5hm443ckCUbaBTz7zIR5qVczmFz0HMgOR3q+KOICBLIhaZRVG4R5gD
MizZAmpr962CX9KaYnbm/EZtMWmZaihCAkO91i76ULjA+7gZ9TxbYKBKNxghENDJ1HfYwvB0sBz0
X21/EEL3VyKdLzXyZHbVe8eBJlc9oE+nOVrnmPt14nKvrek905ZDCRSsH91aN4Cp5D4fVjtdmG1E
V51QA4nEWK6S4sdcjXaDAEPcoRt/MXrAxC4NcklqvwkprR/jFqkELL/VYpL1rUxzSObcsj1nsZpy
U4Qy4v7g8vOfwmLDNTI5LQCUX70IwKjiOj+b1NMXAenorsAP0wsjV+YWIpum74DTHpFSdCpfASvb
HSWlYBCr44OVvmEpDmg66rQti4JRj4pxmW5Bzd+GesVwDIuyeZcSwOHNaWqmdHW1fPKwsRDt2r8R
mJPNtPewznSiAsK9AO95oRoc1PvAejDo1BRhpr6g5q1SF5aDqaaNnPzCu7YwXl07i/Co2nGkhvOG
SZMDJsgtinVTR3gG20ODFwES3qJ/MK59EtIMVQVcKhMb1/W7LQZzgPrC7hVMGPnHDjupYYzizPna
NUZitkMvdAUUFUTuXin3RrvTK/u0ynlU1cFYU0KZpBH/IIzGuslj7umAE91Z5z++JxoRbZyuDlHB
Go+JMM0WWhCh5Zue+kWARzPBoqWXhcG/CGsF0V0QIIl2rwUfVECTHjT9ij0u226jgfUzfDP8slnP
IMncpDdNna18DYf53GqwFL1pD6cu5ZOz0ArudaxNy7EX1NO7P3nYVx+NlgHhhUC/yEKOHnrE5lbS
ZMoXQtF3ic4EYI+Q52tnlwgulgpeZ8BC/Gtj5PQPmx+9IkZuPiI0yWfYifGljGj6BG0+GSLf4tra
XaS1q3p3PMgE1JKrnY9q4RVp0WxPaafYfRW+97u/lQZ8qxmm1PCtPAEsA6lTLz5BHtrYw/vUtx/N
DmLeaEsB1HZT0FSz45r/2vx0d9m+cVpH/YLuWyHtWMmrZUD4g93d4lQ726929YB3BcMBy0hk8fMY
jJ8dV9JDtM+NPm9p1aEtfLGCdsDAa1B7K3hR+cc3K0+6HAcmklM1YcKSDVdBeTnyUwmGRMuEuUT2
oKOCCKYlVmmL6lbQTPJ3p3AaoFTwtvW+4NTTbhB7UleFBHhRhekuK1PSa/J7jqsj3hsEkNEWVEk2
jviqIF4XZFNLJl4AImjVKNUQRqHubuEqqdVepMUbCvQIGTTPNbxCIZsnTrN3Vl6JS+xOJyWEJhqe
Vzg7j7NyfA/w9hU7Hi/nIc680IbE1C7rpoAJuYRf8Sqpu3ZXIChz9UQ5ZECbJcxVFqYlp5NF54pN
Hmzn5/f5lCnsMnGjZpXJjHDZOLLLqeFw+nFr0T4bRjAgfbuTX817SFUwDL0FD34yN2RxIvE1Z7RI
tJBaXD6WxJu2hahAlUSdhybna5ZEUndRh7XWv1D1CWX6shq5SvrizI7vbYFXV/5veGXwu9KPwv/w
DI4n4I7oR+rYFIjX12a8mUFttJjnoNJTNMZKrDFPUT2//iAGbRtpn5i+/4TDFxUP1aovlGPSvoO0
4tt+uM/GPT8bWmWREjbXH2e7+p2B6Mrbgaw0cYm8ObdORQbEFNEgFIEwRppYve0PIBAASmZtK1k0
8rJ12iW4BSrnmdRtsXBoj1ZRXh0BP2czV+3lgmNYaw26z08Q9iPk9HV8JQslmMNl1M0BGxGwK/DW
MSYvUqUIrWeDk77qG63mk5ewguZ6MsTnnxFGO4qReRqYClbskg507fVihf9VZjKPgdmn3SEM9n06
lfeTHfcc5zYQftWKcAh10EPv5lzXlrP/2to3WCjlMAfUzPz8EGcNZXgsgxbrbC9PdyYC1i+k8t+x
/JkR7JR3xcrbsn+dxCb8nO/LTOO+eCJCH1QE2sTVHHs7DykEAuNlCW/llOJxYSrRRWKOich/9DvA
eEK+hydYaPLGF9mTwYfC3TZAdyYk8IYOWdmP3+tzWzz8wjqJfDTc4ibuzZiVKO4MFAOlxkdwhR++
kLTU51/lvyWmdoEkGH9Kg3shnlmjDj6Kbewr7ySNftO6HS3CryeL3VJl3pxnjtkVXkrIOX9a0wys
LMIh9nSlbRC0jQvOeHTTTMRqbnUzb7GTNZGA+EdR8WuLVRQdPh7AdYgRXCVGTDP32EwudibmVb5d
RJ9xXXR4i7Ljs98my6cbarXXcoiP9ApjLDy0um5z7/wf2dgYOCAiq0km2n8otN0KCmp+nWJ+NKL2
K53uusdRJJ12qgm6Uh7DnGq0oEyeUJBhrmWPLyyAQNdsVDmOW+49NIzMwG0J4lDZhAiGc6+26QBD
NTWSoi2y9aiC4LNFp2XtbyYG3guWOHziycu6Q3NcesoYmWYANuEFpyy2JsZ9yI0OaI2VeCqOMYJi
EdKcf/cOno+/EjHRFMuRMG9VqtURVXEOa+Y4p5OasQPxw61s7iN0ZJ9uqx2TwG7JsSYL7VK7qaGS
X4x2wEqYyLH89xUAEo3Ob/TI49/glR1IXp+T2ud6P2W+FeUDslU8mt4vLjp5ggR3ndRy7VgDkfGT
Sd0FKooyF177YOEV/9ygiUbOrmZFnFgMk4E9Nq7SiyLZirtaC0mWEEyE74ksottMHLZLvtxUTjEX
/0MHr80D4o7jZ8r8Sj8XgAix3TPqo/Ig8X/yFWIaFsY/f5F6fsulJEehIZXM3HwWc/KNIOafOQir
nZ+3SctGRrP/bPjgnahh9nUraG1fsm+lLE/3m2oFYnQraGn7fl8+d9VR2FPv53LAzVYCmVWtf4UX
d2a8nyUqSaA/OCNARRIYRiHTg3fzIdPF3iWazI68K5WpOh8+a4Z9iRaJVl17QHjaJ/u9rdky7xxX
FjF3lm4Wrp0dSOjZeOIwp5bmO7Mje8Lu/sbMk19rYtaqWYcHHnSdKj5MqdYi4m9lLR53CJA3SpPE
VYIngNI7ytVgAUCqkrGbj03csnXVBqo50QBXs5/a91LCVt7Vj+wn2mWWOV/oPGtSxVSmX4rOVMyb
muU4ats3srShRYEXoKmcuTLRnEaZx7sLStYmZ+uItvwnclB5B11zO8wbqedvLczLrFVtZhZaeZTw
+0AnNTVXrhz/jOf4F40gQ/eFC9epQrIa4vndWeJI/+EsUj2NGOz5c281fp9z6f6A+YhdIHKID7GU
67W77m/V+vpm+/a/W31sdwFuuktsYRjbprQOd1KlCYJQHUfpwUceC2HAI246LNEd7Zd9MgKnGmai
0neraLQI+bpouOZjxyLKYwKtLq6iVo3GmBOrtVQ74NId2mYC6mBEYBHXicvu1rcJHe7e1XrsWrGO
jXzkpGgY967Tzui5f0jbjRE04JD/QL7PvIqCgp2Z+w0BBacezz57lVBOHjOl3IMStLcniMHxJPpt
n2Lk4Pgq3Fhaj6yh8pjL8x1OEZpV5EjZZgiXnLRhpdS0wP6fjz1opnZDp/CBd0jnsy5G9Zqu2MeZ
ShjGXhseCMV9CGvVyEQ5NJbm60uCsxDcju8msi4eHGZhv+wUhZjKh8FwN4RtQnjKzcFjBrlXdGwX
e3R4TVPSmNpd5dnKRA7kXwW2NAH+XLpEQfdnWjHdepH1bEAIHqyVteduflcu1c8HLXOlU0IC2b1O
0+yuBTh0bTKAvVoh/aexbwXBZDO971JIqo8DpHRwAzhe8O9b6e2r/r9eU7kxhjbY+h2cxzVaoms2
YNB3lKw3svEbPquIi9Pq/7YBPEEotRNZdqjRL/V/3u3kTxrKkQgn7MNDwBPsezfpNohzzSYvJSou
ACjnPQ2wiaefosD3Y+vUcBYoWmFOhVu1Rq3/OAkzveWWYOF503rkBiPged7/RqrGceR5OGFJqGM2
DBAHcr0RFKwYQf8fP7crBvJZ27T0Mu5NKQKVuBvWZhwH/AJpNc7S2c0oI6Oiped0POCWT5AV7v31
JZuWKwM2j9UU/2r5A7/j6fJ139rRE5q5QZac1tDa0Jg2/Co/goK1LHtWdMKfwakLzG3nIbo/MK2f
U4QF3QW5U0mtGl8DqnesOngK4f69NenC+kDNdLVnuUeKjAOoxBD1SXkdwwzeg1egLsfNLquwdyfU
Gr+HsrYsb2XU6xKYUpRXzbZ6ekDVrxXAVWLupGgUUTCDjdLbqTE13lWu+NczODHwzCQpwq5v1cD8
Xl49/1q/UeOhs/paL9rcPHbBpcL+auuQ4D4JSh1gNavzGg+rgE9dnmH8vS8ez1F6lMjnl8kJBS8G
fUs6WmRh33Tx/Djgt+TK3FaLBePvbf12QlAuJWRnHGeFT2RnFHZfZj7oSnvWWZaeibVq4H++1kOT
1Nrd+bh9cPN93BRTm7qVrwX5ZICMXzAZk73tezx5StaHJu/C6Lg4OqGWM0OV+pt6yxnCUPp77nYP
BIgSVvnuhKhIE3V43VTLjydeOSvMH3EIfd+ARHULqlr7NuhxTPldMT23PEwKKgWvn0OASDo2rZdG
o459HlWW99U4lefWdMJPNocWZ3D29HOaqJ33V+g+2lBrCzIySKlBdBSYFfWIj35z0fdKcDiegOmh
7goI/BEeuMzUPTruTIvmwO2BNUeEw1cRzA5Ub5EjKQKg1orSPM0JDULcXJfHNuXAAeQ/LgoPrMt0
Je1zV+sEPsSIUdxDdahPwlSNKnVBziAgaJiri4MCpfifvP1HUSRgVbhDsXFnUEikJBhO0mOJDrj4
xniU+9IpqWzD9pjFbdoTniDKNY1IvFvVC8bodMBuG9k6/iVDDWO4kwUWdgvXARNZ2WVqxayB8Gbb
z4vXcwsBMR4J3An75exKmRQ1HIq7VVoDwrfoFMhKT/ZaP4Po067gXZTVYpVlLDQ/ia+/aQXIE1JM
rz1WN5Mwgi7JueYJ4VAB6cBfJOf+nXDRmJIGf3SypsMd/QxxYmbVJdOZKhligv2RXOzt53Ipp5y5
QkXFu3S5+WSOVkkXSfWhois2O0iKSwulgxEwWsmwDQ55MHXcwMSiEoaswWG8yPmJ2ZVMMsOnSt9z
7l7tqRE5iYz9cTnAfQ/xVijcYHzPLqlbpvjm2bXB0WGgtbePgn3ierWeWVsiyNpVOAbgqTq8IRVj
Q2VqoXAa2ftJgLcFHc8nuahQso3HT0C8nD2NqNzzSDkZc9TRUNY2ehs6y49sm678jq+cBr0BgemF
rzxRxJX0ckExRRHQhdKBeOJt8rmshqoxpp+ngWwsWu/6JgGCdT8gxGCOrpczWFzAQkYtLm6UW2fx
rAWI4OxqZ0mR9Nf2Skz8OKb6Y7KjpFS1vRj/XyOBV5sW5vMjc+OjUaDGa30JfQhrDFL5iu8Pb7J/
Ql92lqEGcJBgwnfOk6u7/aCyOedAucIT9g8BXmENMkYNzXFJ3apYru7kvk0quJWnJEYCyY42eIRY
SViyj9KTlKhkUc5VH4aIzckWiJltJ9hHm7DBP6BdFSvHydQAjoLMNINsI1lhp8FQlVFiMZtmUayB
CHGsZjyThKAgE22yTxkU8oE2HpwayYCBT7XTQyOQdmExVdgrtxsuX4Dd9zkZdsncejfRvFLL5piP
uhCe9LNMGcjuLsji4bSgyrPUh0u0+hvxy3DQ2cF65ONtzzEQEB0lXMhJpFdav/97x+k5zmCVD8op
qqZ+iaLcoYN0qvtoE1c9tHSIHrkQt4bl9yZCAMfMxxX/iE+NjkLMpvAOsC5C0hAX4peHMoFCmszP
YyzRlYJwCs1+xIDtYQb17uOpKFc1DkdX2H57ZoN+ObJJayg0pRihhLllz2970RyLhZbT1uonCafu
4DpfNR26+Re+B5XDv554mvHnwpHaHPlrrcpLgquvRhqCl88ySh8vQyF5SsAUuRrblXL7SF9hZ7Nh
iP7P5qnvsxVHVGguivCuZuDPHmXZk19mnOa9rlvsAjhtH1ONsBAjtZvnC5KIZaINUluonhQBhEV5
UVf9UWuajzEAY7M4s4DHoeVq5z4B11V/uwIE0rSTb3DvehqK37Wj1bn60D3K6bTrFg1QTioieumc
CLs1SPmZPC66kd3B9ICpGK/APzF4D9f53XYjFltv3kgJhLIJKe8r5EUwtxJhZXJ8+9eLgwzJ+IWH
gTrS98kWJBvRoeoAIf2kbXdepoBrD5DU9ua3RCsydT6ncb8AyusGiIBvUHATFI8HGOlGwNgnlFBg
xLHMqexbuNbL7Ce55U7tfJ0ghPG5xeAS5R4XakZ+9GwLH3FrunccAk/FhaTnEg4cLQcBZ1JwsiL7
71vdDNH9h9wRYk9v5XzZ7aKBDLwFF9xdYFUnX6/J7AhJWiJHn1DaHbB2SsYAfC0U1jUTuHLWIWxP
wocAnqZi/NVpeRkHd46Ld749pECEb2NBsNTyb6hGjQYcFUgijk5eF+izNoFtanBh3u24a2IeC78I
pSJ9GVgOCiULTiQuk8EdbrhE0l/MFQ+vnuEeVuH7GQiSGHcfWoOdriyQIzxN0scYn1G41ru0XM1W
+uEFWZZNlJC67OHJ4Xw4tYYhtViDGY07ew7lRPET7+CQsorwdgynVn6UZaDO1wv1tZbuDUYK1vHx
8ub+z4i8JpzP3fAIVQ5VGQxuxd6/en38kGhUkwD+8od7nYXkLnV1vz5SGnsFEQVm1MhUFAcsika4
9850GjHfnzcUJigR9yfXhfhLvf1q2ccVonpOJNJCG29BfTxfXbZEp1ADbBqdU3AL5nXWmdgyw87n
dvLHt034bT2+CLGIVAa5zrI/rvW2nNvNvFVr+YzymZ6XN0KBLysB9Q/6WxYBBvhHjgzI2HZn9Zhl
R7LL6L876n3y3KwZ7Rg95Wdt0A0mp/bcGEwUnz489mJA34hdf4NGc8aJNVZjqGrC7IKQPTQAy7NH
rGhSvIUMhUcu9RrnOZGt+PVUmfaor1G4xr8n5dZv/UQXAp91IwAjuwG/QqZC8dXXrXVXehfCunuQ
WUuIEburJ5Qt0Y/HGa6z0FLbBTRzuNIgMOt/+/k1FWJkzBnnZ00RT/bM9wzAptSMEGKUsv2gx30P
gpM3JmX/UYqMWdnbe6X278WbBwO+CKUj+HCAnrbuI3hU8IrwHCvodLVxrM0sRp5ynzf2OyQAU9Vc
WHdpYtsQB6sPIhCfVmPDee5PJ50GUSSEFnfO86CnoCHjSlgHKlIJ0tNP2y4b7s3QhMtAcBOQ6FVT
LEUVQBC5HI+bijSY5ImS+RiEkc45FGSDU3D4EUpvqaQRMQSilj23kWxznWy+PUSBL5w6b+OYrGFN
D5gw4wj9qCwEj2cIKxYQoFALX4CS88BfnOfACz1NPW0IRDzEL03LnuVH8oR+dvwBC6DN3uOL7GSO
Sz+nsParv3v15BAOgqzto3JqPOuo0jvVVt+uSNDTA2mAEiQtKH50Cs/s6JV8efb3w/lJDQUT21lr
kZ8Sm+vrSr9goi+RAfguOyzh3vSi7NWQuLNEPn57B2rluR6pmzSmX9/vzYsqYKkXs1nzfJcAJGSk
xkNosBr9Wu5hjHM+X6SFk1wZkJiMIacDwgfG6BBirhCcifyfl2w40/Ebja1/AOdhg8P1uOxfkftd
EiYUJktEHLJooMDfQ2B8v11yh0UTAheDxOncTB6UPtIBM1cm4+BIjDFwu6M3bw1zEzkFXsf3U9bA
sSrBLz27gx/XNanMmjol5p8IKhfv1XyD/KQIES8Jn6xvuekxMbLMhFL0fbEVr3W/B18k6kukRlCx
lHQV1QnuxWOyQMk+ZotAmhjd11UWC1Y+hue0J/qys09gxbVhtfDmcIdhFEtSmPzzw45XPcMakEEU
nAZhMdEPyynDQhRpQLG1nMk9QYzcfj6Crpoj5Hf9I+bp5WA5xJkq2sk/oNr86/M4pXs8ZxrOAyZB
ez69tSNXAAA1jofBMwKr/xUU4Z8IAb5AwNlNCNzOft6Ktgmwu8nCNBmTiBpJj+zthKacFdPj+Mp8
ajqUevPgmftYHAkhw21+Zv7FoYm6aqy2hF3UHhaxkrU2IKz2cPIDpX7Fu0K100jsZKarIzM6ydvN
fUg21aWx9Zhw00dqUdY6UwqqTejCe8Z8XKAaIuML0Eke+qlKKE/0z1TF2NoxrzEQ5cVSB9/YzUPv
FZSeOFTCnD90CeduIy/EsQ4rQDCyTKJ0M7VDMIi4tN4GUsVKvgKDAn9vlXzvnkMYzmy74rr1vjhj
s+wDTb6PSQj0P7Jpw/JTXSE/S2aXphyLpxwWo+jwpI5/qmiBlPIMK2IjznqJdA2myTuE/XaMBJPD
zSnLSlcZAPYD+MQrz0xr/y4BMcIwJScUDKzoenmwf9E/cIUnCPZaHrd0mXIXsGtVbmJBseBb8Kcy
jtcBQJg+EbCxMdiiCVNXHQu+IBfWTgIz7rCPCl+52gnG2nl8zT68g+exxWcbd5aE05+K7wZE0ePI
3LdUvimhxZ6tcAPFeRZTZvF1eD7uBhl4rss/ni5cNAWe6mlxAYvlCvm7JQY+oU9GoZU9gj7X2Y/s
GhV49WsfWpLffKQHYbCd6H8dY3Es/FmM5DrWUZT/DIz7tghluFA3/aQrVnJj3pRWMLlzH8g3GtzC
NXPkAGvU3WxgCN01nlvq1FN8yVdWoRp+RZTfpmLL64tK8sl4M+fVp5WEchTl9cTYx85nMMjU5y/k
gj2bhvljeGkomLC1DY3wtBhuU+M2IgNR8IwQhG+DD9yd5ahgY3U9WojiiY0+wHYzS7zaPO54Ocl3
DUzHzaSKu2cTbcMkB+2zgWpxA9AnVzSZ2jse57ygVikiqcFzSnMRVdEJ/ePb3PxFzWrTeJLRmFZC
sLwamFtZXSnZKWJ31FRAkMpFNwO0DHsZBLYWDcA7ZyfitxlelueCafV4XW4IB36pXq3ZpIqjNvkr
eJHwBy9u1jBJ4jB2CXuKEUvHBa6+5N9ZtfusZ4SNEofEB6X4Kd92563ZTgGz4NVkBwHD2NDLiXpD
zLxdNLYLvAklh2RD/kpXWAIYSJxEVYsvtTAzAYLTEB1VzZnz34ni2YMYkWQBlSMy+1sVFBa7qQkO
lC7JTCG78wJY8N25PdQ3MHXlDfZ1HMV2KOlH180pu67UQnIvYvswdC0tCwroslkvTlJPZMY5XJ5p
wHsRTqubmqf6GHY97wFOlmtLfWmqw7zaErHiyj0vYr2mjbWmWAZkw3kcNFceSn145O4mwotYYwDM
ZZ52dVE/JfQytWIKxFp3yFvm8NuiFepcmh/tCPY5JbkbZRgeY/ol68f0IDVrNUTlMImnqZaht40x
jPpcfU8yyAyyA595enz5Udtmn0zyR0GuSkSj8gMkI41iA11i8gcGF7mdNszRNb/A7DiGtZMphgLK
lNUMP4ax5th/FDb+w1oZEGxYbQI6H8q3/BYjsX71zS+YNsn2fVygN0PEGzJiP21QYAysr24baUPR
GJLHLAbyytwTRVd/PlL1fridIwLeocY0u6dzpD+j8JafWY39Ja/pSUabY4Te29Js18x++275M4nC
lcdqyJLn+v+nEB5skx09C/Chx4WCzeU8aZPS94MyRKoXzF15neb/G10loXMUq/69PSDbwuGGSgCR
isKZgZMYRfyiVnO7eZtQk9GG6wCMHi0CzCmuIdgBLDqFjqGaYZ9auaFnm+Mps1SdtgkKWeOe8tmd
V3O+Z4lkIJwgQhnmNY44J996DjUVZZZx00kJVaTD1/ez0dQ4y9JJVWHUxwPh9h7ZHRArHADKOhe3
Lrl72Y+5fK1Z4T+Zao+vqoyxrDSfRaLcd+cY/35o/ZqBddkljcx/tkAYojgpGl/3fB4PfrzNwKVM
KsARlbDb59oMJaVbsEOf/LEPo6h8vV5zTeU0AuUtd4pML4dFe7ZTbtKD3nhQ0yU5gomm5lwh5Cfo
QGEVIGlNCvi2L1aOSjpcPnF7ydaUtTu737muYfRGrKooR92xvPD4c0uabarNrNOkBaz3e9A6Jbaw
7Sch/Ke8gXXI6NAugHsibmkw+Opd67FFFolknP2FlPuAXhzmBAwv+P7GV13n1u1dg/wV8JTdTr88
58gtO2ZV5pW86JxgQtmvJWvlijYxMmcUTl0//bzbYs/ohEOCMEzAIz4SwO++mQfU7dJBD94pL5fn
3f452LBfwxDZSEfbaGiTvFP4psrnDvtoPEMDzNUg4VDGTsC0T4XF46cNgswgZd6JNKi612576WTG
tZNn3WlTAu7c0Vgrce5/wV8o2rB0+IAx8V0794B0hDqr5GvkgA/6bR7wrmCPqDvhGL4KNhQGsmSB
byfdP3tQ8OO8quueM6g54R+jvQVOJ3UfDvc7sU+TcKH9/p3zAkjozlCsdwTCljRHYKXK2Rnbv8ua
FamvueDZD9UE5mmVXnkSJqVzFqByVtXwvrIT9NbuSq8vy8Z0JPufRCDmqkJeuW8TzwQln0BQzxH4
/8aG6Pmp4YxtL9GG43RvBwze0vI2VJKoy4srC804Nedn+viT3HeW1zPZheN4DQuikEYcgrSuyBVL
D8M5JRtU4G+M/FqlyJH7WiN4lT+MmpOKxsWXTdvLzHDIZ+bdze58NHUDcleCb9XuACigz5vYvb6p
Q+jCk86R6LkpR9xW2g1xZqNKhdwZBG94mEd3/kONF1wDcfsMLFOki+BZGG3nH+O/b0aaTp4724pD
dBRsbLhRuWRgQqHTvyKTKo/7LIpPdJcVIuY8oz/diwony58nYf4g33LfMUCZWXcBJSarCOhlhKxy
EUWzrZThzSkYoy7kyUZXXD3JgzKYpNzfLDUuEX3DecIvynNWqBRPwHIa5+9nBo8rehruOOx7alc7
xXW7ipjpk1JL2QUZxKFO9bczYl1lb/JJSPjNRN7Vx9BELOaT6VATiy11sCd8q9lLQG89wyHfSjKN
3qJJbdIy0oxIIm6CUjv4bsco/1Triu1LXgos5AKvP5fQ5zaPxqqbOxigEhsp0byiRnBrJClzB+pm
dzQEnkq/S5POQXffYAMA3hXsYk52C27L/5VkWVbe6Y/oOKoVtDTOIVZWDwpkzU8brQgZxYJ8LIs7
bVFht/kamGAiWyknySb27a0CNa57CG15B2/F0NTPiab5whuKjcBz6PTyZ6nlwzw+oYKD3AYYVpud
hAwWSJvrqnNCZvUgSJbFW/t0Pjc7lCq5JnYmQpgU3pRczWKIJodzl+l16uxUsYGdRDPMxhhoyeiz
hzTg3wu0GJRFdpzbW+eaK6CCXvjYu73SRgkjfCsAtFLtS66YkGaW+LXNCC1yDSJUU+NplN7z5kPG
2/B2xAivrOVd2eZ0ZfM0X9iGzPMdgYqdLGdwfOFRkg2TypFKJ5Wow2w1kbLk7ml47MwWZeoS2nT4
ptf/on8K5jP4NfNOwHcXNpbmGuI+Fci12amqvL9gHuWPJvMVCnPqiHceyFkRPN5yYhlScRTbt21n
lXaFgWaHP6GM//vvrW7nsUKC3ipjBaLuRik3tDYVjqSoLOc1oPrHl1PUUZYx0yV3ZMCh+1yQWKUY
/EMvMaMBkpI0XYWL/VEeGg1Ew7HbRDZIcopY/+49Ct9xZNVmErgLlYcajSbyWUl7MaJMr9h7fCtm
6E9MX6+XrRes3sgj0PxlOZR0CCf2c7GZcvhuoKFKE+chAl7a89sJTAGdM/ewKHXxOf9jw6JmlozO
HIHZ7KCN6hfercCHDSMKi5tWSXq9OW2FNhb7xEBCBs8Oc/3Phfc1YdTZ5JuWZQfeRG7R1oKro68e
6YAbMGcfgUjy6GqBnqJOvxC/7eqqAEOpVpbSXLgyVvcb601ukk+8RyY2vuBUGraR5JAZ1LOf2GkI
qpmxWazDoMa2mhPCHQ+3zBaTHJiqgpxOjXUjDD3viYHeYaxn2WxJxrk7vM4fc7WsA3ECmJr7etn1
tXf8zIQKvtGvCMSUmXBGkthPH4hf5kj2WvUBu7BEjY8JbhDxl3r33tzdMyOCXTrpOFlPhp9d9Vjj
iDTR8E2QkIlNI73iT99x90LsmrKjfaqLeGTKA4m0YhNUE2aTDptuYPjOXmwjIxXbGAt/9xbkHRUC
4PIgo73tLvgzbQ7nHUnr5yuMxKoLZUTHdzKdH6q83Tuv++VqGjYrWI3G+7d9K+ApRnOKtpvyRMn7
Eus8Rch/vKOG3CQ8WqwqprV/V+DgqurPHM4IQvqBac0wrHFshGElNjqN+P+T1jl3wtrjfMfSfd1E
nRM/N3/lW1YM7Mm7+sbcraqNyClO+/7H5LG13wgxjw6GYVN0qUWVsjINh+JRH3wwvMuRcWFZ1VJD
98MMo4P2a0GgYjf/+Zv7JDo0NIliao0OeC7v77ZbfrQxw8otN77XG2to3IXTNMpSdBvPgJE9u/EY
EqvL5DFvQPrQWi38SYwbABUhHevTzCPV8TraISc3ltBRxUhLuudRJoIs4Ix9eajpPfB+XoLfYJlw
zyxi+J0syus6+1VgVrv1+erCQEFrTxVDZlCrKHREENtI1LrJuh9B6w2m3anZxTqi1TN4Mj2RsDWY
PG/qPJVXBq0LGmf2MSk0fwF8HZUayMo9PBqScOM+UKma2GvNusqiN2JQPL4HSoDALd2TKRsKlWST
/Ak5vPygoQRiqpOxUKt6MhOtNrJfWbkwCa4zkdasRH5VS5OtSB8+l+1dNVMLCH+g/dxx5q10ym/2
BO5mOXg+fvar7ucSJb+aJJuZtQwxGMEMQF+jUrLoTVtvcF1q8uZKcUG554zpn/R3vbTEWO7aFFGh
dY14NJ2E6kZC5y/wShrjFNlYhwFjPcZNn12Kr+23AT+3xiimLiwo7t8zcY4xzsi0VcSl3Yt+hTMa
+wb6Ne2J4i7eYMGRWjE7tPBo0zknQnLIDO1PQKY8om9yhUAprFYhCh3Vw88cUusZS8Yxs1dKOlhT
aD7w6GvOOfK8A5R/ETEoWIHGAu5Ds81G6eKxAN1IcWjZMJIdhE3fRRxBk78i6iOpcwUcRZtg6dwP
ZUE/SXo6T0Kqb+MTaAAm1YiazNxUDQGM6SV1nUNFYg/3RHYzqPtpBxMHY/2hIOOpbIqtovMER4pz
0RKyxZP5w7mfktqz1v3WNtuF6jwhjHsWZe/lyAGf8KeCczR4kXej4Iw/5kx5cbYvdbBArY6fTEFH
f8dtgYJcoH5I8djfbCkRWQmm+j1s/9b508VGquI5Zlt1pbgGPhaVs3QVuoRxpDeRCi5tC1JtzHxs
nEzY2ahUGFxDyCA7VGPNJFv71wuQHr1bmZ7LMAmJ6E6TWoCoAAYWg+qNgvuT66aj3VKTAwa4zOCG
wvFLul3pbbY/rnP6RcakKZqPNtZo0wQMbsDggfKa+XtxYmnHk5Nn2lgAGs9IYoPI3N4MO1/Lk1XG
XABmE1A9ej3+HjliqQAdS1986bPgRflRuozAr1TBxbIDwwTD7tUQQqkbS3awfHLG5v5V+AkfygMd
pUa6NWwQ+FsX+LVrsV/OhWaB4Jdfg1DedupnF8EjRmiL6C55MVDtcw6UM8BpJr10cMs+p2msuSlk
VtJrMr2rWWfz3KIl+zwHetgm/qE6U/tDqa2CimN4lL3lpZHNO8j0p88LPy22iWjQ01JdCENJFT3y
UiMh3KcN6hwfrR5uOXaGIGnBt1liDweNXFVQgV5n5Lf208kTNnS+hrIz24aRc4tyBgx2aSyzmmDG
VaBW+ydKwPdU301Z6G+RsZIKp4Zk1YzUa20ZQfWuuAiaDrIYb3J473ggFzXQG1wVVFXZS29KI45i
+ZE/NoGiM32zOSuYE1TKec1WGHvOcM53dK3tbgGMK/SjJSMLYWEl/wZOEEQrqim1hADzKfOUYQqO
0NzHew24YdAyz2rfUKQCwd9NLm5vXHcfNWvjUgAb+H10eDiveKXhNuV6Z82Ka6lpmz2dOMccC6GS
oXHvM2dYO76XLu5jbhztxvODc/NtooS8lQwZXsg89RRReZl0b1SHQn7p4sST8zJqZX6VOoy4mM2H
vHWzQhAv+vbS+n6GbTz/8ibnhf+YK8CaldBztWpY9RfamVgHHMYQ2OGd5d9sRmsgvZ1fhO1d041E
1C9ms5UVsZyY8/TUKOra0H21NfGr8p5f5E0AtKtuX4UPAtyamr1ulJntBCpX8S+s/nf4u0e3EraM
JT4LGBiOmF9soz9FNOobMWVfyZ8AqPVi5SyJxQ9f4UWxLtw4HEs6Unt44oq3L/TcXbYAg022wWKc
+NSwH+1tD8/Bm+sfVNtgYg+vvY/sTvvW8MVSH8e5UoQEPSDr5csDmsynOMbRSVpLaXf1mYbfqJ96
KQtyPR9Jiay72K53fyia+b04cRQsW2lF+vktJQny+KVGD7pI/p/MU3Ovek57u6oOasE/4IoXnggk
wCUq72MwJq0LAw3Cp2dJ+6j9kufrqzGcDy4w3OcnBUO/vF0Q8WnsQGRyICTWbfK/EkdZ+QvlOL1+
E2f9dGTRBaZxUDIOTXIUeh7XrFdEsmlxO7YsvdDaw9NHlocdvfUgaHZus86Q7HAEkUotoAkWJbYe
Ik0r3WRK3Q1UMZk/qlBXTvWieEH1vZTJFtqlbdIJUt3aqhdtWLUAi7z6yC2pELx3sbDKiyggGw14
59Hc6vlYyy3Wq+u0BGVZVFVnMVd8bFhmXqYICcXakIUU9Q6Cff4FPxVSsBpHIDQJ9g7vDjyaOLm2
hKl+Lxmo9n3HC55EnPs2JOSWgzXB+GE7Cl3/IXS4eoxmNUc8ky7iHkknwG4aBvvME74HjMzrEC73
ZNLqW2fyVDLai2rmuw0ZWMDXJ442z0V5t2Ob5bsBtzJR9S+JWi1g1D1+07nb/V2/hBD+58ggLbOo
LcFrhdfd5eUF54uvDaOn65JKMhC8QjKC8oO+Yya7+dX5Nk6QCfMpvxC6oZXK03npUthe6l2xalKD
nPFHKdpKY2oKRIPMBpPjeEhV4qjf42JX2JBvPI9OWip/TahLTbMpE7lUnTLbOMUfRdDb0s9P0MbD
feRGu8tyaoezluq6L3pTI5wRIARt91qV38zrTCreF5rsypAMOy6CviXIDyt8xHXT+/PFWPFhKNY5
JP1VKWrVZAfWvGlskYRqW1Wj7iOMulZ5c8D/heGXrKxIgt9jLHRxj6NIRWVFalPjrUFlzc9xMWQb
4gF58SIyCsIUbfVLIvnk0zCyLaYSY+TzFSaJJmXV+XbdtQxAbH6ox255N65I2S6WzrY1YfSnf/N8
nAn9mWcDJlYckTbwzKsB7rEUa/1XrZHyx50Ab4rVPzGhaz8fwxTyxrGnyE/LCt9T9gbj6mO01aYz
P+7oRZ3eWWuHTJTNTSQrrTp2o1mrNKWUhagljwPQnq5JzKJdSE1MTGRQpOr8YZQQGRyG3EJ79DR4
8JDrB8shOWqV/ha3XaZvlGVoU2xY/+QG2wq/GJgPQSyq5oszyq1NmlcYnAYudEDpV8vBbhqOAmEf
ZMvIco/FQjILqgcN7fcILgrjEYUARMZkpkG2VjqEaokbaKD1HhK6BwIlLCIQ66/8xao/KkAUtedF
c49vO/aEBFzf2RqVL4Ik5b19dPljGJeX9T6zW5IJxWQwmAdvCj4jh9KPT5Qh9yzfJSO1QNNhGl2d
0RLzn8h89KDXub7vD58ccknJjcwx/lM3w+dofkJIexaDSLAS+/xRxFLY4Qt51eqTovcNmWdjm7xR
kXx4W3pZANxjJSm/WPh6d06zbG1AJtMsTYsMw6OSR/2Rm6h9oX2VRLqrTboWQqyqGUxyv2PwsYpd
24C793u7ch5K2Oetty5uTKVt2xf4frGM7In325raOFCU5OAvyZbW+G7ziBBhJKkIRiEMLQi8IsIz
B6DVsiht2QtKBx7m480aFqTpogDT65t1le+sfl420IZSsjAt38NBR68fcHAqAluwo/LULJbG/4gP
PBxfbWHR9iFpEGa9cABLHeQbCPHlb2NIT527UHP1caj2dqluHFtoYVjzku+IeUpkJxqBoPoCge/1
tbBUgGLd3X+SNKNlQaRoWvvbBRTbEc5RQrMesoY/KG+19Hda7mT0WM9A51A4SidufCDLZo7FnjNI
XUEX3ny3i5KFCHHA04VcMl1cQzY875bUw/2ellRn3sufubmdA9nwHOJLHlIpYzwVwxEAlazwGCeX
tM2/BWJ2LsVTl31uhw+97SFbKvIB4H1jVpwl6xGxVvGbD5/p9jH5yiSZKbX4gRNMbhhyzBNfdech
dOQzwg9GXmCokHMxM0DYoucySyWcNxj/uE4Jfo48CLi4Gln3Bqzovovlk7+4eWmcwJD6iJNsXesj
rJDP3BDlIw4ADU+h+DmNIKm6FXvJlC0V36BaGLkz2yYcqGUFu0vyBJ7l2657haKGPEYbK1xylHpL
QBxRIIabqGqbaOhBJtHMoOpWa0CA8HvZLr4lRgObUs8YAW1zOcFQk5hIj6Nk27PTPlFa5B9Kmrge
+wyPbf/MMD1hUmWbEt91skI0JgvEldI6DVTlNXwd2UWs7+TRgbM5lMhcZcA3j3Mjia2hVQh+8/2C
ntErAxOvKeKAsWpo+KVf1YALpvsUknuRCa/eGSEw/l/CeVW5TkZRlHVAMmcCT/nMtseRRxdJImyC
QeJatmamCIQisWKicSpbfLAXbfFb5Pg+3bsvOjCSBRZl3oxUH935Mjs1YDB6ojGv2/+tbVHCFnrV
KKEQ6J0PodeB6FnTJlDrTZKrrOa6/YVGIFRE1mMO5B3tSN1va0MUTPhvda1jP8LlBLzhLFzFjIY1
kZLYln+YqH4PXslXAEEwvPaqFCqr9bJiTU3DX5cR7AJvGPB8Hw+0uZvemyBqKf5ogHVAv64ghzYk
6PXLk6yBlqIFxo2GwrwFOeRQ5h2a8/3qfAq8WTlmPV6/y/WS+e/XdawDlVcC8j0kDEz/kvbML5iM
ADEN6khD1SwMHsS9aBAvXY5SRQgKJur3vwS2Y8z5vb5Km3YtzXy8fGkGiC8HcA6a6CzKft/uIfD+
/67VL07jSxqEF8VwG1+2CQVS+wsOA5HP3u+wWzIW95hPyV3b1Q+LxYmgMD3Q4AemmXKYX5HaLch/
xdyfut/dVfV+OA31wV766LjnxScSFBOemBh8hTROSbYIg4QsfzW6LwjQ973fj8oH9tUiizvJ9pyj
JRvItdBN6DYbtlnb3rsL4BBo0d1MCR17V+h6ChgG2y690dxwKoEBMB4K8GBxnqEaoFO4XywAmR8z
0b31QWIGdQocTNidWhQIzjPVTQWUd6COTEXtJqkU6XE/GdUzJSyDriD/gJ/PV+WIDoWNIk30xFkd
8ZAKzhmQCLROAYAClj83LozpLqsOXHLFxdGQoE1KmP1+IUZodhBjorYN9sIZ9LaWFjm9dT4+9ZD4
dSTo6WjoG2JlWf3bVAhb+CxVnYEL58SAscutidPZLN7efMauJC0sIwfE/onpzMp42wV9157zqnOx
3ghTeyZq9K3USjRLMCksrqzb/3o1O2uvYkq5FoNmWBW4J2w/YEbr4i4mYmI5o/hL++T/uhfLg323
6Vv2IwG4sn3q1af8Eqpc26TGLOGbjlUoNDtxX2NKK1EBgJ3I4Km6jie+apyqVPesCt7IXHI2/8BV
UrsCyezn5qyp+hvKiolTCkjtIkASHqzr2I7CNhcDE3YZMJ9SReunlqGZicCaaQPgk5Wbx5J6e67R
8yIgIkzkYMzcCLC0TrVttuyLkaXk4+u6c+V+3RR/YGzIOZNIrsPznL3vfjqzHAAdB1bP9rhrIr+a
AiyPAD1UjzVhbPDMWxYgdSYLIe4UA0Z3NMwmL0TxYsA5Bn092/Gm9HYxJracwhbm39JOKsT6vCHS
wBYMtEqSF5IpwWTldV8z27yVl8nsx9geKO4+Jn5hHbpgSZUcQ41N5NSw2qPVv/Vdfm1inkQxoD2l
CmT06CVJG+L7PMxhZcEM3LNP6iOyS8SaJFYxPSAR4c/1Uo4e/0QH0VHObf0HCIHcy1IXIUdt2c2N
QHrQ+r1Zt922ZBbhE60P6kAbQmY9iQmbQ2SlIJexaexNjG+dATRvEZevK9vrFXCGf+921neGX/P+
UubL/xwohwy2/oZkZwIJzjeWBEKyL+Q5Whtutz/4pB9xjFvBaoKhzPaO0vmzHIET31vaD0rYtO+a
QbjZCq6rTzLsEsCgaRGHMRzSWjVmioSJgmxCK/RZtrgSfIQKLcbaaDRlcg2QbtT0NBToX/kJZqcB
/0BsZf6YAz/ripcErC1oh83XiMU2NLXKjBViT4oUGxjU61N/m+JtbLnMks8LWyc2j6zba1hHlDJX
1GmeYanzvIBgGf2co2OiUviXHGsoA3QgkbjOKAC0zcvZhFL4uv8ipPV1QLrZVmS0QWc+nTPLPYyZ
a9P8/VgNed83TwGKAs1gYHhVzmo1j6bLoCARsFowCcl3fInhFFVE9i3Az3Sa08viamEoIt0pI8zT
8O7sFJO4L9K24IOYlsUXHpVkeUPUi11PJfl0QQ2gtQorNl26c0ml1OVVrEwLMYvd6uedo6fwZMsz
GrDs4yxRLxc3pt47DuLN77H5y3vfdi4EHY/VVs8kTiPoO1Meb+W+V8VbVUTG9i3B7QUfINpGYICI
lgBSgO/BPU1lX2uOuhwkMgjEQ+rS21hoILgKx8f2LLd/JUbVdhkwqe7Jgh1ljXje6zErRksSoQzT
DAbCk0djmKhVPtICpNAIwVQGSyP43eAUBdANd7ba0pEGoYSOAmidi9jL689UYuULS+PKu4Xv/Ek1
ZX4eiESW2EWDNom1jjLMLytxtALZ0UPxffIiwv5BHJLfV8XiPpoB7Ui+m4BQY87A4H4Sq/6o7/o0
4AZy79Gs0y7S/rrMTuZpmvBibNuS3nL7RhHcNVf0MGoNqYqQBYsq6smcwiyrXwcRTTrVrsEjn1Jo
jH92Z6UcQktREFgg7392LaQVQZnt//oLU1J+ylXqfJbi5p8n7w07nZVvmSWqCP1CLbAVk+A3vlGn
HNcRpKBZzLXoiBJyf5WR+jrqtjTRFyS9In2jFuw552OVnFHzEoAlRIS+CAk19QMXQfZvAt35pm4j
G7U/YHqFeVQCuY8Yqpdsjijd2stPMDlaqmdS7H13qQLEF0b2EVeD+v73B5TwNbUh95Zn4aouoSFm
5Ok29mfdhlpIfou/PXDRohny8vW38VymC7xswRgRMMBEWtoFy6O+nclcCE+rA5gzOdNVK0OB3iNb
UF5/yolQLwB8tKFn4HrInScofnzOQVpJ/Gq6AUHFbKubGjKdDLa2/g6OGWcMnCLKYMO9CkjDctv5
hmklDspAuIFfJ4GMbuywkNR2V0oHH5uypBqEBL1V6cHgfwzCNXldkxxMQHeaXg6U00YdSo4+DCO0
azszcjMrgw85TYUWI/dPysgG0elRSnuSAmMFqszTI7+rpvq12NOfnLx5u0Ix3lDML+yYz+s4vZrW
5i/Z5uIDQ5/itQf6HUOhK+k/Fulz5QNP1XEzZmulw4Zl0n6vj4p+b+FeqboVsx0UlSlPtm5Cfg7l
eYTJUFO2QJz4mnyrFdFe9Ogiv0X9YOXvKVXR3UXBqBOKX6vsgL3xZOF5YVxAvHnOhKlrfi38WSbM
m7tHQs4ytYCmgaYoGRNYvsCVLnnYrL24oLAh/vkULoVdQVAOS8MOtcABl9PQnIF/6+cwsEjwUElW
rNvquz6TtE/8/A6G3Q7y19ZKCVQE89FldwqUvj4OAYbanBspHYRA9IajZj48m7m6otcu7rnhOEG9
Ymh6j3jmxxZgilxEYdejN6wmYUHEuYCGtyF/mPVOzasMzfdVVgHU5yC30FfUj45PXnU9zLIxCr/g
6W60Fn04qjp0q+tlGHt+8DrKeRfCqeNbtZZmlA9X8kRm+9l/kTA+ZM4BWA8PaHe29ctGv3bAruj/
u04cfBzlz0m9sBlK18ondvxEKljjA4j8n8l3RAeplI1GxThnpZ9kzFzTGBFmIK16JPk3RJ5FwpPs
nw8ZFmlmCig7NK7mb2dexrcKFzxlX20mf4zMQT6TJheNGV8bAJIbwHay9poFPSIiBPHbLD74lK17
mDAHIbrpoa89pYWXEzq2NB/KTZwp0OOgvLbU4ShpyZLYWH7TlUaEEja2s6IAI1ymHKN7sV7Zi0xt
GySI6KMtWbqmZI3wfzSf6oW5T8SFe6g0KdjJK9kh3sfOWv8x/4h5dS5tA5tjDKTArUd+Uhe/plPu
cwLaslvvKYD9ZUWsZaEBIvApd2dEWVkqWwjacwdXITHkOMERptE+5BxxIQvJvCe1gWAGP0pfcKsN
YaEjlnNg6V/f0EY9933UVZKI4YFtKR0ElazvnEBtXW+0vLx4TPS+qDEne9+vPmHxU2oyImPnj9PF
rZh8EeH6NyDW4p+UzpWgjhw8ryZC+Aat2mIj9tLeML+1hX2ORI5h+xvDESl7yi8cVRIBgrf53u/a
qQHH/2V4olQG1H8wVCofZkAXdazWU2CeiAwusSRWEtkfZiMTeT2zIYD1G4rK9ZcM2YgSOGXwKYxV
WlTSFVMYbvNdtnkUK6GSQPyVKw7s9yWlh8kp838EmXWfgdF9XGgq2EUeP/EcznsYUJiZoEt/1Lun
D58kHh8HeDcf91MfNKTZwvgmJzw1h+JVLLhajXLIVlKrbULn7vlVPAdWDyPV9DAmXZa28iysoJCj
yod+zZnWHAVby9iqJUaGFKVuNPbQqK9M6O7WZi3b3aFrCAub8r2rdC2TXy8OGzIY4ZXxd+d8MmEr
Ke6rcNA+4T8s5qt90ueoMXBxHDGMdqhKzufeFBq6YkRyJb9FPIWygxnF5hyZ3FGa0DmAmucfPQI9
MgqglY4Rclia/G4A7Q24NQzm1WTTzcMy0jk/REoK2VDk+RrrASDYWGJ2vTwEPxSZcH/Ha+rsh8a8
jqHF6lMaI75pE/trknEvrm9g3uu76dtB4PpigN3mru8rwrV7xcBzKDdOZ4KhZxruxE/tEN2ywJ8o
IFYG8uIJcSbdnp0NWW8Xi4HQORdqQyg8B28DuTFrN+Z10WvDWi9Zr+zQs/mtt+NGzQA9NG1lD79N
v0m1vGG38XbxVaMVo++7eUXWIXBDZvj18g/uELmyFlL+Q8/jrRynn40hQeOq40Qkc07Pl6bKXa7D
gd4kkBEwZ1lt+TzIHvyEBn739Qv4gb2Vf+x+NpuQHngdprgWGMYml98Mv+kGHv7Xy1uG7maZ7cwz
WHJK4FyZ3GuwTpghHb5/xCo+hBlyO+/WkDAm3jMjsKfBq7xW0Y0lHWVwrYcQkXOEbyrnZFOSdeSM
kjGEu0CAkhYGWgZ54tpW7KNV1lFGC7KT+cAPAdQLNKw8rYFPXXGPGB8SoDHjuJBKbOHK8q6pDeBo
xdLshMHjLF4q85FL7b0+kUytcdfN7xOqZR7LTPhwxobSSZ2rDV37zIMgmX4C0exXmYWyvYmhCYwD
7FKG8YAal6O4zO430aNWhbhxP1q8CIJ6Hq724KsZ4PCrumQnSRrh+V/z+9yFp7cuuNYWNn/rz/ex
/+3pyVsNwwNYorwu4Qq0lndMxkQ91w4TEoH+ZPmfpwnNVpcRsqyCF4NTtZmD7l+NoByNutcxRkNA
dvBSD7xF9i8qbC33wmo29PCUa1fvGbQujvcAWCzJgdsCyXCf/rgFB+0TjiL5p91u7bhoCd0Uuw3K
sjTQigoyIs7YQo7IQF7cD98R1eFjBymz/3aFOlzfWnmkbSAmhKtTLFMkc3elY9gnRRJYfpw6yGxP
g8Uzl454TsWqPFISItVcLCaBBBKWQKoLKQJUOeAs5vkaXiynEucCGC4R0kf5IKTphcgOnOvcWzsC
5QFX1wRq7+F3cPUg/tTodlfbYfThYlehPyKemQKdtzWX2toAuCXWtUAXvlUVHTKEQkbTjtEQz+fx
fO8Ksrzm9m9iRloYC72URdt6g3bfGxY/YCXw8s/I87soMUZ+ofeZtPJrBjA4E/gkcm9F89739pDj
X1irj092aoBKmXH/pwxWz9YDMnOOv4u8f6xCXkSjCxYB+ihf2vn5cQQTeQ7Hxr32JTaGH1g8ynwD
8cb0bW/J4J+Jx90O1XhQJpFCLo4V8vQ9DaxH7SmNxxjFJyLORPYjvr+58jlAba8YiuZtYVostdMh
70hHF/lU7+FYTKBAbaykjWY2rU6Y8XjCOzvwswIyEiO/amLbYNDA+/4YxyiFN4N14kwIR21eRtnj
3T73SSzJrKrWqPzO6m4+IX9SdBvKIQpJKlhY9u7eb5soTqlL6/cENXdPcY+7Uvb09wviijslP92n
1wZdIJj8EZYVqaq5jJnCqjcT7Gw1Vbqa/zL72TzJ/O+rXKhUw64B66VB52T6FnIU/Nh0t0gvRSIP
HZFAXkFLMWxXa677kmjhT9L0mZ26rvkWDpUvTbRJfD4fA2HmVoVCjiKwSeo+OsPI5VfEICxLzenx
IJFXV6658zxcClMS78pJUqGmKcnJMdRTKfAagOgooRL7yidDyaZR2bonRgK26bQ3Lc4xuTwpTuU4
5lXWcKboD2/bHV9ooy7KVogym5wnbpLW2MVz8rdPa4imu0T0nqU5C+mxXMKmpjzEQvNJN4Z9PM0x
fjumVwDyc7E2WdXOfr9XJNsQ+w85Rop9nNyWpAHawFA5gh5NZlRJnJeoinYk8zcJVvIu2Ca6/b8q
lASJwoCxrCURUOZQ3LDsZMnHqQ6cYI9t7oION0bkwyyPXkG2Uh0pKxLRD9vJe8rKfi9vO/qtwIyo
dXblruAzS9mmFONPhPluWtbDbZR1ocQ+Octg1X5KV1nXAjN2vpuCZ+GX3Bp2KIE3Huz2aAg/HOmW
f/0zbPyLI8IJUoStgsWGZz1OGRgXnzOeZSvnsIs1Jzw48VKziriqlZzcIoCfFYzn4meGr05mf/LO
Ddi+SoBkszVLPhkBBN1hf8Zzx5oMqVY1lhPekDxWhbMdrpqIxvTV21Fu0AJCAP2a298MxogNe77N
R4r5rfc1sSZdZbiyTcQS5JU9ohk+eksmQAzGzqCuAChE0lVZLFeimETTeuF1aiEumucimYbt0CDJ
MPdzhZBYU+uCDGdxKdg6rPQZMNOETcR/CWKh9js5pCu5ofoV/zT2q+WQad41rl0rLv5jHg2BOrXQ
dBb356k3VlsJVmYW5JJZsbFEe5/h+vMxtmZ4F+HLkT0Epapwfc8Pa8NzUhBiXpjiIjfDKewRwgLS
DdwF26YZ3fZL8VxhnDJsnmeUNAVNbOOKypEKCfZiYglDpi4CcIH8RveaQC3xkOesOA6bT6tN9izw
QAwdHuFeCTGXf+O5d60JfoG7Fo9vIe/o/MKiBYrjvt6UATrFngdngxDTAlIDoM5vRUMfBhuv54ki
84penA1ai6SY15QwRS00cClmEWzCI7Gzf6R91mc/hUpTAP9C8Jc7IdipX5KCja05dWpSEpUcuFlt
ntsXRGIXLbBri4uDLRorTYaF7EJ29OqxuWoMhVQAGSnebrlNMg5OOdxjPKC+usSrnB5KnVMD+RnJ
s175J6E9z0kqVp+lDfJElwuRgfF7z8TfeI+CDQgdWbI2yIYa35myEOveI4CzsEAUGMlYBtGj/Bnu
Qzaloih+vL26S4s7pyg9Njq4OI8wp4sRn2dtOqHEb8q6YKz5n/0WKXyFN8OPl4Rn9TN8wBiwmxyg
PpG3HdlPuzSMEwKDWF0kle8YK940aIYG0BekoZCVbH3v/vpFERyhGqYKgJcPW2eMow45wr1X9VdJ
mq0kgnt2mNUDpw7mQHNjB9PLjBEv77M0Rq3/Z6Ld7pgNG5FT/6Ar5qtMfRF36HJqA40ZsjVh2J/R
ZMItbZCd5hj16nAi6HWSIxGnHhnu9ZsnbyD3TOwyG+bgYEB3r3LNX+3jE8ILwCbJ/uK5Sy2JGtG5
pyZmTw7c+ck0NgqbjS2ONevujHxmovmdPTRyzA0O9eVB5qv2xv5t/X9GNqZtAYr1DnRe2p8UtHQV
hDcdeqpcwxOpPmwBT2aCfOLtRUmitFE3s0wdwFeY7BFSCK4i7g0uw4gsuumfM4AumxswQG0YeWDR
q3vmosSIhh7fQUtbtZIKsPJ1Wr0yTEBzYMheyi9ABafdYjvm6XVYJvNIAEjLCONGZyXTe8ymz0vO
tzS0OFe4/+da4lOmUKLJbnNDRZ75aAFn/fFS3RuVNYW1fDUIWXV77TwRW2whsVejD7JR8rxsW/lM
ER/C7M3J1U24dlteRzv2oDGPRzF2Clu0Y4736RBaathWhhYF5rcg/b+SPjLN2bFx46HXgIxXyPsg
xJYxscvzdwfbGoKLRzC3JTahqfhw7i9Pyw2ToAjyo0c9cwW5DwjlEt5oWkmcyzHr5pte1Tn+klMj
GU894NIYS3i9C8oiCGHpaXXQs6V0cqEo0AR3cByAUyEAVGx7uJXkIJWaP1/Kpnl5mMClS0e//1Jx
O98V8mlRsSlg4EXYJSVWvoki4NrYyNdWdimOhECxlB3Y0rmVbZEFrrvKOnRUH/tX807pdWWoR1QO
njeApAEMOfQiYCxHYhAO8utyJ0wFB7JGeTgrxYEkW0uVxIcKJCR+uS39K4A6q4AdrYOqUnlAlsDS
AgwFwgWIi060U1KTJx2tSvTShXvWY9n8wnxNDKCkAu0FUTLM8FPWIYqaIB5napg4a1NIIkfyB5A9
biufh4Fl5UgUxeb1UYft6F6xTMaT3kapGNVpAuf7WixyGk7w5KNBnYn5ulGsj9KjSMAmJdJSwN4C
A7bjQJPXxsVv8Jwguvwwe0zDl3bm5Q8Qpbg2gzk20Wyg36QG+IWoOdcHD0TJIp5rO4Bw52MhBwUc
zTc3o7byeX5XU9Yz01AVAvw0j067NjuG9Mqp6MMSOWBWdiszj7D1YqtEpsYEFM/rWJhTEQcdwJU0
b6RyCXaQ3NNPZQdcRAGIG59VPSiWUTqpDsL1nzA2eZ3A0ghRKf1WJleD2BUWrFuosR2jJLFbCAla
SEKvmDD5w6yq3naXMn0h8luXocOTh/0RFRZakqDiwGbts3/iolP5DpkXtinPKGZtkBZLNo+82D2Q
zrdgkwbGZvg5aAA1Z4Dv9wEw8HLNzZtXtnEZ/wEZMhEA39jBli92GAX8wsXXWXKyV5bu5hHZi3dN
IY5A39XDYzadpYcR9fDFoxipmM9weF0K8967IIo9e9p3mmO4htC4mrCpiCPJwdo+p23c+QzfQqgQ
mWOvqxFtjU9qkMkh/odaIH0rcCYIhTorI/OV8HvQ1vcSsgFOIPTwVGEctoh/av+vOXGMJUfxzXSy
hNkQXwIo0CN1h/8DBvyRxEPXhRoZE2pucZXsK1Je8KHTbt1ZhEaxtHx4Ua45y4vFpnqeRaWdCcHQ
G6BLHUNQsB4o2Gel119x1OnOdiLnsBnz5mmwm0SM/V+XTSjMev/vCwS8pxxpgO6UwQhP8UdDd2IX
NHqro88SdnJV2Xnj25CHcwvTDFmn6BZScIMJdYk7+Vml0rzG0HMDsZmgdQRn6iuZphM0KxRpcvFR
SgbQLENJHPVuZ/TIqqZMbLqle/t6km62G7i1ej63gDmH7oeFtE/g2ROdhC+QdkXNj3//MEjzxC0e
V9KIR2fpQI921eHPxjg+QjGU9w3ohiUwW2IBF9CW3Z90XlGiAEWKSvknd3sMoRTqPcR6ahULXLUV
fmz5Lp7AEEEmyBxpcDsCUbb6Ze9RydIhRn5FLg6px2JayhNSRHtHBTnYKVU7dE2QKWzj8b1Ivgnz
NpIaNkuev0B4JmkjAfdSttO3Rri+LB+sLofmTVDArOH8GfkFSOyCgvoUcPkCSHkFWFx0HhFBAQCm
o8k5gyXW4tMPzyYn3iT0IRLBI2BhkWAllv/rvCz1+UAnG1YCCoTUlhj8MoCI64Z4VLrziyKEn4sj
Mkj6ERn7u915pYXA+v2MEhYHc2qsZbXvTYuPS4zKBxo7SS1jomrbYKa/Ogt+Br1DXvwzfFF3VZux
V/HPFDGzcgy3Dd8yX4ftN1mHSrZJXMliWTESUZSBxL1JBjmlKMpvrsZscrL7G6+XYOGeqtMqdAlM
vQYce18qOhKW4rkgnaaNvnKF9zmZozH6Xwd47znLqOrPnznzSZpFQvMHITTxiUIDCk0oqzjPqzW3
LUxH3I3OGbd6iKshpx6xlvKoJfJ2QhW+gIdu6mTQeEfItJdah+auNcXVcj/mS3GipWm5r2oOiKXc
FAaMCb9Nwt+2SkW8AuLYhlQNRI1tsulfjP/Y6wY8lHDGYoek1nmEbBVsLJURBNllEC5koBojKlnw
L8XdXUp88D+KhXuYBqJ676PxZxzDWiLS0DLVQvQKdq52EaRva5CtJ2TOmtihkdI9EVfYaavzzKrS
9D6iOEyzNc6tbKe5s8C1OtwrLmPGp6atuCzM2rmHEi+EMlMH08U7+BfGVfL9eAAJfOQFKsnlJkYQ
eeaok6R3RmvPzO74lZcDdxXteoLMD4dkm82GLKM6nSQ4lrOAe+2CcPyR6KpM5RESrVo4/VRLGNTL
bxA12Hp+JKGYEmBO4gTtlFLG61TF50AhMr/j2eUJw03OFFXVX+K1jvxTHPYUPSCGH8FRY4SAAx7p
YoO8zVdZGKtYz5LsXCJG0SPokXAie+6WvhnQ+lqCQhnGa18dBrR+L94IPVT+Xo1/tnBvhto0W78W
L/b50pbyWbE9LzzbchdigglhFriZ1Tsv0P3wNizTxfGeZXjc0oR/oi6EAz1tUhW8kozMZrU9mqT/
DuYLj8/O9PCs2H2gfH9pSWGmbBTcxSrUyWXcgV1WLKIA9xJ3Y4D6CYmJDMftLjt8qZdj53TK8lM9
KR6AG+bAylQAhrBZz6LijEagpn7oz2qrTWhpqHT1clM7jRuXyA69ktK3o9xZ+S0aKIonldoBiSFy
/CD8ulqbW/H4PBPUlzR6OLtOjKoNBHMdUsUNWqF6ZdxNeWw9DbaF0dChSC+nPNiDabrbBRJhDeZN
HVhH8Etjh8M9eEapPSl3LK5P4PXE3WY3dqPC61ZvSrJChpfW4eh1q4XfGl2xhcMOyfRh84nJuPtr
fVplxtdZlsvcc1TJAU0WtYNCOwF+LVp1B4Pyfzxr81f0gNUCOZeTYofwAAA9s9RoXI7u57Cr0EUS
V5/S4JOFXCFjnPD5bMonugp4bft0r1hY3UDy9CdMU2iEj88DGfqSipXx+dSh1f/ylW7evHHUVK0C
5PQ/w4ZWKguo9IJvPFVEIePgVgHKoClgiwfBQKRKJIMqs0a64roXbCJSXQHV2ogcIYIp/acAj4kK
QdPKjGu/We9DfS+0CiEa6RxHTkdjxKc6vu+GegjYejevAYXe0XgPV0jfQv1cxaxf43zYa22HqkMe
03z13QwOEv9JT0qjGkiVUpIwucY5m+aLqItbZRFAttfv3AGx2+y8Na2M2XiE7h9pi+JcU78wEiX0
qBCy9O1dIyyxCkzJnrn0PM8q3IBS0MVS4qKe7p7uB/+fs/aC95TUgkrHF8e9VaZ9Lz39PNdHpUPI
YTjJ7Ivs0kicbInhLyWkPEclzddbWVBoUL3X2kCPFTp3iUmDA1Xbeka37lHvgdCeLbsdIX4ZNscW
nkCaVavOpE7rTEnaO2odnmhkVKNy8htDgA7MlM56w4r9zptgwZz0EUSvVWvs/lLAIUxADoU4gEZ7
zoFCiW+P3qVeyB5S9TIV/Z/Y3j9hvtPql8d6I8kNoISfSBdWWKi0GiLw82z7EkQ3+0PdKo3xbwa2
JClctTwKBrpPJB9mFlAfjU3k86b0cwRl+zBscmPmvGAEw5GRrswpk9smhzzv3PyYWc0KDtVQDdlO
gSfMupS0UDFERCrYjbRL1baa/7XWptBa197LsDLhH7BDWjmJIWA7NI0Jr4q6Nfo9xWCZlMtmYptm
vKWvJyq9naraduvPZS8kBhVeyJxDfNkTgtTFqCHoo9LHAM+mZ3AJS5/ZJC+e/9Kb813P/EBxG+ye
qZ5NkCO2AdMeac4ksy947ZY5124fQsGxllwuLevcQeHxykte/MPn81HRfwDlr4V2vAfAV+OGyeYm
P2OohWjip65eLvBcnOlERi7ff01OqvzUO3EuR/JIj8/AiShLgW1+oHcjopcvSP00IO28zAFURLgD
a1Clmz1ZMiTILfHm9osUMruqM4F+JqD7Fr1RsSCSePG3MlRkXHMRh7Top8K6/crlWkfExbkO/XyW
EDPs+wW6cTwK/xZOutuJSWwu/79WaXxSoco7HxX/OOVebRQLU+cSs0RnOdstGkY0WVUzlO+mX4Xf
EKJwUkWX9q880ieBFDmQh1WhdlwmQWjSThqIKPUgUyEFIHABs5wItG3PRZQ+X1hpS6oY1DK3I03L
ffgFRAxovUOxNHmCsBG6WUQHz82mouYQ/gLQ1sdrTTLUtirF4pRFzDd+lZgAaaTN36Zt9fGOMQ5T
Z24oekesoLmjuGWenCe8CaaW6VVJSO5w22GfWM69gUS7XL4s7o8vmcjzX+wxZfDRvja0HRbIUdjA
EC4eo7HQD3niSDCfLQgV7c/4k0ODSGGlnRtfubLF3DLI8+V7w/75gn52oFBwPp9mNPFEnSxdCXrM
Y1TuH3XVixUWcw2AmWrqwhNHoKKiu22vYz4leOizTlAizow8YP2Vn1iNHnVXykyH1Id5DpbKiPn+
smD3G+3M2gk4QhOE6pOrDLwFeDmceKfn5r0aMMyq+VXfUE8ysv91hVLcCaSFK8ckBZU2aP3Gwfqd
BZeKb/JMN+Mgce0MCzn/8WBzkh10L4mm7sobxwFkSRwWi7eQ+GK1dbVzCNG4+lg04ySuVOHxkScu
dga5ANXH0HT4yNmSjCUePdBidYggDctatvZswtXudyKcO+/S0i5rFDLmmEq7mAudwygUOO4N6ZgM
0XeVIg/KOIrkt8ZLb0soOoqfDe4J0yPrhtVa03md6Ez6/JFZX5T+a7Ry2fc+I6wOH7akoCsT8prU
/eH5BmEG2J3qA5Ov+MUQ6Z0glm/Wav+pmK7mnM7pCq7aTNswp2CmxUwiIMjHdFhOhABd6aUidPFU
bHwoiwfxlH0F3/enOPG4SoOMJfPNJaFNpn4z3Flyv290S1+Sh9udjDN/4FZiq70JtxruU9MuMkXi
d1L9F+l2wSyGOF0EwZ3xx5To2kRjiJo0Vcn2nisZjLg1FuGayt268iCy4G4kB+AxhGcLkM2Pm0wP
M52V6U1iEhDVL8UFgmLy9rKjgW8PRzdTXlF4SM7a2N0KXGoyd/UPRJtMAnWAYC5Ac0b81nAuezcz
CfIJk4hKuAyOxXmzcusT7ifDwN0TRk4xY1Wu9gPzi01PIxNgnm0wRflYPlloQrGtXC63EzjarhBY
WId2Tof7GXA84/+7Y6trSd/DXEUnhLSJdn7Ejjj2c3gtjdHRGhLQmMmK5tofWryLPs4xQTU/fU0y
WBarxvK8T9i6zIvwannXLS11tYDJsc4RDvosH1e9DTvTYv7Tf8vpwSn6PH+kgV+lreWFKxrbYy9R
wx8rfNl0WPogodRkyyg/Vzv5TypAmqrfqGNmEGx8mUUDkhQqPdYOLCwYszz7axV0HlEosWd2OoSn
zgVlxGxNtwVx8G5rzzFMFcirNTqKkTI7YujgljLx2EZoXXhEx8XvvErmcbDffM985tFCHodd7THz
RUy5cxzBtyzkbR/o48lO+YLqt5RwOYHs4sCUZtIQAvDFYufo23hy8J34oKmRTIJSaMrDMyXWPzDc
48miLf79kBgxjGH3UQ4ELcdOyLuOUII++EySKUMmFvJ/4zWVC8eAfek8ymRUQO/QhDxNNouj5ItC
M3glTPszf68Cu6oguBImOc4Ms2vLpTP30v01ZU/DYQrQatAF/19T+BtBwjdbRvwclwq2wjNN1FZE
Jaaxyd1tcu7ANgU9jGNp5++iCoS9WEF5RFUwE6oEPYI2hUzuEUGhwOBpfBJ2eM3Th+X+I2zhFFdh
RX3ttliPir6KCQzbr3tGXq/m/WfOwyq0nbitBPfH6HN8IRXlYBT6AUCF5GXYPnP4LILMdGvb4YJp
P7x6GQIp+cEdNqZobmUBdlq4xlC7uaVVVMNYlnPES8BE/T0b8zyC5TJ8HdQCx7UqONAbrynPsKTj
+DRUQOR1+ualzHMukBl5bFgpsu32iG6Zf8CCc6ytoCbeIjdJTXVL7wGLeqiv7C06UK4LBkenF2Rd
eh1XCdp06Y7kzle7eY6tBJZ8iDFjO4crEZx8JAyanfWEwnGJv3MaBqaCJ6MQfBsoKFknJCQbrCXv
YMMIFfBozfqcsYXdTBOxBTB9c1hsOCb1FsRjpObsktszuCkAob6YdC3SdTK+muznUgz1wv+SGabj
psm0d1je7M+k/IO0ViBR882Z7NG86FRpfsSoSHWfQX8LYlr62gd854YwDlS1HuBJ4VQXFRKnpxfA
U8CsnUZOK+0wIIy7c24kHublKCNbaYnCtS2QQOAUfgb3uI/3stBj65q3/6ShWP/3Izmb0WNq1kdH
2HSKJxBnGa4PcC0CWd6Ys2SmjtXJpaJheOr9tuTBnTm0XO6xqSjOfF8E3Ez5dJ6/pRo9PdJsXl0a
T++H1Rj5GxaDe6F4QiFJkLnyblXJlOtL+zEnqqoZ50WbrGR9BSb3vbgLzKORA5VkGvBvv/zpDFRj
AU97zplefF2AJnImqbCzPwAduoqy2QnQc3RizawED/7AbgLa3FCl/w+gOoXHhtsKkQf37YOC5bJN
SdV5M4yO/voBxL2zkyHGF3i0LZ3SG05L/pk73Kb9mmD0PyFODM3WGwGPrJa7b5z/lqiJa0EVu6po
BCYqVeSxio9O6qDNOjOl23mme7Tt/Zl+rrOXe+v9E8NQzBg3+8vpyc97iw47QraiBEQPrGpFIMN7
TsWzzZDUyCH4RkIWQ5iOA0B12bRodjNONZq6WvKGjZSQWZ80cBUSOhaqwse+TrM43YVFNq7yFouB
V6RQxKnWCflSfqto+6L85UEy4kJzbiPLkFr6f0lGdEtt78gvl0Axovv6B0l2uFnrh12Ik9M1Txqj
+ZSM0HBPTCJplOU/+YE7uNrh5coivK/MJjTWQGS93V7+qiLVAD+h9mC9VJQjTkEAY9PcckOr5B/6
1u7uz/5s9Tu31TiZFJcaWSBGMVWmlb3VmWfw6BzyKrOfcBKFhodmrcd8FabU2xDfiRFD0sRZWkUN
/Gnn0wOiHd8wLL08RfSo4EKqdfiK5mdYj2yrmEE++PVtCFzIGgRESTie7umNQYa9xc0SBvT27adm
33XX7sqcuDDpi3lPUTMT3sh5jZCKmJOHZ/GztCLIhO9jLBw4/Noh6nEk+J0Qo2X/rfoy6qtFHvlP
XdukUlNJmaXzXkxJRSVFD7ND268Neexp2ObF1kiA3dZjQWkCF8wAnMIWWUFoNHQ8Gg+icnIbL2r9
MHTlBnr5+n1mOFySfx79m7TPe6/u3OtF3bnFEx07Jk7AYkXzj57AqGTDvLjDC+Cc139hxLFAhmgJ
0HQXetul9vZW8gx1lSE6n/IFZva0kJ2x+kqZJM3fN0a/dBFvCib9S+5bUKEpHF08NFXu8ZLHlkMb
Gtql2VUnOb3+4bkcuIw0v5A8RgKjDzRewBsHhLK6X62o+CxtoPX1TMOaw/iBBRHVaq32LRcRE0Wj
pq1qF3yTtWAHVdx/et+j1noJKsSqkE5yhtsG6toCUM4ITheA9X54uYJ6WMBjuJlvvrNciyv807J/
3+8+sYbGIBhWSG2MOyAJrpR9yHYsDun7rHzt3c2GIEBjhuv0Rtpv3UJz6z1LC3Oci21cy3MPbxCb
QdhiyQ3GyxxQi2in1hensek+ke7ihzZgttBsM5QzRpl506IUknsjxFSZvwplFEVJX2mcILzHQy7W
JlNe9tZw+qu44XICIVBG4twjWBORrSXAResK3zdIO5Y7WI3vSY91z3IyGOaPqmd6HXxBRWiOeO2U
J60wEcughvd3Hr9Fj7su83dbxWm/afO81CfqXAZUf+iLN7bEbmldO7ic9wxy3CzPdEqNfa8m8Hsh
20MNMXbQd2rgyguSn1FpcS3FLRmLimJA6fhW8FtcZ25hCZFsZX6rLVPR3//bKvIjAQwfig77ekBe
tfX2SOcpaS9+RoxUSV+KDpT8Mv9MZ2g65fMCzhb270pimrsIMFf3nHEuFaX5L4+FgEnwktRwMEm6
6KdGWnk0tPKpg23U1/3uf7ftTOC+lyRuODW6kYbtcvn/MP3Vwaobym39BV0FqhsYTENxm/oSsJsx
FZzJlJVK5brdbp3RgaM2km9JhWgtOBTjf3X6FzFQLQ7g1nZLpV03LoW/q5ZGByg28rAi1hW93VEz
UbXecmCwbps2bLJ0hVNxkASuy953wTjcSRXQIEjBT+5AVTe+Jj7AW9J9FYYMcz4B3v1yG5/XGtNT
M+ANRZqu67aMHi8a89jxNI2piwS2tk3U0QaSQT7KixvYwD9/CN4qP2rDGz8QQv5pps79Tj/q/EhD
9UR3qbHxeJh9rWksiWe5QGTLdk70c5tA9A+bU7RTeJw9SER83LKVKrhh7PnbyPKFsp+9Ob2nP5DU
rEJEny6oJVPz+3SanC8kOzg2wfyoVYuEQv5aA1mK8KxdyCrodqBDTY3ApRZ2SXNB+zBTwLkXieek
zZTGFoPP2ROHiOul76bXbwow3Vyvt9xOVsAq0MrC2jGdtRCo5v+SZuck9C+O5xlGzydbAGzDOvNC
WP03NhIFe6N1D7EACN+BbUhl5okQj81fpNlPlOcAwt/N8OrO6hrRJ6rqTj85uwFlS8wxgh1fc0Tu
ulUpAOTtCUazqhBSP4ixGd8IO6nalWJNzEQizFVj8xz4822RbZmOTietDVlvEbtubbxvBC/o3x/i
O7qzzkoJYibgNpP3sUa1m7fXlkSlYdbglBrq1dsMHWmvuvsu07CFxDZJfQB8UAMRN5wLc8tf0F4r
7fZ/6oazjX0uwQV3UghfQefzbW8HxKIJeIT86BWlHkfKaIfvY6P3sDMzynucQpQe9cwh+Osh23+S
gs7kL45lfd2CD2R524hiGUeEWRxVfSXqbWnGUVHZdWmzY46yLC1DcGMmB+8wcSFUh2iqCx+OpV5Q
7PYm2wwEOhJ1lNwt9Km64H2hmdWXA4VcEqvunTkbgiO7KYkJDf+M1hOTPfi/68lnrqY+rX/zMRr+
xUkko5YfYH0cFE66yoQ2KZ+HchWe2VtWVadc8SyWgoj1VgwRFMTVd3Na9eaFlNpBadtq/eOeDva9
b7vEmPsGVHIpIrDjFlMYIk4pVXe/B7hl/uTMwMrQdiPqSSh6rXCTwZ1I332/F6AZhJfPcmXdAzWf
7G6R4xjI6qeBR8bHptHhKLA5HW20T+4Y8NC2uajq73W0XwcpJofguFdeW8eOu7A//r1yd23hLe6p
B65GHa8wUk6SCD1CF+KwHcqS0JOP4OwDxsi8IuqDr4IUqBbWjjjUu4nb6crVQdsTPCb1rbJmye7w
+mex1aAiRFLyQ1QruNKG0fdG6pvmgMiuWIA+D4lY1yBjFlKqnDYBJQxzYbuQR3UyFRBXyOy4KR/E
5aLPoapAIzg2saq7c/x4SDeb4S4xmjeLQjmXZGICXS5bBM78ZsF39xHZKyliXDC6hUVisJjTYrSr
g/XTY1BsIEkAwSRJYDuH1pob/o3G2d6CM6IO6Irf1mvZb912uoJHyF5HB5fLgTfo8gF1UFDLx9d9
k15gazR9hjsxbaVnWIuxrZLDJl43yyh8nZ8M7u57mHi4+ZPxHuQ5ug/KS4HwI/cQSkMZ6QtKigft
I+hbXbvqRuQkL72X3n5jD+4IGLC6V0FC8xAFCBSOm0DIr5PVaGoIY/xDKBCZ9Rrhu8HzdI31GrfN
+CkwXrpOxz+9+1SErALlKz4kdf65OKytSKwuRIGMxbiFm9phpgGqcqwYK/bsuQuywmJJ8NhmJFqb
X1Fn5LdG1AECX42o1od5C2IGaiFYPZdlVuytPQba2gA9iLLqY86uvKdJCRz6eo3gCw2o61Wch91U
o9nJBx0liGUqTPYgpD8oT63nltD/8tR17j+9mUrCP0O7FUWDmdKpbb0mflnL4b4Xrso/N6qQwcR9
/CPd386gCHNsEITd2h9/IsqVDId07T+GJOqP5j2hpZYdKoLeK6rmE+D3/YDImlFQLMDv1aHWK6F1
3dCgS4BEB9/JxRV55XYE87cEQi/0UeEtQv6PGFGV7b4sF5Y6PJB6ysiw3BvMP3BWtFwyl+m5WdBW
AA+Lk16ICH4nSiC/0zS5DDmziSFrdh5mszz1gGROVwNgX9z+paHBwccHxVRW/xxmV1cmVeyyeGHP
vLIcUSGlBP9TyPq2woKMLklRNn2qs82US1R9nvtLvqn5qq48v2mZCsMLiFXE9QNqUD1FNBb1P4uZ
CSNP0v1NOCHdDxqs2vzX5LswS4W7iTl5FM7CvoJLhlaKwwz6zq0k/Xcn0daVJK3tTvgcy4/HURwn
HU9aoSEBxmS4T+Ohqi14ABy8JHZVbhPgoMTAbjeiI0FtWHLDXNSreD9AzN4t/P/O5s7HiWciyP51
JksKuowZxILreWkMIdrSeG63XkCYmUl0GteBNr+ieraeG0ysZ9SV/lbXBEDBPUBggtUyULYJk6IM
CZvKFPY0PakLtTpZiLhRqu1SYNvLK9GHBMXEfwwvWPqZEXYqJhL8o88CwvMStvSJUsSLB7+PdhFn
4AYnNTKzpJYDU5jzwMOIbD5bKjSpgFQo1p7Py3BXEcZlNDGO6PwGO8VoZI0HvsO+yowgMCIXl8Uj
XVxdo+1AS6UXAYcetE0ZBXzxV8nilVfvMT8HV6ycqR00GO4boqUIgAB7pTN/Wcs3hr66uqw86/8i
BKOb9ypiA5tFk/veUFerrDSU2ssj0T/y21mOecJtBeanW6mAUUs0Rtm5tREGD/SPbQo8B1qQo5ek
hJw4N7l8r5CgpofZ+as8aNnXyeo9lxIE0kUbSyQWtaDPQBizExZflXqrreJJbJOUmB4jcdv9iG3n
J5dqugRfBsuUySzmjby+f6VDfoCuubZprMA+pG7DLowVkX08tYOEVQ+8Rp2VT6ipMm7yFRpykrvH
AF+o/KathSZaDJeUy2Ke6Q6OBXCb2yfm4dRwANFg8ZUHDRZLCbzWZ4MQ606jO9NfuaJ72MR/a73U
vbpm+DehKQ9r0cL6r2nfbCVBnMKUem8qGEYFDsBXmVb5TYXRVr55u+PXshSa4QSUto4gRTQMBfEo
gNC0y8HQlaeV4yHYr/WQtaOGlB2xznZOb5I98uHnlY3yhXS0TLvdmBIq4Fgu7S7Qn/S3KcF3yEPs
KNotwRqTxDPQah6f2AlwwyJfCzd45C1qPndBMVM4oqW+k4y5tdezjyo70pnB1LtCzq30BkGMU4Y+
QJ1ov7yFdKqjosIqPmQpPPebba3aEQ8kXFnB6ONsI7JjhhldR+81tV9HZpD1aUDTMgOcQmq11yXr
lSczNB2mVz3R2z5yvixSW6jhX0jihjWCwLq3fIW0vKFskiCkWqBZlzlTWqOOxPdSBcUqcb79vAY1
SvYKxXvqfnHnowNobfzvaLQyfBNbtSxlbn5/sJHnGRIiWD7nxIJ5GYymrCgqr6eupZAzaa2jkgD1
+bIJuDRagxOkFN6NoHRDaXMJua+nCaGOyFSAqjGjeHaxR4AT2vWYCYydbH75AM4hsJt631X5aqEz
VYjl3IoJpXw7faGuIGU+4a3h6KCOWPT9vEX+t/Q8A8gxUFXIfgfEP+H9rdL89CR4gB4jwZl5/e/m
TY1GGBZ2JbBFQMWt6bQ43i25kgu5Jl9qrXPG6oAnD+Dbm9wWPcvBHQsRZVabxEblvMJWWbrVtSTq
uciBsHYlNriFORUhtMiTNn3CNaD4KD794cI7kyqerdHEyVEIOLN6zpbprhLm0PZSsaLVMA5d0KqK
VZO89Sa7It929++YI5qbRUhNyDQc1D4PU8CNc+EHk/hyELmYo5v+Q4h78cR3hyUx+IDyLdo2JxmE
2fU4DUuy9vBen5ryI8WUzIxSAJuaXLKCeMUei9mb+fWAE6N/3FrVjflX34zwpcPseu4jKTKPtL6U
slyYUxorsZHsQIxMesx2sG3ZHSr7ECCiPnyqKrxH1RQdiLI7967CkWAaznJK1xDt+zuILzVsZIc7
oWeQXOEUH912QKg0urnZ7yuw8RcWGa+I+43iDzvedp9qOJ5b1T5QyvWAZzoPVr7PDs3uNrHuRvyY
wHZBuU6eKPGqUV7P22z124NhZYILPlehVrnlO+ArwlLp+2qnl/tpzax+x6j1sd8aiqaH+3nTWBwe
diMJapzB9UDkDLmBeVKdL6e9jVtQN4LD/A7ON3tqgYJDVEhcTT9l6KBLi7R4CVKKcnPXE3C3jIxA
4x2Ouey9J3WK0gm980SHFlS0GPSN1r4EPXsvhuWVhE4pP5qzPfz0fwv7/pOTq8cE+NX7avjxCE8r
xRaIMLDg+YbHUVC+NY3wF3WqItFcuwaL46Hk53LB6C/ngu3ErFly1t3MNku9QBsImDWDEvZRXXcB
1yuIV651CVI9tW0M7Emn2n+dqwcF9FhdkmvF2q/ouLXpWYJZaGVOnKpHJ8VW6yfx+mOhKJeGm9rv
p12b6QwMGRCHohOupKP6tm+zQEeaUZG+Gncd+3qj3WRe9rfeAFk4xsOEcgcqYVPBfLJzCRfvn3V5
GbeAnDltwDys3vkPjsczC0WbB6VoWYvlA3Yr6fAIz9mtGuc30yB8KnuWl+gD5cPVJ8y5Qky0lwk9
gyprqQbZVQJMOLk2LyXVG+IOhkRF0lJuEYbvzKMkneBijuWGzbC+s9IO755cV96QFWRFiq8M/uWH
jgJajpHNIlDk6OzbAmQc14zDhohMf4DhaSueCuwphaJjGbzT+/Ij1g5W9w743RWNUFDuv3EFICSR
xz9dnvKgzo6XUuqhKMv+xjDTRkb4lj9Rv27m5CLyGHiAlLqfUQg7HzrTMm3qk2TQRUtTsbvDlA2S
9BVuB1n1HXBa5G9qdksT6qE9JXzPg9E8zt/le0ApZNRuQOqYxKBpSdQAJW7t1MNq9VM0exT0xLIN
C1ssqrpD2SS1Zt2P6G8Nxzvb/3W8y9WCcZv29swYzIOtm7tB4MhKOV/fPNbs2rFF7lMI05jGJKxf
7bTTaBkOaH9YvLKKW4uc1lhEjTCUyCWMFSQO/JhrwNr2ue2W99TWTfFzMZ1P1A9df7TD/Rx6bYxX
OuIXt/VyI7hSRh5t73v+vhACIWrMVq/OFmok/NdcrOxdg4424ohvTxVloIcqHAYzTJO8eaMNSvkh
U4jO7sRggjrW4tCXfImEtAC7zrZAJydZxEt38ZlcjDVFJQ5NnTZ4fqPxUQnyLdXOO4bpLr46DaJ6
JdYbJGxD0wjrRbuOhgHsw/qu4nrFkUJwyJojPcREylDhCUwJRK0spGrBJy81o3TC5BK9mVrwiO/h
tbGvE2NgQPqDNeZpPwRFa0uQNA9/Se+Vzq25xYThv64/EHnWxvxbdNFPFL5GFJfLdMC9c5is+27o
Z5OWSwjanng+Zu7+tPXPAMY3oFqz8++LqBU9gDdlOqkNXGqNmaH50oK2n/mcqvosL94Q2ioa1LeJ
PxG0lmMwJhzFCsTut0lhezUewFaz47Rt6MFS6tmdpZ05jqRQZmEWxyr8OM0ph452/wR5AalrNdPl
ji+CaqqdlC5JHZJYcPp943XV2zvDuKOsKzj9HydMbRAFV8xmbqIpok6MxtcTNBTNQ2ra7xzNT2aH
5aJTE36sqUONyQyEbNaLYzZgrfDQmgso/q7uCoOBYIqslK53kYjQzmz9b9jx9rqcXL891bebH2XT
1fyHFEGZP0eSbhT9V59H35n2sN0gxxQSeaaDZvLU6mdohA1LWdr4PZHL+8Fyd+PIRYSkJqC25g1X
DjBEPL50+bOtDnYByEF85tZ5Hpp0OtcKkFif16VCQLxowwQfAk0Tcba4eQ57udXrTI3Cex8sKkEZ
cOy9yb8vyboWIFRe1KyX6cmIPiJmIHbAszAsMnEMsSl2Uc7Vt1UuQcb66OSuAr/jSMSk5DUjyPHD
X7Ql/XEXItkKbArRZ8pRkXyYPD6D2jrNBrnqRuwUQHkez82xB4L+E7IEoRW1asYoUBFHSAdn1o0T
nTZzH+CnsFOqykk3S3EFW0QlbP2eNZgtV6kXejcTSR04wVeXP2pIuKLInO4Jz2jeGDsIQE/0ERX3
Y3gLGIVs73fk8D10ghpe6Ood+LGcBWatWzxSTBuSJvg62j5BZjBnd6C0erOjgbClWWQftr1TI5jY
SdasLo81XSfiF9f6XBsAoog3GPAS/BVt8IFkC5gb3wQdTmBasJzt8a81zyceUlOlzqODgXQ4ugdj
3jBuMvNap8J+LZfSKgKgZdla6OE5PhB8y4tfnDVQk6ATLRJ3TErU6wz8cdo7q3NFxm/92kztNZL5
z6bBBcXFtLK2rVGY2SHlljWQ227J49hz0gQoXKwLWI0wwq6rbIpB2Rg8qa18NVpP8ViPSi/5MRpI
WQ3i0lj+pqTHgUkK8fVV8+eEPXmfe/5NlgBgDs7YQsfdHtDKnKD3MXZQt1rHeS3+tZJASzd6qMqt
asbt/k0/vvumRYk4O97Tg4ZjyI5/Nu/ZkVstVOJnncZK3IRlcDiSuPfFTOBez/57U1EmDdGVRhhp
epfQ6sQ27UeWQ7LKbbd4n+bGpdWjMHBpWsQGLpF926OjBP3f9Uz5lITD2lCZV2R5bGiRyKDoPsXr
MumuHV+yRGJ23H2NvgGrHHWlOdPbRhYeCnJmwUTfo8Vha2mePqhK+yReIkjlakETdMv4G65W/u4a
X+PrBFf0qo/AklIB29Jg88b9gapPvPolCN4zm1kMjhpZWffg03YhXU0SY9d1x2QDa5i4giW76cml
qf39w2lIgyltL56vsP4dSs2uFgMhcy6FkvN+SwqxqkYAmVZj9ZLcQb4n3DIAWKBs4Pfvw63q6Vii
lcVLg5CtVY3dy9+SctGZj7R6yV3QGQJFC28PYEWJLdYGuPm/dNrLR3QJ/gIDByXangeJ0WakOOUl
xQNPuRU8+vsj5n9iMEVNbWsTXsJoJCW19rU6tZt5nC3CpLvRS813CM0MZ1j6rI0zyO8KoeyCO0k9
EmGaUavw0MBa3+7gofebs2JMB0aQoJ2ClbPDzV+maVhDMjuN1JpeSPUUyI8/c8g+9haQxWf6KbX0
ScqbBTzXtghk5UQEXHLkw0h8EGK6esg06z7OKmTNqaVdaWw8Qx/pO1VfSRZS0ksCzL83PX/qmCO5
L8YSIJQ8M2gnCh6mBjK6C5ogbFAB7HAF6v5eQGVhkyjzQTalC4DM62BHg2uoZLeoelIraoN3+EKR
2lVyMUEuDXbbmEGOPteU/5t3NEDiiNmHemLFyJiuY/NCkntKxSuOzrUQdH17TUekgGeh/3lzhea0
0VsMSM8EPpXW4AmEDbsyAaSTqvkwHM76XIduKk1ct+R4H1DJEEEwDjVuifD9HBnUswouHZBJexez
WZqOZqQ+hHo4ZPXoqNJHA7e/+Tsp7kZy0XDtcdxzlrNHJ6kOnzaTMNZVY9x7ofRrwN6z7xwJPfBR
4iWSoIy3XMJWn7shlS2pdrac7Kbz+LA22/P3ikNEJFSytMLYD3+U/Lp/aTJcAsRRCUt9p29KRlA5
aK+FEBJBXIYGrCXLodysrUaXGooxd0AxanWlOFHWICJobkptRMBitkh4gfKnPeY+/eOQrDHj1ku+
5JK/Wmo806sCx0mKtFaB9aIdDgg/QMk902ZmeGAf6YkSBwW3ZPdjguvbwScW6WHbppMHmQP4sonE
uVNm/QYwDs+FUi1qXNnjY6Re3DTsu+171RUREjD1qjdhxFvnhxJjaX+ulYQFkZnVX+Wy9qF8sthl
MoE2m+4n5tj7P45hjFSOUEipiY/Sz9NpB1gV72VlKhI2H45ovwJ/TUMRGLpGqrUFjWOBZSkXfJgh
Nc7ppE/dyfjrfow0cjzZoZBUG8Nk3PumKsUun5ZZOaNiIo0ZCw8VqlNBljPFlV0XwJ4F38/+63k9
LJu7A/FDk0TWV8leitdOnoJzfwDV7sLgRtuTVZmIHm/awKEtjj3uvrstAXlKSlp1l3rInLJ1CtKd
DCZsVwLCou+i0Ni7jgcLocRHZPiN5y8Fa4zUJhMdMi2UTjYOo4G/ILODT0Y7GRy/SYRBfbjLuhHl
K4NIKwEdKdfdzGwCpRhVQV7m2GMYmOy0vuGoq80C42CPpB4qNneFh3ZGjpucq8zJNLxSvOrO5tA5
uhxfu4tqJvr98KWWnjklUODnhkmkM08XqWjqST4Iiup7wdkjHfLvqXH94LzJS64LPVXawEOJpT0y
XCYKq7Y0HobG6cNkhFcrV6QMBCtQuhEXH2xkeMjVorzfiVnrDG1c5jFjKNhyOTWN4DiVSFGTqM5t
V9EU5QaSp3FX+ncLCdWFDzUdaKeQ7A78ceYcJeP5kVkxGv+3i13j50UAxrrfsK5Q1gCgvXlmsEiG
oTFKoKGl45fD445ZqSkTiO4aH9896jH7Tu9+X/IKcrGC1tAnE4fHAQ5unciViNAy5lsQzu41CCZr
/sRyxfp+GUvxV9bCu5cYIhHoK5QLfVpK6Iu+xyh2kLZoj/QXAKfoJKXA364Ma9iq+pDZjGAEuqc0
gTp119dQZq+5w9rCAo6R0iQtJViFtEiqAxwbax7bM8eZuWarcvbppnKNE44kUTcJvxPknYQWEGqQ
zNGlDYF6V/qZJz/OXOaXJ1q1RKH5eAS9/1Dv0kF9P0A26sngTp/KYK4Pneox9nBJK0GMCt31S7J+
ft7GOkVYg9bGdgZJzvaxXQd2pO9JeOr3dNXdoPfBRc1zNSZUGu4vwsPfZv4Dxo+qeq+DpKNELPmt
TVoqLt/OCwtFN0wQ3YyCOPa1SxyATWtbFRpaQ53ZCbjVQtBUuIQuJh1wU6HiU/8VgoPYY30+tiMk
3MxMYX4JR0en1deBFjS5TPWCwv7a3tEO3q7JDPeazqNV4Tm7iU3FmxlHSg4UwXp5Tm2q/Fakjy9z
RHrliMvktMyF4FCJ51LzxInZIB81YjhKV9Uq2UULVmLriYnaa95dg8H324Z69kwdfw9ZWDShLA3d
XPO2cLKsQ1gtzoNQmQrCpIVyre3EZ0V8anwTBw8ZUhm5aE9IUl5q0EX8gbPCrp8gYuHmTupHn/2u
KL2dgsUUAOBmnPO0DxLR9YHf9q/6ndcLu4/aW32hi8bZdNg0e+V6ozYL7qiU4CngPAPIaPut91/a
tQ1adBHY8Jm0AOKrRXe9nvXsdReztgHjIlpqSKUs+ZPf0oWaIo7MzzBbqk/PWm3cDd9U5nQaD9pI
TfJcaYukOO31PWCHatAv6EqKg6H+GEm+qohYLWLkYD/9xD8/qOo7QByILcPYnGTJ4TB6gg6QqxIh
wNSRA/sUe+lm5h3KkF/2gdOwWco+NzWfOuynX6cBsMEOZlHiQsZmPj1tspATpIWbBiFk4KYGMH85
Rh+Ek2+mLSAHcPisNW0eyGb/nLxgORYXDpcERGPYVRlyRIxcXGYSM4OnlcsAKXJk0FE64VAcCoND
+W3ifbeBS0cSw94l3A+tjBwKFREJhw6wg0LUyAX7YMKNMiLg3DKbHONtF08GojBpndtwYLrj9acY
9o1R0UZTgRJBaT+3eNRT0e3aNXIs0xjNs9KmT2suUUisPAmJyONiPDzNr62ZzTyi7c9Y+CV+kBh2
7aiANsA7RNmiiXD0nGWLBh1mVFQl1hP2qmbPcnzdBtnkXT4NnapPAQzMFcynsye7RhmKG1juATef
OocGNLyHnkepPRf2fe97Me1ZvUGUp5WrvkslHl/Wh+ItNYeAUIQ1yHs6RMAHMlpCjollr8cLFcD2
ndEYFSDec0LWYy2NOsqaeB+QxuxYnNP/92dBSvpkDorlrJezOokrqRXA/alI3Km1jaSuuA3xhu0I
84oaKbCDdce9jjy9wFxfBikIhRknpO0Nx9xxuhhjBSJlUVAgN5A1aLhzLLCqzy99k66CSTHdpHE7
ncK8eFodue+ibwJQLKMkvWNnii+L+beHE0fMguTri0PtDKI463cx0N848x+91PvNTGb/xIyAcv8r
UadeJmQMiKIvf6bZ+OgFTLmVoooLyq+8Xsz76LzbDtkZnIMu0/cXd+7WgR/0mIfTYlt2eBdhvjoo
6Bq9m/vlFLEWorAzdvT7WYmSWd3e31mnha8YlhivplM0SB6tdyITL3PCG0WIUhXfwESbEagAar9e
pR6CUE7m6MQGluKncVEYniLFNbBOjsEs3zpxNaYBbsOS5JBE+8h+bvM2CMT079rxnMyZDc3TAsOH
TtIvCnUUXKrXOp9mpllYDzRwtFxb8mGbXhFqj8gZ7UoNraaRtbmS9w89SK1SClJypTV7S0j0gzN5
VuaSzGhOmvvKVo9oFAldzYPTJUiOt/NT1KtKTefSlvYXCb0uLvULvSCURBPhBcfNChDF/u7P4Q5l
u6k/w8JLwZ1YUrUXec9vfoghDUTFTYV3pXcdv8ayMFoErFn0fCyiheo8pyxRF6mpWGeZ1nurP+Lc
pt8kLIFSwyRZcUQmNtcoIGsENLFOhXv8Rc1YYzHYN9n1kyF+HNLuTxeDtAgea5lA+u3xX1Vo5ind
ya1+i0ezaB8kt0Fc8iTLaQFTongbGDlMqiIxTqNzTBZiYhCLMpRpw0fU8sQ8OBt+nkGKbXyXdJwh
iXX/z0KwSgZx3FpVHtpWe8wPsV+ywg69q2TOEUEF4dEpJDI6Oj0frr5cYpAEZxlKth6djoy45qON
12BHXuCSEDZtZFaNDhDQU2TtJ3ElJP6OYGbqWnGt+n6OcDob+/DgoZU9hboB8PJQT7LQ/7Z2b5rx
7FMQNsuHsrQ5mKGg9G0ZZHKA4D+e8YW3Nfcyz4dV9zo7An0AD0FVKmLg8/v7sXtbK4Bq7IwRbG8L
tbySp4FRmht1fp/evbheKjMGVtFn4/DfZfFklz6kub+VBmJhATF0DQ9WWe1oU0ZfjPoibHphVxdU
NImFxCq4UiPr/UWjY2r14p/omP1+mpki8oaZr3R0v6WJPvERgiCH4a9C8vMrWNcXULWMxLOybmko
UYEKkapf8QMyUWxm+EI7dggdzQH7/hHuKXik7djFxfkAiHssQMoNbTobqv28NT5sVpwUPQGIeTQG
d7Ftq9732RtrfJUW9qQlHoh7uw5L3/0b8JAekMMCzQ8Z8qixcbRKFn6YHxgT4TwZFQ/ZhFbby4aL
l9kpbGmuMrslx3hNrLgfPOsEhJytfHeIpR4SqGovY/dzjGkmZByi/DhmI8anNQ3KTJe2owGASwSG
k230kvagvtNY8VtO+S1KAQWXUAiCvJfHCgy3oDZ9V7BP1hWNS8f0Fvl523Xj7HWA8QBlhIArDDXu
NwV37cX5bGTKQCMxXnputU+D56h/v9/TtJslSYXwlQ2azE8u5v80EiAx9y69zOV45KJBPG0zue6z
KNHEvv3tlbstwYCfcec1FgBjW8vn9ixbqfc0kgpBKcBRcLESlGpT3+GsGDf2sW1bkkjG7niigEHZ
SdEoZro5w0Z+Sza52l1xen6dYpSqLo7EcHBJklmq7wSRdYrK6XoQa51YAq4LZNAdGQloqMrMGQ55
8hm2r/2pIRyYgyWteU8fJ98e68FCovbLtU3We8clxZUQ1fXqoaq/n6FlkR8sjvaC9eo30QkcA0gU
VFgFaNe8OXSZYEywDSq9hjTZcXHuvx1xhU+v1TINOPpjLfCiamG1GSLu4mp7n4dDSi0O633BENSX
5DUbDaT9ecw0ubJAuVOOsaOQX4rUbmscN41jVNfum7NKxDffdDsaMmysiIj3Rcf0WsKnI0SMauAQ
YrVdD6ZQkEC0wfPlWH9lJ3jvI2PqSkAx7RsockU0lQ/pYILJ7T43KhNJCChvTRCIGOPe35NLRmMi
o5Oy6Sxf/uSI+LxzPi50L40c1m+Yl7V0VwEusYBLdjEu0FzWYQR9pMIeI6Oq30ZxUTaVlsd54F7K
nBR9f12Oztt6TnVgYojG+oaFVkqcwGVQNjfvKYFipTjKhJONqIDeiA0v+O+0WVQ2eKlFDkC2Y4J/
WnFGkmSOxB0doPusg5K6fsq1dsZPAgyERSX0wmnvJ9pDSkoWdzbTuyE1oiWxvNNNEY9C1w4+aNjV
p/mEpjfGC7wVfod/TTJepInWUe/wLMEFwZtNsF+Y2fCB5XfJSB0sDx1wll/19Ow9gszRm2t4U5y/
gJ+weIKfGsdzG6WrL4iFB7INOJG5yRdm2DegPNQGhGgRykZlxij1bLe+t4gTNvhh7yoCntUwMZeF
8ANULA/1Hsr8SgBXkJlcmjXHZgZ4cWftWjx3oLv1MtlsYi1Pa1BA4fAmKaKtlI8UG+eJ37sqRDe1
7H+ivVrdpjJyrz+wJ6ZYo0C/nmWpD4hxaxVmtkPBssgucr5mDNihYlv8OicupFIaHozpaD8s3kWl
O3Pcp07gbZP3TZ6tZxZA6gpdNVwgv/pNIhRlhQd2aqsGi8WP8E7QtggfJGPzDjq+tzMPVgCS0lf7
dfEesihwtJmyNkPzn49IWX+sZXo33L7++Rq80Ye5JEubpdu9xDchY6H1V7Fvn93KaoZ0rAI6hm4O
UgIacI7XXHC+LYQOHpLPZxjhPefcH4016OnnknxNivs0qPGzWvNzuXW02tzdNFxk/FYONZeGgSqV
bI5D8sjUGNl1HYlnTXr7yx5s2iTWlWiJfoAbVyWH7kx0F6UXRROYWTe652K+mmPE0Qx9OtIfh6HZ
zR7t+9L99rZ+ustRBM9B8M9idW4qSrmFEU7v1ZWZamaEqbnJgUonNlmIRQo0hWYlXwrx7w60Dna6
/wgzrpcwOW3l30U7gXBgE/B+R6cTV6d+O1jyou3+hNteOMF14HKj7/ltgpxQYEpKHRRkij+cvor8
Gm9iQjHIxeJc5BEYFYDiNwoxzzPYy0+RnwT5RI5RfJMQxDilrprTJFaAwwiGI/ggNkP5mpOJlctw
4ilbsP0YlRdPkamb/S36RJ8Qt5Leb2mH3FS42W60YTknMeNkWNQIjBccZgqATZDvH1UEKinC81EL
QJQcqeX1skxRwLopZwi8cx/PwfW5GJqSPCiYr+9d9NsiFyl4Fse/rC96UkW/LBJb5zTAk1TFXCjU
0uvUYUxopWc73Gm7h+Yn97Iip0j7gvqBFEDxBi+qr9ZEVlFfvJ769qKYOlUpZL5WuQlfkTxTi7xv
dElmdlTBRFB4wiOLcdUAHuO45R8j1jXHKNS/XLxHIYJESIsDo/oLrXSDLyGufJltXV3LSuROelVt
rshmMImVqc0xVJvagGcgw61cFssj2Ts/Fm+8yQg3BcNqFjyiWc1jgJeXd2DZ8ewpIFF1bw8Er+OS
qvNXU9Dype/Jf6fvjluEONZXhLbGfaoeyeWYkfn0UbR2rtYw8TWVsC5ZQDq9P0k6OyBloHmM4jPF
JxgrSHhEQ1R1JWOePzC022+0cfaD5ndmWW317FmeGHaZpO9TKwDZ9MyDObmdnjgd+3hdppv9aWJN
7hHxz3j/rom96sUBh+gOcLiJrWXz6o+qshPahqVIKj3LN+keWXhtwHV55u8DEsVgO8UjYU6s/SZI
HTWUTNPIGF/jbB+AoBB1HctF8ts3k5zt0+3M90qJA2VXxFktMSmnsiGNP0S7RkVLT8OQtZpBbOjC
A9TFhjcl5MtZzZp8QqkJS/1toxY9ekt9vdbmKlOkF5jFtfhgRw8ZPNJR9zyUb5nBvsMBL7oxUy9F
6erH6DUoDMuyw9F6qpiYAOYNQSfMSKa1GAIvtQ9AVMec39oDuj8C4vewut1v8qVOzbAK6PT/m7EM
jmEII6xv5mWyruULcA01YPO79kb0Rp5i3zxkRfPOnJ84WFq3LdUpwfkI+A0w/2CL5YBcEPpfixes
o4uXAgfvSltmd7yuE3zKGc0WodINYQMjZFyl90Uf9bXnhc74p8wvu8StqDMOUSjvT46tv1OB3CsD
nKg9oh/g987zDW/f0iHpB4IE2I/+EQmUVA2TTae0G5ZLbOfnIjggFRiETOw3fAYZRtXijYayRTNN
4rwpsYVPOj8Z4jO9aKVmh3ZdKvZ/n/FEX1tQG3IKqnqnBeBbrFn6HLA2ME0QDWR0utLWF4f/nGIl
B9FVCJ07lQjPzHPDK/mRa1e4HKeWmJujsCcmFMboJ+1M1Le5yVPzAxhN2+ESVp6F8mo8VoFdNdM1
DhYRbbm3PWzlk6GIK6WrNThZ/RKSb/0EvZc3WFegOnB5K/cqsB4Ow/ixyvCu4uB2USVg31ZLDX/h
gui9nV4Jt9nN1XHPs/cTeMFPKaPDvMpLaS+EawQOtG4gyQ1G3vZXfqHgQLIdaHmdmsQtXhYzkE7N
TIdSCvq6otN8xO14JkWFa4WfQHcyihluuoEO2GjX93cTomrkVLd5QYloT/wDwCrPZx1vIi/hGiSL
MCgniCi+2b/OtYffYOyt5mDsiFekoIh+Fi0Idp16tfe7iE18IM6y8FmdsfBALko6NJF9/T6814xo
2MTdukZGDDSyhWvcmwwg0nU0/5q/Zrip1nvIpVO1poZfg1Iu7S6oXT45stQSGrt+ibaQ3iBtXzM8
hmuuN5YHsXIFh255h4dZ9LftBIJk0CoD/1v15mirp5pHvg6hbJsjm9S4Cxc8g2kjIxB2jil9g9np
Y5yABDt8iERNN4cfzuhlsrS8eO5OLYx7ZPl1GBx9hIqgYoHiJasG/rdSdiVlhtTMPkNywVztWF8i
y7sVsSL2PhcPZP14fruYI8aGL3Q8rDNV9piuLJRazx/Bc1oqZukJaSIn9sKGbWlwV/0/fzmNKUa9
5sdfnfRirDUx2EbBZ4jJHMRYYEYmFJa6btKimoVFTA1RL3Yqo5NdR/oy2bqEdhYXKZit531JPOoB
DsGI49YfvNUsbXwryyP70ybG2WMDCvlxlcsFqCtxHW8Xduni35/gNdXT90o0VuTvrIsIbaEN74ei
tFMu2hEI7zirAhccafU4Ofxa8MJLGSr8W24mLJjqgBbCBMrXruQSQmIobezyxEesjq3+kchM1jx1
ljvBO1Ro6ZifhRXOYlaoTPG6azY5O3f8MvuPUKsjYfLwP/5HNaz3HIn8VdCAvvNbZPYp1vFXq/BO
y/XBQSywep7sB/V/3iQikjtbDxQKpc/+Vdu7dpnueSkPBcByZ5yENAbq8ibOV0nyD0U79Pd9oExK
n0Xj2f79Fx3aqxb2en+YBe9xz2H1nsPbC3xN8wMgW6/DkKtOacWNtQAuaYlKYSc1psijc5iacmTj
deDe9vQzoeZ0Bx0cSAV6YwHGeWUH9wXX3v8i9KtWnnYX7oOP6YLlTWHONe5bw8DEwxQNOktctSr+
Y9LCx4KXwy9etP54TTL3mXItCDEj20JUSm6m0eU2n6CavCBG/9E51nbYXKtx7Yfgf54SLD8AtW8z
x6oEAr+f8HPcCDz2T3KydV/dkxz54+XF52DyMW+cOaCzXzd5YFAOv3kJc9nC/wjCD+NOwOJCYyTQ
ILh53yrXN55E0dT7hmApeIxoz6ms15SPcnGNxvIsFqeROCnRU9Rvmb+4v7f0tbEYZYYfv+pst+lZ
XV/HFyMQI/4xj4AsV3PMGtFa54gEnn86OxSLzQv7xxJwbeIxJBk/GpZEJRx1RERPrinVrShfoWdt
rH8n6dGw5x6TXnW9UdxwiTO7kSE+O5vb1utuYhce+LbbaUger515c+8HWbNVEj5Tryl1iNXGLUYp
to1LjwFJnAVpSCZ2+GLalW+kT6qam9XTB1W1OhRaw2/0OlvfBK6ZBYYCXlWlJZztti0ungXWLB+v
eqwOzAKIHQkydOXk2jO/orve+LuVPXNhsZ28VKu4gfvahUGSh/VXQr3LEnkeAH4BxPvN+llSrD6r
ssNt5nW7dKar0J8CH3YtO0D+1RnQjkbuPoT4VZ+m+/5t64NygQkc+fHZ74XDx7vXQ1D7GYFqxhOd
xJPHCN2H8Icj41Mndt0HT6iOPoVu5t7t56QjswjIj4rJnAuI2HVHlogUSmihUUnwlYD8oHnD2cs3
qT6P0GSe4LWX6/jxYoDB6pNNtOO6+bK4xqb4IWm01TFkokaK/U0wQaEvKC/2uCFp1bmjAfRUeZvw
YCtB8vClj+olorUvZGfXjcFkhWbraUW1krCU4qc3f2a0ysFl0I3G37GCv9O7bJyguIg+TRLpbzle
kxoWkXPVmppmz/geiS0938XW8AhL7OqOOWczU8lzsyrwYXV3pZnayKo5Y3xBOW8LPZN/aW0XSYR6
LF6qN2645hwZgbbe01lgOVOTSxNedLA0YzO/my9ZwTBfw3F/pPjFXBGNJrdpR0o+2hoBK9GDXQif
VTMvlYKSUG3ubfQpV2Wt2Ic0pW74NfIXB8IRex8qVtbVZY0NxnwYl6ESFeAPU9v6DB1YErHUDkBW
HSVwA8iTZ9mR0P1BuQSGcmxmSCgl8eYWMJn3dhQleVxFLATyaXrFtptcwTlkQDKwec2FrcbruYLW
IvPPi6OAyHUp9o1VR4k9JMTb8ox5UzelT4KnEPz+m/aBZWxb7RYt5ECfR1b1IN+C3QRWO4jIzIvW
LgT/f6LADcWsVOVunOLb3eoMex15E1GfFDEXRYTHfkxcR7G4lzxLLbLxMqYrAzj4KchuXmbF/Yc8
j8fY+skLkX6iygtBOX/SsNp6LBMp0UCJB3heBrIzKMfb+NlkHvM0AErjbPBv441nhmvnyUdv4DEF
WjUPq+sRcT4lyUDhclkJvReR7cAjobgNBjPc+Xci5erpPG5L87y/QnjAdfFR2o16SOr8NQDsWnq3
ASAUccK+W08eT8X1W7WhtZdphOriu0EwkKXlCz2hJF3n1dH5cA2CyOBcjQRlAVI9R98heZ5Du/CB
W9b7b3B04krpPCNggQqx+CgoDcdjgyfBjKiXpYUZFJIXRbGOgnUjsNALWpEkZyxSsQLLMlmcl7u+
ccEhWF5Wq08DPMYew0SQHN0GN6obE0zV/2oqCoUFc+npyrIk6ULXZ3awIAnRAtxfPC08Ntmg9O7y
Uw4k7p8OIR4YPZ0aSkJGe3J83h7b6Z698N3GWghuqIR0Xqm/G7s7eRUaujsiuPlaWZblRe3Wpui4
5AjLcyCTeOjRe38zrpYP61S9LHOKlw1xL0eWrVTFCiFSq5hP5qY5as8oWWcg73EabNvo7++1gG2u
nxkpuO1vrO5h5emCF3OwvlBUDXmRCK3/1vU6XpifBVr7nSCurh0BiP/oSmjbMK/dYXU+ufbC911L
nrbI76f71CyY7PhsB9QE2vxmABx1fScTxbOmqip+vbkxAs5s7aPXEkiXuqZvolxEThVFMPSxxLdK
C9nJWfQ2YWUM0XT6xX/NZT0veUUNLNnypQJktc7SaPT1MQuYV+bg5STrpUT6lS9yKhZgrMiPXLzF
BZ8fEu+PQke465/naInoCZRpXDGPonmFSHk2GeCqZg0LxR0UhUGgPqlXoFCxaLpJSnrnDY8sIMsq
XMRvLyKfDsy8Zva9duu2tcjs94xsFuaPwgY7W/t2tWWiEXTT9kAd9Rz+iKsj2Wx9pd52RIAPD/qd
vekTXRRFrpGpIWZ4oiRV5KgHz2gTAeO+VqfGGfk+OMN76/7synTua4gjVfoJk3MmUlKOtNFA3aA6
Wf74p3Km7Ijcj8fUuO01ZR+fT6sulnwA3WadKFNIilnYq4IYCDVDJv9K4deyIot0IjqlcnseFpIF
F198TBS18waDQF/DIU4Ttzzx/H4Ho9Iqc+cA1MQuFoRsy3V7pHTVkFTfOYjuasj0b4sI4GbS5aVD
VtEKBUZVFhDnF4L5k+ZRWrNlHq7VPWLkHZ6nKn18/dPpHSf5ZynT80mjreRUIjKAdMbuGHIUz4UY
H/xY772PFKvxQGCnVizArw8RYqOFqotzZEtyI1PMXu9VaLanVE8SzCPfgSPhLg6ybTNvCu7YxKXj
Gug6IDqiDICreXf6DF9uvCFpAFIK9CYXOPQBEtRNzC+E3/AAAlTun1NUp7iMwd22GTKoV9TEQMcg
UyUZ+8+AzF0eUslAiITuMoggW/SbWcn2Hugkg702fF/XZkdGnjgojwyRsmz9V3M9V51cOTJjwqln
4jY5pNZXywSmTjnNSxGfXHTR/rYCKF5ALOALxjz7lnEowamI7lgySyar8Hk7sWf72rEeB2P9IWKt
S1xi7YT9ub9wFVMVfkKRfcSO3RDCXJzH+gj0Vx+wr619z3dt4BjoRxIXIbezHkdNyEn4gbNkUPT6
WtiXVGPeJ/aVmk3lfeda8XdF5yU43d5o6MT5dwTrDD1PoVQNNhOwgPlOptOFcl6Zc8vyKgJ4hbnh
+uLz+tDlPZY+AS8Rkh/0QpAQx64eeqD65a1/nRlwbcYoQlaTTUmGrcDq22U0ljw29YyN6pRnFR1h
B+Fle4DeX3LscNNyeJg0QxD9iYXH8N1zJV6kA7dEM3DdMmMuKRQ7xVX+4aWSEmH+sEi+NO5HjxOP
/hIWV5T5rDaafMqo1nIRa+QDQ4F5R71siRtyUPrrKtdkdczawIKm7EbQrq42qeZ9mW/mcUTZH3ZL
EjynSAdw5Xd4XwBom7bIJHA0w/CzxmNJPGIamxF2wgfQsDFXVNVqpzHK46icEHqk+Ua9SAoDuKmt
ddT7jukVk0LAFWTPfhy+utNclJKwW8gIjpAHBMkNVl35LE5+Q9etwyIg0Y/xHwhslzXUU70dPdNw
lq311bAQCG+oSC0aAcNJNxlKAIPUIC65hYgUljn/AyEqB742HVqjgVMKzpceZN0/huV12ySgz/tB
zQ8VL4vP/Y+8yb1qrycN0I0Vpe/5589ODeT0S/khUdEbrql3oX/DOS9rao16his+frIg0CgUYKPu
yPNPVPKU1oOFjOvv4LJE2U1eqZv3g/zdNg7qC2TkN5Xw/JvmVFk9CUOExltLUBU5+Zj42xYzEV9z
Ov3lIIkObrud8tuNT9xFnZ2DFqOAuYqPapkvWdPnLWbs3wml6L0Qsv4d0MKB6XhR6xOQPWTtuITV
BOzwhTNvuS6fSe1THiUE0Pe2YrqJGHM7siVKI+rgUCjR5y6pWEBpYCRRN7M51qm+pzi83OFi4bqp
KlE7WF9nnW4jCx4K5ccyCSRRHunXuI7gWB5g89yAMfl6NZ6mY+Ffmro8Qho/us3ynawr38+j2fc6
SuB4R/UsDdTwdNQj1KrzGs+iCqTRhGXdXu1h3bcNZX4N4dyRcaOW+GaAV3cErMHkB4+5Q+ddcu7k
+jj+s4MiR6SF26A8P2DuJsTbg4xW8mYuXFg0cmaX73qfThmLdgtOB4/Xd+Xka84ZFRn1ovbyLhL8
Pfs4aIFsfSLCrZhxmGLTvKmwN95xqV+f0PEK6UcNj0xgdvuMSWlpdAgt9uSouP2srTJN/UfSutwI
9s79TRV2EemKdv90PUK3Pay49MA0T8XvK0Fnb3ldjaFFC43C3WSMN896j4f4x5JWpvujEF2iL7hL
uLfVUSL76Y+KYsrNbIgdi4DLxE4oLmAAir5Ho/J8QrYE5pOZNj700AfHwrlwJcv0FBs8pzcVtg3z
Yq/tCE/qKVhb0TRcRv/8azpWpxnuN5hMgPiKSpz4mulyilAjZU2kBc8jCKayowHn7o3rda1x+5rO
q5cwZnsCP7j3YCDVRpSmq7/T3d9lIFWYwILCuC8BLM8esHjlW/98WDkHbs3KEbkKKEVXtuTRbCJw
4VQRuzxYSPhxFVuzowywMUxEQrfrwOUTjZO2RwsOtbljXZ0JLMKgEg2aJZLxJSFsBmHDo24l3ggK
qaZnzXunELeEUGvFm/BbbbbNDiqJFxfYf31h0qGCMMmpZdj/hDkiZVlNxj4doxgqZVAxFMAgRQhC
hIcuNqFu989V8zgI4vUmynJJ838P5eManYzU1Rr1doxNUuPLokYb7Ag1Z0yoq8CEJqxStSnvs2Qf
IBePA+WVxjjjLIKtaGJPrLFJcYMOrDsVpulw0Pc1rg27JTmVRoBcrbSxp1YWkKqmyQ6KExsLA7OP
64EeLUILrcUvOh6VpPfnu2DI50P1vCC2JU/qYF8ucvjIt/envmj/beNstj76dyj1z3A2Yubq5UQ1
8c2YyKg/SzezcviAo//f2bd+fnRcniHXqzTM/2IUQpdmzM6CTJT8I31F7r/r0Jr1h3dTPGQJPhPF
iaW2ga2fWE6CriT0Gqb+sd9LJC65zr96BnEdVt+KE6IyXC6gfpVUIIxYZAXbKDLROGSaGApIWAR8
ylP7wy9HLi+2tPfVC0CzazDFJTDJ7H3V2M7eDh7f/t59ebid8FoWr320mfPH0ltcZfXN5phE372Y
6yEyBNjdm2LYlKfHCdVJXh92xSzljpd5824H/3A8HKKHUHo+A/V8ZOb8xP7knfZWaRyqZSA5x2oW
9/VOV1mVYmL27zKi1FE6roREgoQaBmG9S1LvgIprIGb7tI5BXOu9CwU9d7XD2GVLJjDGM8hx7odu
b/YFLC71sDQMmZB9+suuCLzMgCWYT0JLP85/JFv9QR8KH44YoKMuzRL4/GsYT55w4hNX84nl0IaC
U4A/q/1ENrUjBmp65qvlTlGAD7w3IdtNZENrEMBdWO11vIVhxSvqahl8uIV/1feGk47OQDXFojGx
VxIt0jLV6mxSebkNwI2gucO/zaKIMg6pF+9KGi6oFGgEBACBnlOfHU5GKf0CxCHe5SrGt0g6WgXD
9XHSiRQwCkDERFRe4QwEJ/H7EsoYyb/Ieyk5aVNSQ//jwByzkbhp6WRY4wo/ALW0l3d02ESkpq6T
PzF8GLABaqs72knKsom/1svvQmcU/kHLuBH0qa/c6c6uUwJDQ5uAwZnzpj8LBZSnF5QOlW4m8Dyt
IMX0rIqdqMIF1r8s/AgARkRnzWwbq/KjQv739K716ztulZG7b8yU2pl1xeowNshxDhB5ewVymen3
DWNw9F1vi5TBL3h0l34/JV8QEBj2dAmRLWe4oCStpDyonQrH79bo2SLlJAJqSvWldm6K725/+Y3X
vwarVmFOOj7mCckN3/kLWsCbUuAIxAinCULp9Gg/Adu+O3VGS2Ip4QdYm1zl5e4WOMSzAyGCgDcR
sbtWfj7HtXvUgfu5aHolIFS8FoOG5La2LXN/UAwDJKmB966eaf0Gdlp9uOsuKCLJ9s6LzDdeuoPR
5ypgFcFdxlcGjrpkZ0va/+elNHHsIN6MXxiv+EVSXz4KCw3tBsZ0B+oZEXf0Ikemoh+xGFYrXpNe
2Vj2+i/SLiyh75aFlPswPEiHme+cJ0SukqJyJ2FZ0u/DWEJ3AYaPAxbcDdKOwnVHNVrYJAzfdfDZ
6PqQTJ/fAdEkA5PmtBSIZhdwQd8ZhVXEtPRdox6k3M8B9H6doooCxsFRe1uif/ILw2mgBbxQewxp
xJAkHlraf1NGSHcRke2hleFcDj9fBFJW6aM4D1oBDTkoBlvqM1R0neNkdwOOcx2E+Qf8Rc7MjRCj
Oyv7DvRZfotWi1rrTsDciFBseqVHIRxsRTEYl9BOnSzO4ogF4ovGP5R+uFDZY5yL5QOQ582Ru23M
/ZqByn8opj4/YZPjHvE4t+LfIIWHL16M4ToIKAupwoa2UU5mVHZW89+2wl0syCnSdm0/2VE8lDOq
eH/0spWOIXcFE9Au0n4y3IoSMTc2GvODVF4UgLGVn8lbV6k/ixDo+3thcG4LyOzM10njNa7wK9Hz
YkBhhyz4G7xKsDGSx0YofptGB97ciSObnDXdTQV588kqP+G52cUWI/v7N9Or2yRvctwfV/fpsXWU
ZtacE+a2Ga9BokzXZmr3PtGFBBsfUWhGNDj6ZB8aIWrhbh4/rKww5HAyA9Fis++kKOKNqXpClq6D
QOoWFMSoW2aA93oCqkpL/UezQ5qIcTk7+ObsOeCBUe4sTNyrdASHLqS4oWJt1Ri6FOY6kGkQGwz0
F3JulTFOWdYBvJI44aRsxzBDhXQO6UY4QjnQllSPXaPaIwU9CDrxIWRo7bYnW5Y8HO51zIMUNPpE
2lA22p7tqyri/X24GJnYXZL6KTAPxgPbX+V45UPXU0eA7+aexWWVG7+qBBWdv61QaQe802k572f6
2a4dJEYSvYKdGR5bVKAKv/5sLsHBwDbDhzs+erUw4pIK+CET6D3Ac13rvEgw/XZvYReu2bjKRRoM
DOln+sv1tJuROU5xlx28+A9we1zKk7bNOiJyJh1TZ2pN9+Fk7NEUvYvBcNHituNAH1RxPpoLVERP
V/xRJLv590rPuSWemQHTL6p1BZ6/TFCo7ZleKUrXjQAVENx7BNe10Jb7yyyyN3uKzxraGEQzMhRm
MxkvneSTte11jU/Dc9ZJf8P/7KeHH7ABcU0tpPSLccy6dqxjWtxglh1G+pIFFZXgYbD87AkCPAIE
zvEkHVIwkjtH+ns88ZRNP5RBwQAkCz6o+qH1YNYnjKKvBeyTguwVLpN3zPeQFJz8AHLiQw3WBEaS
VXUG6mM8qKR9mKeNLR9limbJ5TmtZoH+atcqy/wlCt8tKdEXKQ3DjvDdaQxKlvqRVFoLFlQe0/Xe
jP0Qf+A6DcmqoeiTnXe6k4+QA8+OMT8FA4RgbLBbKPrIrfeyMXtyXAxE1GzXpmR8tLG+/tSStaah
53qjA8R1CfdSrb6a6VcU7lFyF3ahLb0qvMBEn9tCTptCz5gvLmt/1paBkULTqKGl7SU7u/iMy0Tm
6BotvWHkJgez5VUws96gGiuZ8vWVv8NSqLSFCoN6ElFSU6RxV8JygNXKGZCoNnYdTSyuJT84cdcT
VDUZDB+GH8htD9tDhpyNDC9s+GwnBp40VLNyp3HqDAMdwWF5SssRU/rE4ps9VCqgwPhTF05gd/lC
382wGk14WcTNcBiAqSgDU2eUD4mcZ5feu8R46cQcNPoQ6/i2YRua4oCpA0/quTx8xH7c3dCvar0y
DKFqi/mglvBag4SQ/9szMqy2PeqTv6iNSaBeI/oS/zvLVvbN6OL9aw03MGovpXHb/aKHPG6doDUp
vS7ejpDdLasW5IMecTgLcg34tUA/r7C74mYmyJCSUqIpty4HlWZSoUBaximtGNCPLg2pZblADC4g
hnqmvvJCzHS6QYpcjGbNGF0plwaEzcEzN5sKSMZuvUqpTM1mpUkHP/6EBM5MNXfocmEbYmhViA0v
KmZfk/FYTLL1NdpVvOMco/iDhrluFQKopBRcWnQnK36c7zHD87NZEkwowcXNlc9I+ETy4++1rKBm
3NHTkh7/ao4FyH1FvC3SRoonAF5z/f2eOHUBAXnLDWSbXR8lPoEY+g9XmNXFpB3Q9SL5AwCln3zT
HaGpvCKK0okf1EcAqT5aQZUxqodKdscNNwjQue5XZVtLaU20v8VDuhdonFXNT96JdIDdu9dQLAxd
DaMVtJwZziw8i0WJSBq+Hh3EsoqkyXW03iGsArjC/0fhdnGk6n6chXQ0gV91f1zdiCD6BQbo4tGs
Eyk1bkJPqLcBroL+gRSaQID2+ciNV1I6B+09RuE0535qWsEEEGx6fiPfa52VRaQ3cOMYcn2cEmPr
mPJ0r5P2LoPaJNh0H1vjcrljke09xwLU3phWsc6ncNhnDZn7DV+LjAoi1scaLkQMRmiaOJMRY7Ff
/7slV62gvVPj8Kr895GpYpUb36ihfKZMOHUOdywIN5y0420BNzfdzx5iqrnFzQbVObvFpU4KC/An
m8xWIVe+UHmWhrestwqKW5M/66LaxPP48cIAww+wRhrFcV4lOotgzva8ZwChn5r3CFXfq9fgA9ma
VbUPHMLqY109jFsdu5imCLpSAYBCdKQDbJ/afbeut5jWqb3Rn2BVsy6FUMAVOXXKyMxdLmlXvFSh
0xtHukeF1XwhMQDtf0gXE2S5qYi5A/m78zEGsZN2HmMQ4G7kuT+DfsJX/C3hzMDe6pks2nCGGFf3
/OLjz78YGf+QPyBzzmIMRx97PWlasMAtA1bj0jKbLTEjYEODYy7XJvk1xWbDVH2cfMI/OgmuHuJz
148b59xdwj8dH8YxY0wAhYj5XVhSB8PV85s38e3jg9yFv4bKsokNDY6lAeGCnJoBGTm1KpZ9NsAD
EwbzHUQ7GI4hREbj92Q/BbY/YUqA7ItxSBE7f+wilnn/tEqn4SoXoVFN1CYCNAsyZ4gWXFgwk2/1
5t+1oZ1oiocs6P/bCZS1/KINg1cdhOI6PuLXAMxBb/Kd5YkAM3Il2mTDDIuYJG1HwqK2GKM2gWIW
YbezE1Axtz497k2VD58Gt6GOxRjQLMnI5aHrksXNCAGFEKHferGpkiaroqcwIdwq4RP9DCdNl+Sr
EB+7e/Kl81KAmBWw1IHmeB7Exy+4WfyF4j/3ljGtfvvIWwrN9vaJytFSf9t3XdfF2fr7zCKYOdrS
v4/q+71nUKPLu1jl3NqM7KdarucTR710F6AHGT5uT1tkIEN1unnP9U0u1EMDnaApAoJlv/LCrlD8
Ryg6KMQmSkodBoRrq9z+3hvp5NPpACw4Ds0Yrsjt803oly+Z1/lFQvrqQyXhLd0wC2ZI1zM7ATXi
mnp1pnEh3vN1hIDu+uaCANHkPWH4U/BLMKVITWQvyasfbapp4F5cR6JdM7xpdRy/25+gBY+EzvKa
zcbsK70VuFIYeWj565oIIfkQgXtOqAyEOxpdeSQuraNdMfMnfmvYUCbzrOiBo5e3l0SBDqCF0fA0
3fxQ6jeJddyU9dCSrq8AkJkfnzMWXU7GJ2kyw10mCDpMfdovC7+37w9gC5g4CUC3tltHC81V+VmE
uS2bpptBtXenME7eqstuecd2neqvRwmzOqn4K4YMeAm2Ndpn2fsWugPrx7TsrX3PTM8Otjha1u7J
Uj2oypnPxzXmW5oyUbK4kuFakVtaHjMa0Q0oRpb/nDe1xBQk8eQOS/qqFyL4Z4QCi1p0BdzXpwun
jlyNYfn3WvCOM80Uz/qtj2poriOrQF2ZVBPMUTNa8rVZoKXGgMLxUq0CUz/VtJyqwNFGLP7GpqiH
pDNmc5wpTGaCCLZi8RwI9Wwcs+72JH31BPOw3jH90hS/bAfbo0hzzep++KY61oLNj1kRp1R8bbyd
QaFvrdYUcjCqtYVTGbJJoqoM8mD7thxFESqmgGLeGO+xPGdS3+GVT3Oufc2KtZYXsyGUQVO3Ti94
EgFgWHJIHibGjs8Y1xbHjOT1/WJRRzwCiWLHYsPtH0PqA/EwoS3NN3amenV/5MTgIiyj3dX9S2AO
jyqGJHINslgL3GB/KOGFCo/m7VYvRAI1LnBdxeOAMAPs08n7NmcFaGDPKecFsqZsrtTKfM27m5kI
kwu3aY0QXSWzYNCtuUpFFkXwD/nQSI4JqoR2cRsCDofnYRxC/A8cyDLZOgzTdvfFWTNanuZ6bbLV
FakuK3ZACSX5mP3fRFxV++e5BjgjxeluQNDMw5/2UsVV+CVcYBc2fyO/OadOfgi/gDMXovE/nu+P
3rWmKNW0SjOaUMQeNrIs7jZ6ZR0ln2lQ9DVLvWfr5y90zEh3ZEh88sTW7kzbnSSGSA8EtPIqLg6B
hr1rEXNno38/QDyEk3UfDBR17KnCV5tYpBnrIvlFxEG9pkzp97ksCKCPxxqsuQnmeBhS3TH6Z/HW
98du0l9T5GAGch7WuNy1QfO52GI7xM6I0uMg65N600eEzBCLtGgRf8z4rEs2cg3LCdovShzAV5V2
jjtZLU5THo1EmDvUefdRDuIbxTmmGToXiaoEJPUkRMPdYHM96j++RXuAjPQPH4/i3n92zA3GiTAy
zy5sVXuOQ4NKjLS/LOggVGpeygNKia+Bn3R6nrYmR/msJ1fRPzL1umEFvXtxyK8VR4Gppash5TTr
11nLXWOjJJ8O47uwTT6oId2CGMB2B6/6bxBjxA1e8G34RUlquTH2yfum+A/AZvVi7kq1jZLpDIBv
xXm4r0q0u7VgP5jcwarDLJZpWWXyAh/f1kkOIvxDw5SynQ75j+OgnHrvyjCdQ7sG6GtXd8z0Dmrl
AeZFAp0DQZpZVRGQsoGBI/k+X2cl8UQwAU0x9Gva9Ir5XQLWqBeNHAFMSOtAQ20zxINKvVL48+s7
4XpScqqcyVmn3Sid98xUhDxeCmYfzS/RP7cvoKEgJhulmKPfLCy/wEoMLK3yEWLAniBUxRnPXLA2
1KCJp0iBQ0RFOVsOhxhvAIUukSnPRXrWz5HqkT/3fpTsG9RH3DiD9Wlkqt85Uwn2Ohvditr9Uf2W
vqjnBJAtoUfL4gcjo+DZNM+gNiDdRiyRTMz9Fde0XAjh6Zn8f8f/jRnVXp1hbb9dLb+Os5YKVyXE
2pHELlk7t79JBfXI9WcSAxkzs2OVXdRMfyE5oEEJbyV9a8X4SQ+IgaAjFxQCCgZwFM9Re/5GiX3/
FTzIlHQbnKOByLMr/ziKRpWDvdwgrkq0eBwjSwjF3NUvqDZUp2NqRMgJcr5r0sRA8PXyeJjCDIi5
73JxPjyXcXCvbbF7QfbubolF+NL1R7/8RH7VtwKoo08Fj0m4ak5Ll8BE/sD8A/hUmphDRLoZsk1H
oHiG2C6/OxIQ9o5GcDcM94/Mcusciw8gkIwBILnrumgl964m8W5cgz4tPWbCExOZnLKvWkt03+i4
Lkr1rqv2O8gq9Wt3FfBjXXmkgryuTGhYpNbd0uTfyqEiUCDU1XpImsCPu+58tbJZR6lg4S//E26r
ciGZRQ/udv0ddFCqv0DYPzdL9z9JDZx2WnTQvMSpWbn2O476qmncTkdDK8y5qPGPUTG92N7wugYZ
9aPh54JSUnD/pum5FgGbBRsLog6iAQMatJaA6uyf7S8xwNUG3YOYkMUchXEtyDLkZseA0HS6YvIA
0ctXSWusk2zd3u6P1Oo51NwwgCcW7tMSbbw/nCHDXT4v82hCydu5DPFnIGpy3mnac6/qC0wqdKnb
ac7t8QribfoNdXOpFz7OMU2okCUlTlxKgryGbInXiu3vkFF2iz5s/k1PPIhwW++QCvHccXQ88YcY
YgVOGYeGrRpaRuNn0Fq9Ux6GR5WHV+M1fNloiFBPE8TQYEEIX6b+PQ3ehBF7VH2Mm1CHstePhIdi
dRUpfZeJ5T2Kjm7N8zFgiuPtJmTTXlZIVcarAT4B5j7nT6xc9XpjPQRJgcci+jWD1l+mlpT3SruW
JKRaHFQEqrJ97uQmZu08lXhJbFglfseLZQPlL4Ukqblu4eP1j0h9pLame0DDjyq/RuwWtVtgD4xR
tKCp8cnP68w39oMeVkl1SfFzWzTb4adLFBsW2Y8yj85M9798/3J+0Q+CGQXpdwXH5VoiTUSiHXky
NGN4G0EAgM9oWxYnUw9IbnioDPkz0/76ev9RENyZoW2PqA4B8G4sd/YGGEXy9OXnJ3P4KCJ+/hSv
7E04F2/gYAsnmuuNetZ5untL27jkJQ0gR6Cv/vzzu/DTkxbT4UxOwB2kk68PnJqDiN8JY2AJyslz
t9bxZ+nk4BuOClzzff5ONCkfc2vhqGXM0fZ1zkxm2RJaQRSk4Rzp8/ZhX8FXBBg8p/XN/anQnHN0
nisLiUJeONnvn9nBzjUa/9IbmRq6Ht4XOSflf2H7sEyiDleqhNJGfnADQqR+RycLNQzozf6Zqvht
vHQpm5d5mQ8RkSNk/oqE4g1OJebfoQNWiUikYIrPDR1xuIUCa/iYa50CO/0IhqPEadL5BK0rkBNd
w9HZ3eK4nw94BD3fR2/chiqdRUQ918jt4MZ1WKM5AmWhyewaWW/B64DhXpSlGyNA7oViFWRUn2+d
T+dIWyrgyO9uvdneyV8ZH9YinAZ/0mQpg3hzx7CQaXisMggMOccs+fEimYf17jNJaghcb0kxC0ih
JXpFG9NKKHv3VX6dnMvOaX90homzE/lRci+FUdj5FtEiKURpyy3Uil6zioF7SjypgXsNYjOaaeRW
bdewsDFwbQrLUml4F61PWT83WXJdMjFJnCISR/UCHBxx07Kcp9IVT5ryA6ymUuTQ/AwYJtAASXv6
q0A2jwggxs32X72IaIJQyQbvMwEHaNbia02KnXsJxfBmKWAXg8eXG6PmOoswrRe09AKMzpbQl8Iw
08+vkiERVIWxy62/UBJ5QFJA9LiTACrupE25FI2Z50MNq+MKdJo0aqubBfQ6ZHSvcoWmCmZRvcsD
7fM5mrvO5YD/m/7DU76oHGNB1+JH72jFuIdr+4cR126aWwqRAAHRG8dC2O+jlXxghfsr6yqvhhwN
xDeEg3k47GBlyDyW0htNq+Nc1yclAiYA1aYCRCtpL7adHzK+PTpfpdc3X+L4Te3KsDZj/DxKiyZp
3Bc7S2UPi7peO59VyDC3NMQxN+LnBuJB2Rt8AKMD6+z92YKJ+SBf+DRrAS6WOFCFdBOZOmxO/Ww9
JM8jzNhkfM4w9gSfBNIxl/eebll1yaO/f/G5SZ/xT1+KrkRr9xJAeAgcu0LAhqPRX+rv5yx87khh
o5IR7YoerQeeY9di9KtDIY1TYHkdYoaQ6SpuLul4ZUhBc1XZIStFaaZp9ikwReEsZoLxtVQKmeTN
3r+OwSRmnuk0y1eXMLhu5vH3tx7gRWN0gKQi362zBnLd97dEiIce9ZCHSf6CV2Bkiz5ndnkamA+e
/+HD52OoEkqxYTz/u4fEjygeu6irLb+Hs8TUQxJfrgIlr3J5xe7XCHmUKad+39QvVuo5bMAv6RBd
QFif+KNxbfFiFyEiSBGbvo10cHdvZIP8a1gySvei0eYf42HrOc+sr7BLEpeoJQ+XK7OKgAtNNr2G
3bhIE/AIn5G5DgvecYqC7tr8xVKi27o2z3+vOIoZNgEOewG5yTIydKkC+iCfk9P0d/pILRPsIU/W
acaXMwX5kznPzsG6XabfK4pSIkiN2XqEmzhgytliZQ3ObZqRnytn0/VIo1Zs19JmQwZH2uVbRb0f
ljR/R3gBChWGrBfYwvFSgjPsAjs+JdYgeo7SJ3yHwSVytv/MwdB6xqObp9FDmfvY+9hQ7dyBrX1R
ENHRvRHgyNFJrJy95A//g02RMsvd4ZqhF+Nm+SKenXsZbovRPVa3DHdEhBdJtqWK29nJ/hZbv9cv
x5gxO83dF93B02hd2FMudUa4fhxoVqJakEwqU78xQqgclv5gPeZyGOL4Ojv4ctchcf9bqg0Q4H0v
2PbNoDUKfrW0JiOnRg3SkKEieUHmHPAFnra1CpJ4WJz+YCv7cAqKsZ+A401cyaUAm30P0rmNPy4U
qdGFPJOC6awwXe8Xq0jNBgdg2GkOM0AdsLDK4IYg0BdyV+O6UC3oHCom0h8OwfO6hfSBKnD1Gt6x
WNU3FDvBXHuLuXa/YKg2i9PvLmnbce9L0GCNVSr2lq18bQRexr3WPAb+rOXZ0kddJh40wRp5J3bd
4b/Dj3lEpvS3Q6pOlMvKHznlmUBNdJrT9VFxUNtKdR8ErjGIzo2O22F/PX/1MIXg2wK7Dml1yRF5
hzvv9pkpnc33iNFH961z0BTrBc+09bpeysvK3HoxhAmFhvoefNEt8gQ/VSlRaOgfzA0fu4qmu6hr
yd0J10nmbW7KbS2L0VSj74LOWW2nx/BgADcLIvRAeyMwZRtv+KMo/+k+AN1TAp0ctmnsJa2nYE1W
2y5b4oLpprQK3KpzilTVOGFYIvekIFoUswN0ac8FKCUBb04+KLsuGBF1q7LBHrUuJyB6ccPgCow4
xxeQu1XABqsb2efD7qrvALDUD3ilFqebhzCoCoiDBTuzNk9lIcxDyheaCkJaEhT/wxWRtlDg55Ip
i9fiDnRchsSnqhOCXawH1rzEgfRRSum4Tla+BYGvjY+/4RdWfeRT/I/90+lH1iCGTLt4AnkXH8pS
cc0k0v5eGpqILxPGNNAJHPU/xg/iE7OQokGSb/9L94RJbs/12I1lEj+PgdDAzzv77u/0jqpSVYEu
zRen2hidWdvmk7jBZz67RV6A4Lv4i1clJFsuZfOPl7IKP7UT5wJge6/u5T1CvbVt8iQlBSTeg84y
61tStAJ0y/4qobWo49io2KcnbexE3iPLwSM6HnF2+i4uyRjK/MjkXI3U3ZPmXSoL0p7IwHOOKxzF
E4ed+7V82MLKSqxQSHjstcxq9LzUJXHR3zJwbEet5/qHoT7HBYKv0G1NJivu5mlyyrJL0QgrzXcV
jTAstC2jArM1q9AZlVRZ4MPWPc21QsHJ+MjepRm4i08wQlsT7FeY/DyueXEjR3Rzjc/g747NgpAO
QuBJ0D49Nepwi0PSkGjMe3DjSMkyHQFFOyQ5IFEhoBWK0gor2fmwHTbiauECXkRevqy5tN1eRQ3G
WZ5QoSsfX1oJJxllK77w88iam7IyTvmaEoo2Bn6ENrISDuTI6uOPVFYvdnw9HCizHaItC9KQu0LO
dY4jtVrKWElMlJ1Lnzg9RUforJbZljknmWi1R+Pig7wC+XgJe6RZOheC6qUzDe8HRIFystHka6kH
iL4LFetkF7HsOqA1vMdjZYZen4pO6OhUV/4s7yG4iRQEh6loAtVJRJ9SyKBr2p+AiPoBhc8dmxQd
Q6w6AMM9IoX1LkAR7HfyLGvozIJL/O1eEmVD1xt3JEN9JHN8bwkJ4Rux1qKlEfmZbsdwU0/4RDl3
GhIfK2Yqk7ci5RawCRFHPTZ+ei15IOr+Rqr0rZdwxyDEGlK1NoaTDyM9CJLS7sg5pHamsOw2eDIN
T5bwbM7FeZa2PnFmssNrTcDY3086uIABN7JPPC76g6Qs5NM6k29+9Z8WN1sWFLa1YlbgkjdJxWX7
ndH9rObpQIe7Ttr5WCTmKylsEXwbgxYnyvv1Tz6BY3XtFyIfuy0AqgOgguWdiLTu6e+8Sy1eEyfd
7+Pk0l8zdm6SqMjpKR2m78lON/24m2Y3eh8tl1TJ9ggQtEFygpqaMFfM3mUOb+rNaO9pWr9plT7p
U31WgR73Lnk2cejYeYZdL2tJjoqssjAX+NnADdOfAkwEKJFWY5PLr/MBg1Q7KtwSjGiop8t2XDUa
1A70QcKEibwsl6sq8LQ/THNYqc9ePRNx6+iwysRTjx9Th/gNS36wDQ9o3lrkBnmqfiDbEs+R8ZCp
Uw2g6EKx1ckkisVGFHSg0SQrnks9vu4wJwTSjgD17J8i3wmDq0NXTZG9VNQrd3TT0btPMx6j8YPc
o43biE0eNwpdF3PoaVBKo9lDW0FpFgQ6dQhs2lMR7dJvXMI2h/2ZUb0uCi2DEn6YY1WQJZdwEyNA
CbCPnGCP0HY7jOGJ6kXBnIgxDF/SwTk8VChUvOc8xWpLNK90wCmanFnQDzBB/LKVUCw7gIdjKmJH
Niw/EnSU7tDGPar/6xEJDqhAEFRYXtgr/5lZRGDWRuYxHqRiBGfGDYHCYfUDWeQdQHfahUQ8Itr+
CZunR9UZ4qY0hkAXGkasXWYS1rd2hGTgSjTr+fqdeMslrzVC0wSxVstNObphppVEQQjej7nUfrFr
L7a55DvDSFQyKgut1spwGsyzAC3XBUn1CIp14mr161NmzFJ4O0QcOtFWN5GFFVOEuQxrFDoCy6lY
j5OWyArvf2BBjdkb/oOK4dx0I2x/D9g0FTiUwrLl+d8ojVJvQlFljMThNQ0B4zNo3ioHCi2zJXkw
682UOV1RofMoro5ac0U4+qZt8WXNNNSmykAdazMeJiwK3AOVPxJ3kIuVeRcm20fkd+zSeCVDdfp8
g/Vkek5SAW17+E7Q1Z4bYnQ90Nvkiv/9WXe4OBnCTfHrthiTTlsFAAZw84tnn2FtLN1X8sm7G7C8
cpplCz1YOXmcujQvWPiK7kOPkE5g+sLgi3IfR6/0Cr1/FB4HuUIw7ecUV63XckmfA9PvYTswswxw
gqZB2dpkq+mCh4pAooAddaMXBLFRh7YNUDfYp1Ui4iSUmPQRsf/RmrP69yjtMeDdrICilEJSaCc+
Pe5m5mFkmvVftVKxFS4CeuPjukD/WBGCaAhueiBhMiiZq9GvV93svG1eq1r6tNlunReEDbkEB6F4
+KB772kNapquvf5m9aGdja8R/dmjfiIL4wqkwmfRMxJ7CjeSRk7wpElvsf1LAS4agzWsJDUc70bd
SuQCqmJ3uBwI8DPTIbCqL9suGzb8wsKAJ8FyoN7FFnPxOYrfyVNzYG2VChADpHCo8G6Jxk5DiXv4
6lENxms26xhdu97T/lD5OPX/QtzcOtr70SC+Cc5sUtZSKvDNKUekop6MAlKdxJlCAFg+CQpcvG7X
BIAKm0jJi8EZPR8ASEh4GOWlan0SpAvXF7w1Tw7E9H/HXA1NcS1gq+wErbyJHz6lMKYL0IWywQTl
AJxnt1uZd1Xy3Q6HP3HeQZ34f7QFwkKUmEfP53OI3V/STaFNkwxX1FhtEt6KfMsEu8yEXdPTxIG7
MQqNigoBPfUObPO49jSkjeL8eUqJ4190Bbhv6i25F41oFk/IrKqeVcwMoJ8jZ5pd458qtDLwNRpI
YlzjABAfv7mhUvaNC17T/X+97RbFOaUQ7dz623H5v/m4g1okkX5ROpZvULnokZZWTp6g/G/cWMm+
HEwBAhAUS9+GewZjFstrg8LNCfoLLUbEBcbyfl6lfRPEUWGRMvHf89zS2i2Sl0BBdBDnwQdID7O9
/3ScUjxGVdWvCIac5LPQeoblgTKiLS8a/qBg6Yt6wo9SNjMcau1dt4i0IKFP8DuC6ZivDd1WbVm0
HMHBeSUT8g3u6RjW/tgIcto4tp3nEZMLoXzrOoThWsymW6szVjNInisghPile0AYS9Rj2pPG/VPU
4yPdyVxIA1jpMyxy+mJH7xNOTGy+J9hV/HNqOOs4+ucCHRKY7uvhsbC4Sc6E4Fs3BMI4+3pAoJug
D9VTAXOtJF9EZN04SnurVE5SMRqrHbC5ByiUbfrzwmHd1uFO8ApOrlByMyZHNEhnN2pF4NYMoxnJ
fCYT4qeK1z0i15/su2ON4fAZ3fOviaeSYr+AYECrDN7jJIaaaOUO04+COgdGIIu32xcVBfRlxGqp
+qFFfPmNVMyqTcN1r7J3FAlCWNPs5FYZp5GvveUc6YaLhqZptwNcHX7WNWk0r8rQ6FwRPrk4FNxv
UWvFGJHUKj1DJFfCZNvczaia/uZu4EQ39q8gGgMmligFb/yOw/tHQRBkpNQ7TivTTJ4zd0rpSATK
nQKcxGLCdg4TsqmBqHlEJQtuLc0nSufUizvVWIbX5fvXTczjC7qoUwLi0cKlr/i++D3oN1IV+oW2
x3h6l2GzEVM3YZW6IouwA6oXhUbGSCGXq3TGMGn2EN/URYNfG6JpL1XV5F9/qW7721bIDmo2IMbJ
q09uOlPMzy/NZJTMn6V48s3a4f9WOp9q0lfgDob0PHPEnIglmiLUsU1UBYu4/egDvVg287nRrHoz
swgTBiyqe53si9k8iUxSXVA6mG6bOQ518pqZ1LXZW1FX3rtNXi/zuOfDZdgioI+WplkNKSbKDToP
MglN1ES0ZXseyas2/+d2pxxxwc+8xtXNmycl1jFW6kZhlwy+endXLVH7k2iSa05nIcgmtOFZYraC
Ax/UHSPsAIhw5ql2P5yL6TTjE1aRwdrdY1AC4Zrumv+VpxAeDqaeC1eGKFbWr4+j/XkjrPkiNCiZ
7L8L5RufRxhUskGBBUYtNe+lZjyieIeizGeXulHteglVgf5w2aVbllIBgphBL3zHBHs1KbVij4ec
39r2wWPE2dEBGIyze50VGmYQ0LF3lYtXq1f05cZZ292VaoD19FwEgYuZAx/FU/7AfItKYMWWuPkz
w2o0QM0KFzZeYLDhbRD6qAbXWbD1zwJIknKFzmYu+iC+Gyb+hFxHm8Eu3uqFtWU34FC0hPWFOTHb
z9WUJ1EWmJLkGdGE/u5aXOxhItSlBa2diZ6bQuvy5V5TivgI1BC25mKwSyL8L+tNw0LqWnq+5UT6
qYxl6sMZ/S2Ovna26rS+RhMyf7huKwQ4ehkXwVjPh6WT6AxEpm096MomFnFTF/XIjDg/DdaMfIPz
edO7KCdmJSP8itBaiQ1W8GluZB8ETLIyrIbea0MNgDQ6GVUeGyW5fpXG2Bg3aAyLpoQnwqRkHev/
x2/b6jxtfBUj9uz9y6C2+x1R4JvSyjx24fUnArZXugtyvK/UZC6hPdJObnn393EaJe9LpiYw47CZ
HTgt0E+33bvGlBytIKCLYeybRRx6pSDMl4kTn4E43MsNtjwN0H0KUE2LEw9vHG3wD5wKF9LGSV4c
bOPRzt5Af1rURF1xI930/0AWzJArtAEemFOBydTknD9lu4QIRhnMscJtMjwvaFQzOXRF6IQcw2jY
y857dIp755PoHKHY7mxD7MUgBYQDHRGY/EW/5g2g1tehEzR1IuLAlpkhe/dPnI499QEj7MIROxt4
m+qbEhPFM9ah01T/IDtLu8xBL7kkI+14XuIP02zHqKwb+r1pAGqmXDqLHoD1Yw3eI8Hoz7clM2mA
C41JTsxZ4yNL3pl9K5FPoUn64QMhbRTnlOQkJH8Bh+u3OatU3Einjx4aipfhwlkrOILMFk/cAfZZ
Ih/DYvMG0VjXqz4QBtHifBPzPn5eCUV60Lc7awASeZYdH6VsqIBrpY2xkuqga7+8xVb8pCPUzein
SbP56nFW4YaqdRQMSDm5D0gpgaJ1fK7MAkIO5c8EEWKTnXTbBP1IeCmxJlZNhEr5STkeiUvnuzIl
2MrbEwLuRNk4pXz4q6eh2QJGgvU9e+w6ZBceXLq0yOPeUq6Q8rO5MYXOXrjt52Hg+3UB12GxZG8I
6JB77IR/sCdoaaCe/LtRArBnaW5/+iBeJHlezqaArSysPHzzIojApXOha9hG7W5LYfqjwumdgfFq
W6tVyFmDMaOfdM0ZfqjZehFmlGihTowjclN0tzjJObYgFYPFCLiLFZHoOQQny59i1JZqFIaPFCMd
dxGb3RolOmBd/0sZTIJ+7ApQSP/C2eLFi0yFmEeOig72fqLOSznKCsg0398ETFSX8qY+OLXbfar7
9tIxxnVt3DnSC+iUDTL08HEeOt923SEmpLl6IGMVW5VZxQPcc+xDObdnmRI0su3yY8/OlRI4fAQ3
d7lytlghB3tL7xUe/3wtc/4winyFaM0rTXqjdOzVRPgZY9yLuN53saBufd/OQPDCpvvPz+G2ebNT
11xngY+B4iAvxnVWyrQpR2R7ER9dtkawPp9FVtfE2vLVzfHT3/2D3bHVfbPttF5jSMmnQBTAtnd8
AIML8ryOUQSzNvRtdEYOV43+F2ZA3c6KD+/bMuNU9ujAfzkXn+4EJdMMns/eyTJlj7aS2U46iFLn
Y8X8jkyQ2YtZAWj9yts8f7qRf3xx+7X0p+xhVaYVEggDV4y6K3q7OIytNoZUMLQRr6s6RmL6Gtul
+lOYtrlz+IhAIZNlIq7HC6IYJc41pg6xeMAO/bBLUQgau72+2ZjfuiU4s96hwn4+paKlhfqvVrE8
hLf8hle3VH/GUo/vsRF9X11GO8+uh1j3sX0Iruo3iE/dkqKDkZt1VtoYe1RxuZIKg9bUnGphq4oJ
XFcVX9NiXkDOEuYXJEnoQcoI7IJ2jmNnd0+ImNKcbZlIPDbyYx4N7zkNskYhQPHqsaEw06rDbFr3
pCrzIRkyFq8UZXyosDFLSkLxpDxUoQBHsx+gWBAeIhv7FZeL42n3ps39TaC47U3tIopBqbon3Aq/
ccEeHJMZP6UYMNxWH5TFsQGXu3uWr7sUWT7Wwt55yMC+QAvk/ghgx8DYojFKL8z7i7MrLMaO1Jwq
Ux2qnoTAABVMDolruLWl5Uj71IK0IRirbbJtgg4/ooP16LIvzzwEnn0a+dFNkCXO8FFx5+1nJzhl
JGfOwoPKGyMiaz8v6cG6IYpBWPR71rdaOpaUVgeZTOQrBCfN6VEgdKeTbAKAWcChT5prcTfQWcVV
jLb7uMqaIKFoUFB0/eElElxWh3KHMg6k6PDUpZAnjY4MD4PtBXLJo6fKF1D4go/bpnxPnkiFmnOG
ciQIoSxj9Gv3RfGjsjY+fz8/DDQgAI/Y9RPCXhQ1hS/GzTWv38eldrc2tCa2icax/cESaN+qfmLY
afWbvHXl+z4gVvDoTNbQiZ2vByJEyDmES8dO1mLPl6aFGE0+XAmg6OQIbJprIPNts+ywFlH0EdiP
JVqiHprvVqiYZfhS1Bui3QFYw0NNSaTfM314/L7CMFUkAKQ4W2kZcVWE1qLcKa/7mo2/LV6NC6Tb
TlaghDXb/xBi5NtcsMi1L4MYtzfsLKeNq1ocX6YIURwzMMtMBJ5mIlOzL/kPwcUshSPiCl/aUSSE
tQ/t83e2Vn2FP9UCRWjEs4VKS+TzTyUX96P36J38MKRVRND7TkIKcm5C7QZsix49kYQjCWvRK4cG
UuAAuaTc6r1FO6mOveL1by41ak8nHFKRhdSUxg7kd/KNtMm+4UgYFzsQB766ZooDFkmK9Eagd+qa
cwq+ZPVaTWIHaVw+AKkDaSuCMvTkVeesqsasgP/cYGSTJMLeDPzzDC9DzDXLSj94ZFmS5eOLG9zh
QVR3TbKXZXNQvHDp/mpQTRjrRjiOHtjGLa31V/67nL3tZeZv6PgD9ssPLoKPyvtziP31cxbD3bMI
VyV0dcKjbmr9yvhISuOeyJVRI+c47ZtwPV0mIiP6o8U5JGWgyUy7JnK/PkTrzdM3dwgXU/M5jBDS
EGqVHJs++PcB6N3ioU+iOB5YkW1RgkEV5urX2eWuvP+y7fSd4PHMjfo1MR13h4jNvqUmMg4gSAS8
o4B5ErPwgPsRGrUjjNBf5BPZfNhLcBAn1r74fszHskLRR0ptwucEHt0JUJqm9YoQm9jBwL7inryK
DHBOva4VD/FVX9b7LB54c93ribDm0G4yg4OCZnNdh3QA9EubCW1/YiKlEtkFN6e3HvfAlfglZ+gs
UaefTojYup1+4qoTae0nqMGIsJQNm6h+fh0lLIbxmVa5HxUf3e35vCFOBYjen5i4vNnz2Aubm/49
TRo3u8uW+UOr2fsDmttmWb9/vF4nk6z5LYTQiw2ZanC5r99IfdIBrU5MRTnSbZEHy05V4XrJQ/JX
J3HZ+hoPeARY1qCYL/bN7rKxrekKPnl84ysbekieafQIpM4BLHeruviBtW69LvH5jEaBIk3b7+IH
ToP08NFAqsYV4gTygSFGth9yFTrMOJvnr4E/rojNenpCUHIrWuq+FhVoMxZKglNJDO2PXamKP6Uf
YNhkx1wvv5eiUG1eT48R9ma8y0UwXy5CDItLsSE+rVXFV7rMCf3TxNGvjNbCDICZ8f0qnqhJQQqt
l5Zuh5fnOPh8HnTCbDPNvyfG0n5IW4WPxTojBbqkNpJW/vM3F0DNoSEV59ueOCvn5I6/ZwGqIl9Y
8hX20+5XhLgN4Lt7/5RND3UYxcfeBGehRTXYZ/YsnFloz+Gajsdjgul+mzM1z78VCrlaVpPmLGDT
iXRwzgf3S9ivkSu7+9hWjhFLr9KE5pyX7Huv4Qu/5cLurF2sGYC/vfo+ECV+ZYZFkNakeUl/dIbT
Eh+XUMv3rGy1rO5gtrNE9x1taan26ytkAaK8csOE7nnqh9Y02jVInh8h+bbdaCvNRT2ibCICaYqX
1pynxzzyyzy9uWPQLmiUDT1GsawZI8j+jst5SMPlh/FmbTtFan9GJreCQnzwUO1luoah9wGkdid3
gMAntMq0ojY0quICOdwNg17KTe1spdPhdEt4GCUOTVF0rtcfD45JSxYoaS7Oj7xbhtOYOF1mWguW
vVncxlZUD9TthohRSzcbh9pBsS/SaAyHJqgqzAIiqGgdKaNcPh9W3DE/Fhg3d2UDuqGXjLGO8jUN
vZCnmSzjqqBBYqvjeF5a0o7JGMt/RVbNlcovH38TPJDFN+JjQp0AfRxlT4+Trqw80mrYnIbqMrJg
XL+O9sg631CShc+XBJvOVCXrmr0YFswnpOOmiR/O/JzD8MaEq5Pn+RLyQ80acB4PLKn5cO+9bdMg
N78uFReqmhVNCkTQ4QfK1enTqYM2a4nz9lK3ivgGuNOqKcsvXVnrO3R4reQ+oxFqJHwq9S5Haxou
9SB3KM7VYgi+mGXolgPJaZMOVkbNnwiBiqNCykjxgssfnePyYCf+Ev/c8xO6pLyxrfSZ4NSlm8F6
blrbUDXLF3d8u35PPuurXN/Hx0Gvhj6G6EWhPKRsCilAaMbRhRHKm+Tbnq6M0o1wXWIjMI6iV4Lf
cONP6QjOG9aycuqxlnQozehHIpqCl2gP/g6q/2o9W2D/+JMAIQHk08yYJ2lWmyNzZTTr3ZPcd/f7
AObIeL88D5at7intcnB0b9/75ctZkdaioOSeMK17Z6AwW88uyBTh5ynBmPtXXzi1g+iZrQA4CkS5
xEDEyOAhL/Dj8DeIp6aAXIYIE5CFr5DvNYyeoX4XCor718TjN3ciPP1QI57wkZT+0JIbEZX/BQrc
Dm+u4isdzFUPi+0Gxq3YUWQOFfq9n7gkRmXi08yZmmpJvy1mugwjCvqBSQ15BhEYmZl1y+kBz+tD
3bnZ8WTBbDMmmi6xiIYEK3b3pa8V7PQv+pixPxW2zrgHV1f/K4VjV7nKhGTddLh2alXaw8rBqUr3
2c8zWdsfhxnQ4F9smEPFVz/Sx9VS5ABUhMwZ696CBe1MpTnIkC+KpHzENvF2zECoYowi6zcF+q4+
ENevup3DiOyQKYdhV/9QlAsOKBYfil545GKQ8D9VQi4xorDGfFYOwPZ3jKJej01iFRnn+eSxKJOM
jX5ZVpSpW0ucyl6AGcSgXNkXhcZ54mKleqgsXVNP3j/kxxkKGVGM2Hm749vc5va60MWwaoDHkzuV
5eSHhLTFdI+0NgMGAcrElvmF1C9X4UIbf7AYOh2EJF+7UkQ/nUixAOfWyV14k1vbI1EM5mRPRDQY
AxPJuJs2uVGtA1kG+jN2jaLJpJkr+nTxjHc2Am1lIwDgsqM5rMnlR+C4t0XV213WDbPjoxKwqEhz
Oh7epMHFiB6pwxG8WHPG1NcotJ8guAl2jC39fuNp6vlGK0rSl0m1G7W4PXQPuB/ER/zxFaEYZN55
qLhIacMtknw1psjUcN3xQDVWVOurnGya2mhTkSZogQ+fTOuvELtdo/qNxOec1syfMZsaBdjHdyEk
qJh9cdT0wjewo/20VuTQRinPtvWrgjU8G3mnxqcxlH0T4REyO4tDbl7zj8N2ldE+bLORT80HAEfZ
76gMR2HYol4f9aKxlYVFmwkPCwkRO6ljFN84TDjtY784krfOMvAtg4YH9W1aVuqifWz4GnZxtOmu
T/ia/RX1jG4DYDUgOVtJZqGeCeJtvjMd/vxBK9HjHP7W//mOZzGYZVy+ADR2Kp0ANhlgNuAQ7Ey0
RCxkn4nIaZTzWLqQtcOUBz2eTsoFCT/ge4/POFwaSCyukc756ZPjvp9SUYr+k/MmxPZoIeh+fYuy
YpHxvtwAWleCI+2rQgid3cdp7hI36Ql/3Vy9xrkjcxDOxWvxkRf/UGV+0dJhpe2NLLm42ndt30vh
jCG8XG7YpbzLlajpvtOaxMeaFOvPdIpPokMwlq9lZk2l8TYSFPSZFxOcX/9ekr5n9VCyqyxRwxLc
AyMAmtL37KKVmiRljZteCPJRaIF5EiUR9wpDwT5slueLNWRNlUhtP6o6oMc+WcBQst3bs4LIkPRc
86hwPvC95jgDLMYODKh9Ub13b4xbm6bt+/sFX/4ejpffvRsz2vwWWQoUophALBU0l47lweiSjpAG
ZqgP+sATk51pJHp8jjwWgtEZaxf/KdCxXi6RBJQKyCTph2gZ3RozrqZRCW0xlwmXNgpQuOy09gM7
xUS23xCimzLgKsoMHGOijKtJqCgA6qFlno71HUWqm7DBxH3AzqKKVTyVQoRBvNZQhRx6eG8uQt8v
AWrHsEJYJGV4qWF85T+u3qp7iKqrnI3RjEvUW12iQUbAwC34DAarWKOOqSGiPTC8pYfXatQNCKav
AEPF3NPqDRjnN+G/kmOwlwx53mQjKanKAS0O6woBF246Y76fXhVxs0gJtEHqIPta6bqaCjBsDLqt
uUyXY2l95bYFiVynrtZL7nMPuzAaWVGnCbqw2vJqg98DNh+lKoxBGj5hW9QRKdt9yD+u7EG/ra2a
vo0YMk9xRfiZeZWrz47rteRgseLvQ0Fst7yP0SQEQMK5BTenKwPix76nKpC6g6Wv7GAIHQnIBrP4
i+PhvzrfiTGGmAzOH/Paewf2rvfRmXZzQkppEcTlZ8zbZPiJt0P4UhuZgb9nJtYEDL7x9yYqbV4M
MuhrYjQ6PfI6x3GXXhNOD0pUSGjHmlwzMbG0HgozWuattiOj7aFQUzvetYIe94sbOnMZQ4yFJclk
QBtthM4DEPLWZUi3+VVhv5WctaBrDPWMYnF5aJwbixr216pzZaHHH6VRt1D2+cWvn+ugHaKm/Zqq
BbFpvyt0LGZn+wF/8HQjn4ejKe0nDq+NTO4JESNHRXOwfAH4uZWQj4Ci3ZBEGGhXxCtfjCDqvayY
aRhZlR7/i9fXtnNrQFI+pq7elo0Bzxh80nv9fM3Cc/8Grtc9roYTFxCzTbCL4yFjF8OP5e+QmF1d
UzC9RZib3ruq0RPzYwhlpNVJOT8glee/hvM/bBE4hGqFonJn5SdFIXMLeqNmxIR3W2cx7wHHytfo
uRU+sf+I4cVnw+aqDJJ+RBaea/FaeoX/DFptx0EugQ8Hq5rmbcvKgSWsg6WoGyQjjD08gIRR7mkX
VFb+dytW1eCHhcax2biOnH/fZ9we6TJUwkiTiy5B1iFPC+93LuSLMywijFjy/4tH0Kf/ePOX5KZq
yRbszrlYma9h7FhPfrLZRSo6gK2Ac0u5+bHC8EkP0Jbo7TD6kj10aJgYg6bWTu0yQSIt7Q77+MEF
eVtqmzGV0PW6iczTckGpXpxP0ETBtzDYLXX23rjhF+d/+uxeukmFUN3Ii1f4DTlGhSBQE1AOCTq0
zxQwYl6c1W0Kg3k6SU+gF2dZLZaNNsEht7TgT9ztdSWfExW67oAPqcClsIxOE/KwwAPBxRrVtzfS
L+Q/k3ZjbhYjPzC1hGGuqCdLECeZzQmnouGEeawpA4wr40t972RnwhYV+S67EwBmO7zPQlFdZlgB
fn9WbV8zjeknmCb1lkMIuXFB+icZHYjKKT8vsNtv/f8zUS7NJZZ+N28PSjnadJU4BMj3/IPvUs46
oFP2tW0xjVmBeQwNtGQUQJh0sLuGgIxj0sCDBEeXm+gh+o98WGOQ0Q9xl6czPD1V5+AWLJdFE/wI
8sMGv78YwM1VdgMojYTrRPZCP+UuJe+aYSurSpdf3CEH7JszW8pLesREFz77NLxe+74+1va/Of7n
o+b+dq+oOMVoFPcWX2WuJw2QGKdTSGKbsXJI+LjVhXpUfLt5B9R3wyskuDhnwML8xq/L9IO+dFLU
R8LUtNtwGt141mWjXFgJTlzPNxs+STLP2ZoML0h/tozNuHDAHkyM0b2sM8Q2J2tkqMkfymVPqpLh
IAQzDv73CNMU6RLX+GOEt3ydRSCxTNVOJY43R8udfqxLzMLnEWzf8zEQ2P3JDq+iP5MLaVKT+i83
I2gnaDYRSjCKatPZoqc9JPb9bgV83iCq9HgZTOhe+hvQumnD1nJifVAJDj2gCM77g212glp3HALl
Y73k/1eRG1IB4vYU1IAlsG37LT9nV7t6aGmh14IxbLFsDktXJdW1LruFFioUp0yVBqX51utrMW87
CqhVTuGdWS1oqMIXLX3Efnvqrx1pG7VAflLoGSJB3pBT3cW3zgy5IadwhBh+T4x8RsIYJY6oNBhh
cnG8p58gL3sUqa1mmIoYdYdewC5CRCRrK/wYYRMnfcYLdJYxzT6Rv+aouz1L0IpWRknnejjfcOMP
Peebd9fWnfSRBtCSvvRX7Q6gq90X5MIZHEXb0T8pcMh5b3Pz5ZtVZRPjtjFASU6rgXlYzTKpPSN9
adqwWlpb8UcX5nD5NjR+95HXMyGggL4wHigLr3Z8hIzEmmvFRR7gwwzWyJO862TvSEewBE+SUIeX
mAWiyIzcvnb16UEvyEd6f1EYqeIo9b0r8BWLLRpYlSle8/6nt/oYQWUJCyLhVHNdM/qhpVzd8ag2
iARRXXbAWa7gp4uHXbOixeXFJCQuaZE6OBkTymVaRonjT+1ZseFll7Cfm7Rv5ryqjJFFV1NdMpho
dbfJ2UI0vTNb3qQYicD7si749mjC1pKlAu9fmsE8WMHZQBUOx6BbilF7XzxncCLxyJY+9LTa4+hA
E2vfWS2rupTMZeCfFmrA9Xmpw9s5DMGQILxdSPc096BGhm71E0ueaGubr36lB6MOeBDaNcgoHWxN
XjdP3Fl6MX5l5gI3csRttjyQ4TfRSkhEkfXfcsvJPLZU2EkeDSIdlFoam5rTHziIof00J2ajxK/A
6wSYe7Ip1v8XAXUbtfRC/3XZGzlmyDjM+z8QFhWxPnyXt5Wg24F7lVddMAcZNGzxWm63iX5kX9NC
FQETKyPV1uDfRLMdt2Vh8uo1gJxGSMJtl4p5dmfGm82LidUkyTKVMRznJK6p9wa7930Pl+Jxg6cO
wUobq8BRZQJ6w6bxAqqa4UKN9Kx3qmo7naRmQ5GbmmDPGKKXmcKGWBMe3fPnMlHCPdYcY8zKSKWC
IydtJaZdhUqxr2O71QAzkdc0hnzT1a/EVi+/uHq9WMQJO7dOPrFwORma8cRRCuPGOr2VceZwthxo
X4JjuYeoehAC0sGbIUKJZRg3zyuUYBUP0K5yYUuTQkIKJ0uD/Px60Wp6ZAqqy994o9eoXtfXPm6J
qjrlq9m+dCqnx1JqoXfib1UQHcZid2rKb80YX6NLjzuA9JBnqUZbsgI3Aef1O2RtEp13fGKSjLZg
GZVgvg0Q0oDS5ArlZUC0ZhP5yrSA0NzFNnY39gG1JNWEQku1owdLG6YgJn1jshejqiaB0yIHWldB
uFii8rWHa78jjQ820VaNIHVbqW0xsCwLtCY6qcuJWmyJ/yl3NPyjZEGLql6P+AKNWs3htzcvN7WD
mdQdyrNDdvYKb60QkttzBO6+deB7VOB5LSYxB0lFFcBokANhvcskWomjbmFyI3wqluqnn5umgw2q
wQtHvDoOa/FYg+a+wI9web/2uDKmC1UabC3e4Tj4DFoXtAeBNhFGC9Jl70m/r9hcrwvg4kmPc8sr
DRekpBgGewTkkgNMg9IOdUxsopwf9Ic1igXljkO9Vpdnte1JLDrQOKSa8sjYorXA2BCOP7urzycD
qWDwPCHO7OQQNAzZXtLUPtYGb027o8HJawnLia5IDqjH2jXzjXQKQamhC9PSiIH7TVB4s/yIet9L
a07LYDH+zHYN40uuEVngutP3kwZoNcIOHbBuzqrIC0Co7985yknDcyX3UnqszMmCDUPyCkeNAKI/
5Zug2fGXt6GUZBncEjbNdCnv1drzdJEQ8Ot0A4dnpyUWjXTLQFj3J4g/DLazpZL/7wqxjbxbct8U
4F2krxY5DJR4C5l/VPDCwHllt1gR6Gd10+ynRpORZga5fbU+9eclBzjalqfcULTx6T69pFM+D2yG
65DmFNRILox0iB0+nJ33Cbx4ULehLDE9s3w0cInp4vrLjW9Pqta3XRyWUiDPQHz5qbbdnyQF23pn
8cHOR8WLnd239BzDzs8MPFloK5V3xaHeWBDO+wxQtPxBpKPBdoc+PeqKsqiTEeRleB74eqcVjIG+
IkRQeZNLRm7b2Qo2pu2A0BEsSUFkD8E9NOnxFwIh8K2kbZGZCrs0eS25ue87nxZoEL01Gv1fB4LJ
IIgU5fc68MRHDFM6Je/B0HLdA7JfZbnGnzmHujOoL/tga+YCpqJsS6+vh8lP6nNRz0cs3e2ctyUx
mDSSUaMnRsVrTRJDr8TcI8v7JKHh7jbfJWHpH/B1RpqrV+e8Jm9xzv/P3/xNcTLcs6S0E8mJ+d4m
aBb8iJKOTTgXuDSbH3CnEu3XVzdaWyVyfC+ZHsiLdTQ+9e1p/5sXSnU5T7EMu0HOmfMoLkrsdwMs
+WQjPxvio5QxysPj/PJK0NPuKcEjw/q1xq/DrZs1OWvqJOQZbQxTNKbgXzFaqVXqXXQt57wvCVPb
8TaRV6U0VLRgHwPEf4Q06QGyF8iZEB5K5bmNR85UfmrnFNwtfULv0HpQpmHSFiia4gidRCm+X9HO
CEaQJCGShAiP6DNsNWWmxPIwft9VP4EXMwJ2nFgryFQAaKrI1bUfM0B8o4Qf8ESV6s92CMEZ3x7y
7M7MACOh4mAS6e7sb5JhlnalD0qAqq7nT4eF/z3cr1yaev/r9kGRHdD3acaQc2QyoR/crWDF37Gs
U9nef0LUAbxrRleCvXC/oRMwu3TEMBbxxjjEdOTDehzSaXmfP4ogL4OzG/8SsTWm+tlqfPqfRLMZ
AjqVItOxW6duw30PkqyAhjK4IRKVWlRmV6z5Iy8plQPDHtauXR4Saf0xnucbyWYMZbIlVMgiOIiJ
sYqtz+yAonLoTFVDmNx1zbZUpktHJSoJrc1v1Snqtwuhp9rOqhY40F6GqMqZV53K4FLg6a2PRH/q
veHaEHEMg4JZE07BrLZKxCbjSHeCs4SUsiZpvbGoS11QJQ+BvBQ1mLx30HeAPG2pQ5nfVUivkIC1
ypoxegnjUB4EqFCu+lVmsrB2p96F/RwF0C1d+hH+I4cnRKxNMmw0TiDw6azrKUuGgnK8mTUumHj9
aCQZ5kb0gUuErTn4pOT+9vKawn7JEWcJztSE8CNXj4DJSIb6PM5KI26aSPdiprfCv07q8ZLPxCNI
CBj//Pr65jAPgvHccKCHaZ5B/hrLMmnjFZp+zG95H3M9VPbCJwR+/YVSf+Nw2ymBSQZc+DGlWoX2
VhEERLnANYRPNqanKjHEvtvLi/Wq4uX8cjkmUSR8yCe4hb56WZ7bwUEi1RrmfqGjZrr3dVRNH2nP
0lsz8wBOREDD99U4AkMM0JMII0WbTZQjc5xwlb+UPSc+nqF2uQmzLdpvOh0pxj5S1rrrH0NjwIW9
H/lYbaUwzUQNfQWpIbui8fbJXXIMJkbpyfUicnD/V1ac1IOuDTO/XJACdwCKZHiVkKWsCcj62lV6
34rVJTLm6dtxeBoJRQD5V7LCTZEaiBwntt3nMjxOn9fNknbc2n+GosoU/oGdK0sAAvXKw6hbCngR
2Q/kgeaj8Sro1YvORrMiN5+qVArHrnq2N4DLxGe4f8IWePsgTwFoWoHMqJHf43iXb2iBQcNuHYYA
YxNPLHvJeIwEx/S7opm55EQ7dMI6HHdiQNusTmssIyWSXcowipSmSslfAju5KtAAz5Muir9v8dKV
XzKkFoketU/LFLx8cZFnzH6Je6OKE6mOdUASgIV3JIiEviR3AdyZd+LH0QOOoYjYgeymH3UIr7Ds
AuexoqsDFyCpUnUa8xUUQpIQqcp8wNBVLdCSTtwgrQULNgEcjrf+WOH4++bL2Zu9fkYF2b6wvN+8
qDssLo39Q7PfYKr4ttqVzUKmYelqOhGXbvo0UzEAmmpeEwpcNReITNuEY3L1Q7SmmePqJkt+1J8j
nQygm5mkRlgJQpvzlDmEGRGl3AcWpEK+rGJSXuoeGJbkvvs2jVXvak1Qcjyo1fz2yCT5IoVuEzdj
BkTANxDj76LusBTcENQrsYjQnsELTnUZFrMpVLVnPCWdqc8EAZlSECVu+TtA69UDn+yYS7N6mKfJ
8kYFYO7BQXSooiMTYpWOMh7YQwevkivECydDkvJn3T/GokEAUhuyaNI+RofKZ660rokUaPBnEhVX
OUmYvnuoN5m/OlXXxBD5v6YzFHzDtC3BXHDyS42d38mJ59YjKmBDz+nHVB/kSLz0PUYH+471jz9z
9Muh5MOPwyhgZzY/uOQAOcAayx/pxLkAHE6X0du7LBZfUvV2hoNYGfStEIhVA18nQ+Gnkki9iYfJ
HTriWKrrkBiPRluQAkKyDaJF6Hox6pctve00HuXimMgat78WdDClOj6+Eh76C+YrO9J/wRRdYCTt
YTaZOQnmM1C1NyhLSy2yBTu+wrhcW0ASQcSUHQoi6aRxIQcjoQmDtsqWMvxTbUIt05FEOw9n56Hs
88e3dcCzA2vAWsPIfMx3pbAoK+IeVgPB6JIAsT8XJeFDl5+2N/TPAdRpiAC2OREYOTiaBg3fH0ye
dMUAqhKrFQKg4PcQ7xlXl5abcxsJSRaaT+Rf5w4xR4sQg4Df49pMAh3mP5o/h19IezWgpfyWSzvi
1kgc9tZbNdQ1HbUUXDnpvb/KNPP0Cid0sBpIa8wm/tfxcOGWfLWH3GvOIMekO+pVpLtxDxuiP148
Z/E9BqvtPCBZOFszzz13lLWuC3a4Og+ylBN6IuzlNvjxzG5uw9jqvfnY9pPVm6X8P+wpxfwOCzwd
v1KZvSwfRu0vGHWS+Bx7JYLbXS0Ua3iSR59TgZAKZtHqjJbux+Um0v5XbMYsADfn7QaLdMbtth5O
vtNGTf5LJdxAQZhZGxUDFKqxn+xI0VgOnYOyLfJf3JkygSq+lkgcLa09ldjEdLXLpGttFzqZSVTK
qbM7kDjR2V1dB4zmaGzZgGZkpXWuL0WfTefS9iPljta1/5V104sd5T468DzYpRZTaCOOWqXT7Mme
L8SJNV71rrFbmBIv28FuIlpy5hmr91QiZFJw/tStGT47RuNQT9v+p625VZ/an5q3I/QZJDwIceks
PRAuqhFjd56SGdVC++kEt8vphczfkGQtIwOzYA9oPS8GjOsbzAXg6yVRg9XNMwnmO71TG7RLhVkY
pjdBN2xXzRWDWlJ94yi0hmCXz+2r3WWn6EzjJiy17vWcOWBBJpIAnnSW8etpzsgo32A7G2ttmjx+
RVadL4H1pTSVwaEtikA4ONxvhEyfzv+hNr9XzVDXGTokuIKclBiTd4kDxP86NbjIuD9KQJPSeSir
SypTRQ6QB/e/zmAUepauAphH6xCDMntQhpC+tBimXB9VL4HzdjGQxofbn4KrXrkXez0WWx7Kj0Vo
a2ov9ZO2mRK+TDHH551IJQaXy8w+Nmfa6xC48bQ7L5sMpNW5qUb8fqZUxzyQHpmmJq2kJI8w8wdI
F44eEWEiYGIy0FXnfxKx3w4XiZ2KR6loa4LcGT/6d9enj1RhroX6GbJQ2OR9tlWb1ClD9mEBlOBe
kPDrG1e+CEUfl30md8pI94iXzi6D94NSq9fNcYyqyb70fLHiJgfM2COJdjv00mwHFIN7XpH7s16T
vjegwMGBaZxP5kEzjRBDUOaMqv1N6qC1zTOIN7sfd1HgaMpRUKJYhUQGlL0s4qrfwGUkvHekjlrd
+gGJCn9NnX+nLYJQqx+cWi7Jz2ouP6TuxWsU533vOMJDtuUGMzmDMDeCVdefoRuoYii9slNqs2P8
a+m9AeF1sStSO7g/Jha1sFp1ynXzzvmntrnrV/zBecAtld15QY6xCmLBnRzmGaoVh8MAIYBDXQq4
xsaUyweILwoRCr558YlfQTFB+rPytbdS3A7z7Ka2p1MHHNOlGBsRBsSe7V4sKsdyyMxTk1OXcFrn
AS9b2ytVpLeNw7swSLDXOJ/SuwQuUElVDmycLaxirAvcu0tXSQ1T+k+DHnntlRQb+wilj8/7PrY1
O+RFQIbIsrRM71sj051wha+3ikXTr7A2rCAjvIr9eCgRTtOjIyuzOoj+hJW8l6F0vOaABhhzktur
tvdm3Fmr8tHOiSYvaY22/Oy9qTlao+S4BeVoO5jm1y0t9eCa19JnJT68zhqhcjz8sDuiu2FhG78g
OVTDXDdct3KDsre8iNKve/+TIeIGdNgQjDvA20ux6NYtvPvYaAW3+b18/6ZQQrfBX0WGxZsRFV9a
UXUwcmAu5SQwSHQo91u+MSUYX2YLds/E5PpdKMIg5Zr7hg8IPJX0LmUpJU4r20PAOKretS7t2Cv5
d/P/P5oosTYJYJBlP+Vu/mBf7oQeUHrv6HQcVg/tuTnPkPHT72pUuK98fV9Fc8zRC4AfsYd7SCZG
/rocQ3z9XONZHmBp7bhoWZF1hEGrxtvuc1T0GlyhZuKwp6mOMu0pEtVX4/Z9QiKvQGG33h1OKj8U
V/gNHVqIsWFhG+gYVkC9Z5t7IY/6wirL1+AMpBectx7F0l5T9ktYHlxfSb97Zg+2PTpStX02LTiF
kN/gVSMYDC6mooaiZ8WlivOAw6Qa4kELomP4dR6HW+qYam6/jlRWgkZPOckdg4Zfn01K1qkl6GWJ
W9DdSJKGsn4wZG31vC+VbqP5LS8Lm/6HrFs7hsqDuC9Hj8QlDlMCl6NJc6oFDdqdvld0j5Paql79
giJ0bplyiLVE00mXc0j9BMza6dQBbWNrxKbdperYGP9C1Jr5NtwxIREheSQZPURcIs0SVkl3fhJ3
Y2OffX2fvtUTOsvSXp6TrVzXL6FBbRSABnA4ZDnXrjzWae21mVCxWF/CLXszQ+CQl/baOSsacM0Z
wKdcCcow5BTqIxBOIV1Qa+aHSjnhpeD/OED8Wgv3q6Tz+dwAwp2KFEwObaG8+/sx6Rm0slC/nffh
8yfsUwvQ1bDBD1jZo1FftB9VmltvS+8Qn7T2jlZiSKviYeUYH3tO757jNfAywh2S6Ro1tUXOlgiT
ZHwcGtzlvUBm1OPGxQqMOrpDdTGulZ/Wdlg1QrachYKNWhoXIviuTLoVeQnHKXJf5zxUjNE2/9CB
B8rFDJSVdIfUWdbXfVi1OZpLTIuv1uK421wc/Ujnd0DU4HmG2xZadmGrrbHr3AEdA9EmYV2Foeoq
S8bNGvJnuVLX4h61YqgvJCHjDsNyJAoYVVp8GnO/8sti473taUraQ8al0ErcYIPjy/YMYmWoDvQv
II7BYMIXwb45P2QdUAxyU15kGT/cAO2aBRGIlts+4HdnaQCzM7DIV+3PLRNftLIRTqfbq+LsWUyt
NqGRSoyqgbAMi/SvwekJ8/molcqVH+5h8AMZDY9kyHZi/3CHQKdIBGTyu9oBUYcSHx4aMeM1191u
2Ah+34XnyS7clVMaETBEiDxT0otbvBzW2YhVxPiph0p5/8FlRKmP/jZWl7Ge2NuiUeaaDg7S4hyD
1YRxtMsEYTG4/0tQfSUFuZUiAcc6QsCdAhxu9lfoOVpDOq3E/ytInSfgQPxEVzECkjswyPF/F/Sm
smlp6AwsLq5yUyx7HdFATZiiRX7s7oo+H+Jmf0YFhjympFAGTnaWIzXjDd3zO2XsPg9nicneG8Lv
JiJDSNYokqzqJfwm+rQx3ECcaaONUyj/5HUcc+8dYYAuZRKnjgglhtQU0NrWhBegrUeYRnhp0gYg
+b5ugp5Rt8kkSML9jRwonUm7nc0Gh09K6g71h+m4kandxZTat3JJpVlVbWhSefpsYZGxA0nd4HPc
jeVJsJUxZmSEngkt7i9TDKEyXLk+oyUyi8ZkbAiiK2fivq38QPB+zmrrDaH26A2WOwhCPOrzl7kh
ZY7EYABr0mjPsCXsgjy3aCXbZ3Nr90G1LD/U7lU387QSXbYG9TzQqZrdNqXbVPtUlpWuXYylWLj1
9jpu2anMYqHXPHhNp1JljQYMYyoef2dqQJcbmRh7i8Iuc7MNV5g9Rfs/7OlFkKnZkBteJ0F+fkP4
Cp66f9Lw8ovwEQyM8LQFLJMTKJR+97uNiak1nsyo50FvkkE6cdculyKB4FyN03FaWVnHgbrApOYg
gyUf8n+vw4R3AnQ9Q1vNtdRDsgaSKX1C1d3zis5BpSBJUT5tkorsiLwjSFcMyudBSglMFNfCd9KX
M5FogjjmZ1CohOgkf0n1xEwHHTi3UafzSVZpUm8Gjx2Zvq9Nj8ySmb94b6Glw5/fbbgPqBlLtl0p
SHm2drqvDAeB9KDQ52fLTwRG+TSywDkJBrFa6Bv9T25mVZQq7nKyAyw2kefemhV5/Ue2OQh5kxUt
CyrcOokC51rOTDbD3x4gskV3ufgd3iULW+AcQ3oFOxPl3XEuTquAaeDjgAV0B+pX+fuqvP9++K3o
gJKnbZgXWw0tBMCeOFSKmWjoacZtxb2/sqHJlZAXtTejO6ClW+6stBtRyN069a6nZYDw1PPii83C
AVbXQaiuobzJChWsUGcYhjIBjBj/7wKG0dGsaBavsT4sEUL+XjZ41eqrSrDdRCx2LEE05xKKOUuv
1C9faAHB5RNKoepdY0JMHg+iP0UQYZ3uap/Qw7Qt/mp9+tlD/TvUEcRSLg70SlSS945wIoet7KjW
t4z7mZIZgAYPaCR4BmfFwx1xaCP/txVLFCDsuUOtf2dSkYFv9TORHXIPLYpF458uLXPOG0AHBeKd
6BVFYENZEbaRnajkSeHgMcDbdE7vXemiAKJMzrvBRvpdhCp3RAdqGEpZKas+92DbbM7GWTltdqI7
8oWPIk6WzfhNifaYvXOQdnJNBVKkTisHWpMRRLPQM9aFkTsArTvEyvYjzbv7BdwEIdn2CXA4f10Q
zEa0QKZJRE8D93qx6JI9Oyo174m+jmFDHoBd+YKyJ2FqvEZA9UDeoqNdFixRJFx4v7W+CC9PNDwh
p3TMG0xYcRVaSXyjQVR7LlSiG5HXaI6Hsss2+kIgpAFHNJxZY85jbdyGP7cOmOT/AwdUktH3/79v
4Qc4l4W2wTMBJiqYRlF4GMiyzDMLCCjQzmD+/fD6+kQG5kmVc5oIkuOerYG3/UgQowgmsWY1CnU6
yaWvIS8atPQUNgMxjGCnXT7MPyqMdDc6ehWrIwll864IGSIZJaMGB09OF+cm6H8mZ05YBPOA0tfa
NZ/cZrVc9LjLbHgnuAgG+o0WBhPsrR4+052cSF/2gJAGE53XxebYmKR2tf94zoM2VXBnQEUjGm39
GCNtmgJAlSyzOQqDUBz0AhM4cLn3IVqQpYKI6Rcb91KzORiEXaHS8Kg+WVECw9dT9+rAG2zeO/YZ
M01d0+kYEn3nMmU2fPoLgV75kcRBDQlgpZAgP+AGIhihnflCcbIhFGCc5brvnAFwEz4R1k7YHQVv
wP+goawvCcYaJ0FnVI4bXh3M5BUEZ677IMWbfMRVj7/RfA/b+gpN+uRghHDiYVRZ3MPABkm7u1kX
OC6adLf3sPWY/6MihvEj1aFesF8ynmwT1Y9HQZyePigwUPI/C/GuY380uaFYBNh5NhCvvpqs/TSf
q33TWKe2m03MHIcyjiGeeFPoPLoMRP3P+rNeILmxykxLfIYhSJi05svv1C1FNRB6jLsjm0V73r9l
B4bcQsE8myZ2fK/SNmSgun5oahTZ/FA5YB+3PpYu8/kVE4lhG0+h2EvPjbApGhnJgIS0wepy+2sX
J0zviACk0gME1q4fI2G571ak3SJha+o6xOL2fvlKMb/XR8pyFfD7FKV+4PGvkYCBGzAiqH/9AGZN
5KluEjDgEBUWb3sk7QFFqUL1TuArFG45hHtmLuBK9PRShsrf1+TJu59WeBHprHO6Rxkcm1UiXv25
RwrOmWDeRvjS1RYZWcRiVMXUfyu+qCiizgv0NaGNT7Tq4aU+N5VM4zlJt82Zop4sLcvYmTSrcqUa
HTUpsi4ZvwFy15sv7yEwgQJSaup04RNYyC/msrxzG/AmvZPUxnhIgvbVSmqOJLm1a07HeIFdgAGi
adwPEimxuqNj9AX+5JNeDBBPsoDBxLOo7eiJxRocvvw0dRklNpqIG21bGCYa71EWF3P342zDSGnp
/TjaYpTa7mT4FtNdJyaVgEV3JUyfSEw7vxssgCwjJ6HbGthRvvn0R26l5bhSpDxIErdNrvnWoyjG
7ZaXDw18D6SVXAmvvURuzrgnCJLFbLuqH4lZmu7GngnRcjMGFtrx4YuBGsgjslCfEMQWoj/nqJF1
i5NAb4YQYnIWUUM7V5cDZP+6Dl/5RMJscDxpclx1uW1vou8YdeAGOog5KHvxnrnGRhNZspoozBRn
/ZsvfEhRwqgvGmMQf07CVmanfQiJaDW5jyMx8QsblEcInrLNYcuv0/Y1q0fJ59gYg1yLRgR6NfH8
qKukV6vXvyITPMuB4R+LaoZ3AOAMwc6H66nfIrQNhGVCchybfIrGAP4fU9ZMGiDLOiAdbNOXLC+r
O1rONWkLF1BtWFtBqsmQlxJyQZ4S3Y2qBPBJMIjWHgK18yuJHT6JaaqJX2l4t2TbVodGBM7n9rM6
JHfmROtVhkHpQGM8/GY+p1R1v8wod0I7RV/9+9dP0n+QwghU/D01JcrWbM4COX9bIzxqC0aIe0mg
NbywHmC1D9ASWNpLv9W2T979zCmgOOm9727VJVX/71iO9Vqm4OiFXNp7s7hU1zHKA5exxs3WN9or
fUsdZvy+WtjM/IBNjohJwm0x9Uyib5SeF/SFGvVemD8fVmlTnE9i/xvyshTT0UvZL6X/bsc3aeSv
QXS7BJQV98Qyvm+gEjeOWpSmTz3h99ZB6q19JWuLu28jbM5DSSU1niKVf2NCErKXy6WddWkFjica
6OyU6NI0JAaD8g+K1qQQZ7o+vpDAhPNvZsf0YUHBrM9YzGlAI+1tDPDZKTqTvYvCaSqhiwDhlDxl
/JHsgiUpdOjBPsbDMKgoTCKh/KVnfXAZo1Y/hDtlMhx/nqOEhamts1kOmDxD7UDq8vLK0GhPPtBP
MVAfjnSCDF4q9mCOdkxCP//RiZssYmHJ0/WGjaxjvOUUaD9hHxRRgqfVMpkruC7hx2E2HqVnSL3x
AxqbV/WUmZm7SInhyULZR7CVm0P4UJYq3kEeDE0iYtTcjOzl/3UHwz2TzvIyGMqMtfOldBgPCwSw
2DVq9hd+i0Z84EX5m1D7EZvkutQyB0FTsFD2ChkSm3BoBIOvwViNxemLwh1PMwyckSVo1uONXIxO
w3/UVMdNg9bFmKdOi1cCwW0Bbbaa67Nqigqm5XaLPCvhw91qnT7WyoXQinfndfy6r4uSnKQ7dS2o
vDZeSKR/ToTVL7a9P3GNvni+oYt9/xZybJzJX/5Ee45eaYzDAYtmWMOkjyr4z+tfgqCbpm4iMCom
eRkW2bl/aUj7uWQOE2C/cTRHS4OtyBevuvH8O/GMZPPbzxurXBrLYd8FJXO++uMrxBUL1nsQoQYm
dF5FfF5Hm4vdHwFYyWPSmWEu3jpfC0qUGKo94UsajHIn3V5uxSNvKPR0XGe3beGGXYKDn0HbnZbH
VAqt5cuxa9lMJ7Bbo/Ql7/pTC5qv0oazuz6jTgMnQuT1Vpm22Pe1z74+LzO9GfLFWcNbWhhbT6+7
TF+dl26yJLfDGw/rl2MHyHcBjEkUAd0GCgQFTVmpG4Yk9vmX1DKJRw6zM95H4E3zJtg4FKAA90TP
gsGCnulq8qnxY+MdOZmsnr0eJAS3zUp2+DOXjD5LP+ejkgo+awwmpFlqVSBcb4w/f7Yejk3/9ubJ
TwLwxcKHPLOEHXafw1I/1Xs8CSkSbr8cWQM6+Lj/x0UGIiZaX7IMdq7GYoeIas86ViqI+lTIcWhc
P6o3m3nF0n3cGw75G+O5PRkaTwVIFnYwHh+xkh7zXL3LIS94rvxpJVZYBZZG1W5eSzqFROAsOIbE
E7YMWZJhnD3ja0wh1wko7Zy0ripIgJxpzYGfsPGx3gYHRYj4XKaVQV5kMqlaTjFWLDneefWXwpZg
XtTEXmS5IW061bz33NlHdD7GXN50/qsSQzIJwlmxv2JQl2NnFCWsU6tLHZ//bXJ1fK/+tpDmek4/
16FJsJWJnHsuzkSGWYj3GNpex/693g0liN9vMYKkdxxllAVmky7dDXIiyHjgqqtajUrUZdaEf6Es
kHZqIrDVcaXQaCYPfBWGhheMEja8vrmbq2DtmEk27l5deAVbxY4232HXTVmQF5mvTAockCQVs/FV
SYyusX17I9B5YT57jvshN/Ox609EkEfcJiPTZE53KkbugcJRPd3Q9KAXt5zk0QFToR6YwZ8evhJp
dt890Iw3NUyUt0cWmZwS8BI+0gKQxCAyX3todtTscGvz6w4maM1QtWVQAutYBOzteIXYL/s6Hpez
vSKzh2OYmoe6n7dvFErExo2J71+wHBtkYJppibj4BZxqUvD/pyBx0EBb64S2UK+AxsTKsqbReej3
q2+z8TjWBOtBwV/HhKKNi+E7WJJH9ZBcr77cy8nKXacZ52eWSFhGuRnXsZ+dOIabpF7+66dHVOLZ
y5Q6XdTnBT6Z3UpeasKdOraY+lMk5LG0MtnDJoCzfBtBXnMy4RPdbpuyjTI8IFV5bIPgJhVla7pG
hKmXK6P/yJeadGqvX6oyKBN0m9LL6eBM+4bfLjl1FF/N56Q3cyctCbn9AA3mL7v+zRATAwAXRgVn
+lXOOo9R4OCLsP7pGWqi0uNoZcr7qtflYUyhTd2fCbxPoPrCpoAKM3wZ0ZIW5O2KsCte4eVkXZnX
1Emn/Tl9HjL+9mL1HMcLISZXtLPDQ9dy/Z6XVKxyWBDCJxkgEdpG2UW4K4CJOZc2GpkvjGMBHGOd
0dg4P93BID+PMEdr4fs9P1h5Gyrs8sFHpWvsHkTiU09F9u2Hx1t0cpIxjlLk/B/4tIdm7T8+IBS7
gB1ylVpXIXWsahuKdS0oWUyGr0cnXT7+OxP+DYqshx1j3H0vv1mrIKl2NxhycIRjvb6FJ6T1+5+j
qqPiTv7Ki33ptzHyoiyNcemhHkKbL8Q+5/27Zn86t3TLbjYScV+GSgPj1bwrzDPLoWNDRadAcQeO
qM3H6Kh7Q1BsHPW0LctNmhSXh9E7AOCmbNHYtqkzjyOvP7bqMYCYqnLL8FDd+G4kO0h0bV5+i9MQ
+gQ0ktKJI/pi2X75lYh4CPcHyxQW4IO+GY06ScBhRRHle7oy9wlbyWg4IAbeCaG+DeWoT/iqCdvz
JPR2s6zuwLenHLcDHRnlpZmr5xW2YiWVa57Yb133EBfuL1ggpSbnvDvRL03EHX9Tx3IxEwb60miG
6qMXBeS+J9n4k2pBjhZjvK0On+OgK2KC4wqXHt/YT68jsGxyXgN4063Q8VFe20tuSqKhJiufZku2
XvOTTK2pBECyG+GlbyUkae8G8SPdoQQ9slNqilu6SNYRSKfWE2HPzImm5xm8FI8PS8CCtVKh4JQw
l4nT84b64nQdJxLgyIBcbP2kvDr2W8ojNS8aBtPT9WldThOYHhWaEhNahxsRnaelGy4k9BWZnAhE
7mR30kZvkHWkC0aITsi1taK8bccyPpN1Hhe5s/+/MQ1fuMxr9m/Uv/72MipUKgE2jd3nT24PuEuf
aibUSUN0g1lNGiNpmKYxLtnsOCS2RUgLhRzEHqdcdlFm7w/5vU6gRXSM1ss/cVntN0lfgyBHpTer
1GtxvA2f2X5Hnf0ryR4g98ZmdGcODt/d+CvreCL1COsKL6BoTMvoYe3H84VmiQ/DXW98DhyE+YrW
beTb/WT17po9DyZpwe7eLtng6X6GWFX9qUPGgKk8g+uKw1s0wiqn7+QnZbwhbQajLoiDsgUSX2R7
DUzbMkXirl3J9DrQqPWlwQyehxFZyFccc8Ixad4o6E+wOX3PqpyTLrmyQL069lVvwB4PJO5+k5Zn
Kldhr4lY6j/OdKYaklCiKxdgRMRULK37WY+hWWSwHBh9iwuOQP88RPwX+1AMARtry0hTrKgFwjk6
s4nqlcqlUjiEnCaCOkvygl4lJxTP2zLVRJ7JR8lyZXdciMf3wqa5bVTQw8m0ZuQSfG4y6GXyvTyK
DU4UJ849nviyMItxQL6TG8Lnk9w+sIilc7VBCKUrwcXS26OSmo+9gk0fRH7kXOnMcPBHnKkWflZs
R3F8lR7wepgydVamVQb3Zx+JbbIAHShcwwGNB6lZc6D/VmkR7BLkj4J5FYmqozTXn13d0SCDVGz9
f7FCvMgwvAmb766LFGyWrMhASjjDDQPJ4TQRnimdeyGFx8KFKAx/FMkCfG6tmMqHKeQufYv0jGiy
E0tlIs5bPIi1O14o8LYQFRWzQTyVTLuKntLyh9RlHi3JZRBV2hnDfH7esrOI7zghPCiHmWzk6QJX
ki7LaRBfZDrjTU86R/xQTqNV3NchWvixhApPtzho/5miyf9SEAMDfNZ9TMzagDZ73Dv0+pjQ8ihE
2Zo0p4Op3LQ/6tBe5Ygs2Req0R4dJ8FExEDTGat7JTlCs11B/9prNnofLr58WbsVsIO/y/GdrGcU
x1G7BvB+eQVC/dYAS6OaclsxXet1DKJbnEPOfnwuPYYvevGGcZEQkZ9yznNAi3HSOn0DJTq4UHh0
VdJCq5pvi5Fsc2ucrTWramekcab4Sh1YSEsE/sDFKqSEdot5hvtz069t82SiM/kqvHkLSJLDCbQE
K1ehqs0bQ3Qo1NwCjxf+UWxxqCfcxL+aX7mcoxbO5tWw/tAFhrFXTTzsWpWiyoFYYatJwpRnvECw
8gizSsAbHxQHjE884bGqxZUC7Exm07awdS3TAoCn1nzgUHIJAjIW0jIhzJaxPQ/YInCG6BCZ7cxp
crKtCho6JM+W7c14qMdQE1NlhxtdEXAHXCAytpQD+pVuYU0nGkZorNYH6xitWbeyyuPhDDg4TElJ
ZEOw0Hrcv0apUIjVT1z6rrFBVUmUWLBv6PYdcLispUuwi0AAPqlnZeN5oHL81bYJTwiLJwTDGwFh
+zavx2KW4Wo8d4b0bEvn1ElpQurqcryxXhNeQ0LERMfLLdMmaBZtCJBzjtMzP7cnsQHDpDfrJsx2
CX4xXRF1zaErDn8f0bXd9uye9wzzbOgwHoDayNZAeY010h8MiGy/j/L+rvOPKHWFvJFtNaZ/QYIF
uPZsUIYoALyudxir8mZfsW/Bl2vwY4I7pPMWhmhzAInC70p5X83mT7DoYBsvXEzkHC+kphDQbYfi
i66lajK9dOtgupwKK7xO6zjEwk4SRoMONr1nI1ESrmmTnNj7TFt0cpMZ68F3ALvr/LsI9Q0TnuN+
KlZc606N3/E4enEfqfm4Dl3DqWydNMoSYqvV7YC8b/JVhedmquRHDasgPfc0IyZEkfztk1j07jzs
ULYfBzi2bt2fV4h6JZyuuOUmyKJbWfXAHR/9xRi5an7JNdWVqEg1kaBzQgElxIEExqfT+Z2fJWxL
4g7NYBDDT44Emu5i92V6cmygiHhJGwS8rXFrfPwiO6jqnPhFt8CfiOdcJfE/thG5iXlQJSos76Uc
iPoUiT/oklC8WvG+QzoTncLRCyzhTgqTV0hk0/hKr3d1Mrj3zk4SdkYy2xAhpUewUVsscN0IP2fk
5dNiaMorOizUdSC5w2RkpnMQbEbHpPq8swtBAR0U5Cd3rj+sVJfoBuS+491+9ARmX1lo77UqpwZu
KXKQL1QOtU2cKUY1XCYhVrp7Bk/LRIyVk87Qh0EXA+BE/pgxb3Xm5q5+P8R0IfjG5YZZuKFVrBwd
ekg1p2LYip8mwGginZtSGc4hcfrmBG4QgR39LGRUfFYW3dfHLZ6jcxpD0QMux3DVsxLWSiL94R1Z
P04lfHUNZ6b2LN3v1US/pUEJXEKr8CX9ak4hI2mOdiFwXjNZ6BpXAVcpJ4oY4jQJ5xohN8CGQojr
JqZLTjQ+yL/2iXwHGLrzuvTc44tSDydwwmyncOmPUihYyD8dkcx93V0yYc5+4ejooqtfozMOhueh
xg9oMXA5G9w9ODUOHmR8Y+Vw+7e/HN+RWSET9a09BjBkY9z1CbffEUDsWpQNcB54pM51s1Ry67j6
22+J0faIOuS/29vmnNNYOBS21/IX5n2LTvFZiIHUtYHJkIPAwJ6SbR1cnHrdLGpsHK/JjOa3cQqd
1Rwmqo4rgZ9Zy2MJts+TF3AL+Krbgktyy0nsPkKiLgynu1ROogXCWbG6N2hDe9jom72F8TIzHi8p
onb2q9eipx78sTvlqYMzQQfzA12jkquPBjqVM21YsmtND/Crbx0p0DipC8LvUpar9HfM/8zYLlW3
UqVKWXsoTxFwb57nSNnzsoOxr6p8KUvbJfcD54SfB06x6rkdxfNNiYCcTaPNkPTlM/PVJSlqTVUt
77zsUFFW9fWHBxF+O4pPUOZ2SNTEStQwX0JPOaRq+7SUcgDpPHyUzS5YexQquWcNivn1UP7IwJU3
rLqJjWAkrSiVPTNpwv3TTtqQIVFifRbuW66iSEY6YJ++o2vaFsXDqHgTz1u6+LnjH6sK/63+5mYs
eLUmXYVnM/HcyxJXyI2rYqDTLeN5gbsOPIU3tMtoApo12GiJZ3wKdl2WeHCuao9xgBkvHXu9ohwj
fD51E2RuCYGcsypYNOtEawA/I2/60JBGXbQnNuiOTRJgaXXh93iY7Y0a+IeCgudey29vSztDY2qa
SRzZxlHZmfSjP2AodpJI1ED93d5/a6LtbYuRbZlTJysIY6UCsjQW41x1P2aD4PXVqUndgpKePSdl
cSvtkQuhesbkzEej/TqaiKcgRMQf73hQX+RdQCb/ClaCCRsTveIOC+CTuEdLL9O73D+zDnm44V5E
/5dejLYrZ75sWVhJ4HP4dU0h6HtthSome7jXY6ILTmPZNvKvvQNHlJwhrj7MDrrTodzr8UJuq2fx
TxYsgYHRiH+ZCGs0dusH4PVEs35B6aydVe/0VIzqHe9LDiJDaQR+xnU+t+9AVWPLWdmOWDwJj0WB
xT1EAeBXHOG6PBJL+NFM6iqORGEONaBAKHwexhE0+3akREqYR/bQuz3rMOBf7pLvmz9oYgcA5+Ud
f2T/8CUjDhev+uOdkqiADyAXzQ3RMXEKzGi6xjmboU9mDbG4v/DJVxiBHd58M3vvuCWdvNt3/l8r
nRBEuAt37WKti1SWQ8SJFg85rCnxPaItCNJz5j4J+plxQiUf0mes93mEJ4WCGVLDbY1uSHEb+pKH
KQZKIKEFUj/5KTBaM+nPBl8EUQ+EwvevRV9xX4w1S6XKBdVrEsEmdHrRI17tyDxD4FckbPzqxinD
Y9Sw7QyXwCr1F77EqC/WibA2AOIwE0/DdOGezns7rr8X7+vZSuiwvipBvSZ5df1tPuXq9bajtXiK
+4MkguSscoBPgaur0beU/Dskw33AU1rz8ZMUBHQBmQp2hwFZvjb5ybqkid/PNwfXAYfr6YYD8Xj2
8sCl6DhmRjlb/GZT5ymfgqsdACxEHWVaeakpwvQU3XMxbVcg6YikjwP2s34Q/39udp+TmXIDCRNJ
22D/ZB+IRciYtJnAV5Bt6Zlxm4P7nzrO54wrKMZPzNa7Zgg5VCM92f03hMYpsozpZKlILHVOyywH
40Prsi7zZTdvtZqr7/35WCUpY5tr70HItu/2n1Mr7icIwPHPcvagi58RwfIjZ50UNBHGXOAICj5E
9dXzEuvSB03Vs8DLZwi4Xr9onVRZF+dbXZ6ki6JS7sGtaStcofmUuBepTlh0S/PA8MI8sSTwzHdU
O2JLx5Uctmgt1xcLIKbKYUAGQJHLFBmOXesb04NYYEt/MNc9/AkESt++TRBrSvkF2eUHJsz2ji3C
02F+sBlzPhOKOhnkdn09loZojE1Ak389XJN1Dp061Pp92HAgtJG+/ypZ5opproe48tfUd2h2dbeI
sxvkh3QX0WoIiVXXXVPjzIjOY6nIi29YemQOTwLFSJAo1/PC49lJ+7Q90cPihGuPKJEv2E0ALJm6
BEPMSIlcoI4dGKUdA5QqODo+HxXLU7HnaPEM941M+7/kwh/pQxxWO1cRuZa0sycH9pV5Go49AR7L
a0c7o08KqyBC46RYSDQUKnqcmG/RiGMLYvtczUCtQXwa31y/JwSg6UybSlM4My6bmaslSSfcUnds
2v+ZO1T8LsHzvL4c6qNHjiFIepZ5bqSioE8LFuOZDLBddQhdGy78KjvSbKmiFOoCtwkI5Lw+ocLP
NIPc21WCuF/a18DizR8mBFknvUXNhf6zPv33Fvq2FH2BSWys6JuS75b03neIRCtOzMLnD97tRiCl
+oI7557MS2BnfkkgbwsnePuJyEFZkn+xpsto3xalo22hXSnZ/u/l0z0ZfWxkKDrxivtyK4uwSVua
rGTLusYL/y8oc3lQHU0lScXvRZAh75xrN4Mm6u4DJ1vOwmkWzhp3oL5eUh6Zuyb3/aw5tFXG5c/c
GgtWOT2cLJQthxnZGHF/yoMIocmrzEK14GQZPG39aj9a4AHgAnizep+f55Q4hwF1DawjTIHCQ1AW
Ejwx5g3ZtvSqTV+BB/pwLtO0mI1B6xMJeJOGV1QzD8xIlMqn9FU962cdu95uNlsP9CgfxP9qTijr
XS07PlZjHtJptjmXwNQonnzchqUSkpF2ys/pxRMfNvv57/tIWwWxUsIlu6ZNv+51veS9wDyJe0dz
AlUm7+NBWjnlT4gl5CZyRul1AOY/91Q5qnle5XslItSi/n/Ce1lBddb/QIWKDy4dwl2CPYj+XN5a
w6EhXXoGnY3xJ+VT+32TLOoPZg7GNQXp8IVxXRPp5V5QtX7RxG+PPrJjcdo/eguZqPVSJVQlfpMl
s3VEALplAOxjXUNEG4EScfbjFdQ+f5kqjYpROvokccxVc8LYsNYPT7CDkIc/7CR0MWgrUijHDzHi
+0BEby0A4z26XJ0Hj5EW87xdhVP2pImjHZyrPjTh44draZ5UnGJtAm0I3wifNrQxd8S8SlV4lN8R
qpK9XSIbaoMqRpEEID9mWoBf+MkASE0u3GI+FppsJuHoRGWT4hP0nSgqvsXL18WEf1ARDpurlQPO
cqdE6mClAphXu0PkGYJ7QbVtq/0dtZUPhCFkoPOnjTSPunQ4qkN5Fxc5sdPxSjgG4UvCfy8KQrRV
giD5lAk1c6krx/3lHfR0l8v9+gpgOf4v89PjYnRAtcf78fW51hbKVoWY+wmRhRaZ05OSAmK5NmnU
XyA9FTY4idNZIvSh9EpArmy0ecwgzvBFrOJBEFU6R3MwssMyNUgys7y8wDAsipDPPTv/DMHGsZNZ
U0Gy4E7bnhvbU1sqyiQstK7f4GRVlobxn/0exHnl7MeuhnLPvKQX/pQcpsnFecr3QhkoVRRPX1p4
uTqYVTIof3jYKuBs5BLO3Nwy5g0EoRchlPeNLYPka36CBttUb7cTQ/cq1Ruo5f/TL4W/DVU1TjIi
NT/PHAD0oixs1empXE/kDPcoryggV8qWaOFHrajLAuf3k0cbTbWqUNpf+A67sGX9Qtbs8aXPZ2aU
oPY8mBA97BiO50DdVtVaKIrZS8QaRjPT76LcYNBg+XV8Gd6VKA+dzUjXqZEzPDCu86zRYE43Pxkm
O7ujCmhVOQp3RJM5keRX1TSUqFrriph6Qdj+HrkexCThkJLauzf7l5RpnkKGsd6HN23ynpmuaRC+
ocCyldGIHOsFwpjk/dkw4nZUIxfkJqvHp2RM9MRY9YKTbU8OKpQhzKtlAI/B7ExQMy8up9l/ZC0M
KiwttcVwZIbV++o4UMWoX5ccM+tnGVM5OsGYx9WjGOo4izgPDb3/fTSqp4G6NgJBxPTXGoLwrXP7
a8dBWoGDLdqZTf1tREV5LBXHqimNyt9EzUS6BntXN+YD6+cebuPVjqepQ2L6MjUMbh3JfLiqfBLj
vDye1xw4KzEH8iLJreuNbU6Y0Y5vXEsDoG2sAljs3IXlnOh0YJr9+Nr3lm0QnjhE4EVjPesNfqot
ThbUPl1dcTjxrJMsYFHBcI03dI9kYigXQ7oHWK2PmRvXKLOnRpv3R5OMaK0BKUiZWHbxM+LdSkkd
NM+Fp3ZC+asDwAiOJ8yfsUK7GpHhLhBTKdmhVNiDx20/ML/6tM9/7POMzkpR3riux7aaD5TM4iKw
Lq52/j5XLRJC7NROPzxlVU0osnvX5VM1QbI1ZCj4YW17sGpOiuNt0xuopHqNKIkjnL4y0yZIcm1U
VW0NXn8DC1/yUUaSd/lBwIXmyV+L24VdvFwYwtOtWXO5gL1+Pfr5GhVZsCHkT2jnBRdbv0mqRS1F
S6bRchjl2MtJRgdguR9jXpy2UhxU2RCvhTG5jlAhGTHcHZ4XjYzZiK3D/IPUIt2F61Opgbj9xooN
UWD0y1XaTWZ+ZIqfJ1wZ5VdvkNfceOVm/mJid0iT8XP5hsS53+B6TPzv8dC5AmjCCwubYmA93Q1o
Kviq8hM9qyfdqdbFMNUvhMCS4D+PxFQuVv3RvKSJk+4/yW6RcBVi6O3ernnREtkzEtQsxzQpMS+i
7JeOqSFE16l2itUU9e3emDdyT8ZCpcj8UOIydcherLBgELg4c1BRvvVfHP2dRHJlfy615fGDtxUZ
KzzmLCh6CzLYn3RZu9OeSt3NKo/hgGpWJl6bc1zyDmSD+1B2RzrBj9ztS1nbzkoiiB265u41ybo2
iOjx1MU2ibRrTLR3IcSEJTmfE4ZQusfIgVZ9ZoUyE5yZAW/7qVG6878Oefv9d2QSmslfLLQTFJVF
cEH5gFjEFbvvO5xBzb/pxsNDr/uDpK9v0K5LAx3z7FKejqkFluHUPQkb1exN1cMiCgXs2MtQxwv3
aZ7YXWwJtXslAysqaKJBvaz9OSVDRXwjPGy0fav9541b/x57/vGevA3E9Gla5FPCJmllNFSfxFGY
D5T6uNYXJ3Ole5dW3f/pfqVJEFCHYTs5uqzL2I5zyZ3xu90udDEB81sXDGsOe+5QYCy2o/pxK/0M
2JP/Fw5E8v2El7E4QKWvUOiDQO5z6osFwX27EzilSozoLoXnOadQQHx6tzrcaqz9tH+wM2bCrVem
/DMzqJXTtDhmdSU5VLvFulUmQM9seC8uthKzlzope5v98GGVeoQufNfRSqbcxQEhWzmXh+0HHoAx
e7+HpjxUDQbLpJmwW82R19FX2liFdAHrTY4RDHZNV/8iRRvbvyMcBGH5CVGlPzopSyq675hnnl+x
0AlgT8+IE7Pz29ESD+qSwr7iUJUw3eeeF3msCKPCx/toi6Vyu454mQseIdGnwEjVpLul3ZDytSuP
igCtUvB9SR+Z8RPzqDlgXp/wVrrZg6dZSUwVynL0JrBL3kccH3Hy3G6s63/vRIF2+L+PUSd3JpKl
lqpbAVoY3pnaYwtGAr3PBv+Xii6G7qh3ZH6U3fXQoTvLFB+iFszENkbzH9P7T/6XEzg1ZJE1EQVg
RrG26/LJ7onTqAlGOrAlkRtosoSzbG6g7wKVRhco3iro1ty0ZWS/exNkszS7VBLEp3GZAEJGcsgZ
RL2ntwAkTjZ6GqlygNKU3GJDTb1ivZX3EmcjJZgzt/hPUlwC4lQo+tkSV0Hg6zAYOd6C+Nnjjccy
G8im0sYgcBfrXXX2F/suC4XlTZpGZDuW68U6vguxiCOFCOxBMTu9EuhbsoUEjWYJ4yqKxQNOBrwW
bSKAg+zctsFRTuiJNlc1UViswytMAXW3Gjv7sbdr1izlztukejRzaTXcSAcOKeKE7Nkr4JHHEwkN
r/UBwsUPwnx6loACFFdin275uSIP1wIDWFPT7yyWBav22i+QGthk3t7B4VENUX59kTx4cSLbSrz6
YFNuhrbmT85quEQx8tw6X/uF5imWtbxaPUP2/PvdwECzQll3IVaVgxOMfS3kzwgGolYTGqGA99og
Sw3A5Dt0UMqKAhSNW6/V3IVzUx3Wl5EbmPBDsPiygKIgZKNiQ6Symqb9gXf7wQ2N6aDB0t1a1F7Q
jkLJuXQa3Tr9iSmvfBC+3A+ykv4D5jD7IR5Y6JIborlDvyRvHVe8SzHeDwjja6P6fdbQNny+wWdB
uZsYXag0YjpeWB9AFmmYqum+Oj/dcEwBtouGviKLbvR2CT+5zOk/dfT6VKdpHSfGJryHEaoz9gMn
uw9Nt8/vhaWIfFVVkQIWdVkrwV0D1lT1ahdQZpcoO4OUGKqOwuF59vnOIPhGb717zBQB15jgKFX2
LMg2d3Mj9fXaVRr5f68DYIpfEcm1tA7KcR9CSzID8vHZwYkAsmilr539576eS4n6ZOIg6Q+inKyZ
ja4rzto/6ELnW3g0n8rKjp7NBtKaz5dwyMLWSVMC7IIqew0/mQ+l4DtclgsGRZfQyhlQLDF33CLf
5IbHMC/5e9YqPhx6ynl4nt5toZgP6g7x0dqYzxz+rc+JDzJ29CAXFfITUA01qO98i4gq8HhOsHVO
/wAj7kIJVu70TDkli/ppbbKujnvwG2M9aTsbQnOxoPxaZMsmM3z1sbiaLPzIpMYeYZ79ispL0WUs
VV87RBaEKZg74FGtVe0qF27UboPB0SBu92IyS04o73NdsFbnleUPCMIYcdtYwJFnV5UET7Aonc1G
aDEDz4PuEPv/Gik1oXFoGjmvjMeLDfD9ZiQaHFmIBJ8eHXTca/rNqxHLviMlK6LS1LDHBGbSnWen
A58ifZoQxES2CFsd69Fi9oRfKUPImnnA17wFestzfipMq3yjeTfrsxBUptDeq73VV1iqnWnbt++Y
hLhp4Yq2CIVhB3EyN+6F0EDV2p103smTuDdRZXgM/fIUIuLnJhHKoLlK9v+s68GHpdF7UCpYDX4j
nUlM0CMRvCAVD5A+mpWfhMK0FUuSyZeK0F+lijN6qBJdtVSim/8uNwrOiZB9yb8crj+hsbqaQdX9
GFMNLkW1qi4YF88nIJPfnhBMpAUSqQF2B4qaAwCjghXgwbyw4A2msdOAwAqlzsNsjVA6H3Zt314A
azIOt5LfhF6dE61s81zNfxSGHDh1Qf3bhlf8UcjBnIiBI4ZD9+vZrymGXJvJbhn/tqiAkP5V96FW
UoMEm7DhxTLE40kQ+XLYtmRf8UDdGdVqjdGE/Vx+hnULCmCQGQir9StuYYl19c0cBKwkiR297vwL
Ojjwzd8l0V82bsReJ3oqhxipu/efR8Wvrx1aXFMy/WbCJuG6zXsNELpHiCnV5RqfH1VbWNFBcDGD
injnP0jmRCKqUQxtJIh0YjWm/e8+nQHtpMlxpa0CZ+gPDLvKlthf85kHFD5+DGcuyNv5zfOY2n3x
n2PYntJ4lXWxk1R3+uIdWW998uh+SMQnb/7OFWuiAL8jgd07B5CdHYW1CK6u4EzRX2wq8S770MvJ
KxYiQlHbQwT0XIGJ8071fV1PTIk2SCYEHIcb1yN/zu4YdeKvdFpprKUiNENV58+6rjMfjhmwXVBj
nnmQjsG3/CjWxo8YioGPMEA3AdKNswdf8v+jdocV8vQjPx9aAoqm83zD/0+WZcBbmkHmN0vRKuBt
p+m3GgOCTMh6zkTFAfsCQV7sniD/HK9Ci6LOz4+/j+YSTGt9JLlavA0/2SBf8ikzlBI4kGgGaBys
quU/Syv2CT0kSPI/8CDZ7vOZ+8WYtZvt6N7Qua+qTMeSsGTYkjPZ6edHrckJulpVLh1jizlxZu0b
niBnPUrMu3P4iUSWHAj55OAqPf47dA+C3nRDu7hvjwBdqwZ6w+60tyb+IGsBK0Ukm7nRi8E4ywT4
bJkuIonXZ2T6SrGnogiqUKAoy0+vzbcegCTXPMouDb4FSlMw3l3iotsVszeVl8O5o7r7RPReAxYf
JIROkDCUexVJAtDy+jR1rIpfneFCN2u3JOUR7Y3jKZPvUeJqAKn8sa8Q22XKFXMKQHH0tzACi3K/
zDhsyHHK04OpihFFQY/ZlBl9mhmFHBKNf8Ht92y/+RnkuaaKa8vzTIzq6BeIwPZzOx01y3hTfhiK
o9sMFRdykw+8EJf+vjCnfisLx8w7L8w2+2YAuG6xDkBGmiNUxthwVH0V0bOl9hhCh47Bj/X7xvcy
bet8D5s9PwwsEXDdL2Dk01AwSer6SAfcEYQYBNA5YVT9Q5c0FByrnTvU4GS/1Dij14tY/1NCRXjF
b834/71i2ffGFKq/XkR8PC9turAUB4bCEpBkzfyd3X6VXofsoY8/y6FS1NMGY2IGl6N+hlOEbwKt
XvJHRh913+p08wJovPciY8Npp/EDVP0B/NdTgeJArCxqiJqbk/hkZ5fFr3g/udLa8ETGiEEDGd5m
+E8GtXTWEmNc7EOh+yOE3fCJfznFndaDOLtl59UWBBqmCMXC+r8hC8Vx1PY0WRv3FlbyIT+6iAi8
n5vPDSGvxM7DUK3Wq4PnLCqDtoKZKMn/lIPSgb/QuXb+y7YVWzc2OegpLOhilryG7RhTF/eNO0Uc
TLaaOy8gp0dGb35ifYMXFiyvIotLKodQgcOhcEzVLmax3SaZQ3SCNCA9a5UpNNP172oscpkG8mTZ
xggNaAIzx64ch89NMxsY5X1bvgPneO6JRHLLXrL1V1Ol9RQKTO8+wCRx+tA8pAq25qye6JQBxhhs
AX8kg53KIiB/gmtDJJ8STXjy/NaK2cMe+ka4Uwn2vw7SfwbQNWZ1n4/iXqCJizC8H3dxAZ1s9x5P
Ofs75U7k7b5bliecGAdEXxfg4XtxpROjtGQqE4PE1xEQukAdIVjIiuG/1s1X4pfjm94ceuYliklW
AdhpKAaYi5KapKzH5+KgrFrI9JwDFC8rAoXOiEuicRBxFBpRr63f+8G0syNyIZtHvJ19mscg0SJn
9+LEAGjFEk8Gei4feyKcVC9VVqX6/eBEwvYu1tTioOq6W60JdIF/DK3jes0/Ualp9Cb4T36KJ6HX
QOjUQMHTTn3iCy5mDy/mabX9CWP0Wkh/VYwKrN6xXC0UtavI3MqR+MkVS3xSTQpNO0qZHoFCYdPK
XN4EAki3qc8bycf8yJ5yjl5T+YCuyGP929cRk0qE2YgvZ0pWeiccdV1KNSg1h6oDsO6FZJq1cuwT
0B890DKLCQA3EfJau8peQZ/pI+xd0OsrKwlQMUXbl+Bh0PmygXZYOIUejefrCHtS+axwaa28DYG4
2kwV9MkyUymyQ6FETqyjMXHXzcgHhEf06NjE9SJ2wctV2Zlu4soRmAU1L6obP6qMqXMKHRMeADTg
TJtYYXvkhwIym0yaR7F820CYfwyUlSDGy9grtBT40ysgpAUU2JcZSr7VsCsqC/YpF3lwNS0hOGFc
0h6xszhVk7eV/HreAZlgqt/QlM9OHeEm3tycKDzNinsqLH0Ia1WPdeqLXpPg2iw3xVWsfIbvngdB
s0E96DOPKKm4WbveIObixvxH3WT+0KAIkNj+jY5ZTp2fmIiSetHqOFV0BgjsuDOeYnXn1j4whek0
cuOheA/i0JWiYtrUpgr6xpdDTNLZVhbFcsPyTvOnCj9uBmPkPOCIqRiz5+JPL3/0NCHZnAXn2Qk/
9zTJhe1xu+IpWEjOhycaaQsLmZ1SYeY+hMXWvzoume8knrR4eHa2FA0oWj8wNKqpA3S44GINALtc
9Pd9XQySaMQ/pG2mP+h/oLozLgA/QapnWPnEnDWM/FACHnfUeNvr2X0o/d0YnR739XE4L8RRmHJ+
2dDSCy/wzNhfKBEEH5CGkecAAgBMVu4ZWzsv2MeBUJKYpZl5jN3w0d+UPC7vkKVmQqqPE5O0vvo8
NBCXvv/CtfCTpF2+XK+FBUSQS1OORbTOEb7MHs3VIoMbkYQFUnfm/HlhJUU4noRQQYhfMzY5bmUR
VRVb6bMtmpawLMlupAiTpwd5Us9qtJpHR53ekNUd8wmGF9ZQkl1Dl+Rfa9FX1GwXtb4rMbOxsBTU
0NTvBY/t1CD6qd1MWOlu83UvKXgnXzMSLWk92SW9+JqkewiDQDmoSlJySttMFQQzGvq0WHAjR2zI
H8T0pydO1LHTUNSvLMoOWApKrAqG+qsECbeAd41dpuLdYk2u77Y2mmq+UgO0Nyzn6sdoOxPm1y+s
O+CbX2QpiKG6tS94em2hoKQ9wIyOLb/eEANMioD762XaZnkMqOcJIsVfKXreFON7n/otr2G905gA
ykOaXqiwRLA6a+gWudENbhd3xtFaloW+9x6HP6YDVgbkSDfNplZvRn8HxWRuyZbAPX3QjDKjNd3E
8FxFt1hDKm1RaTdFg4DY99oal07kGCHi0ZCNmXZ+XZwWmILUA2FlsfArsLdIjNjx3wKjBv3tSsg0
0ARVjND/nCHrFYPSBBZAcNflRtApKS+g0lHRfl6K+LvID2tKlqhFMnUy/q24h2mCaKs69/ye3dHw
ZpdT65jQbMoCbekUJvAiUnx/1OGm8KeABt0qPh/Ur+cuKZD5MRwAcia/Vv5rY8JpJCt1m+/8QSss
TTomJQYdg499IjWYDffRy+SnbcgcIj7H/GjFH5z2XZY2pQJCW4vwg7qQzMFcuzglX6+tkGODywJ0
H9FEJcZi1egI9aLVhDjPMDgZMofHHH25pwsMnMJsod/mM4x+xttIzwTOyVw6g4h5+8ynTz5BcPEr
K4A7jcgVqpnkInCkfPVWD1KogipBVR4DwaHzEnNaBt0H5baII6AFxU8/uX8h6pH6/29WmYacnntV
MEhcz5uUZI0Fakze5ZoLW/mKAVbfuWgu5q/+FP+zDjBKKJgnLwgdItOmwXvwPG+qAk+9DdkKANai
xbnFhBY1hNm0BT+vEb1MdSprox+noDRq176x0hm9Z1UAcQLUOO/g0MNarzAT3WZqFVeELa8fGzzP
iuMRWLRj7M8d1lg8uJ7PXNyvqR/lTSR/aKAfWqcEvE+1PAh4RwhVBVQRsEQPeDCbFtp62QH+FPh7
Stqzy3y+4uGVwUPFqSzOay9AJL+TyHyUVdLIB3iTWUUf4KwcKqha+RvPZOIoDpyBhoSjopenGtGu
S36sdxTXXYQVBdd8C/Lt5WSXzc+sASYIfFqUDkCTgt5qdL1TE1d0cic2z5125UKa6CVPvdRZdvot
b+fuci8uP+CPbmrbfrmYH6C4fl/Ko25PdXPJ7hYKhnwyzq80L0OrRMV6X7vO6YDhfEr3EsTJ0dip
4wkiTQM/MYGWSsmLCO5nC3SNKHI7qtcCke8Cg8TDfdg28fFaRUlZR9N0Jc66fijr8lqfOBUdFQZ7
bEVY7Zr+Znc1Q3pgXUNKEqNJVSpIx9Z0kRi7yQT8CEP+i2HTtD9Gu260D+GFrgrEz35hkIyHEJJ6
MRvrKB6rFTlJMht5P6ND/5PVb2/ckdOCkXsZxTrZ2fdPUwBUdoHzD7YxGvA22ElLmE/T5qdyS72Q
2b6o0xO2g10opDZlbK4q4TM8d+GPXCgYex6KvM9u/p4QmFZUiXylAe5+1olxKtlL+Zx/GWwK/rws
b5+1LbpbVN68arj1pHIajBpHHr3ZFm/ZbDJ5tWOuEgcpSObI6d89I0GpYQ3OgapgifxMzB4x0Z/c
U3itMj/HBSSidnJozxmk6Y/uho8G/XSSxBD0rIxaKKfWV7YS7L4RXuPTiXD/eQkzApewTCcmv6O0
fJnNxEQrg2P1RFEEmxnccTJK4+nbWM4RETJ7yNd3LCryaCSvo/q8pOwazNcH7LrXNA1xQRKTzL4T
g9cBwVrOGpCFVetc4g4pC6Zunh7akderu9NDv0HPd0JkGkxwOeMCFZBUicOVK+uVBZVSYSZt6PN9
ycA2jArbxQTSXKzRpiPHSqdVSHgtUFyO6kM+nBCOxkhiQmlPLYv1lOjygqzFo64plwPPBwFV1R05
ZCKiy/kki5yWIgmOLHpDS0NLkoJE1/9u3X37E0wCg7MAVurvq7My97OG1rh+6nJBWPyLThBx30xS
59rfWXUvgFs5xvIzqloRDJ94vyc7eNWJQUZJGVCx/qHqEln0NY7rNwUvxkdDZTQxVYg7FAv70RG9
CFcIsEI5j59udiUy/nO4WgQMDFvagahN21rzJ76jnJhaSQz+DpseoPX4fyMOUy71a/2RX0Qnb5XA
bwt1EF+6oGQyEilw+IYxtHDMEgctykoJXLhUnsVFXLqnQEYYOFApnNOldOE3deSBUUmFALJaYdY9
gRCMHZaCrNBa14do3lTwDgAZLwzd7jeqPGstsQQ2ncIcF+ti3onNc/L1pUsRHvBsWR/09j5iM3hQ
fC11mThKpuR/okpXOLniq+/nIqsRGHxi/iSAyjd1SahuFmFgEUCOaVJ8cubZdyy2vUsXaK+Gr4Vi
1rz+KUI/2vHDwZJ6TYfIv8eoXX87HQJlK7pAb/bwd0Tz9pfejFohRx1TKR6ngG4pbUHyBiXSInhD
bwqv6ASbhBA5ynFIiVhI8Q5QtACCKdHtY50wom7xxHQnY5uaRkllaIzXZV6sdg+8iJ3MwGnIx40y
FDoWv8hf/UMjd/uYyrhYw6zUPn6uSAiy/x/2s5FiP5Yc55ucOrur913tC0rPLoQQOp6s0twlikei
6ABl3gEa27/rsajTtlYMdDSqKMDGmUaRQpqOEhJuxrFpaVhIsTqTW0im3CAUQATxJ/qUBNymvbwt
upKNlWSdxgqHmC2VzUJe1COoYUu5/RQIsp63mS6P/khSxmfYrc0+04oHwD7S04B3X4RnWC3EUE31
rEMKkInho5ARG40B6k6Gf/QDN348ElZTWo0ukRg2PxSifb3mhZNxB1VgiiKYsyPH25NqmVzXA3D5
vVMoDUfjlSvxiioeX8BRUyAw7rZ1wzOVKBLWcpc9guyVIbf297OdtlDwqxaC2yB8uTe8IQc32VG7
4IPshK0B6sxqdRkYn9hBL5vJEwmMT6iuOltsTVePXzsLJQ9pARM5JiwWVwQSkpXr2qlqEREZ8Qf0
n38jnGLFSlXRW9TusUTJJT+uLyY0++zYWu4WEQggQeoqN8r/bQplemzuR4JRAw5UaS6JOnpskNgE
BCOGYR7ykrQ4aWt3sVtjYLaP4FLEPHExUqC+TOrSXQrWKQghmc3pxI7UMsrPMg6PVSE/LmdDayQm
GNFH9nmdtH8jtLf3Xx5mkMn9cha1y0XRQlv+sBdCTQbUzt0oAYAvNOnbbPqze/5XxFlvkepuImjS
mMw28GR4sc+1zUb7+e7hGkXU9qhoigZMOHhSXk9alU9+xILlviq9mLk/CzAGR/GcmQdYjuboyrlR
ML2tZjLgUoV0TfWG7cbmS3WC8FKyY/bRzOsPhrN/sw4WSyPIdsE+9ZZa8hpoczsGVmtNJzZM6nfQ
qxM/QDB1cPL9r5rnVTcb9z11ddDe0DyBAR7lJZlcXN6AY91/bM5rcZnjzIZjJex8oeeaUnzdK93W
Ercgb4G1OeWrr/4kMYqjXfMF/EDlRK/MkquBdOL7KrvNbX7egFPaDeOC1F8D7ItzOPtCYusL31dV
WWcsagb+wB7gE2KPSZGSHrcYSzYwgAHY9+/tAzuYIuGMUiigny7OrmZU8vX+NLwSVVBWHMgkhSGi
cwIYh1cd0zB3/avOP13kNteyz4sSkzhie/9fndH/yzTdJk7sOXStviWXwx1Ex+aLbjuKViU/EAme
YFt9Qh0+qd1JLMBrUXjWrbsI6Q2NqL2uTdmjElqqmiZFgJfZ/5H2MfxWuUyoUMQJ/8i/j9RTFDGq
67fH2xKtEt2xzc3a/HKV/BvXW+GbhKWhBDwuD+rEHqz9bipn8/yGVYixW5WsYXzqoh+1WOm1uF4/
pm1fpjqjijDmjJ7iyI4iZF+45+48B5H8L+LWYs3ZqYr1fi4y6gODt1D4+FzbxYy/Fyj/uoeIK8YF
8DEPr2JzdL/0q6ulh6W4hbgSQKQagBtOD+08o4Sexh8dEcU39ALe/Z7KKwkiQ6k3OkMcYxah9VKg
+lsormu+0KU/Lqj2vSDlPOPAiIwKQpktaEQ0dQgirFKAqSBAekq28H3tMJ92p15J0eIzTJNjzvsg
UDPoeTGcoH1P9xQTbMFbyuQWykJ+Iju11xeeFK+vp16/y5QP5junHjLEv9gXwrKDyN9g6GkgKF91
IFMoNETZROZgkXIKrFFlT/UufzniRpHa1ZRrRkxRXdMbuXQlHZsPc3mcQVd6QTisuJ748QepEh2I
55khPRwdfDLee1rkGkkb7I968ZGvitk34+tPLQjs/UdIfEfaBegPfWb6kXwns2RslZUNum0uLevC
AZWhbEhTtcoM771+3Z54NB38hoCOT5Fj64bcCX8HJ+7Lot8OSP1yR/AynNfDEBOHWp6ROLzAhWOs
5hBGUBVIpHNeXUV9+crhU6h38hJY8U6dEP1aUWi2OLg7Eza1uKvifhmLMRn5cKNqQ4sW6AWLk/xK
ONV4vtS+DWHkjVDiun098t9s5JKgtitAKSbl/jaJIiWVuRqWyHPofWAnGP8ybRDGlv4fgQdz/Nn3
bDt800BHRn7bzW8X0QaF+NqvEW+QVMjkIGM8voGem9J9RA0pi/u++Ojf6rF/v3X+pM2IrMc903Wt
oSrBCBvlEnPoYpIMMM2V3xZdGTef8z1xF2S9bQUSsHEhXcIabZcxJ80ilJSOAh7nPBHrrzRTrRqI
WCjQjAjmbo1qBBSOEnvoDU8uVc4k8zQ3nAyUG/xGXYK3+FXrZoyOHmWnlqjjdr3k+9kcVUnsNylH
C5TaMRM/8kPV7BPW4jn/4+zNk6rwEsvLzKAoNmPQaH0s2mOa/A4V78b8Q6jW86On7oh1R5A8Mnr4
JSdXrP72h6/IIDos2U4vaz1aVuCJC4LNDwJYWlIlvsOd9x9ERzP1kcBlenzI0qMYdv88OYVfFGwu
8PIBsW61MI2RdgNDk5UmYj/QFzeGiuf9Izwte9CJaCNGnxc05ChpcBiz3pX7CcNp4deEVZLR9SEQ
wuA4MWKyx38smxRn+Mg4Kn5NRo2ZNg3jEhldBpH0Sx5GHkxeFrhQarolERCmrwFw45orPDkdQQLG
VJyo2Ry3rn3sGeseL07EjV7RYRtBZp9hZEtI2MyVjEtJctzC2awMxOfRv3+5dIHaa1OjLEAzvKg6
2//wiAGwUKIFqRQaTRcdb3vUN7SsEAPNtTdYzrMmqcQKNF8AKnvj7q7/Rafl3ta/LiUWmkTeRWuU
aD6gstv+j5KZqjTLOy8x1QqHqSYeYb14AhIwwoykMMJlPLuykjTj9hwHDI5twFQTQ6t93FthBzvc
Zu0lpM2L7nGhtVB99tdE9No7uYT67vFSWHgb4rLkgSbZFJGKHhlg4HfUZ7g/FImbMZFtyEbHKIWQ
R2d25aNV0mE+yPvSc8B9ivl6IXdMJ2iQJQw6r7yuGOCcN6c7JwA0Dn68eblOK5GkI+lkkpzERAZd
CoJCVjhUK84wUocwryPELYp6t/xhUb1DVunCBR2PDk6SXfRLK+8ajkksTyD9NRVh/pu7D6CHswRe
mIof9BDJQKVaadMRNBZVYyaHTEKDhHnwWBhnu1zvxhYLiakR5kHZYxH673bROITClo6SoIXKXs+9
jlIER/13BH7Y4HjkxE31U6MFRwWqMjEjJzPZTDf5qSSbSZyLzGH7epO5DK0AvAW4gzni10ebTeG7
d2WOjnwlh1X8vrW6Fqr6DqPr0cfdo+LYr9zPSurvAb2qtVx6v9RTNbF2jdV9k+gV34C56TNGNL7x
ZHlv5m000e4OXKVlQc0fy/wueja/yzAr5vpHcdoTfZxrBJ35bhUp3RHUTJVRImVkVYGt+Fqgr9n9
BjB3br0nD6+gACdHPj043gwuBT055kP6v1jwzsweWDVJBOwW7WbE/zC1XupRl9Ix2RQE7RTN1tIm
vjyYbzLv8VSaMkix/Bt8XKPAMDueC9h1qX4b4Yz/tOn4bySVzbY+IehtWuRx9AdTfPK7YEY+SJMS
iYninVPS3nKCCkmJinBiqf1c1jwOBw0RkJFw+4+EH00xU4lFVzHTtedhLvncSp5ir/ZA9TScEv/k
m5QOl/wxY10VIzVOZb+PECZrAwsWU9ysSJyji6kl/gDPivXEXunxL6qWHce7ua9b8S0FwTSkZb80
t7gmcTcvV4YAS2l7S+8ns0rexgATLYW+pC49tpKm//nTbhMJYSPkwNdOUtaWUg+ba+dqJL/D9mqa
AzF670Qs8OYn8e/xkVDKK0NFeLElGV57hOtOAGmCzqWOBul3UfgcMfQxqkbEijykJ+AJgaM+VOlT
yYEtyHCdGMv0DF/nJzH+qU4YrI6gJYx9oBIHh8/ugt7MQ47qF7+KxpNl35l21eY0NBV+qvMn2e8T
NXfGiu+bMc1OsyYnMn1ikkWjp03Os1x9Z1y+Y8Q2xiBsiHIrJmtat7vQ762h4UsA1Ce98dyu3zju
I4PDParJ2hzSJ3mO9sfbtmSu8v4MsMWXvzsgHyGkyNFW9j703T1RIvKmahbNXsxcIcqhsJexOO2P
neAbV+O3CeZY/uMIz2Uu3J8MRkWyGqh625aHgtKgaYySr5D3Ynk0H7kPio4Fpxkoo9gAdoxz/ERQ
yQEY7GYm/R4H6OSpkenoF40a1CU4Ft0g4ihTgvT3bsItv+3NQKugKfBGQEz7nTXHNxPpoMqI4uD7
7Uf7aiME1N2LPCUFnlID46M4DCvlcrvo/oYxJ52jVc6EmvfvuTHh3L81HawhIR3W9JsCAOJvbwgt
n8Tcxxj0WFkASOV7IcuHYBWbqoddAsr9N5Bt4JG6LitSgx2GVej6TEkZ+m3mK4IlmruzZTgepNdM
iB+6PEaurcm4USYL6Jkq5w6XhvXZcWOcXNOU/5ZOtEgpOFNNrt2XoTzdIAoz+S5spjdq+tf4IO03
1sImZD9nuEYCCYTSzhWPxdLjGzaOKCDrRw03IO1/5Hc/tv7VLo0DwpCz34WIuQjFVKSByiPtA/p4
Utk8zy1oB1zLVF8RXhiTb6G25OpbIvdffEQmUy8CUvW4S2oCMv0N+0OvDSG/cbw6cvbbzZQrz9Os
fPTDUHKMg7uwI+xU3JmN7TUo1qw7JulFbK7ktBLPh/Ih1X8CHouo7QP67bDsGB6GX0F+TSAxCNPf
XR00T5R/kgmLPgAZWdFj5lZmd5zyQ/uyJN/0GRhUBlYMd3zagedkgSKO7sMhwDDHHfJtG+oeljBK
QDgjAqfoGXNN8blunmzTNrHkHm9sY1m73yTD2N6W/Lwcj5D4SD8NvOpiEw3x/TG9iMCYZtM64eVO
A8ipSaExlKz8wPK+8YRM9789nEaFp2o65Ne9G3iFY9/XuY35K2njx/7oQTRY5XhKttpc2zUUELh/
8SbdTOQXARUAsGG5E5Q9g3TYxOB5dflodXOERtpeStd86PQOwtH5pZ6jgzTWJq9yOdnQiw3ac7KM
+iNsfgbYNdUa6NBCjxM+IuTUZvAfcK47cRvEgwYRYLlQuFr5W+TItKnEgKNmGtZfDcyPMu4MtT/e
J6Y/gWiwGyUf07XeYvppjE+KRqM/ecQNHl5UH8CJuazRLeuyOFAXNEQck1DfYw1Fl08jXSwNcnfy
RgalC1j2ndNs+qhNmJcptaZvPIylxnBhuRfLjt5wbx+nBGsSR/rQllHmaaa4akRH18vH5+zKOIuA
ahQjKWsP3a0VjnPW5NdNWSAKKJZtc9K1/mpvVYUAfuKKU3ioCNfJxeTDy1Qkdvrl4jt14TsdtrEd
8MrjrS2P1nLPdkOu7UNuH/U/10lPmgk5gdes60hh9FY2TYgBK41cXVUUeAQCT8CmatcIvABZUGEJ
e1Dpg26otMvit81zVC+xX+9yXhSfaH+GmijcOrQgLkxxXIueerrooTHwuEHzzISboBic7bobXE4x
AhuIvvFZaBid4dqLtxNJXzJSq4/iAAQ3fGJuLfvPqyDdbKRJ/lEltomOakhN8nnB0oFme80CYtl1
JtOn6xQztLdoP2UF7MbE+I2E/z3/Lko61VBdKbxqoW0DjlOf+S6N/RX1YT7A9rXLmogb7kXhE8Wj
5JqLXCOscxHRAxG64vCAf0RyD8DNbHLBAMszU7Z1lWRepGo3SfZFo95IrBUGIpz3hD0VTI59ahZQ
j8dhN/o1qKOkSbpmk49ghozzVzLNP0HE9bdg4wiOjLXg5Qyhag4HWjgFHrPrWZb00XbuhYe3OQVa
Cg7JFPSvudVijf8ZX6K/Nezfr21Yefj3OTSnrKOGwL3vqd+9PpFY+jZS/A4sFKMWUsysiDWFLn62
e830IywlXPzpJnpJnULhgTbvzgLwcBKOpazPE2yx+bdGbn2XbF1hFJq1M+FJ7A5QYbRzfrrlZXXF
EGcx5qFemF96m5+0MpVYrdj+doy7NKT3v312S06/GjXJfzEe7xUxqjCnvuynO2xK29Ld9AsKAFC2
1I8e6RvVVE1AeSvwLwDUWp4E+vhRVi/0csSQrTW9mLV7J8gLFIXfpD4owjetF/ubZcusfL2+CNKm
SH/ZE4cB5cyHO9w7sr5dwbC+ZuxRYLRi5Q0a0lCOL/Bavyu5GmSROJ5Ze1fLKtAR9/3ljPNwkqmP
iX5osKm5Oqaabfjzi8ld0ksn1Ad4a4uS0LCGTC+i9secPn9tDRnApOgKvnL8ILfzJJqTkbwa7HoV
PDnMEDdATT1osp+U5eY05K22fmVvN9+Y+TXljUsVzxbtxqwgrSIukpYUDI+k5qxcqPjeqHkDrUmO
RfptcuhTGc4KRY0CBpHjF+oEG4B5dvKPFzM+5vyLZgFwa26xRvBZycdVftG+t+qiOAfq4YMVr5D2
RnpVqPsHlc21drOFKXWIj7dWrFreKB8+J5ihwzdDjk8zeB2mYZ0j/DOL41zsBA2AuAqXWaY8GxEq
aVGf5ZHzjSN11rH17s6PB9aYkGoWRhob2lOJF7woezyUcv6kJt2X6HDp2A11/AhRXVUYgkRvs/kh
Jgpi4Ow7NFdQbeiPktuBIhZXfNq3pbBuR780RlHEBfXw6yZGWeZf82zarp6o8taDkctVRB3z2m+8
gpiUgl3g2nUELF+LlKm/3EEpqcG99fxmN36Or6Lm2wz8b1FIkup8YJTC1+2YXmgeHqxLLIKlMWDW
TFv8P/3x4aI7sO4W58XfT1SBocUPPu7WfVw8U7HeUOSN4w9Yl96PM8h65Ma7ZaiRbDiYZsUTFdqa
VpzgxFP5Ii9Bjbvme0JcwRQuwA2THc9P8B/seqkbv7YLdmJoY8aEuCYH2PAu6zuCD6K+2LTjZ+T3
LLnMIFZHo+lvcwTLx6/0vAyUFOJcrkSC6W/LiOXIsAbjDOVmFP/1jObBH9oUtJbJs9PakMzBwlHZ
DgJo2hprDQ7E8NeqUVSkLRM+v4OQ7vYDyblMPW9p7eDOjDxUpHLsVlKd7dZlYagY8x6mz+G38fpF
zcGi1sEYznOtKjxq15sUue7x00IIxGUdJ/vbrucHHrUDiMal9u1L91J/DVkVECBbvbMqoGKB/VXV
MdcfZrArNt2ZKV8A4zMFz3ZlfV9E7OmXHVILx8PutcWWHWySnwVH2aO7Zih8waLQOZHk+LQIGae/
dS1P0sA1XmtyzMYdsRB+NCYQOgH5WIEJAShL3aZbcLZ+GVTY1f5p1ShMxvjjKllvqN3ipL4lTcTp
eW7YVmNupyKhKnCQ50gkM5tx/+H3XCMaAqZYqCTArY/tUM+bPlZWGq3bJ/V7kIap+hrrYjWXEVsu
+h/zvHt4orc0+NrxG4D0sQOWMrBKc6hQdlfvRjU9p02Tmjh9dfp2GMdQdn9mE+puCv5G9wWKZxBX
HQYcTPZfAEylbLT/yyA6Gu7cJuF6QWwHumRcp0DFk59XopzPLxkE27DBABg5jYXQ4ZNwrq+wuKHd
JyR4vI6jUSkZ4a0s+8l1u2wChhiIKkzsnl8LErpBjjnVhhhLB6TIS0Wzm8P0H21+AA9jEhYcQLxP
fPQzsIFP0ooZkMX26lGJh0n8VNqtxwrBNWE4y8P9PJ/INfdfEOht2Rl1tHtt454GAEeqccVCOby1
0hPJiMDWlWLY3AqKqiLuimzdG2tSZRkquNw9ay3DLusQ0dm9YsmjWWhK74dEJ2qKB+xp4otIydaA
BmzpNgZACrARaR/MQc1srD6G4/b4UPxvv633rKYFQLkwxqxABdMRxhVogCimTGbYC7xqd9IwFPpU
qHlZtIIst0KZscvaIHCMsMUTuO100KPUrjJQRjVB+YNAUM9VPHTXb+Qstkqh2pJXYuXsFiGzkuMx
e6GMGSMtyDdtKNBOLoOjzN4PqeflXGYocjbZINuezznMgEBckmQCN2MQABWPWlSKko3pAnT36iwd
o+O3Osx0qPEnp2fZTVhSf4HiLmxpE5SZRm58pg9bJzXMBVljIFC8JtQuGgfLAAPeg/Tf/VPs9MDs
HEMe6kCY0p/Ot+ZANqo36NflA+W82w074uaQkdJZsnqrGw8TKromyeratGH1NdHNrslsewQ1JnQL
TlrgrF/hHCBe9zzxxzgR+JaqxxfDKvZ28XDx989x+7rOSIDw3ic53EB+wgGvme2bf5vlS761jjyb
cXQA4ZCL1GFdnmWsPKnk4k21ZIhJOU8F4NDAKELhlZbqsWwKyqQ8CKbtm/hU/gVDQ+qFy8KaSYn2
rXPLo+lGC1WWeOe64LaVTw2m0pjUQNeIixwUq4KjtiPjz0hwcs6AnweCp79BxjHBfrnMRGeGr7+a
+C09JOopk4+OEMpZwiCkO1IDAIv2wwXP9UQMRtuL0BD2U7LO2lN3FgWv0Xy/e+b+X1mNUg4Hzb+4
4FmVNwudAg2kd0YbgN8RCmNhbKzDBbfp3bO3wPcjk21DIpnIlucz2o1GPtivMdlgdu7p6WbesKkI
z+0/dsAGklqLX0jgtboKTkk5DU3Cu7Q3YnZ4EEn38TsfAfF8xnsNt17rXNOg9fh8tj6baKBRA6tV
zN8IgL5ssyLVNcEHouPj5QmkeRTUKYqCCBIPC737XfRFmqY7yc86GVqNleXHHf/qtjSQiwc+rX7O
SKQCuDV/hTl83YdtsZrISZgydNmqVpVA/3WCigu/zNUPCIEDnFpUbenNNb4VzpyjDlJ5kge3boJ7
ufd9IoZhxwXuuIXUhxsi/Dl5qJDD0bAa6yvtQIPUM4M9voQmimYhGV3YAH/wRavTEaiec5PgB5rC
urBni7ZS1KHs73x3aGFSQ7wz7iOJWxGf4mtGq0lP4cx6uPkHT4D7ZyvKEx7ISgBZ98I1y1YITpCP
Ztg4Yq33XGLHX15lzjOpwr5RtYthC1rSbNgCwvhPiNzJepwGfDOZVXDB3CiHQPU93I6+28AXnn+S
fR4BZWweGgYYM3Sv6283HH0726wZ3AZpBn36BypKKM43YfgWOuuzrCII5+XNoC7fK14D0etSFm91
su+POmLg4BmjZ55ADg7+t/is56YyvPFIDBvFtC9hiedsvV0cxqglz5zVe+Y5NY/HPh/XK7gDLmId
9HgkZXOKaUjOWGlmfgfq5gRTfJCC9Gbl0ERbX8wlQh9QR/0/W4nYWHUVeVY31JdSq/P92GwfI5dv
NjMy4vUwPX9TVVbTGjwvh26pkRBHnmwnwCfWJ/wUDxw5AFyVOOx9KLgyy85RYjivcY2k625+AROj
jPoSa+XebeJxO8omKDEtknMGNtpyInVDHZYejn+sOT4LWLrgy9ES9s1jwscz4ti8SNf0LewE0qGn
rIiwBDahSGp3/TlzGOqhlvmLY/beiHRTf7m7n2XD2Ik8JJYRMOsm/hPMrBQ9pwM5adVxwcavnes5
P9IZz5dgrPI8GcDpeMb2nnilW+uXWsTtr2wFlFmxmLBP1HCV2aYKPdB/p+64pVrDcmaIb+RaYiqH
mf3m29KwqlpmUtEuncSw5E+djvpd2TQv6VSn0QBFdt5I0EqXb+EmeeWCq5h77++np016T7lLb/HF
j7c9ArumdlJc9oUeSml4AltM28WzSQAv5Or0MTDMCVwuAQsgCRFbYrdVJVn7aS7enB7cQfAqXq1l
y2H2s5M+rp4WUZEpbrb6FUCaWrNvhiXvxFQ/LoizT0u9Bs4bFfyZMeuNdh1Vb6tY7JMvCrgzLyzi
4Zpw0X5omS4Jlpwah3Og6LWNlJPRZUt5mrlHNtt208OGvbuNyrZxwqFgFeNrtLm7Sh7dJXhEZULc
zjW2vuwym466xQHaDjFd0SknCcb/ytvfzscFsD5GdWt3lj4HrcHHcNDiES8YnG/2N7wz01q1k2JL
ZO6rUQlGNc5tNERggTdEXuLbCyejHamlrduEi3tgZruk6tq0pyfcsXJ395AO1o6MqRpjfLr3BbHw
Apc9V7g5FFoYjXwXo171kx4K+mpVLF88jNc/RkcJvZQJ+YZQ5Z2HetGvUKwdEATIQxzghsrRGMwm
7dGMkG98HuhLPVX+N6K2hZwRSWMxe20T9vDwsl7u6V5EwyLzawU9X4WDfRsVuQa5ZJ+ZRV2uwIU3
mTwmdR5+00SsvRu1IWhwRErcMKN5ydwibKuyjYLW6zT9PtS+x78//LdfaqlaKL3uJDZzd/3unrei
C7mNKD8BGCAamfiDq0HSNCG+8prQWiWvDhyQij139MZDV8JPqpi++vI8KivfxnpedrMJgzltdo15
ZpeGnA6szJYODoJJvThu1bQ0n1Pa1bS8+enerZvY56VZHLmauT0DLM55Fk7uAwy90GVrcr/+AiJK
6smivnqqK7jBTHfNTkCvq4Q1+Wv/4mbdxhg3v7YtGXYd4SwCDT/Abtive3dcKLXhPxsBKck3TOaQ
7agtlCsbz1wNFEqs7nXGrC9iYSDfrWn8jQqBq/2UrBY9uRX6CP+Dzj427p0PDQQqqSahWYXdHTlg
RKmygalNC/FGWq5u+coq53YzPhRaNrtgAl5sz8RPQpQjJZkIAQFDFFqGn4hrdLggksCJK/pY63f3
MXd4GxArdUte5hqgt06JMqFqmdSkHivIqlR9QCgyem6zkMfHtgYwyKmJv9e9U3zOK+KGhKWH03JU
4/oLrT1VOh5HmI3Bhl8z86Uba6XFEdc1j6NpN/3gbOU49LtB/UMg+VbIiPyZnDGZMQgwqqdYEFwu
47aVMADPxn71N3pVzqXd2XaSbjnWl6OONgSH5XJnI+Yqj2pJP2U4F1Z2NYrBfTE5eDtAjb/9TTng
6cvEmXCKJS/xK8t5cM09/6u4Ywlwqb9ckDMZOsQD51mUmG13w2cbeJEez59tLmJiEsPvwFtzTIYe
RzGiGb6BpHg2fm9CehU99BRAe/C4HzIVXg6hqtd9E69/sRbJLzCPph+a8HE1UzDa88qBIB18XSYS
VdXh2Erq7oHnBLa9WR9GmbnVWlVHS76kNKSJ28uu8uxYiVIXa+BVMCGJQQDaBLPvWQmNRR3tOvRM
Zsl+n6g4YOLq0pnxFQGryM2uQuZt/7oOHKTJfNvbmtNh7JdOiXnX/ZXkxCFfad1wT1AqA74F7FEX
AdRMWC+lxvfmHSmEelTQl3uUR25aKBfAQjlU8wHgjbBqHT9DhKs1x5kOmBORS/QIA7aRMX8p9wT4
f/u0aeDC9nJGDMp69Z5+DHZHfK8mP7Tpf4eUkyZ/1cobFQ80NCJ6DpdWyGDTm2LhcVR8GxECDUI5
pteLYBlLcqGNBaazj/hB9c7oWemRJ7PeZRBGkOGWSZPqvRhCLY9OjEcOSNhjzE2/UeWVkfbaManE
gBp0OO/BME6BCwwTuWIHdkB1olavVuDVrdWwhpWIO3DewQYvaKVL7GC3v20lHUxDAxU0tsuDQUHh
QvGu0rbfcchDANdzaCKGi0DynSqXtYSGTvESta4Msn2b4O0jgE2GowSs+wSsN5pZLq2XLs+pfGix
WIXoXJjr4T4+YBNTtcOlb6Q5dqJ12JpsQGnVySgT9QslyfRiQiS/MNP9G/rt9b/QNs4eUMsaU3jN
eWC98GdPqALJa7zXEXvklGlol05yqnT705ucL7gS6e8OwJ71h+sM8GHROGXYQ11DdPPHf5Zl+6nR
vvgWAlF6RlB0HJrLgEV92KBpiP9M9YUsWDNZSZl1s8JkaxpDsEH4+nw3VmCipbmvVfatO6+v13JL
pF/X6MJ9MzvywrEMNyXBjjXdAlOMhjidIg7bVinyICHZ2G40A4kJBOIC3h9MMI7dUB6C2CuLN4Lz
dU6X/g4uMHW7b0SfxHFc8Acq6xt6v+yUu6MRGRpL5WtxCFJ/LUIcATPcSGr6h3L7lETHjpwuWc0q
OBo32Mp84UzYXwOQh42jE0Tn7/BN9enXoLnd3CsotWLmZSLxtBStpqY8hmAsXk/XDGLHn56excYf
LaI1Y22A3fcuVW1h0I2GO3SZg5a5IVwaWS7tEH4T2Syglq4+lfqZeAZLsgSoiE+InN8Kh28DaQRy
X+NmWh4kxt3I7Zov4oje+2EpYcPeOFOUDhvx9OFri4bJOSAPLyAmolB8F9Ms2ObAbL/GHCKb+TzK
tGmDwJRQR6bnKm36OJzM6S9g8n3FHGReL5vw0wUBSIQWWxabvnJWzUSFDqWjx2op7LltiMUWeYxO
dkS1aFrl1arLtDA3/DgFAYRG2fWW5p600F/C9n9bXB04jStLplH1ET7O1hWrXLg5pZaLJDOJu/AS
hWLBDLMZeuAW/Qo9qYs0a320qGR5a7VK9QM8QYrfOYbHLG2kGJ3PTtKjQCu+BDoQNEpNjq3rs8Of
CZMESebFx0li3HrDKA8VyikEzC1yoeOJVaqRyBJ/p5wbufdGbqZ233EVhlh+qv6UwiTSuG8ALEQj
Q1j/fMZnuVDzyzGxP/U2RUYnoG27bNLeGczUQBpUk8QHnXHRpQJ4+LKweZ6gvXsm0znW5/iv5IkB
YuvabLZBQsFcZltGpsYlL/am5MieEHK0w4nJ9HZHpOiXxOmq3/4HM26uZBXcJiPfvSf4jcer9EXV
AsIpBqwjudWNjHfgowRNrtAwoU5FOZLUxZDCRp6hY7xFhf2a6VVY8ipUv/OodchCcA/1sUwOIoan
yvf3n1t+wyJo+8MnxxPGywZIL+fX/zyzBobULODNcm66819iswFj3Wm8CVbCGt5WD8lB7O+9Rmt4
Ptvbb1KDTbDwVH/uZBb3nRk+XH2CJUEXQV3fosTLIPFtRaAStEfdkzLrJ32boOjGrXee23wZhvrQ
iI6WiTz4xS/wD23RJTL56Fx86jnRsOHsiEbS4e/xlUD7EWiJVPsWnS6H94j6rzrZ4mtvL+1+HGVA
+a/fQLRgEArQjX73JVCswqbWaJF/2Xf1GCOU+2nSRWvdpGW+GRunTF43rI37oQq2UC63VFnsXU31
F3kv7A+rHpXfyK+ELkyxvwuIIDdxFp1rMKVIgCF/ETVvWVk1l/bR9hUhk3fmWQ0TZuIRMYzFh38y
cqNYKuzgUNzkmb+wWQEr6f+Qu+U/4330FEJwGPOOsJgoAREoSReSxAEPldnn8KN1Ukay152/+EEh
/PlG34qT7UQkYOKppYYIcVjbyn2SmJg0NR9Mfy/MoN5K4mJ3FOVOD8T6wBcHei2LgnZ5r9TES1x4
v2b+7Itnlfx2ICW7Q/QgRZ1u5GMdxpn0SXG3tlOsCV1UdyEEWA2DQq7U//zxs94kuNCtAR7x1eQJ
iL3naEGQaY1TDRAxTV18gBbjNeCL8Zam1I90GMc54izGEmS817pHhReefKoKmSR8CE7iFdPkzY84
vTxTB3zYIUpHG+7z4bRFbMgc6KzH2Hc9JVU4tNvfRZCNQ7K7zXUnmD44G/DJSzFVJTab8F/6eAWy
A3t7fq308vUjsngMV2JgYNlF3tjLZl5sLcWhH92EQ7oIM9JlZhzQgoc5EX81G/X6hHhsJSe8Bn0J
2+enx3AmxLiqyMz6ZcRnacmxPEhhkaRtuIjxncbak761L5ij6rpW+qfDG/l4bInR6ZEXd8aRrs35
RroIgHPLFkMwh6nmeYhVPR61/3bhLG3vSjJFTi0OnCjRe1ndMJN5ihFySrGY6N0hsvu9o8J05kKs
gyo0EncG+GZt3zEd0N72LIl2s8XaRcng3Nco+DKtP+WqU94mksDctgUZOYeRFci2VtxGc6zT/bmo
EweozqMHruXbs17ipavczdycof1glxfiNt1FWkWTiSpGX73lOXupR1IZ5BnbnBCsnmOcsIxKK8OD
0VD5SM2dkR4/iJSmpgG700xvILy0hhlpk2Kp+abAt90sN6eNOXWne1QjIPA23d+ep40SYTAzqPWi
zHO8ZqfuhxZvxP9WxZz03k/Kke83Rns5n0oN7lvR5QmpbD/28xci1hS1Ml7gmIwQ6o2h5Lq92fOp
bgsNqCaFhgW4WPFAQZg2DnzOKpb0rxvnB6hVrOqRwbWEgLG3bGZSC6Rvf41jnekHl2pMU2NEUwOj
y9Ehue/xj+b+4j4SrW2wZ14oQhaq6FWqvOLg6+N7qLIg4rpwbwWCWw4hONtWDX/SbK1JaGNZHeum
XLunfkzrFrYFgjqX532p6aN0Aqek2lcSVc6u9gJdTLz5W1UjrHkZmBRDr0Babzaqp6Kl45HOqoMO
+r1lHlbu71lo6Eeb15PidK+bmZGOCsboFegewBJAgAtuSOoTcUSnBXIsIGQU20hV5ugtiMszDNq6
WHWUaTQrPum8Iw4kQI9wLTo7+Zr/jDIaCl177SDgE3msL5jbIaCI8Kise07AzVnGHbhSr+ts/Cwx
X6R1eDHzXXRWnJyHVR24a2M3uvJZKcpDp1io6BPMtMQjL827w2+Q03p2OEZFla2UgzXCj2oFE9PP
ugreKv7Qqnj/ajTO8fpvWAvbHGxOqIqXW86XwddNcwuF+He0/ExuF12JZ6b7wwlUdcmc/38nO0lc
GnsmPb896acQDvkRP0c9jhXQfbbWwLHFA50xdtEcqLxMGCI/19NspFiV/EXFto6jiU85F0UrCygm
Otk6QEf6cwJA15EojNaFCuIcxJ5+dPi8DztSyiqy1tg2y3ZWJ9mwZitqnh8BBToJRn6dyyiy+q7K
j3Z9yHAEO3jTcyPpe4aqHW/FRVQqXd6Na4HV2le/INURhGR2j3l02Bc960kth5kzii5W6KU5wguN
0VHa7TF7E2iL69KEBzozzwqDyCaH8n+bjwN0TiqgxNFtT91t8VO78ZIxQTWcld/eIjsZGNYS5jr4
v7zFLIdCkntEFRcky7IzW7VuetkUyAcu9Do7Mo7czw+TbqKCu7n0UhHKBJF7rlF6x1IJzsesjC1h
3ZfBM1zYquMyX0Vn5IzrDe3Rp0HX+gMd4jAeLZuRjfI2LfDbiyfvDk0OPAC3fKPoP7FK8PqcinR3
SFNhBupLB602Q27BmVQM9pOeL/soiZA7Cxru2hXDjsT0HCHBMIsSuiGiSG37SXfof4y/PCEUyAZl
AAbxv8h5LoVyH8ijjlv3gcjDcA/HnbAzr94B4x0/fp6PCk99ijzRmmkXHWulJuP2+6JwxzXkTu6c
iYqTN2SdpCJIH3/o1r27ezlVGkXsAQe5iFm3hunbi00gJAQ2y44Dwb6vKRKbkwPSnNgAHj+/wB7K
dP7tGsfCZ1L7g53JaD8vUu6Kgee5X7BIDTgkinpgrWgUiQcjGqcI86Q77VZr5lgArm83+MJhXdWQ
Y6MaPRwYwMggg4DryydoUchRxr7fUumNq/WaJ0bR735/Y10Gvzt9WVcXU0Ow0YbiaKO2jlO7roeb
sxshKJWFLQ4qJ/SFrmFUAkCzq2pl034B7ij/67zSu2rc60cv4R+FSbtAg09IRYCVwQbrPl9kk4SV
TmIOgqij7+bH3SMEe1v/iB1qyGxVmXMSk8wbcc5KUacwzG2n/0Wg+VVhmWJq6eUBlz7d8+rn238K
1zml/qFeVE+L3Iw+LYbYoWZxcbEGzd5OfwIuSm3hpU07mFpFPmKTNTp32H2b/1AmAanYhNuI1s5t
l1Y305zie/qQfbgY51nHkWV0B2n5VYDAnuHIFYW13jPD+EVlzYLrMQP3m5hf6gRcYK6tTtMxMwg+
BlER00gock7PtzdR8IEjkUZvHV8+ArcQNiE4sDYGZhjmQlz658RpsKMd3xYLre9wfQybAieXtxvK
LymSeIZNsqCrGtX3dQS0FmgrKtLL0qINbhok2L2d561z04VUGDg3S7m0ldztBM0C2tUle72f9Ncs
JGia7nrBSJa7DZQqZI0VShtX6wHc9ot8g1IxjY+/75xvR91zXqrB6iMKzhGyVLS+Sfiij8R6EqHc
eRILj7ceXbTHTThIez+gplHCshMaOzpe5UrDbABGbCDalAFNctUzHhjfh6cBezSWTvU+wvunYdOP
UhsxTUw/rUWNmLE3ZO1IxE9SJJmwNG0kTz9KnwBFhu+ls/6iyMz/ThbHTP4rvAt5AIJHjjBL66i4
PM2fXKi3TXVfnH7MF9HAgDcbd5gGE806DphkTe7FFFz07PUYPhDmdEQnwpnhGze32+8rh9ZXOd0V
wULsLm33bufcuPs7/6tv2fTTPWiTwxUjB684M0K9XT/uHTiMBfAYqe9ia46cPSghmlobSgaB13I3
+kVFtIHwCRCBCSe10vfVKDDrvraYoqLYX1mXR8IzkxEMoPEw8ReucKRbI0gaGCbsuviQONM6ijtU
gK8YvEDA9TiA+dPgR0dq/+rIGHuKn2RTvYt0tYoRC/vRXkz8Dh/s+WDLTuKDt+ldTrltrQT2Bael
0Ll0FkmxvxhdQN9W76c6woD3gWL5u8HgdRDpeZwA6FXChmVsb5iFTDM5wvx+Qb3CXP7X8N7feF+L
tFmSAq5u74WOrUy1x0Ry2gfKpZ9+qlB9eE68ghYX3EybA6HU+AMr2xoZ8HbloZqqoYw8AxF2JZoq
BHKu/aD9Y7bnP4LpyPS9vclfQxKyjgHDBg7bn25ywTcp5Jg6UfpRMGTEGlJbekukhTYSPivrv3+V
IxWrAsVNpkfyTrkS8wnRdI8+jCaxCHGAG/VWNm0jDrU4wL3duTWDMy3Q+5Sriyu1DvGOrSKwCR1/
s2zuIxbo/pc+jnBrTh+V0t3j7z3bcMdRzdpY8lLJrlnYeBbI7IxeWfNnF/z9f2Sg40VfLskgx/RT
itn19cC6h6vpR0OXZ3ZJEm1tzhoAfogXHqp6eLclrp+gshnMxyGIvCvviBnmVucBARFvtLlBvVki
k6JlwxEuZRjrqzOVNQA05/RwXr8XeGsfCHTNzkove+s7O4Yl+Vp26jvFApV9JCbAEIFWCsrkvXFS
4REKzzjFBoJ47momVd2v552hlZ+r35cHxvCmDH/3VKELCkaHJy9pt11VgZSKnIIvRv1EA1aFPsB3
dZRmIfduoCnBs+JflLuCdWn9rgxX4qjyRq//tZoCMnPMsgSiEjLSCBcigHIa4s2MKJfxSYLwPA8Y
nEyQgptHD/eoeNb4eacNUCuJ3rjxQ2rgQtDcmb4pJeJx8mOhwC/dOYONeTws9Iywdzy46qXokXgF
YFR/JTXjAtG5vAocGxv9/dbEUsXxfSvhYCdUlrHXxujV2SFt+FWjNCmHep1QipuOSySMuejFMeB9
JwbMJi555tv28Frjy1jc2g9sEoR1YDFszvYBG40JM9B9lBiWOZrgZI208rkqrfZDrft5K+ziqkPt
+k59gX7C8oKLIpDX2v4K7oxqqkVyZUxh2o/Sx4RGNVnryUJgUEpUgMoVP+WR3SAb5f0Ec2YhNNvA
Y9+4DQS/jalNXTlHds/PUti8MzWsaQ/hGKNiv8dNL5lO4SEefY7OAUPX3XjRfOzDLMRcSYW2v/SZ
3LPBk1vVy5mxlv7hETK1BM1ccUVwH0eY5BxC8HuCJ1BGdl9m9WTb6KOJXfI+9KkuloZtjZmyzmyz
0dfQsYsfCaSELCF7Bhn3z+oeESlIwYhP5AmacSNQIi4hBNH0YaEtUBETMEdTQuX4EnY2797E9r/A
e4q+GQeRpJRBCtZy0XAgmx01a1r733pPFnNhYX6R5+xcD89XoRqeC2lClZTO0CTKUvae1X6XDs2j
s68Qe/p0ubKsEAYfAJEjrTf8Y+BSZAN2cNTl1UzQfIDEjOEh1C+8UAFwJfmX71I2epT1UekxiXM1
ieLIpbWFFGmJPdnX4cAeRvYygdiPY08rphcGH0WM3wQ7Li9T11dJXAEcNmX9rKGToHH1Psu/lFhJ
wa89yy7Tv7UQ1MOj6wR/CFiy5lGneRO1w7OL3ZDB8RfXkWhfwhdZ7g1GVzo5aY2OY3UjzH7GHL+U
8kh6UWL7UiqYlWTTBJ7QmpS4bxXh7fbRM6G8EKAlnvcziOZPBBODhexqoJ8/5uS4h7XV9xgiNCrC
4H/1hdc2v9GLOj2dLDwXNQFhL+ru3wLSDINuKadeN2T0amBE1Lmdl4Zsop7H2QQMh45JTKEYrioT
mOszFpq1VXGpzJBvbB8p9HE3vjpF4b0U1e5XPk7zliCYe/pC+x0phwgvdCLcEAEuH8VRCGU3rfKK
7JvtbfUxmNdLhS+OiDuzHi8dTicu5ceLb0nNF0ndP3bIV70RnX4nWkdIFiumCM8oFEw8rUcCRky6
m69XYebfolgXgMBUHltJ5Zr5BD5SXTZr5LbtPGxnhmD0XBySISUFHXd1uzqyV/yKuOEa6PABJzZm
f+8aHidid8oSrkZ13tU7TfehEcTGWEsWRLhSQc+odTOBxKNiArdixfpnGjOojJl+UchuFI05k8n1
DGZmSJnCjBs1bZEPFbnE86g/GFgaKTfH5Q0a1AE6+4tabTQJfhblOBFjk5O5gOLHRM6CNAw8fMHG
eIcuOF1sPVDQJ+ujeBuYg93esrc0KE6n1f4cY9htr2CQlrHCzpnrajpI+8KRi+nmBMW30Y7j5Kfh
YWXlcRqxedts3Q00qdK9z2zpeRDJuQaTvLse/1eYnWhXgkjc6ewbxcQZTZYU7x88eby7we4ashe8
OOOgTbS2CWwuHFdL3EatcYDgjH4aE0gKBM4629Jfdvu9oNMyJZHTAZ/DYeSAEPD02JgLrHUIF32A
+slaTYUz8u/r6p4Jo8iwj/ceAtYtNOewdsXHT4z6dSu/AEG+MbX3RVGkTtrvLgTNl3xq7vh/La5G
mTZv3SrbKbrah4cEcSoQeHY/6IVZTILPflz9cy558OvWEWz3EWJZN199pcQUV5UK+TfxkJ9c7i48
EglxipnmTaTHePUWKEvWKMOOjVsU5h7d0n85QU4eNVfEt/Q/HvLU1Cm0BXmWmV3x7X6Lq6PsCUfa
lIEc3tCaSMqesPdy0PZeBORZKMfK6l1cqdZicYUXVruysk25+mWCpOxvXEMQlSGvmz22t2xn34cV
TjiASEAHJGLtfTFCfTVkUy924nWXHydf5zZDxuBtyV6AwrPeOp1eHEOPB4aV8SR+vogXXLhC5FfG
41PNlWVgzxoYrhY6uJ+KVqpvg+uLuKM6CDZ70z2kJtXBojTL0rwKhUbny6j4BOOojt7F8RV7ozNR
rnd2RTXwsK6XI7cKhtzGqW7PFSJrjKLF07WHBqdT8VwaegMhF+We2to1hUlSNdoFnUBvLJ/JODJ/
6Uc3/ZIXQ6UslqUFqOA3TAxpsARh5I4RzB10Q5WxiUDacTlkzLso+xLrFz6geFKAELDTGY+bMFO3
feygM4kYiHySkYbCMfiSwHYy66nn8gvY1S8T6bOupT+wFSJUrkHQCkl27xktL9Pe6Zo3YZaGUVyc
MI9LlK+h2y5hmVbBgTQiU7pnB0MXt2i/L7SopivoNAZt+OmM2RjAETBOjGiv0s5aSsNc+4dwZm/J
RWMMCNOKA2L6rNYjh3wQFJ/iQ0NlfTeTYNkDFlUGsNJK8G3GMmpvS3FPG1Jy5QAiLFgV2O1AMv41
h0dHj6ADO99M4WDlSbzD3gr4uzK5Nkny5DuA4es2xBZSylzro6JKTwF8smQ1HtoHCJxL3zQv2Zx9
aEYjWIVidyGmLAuM3jMX3Z4uTv7fkS6eq4CZiSJaAtctwKjvP86gQ4cR2vXAgU1uhRwyRuxEMfKq
lbOQSpT4KpwqG5pyjHTFMTEvTbnsVh3xFBd2/bhYoQpG4JWfT/qXtm+8JOPMBiNAMMPj0rKP5mYX
aFIpgWhRNRgenktZAxGkc0ju2JIyDyu0JCP5IqccBbDoNOmWPoQBEwBn2Ihr2MEk7fbqPIzaDcr3
IABr3iH8OIOyqQaKeDaha/RlFOE2SVh8YJN7CbiBLB6ixVVQ5ws2UMMUB+7BhV0M7J/uvQ1hQs8p
j0a7zbgPKWFmClORxEmLu68Juovksz44zS7/qD1ALGR4NiVeohnUeTiHa8aKRMY5p40lpaTFZbP/
yXZDVHHoqiqZgtPdPBorXSwiOv2rZ890bBN2lGvmKEAJE3yLX12ZMeG2NcEIorU7p7L3ZCQ4iZPn
3LRroZEH54ay3upYiKqSl2WYUMbwE652U9BpCZthC/blFBiO12RFLuf9J3jSHSnCw2HPrL+P4nfA
D1LIxbWembV8ozITpbyJ8dZTf+KlvO31LrHdUGpGP8ubMkEDwQM/uneOWeU5hq8Zy4j8ZI0+sNbZ
vIU/oCGlCSvP7bGvzbC4vMD6ch3qPOQULVVVosaT+Wbxa0Xi/HJUTIyXEtIM9+88DNKTSmctT90P
xu+FR5hCN9fxL6ScwbIYruLB5U5Bf06JGrCXLsom/ujLswf/bCz7q5Pi3jM0/jTz6biZ2NTdE/Xa
tyjqRntpr4weM+3r/W3YndYwKXeZsLRo8LCiG+m3srmMBsHP590GdvPqxeW64CnXzd0aP1D44C+m
emyvVKMJh9BDU8v6hv7ycTRcTqjqIp6c7XU/4dN++cljW1QCjiGdRZ9VXYcW06UGOV4kom+HNeZR
lxEY8qV1QUcczd6f/WS/8AF+MbMYFTqtcGaXTDpWK2fMFBiXjH0XegsNIYZaOxsqGqgus+P5Mkcw
so5wXJV4aa2yNCa2aA2uTr7pW9dXc7IDRydI02hn4ildqFiCvwn4v2cV9o/qqmHor09cRCYX08yv
G1S9XEWPYgdsJOatBetfcItVbiooI+ohrEb4dKlvN4o+jvsivgwl5jtfeXsYt/U5hrV/9f8bhV0u
sdCN8qfpjLB7pOle8LvOQ5zZX7IfcZD9xl4ob8UYbdQwdIjbtWmTTv5Qp/4dDmWFNlESFr1WCOp2
KHaTB9Qrly9EgHKr5T8BnVqu/3dzfXYE2XQDBrcPvXm1YjldA0aD4tEbPbMyJsGWARWiM04KaOwX
Tk3FilpsL5+10u+gchuBaQR7dAQmiqJsvo19llNGnITPvfmACVwWuOjVogH3SgsTKvxs3SILbTrx
hAe1LTe/Z/1D48lE8+4SLDo98/IgnnMGvpv2uuX380+CiVIvtMk5jgLV3SOx9E5p4UbpTVl/3tR/
h1kM81V/nmkRepVuM+ARvXgNoaHjHHBFVtwc4FhpH4uyUwmoE7HNuzYwOWriyH7PUFN5CxpQgmwx
mf1bkG82VFsuUA0CMurasLH9zgrmozTlwoU9OwRo5CvbvnReHADo0nINDtfUFzVQSoU1GQEcdp+M
7Cj12xqaQeyRwafaWpsONYeCHHrn8aAj3gXlLRbWSxd2oyDjjSTXoDRkLxkIukBKpZFJRxZiqaWU
xm+w/NjQ0BDVpgZdSXNwbFUMHg/jyWUgTEeSFPAzRV8dKelqTNp5CMp0TAB0r58skjq1ApOeqL9V
UsSo5l/b2ieGgQjfHeVKuaHdIbJ7W16jsaeN/EmQFKypss2TbpBwuCJBQGm1MneP5QgQOeph6I0B
5mRNt18AwfGdMzx27oGtOx03ETXjZthICGGhCq2DiyhRDXkkUyzRRhkYwF3yxcFytatT/FJf6crE
dnH42eNFCVxtn29QxbeJUCzyh3HFDU8zY4J3Ttyg340oWuMo+pZ/mcqRrjZZWItuUxDzquIcngd4
dxCzJYhcLtKwwZf5HBEXiJX25ldHn8UEBMBv4zfX5DYZ9v9dO/LmLrdJk/NRQv4KQbG5NejGDzuH
gHFcnZpcPoW2c9vnTFMIIS4YR2t/BRDXzmKvT4XTliJtHDjw8eZCb1uU6dyttzjAO4iXZERsRQ3/
lJY17hmo2gLMqYD3X/67GlgAAAPMVAmOo/KTj98VVUgEUeBSE1+nmbqhIFEO7iy+GjcGuQ06/+dp
P1Opj5YTpS/FU0yeqPdOjy+73lfZJ6Ce7EB4IPJFIlVy6AXIerX1IlcqzBM8RayKHxN4iN+Q/vr1
XfY2ogp9bB7cKxPw7qrPWbbmVNUpCGyr94GhdQ2kF1zil6M4mkmzRG897XPVLUkL6zTlXmMOQaoD
eCDq9fnOPEmbabcAARtJ/sL5qBI0zVOM49t1sycpZVaZy8BJjHEEANnu0tpOoxYgf2j4asEQE4Hz
fXH2ajUkpogYnPj7HNuUHphXL4RINhhepI3aUSaSxdVCdyWUgbk3NFh/0c/i2xOpkkPOo9+q2ArY
yizrTRopDYq2pC2GrfRYrz99A951gjPpnNdy0IcEXoEhKmYgdBNnwDTkq+SjC7y2D+fI8l0tBLFw
6877iRgIq4yx3uy6PjN7awIgf6lBsGEj6mACjRlrEgA5OymcokupKQ6hnZsMIy1K+OAcKo1fN22s
4TSggSg/aE7k8/NeR7VH7Uj5iTi5Kpb4cKZn+Bs2YeQ0gXAOyrOuTjA8FiNBfTRu2Nh1/8hj+RoP
hGojAsni2GHxxcTAlyRIyTxMBO89rt5njXR+pPn+h5DjbYrPByOen2pKUO/iBmCTviLrnkRwLFen
/m/1JSojrO6YZat9pDuSiNal9zSXk9ImEd2DP2VH3Ee/eaO4iuAw590HFFD5NJrvpJrra+mBoWBy
KjRNgs6HX8wfrFRBMwU1JbEFrJX+V7ENStG7gYZ7m2PvFOzKPFob0OelQKATPf1W59UJxW8jng0y
Hw+RbHkbAPqezGY3RrRHbJjXWXoT6loenZflsX3iBm/e1U3eNyKKdI1YKrf4QtxtnfCeZe1RbEIo
UksMiAmKAMk+J2ASFL5PkSOeuYGo6PPCsMhd2bJEK8uJi16q6BJcj0J7Kg4w5UB3GNmNOGHdFR0M
b0xj2RaJUB6VWMI35F6llRZFm0zOUBcVeACP1v401BKcVsodzNNE3PnVsOc86uS7/QgyHhzv374H
VvWjVRn/6Pz9DZ1xllGLYyyYnrKFhmyelnpLf7TFq6O15rvGxV79MGlu9XOlJI4KJwqp2zcR2wN7
FdczeQnhUrK83KGbaKj2ChEFRLbfkeYXyuco0HpN27EZJf3oFnqOt1CvslAWxUfecbgR0z3jGFFz
hJwsEBtp/n2FeXcZal6/mwT/bEgWa78LNdTgO9qj9tusWWNoQIuRmVGGk7mHPO1FZ4xSDml9OE3L
3lvCnF49Agvb3reRf+8zCfeaj20Tnvegm958wa+4SCV4Aa/nCzFQMsCYskOyrZdlN1kJnW+Opm0Y
ltlWLEs23fjHvuYEsQ6uEGimb8U3/3bxC5UKDVFxh8/4MMYym2k0c6VGcRL9rNrse8Ap48A0+VC5
TjaAmCARhJ7AAJE3qb9TBe3IKVA7EJ7ohtyIDvbNRkOw7OFI2UvOzPoY+Bf+4PND05ZbzomjinjX
9kMpP5z+L5JN+7wxs+FzcjxX1kTtQrAOqSUDENx9F0qVKWLQ5cWIzLGKTGrKw1nOMoUPc5+IyJn1
ByeNN4er90WikF/vTTL+ulxXMDPcR10duwtyBcutGVIaGaIc8LVaAmD7X/vSsJRdbfjIfRJSK8uN
8Z0Z1EFanNd7v2L+F8eAGxM+SbHwPTJ49AiFXeMDs5cNoA4UmE/etRWATfD9fnxFqdvXzx5LzPX2
wtgLbpobEL1ljbKXlWcMgg6TpUP7nZSWBlf9iNaK4veJZHfyL0zAowYviPP9bhlHrwxu008qe2yf
D/9pGH46tR66t5RaIAuSHcAzpe+VapNWzeeqegxSK2bu/p1fDQ13Vfc24VH8hsC0jbMTnoPzwZYD
+Ikc3kxRMkpmbbQeH8jCWEqccbvD2PSpcSjOc+dum/IwjxTOO5FlGpZ80zKGvcdrcV5FWHOgn+fO
CuCooAJGmI50wIuhadxgaCCmTIUz3JhGEYkG6n9XXhmqZM/QEPgwKyfUpGkQpGnN9EtV7swH9ha8
aLCimdzv0YS1M6iRwMQiRCrVHcErl9Zaw1Q3i6HFR7UPWk/hfvOBlltUJesixVm/OkdTRcKXdN6k
YwVSTdICZyXcJz93YniofdgyC5AZmFtfmwPOQMfKFRFG0pX6FfvKKANbjyPebZmAoD6eNDEqT+JI
7b9pWYVujIGtP6oSoVBSR/CcGP5zZw9LEfulx987rLJIIODXJjVJnBmEkSIOxol9zbhx7X8aXK81
+iokePwUEeuvngpvo/kuBrCA37rBOuUbuK1DTqyaNSyXf6a2mgUJ3iVVs1faeMxDOh5gLKxysENX
iJJ0OYyFJ2tjJgqJvzCXqUcDaygsl7kqWENebm2thzXbXSSnnND44+OXsnZUH4rcJggfFHCE1VDg
pJM7Py98kq0LkNmU/HJvT1TpaXa2UEmR4x4HXroIz46P5cN8maNNY/RsyEJkE7Nf231Os1zAk6Xz
mxPxwk7ZDkTCBCB7pTWsbxgWFRq+pboswj4TqACp8xOh3CqRAmgZ7EmScBP9GeU2aU1Y9OcciEvj
ka8tepp0Nwdwhcclat3Nx9DUULSCKzLLVun/VI3RnFxA8nZ+rlKf8zaRgpzXiSJPruXJi46Gmnhq
hTwKw70wpc72EsiM1Bg9FCp6poaMnvoIAw7jxmu484RjoztphyyJVgyfH7aV+dq2/DH1QGz8Ndqu
F2m0G9jLmOXfO7gqi/fjxMdoQynO4Ugq4ER9ESYwUQTitY/7odiHU3vnmhOFHP2rHpEmGpJQ86VX
hhRz3GZQmVWtwuEVC5F0KcjCf6M/3cDmlHkl+DhQEgvJ6gt0hA7qBix7037zgxJvmHLpOC2kuOsH
kiplxjj0PORR8PNRfqGWKDIaJziSPZmvwcLbXwgzMELbI8OkC1vq0b98DnrWotuLw8Rf5v23pTlX
82Pz5BUxvXdOkgGGEY6k/Roz/FvYqUaoodzTQinESPi7sVk1d/gqb18/fshwCifgp5+4NR2UcfCK
jzzEBL7efTCBahIG08mDhCIl9o4UiHbB3FpFinMHFAobJfktbYJJRzPpY8N6RbrlpEUT/wYrftmu
mr4/KatCogCeavzo0sLgBS8Gk4yGAILpT57TVyYzZpmaiBrFc0fyJX3gcBEbWOvGJn8jAYHsOHjB
25be3aQUV3SzciQnLn0BQWmnc54dNfUQW7vdXecc/D22MmPBzPAAf0XqMdGHLRcQwnfmdl4gS8DP
i6zMpa14pApkA8a48/3LGezH5LEizeHJRAgm6EUYCDunMzTHk333RCp7knB7RKa8oMIMVdTZs1N0
m0PIwayQosQav0bgLTrzrh0x6Fi3/EFW00pUVMMJ78Rq6hmllM6UOSpTC2OGNgwa12dUF0dgKjtk
tgIquWrShkRY/OXfq3268YgNHj9gk0T1maUO2PP00HDQH3UrKECkBKPPeETlLRiQy142BSKHJqgo
z+iVXoFVKUeGug97HVVG7W56js3nxoRxBW/hETgfPJLkYkHQXrs0lhPbOt959y2CdoGglYa32cuN
kt2rtcact/xIeExEgoKSqIfTcaOMRyMdsKjRL0bqrrNKn3S0TDoNAtyeBqOH5hVwstdoXkIkYVTC
EpWcAvaum79kisDAbXTR5WRKjyaCxVvgizSggZ4VvDU3L3/6lS1Ht8NV4x2dHHDRzMlMXC2iuiJG
WEFtZ6kySjigY6nbrp9/6Ohq2/uhefKj6iIdC7U/H35DII9qjwU2sEjr3U8dcruOMX3/XBvUKuXY
JjuTd6sPtef+gB28WkAdbJ79D9V+kYZbnEzgOSXsyafkCKmsbAC9OyK4+NgO0mtKfKrP1j/4exTj
hbGLBvTNFRI2l8gtpcd/5Yaoqz1Ir8nb5RwIHsnR4M3z5ilLmnoxx6EItIBZSLaNq7ySYUYHyNHy
7L36Uz2hXUWYn54jnNe1pV/BS1oFptFVXQvowjc/0F8hPzdXx8eJZbxOJczgTFaNtcRcv6+b523r
ESVfmWVHC0/FlsLZju+9DBCuPuXaYnYD0yOFBigeMlKRn7oRSmUVQirVhH5xKk9owdTvfdRbPUfl
kGeERlaGQRaSAnxNXKlo2UpgbKYWpgUTJv3acOndgmR5lrYReX0VGBNJA+rISD0eZs5SB1bSmeLt
hxDLt3AJZtUczT4y+56FvrE/D4gyln7C89LSYR326MlUWzRJnujB0yMUuGKtvF2vbE83OH+9P6D7
oQdK5onQZ5D6K0TOB9p4JnQcQGXlDLe5zF4zVmKdD3wjDHi5mO6j9kodszKccSg0peZRf5SOIzMA
mTmOpYhLJBHed67ulFl3LBHqgWYxDQTcwls6BUt8S3xgsdF9iIa7dvlpmBXP1v4LEN/WPiLUon/F
kBGGhOj99ld8egXPPG012iVnm49zduyZeW6RxWjqiIywDiDn+ZMdQ7qX08q/elj3YLIAUXuVrNqR
+rjQnxnGPJ0bAabHGC3uBB++wBHwdrJFLujAG4idsxQkLUOMpLGqxXAAn5GnIVKQN5irHDTE/nPu
ULG5QF37j8KfNR8xT7LSbOcbg/u+GwcP5Tl9Ea5y38u+wox12xnT6F+oDka5fExdr9VcNun4N97k
HS7EkdXXb9Y5968Di0z9tXErogF8TDk+a2CI+VgI0V+pJPkg8pxhKJJr+5ufYCdNY/Wff0+jCDPT
Zs3I4+ydMs5PGaa/WPEUVrYGPIpmDy6i+65sAlX7QRausGjDIxhl41XIdVFXhMNDqUm+qF75hjS6
AeaQeDhcnKz0q6ut1Xo39F/w0Na+dL8EsSTY/5TY7Xh1GaUzKirb2JKOX6j/RKVtpEROr0miYDO8
CvIJxjT4XwmcTKMcJIrFcZVKnscGi+Law/Cfy770OAsShxInVrpQTiGFUHqt3cHWXsdvIZLLhZkf
2uRw067NRnfNMygRgVLxjWLKq0o6Z1q9a3A+v8cDCaGGtMa2k0H7xysjSADzjnfp8zGuD/8uyXcK
cwzo+9cisoL8T/VD1r5iu9rKTOkxOkKkpgxvu1xtZ/Vyd28I8AZuMwKSwGP5zEq5+918/c+mdvZR
8cF1VWGxhJ7h3T6n036BWMrCZ9T9V7TYnKFGBTydJ5poRlQvwkf++aosX3j6ZdL1Amlwb1VY2stm
nQAqK6FFUVlVxsYH6TwW3G+Oh4+XVrz0UOCYL58wrTQua6dwNrRr/l1WbcsJZAR5Qdtfdx2BISzd
ERBmkIg3i3pnrbkH0MeFiXnXaZGhnXtqBSKg+VZinBdDLYD4DI2CQtqNOUrsZLZGX/323oYWOCCO
R25jI4hqLsrFbfm/AL+agk/MxTKIR2hM4sxjeq8ui4qWWrpxEqATu/lTjN8WbmvMY2i5Qz32JOsx
Hdmn/LsacbY74LvdwWYXPu39tbZ3QM14a6kax8osuw+YROmLYVsF1OvaDJ7TNZxfpKnFW/SoO9sl
IFbQ1wztX0a1Hm4ObKhBEmU8fHcA0qclXPsl+hpCGgty8TdKCZCFB8+aLLv/RrI9h3WF70Oiii18
wNr/QlC0oa1zeYz5XT5gaJ11aEjgQ3aA4Faww3RG6ZUyM54aembudyD5pB95YFfMfDRRjcgeNMlE
LeacQReNyIiJPXvM9U5cpUVSVr1Rc/wueGkHbDw2kBfiHfxrGoubcW52bnz710iR4xgs8vczlyVO
CrLmKHqjoycRA7KAd/7VpvneX5GPOA5mtv2ZMAcJ0258HU7sq/MLmFkyYVTUiE3RonrLgJEtnP41
5iAVIMLFjhRDTJuNUS9524vKt+ZOxJS640r+23WwXfLX1vgeRCKG1K4CIQPS+MRjWVoa+N9/BpJA
aBI8yJPVPZgaPpZsozLX7zl8P4VVbWSBd05tuLg50KTmkLaPm6JFiSjVPbwKFAqrMv3/izmWZKNG
DwY9bwQY0GOFdCoEWu4JRXMGOE3VvCo6asfFHBMyWu6HgkRwe2qdeOGAsFhomIlPtf7NDq+0heoP
DWqjww4EcwNzr2UrR8xSI6yxXg4VeZB0CkUiw6DomNwnXkBVsS5sV956WA05VdJtATvzQ84pZ7xc
K2Cne0pepqBUoF+IPG08+GKGqwyOZr70oes5ncM25cbtdZ2qPHSWXEd6Pw2QFmuDUC56JrQ7JrfS
2qfNJsI7IyVTQ+5XxHkasLIRWkzXTBdsGDXfZF2dV+VqkmHLRiBwic5IgSz55PQWS1g38ne2tGb1
6rUa0s6yOfRfAHzXxyjPT1s5seRlx2Pz1ak/uXkWpba1terwZvO76MAcxtLCDi1f9bFk1JqXhDPr
x6Nhfx5/YvsHURKDoIlslBeh2vOt5uDdfupfhZxFNK36ptevlcpWA5QOnzDc+kQrYNmv7PwYu1KK
w7UWPjMNuUVXEnXPUGbyaeKPk6cc19YM+Akef7K3bIedekWxG1Nde1tJL+IgrO4oSTgz6Su/jomF
tfcqaw5TCbrlE/V80BvuRjQXf9Z9yNDN8xT0WVyaNTzghpmQf7nrBompddQoser692ZQ9dtgBuor
KrQtvBeatOLsAC1L5eL31cRdh2DYYAD0xGsXSlMURbpLiGnEpjFr7KON61ohS13g4yVBH+RvUEsz
ye/w2RYagJoe/ikxqO93e8fiVXSuK2eVRuOPa0+AuQxG7dVZlthH1FvtblD3eThFVNAvEzm9gWN9
LLYUT/wsVUJ8ubHV3IaVXvlsZOjd6lzbA7Grg+3mD3hY9lLu1cb/9sgEWEAQs6FoxBZak89O05st
TZNnY5djtdMYythmJYSBn8+4Rp+zYadVb4pOixi2PJpsfDpLZp3y5hUKJ3QtSnGYLKL+J95udAOY
HTA1n85HCHKJn1KprbBNDnW/mSWN3DV2gnjicMDpN/ZRGcDjOXnebyvaek2G6e7pDE36tFaBOL+h
Jzu/a9g3RNz9XhslJlbDL8HtKu7MRwdwa11oRWMzHS0Y2Nli/DvQaq862HvENoC2SAP86Zw7PfXC
alM80tsoXzOpcycXqWw/Z5ogkduAJaOvXr3nzjpKLn0E7g2qRQb+4mUTA4WloIFcUOBOiR5ceODf
VAn2aayAjejX0eNZEyafMGyv6h1Lp4m0TKI4SU1o7+uvu5HWXQIZZPaMdAw5xym6xNuBMgiIAqgE
peNtGT+LhzF2j3yNvFObfWtiaR9O/yy2rsclZC7jCz9vbPPpa2molQ9ykjMovrxNlDDtX40YPIDx
XYwR6nsEIqNzoQpUkgVUHfiUzNQS6z7ZNrmxsn9safNpb4YxrunINcPyOCYZiGkQt+xMByIHZxwI
ZErwPR8h7KHsvMiVHEolp2jC7frqRUCXRkOS/fDREyB13/HF8mYSsUT1B3luzGxCwfi51zR6Fc8J
2SVw9z8tMR5Xdf+UMUPUzm1RUEQN1dpZRI1+nP1hp0KFiVyXDNT/YYbWOfUM5o4AeuIp9/2y8gux
s4XRWz3gsKJpOa7iPfYPAMNtiOqP/9qZ/Y7UQc2BvlHl0+qdDolknITCfKYOlBNWvGwtYbT9BuVn
zrxSzwhj/SSmbWHn/FCRCphjeeURLx58w8/B15UBGspo2IdcQ1ctiz06y3kePp7+k4VgBl0QzSAm
270NBaOoFbHllS7++jrIBw9pz8GjUL63lvKuhfMe13Nlmmq3g7PRJAughF+ed2y0Pobugs2y/u08
gti5F5sFlAKWen3bNkRWIRMUg/d1+S4FqSRqBU9EGanIvSZ7XiNXEckqmtrn5Qwz8OZojIxCsk0D
3+I+Yg62rokxYEgbt87N07OmlMc+BNzeOjuFWTbRB5+K5jjpCFnzUOYGgSJvTGb+eKFmy9JNnM7Y
gOHeNZgM/StgZL4Zaz/UFnzOmbbF/9+QbamlSztimMVvF5yQhR5Uzdz4EGCEWFi6yarX+BsxUrFW
ZrnIhXbLYlgZRvgLQ3mvOEt3fEk2YJP9xEOpOkEy8Ovq1uXFdo4XkqlyMqlgVG0sxSEf9U5wxuh7
er2D3KawcZh+F08DFhr5QtabjmFOL4ALVMuNqLncvZ88P1spp2ZFnJdafDgjmDrvx7XOZKjQqUVq
yPTVKHlNzkaRAuFfOGUXKYr6RmvAFuZOW4d6KG3TKvKf4ZpbKR6MTJkanNdh1pyl7zs75bb68F49
pkelN0f/xURLVG5/yLGGshJ89C2n5w4iZLSI3xLvvVzlB+xPV6QFww5vejSnyFJY8z8ZQN2gps6G
Pa1JG/Q3CsmDJhbWwQQ01IsgpiRRP8Hwa7vH8HDm8VJgd84F1GhSq+VoNtOnYP5JRsWsyRleuX2q
FSARKTJa1OC0szJ5kPypvsu0PeoprlLEXTwgGuc7KWPu+QYqT04vMINSwgcBa77xXg5LswRhgftk
RObR+82LDECC6RkWBPPjtCJuea1frG1yWlZOqrtTsf2PDcKshTeo19OELSUrj3GKnwLsBSbcLjUi
XZWzjTm77Z62L2X3BotGOEZ7xrKlcM14Z5krguwBLyjx5KgkgqlR9PJ1qeh00nerwALuurwiOZq0
bZjUxDK5FYF903U/orU6XOysWvhzXpnIvXWHsJFiqhOiXnfXLzUp27NE44k3/HqJWmJVzikthPws
pO13zbHYiR5+pd5MDvgEMDL5XysSMXShDfDpPeA3rJ36XJYG01cEU9vm/J8lpESBJFyy1GhIEdbP
ZFfTm1eRoiVa6SdBaN0PZUy2+LjDqDHaO01uwWMSGGcu4QR4r0Esrx1G9YI7Btlt0lh4yGwgttz/
K8CkCVvKFLrjo87mv24QGK8IG94iD6rUl/gFSmXr81QYNrKJ/ktx7cYfgU7sUmvf7MK4xV7UgRw6
qnK/qY/HPZbG5RImPd+QzW3hQ+wVTL8fEmWibkoa9Lj2JwOodzG50N5bj8w0BXt98rG78Hw78U+L
k/yNkatkDTESAVl2lQFw+Rm82iQHN2hSSb7B8OjQl3UyfE/0IY56rYoGvQp7HeqfsJ3RQ+OWxiuQ
T6QF1CUnkbsE2kD1hF5E6jgrCFsozcDBvURbS5eysf1c0jIxzjQP7UKZbV8YjQEIA2+51jpS3yUl
SXVJqnYzGfCfJMXpBAshOQ0VDmgZ3jwj51ishphovOqnAilIyUIvVEwsLrWOBVbvtZdYUPIrJxBM
n6MMwmD4kplr92E7hWraom3xcbLABBEz/EeE7r8pBewPijFulfTo2XmS5AUtmuE1a+nVuD3SIXz+
OJ8A/a+Y0n405x9/BOffOUZ7XhD7kCmc4uuBY8UEXMkwJo/NV8oX5qJhDe6cSBHAXDaE153w6Fz/
LTpKKY95r+V2HxcudfhcuVf2HB8kVr1gYWMvJ6mdq3sDlW7ASIf/Je3O+AlQ/wUhvXkGHLGPeza0
WgClKP4rjX0Gb5asJrzAyCc+ZZWKPhqJhJK983UC3NMbcUnOXntH5XZg49BGLzrXkYeOURcbQIpI
wvVb4gkEQF9sGQDs61weFymh3n2s+zysbaRiIAzEsDuFBGhlvtPin8XHwXi7JcZynUc9/rufU1cW
wxYZQ0p6w2OT1zVKqg5B9sG5RU8IfrCBOvwzKD1fB2oBCv6y7pc125fR4NPbvc7Uupf/IKpInjPM
TbolhtDdSjyxl3c17oUXMV1PQv/+8JThHEXrpaGBUklgQQZbZAnedl9bxeSFeA9DyafqYzCj17zU
2rQ1I3ZmvVPseBJd+QIUxpun7q8z+umtgXyDEzVOg1JAIPe6MgMfNRblQ2m4/IrAQ4RR3txhCCkP
Na+qMJZlo6Ps8n7pyaqQoQkiDhygLhFyc3t6/MPOvZb07zaKUwNEGG9g6K/gmVQ2FsLcAvwT7ZW2
X5UXvByFr22kBhivC3gICExrrOkLYQh25vVEeVAjl2TlxpiNl3p3haIXigvfHdIiLL5jhij3lpvd
6MwJ/3X/t0AkHRUawWFhRvxx1oZVyZ54e0LXKFAPDlvHpWzVGA1cGXgDp0RbLvRqSnDlf/6Q9LKw
oyj1++NybqoJ/TglhpYLg4FsWJYpW+EPXRTidsc97+mEjsOZ/hFGtoNgtJdLazCS3hgUjHNTtiKs
bVwjLsXnnGly3LJ4b52YgaNZst6aR7igDR87oZS3Fq+mki/d48r3aLflModj1Ehq/1B6q/1mz7+Y
cgDg2b0TW9Dd284QvScmNU82nBc81n1h7FFpIiqugjLxyQLiN/voHFLSuW7btOYNXl14tp6yxD0w
8MtWo3j8m3d2WR97jax2/QRETfsHt9svk4oSv8iqpgEZImTyf75wC2ptj8Bm6BMQILYlPBbBpqsB
lAse0AfV1rJvZBl9vnMqSyKmQCVHiOlRyoEvaeZwVXnJWyVDByyIZJp0gxk32GHbyusDrtscmMks
h1nAPoERGH+Zr0oS2arOHEKmu/4tyiI5bF3uNSXj5gAcJSJVKZBzyI1j3zXSWY1tCpNxeD5tOe39
w/7HBUCsRbVGsCCayg3oBBaSbJ8dDf60jfeTV02boUNeGVg61rrY+3kI7MGxOyikNmsICqMJM9ke
LvuR/TdpXCOz0g9xPJVnozeJNVS7m2ySJXYVpcyWuSmNIpNOeIYvx8P07THe59paJQJdFCdj8vxL
2YM+C1XuMiTH9fAnRI0Uo0qCAYGkCoh046YZjQsfzDE7qcpYYZ8uHWm5kkqT4FLGobR2F56zUa+R
QODSIPPztlZCv/et6Ef2U9boGJxq1bz0OTcWGfuQ5w8mOS4gtPeAfRogBRr8Oj1PIZP9V53IoloP
qmWovgzX/MQSW8rN2PsMSwldRu/tSf/zxn6tAeFL/nMw2vAevd2OM3C6yhUPBvlXyZ2RkLz9jMRN
kfl3YN5O5qBixCsOvNobt6NSgb0eWiesNV5FunoobfgVYbWTfp7oO8EgYDZW7kNNxGXxdpffIB72
wjmZdGD40JAWF3KmVgl7CXgvpIsbYF+XF0GSYxel+4QEDNLu1+sW7cNBaj/4JBjvgAGJZcM3AKJK
xHnh2VngnEZCCeuO6J4d3QB2YZaC49n9smjq8kgWe79q3elmVCB791LGdIFks4AZw+Jpx8j/rrZJ
gTmKYusLJjHQ3SEihSsT92vF5dBlV7T7sjxn9wVQ/FLMSYjUo27skDLeTd7AB9nL8kzquS9Vkhih
4atbsU4nnbcChTqh0d7MKUeq0d8NgrahaaJrRKPt/qOyFVFzhxZA88wHFMS7qziKo5lde3jTOCif
rsz210NYyZxU/MznlLZdJ219CvlVX/XtzlNCmtVl//Avju0lsn/cu8+XiXODOFmFlQM8d2r2edfZ
HPfmjtaivY54YVoe+LqYyqlXcyOQsSSAFSTHVNP/prxNlk8kS1iHirwFErTKJVSQKQGLG+wSea9e
XiE/rWYbY2SDJF9+8cLI+SN7q5zIokdByPm0QllIsw6aGRBjwD+hG07ulMM3/tFvrPzMXqXOj/g0
P/l78IXUe/je1A1aYODoHU3VpPchUwdTF5HKUmnAcJxu5CLoh8Po2BoqlL81mFzEGVf/MAvJv6L4
IEpNLWjZxKsDz9B4NMZHWjixlNGetyxuOWoG3hEzyay3B7A41qDBQsDSrk4xsDRvivv28+t1pcF6
hretr6Q3oYcgKIfwErGXdQSmJW2Fy2Zpx/t7KrA5C7pGPQjYeKM8LACft0DpDLvrtb9uix2L/LsS
fYquBg6GoyytUNh/g2nf8oIND6FRqrf+aRDWJzJZM0rFGTuPfQkOYSb7SCaFg+pqddCWIc9a7j4U
FlA4haYV/c5ZnUirO64S9nZFLntmTGCRlpuPO021hbT7RBIMHWgARZNhhGoe0mH96VrK7UPbZGnd
4A8Me/swlcqVbLrgNh9XRMzj7EbQIe9Sgfj7yAEzvVm7dvGRdTGqQWYJ/342roUHykR+U6LTp67g
dUwv5r1pw82U0hrzuGccvmwsbgMeXw6upcaqsBeyFOkEAs/y+p0gSq5hylvQLvUJLoC3oSWWXXkE
rDNvDLDMXLi3hS+X0VC2QdtUCfbi1FBP3od4sTINHm8EhfQ07dbrGJ2oNAIQuVncDIs2Z/2qy2iI
2PqDb/uZwnrmDRrRwoKhe324P22ofAlZlUoi/5T+Jdt0cD34yp/QtDjfzVkySIEjnMXlUX3zHM11
FukMdHJ+lxZURevDjKVpBySnSwU6kuTzRurtFZgDygpz1TcIebAXVHRuh7EvrUzY0SXC7Irundx4
xg3/BFNKAstHhH9QZHAl07qW+qgcF90cCPiQ53uLyxhQrRA1CVyO+Uv1d2t72FEJKGhCfgyhtmGs
CdTxO6IZoUGe8nIySfWPKkGfsDvYKxk4MyiG6VXlpZdjlP6ein3AzCBwgrsGSUZ76cznkjawJeOU
jEWleqB2fcwu6pCHnwohmv7JJDIKeQR7hWujB+CS3TtTbGDYvvu/L3iXBTS3LVy84tagEehX175r
SBNXTo7W3klSohxOzm8wq80qH3oyU0B+GJPCZxs/+7FbD9fKDUgWzul6KQz9RyCprhiTHDGnZjeQ
0qVXa4Wvb2ObsZCEdLxBlc++7LFxuVePzpYfL5eZUNlw+Ta1Y6ivlBzM5kuoiCqPupE0MBkLZjWi
3Kq/Dk02k9/wOndi6DL1iNWXSg5UB/neYXNZ7CEVdiw7Bo3yRaTAGbYj6Xs2rJUFsd48jTlG/ZzG
nTIdln5KD69TK4b2957tNUHgyZxbnPohn/CToDLj9eZAy8gqeEfZqY6hNtzcDUxuXjHtaIz1c9gr
Kd7vvrBCXFBcJm6TS5V18AkytMPsFDGRvCVDsyVlHia8RArcUVa5/b4jJrCyEA8jQoyLicLvF+hD
MMSOJBjvtCz72lnchXSjWrGeeXahxhqdJVqj08idR80Q/51VyfnkA3mGRiANs5lyyFBxoZkuZlAg
kMYyS75aKlgawG9l3X/ZCUMctfWpFbvkmWPuyqHHYLihIg58QpEq53cEHEyo4JrnByjhVOmnWa7C
19wVIOatYERUVlkeqVZlIqUjdQJlYWOJdzPfgCY4bExDGgibQFkOuiCO8W+AkJZcoo+35/to2uD+
IzWW12EE65W6/VkiE3GIMek5phcIi2VYizs8FdhBnCDyieCWitpUdmIQPjvWPZkBpZ14cg2yOLLP
fP8D5DxcrqooGDFqfCCaaWHveKOOgjAmlHtW0ZV/g3HctOyd7XZ/VjnMifntZIBvuFIAHRAev1Tx
8PJ+1AAydjDAqBBLqWnw5wCWsa7JASiv6zhyyuLgbS8q8BU/5kkNqMRV0Q5Tc9LXk+BfCj2V5KoB
8Vi8RRAnPEIg581nNgcFn1760R41kF6Yf8YJQBFy7tCU8byx4Ri6xuHd617OakUVCvY/ldvYDUsy
7zSmobOmhokIX2yaJDZxS+9moR1PqRA+mVwnm90BqkA3QYEnEgXDp2/KXwsCXnGvmFc6vcD83O+t
PRvW4fq6hTSR0AWW+orfe8UtK+VSvOsfHLQVQCs9jm+WWnNYtWiXNsquLCR56+KAFfiQ2qTOzTSY
0GM8PPTT9ba4maU1Jow1xSV11qcFrhhL/27fg/SbIIDPJEQ2S2hj/IsoFjcUT/DwvzKy/oKxA36R
5kRem0pmH5CEUVLpg2Wo+lrDgx+3tMK1Q08umd3fGKSL7CYnt+jUByJkbODK/mKQ4Ynh0JAZiNtG
+qF8PRhYGgL0c6Vc1d3p066FLkQC/tdD+SmxNdFSBCByOlfY+bvpyriZ2cgTKgrVLfj5mm3gLZvI
czylD75740k6AS5Avm1bePD/wJW15ozTghwzF4jaISnPcxhSLu5LqAiaDw7+AsrXNH0xBs5Wpqxd
h/jzkX/q4uyMVDGfVtL1lSmzMqYJqy4gUs52cxpv1TMMLcNrL3MSIPUJzB2wKI8UVQ3Q2U6piZHI
okMcbYX57Gmm1wL0i7jxvc5r0r5jvk8/Ru62WINrU5IsLWZadGJWRaEr0V6BL0GdHPv08GSaKp5o
2T8wyiiHB0KvDS+Ld75hbkgVsSAewFvNN/pgJis2hvhHanh5ejsUDca2UVWUQoaTGqcJ8hZvC/ne
h/cwykHXgDZ4tslmIcdH1FbePCkADZNV4IbIPejfcdaGe8M6q+PqpGO7L1iCstftoTfWH+jbeMGS
bSPul1x5ghpgI80Y6M4UnJHB4C8ikQGFEtDR5Mn+QnBkgZ75fxGQxJJp3wL0h3RQpLzNq/ONqjto
laOvh3gegg7vkX3FlA+iVCum/mxtSeeoIsH6Gz+HNVuW/m10+q/okrNP8Y1LQubslr6odKAVlWDf
QNpxUawWJJkvOSq2ImjjoKHRZanqwUDdMtmg88zqp5oxbjs5Tj2CaStzhC5uhsyVvTuPPbEHXgB7
lhdm8V89fGVZriBQkbHumyF88htqavmb7ywfAg/x9Qfe5vZS0iiIYIocpC00ucgB6afJUVJ+LEHn
bl3iMYh7IPUfbd/oBAJQ8/t3SPAgFA16MjoKskq1C/xIRAOu49qyBsvCnfQhff8pIR1BoE0obtSn
JJO6QRKiiFQDdwd8eGt6JI2p6WKIN+yfqVCjL9/LRQMSNOz+B4LWoRnVE//QA4xVDaKcUezPfVFN
YrjTpPGpeC0zWNKXt9URNomQsACMz7+nyfRUNqISNRm3DJW16icKvE8+cDk/wAHKct7ufL+DccRK
ToejboFwPPU0z7weyiIm1zdhV6CNdaOdEunNgWGGdYNiJHC1g4LG2xAGK19QpGLDGS0jShyz1pLx
+6y6ljfV8M8qiLk4XvLW3tl3FOckUVLOJwWQJFtb9i8+XzI1lH5XvQEXHbL4+Kxaf2BYcDOslnGS
9K/iQ/oNKs8M8lFlwg8m17xk9p8aIcx9XpTZSukzY5QL2U/vmYwFC+6BvSWMhK5/D7lr50ofW+77
VHqqoiz5PSgpghnehT9uybw7zfLp4Z4khDgM9pPK93SjWdjOt+/W4ZCuwIC5tU2rgtSxU453bqU8
+werXclI1MWsI/SUFDveKh2cAJTcZT6+rrmaKJAPBqIChw+G1qD3C8Njv/rnSoS/I6pzI4seCCod
6VWuFM3gnESgSYP5e2nVqYdIW8nyH/e0GLKU3kDeV2lvlb6/erfvCzYipZ7B/dh2Q2JEU5bU6mB8
XX8TJNUCkKpk1ftcjwUFENkTFZPY0qIQ7Akoa6alDxy0SoID/WOeLJRHQjINu41HGOdHfb585DXS
kyZfZ2DFkMP27Z15wQOwOVo0XQQMcv+hGx4DTMZZygKwXkkEZGKdaMZi4uabeQGjAX8dnEk5eH9q
5SGl2grp/cL+u/HYUSgJy0+NlfiI8DHsl7OTlfklCQPFXrBrEWEPK8QBpLmFH5+49k7spkel5XbK
2t4k0vZPH+dy/CMv3rQXEq6c0Sz9RGrEXZ+MPDt2ZzQTVgQr5Zc/kIMY/pGlwx1AY/Sv6ZeBi+Oz
BRNIOPjknaImndDaSCWNbWey2+ocgHVctHlBFjsnX5t5Zto195Is5F30DYI/c+oImcuO6WAYBtP2
+qVN3qVJHbaXXD1w12C59je5laifa3BsRU6/DKw/n/szJbn/dJHb5jqZMbrRZk0s6DlRud0LwIeJ
MVgK9SZoE8LJ0NrjbsF+vfer2wL0GokwlZPibfUFw7+ZCI1t+HRKf1QHUJKoSExeM+E5dP6Nc+Mv
0y8TWGbCIhNsSjK3F+fu+RAJs3/m64AA36mOJFFNYTWTcbC4a+va3QmJa4DgpHZ1KK7wZ0NIl4Eu
imf/HAxh2P2k3CsN8L/O9RPNGLUv0QHhHqCcTtSsIuBQ5fMq0Daq3fX9oWrRfxMYNhytGgKoVbEw
03uw8OlTLKuuWiT50u9wRixCPIvl+E9/nz27yMVxRb0Mxi9qIUog9pdw8uCDLXECF+0IJK9ZPw+1
kA94Nj2cTBZ57SGX/owjnamZ8oXmqYh7JzxkPwQsIKC8iGhsWCEe07fJM+OUCZnRI2PjQ4MpaqiU
LThr/JmK4vroAn8Co6d5kKPlQvWTxBwMlEujvW795R6QHGHJ6hlkwZd9ixS5p4nAixHxQnybUPdN
/XgVoGmJB9d2paZSuKm23wp2ISvmIRnrv+hq9Slgf3IxCvz8lTHEVwxJyXEz4pFKyn3YD2n14rhF
FfugFbiVjy+I+EISK7LZ8LZPjyflnnfMofgi4M6EEhuJRuSaOPkf8WNxlfkmQFYuyZP9Ot6eBd9H
oJ73PFsAF4hkngIJvqFvxnB9hgYh0FiA370GJdg70pz7BlIX3fZUtx713BgslEK/f+C0OQJCqmjh
tVik3JJCKxxBu4fxJ72CLOFsY0Bvqpq5vWeyYWgm1SWNWAraSCL9+J4lwP9XQDC9K8ivQc/7RDvd
OwkduQHHIeDVxhjKsuIiD+WTt+Nd1JufTgHhek8d5TSfHKYt0qISl2WrW5yL6T0hyYB0QGDHM9rN
iD4KqVvtlcNqG5sMdx6VSq4/XKzfhda5y5umlaqbMTQBQ9ubN6Yud1KsFphRML2gDiDmV0zy/jCm
rtlN3MXCx5h359Q5na69IK+AnIZ/wBV3Jf6F3Z2r7l0Z6sAzQA2khnclCLA1Cr2OaqKS0m1Zg/qQ
dqn2GWflPeN9UjhebWtoxorL92IvmLztPXkKIcU+4E7DQ9FCto/oXM7Q9F5XhhJinK7sS7pZFi4J
DM+AtG6l4slJY+FoHIlcDQzrT1hShdhXKW4IYK6SI79AgosKtQIJBEWOHQmJzpVExnQ2ibbEzRdR
G7S9xbe70fHPLiZ/vNrWv1xC5Wh8lUVMVhKw6drZ6/9IO3VIVqeNa6zanDZl/AP8tMwOVB3eN+Pd
kR1wvcaRtKqB5v1fhoGBHar9Kc+F3mS9+43U8fFDjHMBP5nmO+PdY4TUl4YBvBqPUBVHdzcUm1W4
p7Olece57vHWfmZtx6uZFMjF63HDSB7k4u3IVcdZsCcl4p0z9sIo12FvCGIwGL8z8HjqmP6K70co
RQJSgb/F9gJLRKCOxJjuj2TiLxabv0/fUd0RfxwLo0zurjZyOJIvbtgKksD/DsG7myxDDGZYtEha
j5SiSHs5Jlj5Hrih5Bvg38D+RZyISyypHL8vrk/S2R4fsce6u4EEAcvTu94fOOiYuDxFp1c3HmW8
OpSItJqQoUAP6h6JarClhuSYIkbAc8MD3QvBpGfknuEaMtlz7r7KdY13WB5AuY5aa77/Fbv67jG5
1ZSSqbo480YQG6N4hE7mINZitRynS1dMt4G5etHMvgSyN13pI0qRyiKMt2vm5AQbcEjKhKbhJr/1
GIukX1FWkwRpUUZxRY7gdoOMijy3lNgof79JP32nAtTSohggoFSkT+h6XnJzivUWC0Pa1W0xc02G
mv9bChv30lSW3W41tHFtzLxXvyNGNsbmZiZUUdpaqaZH6mOOvK5j4fM0h8dYHukbXNQoZvFK14ba
aajPBocbtOISxAkp1SLuprpXqD5vFn3VotEJN3SDIZcEMqnLOW41CXOaCDu7Z+MGsr4KrWFBl1xT
miv3Ehltq4Al+mx4CAX4IMoHuParh65YolxqwD0J2pFy2X6+lkH9Lkl1FFxfPnCZK3En7NPXbq7A
BFbDBr36EOExe2vY+ESTRt3gU57ZPZILkIUJTMYqR2qefsLQOlhe7z6+7SH7dJIbZcb6Vc3kzwg8
69KpIsiyl0zDeR4A8zgrqKHBmd6BUCrGKhX1IPXSCmLd01VuSpCoyoH0HtEA+kNMXmLhw7nWadzr
uHK0/qMxG4xSTXsoVW27M1ofhIJrl/7VrlAkpxhYo4h1eulzW/ZZDFlllVOVzgkCva1y9/75ir/B
xFqavBCDCrZX2ndjOxpbsY0MoXEJoYJMrneDbl2LWidBMmnTxGpt8nUJ8hdRLDN4l8TLgfs2fqLB
AJ6T1tO5QsBk+VL5xmOyG0uBDeKOVKcHDY3ogbft7ITALbfLPJn2rxkUbVtpyy59cQxQue3HdXc6
YmASzEs8C1yoRIKFKQcoedClYhPdguD0bbqjDOW4bXfBFVOZ3pwB6j4V30yDXHaGTfA63zDk6uzi
8N7XL9FeSU11bdBmUYBd6ab4BzjE6VXLurYtaABnDchR6d4Xk/bkPBp3jtjyVsT1igKkQdzvSkGY
aGlGMauBekOoKpCSGP3cfBQ/H8Bvx2RLdbIthFklG7hY+JxeWCa4+JatOvG1n3wDbWfrMc7tAUgK
n09pa9P3hUYo7ENxIgI3CndSO/aOL6TGBqQzeqKQ3A540q1qRwYh5gHIBrrsFW2KPMciDARW4oOm
HgRpoDvtVEFXbw39bm7F0GhQlxN08XdhcExISykfc5zXGzWUKVkauOPZN15rB24dHiyXKW6a0b55
Idali8kTjRilACqCkfChiA6UFIiS/CHvo1vV6dBk0VaEjj+ISGC7jlYbZ1/tbyttMjmeqns7WQLO
YoBg6f3ebD7EPqCyJGU0p5pGr4aXIcArw4qrGrcLxKurvEQPzygINUW4gcBgdJOz8BTvz1mVgvLU
e8uvaCNPdAf0zw3zMpIX+HafHbdxsQ4Dzi47VfmE1spdw2ggb5Zqv/kSol6cZRQZa+nLkmZgpB6f
pAprX5gZWjE+SimDDzG0kISageUhIc9DwjDGF6owS4Lcoy05DRh3j1A5enpfor8Qv8af2+bdXjNa
bpHuYX1kFUvmBk89ZZCu6w4fDiizyAtDbvlp/TXe/fAP5SjxSrTuywcf3xX3U/9e9cTxrGaE89ML
oUpdHXlfsS+d/NRX9LZAL/9YYLFP9kO9PzaJ87tY060EpT3Ei+QwksNviaXLmo2LJ+NZFHeAiv7m
w6fGhIZn+6PUV5tOQJkDwwxI2cwx8pygh1Ud6+yumlMXLjtnU2FdtIU2JWTZudK6SB9Ynl7uRE2t
Lct+dSmoJstjABD20S1k4Zc4kSVT5MVMqpz5HFCFb42FLv25yOxl6G9vND1HdJigQ9xRP8NORVnY
gozs3RjnNdzGpKEBhozDIqmdzfv2gNZZ8tq2q1FKvZ1NUEdWwEIspz7HLWCmYXeVLs+QAC+eEFq8
hDNrY0NjkbvTMck5TFzq8dZGNBSVb/KwhEBZ+yhqhogxIwrRyLGPEkmSs99z8i+YzcH+BB1LCsGy
HossO4tgCsmAeXGTqK1jb2kTXylAvECl6bi23RnjCtHtv/M4YlAutmv6ihoGVsfxBNL5ei0HSz6X
SnPYhipDWOKFE2wL+5XPvtfaZqTj85Rh1Ztl7Wz1sb897nfZmql/Q0EgFP3bNcK24tzeozbM+h9N
mi9bSZenUXZ/qgHuVfy192wdNHvXGVgEx81Uc0bt3pzmIAsdMZ5gEWGoVHy98U85fNrtx6qYc6sO
k0cyFt2uFFA7tpO6rmhqB6nKq9cio8l5xXBxIEs4dRMnGghPNDJUi44WAu88eMKEI+JxNkqv4Rwo
2888kLsMjTEh8QGYkVw/awyWHF6dXCP3u/7WJ+6xFyetjldqoP3K6R+9K8RLww5g3x2gksTWnFI7
XfSJ5J2XnmkN4AR02mQIPHfXlG0er10syQzd/TF9CxJ+CF308hXTVprD421ZjLqlLf6yzfu0vPay
G+TCgt063U8F9gORhNwduEftyM/7RjwcgJPQA7l+ZWiBU9fXzPCeqFPCrePxoqF12G8ZlVP7lhGz
LvOvNGxyDCwkeaobxhBI41fq9R8b6epzyGG/wgrJ2OCHIbUPVP6R5y9pUn0qO/iW6+bhbEXqMwjX
PkO+RDivH0g61QMwgLtMW+YfWj8Ixft30AoZRWoU/bAILvQzB5tmPaBq8R9XIKTfQ8IEHe6gAxQP
XQLWjM0YbMKaX44y+F/9Q0T1wUFT7TNPqEWBBO2QoKuLKpBeBBYnZ3AXLo+6hTgIY9DMDQIUeRrC
M9Qve+6SlXa2ZAxHQxUIqnlrvaooEv3qWdTAwquojWBT0g0hKBHgq5qCiLBOlgSLLFupRkKJNPIA
g/BguRYlHigS0zMnEyF0hpt1gOLuX4olX5+wlPwQJegP+KppflIkSNinz53s+lAc67nBHDESqoHR
cDR9ciHuvpnRizEziuoOTwGAWFve5g/GmV+bbHH5AWDpo2IUG5jO4UyVBOBbP/lvxlHriHPMNfxL
0gk1hTEOtDy4p5Oqc3cNDmlQ5c0bJcNZXrd7YLydMujhIVv6e1vfOqGtkHAZRt88Cmp/v+dxiNF+
VOPDY4adp7y6Q4gxIEoiwHDvj/Zr30E5NQi9ZYbnnmckgUGXqimGGTXrOmkMdSnxG5oDv9sWDUPM
CwLt7sMDPyGQ0OYqhPiOpybpC7EDoVnGjP6DrOcZ8t+Xz6CqpchCOlMqaEHp4huviL5m1jf35CEy
4Mcty3nViMpuu8a+naJBqD/BvwAuhDpXMffNm4hBi+C+93Yb9U6J11jAOC4bxHuyPh8XbgCNIwsG
4G+mtgsPcPfZHjoLP3lVvJgXgebu8a1p54Gf1GcKOLnL8Yk2mJDmO0vC+VdPM+SuGu9oSm4cx6ZO
ByuvJaIY9rFN0/ynzIxTLUzB5JGCvoe+5r+IOT7qDr4ItH4Ubq2Q0tRtD84HVpw1rMF/ZU00as03
pvWWTPHX+gzHLPeit/w7VAmmHj23Ml/STqx6of3Fg+IWEo+dzWtseQe9YkQCq61zSRj28igTRd+u
VsLILRNlr4wLjjmUiFayxQbKtP0ZA5knGe2aY2FvItCeRrSgtCPEURFJPgniVeXZaUGxmWU6+/a6
SiwJutjdq9FIaUgrbrafB4XBUPnRJ2ykfedvRQ8Ry+79zNdTMPusMPT4ZFNjocA1M/ZOc9oJz+CI
iMJXfS8GiiShhz0ZM+8urR2ogqRm/6Aeb5HtOO6TFcYJTXx4EWUgROBsMkRHPPVDRetprDPCOF94
CQRS22VwLJU/u7FRxOBE76HFSrfuAQ3FWco/PQpxcSKyZI9nVkYkY+L/cfY1VJIWqTqtJPRI0hzU
wLigEmQw5JLamRO91sr7g6qhNOnOGiK1mu1S2Mxnw2lewwnyxpAI1yY22Us3wg5p79LOtP3eM/I0
5fFDCAJ17aiw4ezIvN1ZwdJdAG3gPoeWMKkPQDqTjM61t2YBvUYKT58MYJJy0Sz0MWDaB+A3Lmje
Xm075Uuv6pbnCBaXHIxdAjKQJoC4ljctps7c0TEx2QS+yuXWS3GVAPHxuLp7bXMFNjGGZ8eLLm8w
icgQwU8N0Sg3L7OxOpyJvqwHe0IGnJb6SMU2ecgcxYJYWSfkvNvqBYFtO4oO4saSD7ne0t2Q/BWB
SdkHAuo8mSu9oBYqtBhBfCA2ryucGsa5CvEoJa8HSZd1kEyuci6U27mQDaJkqyLLzJLvYEKiiMh/
Tp9n2M5Yrg77IrhpF3Sj7TGY25+yPdG2tTS2psdACkWK9Q99jeBrl6odwmgYq/44GXtEe4gZqhOw
bz9G9SG8cwDML6rqlXUh9Nvf9sj6ZMoiKnbLQ4OSyXdjfTzwfNZPacy3CUkfq+4lwVv3x4kYxo7g
NR4YIR968kFw/0LGtNcEVb0Iqvc0zXF1jzIMj1DhmN7C4lG/GW3pB5Cxsr8b0frj7xXaQeNpJOd4
sZ7jGJGgLqAEwVc+R/LTmnuWrwrEJNdEe0qXGhyfSsxtFdMa2vKoYcb+qWyrlM9RdhT+Q9zcpWDt
qCjzWdiPuxC7nHZvOzUOdDKZ+Pn6GDGSEhYHuQZDdr3yAkJ+Ysi6KOBkWkhpfZUrxei9TqPOQeGt
I1+yudoiA23QKXfp+xXChBlKYswCEYSwiEFiijfCzUlakqVf93Pf3ULQMX0OvG72QvB53jEcbPLN
9IS9rXTrZBlGJQ7jV+w1jnGaABfmB3frF1d7yDqlFec6jieBlNJ7bi2wFTcnoHLvsIvn/ouyZDOm
hm+8BDkyfkleg1AKi4URekMPIn/YeRUrczP1UNLcTH9ERThBwTkhmm7mL/Y++TSJHAhE5Saav1TH
T+eQxoEaGVXbrlKPW7xMZSQ96IgPZUzuq94xbOTZXNCUlpc0l3Oyp0eQe/GAJr3z+4adU4CUsSap
KWp9JVjluG6ubRFyhCbu810YJADNCeJowUXFJ/RfvYWaQVBq2fQu+6BrR1vlg8TGcyAeKKqpptMs
Pvs7OFMzr7EtsA249UrxRHXNEpQsKvNqQABxmUu0Z/Oh2k4fdWWCLYw++YDSMbmYrpJGRytN26D3
b4faeNGo4d1l6V0L3RurP5MXG/RrAnlBTVes9U7OxLAlUk9OAZ0vaDDgMkdyfG03IOLmQ0BuJqaJ
51HXRjGH/Ph+dBUUVKpEgPRPyHry88499+C1KaK+VVV/0jYSnbnQ9wd73aW3+TKACLvpSOenvYLY
fSUT+kxzwmCofwoOSbsomWC83IqEPM4/8us6iMLXfZOmOspY2Nv9B94AT0oRDeQ3lSUD76jiweRF
zk6cOWyobkogoIGLB0c+ANzs9RrmZw7ojg6sW5XcErH1fMhgVL2WdijJYC0UFTEqBOFM1TBx5cee
Ivh6zQWrCYj8m9Tk8VKD4w9Gscot+KLwJ8mDe7o9xh+gCBbyGuaIWKAKEV8lILMw2J/95ziTq/zK
jMHrknMqhl+kvhoTIWAJkIybRVBBs8U8cpyNZceLAuJyZptpreUkyqcSZQMcYOIkz/v/+w3UZNdb
zv8DpUqWIAv3Vdy+aJYqESFqKFakH3TnnYXlNwv28MLlFd2u2H19FyfH1yFVflUwAU5ZwZWF5oyz
DPaD2fDzNQ/64/aY+lIekonzbBMLOspwj9jYeie9zr9C4P8eS8nZ25umpE3IPwZsPSgnh7HLv4OC
zZgFary6vgT5JxaXB3eJ9b8TNFLlD7HxfQlVMlAuogeyCjA1z1tfWZH+xqAZCLGRNsoIs0UJv4W9
Trn8vpV1bOrCVR0jmoOQtWXcnXMKCjZjVK8++1i/U4XKCobJPuOqgLN1o29vvhywYpP3ln2KjOCk
Cb0u6vwSeT2Owr8qR0s+5hS/X8FKDUfHOGf3oUXlpFwkoxu0pKy9oXVh9QRIRE1EUaRxVmGby3cd
ZXkCClPAftP+rXaTLLH35ZU5p2trMGCs/6VfV2ZmcFffGmtDuXm95VA1PU8XKKAdSJcFYgfruqII
EAZRKZjfFCfueFboEk4wJgnSVYeV15Gb1/OaSYMnVbwTZjJYB1dnmYvaFW5G6SPXHOsU8qjRxyvN
xImaLzLgMIneMlKXZideFJL3kv1O6v/juOQNgZrpFv/c7aJeDYLKeBtWRry0U5SfEND7So/6mge7
boBe1nDfLIDEQKN+r6UNHyRIYP0qTpNuAG+GrYl2eLeWlLLNIqZw0oUArDHOAbzRJ3oPfpm0feuN
1MDpJsP7rEnQkeGxPwglWbUZTpyg6qNUWoL3DeOTNIP8pu9etaJdhcEj2OJi/fDultsXTORjhUUD
hn9GfoDb5ql5Fq1KFifvEr6MEbAjP3VfC5VPwrZTbMtRTKZLkY9AKjB13+ioJmSJO3ZauOP/1JyI
IJeqcB91AJSIJj6ADYscIj44CZtiqIbtMo9p2MghcZCjd/210ijAC0U40Avu2WtV//O0n9mtKQTE
KdkcXNPcw9kqQYf0E5E4qgNv32RBPGshqR7SDSM03Ko5yt6zJc213uagLC71Zif/4C2IhhHhkSU4
AKKvNnKhK8wkXcomVOQH240ptsOyB8toz2HhQDf1Nzr0724CAPpW/xhg1TO9r//YW/KZcFKf2Dcb
GCXTXx5yFo1qQasJFioEV7WLGcZmruu+t/4UCePe7LKg48ESa6radBe/iB2s2sEyo6sIJ5TJfl8o
FrOUVhL7/W1Z0bnwoMlQVkOTprPa/vZNLHn8Taa6D8pQiBaS1QaJGCiVmYREIuTLLvsC+w44PHiO
jiU1tBZzOT+pC11oq9EIF/X3HjjNcCb/wJNoA9ejeOv0Dmr+D+JdVz5XA+vXG3Jv1HSZq3o4j7rG
40+nk9u83KyNfLHuK78m0jEeX87CR5MfI/+IYJHtZAHVLOOgHy9sYKXf8gnvJiUiU8d/BV/Q696o
J6drfCXiec6F1BCxh4s4fULPFMssSKVeGIo5f/uf2RW8fl1X677hh6Q0AMEavxzyAzqVDkKn94E+
0u63GqA4zeUfNcOiZobIamEDW/tNxUfKIpLbRLeun9PQF9w7+ZAN9qweqKu11igeTT0VRgGaOe/o
yuxrfYy4Z8SsyMLJ2y8BcGYCvesT7p05Wnz0ZJctH19cwXWrVQwhtH9cVZ9pa9y+KC1ZPm+7V1kc
A10vFtKI9DrpAWj2Zx8iL7JzZn7Nt6BzmbL2wjt72eiPHx24SDdWueuSAK0QTbCWKvqQsMLJ48Dg
Ir03rioFOuWqQn1wkqcI6JUFLmcywGzg1LWagYK5ulzSzqL7EeEsKVjlijgAr70l/ldbHT9RFCs8
Hy00S6dtTz6kLBptyvx9MXjfP0IOLSgqZ/AJdLGvzt472HilpecOU7xiCTCnPGmNJzIVtYEkKtMK
63GpeIh+IFMqC4Tf4BKNFvbOSySa15Xf97ICwhtuKafieBJ07cHIJSpkmJEdPZcz0prApAw8qQwd
e2yKLYqWMwp7gltEvCKUz+nhqSO6XdJ7GpsahRdDtHORAj00R6YBWg5Yli2e4HJBIfUVsw7qgtb7
RpUAotoA29h48hs9uqlHJ0553W8VkUo53pYB8oy2stnFvdEenJvw95XnK6ScP4iaCqBr97+lQyw/
6BwBIBW6rCGV4yimqL53ARpWz+lsInZehMJ7SWBfrbDgrjasJlSoMv4nxmTKGowZ0IkgP27Pt64J
ejB6AOLdvaVH0yNWtOi1c9aQvhGLDW0cF5mnvZq9BMAiPU6UjijYTGWyZGeOPR58wQDB8l9Cls0m
1LevEbQcmjRixQ8zJ9AhC47zET25NiB1nDqqYw0ILrUUqXOR+E0mHAoiQX4/lh+sfr1Cqecfe0fe
dTijXee1wgl3xuBJF59pW5+A/sjVAhdTge+kJaPre2TEIU6qfCy0Fi0muqM4Gxfem4uyxTu5UiqC
9/M+oO4jA9MEPKTx6dzhcTxKX4jYcA0lKwIIvS51NdsHtcPJRDPFy1n1evqeOJ31Irefa9GmVXUB
Z3z6MyZ5LoG7C4EYNCdBqH82zLfVoQbMDUMkii/gVWSuKSu0WDVqGm9eUm2hwTLoztz/1umqjhfq
/My9vCs/ccNPoS77gx9NDZi50z4Bxh1tHYdLNFzJ5iB4KcBKhu4fL3mMiLblmtc6YMaLKaTeevt+
iSHEFZOOc/N426e8c7ZB41qVb7PKEqUR4OdtIdRJ1Jt2zlRln/VoTw8U5smaM9qOimrnXSeFQRCO
AsRb+juP+DGzrga85BAobOTafbgTUM04SwSAghW8TeUCc9XsqNOpPDYVOtuwg94tHCiEA/YH5a6j
LEJg7R0gBM40sJ+2FOsC4xVrOjg2kQbivmeY7fAG5LSXPX5cOeDRLUldMlC5XLBgbwTm0pfX1WEk
6HYuY1ObjAEWZZ0kUdmotfC0KUZerEnL9kt3ru1kqBULEl3jdjOdEfOF5x5YcGeZ3ELFrXBlnowA
ztaFYDzMQDGoya60ZhyujRYXmppBCe9wtQ9dCv14nlEaYAUXte331QHKmX2XyiUaOgzKyCkP3JUb
X2Vdy1a4beTQh4ytCHjdMmiG6Ne2sbetRa9PRUmxjxjv59QlJwIAAN/GQlpPpCnpQhhB/7+lmRie
rbkQllwQ38WC/qZVn+ubwPL5FHHone75dhZjEaj2Ep3jKxBAyCvqbPP+GUUM6p+Wob84Nw+ZHGNG
xYlanaugtv0bzYhYPW1lY3Bow59gdVq0mKFRHaSXbyXkwa30Oec27P05VCVuP6zkzuv9QBeDX82f
kQCgNy9AzWl5ehqfZn2yOFpFzeRoGtVoFIkYxcWoU0PyPZRe+RTcJxesTOsdteri3vFtJ/5a5kFf
vJAhUXjnHVE4NQTgsolOXR4v9hx5anvhVlD8yqT400FlNPX3psNeA9rr7CimfTkCb1X9cqEV/qAj
wOz0k9OgZVld79K9pAtJaR7rV/d3SnpQ3izUdk4F2snHHOqDADf9kq+Ll9KIRzCatn9OC+WHlbz/
TBzelVK8lLF8gmqdXbdX3ir6h16LzodOUi99zueN4s3I171hzLz8RkqYCE4bJXdFJ1xqDDzdk54s
kiNnfEbSQ3hm9jV8RDKFkQeFOPFvWVfwjEtaB89G1iOBt3cdCF9EYOQvxtJn4OtzO4z/YkYuuKPF
88vX8045q+syzXb95fDZ4+ntkt7Y0MTyIejTBzlkDzJR6aOR7e3w7Puyd1fkPO09cUUQ4Bv6aP7C
wH8Chbte+RohdmJuEHtQVCgyEB1Mbq5Jc8J6g8P8QEuJCmwvSWWMfRYgCC78EBikL3pxWzBseiFa
/oTDNZ0BkMXGUsqLp6euFYw2vqJbYVeKo8k4WTYqNL+iFV06PckwFudYET2heoUm30mFpFZVn2Dx
x59UwBUJsEr910GSf5J2SF7vcBppeRZ7Yjf7HUyb2RVU4+QrCPwNYdr4OeqoEoMpdanWRN9D8kNI
PuPCJVP1UNxLLkLc0VLl7xSijZ/LcWMgZNwZgUaH2paq4rsquE7nyFpjEJHX9j7kNW02QmpDJmyn
+VdiZpvXCDpFCzibW1YYYkhDEfA3j8BmYGXZ3BbM4MLUA5HQrkIEWAd8O7gJz9n/gnp2X4HxynOj
6lQPJYPu45wo8vZBmYZ0RA0uHQ7OqYKugSUsAjWXgjbV8C9A0hTQ+/jeUwiz418vaVlOK3j5ZS0r
CJXLBL8yXWVegXAjJXRLvsGRPax7iwSMEXRCJ4lBDk2L+/2mDHPfZU7ZQPgp9fD+cgRFjGoUkW0p
yKP0HqBueli/uu2fBXENJvBGkUKntoVzc4fbqDm6BTzEUvaenvf0EbXX6R0yi4HGlhCquf11Fpk2
82I6imeqRhZEs6js6+UjP+q5OYwNixdLP4kNoPCaJrureSQlEjRNHe9zMgQPSFRZWyYYRRcj2COl
511jECBdyX73cwwPjSuel3Eot0dW+6lRVRK/3L3ny2cVysyogm1LFdgiSpbIta1zFE8E0k4lbsur
dhx75rSumSR1r4R4HZEfMdBeEmR5ZlHOgtytox++09CdlLNTrEZZdhhsJb2VZKAsviRnaEUsTyuF
pDgzLKfRjEx80+yYrIw5ExETgnPKmi0ootCafDLeUXItuzniXz0PGqseEi/RIg8VN8tjIbmW9V3q
zUhfcG9BYuAdDTqaYRi2jNNwTdhLmN/RQFCuWDP2ilSvgOEYDy8OeTg5hRr4wCvGLlFUPaD+g+BB
DNYomnRgHgBGA52FIYnYjq7wtLfbvBr5Ep2eOmp8odDp5yeCHMx3bMnenk31RRr+7PBFYR9EAQlO
dF1pKoly2/FETOZXuLDn89Y/Y0R/L6J3SX475gW7olZZdj74B4lYlKwgXezLwGnqtE6boDz+lKRL
npu3Uaaml512b6mzF/Vg7A8t90cSDletiuWeTsx1BXv5fXBFmStCnYn6i5pnx9uwKz383Mil1jPf
Nc/5uXFKbm4cPcZBrQPkaJMXn/BC0Zp7l9fOjLRUrSYgWzwqkewwIqaFcCjYk0/OkyIROnXPLp9x
hNk1pYbydesSumdotxIy+d0M93xgyNCJb6CYGZaCRqmGXFkOD1sBvRhS2IdNm9H9P/clj1j7/kJg
9jKsHjOtDL5AtojyX7w32mcX2yYjO7lbMHW/TPf2W+ef+ZKe9XDfU0G5LUIXR1/Xq6n4S33Q4ugC
9EjNrSWvGJvFcNP7RWl0r6aV/wCPXTRTfia1O6mshrDbcPTluZLUxPF0gzH6c7cGiMuvVVuF3D1w
uhOzzwSoizUVgEj+epA2+OlLyRTsC/qR+FWbDE0nlZS5XX3vWLpJHdmGHjTMdkSXK//3IzsNt6Dv
6DB00dakT+Yr3tcQa2/mfacC6YCR9tKPTKn0uLpMtAaTShjf/7YYrNs0Ixyqoyp7V3XmAVaFLm4j
Aw9wbnbb+OhBDKzXrSlMxljy8hqbpTXIX4YU8F2H9hwv4ZFnoANnwQYkSBJFwuS3Pqrwwtn6Mpjq
NfAqe/K9Sk8Ol1IPNgNs0pY6p8lImlKNlVCXqGlTqvZ0uRrc98XrGCTKMKczydraOg3BhDxDfDXc
onCJ6QoWYM44ESjII2tQk2xhFqJmG8t6swytSyjqHjsnD3wNwFf/uVw7AxruEygRoX4AcByvF5HX
i7GFuYed6q7nqqa5z8O0+OWqaZQu6oaB5fiKFgzQ6cOyzsDVij4GczUpkEjde8S1bVlClE09mapB
FdGMmXLAkFSVeNm8VfdOEYDghXiiHxDw9DF8rghfvSULFBwqZsH8J301xtRd/9xP6PbjC41mJjL3
xop62y24wmzt0WWilV0bu+K3XQrJWomEruiA5RiFvToLWaD2PzA0Z7I8+5iykis0Qt0ovQJx2gBG
V3KEdQfz3uutyK390zQWXjrNZw1WX4z1CKT6MsDWnHsUjAKysCvD859c8UKPC/BM52q2DI/b2ZDI
iBcij8cqdKOZ86YcvyDJ8UNp4gUicIAj3et6izm4n0RLDUEm+9gdoEBx6zUS7Wp1WwCs0GG2xkY4
0ggxmiCXBmOA/a5aSE9wiY+tOofIPhQFhLU9Vbf3gZ6Rva3C290LGdxR/9ugv9bJnb692D5evJQO
w4WAyx5x+1jKy6/5hhkhB5hrc7XyZaaF2Ch+T6wjr0VLn76qjcvIujQZ1CtT5/Ex6iJ33ndba4KV
chlF4dkTL3cVX2QrLMR5GV0QObz3cdi4nLgXsIOQv1aY2PH/F+6U0fRo7pagDgwgheu2z/kpuul+
UjSdv5Opr4Xl0bqWRWWeZLR9cNJUMLV6HixRnRghgk1sahY+Fwn0c/Irobhn14YtbKk7W/Lmv8PD
JwfgKnDvRQy3Mk4gxwdYRE/Gsiu+AKDkyPMyHpyscragYcrMl4fKNl8d7I7G4vDadK46t9Qm9lqx
H5e+VphY39XxHZrqY8AXLQlUSR5v6p0AxwEolMOWa+dcrvxj/yaRs5HOpvWx0p2Qv+ITazZe/FOt
yKyvmXNrjAIX2aCp3vpnkbf2Vtt8QHoYN+1JOU206SMyGbyeIfcpApff5psPkSB3eRwsp7hkeXuu
M1ek/ULXVOMBKP9GoewCQTly4Pc5wMYaGenIDs/zicBuboV80uVVV4l6tCI4ELO/6U/79BoOABIe
9yS6gaOvmg4BZ3ZZfV+ym4/fWULrm4jWdydi/uKaWkxCWDiKcZ3uFwhvx7TU6irlWIyqp2sUgd+d
v2FhukNzBx4W6QMaychcCPuibZzugO46wi98KudYkYbgTvfJ1v4fWDOIvQY/3z9eGAbzLPvIN9L9
B+kVpna2n4VaY61c+gwJKv9OzlF8Jpgcow4J6R3uR6UEzr1nWNY/3xr0M9qkFNAabqauB/RM3he4
hSEMmjj2nTVLJ0yjmFUSf8jfG55CudqCtUrr9NnQLGhFnqRADnyvuHcjmdXIzTtCDlutMojK+q7h
J+fQH2Vj8muj5T1ZxpX0RkPKSnGEjMToRUybSGm2+P+l9Sg06qSOZSFhbgWo2kVPb6NHyZPlDGNL
ENlqM6hqLGwdqvbitJpLY5hnxnaVALEtiYVj+vDi6TVMCvN36PzwY4TItONRJi6qprnKCrV6oSaU
Cvs6gKQWYoauWXVvSyR9NUVN0EfCXsGfJybSVTgQmcv45NT5C+zIR8PLDYDS87JyoGMDIilaHDfN
UQQEaVoXsk4FY/bZ6U6C3BeWyS6Ul6CBloamqKWvpUCyFMjAh4HyllXjKMJ358AjwNPErblHcXoO
ptxuDp6jxr4HjZOEO54+yaAxui3AgEBl/X8RTvaBrWNVqDo2tqixa6CA6KOhUR/18X6kwwJwwiF6
4Sbz01G0wLMiaTRFg2BnFXifq8f34V+4yaRjwxmvUKCRo8xDrVhQL3vGOwrD6fEHc+ocyd55usvo
Rc8Qt9p93WGilwDDnKELInfvl3lK/TUxig+lMmble/5MwQZOB47pK30S7wobOPYe+ON90xslbnfC
fojvvQqBgwOdjZAa2M/+CNBmnT+nX43TYlIOxBfTu9uWO4kGWRhowIfaOaGLZ/JeTQiIb2ZxW0tW
bo/tAf+VbuoUqtn5TFaTOE748MYhST2pyueKMFvF7DDi172w80K47l7Ba/jHHqfA/uU2T/uccGJR
biXPo83CWFxVbYAq4DKj3Uvp88iGkLjGFDnPrzijVATr8oegzWfGCJyBIau4acSCenCgMDTJe8Ed
6pSECLvyeSIRhOUGY1zhW4Kx6Tv4KtxZJgY/AHCeGiNjq5OaMaiAZ6ml+TGavk1vDFLlOtaxv6j6
HLgsQVODJgvIZsjedRJrqCsvWyBBOVzYtrY66wcqsixVe8HTVFpYbCoaNnhB21oskBw93Fn2xod0
FrUGOXLb/NwwL9xvOJm1MwrJUVQN+W12TPLRtifGFQByOYCMN6lsxXMUR2QDCVdzNpXSmF+2775e
40mFsHwgkpxxaT/EwQ8IZ8wZ+ETr7GS42hPO4f21Qz7FvkEN/WErAq90FzwS/CNjVxVIijYGpv95
bcrPSJa62PQwEIuNQKHg/c1YRT/lHYt8fF28frFrkJVoFOphFVQSSor2dMJk7upP0b9VTrGdUehg
VjbiWGJvkPh0RKoXNi+UUDIQfKFPtCWR0ZKKtxTrXm3WKZGQ59C6yljO1mk68zcghSwEi0iWQuaN
HI4fwDJpHT2B74FVFHy6+mIq4poHpPsl1V2taE0Y4pkS0C9yzhUOTvK77gSB1HrGmWQXlCc7n8Zx
pHsBayUaj+oigo7NDuovff4lMvT90UVD2HGhmDPnG0E/i4fZP+r7Tnbg99acBEdraDMMnkwC+e06
olEaEqFkxx0IL90FvLvvWZVRHIYVuTCem720o9ERUwHgwnnYOOCMi/vhNZK3OLZ5KyA0n+2gWdWO
+s63+1h+PEBZxn+svmf+0KutGFJF6qontJyo50EKiEE66s2GhcYSIZAocCUuoyUNt7Uo9MJdtqCr
E9dAAn6Mst7nxxAfgZQL2V0KCImsc5AbiaCw5S3WOU+SncuAn2Ttr+e7M+VHPKpDcwqNYMkMW6Hj
ALXKeqY6lLY8c3OGBnFJ+VTb8hsSK/tgzRppTutOUL+gXEyiQILa5HCNuaVySS4KyyZjNa0vqeMn
2/wYXMWNN3XIt41Jp7vp4shEyTQgyioa9FVYvuxlz/cqD854VL9J/v6WGHjQ/pnv60gu9xLhO5L5
9YDvTvY1j15+mEVbKhv8wwHjyWsoURQfcc8503LjzrPcZ1XctNf7plkl6qKfy8+2jl90miBIcsRc
owU7u5yBmz0etKRctVeayjfUDWeVm95728u7x8RJMJISeemB6ovi8I2MWrh86+rKpijTdufl/INV
xeayo4NhNaD8BshvN53QjnQ0EhZOoP4XANsK7rIkNp0zK1DzklMm8GCOb9y9WC0eyeYRY4+7NkHf
8DPAWrTBx2lFoUIR+SERDCyWRxSP4MPpbdXRot8lZxpMVWsJQTQKOiOS2Go1DV6gJGxU7tLD7ryu
31nzXRJ4hQWt5GAisHKPtKROo5tereeiGmTnAcJMIh1/EKHel20lASdAr6ii5/tgwaiqgK1/bs0Q
GuRKMZm460eKDq3C8Lb44fRgHCMguQh+J6ucWIIu2/Q7kOgjV6E5ys8p5czY2SN6Rx3q9q37Kr1t
AwwN790QEvGhJlUoLjH3Y3k96p0KBu12L+eIXiXvnJ5h8SS0sXD2dRb9ZAHY2O7Glqpe5KRdRDe6
kN5l5jz11rFz0ObtY5R6iK86vmvO3s6zx0IqeW4qYoIUxhS55ie0Pta9OPbXLw6Rwfvz+mRKotzS
Hkb5X2gOiliItwu+s30Gmumiqbf/fJRYPiIkmPILQc8gar3wW0+sAYnWKYt2GkxheIilg2Ki0/Bo
XJpDjAz0P3/uHG6ZPDN6jsbXipx58Hs6Atdyp+PD1VMvIPghOtqZZ7aHfBqGCo/MvHsz3ykxHMy3
ae5w8PcH/fB5aUPt7Sp3JEXY4gVXne54CEEBQ9fDP/K/d7YTMOwMSbS+zwGxdIvsDtPoiLNbWaT3
eDYbiM8o65Ajj/TnTJvGYsDZZEA2ZYMDqbWMquMaJMixDI3plVpaaJOy8FhOXTNknZVRlxzmawIs
7YuEp2OwQ1t1okz4VmApI9s6r4eGuqU9iSQosPxa6HbVzqopcSVogqUCsMnxqfxLUMw9ge88rpRo
0JSGJstfYhl19KsDFafs0L54/ESPpUcdGdcxAuOnovAfBiPjerkPoz0aD3cK9KWNa+YFThPCDWT9
9EzixWmUXVYzR5LHhsqH/C2j/yWzZiTWp7JLc1X9S7asuTiGnDtfspO7LXqUf+oFuPWsmPG/KEAF
Aqo/v4kWKAn4rR5s12pFwa0Dyh1GYgNOiXJvE3W9vKpMZsljqnpSOocQOm2zYuWjerj0aOU0WtzS
nG4FwSH0ZYCgC60CRpI9Wn9bMFvccOoCeWp7QuCD6MYNp66OSmyMorgND35s4+IURXlyCHeeg6/9
MvbiqLMXLunhavEa0Hb8S8d/4bKMZxZm41JxT8ZITWZzhgzZK/nvhKztuIyoGkFejX6X2Vj7GYJL
oC8t447n6QEojF8ab1mo4RybDlR++vyRh2QkEC37CkIprLW151fdyE7zeersE3X8m+e3k0LOpH5l
XYoYc7PeOac9nmryV5miZs6FW03hNt18lfiCzCEZwE+zwISMM3ywXh3SFa4wHxavevm67ccKuJ89
TnCDNp4y1gQdVgaToYRoLClwJlposJiWnkqPSW3lTj4UfSHdVEObcDCb6MM2gXfQLciIGUwcawhE
hsOeVIEI6I4mpuxoJKQdyFzn6ihL9Q2mj2minXTocNkLTBmBYN3rRLz8hlq5hpAnhoZSPmVD1WSB
kveTUH6wOyQIg4X4HAcuCFjAKWHA/HDen5su6Ab1PTdS3qBjCQ43CqaYVgl8ctr/Blcmz++mzIXO
R+/vnbu5chrBW9IiYxvoIO1uZjSZ2l7lE+D0RfspGEnER1ZZ9fuFTV0CAER2Sqc3hCzfEkWbOeBb
2EqH/hOVhAJ83fG+XZqUzmsPlfJ9k+0DoYgefDswPUp48B6gXcM1Y5PiujU7WowIzZGSxDPLyWkK
Mdy7jNpjHroAoOkn2aV8AdpGFVFCBpeIO6UaFTw2RT7vy7GoIGLYq3KscumO9pitVFacyT0dkIKM
G8ZCi2GP9U6RjhgNi6gM+H6+1qhvjzPFvkAROLzrEk6s6SHrB4y1Iz8/lT63kvmQXdIAE6XmV81W
6eOYa1VnQdG4NHSiOXeFXbgi8JID9F/TWQLE+VjhXwrEiZkIMuk6KMn/ESXkQzA1FN8YaeF9158Z
IwSQo+RV1D6fhvpvQATdmNya5C8+nFpcPfb4E/gKLzdwUC1cOQFZGwQi2x9nOfoZoWCHF1tpeTzK
roPiQbcIpwZXASxqLrFHD+zUl54OkNEDgstqVynmiATdZZLpc6w8vuCJlnaBqFQMg5ZcCDXsJxh5
WKjsCRt10Jiuf5OrTvBOSUym0QoM2UbzUKiu82xcMMIn0VT5PxrYRURt0Hsj+RsVJ1R34NPl5Z89
4glZLu0Ku+EA8365BzSFo9aB0gq9Ma7TQYSuu4AD4XCiK4LbmpwAHaqYqS4etVAinaNyVLaMVeAM
Mxr0HEwPyJY0TxEpy9S7g1vsydN0m23fIsMMngtZids3q2+fFceRcIf6oFH2CfVCSJX5WFSn/HOR
kp7MA/onFx+iR4yA0Ps2UIFYxHuH50EYz2R9spAesQ4IooWdt8+xVnHL4QsQMl3gTeZ/gFfCcv20
mUYNUyHu+zgZaast3+UQA5y57TfnRtr5zkzJDT0xl6Y2IHGdf6O2qu02Q+P7PtiIA/9yXqOxDdCy
m6SzVae0QAIKCFDaM22vUC39fSzkOEeWhVUhXsBQZrzyJ67bXmGn5Q/94GHS4mrPyELGLteUpvX8
OAh6hDYZ9B1wu7foAdn/DEZi4f0OL+o50iwhJi++jrxVXFzkYhw/NxcZutByyEkJX81oMFQqZHH8
apR8qO3DVzKKPpll1+k76vfXpACaAJ0DRmoYsAqxpWL2qWuBc5vrk5dUxSVMoDg48Q2NBGfy47z+
SfEN2/ZKv/9uvp8YdltMHSiH4MJtH58AFZiRByQ6Kyz1dvoJViK1woeo3/MTIvXF2Pa9DXT7c7Vb
QA5OWZO2eRN+gBxrk87/ZeTTsOGJNSSQEAtLH8xIwYLppXJLUwGMB8joy/CCNluSiTB8382HJGCo
jrsKnKbaYW/FdCzsBt7Zz/UCypEf2pUvOxcH34KjFYbGowhhsKe4J/g5451oAQFC2vHT/xmqOEX9
v7HispbdTswyhuHUPt+fCo/2fMefuV1wPZYpR1xfdKMJN0i9Ma9dxxhpSBW1ehKk6Jv5rVN0u/FX
crsX0e/H3itlRV2WakVOEo7rHEWu4OjFYggS/IVTA9K9q3vPkW4BmtRaa9BonXnMW0er4boOlhka
Ph6PgaaOOJfQbU4WhextG8/+rbrgIMABMDDom4IyahkpikOeuh31Cc5Qi4jlPZSz6P1HGf/qlPvy
oNudIPWjQcBkZ9Rvb6hxmXcuNZJpPcZ0Sdg1/1i6xedPl/QtX7avfXnKOeLfi5A0+f/RF/3sLxO7
V2M+JXMDj5QVydWGXJuTerAsICHlnw/IyEXMf0YE47JtOR0NdwXn4HjH6K/yi8zvpGHgEBRsTqOR
9J1AqVQXgz9AflpTs1ry2K6KQeOrevnx+Vq9wvw0CX5Pyz2xgMdESEXqGWvablCObhFqhFKXX7vy
0tSoZFg1vsuHt3bB3leHvl+LTGifrQWZf3amvQEZdLE+9HalS6UMhopuqPQ7p2R8Bnsk8IjAA2d1
b2LCeUkj8JnPWJJtVWTpQTxrsqZU8SjeJlUzCblEnHo/zfVp4GjhKdTAGdoUtSkOfBU1wtU2Y/m0
VV6pcn3sHCmwO3sM+z7B1qFrscxQEUGU+JS7JZl7r82IVcgDaRXElesmhYlO8e2i/wDZVoAyx8Yx
r43EXsd/A3BR3C/TF8kuTbRtDEQs6x8ijp8nG+NPlXh4GUTGPVWvkKrWbVavM5MYciHU1bH9e6pq
c7VSQTKpZj4TaUF2XN/O8OQVdB8G6QAg7SLLC7vUul9Ues9Ni05VrkHgNJgGSndsan3ckl/10yee
U1DgY+5DtKWEIJQ/VEnSLRZ2htKRlBqzRfAnDx3TkUZY1LjCx6Z33ZZAn7kRI5KoyABgvDEvIXLw
wYECGn6hD2VhvDFRy6vhVBjvMtzwvbohVONQLM1gaGyTHSKpxlIU2njL2nC4edsDyugG0XiqccHI
hUYZQO1FlI2J/UOwzyiKFDM8xoO4HdTiDr1i+H7vbxi9pYn+ZujFiIRnt7CRPYNIoGVJGmnG0SoP
l/hMFhWM2WqG2DNcbYU//7qUB4xpYFSAowyeFTBcIgV95TDLOHxOFI6JMdU9atoEmayFnKlJGRKe
SSUMlGu2PcQGvrF4vB28kKipCCGQ+oIcxi7vdNKaNFeeCb5dT1jKbHJqliTAHkMThYz1S6bzM6wv
A3hQUaBhrNcJKvtbJ2qAOzqw+oBCKeceQ6+Gnjik60szRDWtuEnxJlZVIpui8EYtxAAV0RE1uakV
Th/8i/n1aJb6SP0LeUvo36cspzdWlT39P+JQL8XrccX85Tt3jIGrJrlgJxcOHR7YyPoRcie42M0z
ObHAKJ7yMHtYrN8YVxr1VtLmL0plbJjCh5ikJUOySFxG3EooXIzFFogepbV7dswxB4t9ms0cBjcp
pydCgUW+oNgm6S7YWe/klaALL6wQ8+0lF36uTHjAYG4ZpDm8SmW7yn0sll8RQrHzN5lQzwZ1ZJwh
rkBdrhnLTXd+p7IeaXsrm0WxFe/JuigLFAoN4i/mVS3cVdP5duupo26MG4dzqV5lwVLb9E+DClxJ
TuX+0tYx5hSEbNq27uvENMIf+8OisVy+WHkMQ+wYTyM0JRCpdIGo9AY9vl+lWsTFnGIxzpSEWQvh
36YimeuzBY92MNJ8di2+m8dw4a4HthSvlTKjaDa5J44920IBUAtauIbfUWWCpAe9crlcVsj6MvRg
g9E44/bLWPQWuNiw5F6iktUbupctAn5IYxWGIxc+g70GLBBGoaIsn7NSehhtpxSOUyWpm2+I52+j
uhTynjyJr5tLq1lc1nPiF0hQQn+yHCvNbumBfCVc2xDzE5dvs8ht3v2h+vFmXfWvxV7vuDIxIEGU
ARwA0W9nhpL5pguTDiFdEVDrIFXThz3aDIuGnvJ+HBTj2HBm8+4nUOzOeLhcyp3BJPal80gXxewJ
WxdoC66HRgsKRcVHUmRLCf4BT0rFQki+zRwYcEdfYV0j2qb1D/q+RyppJ5vGzayFHMpox8vUUhkC
5urkZOfb9gEz5z4+NdBbL3gz0B6wa+WKinncakSlujyAQHvjhvfSOfViXbEvcmxqg3Rn6I+bJMhH
cQt2oeQsdpbJrROEDOqJZiThncAMOqvFVvEjYCw51+dxXWYvN6YOX/s72IcVT9OETG4BNKK3rBK7
18wekx1i8nrQRgQysbmildiMHZuOU8+7ivIKu2mGHpYr/Ic91180BBgiecLRloyJfow7xGkte6AI
ynBmfi4KUkRRJh2JAGfPR/pQBVOsIVsx5jiUu//AHGBOjXVEPMczH0hxQEQoBELWFUchXZC2gghA
8ltyorAqGNy/jdLfHkc3jxKFgvvdZXL+lPkjrqliZIAbdHQcRJNWMrINn2YO3xFay3pWys3i1Iea
SF0pmSDMvYuxSoqVO8wSIJsJ1OGDr6Pi5Am71ZFtn7sh0kJ1FeIaIHMdg5KnppBX1+NnV1aIP79E
4QXJc8o7r+kWNNOPF9vvIcAc4hF38JGoVbS1PFc0w8TdOwyKFEFokfhTC4SNQ/5Wn4hxO2Zqd9Cc
AO35klFENyuHkqPYt3nP7uhzjdcqD5mB3O0UWs8BRCJ4N6Z3TzER5uoXsYNjGG1tYA7uM4UrPwIA
bL5Qk2AoN5I4CNmOnWur4qQW0JSmrhM7cVJuTw6ttTuCBMZGqxdZvnSRan2mkXqUkOZtrTIAg6mD
k3716EL3Awj0JLMRByzh1bajhQu5IKpi3KqzkHP2KzvvuuW6CwayiQ16zsRK5jnY9uM5Mr3/iQVi
oYWQ8racav6cUpIzUFlPXG3u+pTR8EzL4jGsa3oROGhzI08p2L+f7F8/aPLD3zlnE5iqZ0IZwUhh
yAhMKAPIju1qQCaeA8KGjxbP3Q37OuxVFZCDouSsOYII6RKhkx5X206I9suHJN8no/Wcwc+yIRGV
sbK6QxrDaxzcBEqSj4fepm5a5AmZ0kcBshuzJFreuFv39cas3lI6Izq3zl+Pk1Cf4aBghpHxbeH7
JretqBjFNKqeBdur7MfgmA97xi2M9LST4Ey1K6XLaDc/pkTRyYshXNsAbPZfH+wJR5b0ptCaR7sN
gzAQB08BKZIHC7vPLyYnIB44BJw11Dup/bgFAj3o5PyEhQD/Gbic+DeliBkw8eQdWsCYDVai6OQK
7hfcxD+/2AArezpeRYkVdpvbMm9qgQPe12cV3ZosWoQaF93ofw6mrPTgYzPmeFBGJvfphzBENll7
IiJslN9MiR/s7tPP0HA+sqjw/uZmplvKskqwGpwwQAqYg7+Yjs128w1KoDqc136bsQhT/Uiy6JCT
i//1D5cvrUXnPrI4Lxi9sxXlCTQk/vSX8/4s4Pc40EeWltFqbIOi7NmtBCtGnpAe+WolQrLaGhI7
Lkiequ1DwDGMVs18jRqibU3joTzUTHBUUfJVJWAz7bc6nx6/17f6gIcU0pPl0PNgsc6sEEXEASPW
YsicdHGDptC7zwPjZbEeDevoW7JjWYMzZAVulRXa79rlxEci98z5YysfbnjsBNL9X3tiXqLbIbCp
7jHi0iPt1k27nJiKZ/SfVDQ8ARWxJiyMOHZAsNA4mPoByJRLznfH9UWHnSq5Btb3LPwtcfJw6A3q
MI9u4IHmqz7HjOb8HuwTw6yW2b2tYw0t1nCaV6GLA9bxno9JNoeFT3WxbhzeTZwfmnmo6KYEcW3V
P231i121Z8HeTVJlHTg1b9dLTR+oIRwkGncSJ2aYXd+4pcRf+E3a5rtPXgR66AxkfVIx05rGep0J
y3fsU3lgH2AAj5kJSUAs8Ye5GsLQ6yEY9zG6hLQVAUDMYZmmEBWOXGcbiuLS72NeBYufwIzmt1gc
6StjLsBru+n73Yi775qFUtg5dwE/84Z4V+3Y+SdfY9UiEJG1QIaTKbqwiVd/rOUlGrQqQ9AatSbT
K2FM49QAwJR7no5kHgn7ZcOaYefUej/ONtvkkVBF/o4ZbwHn/qAzHqdi+iC/TkF8AELH1+vlelcY
MjW1YpLsbTALhouDQj62O7ODPt5nZ3Ed5jqR9NKbzOpzybpWWur7Y5mjlRkuvElyT09C53Aj4QOb
W+zsN+m6MQlF9xMqiRcejpvs/WJW++B4QDezGVe+sqNNGBzmq0Op3RYVVo6S5RNoE25mVqW0Ix2x
j02/M7YIJDB1aipLvKFH2S0b5tGCBunZTtKJ498iCeiKxj+9oLrs8hljdnEgJagknMuTvKWUGrFl
RLmHSWOtDGPPy3BOBYsB+I3YOOD5kqY8ANnpLym+yFqhOTjL5hnvxPsPv9A0fl+QStjM537C0k6w
I3ozXfmheOC6Bzyqyk2vMAiJh7ZFvQkHXBOYovFj2vzR3abCvZ6g3VGWCX4VGoUGeRuTxWCD7Uqx
Rlfn98PNqC0lgc/UVbXJfaKk9wi69j+i7hG/8i6cA1mCd+58HnrNAkAJgB6WJ5W0AIXvJ5NACSGE
cixzFfyGkrlDBOwC6nLBYFuhzbjX/6cryhxrkjd0li3WqYX7JYf70muBy7slSwMnN9zY6OpIMVsc
pS+EiwFyN9g/U0RxnVuFoTqvy804OT5KYCeWSMqeWzx9nWLIKzqegjKfTxq6ECU9ZB+FhjnhaKdD
Y4SUPHvYoVsKQ08yLNAjKWu3QFFav+Z0ViFl2Cts1XvS7lC/OxuWH6VUky6D4U59udlHXngIORwh
G2ypAaBFsIrI7K7798uvuHydMc5nSx2naQGGykbYMgWdr8lIioMaViTaO6a/z/kQABCvf4v42PfD
GtTb/16M4v8cEHk1OAtsaVAMsBaHncVb3uInbBXiXUESIYaWdznoJwG62f10rV2Souhg0Gn7dY5D
dDITj5uYvpc+zl12f1lvTlU/CJ38g+E+Hv717PZ6m5KX8rS0yUmZQ0dl+gDSRijEs6Vvsd8Ujd1U
hinFk4GIYiSI6WRBJXBUGG/PBitsSy7pxZovYhUzkvWFZq5pw5BTO97aurmvM6Kpa2BUhoFZ6L/f
+m1ijkt/wW5jN25qH/vhU0BmT+uWApeGR400MBFtnlWmRe6K2M86M5dRqm52CxMVStKVbBv9xZUe
ExdU4lBHfPLeWIrAN+NvMC9Ddh8iCZld26T0cHtTvK3pRfOXR8DLajf46tUreJ+HtfU0Vns1bIyD
0tcgPAm0Skw90mRZdBDFyYjSOmfcPZuSoOgs8IEcfMVxL0hBHoEwLjd4guwMwjrnMcfhHyrc5zUr
tzwUiMiw04mHxefZWXgoaLKeYhf9o5zriKPPvRuY4B2AcFTKhBkCGlz9FMtlMLi3P/5bEBTxoqfI
E/vfKfvf6ngUCOZF5bYFoqS7ePJjTU9Yysj2s0QFay9wHiLHRxoHcsNNOxNSnVulGfEhoTLI3uB4
kDDx+4NnYtlUx7FgpJ9SLy6Als6WV1+5n7Bhd1l4jeBKqtfLdi1BcPWtsln6m0ia3rxtxSAfs4dj
XGUUbnSKfYRWm+8wqfVeKOBQeIqb/ie8kJrhte+4s8ayprnicVHTy+EYlKTVkRC/YLpJhrOcOFs7
2uB6B3KHOhyFczu3LxjykF0hiOWfaQZ4twFNxRjXZgrCbNBYR+R6o7A7qwdKJlqQW5ZUHryvQxnz
GaRvNYKpiRpn7rt29Af92LzlvC+HAth8DiUjr130+4TVPhmDM5DMXinzudTPxibL+lLeNZMFfZET
ajlb2u3bo0IG3wPDYiYabEjh8cbwyldG4v6CxPohYc9r+P0212Wt32e5Tp8TUYFJNLmovf+l8lbw
RKKrOwZ4hRtcTflZiJsVjh6NPJijr3oAA5Y5lW5v10/+YUbtiyI2tIx1U5oA/WfOPptWBzSgFCYK
t6xi8/r6PbubXMYMyz9YkPAqjkf9tPM3/Y0frTsWqol3mOEo05AADQdnmIEmvtMwzvC7WHs1K3zq
5q6nq4FVLnGPXnWmRdYSCbRdE3xUW9zQK/z+TLN/4+O4gENlrQT7LPLAY5PzTqOGXsYvy5dAhmiA
abumINiY9A/CXxGDjIwEyow9BKJmdbRuV4j3e4mch7qcCQFtyaSV02MvzLKh8R5GC4qjoLazoCqQ
9sUwKvu1/zx7cjdeKIlOC6zthZgstRqza1+T02k5KKUjSTDfAMz5NhW92GMm+kIJt2lxIPaeRgNx
5yCRPMS8oeGNfUKUWITqEmJK26hMUTwDNFXIGaNwUo6uiUdCalOdQwIHGfJ/N2d7MwUBJ/lgE5W8
59WO4L/OJ+63adqiGz9MUjTnxVF6t7QICHWHI8juaPBBqzj0IONk5wqHfIVxnwL3yWXixy1IvtQt
vyO7thufWBZE3knycKME1qSAGOWQN1OTtlgExmnomWd5k60UOND04tttNCsZKPFrYWvB8l2IYXwI
FvQjMmKp72K7IzByjcQQRTh7wl9s+KuxXuA5ivnuGvFcvZQHLsUchkkBT8tqqzaA5V4pfBOfpMhf
ryBmg1doFjOP2NHrIx0XeWBUljzQ3xKdgegXQXS8UUf0CgrbUlh1f0pzkFAq9FVLPRTrF75GkA3t
q4VVoqdo7EIwAQKmXpU23peCbIf2putfVLciU9F63PJJ7IiC52ebAyaOKAXvbM5krqCda8F4wpib
O+nJLN5p9phpcxmaiGLDjgnozUtGl3Nkn8btFScwDrkEN+tvi61j3BPPOiTD8N7Q8hNN4C6xNS7u
0m+4aPF0s80hXH6Q9mVq7wVBnWjhA79ilHzSblY68f3ScZjnsBC481U4RkHFquXCrsHpOoL5g84Z
tUfYDTJjpo9Gsyonb9ewDUTvtmTmptSwtJpe11w5FWRFaS/+Y5kggVqNZh9+8HisJ6SbqnhnPlar
FzAxgyGOSLSLmIAaQYG7nfM9wjEhKMVwN6kRS7gg38WSf0PEdTCmgDTKmuhygNPn3WHgCvkVgnOQ
7UsujUJhV+1ZSEbahaHIQxtPrKOwLDAIPP2Kz22Y3DWmFk8Q1G3WDQe5OJe63u5Dq10/NofkEFI5
mSRfVaYL6EwBZcb4gcuq0z13UfMxSalXZXQOKIm0+qFq2H+/IA9qczHjqxH6GfAUCOqUX56rCJXt
hCT97/xBDQ5R85KYOwkpZRdbwqN/C6MquxzKNkm4T2gHfIwXwYX5JtJC+hX9mOj2SHlviWI8lFrd
wNAG/AAspfHvDmlOVfUmpZIC+6/9fNRP9vLcynMbIRkAzhAMdI8IW+ElyLvY+xRlJGzR22txJHQH
zi+PNqF468Zjx5r6cVNt6VrbvEDsWFbREsb5AaqRfaVkio8TdsD9WXVud3z75OJBn+zYCY2pWHV1
LpQ7EUS9kEwauLxnjD61Iu35OC+mntZlVZhENzzpIbgwzJ3CzJK46CeXPIYl43tkJ5jLllPQAbw7
ae/aBaeKaYavW1DnebH5HZ7tvKsl68Exvhcr4K0VE8LMQR1Ylq45LuIryZVRUBM9xvYNbCxNs/Xm
oH3T8fZjSQ7qHfJf2djUFKXJbFhQcREkKOXvSEhD53ZBGK19LLPcLiUwuwabmkF26O2DHtcj63jQ
j9QFnB9gg6fbCgKcT+K0MFPTql9W9f5VhATaSjT/v0cDYzaWnPosEHFXuvXt6N0lt3uldTzJfIKM
IFRddu9N2udWB5XbQPKZY1J1lhbJpD/1PRh1SIeLIzramqpm7hxf2WnpGCqcJ28opeDHUUutM5Ak
qI4ppdbAGlclm6ZWBhW6tkWB07Cix8uxFzllOy8eH74NXAAR6rXT5lvgWPd96PiaQ0w1VPWjU9QY
j1xBfYXnNmapgp2Nrk1WDEy55o4FQ6qPgZEAEMzo1Khc3A6cgmPPoRXn8J2P9+DsTwonFtshk7z8
xeVCMtUL0mHb75ViH5NnFycVdXxoLhEsy7KbyQYzl3RWwlXm7LvUfhn2JaHidLqtaB2ADQpgO4HN
YdGSkGDC37vZaY1wqR9XUBwZZIfES0AdTC27CUMNzThnbiE4G3fWz3kNIg5kiY5PjmykEHXnoe3C
rRbkKq/c31r9wF8lHlbsOZaipex8iql+wDX/REF33ODc1zHP7+9H1iDm5S1W22nPdzLIOuoN0YY3
bIACrPonrZMtES2CUEdO5nX579JqA2aF06h3eucN+PxEbSUrdA/ztAN3k3FxK2mpiKDGstE1djZ5
KpZ7XDaXQ//JxeG2OYTQYwaoNj3f+4Ake3nQFHtXL2TpHlXFwQlCFB5Nb85S+oXKKmIju4Gpyumm
iwM4en8PfE0dnguYAfrQkPWLBHXIrfXqKkfXIHayZO9P0haEQeO4JRLbkYrzDiktKOtk7S0qh35H
wTuH/Wk52QOv4h6BAA9gwDcM+6Cl4RL0cy1qUnCaMqjB14MuNDbcjCQKAzkqusiJPlIEPfCZd9BR
rzLYmj/V6HTVI1saDVosUNT4H4hm/39G5IrqLQ+QHv8sStH2mhf132UhC25r8DgZWEZWtxINofaT
2oLIwao1xNLBL4sprKPt0R4TUhu3VpfbeExM6dXUC1nykIpb2/B5J9PCCtsvYK7bOwwVVn3GOCul
vP7Pe5TOubdH2AgQZERDDocRLw+iZylUOzWFGmJbUGS6X8lXThGoUosmBwRQYoqiNB+c4e7YdLEE
F1f3eXav2H6nHIDg6lpA+02z5UHF+i5AdFfjQWOglBcmTjq6I5HC49Rri+qwhhEpKljh4WO1OiZI
YbgOViGWrYWhvZ0nrpSqwacIiqDzVDG4h3FXy9AqJNamvPs5fe/PoW2SVcnHHkfgV0RwOjNrgVBw
T86JHhM9yzZZiMA8sv29qQqridsOJQVavBoqvrSLmOtRPc8nuA8CM9uSNIu+p3VZdGFSx0Gd7TRj
2kmb23lTf/HKTw0Z8MXJW0j15gE4bC77uZQTXYhhLoO02GpC9dHo2kUmCKghl0gpxlDolwO91jVs
vRyJPpQRkoxZG30SASgA02ZWaZ+q2bZmhSKZO0iFtGHdU2mvf1AUyf8ZX9MJ2G5o6w/TOM9UTaVR
+eAoXwpOnLzCoBoZQESgbnwzpu3r3hRAehUqVL57tfI9tVUSyC0i9P4hvKbBmyHwkgaRC3n8HrnF
F05WSMosNjxZrEmh1qmWfpVITicv4ikrAXtMoIKZnnM7panXf7kmkzdmjVTMDpg0jRsdVMlFdu6d
+tcs5qdx1clZyvQZcK8/QWrfZ29Zr58zILIUp/toSUTBvA5PVhHOnFFyGf2YDM01O8oGZi8WWm4Q
YCr/NElXlKdWlJKF+oQY4Q6D4xxjBcrN7iwSPuhAJNcJzs3AEV7SmtXhzu0eSbTOW2oWaGAq7GFZ
Vibihqn6a3Ug8ymUsgMx0my6/gIzi59H+PvvD3QlZK+ktxQPyRRmR3Cqp1joFw5NpGE5qsl68s10
xwpYUhKSAXKQAvyVS3HAp1J2rmWF9A6488X8q31vvKtYB6ZKA2Xq+vGgomDsHaMbp2skKnMv3iEb
lx1Rx2UwVulvyNrO7qX7XfMWcguOjlGPfb+9d1ctZb3gSS5IjUMQ/ouC3lFNT2JoqvGemFfh7WB0
AQv1t+OlhQvh9FPVTsv69DKcHIzhlBKfsK+k3gQdYVBebSqbw8d8iysie4g6RhGHpHGm0/nnDFhT
xHZXjTQ9kyrJ7SlZgHLMlNM7lZJ/Bcm9jm1jkFGpZXiE5HLRLF858YbA70w+d+4XsJHf05bRi7Xl
WwEIYOukwsXxn+L1+ja9zMXVqwYo3ha4ZXIFC+Zv8l59eIeO3t7IpDn6wF9IiClt+WfzusgQqN0w
osqc9oea+116ErDBSUCssXvHBIvXTHsdKgJ3OgENxRJeW9HnL8roqt75g4ZSNYtOa1lmHvgqBtlY
h9JQ0kvcqj9zGwHpujSmH21aFSeyh4yIlatlrwD4X5P/x32OG4ewW8e6YI7Zot7QzahFO3tN8kpD
ozcXgmeJW/2bmOnCMeFMHDm2bTyIEDzwNe8+TNOdb4r+va/0Q1PS8srP9wZl8fvEKvg8noxtt+YN
ECRanN4Newhqq0iP+uCveMTpO+DzU62SUCKP1OkcvaOaJPf0XmrGFUWGJPFGz3xHqnD0izfYTEoS
vazQaRywtUPXkYmRaVo00X0ZzeW1RCaOALa9475qOR1YFhx4T45JzZkcR8Xq46eMt1JO1X5SFwHf
WfczktTsdTT/UrrchJDIH4tdA1itXbAwIINWhIiJ7jX7AwcKENrPNEpvsw67iUob7az/wkkHELAS
vG5jdI4nCYSsXNhJggOB3jLIOFNvesTuLVUFWtRvmAOqZAmeM1/b123H4BRMZssKR/wBf2psrnO7
yfoSvnYvy/pne3IRzOhDG5yye9N181scibtR8iDM7dI/U95yEbzZDgx2RAevFdJTqTlcl/f9hG1U
QtB2puxAa+gVXt1WbOB56M1WvwLqTyK1gVazIpE/GKn9BY8ouOj33CEEs3bDkbFFDh9ofgZioRZp
a9wjyETbqHjL4N6XsokjBWjo0Mcn64q35cDnXAD0UdA672Lm8Y/URhqlUUI1jUxUVVEGFrQ/B2xa
5JHRJQw4A1q2ZTxU2eRXafwWnYx375iyUvMN4Z7A3Rw1BzILRRGZCOd2D2Gn9dF+uJ3kDekflBQc
iOwOyyVpKGEPsd2nsBNeka4yxF9OaW2u4nroQCu53KoZJmDWDixwblAG9M58ZjyQGAANUHZtgJdD
ZPO2UultcgIS9YkDZhnsmU9iHtIuqktYgnhmL2EQn3T5WO5+zcwKRwZW6s4/6wc7IEUyP32ubKJb
6ZSRY46Dh8fmBbz6bBcW0qn8YBAONuJIz+QEcRInGJPnO127ol1EXgZsqLX0gKu4f4bf8z9j+VWK
D16fYoQ0oyfQ1pRDxW3uFYPDIqxOepr0WaM5fot80yvUJDi/pvBnM2fvAgDL5kYBmMWp4l5KzgNK
JJcR493lCac7RJi3YG8Zf5krvDk2xJxv7mqdi6N9wm27opwT60jNX+N40D/wNsfHEAvq04ZNt3Kd
iMfYnC4GJi+yc3MEJIltxYRQi95Uj/tcVQa1kxTK/0tPaDbjufmyL8K11wd3mqpKv6lGgYT515bY
iyoKio8YKV4H4JAlTpvI8knFuiv2qrDz9yzVpnz2uJ1ihqW6pujiOQGkn9V7wFF9fUWCd4ZafCNB
q3NqM3UhCvdi5k2/ADdVj5RmrVtapMDdZOY8SUd8AiVEieC7NJYFuDzOcIqz52VnoVJwqiXr/f+/
dg0FcMlZ5gEmd9jTSGEQ2G+PJqjOJrbiwjYeHbfJ3WOB9/S7O7fdkE5zCFIBQSAJD00n60rb0rMu
UDaShkV+bciXYuQkJmTNQDdPxkTYPhOw22VGDlfNTT9dt9doORLt2jpnsF6f9m+ZC37xvlpQVgZY
t6kFP1YZDgaJljOOvA/HVZfS+JzLce27Np0TsSLuAkZ/iRi5+LtUsPKlrEs7HvBtDu/1T++EA51b
jC2s/5kQPT7n2xWyZbkT9TvMY4FZUPqAy9rqJzYLTSqtF6wUi80WV8SE3zFTdHTh9fMZ6/sB24FY
FfV8B0abP9NWfJZ0oEWx9WYgRAJpyUZvSruEQ2lOpEL42Of5oo1OPjjV2RUENiaZSN7vsKw34t2n
jrmz/ahqYk3AIAF4J3eNlgjvgT/EFArr8KMamaO6neIACwGeeXp8uyIMuFTWPD2PnEHpRC/+ue7G
BUwsxKlirBFEQUGGBdzQYvgxwzF+98S6GrH75rOW7At7FqvdkGjcv2Jd6jubFYx/gCRGnHOjY8Vl
QIhgj/ifmRXQC7ZdHaMrbwPWkU/ljIcVfnAFJhvojbmHy0bopHzlxKi7FU0llrYksZXGU7/gunrk
TKHfN3GmDlA0Cq4/2Ef2jlKLQUCwebWQeh0k7u2WNUOsL3NAaxjt+TbUsLNcobhQfnJiQ42YYw7v
Ei/gDr3WzEleD7a6sbzv432P/uMyrrmBFHJSpLIFmrd6u8lfMpLehc8VPfOE/MchgBB24sDUfnaD
CtvordJhn36xb/B/REjAIV0zOVmTr2nfry+gFIF/ZyJ4XzxfGiWF14bHpXly1LbFLjC3N9KDxXsq
DooVf8qrN2+SeDEw198Bu0J45G4XHkr+FdIimTu8IBfk68ahz2N9nSnQTEaPBIxFM9Gxr6BD/Oso
SVuJV23nC3Jmq5Tw24OVdTP06VOnVKWCY5Reob8CRq6Zh7DlOM1W2NQGyYuufh5CDftUvE8hd60p
u6Bo/xHt1AHHkgkrHppKayJQnDleykgp/91qZhbW6at/5RROLjhuaEDZ/sqdPvu4MhCM1H3L4g+f
ilhSYlxaHzN7Vs+U30Ob8PdVP3GQlArc4Ady6BkHR6ss4EFPsh/Ml3StXJJQd5EXPtndVv2a0aCa
kjJU9h9ooMF2i0EUGXVSz15jeEXrsR/1oydudelBEgaGWy3ZRq9/yDkU8p/vayVqxtJYnHGLfHiw
W0C1Tjd3pbmAFY0pz8760NXz7u1KZJwSKj0PC8PHltYOt8SVQ/tyAj4kdq3wme2Hfnn3hJaYVcNG
VbMDO6aYjSKxgMgHSSppaL1LLqMRf/6oSvSCEmEhvp867uAea/fW2qL/7ht6Ma1ZjbIKrDtg4GjF
DLRnyKPoH8t0YwYToMlEmnt4VC9EmvYzYyu8FQetjMv4pY1UcO6pwcNSKDUHndTxaFeqFgRGKz0t
9TlfPcAJ4U97j64ehHT29LgMDJQ40IKx2tJcrfAx0qlbx8DTajw9rv6Ls/CFrrSKYQYkUMZjIYpf
2IyWmQdVO19fqN2/s3y34NEtynEcGH4KWlPT+LnEzLa/+J0XlpeojFqrHU3ZR9QH1q0LBtFCnN3P
meia4K121dgIWUzoDq5QeEtauYjYrkNCggXWBpR9IgpSv5FSnpW9nGKYWiQTj3IyvcwwqS/Gja44
RhbKTQGQY37CD1MEUka8qKXufNJsQEFEc8aIOPO7BQi+qIA/xAIyfmQgYpQI71vbIIHPkswtm5vg
pUmtYI4P7mrmO9uvPhFsL1GbT+Qgjs3RgdmJPEGrVw7zyekCi0y6kBhV26PitUmSDEQT3HZhKEhX
gc/HMs+ixNevppw8MUUkDGHb80fbZ573tvRcE5MEhpaeJUxCzE4XwtCB0kFbdyXBp3C6LzBNAHQ4
SbdY+U+VBHoycnj6eFG6x0bTYZK8QCIqxsA0/ZYpgqvehAorwhD1sHBEBjyJjRKblHozjUxx0h7G
LcHXctTJH8QYy5lzDfmthMSqkr6AuGYFWnQuy/p4fXhu+Z75hU7RiYW+s1g4tdt75hS1nyZh/VCH
sihIC0TcVn31WnBBxxOdLG5E8Ag9o6axLS+ZpJH+MnsVUyTedE7rekO28Qql2Rvxz1Zt+4eAa5GD
Rj3470IevRfPQYmE5kzEMVh+yZ6q0gfnAG5+IbqsBGRz8HsDvLUtzpJlRJdT2ckPTGQZSyG4Ossf
dh6ZEPcMr8hX7tgiTNvUqGyQYS0N6DaJDxUIezPQm88FsGs2W0SmjN9fHZmgynP4HmNTJU+rkY7x
tlJ2zWEfD/dFaR0CoGBDz8dRYudkfRrE0Ee3AC7Tpg3SHSxIlR0hkWYShellYD9UeAaQsLQhoggg
xFvJQi8iT4JimkX8vQDRx4w/KZt8yAcIFG9tK00v+wSt6zqLhCH7EdsWwwovvvwYlEPk8gC5j+x2
rbblk8UwjYyR9JR2F1JBtTGm3jLt3hRD/Jn7DJNGUk9NObMsqPoRcwC8sCUngowJzKJnU71D+2xk
mT11egIqXg3NwlsUSMSZ1flTK/aI+3Vywd2FBxFu/1vdDUL3jRIhtnA6eQgm/vaDchlfMupDtAZh
NLj4ULzK3vRmoN794pxxf1jXYGRGhlh39a2Qd5jRrDWSIOqiuqCBH2LgoNYhMe23bSpDHHVCDDt+
fbSVbfa9odWYgYIcds2FwDwcEkVjUQ3J3V4yQeR3sg1NK9qwob2xbiBqLTtjtM1XI83wBv+KLb+V
wJyDIQ8OOFRGo/Wpvi/compshwWTCXuyLM6AC+jKNVKR+2FL9LfVh+0LpD3a9dk3xPl9+JBdJiYl
I8pf1J59dRyXJPq67wkY7Webb3zh+UcIqsnlo7PMAhvvByeH6VtgpOtq4QalUevAPuicWz3IuiVn
Y0MusEQhnzUA0I0wPWcfyneBnUgX/bRPU5HODur1llKjXt/p56EgslELVza+qOWMOnSmm9reD25V
l+E1ezvvD1Czt5KETEV4xjVSiat2I71wiPwW/xfBceRBrBgtvtvJXhSkfOS//MZE0R1IPu1iJPe2
vnuzd6ZAhUZxzr3hMNjvm6qwExZO97yn351FqD6AJ4taaTkv7TSnOq6/VrPHeZGe0tgjlkC/k2qk
U0Uflk1HsEqnG490fZ2amzj1XEQ5ysa4Ol7W6ADO+s28wY0Geq8g1armqzLd72LHm2pELeC+iJgx
iEo83N/JM5OqUeUiclpmMHD2e7yYxcTPYlRq8Wa2BX+6AFR3KarP23VKpUdrCuZO6UecLpO/fTXX
RohwEC9+x1JC85+HokoNQOQeuXZ8XaLRT/PQHIHJ0jmuIhQdYz6QgLRrHaU6T2jVaNQo1zM+Kl1N
A3xg1Z0ioWF3PzPaltm4tYBuoQhTZXXUZgWZDT72kIiqxDUzfeHhCjybw4Hb7n8dzmGXdY63F0Fh
uodgeM5Ls/fZsmA9qB+rdPCM1wJiciUGKCR2JFVm/2DHB1FnjG0dalTylpwzt7RhIIkoPDxDQHui
s6uaMsjzczhL6RTa4rMvl4+xdeUtZUl90u+YaKoQyRBD9h68JDTY/EkU7xCTYI6JsDVcfvkb+TUc
qkxVSUsiVw5DWySUz6o3JHkJCl1LY7Cd+Hd4aXp/+on/tSS5e1Gt+TbhUYx30Rat/kkhdKNEPbb+
38ba4ItoVoxuLQtMKmNy4mTJr9hutGbFLES0Kh8qPYKB9EAQShFmb5ocP2eY12vtYSo23qBv3iV4
C7PCc1lpgiFfhiWekJ4qkHQ0g1XrqisL5LrTaVW5PsvdxTcGC6k8AqKKV1UWDlVeLlHcKBoGC7dk
OtTtMxVNU0cdbRmrScb3YbT7iiVNq4inyNnVAUqvcxni288n9uK36YsISwW+xXr5mVfVHlwUIaM6
QVe3nrvAzCj0TMaWl2V3rIIAGM149MC0XN8gDXQICkBohwz/bFSnerApJMjiC7WkT1JFW5oqxsDD
bB8PEUxMDYyR36ZCNhIC+3cHTgqdruGirSuU54H1HeiEIECNPKQJcy4MoBQZMQlJZ4x/h9RIOspq
Id0XvbDeUYtRHEhV5IL8ja2Qk7PYVa+2vTIuOpFqcEBC9scRhbItDcbfUYJVCzThygiMBjVaI/Ly
XSBeCf3NVsv/md3fSmE8lOiAgqbZJDYDWzpk9a+zuUOHSu7/86PatSkLE4fLMWGt1OuOdAEvoA8N
NKve65Nip3MIO6Dee6GegSJPQbN6/XQkgBEoYO+T3RydaJf/FMv/LGlTsktYmCv1QIG58o18sFLp
TDvQ9AR+I5I5Ub88wzNl6QiT/fAth03DDFr5NPw2CQzjutsLNRa12xzakOmkueouAZEy4IHj3CAp
XCvpDOGv3jGgb8F7ceVyzO9QLNhJ3Ubs/iwWZE6z5556m8Agf2WjCNHwoUC6CVcJj76LK/L52z20
hvbH49CL+pWrWb2tWFkyz0H3cwwEVpvDMqfDOyY9UDrIVgR85Gi8XAcuU2LWFwCVsdgQysvzeEZL
qBU53KaiQkUqpKGdWvpuomJZ4d/dWEXq9BVfmnG35RuCKUx0UPB8h4ulECDVzYBJZJ/FIUnjqKgS
TuF6fbuQr25FWl88Gt3/a4VvYrdTlmvoOmZD7kTpb+NfKV0JZrpNDjO5OlOTamApapGjsYwdC8Ds
d8Smd2r2ur8X42MYVvxQX0h1lS4/QMaM3aNOA4CiglV41eOkTqla2F5fIW4SEgZFT88jIZedCTgQ
ASLWER2coo9lbF/bYDglA+tmRznFMtYz6pQO+LTGOrhBh2bmFZuKBspog9CpMnfvk7xd1gGKByNz
VwanynlsTeTAAFXCsvwIcSBjsuz5kkjyW8FTwgHpjzaxRrYb/2K7Wrp7VWbzOtIJ0PtZQHvcOz8q
tD/vMS0hIPRRtLOVBP6SvsMT1raXNVrRyP1ssJfCHUjv6r3JtATQZq9ArcTXRtVwMsz8Gja6pFkM
Wb+UBwcfT5kg3zU7oqM2MM2Mb3tVhvOCxr/rNF+1TQlzmGMPCVtc5+42nus+MwjqWKoRT5kjcFXr
AldqQRSNbkQ5i7cGYhUYthSJ0vIE/T6UYBsYbSGj5KtHBwYkUEa/X9uSpslUAbaPKdttrrzmLDJh
15UgAVp6LhrKmTHihlnjthx5VJMICydJ1o2AN+KXosI/pOIP6okuagKoj30780Q6ykrQXGeoGLuN
0sohm48TqLpxh4Rhoz7In4NoOBX0TbJpEPzCIuXqAnpUX7a2Wfzdv6ob4Ix4xj9AT4+UjWkfOC8v
gEXyJjRXGao/krLbxsOj5rnAPaMfk6nwjvY/Es1bEg9XP7Ml0HZ86t85GDgo21WMQhBCJGIzMXmc
iaqw+gXvoz2d8nfu0Vr/0glrknHOvflYnoxRgbVa5ezkqER/AhR2RcAXpoB0qRajtWN03cONBXor
7BiZ5KCrC1YHRC3rT7CbWJrKLXf5FXCXlgqXUtngF4I2pbwpXnKtq/ZjAMuUZeVnLVVNrwdsm3KI
36yPXHw2qx2VrrWLmmfJeMcFh/Xg81h8S3+TA6+/oXiqWLC1gBVu8QsznHLKdKpt8M+uZQpR2f9r
KvkO5BhOqNkihrH6sYX9TdBG4AfPkYTZUA9rjpVfpS9jJbj0JPkW0UErAfCGSdAkE84aJhdjD3uO
3Q3q9Kg9VFtSqY4OaQ+VyVcpuh6u2NB3A52OJhoM7e4x87dK/LrSrZJDWv3mWvcRHLPUokNGGcpG
5VBRkBq77zpXHhJc0vq2E+YfxzIl3MqPSTXB8Ow7NxZzthJ700nrfp9j4b/Pvk6wPUm9l7p3+v5K
D7RwPGSW+wYJaqoAxXD/TBmadCcVhT6jFomJ4LUqX1XIJoqHe7Nre12UhshE9uONERVyYUe+YVUv
hA4xMCP4N69OSrvjHUlQEVaQZ2ZSuTQCAEaO5SthEhuWtsDBtmzt4ASFJCXxNW4ov8gBXRAhl7fA
+VPM4u7BhhF6GuFSNOx3eY1fefJEYkeFTRwkmwWbas1XCPYWnnaRTHwB8Ke0oSkmVx0L/uTbFgJw
0H4cHbKRbc4jPCkF6zXjtGY2VPRqbDNaTGLR9TU67kgiTlDi5oMaNAKm9ceHqOt8wepM+7F0sLS4
+zJmP2wexVaKBSm/tHJ+Pd1NMNZV6VJ74BzRKZsVktzk9AMLLltjHxXxzePS/GIDZ8vQmDG0itRa
5aD4GGw08Jzde+l+EIRLMnvUtzm+kDONkY5axFMeWTXHl1EbNiaSvJyzxbRZ6WeReZd5akrgyBye
ZzXbVuhQLElsKeeBVyL0L9FVQfAXWFAxUoN1MxnX2ioir4KaJWBOKRtbTZHstTCs4WkPr7ZHI5sZ
ephoBAtcyZ/q3El5yPAW8RMhAsI3qLp/A/gjFfOtWwE9fRGji/LVeyqLklGk2szRu+BEgk/5+NTs
HInzApcZSpX5lwvJz9MpxTpAWSm2LsKISBGCpeuXVkNkdmcE/O5pZPNnO4stfouDI7719Dme3h5R
OxtS4sNdDW2acOMQVsxXSOaguB5v7Guji12HGLwE/u2M4CqUBdLGZCCOlCLfR62hhS9Y53RHTUUP
CytQO5tSJ8VtwqihO6Mka444hCbc3/HypnXrNHvgKAf57U0rlsTmRMha4tDEWL1kbBa0jiTmNTLU
rjr/qOpsJ1oOuDgWvgUOaSfRAoENTi7zk/0v3nGuFTx85kspd+YeiILhbKy3RI1a5/+KCIQ/e6mg
5BOvAPwM+OZSneL5kBOFKDTjU1GC71/AQWdLbp5AUu81x+Kv2NEyGHZra+GtUd4A97dPD0bLRNx3
on3gjYYeVoQt258Tzi3YF1O+N/WDBylLgfQTIRlneA85v9bOfh+/5410K9DhFZVY10gRt4c7W23t
Q0vdAlRTFxYNm8HZfhLm9rRqTRuxm2b1hMCF3CmhTbj8+akc7YFj1oWNemXs8TiTN5k/4FYU62hI
xvRyog64yE5v9b2EVf1rQgC2Ezoks+59bzc7llMdyP73o1Aft9m+aLq21IQgQEDuYs4WE7wXa8+3
hj4vZ/cAyj/J/QFHyQD0vW7C4viITDJpoyaMiECATTW/GEusc/SJOgYH+E5imvqYnB+DNCfsY3ja
GG2jY4jj7iTV38YFRYP9EEpJRdUO/qZTpX+eHd2r7+H1ERQ+AC+sgWlRMYOgFArz1k9dA6z3OAEk
EdE4d00AgF/UiJc1lDkz1luFopvspJKWAlXuyxKM3ZWtwzy17pIrjos6fQcsrpFHEhNb2Hm37U3N
kjopfsBx69bYo8fiBeodGOIs2yjDNb6ujvX6qD0qK/4HfaihuOTgydBMpfPVI3U/7+Hv+y1LbzpG
vLFajKWcNjQXTSu0dOIV919TJJNFmMqIMTxaKMVxPCUqKNFPiMPFgSPGCoTiLyiEgJ+4bxnj2Cdh
z5F9wFb5NmpAJhixMk4q+CXjsWt7cjwTEh8ZTYqPiqa9nOEr2nAMYurMJc3OseRkqmsG5U/ugO9F
46fR5hs0EVQhaez1+UTdTQRFk57cTqKj7GJxMOj0tYWpxPYNgBPkmxc0qRpWVqqj9dEQgod1vN63
ZMSqBvVW9NIrEdzWvCQwJXnFGHUzUHxoMWBOR8leSO5KEuCV5ZAOTOiP0RVFY42r/eJZd6KLxhD3
HR6cYTgq2SJjiE4+uGKBAUUbKbaTdncQCm+9aWPQqjhYFnr4AGDfcFdCDYUVTd3AUCYb1LB91LA0
yMp4zkqOb663WPehd81/bMDrJ4zLRM5YIQ49TdehfuDCCq3Mf/zf60RHFGKZe0leH/cZlPX30wN8
w0JsAuhzZpx6zIH5/uq7vd7GB3xM5nH7tvlqCisCtoGIf/zsFzy/+CSxF4Gb3nTUIT8/1TYnbXLk
Ojd0T8RR1w2qvz2F38yoPfqfJKLtjufSjTRqqqVU4DGzxp4IOAH6o8I1MDlc0fkWhkACFo8O5jKk
SiVsFfH4k47Vc1MF+z7fReIqNJhxpOtgFXy/pVxJKlKHJnjjOZW4wtNOnl8zf5o30zAyw4JlbA5p
MWSH7gXbTnUe0lh+WCGxMw0X+yqd/hGR754O2f2qtTtcasJuqjbbnNXgfLFClF0oBoUrE/lVfJv4
G2yi0Gq8cy2Uls7kSwCIOaMGFo7lIcWZbnXknAnNc8lABbOGbSZP3kYJVm8EyyKnyhxsyLekauPl
1PtzNEZ/BCFlV5hXZ3SUM5daIhfRFgP6++gO73JlT/0Tcq7r4X08To4f3lUWDTyjgg8/Y2whlr8m
zjOu8arJq8vzaRL9aT4AaXRIB/aRE7+D2mLdiPRUjwZT+EQM6FasKFW91NzpFyvQchAsVAL3YlDO
BjwiRh83t+5Wxzi3L8iGvJgtojLjU7gywy2Gh1JPzZayHBIJtti+Jz+92O1q1PM8uzyXNmICPC5Z
NDYOCvqltefAa4rEVYiN4iVQtGZyP6T3kgV7zfeJJ81R7cg/IOZNxAqrXvEayjWyL5BPRN75lQWZ
0rMSBX7NmwF1E6yVeqZrdYA4c0OB2islmF3zQdAonVwmJSBmMAl89/oVkZFevxPL7tOy1NzhbOdN
WnAlHHeNokTsaTb4pydyptQmHbBIaWeKboK7BgpqZRhar/NBQEDaaCNQAjJgu0HOMvD/IjTpQuJm
rGFRobjI0AlKh5l1ttrnltCHgBviiOJC2h/z7mElPKRBaBPefBaKPRqc7gjlLDfvCB2PV0+Jv+LK
A0wRIQc8KiHy/ChKG/KJHmKmT48Gx6cHa2T3lj1DNxME+WLeHqXe503doQz6cjtUXZCxprNVoadq
r5g6ick4KaKY9+xwzf0HM/5UvlOmP1aoZkC15jvDWMwFfY2xYe5VJXcE9timTkHWwvLQ2WsFhv++
eaQPhFm0OHfTDUj7mR7W3mGxRr1RV0x9uLJHLh8DTn1cziaB60R85PJgr2w7F0bAR1+QyJSW/kQX
lUglP3B9yfQugQZBL9vvJ4RkgpaE00K1wgb4qAsnS9zYiiW5LVDPANPRDWuXgonFYUimlb2mEnPe
0uUeJ2UzEHkxUOFXrf302zBNjLYFHnNS4JFc9QVC3RxLaD5dl7CX1Avmrrb+fXhazqWCvt6K+uAG
59m6aM7meUF7KwGR9sE0MD87+oF09fsOATUnQAwgDe9V01P+yLMAOtHAF5j38doegfqXVPhEyqA1
rVjaa8We5Ezv3iNo+b2v6b9iQtpBzqnKQr1ECEsf98w46FOhetwLolKWK3s3FDz5YlAWnYPREVVi
l/XzPbpCB5tkBsmz0742H2SYINd0imCe+TvVShoZpl+jYYnhbUeUlWyReIspC2q9g9IpD+7BorNk
/pP1tzC5o7BfO5lzQDdZuhMuRTVnvHKUJP2xzaNYh2QNK3hdv+TC3x0/CCFkDp4gFSGHzwNQbJH0
2cqUW0bJc0v1pMuTMikFW2G8NSiyFw5Q7b57dY+d9znFGdPE+b1D9gVZSJ3mD1yf5nm78Tv+cyAL
nDvSqUOB829hIJj9XUFBjWtZtDiJiofLUgTKlsMuTw9mxoO4xMbS5cTqsHEIcrC25yGemtt3IgaA
Ech2pskj0RdfZCKoTne84brT6YolCnJjXOTUJSbnIcFV/wiuooap3GO0qEO8zJH36MVM4VolNucO
Q6l4/3E1mYALDnsALk8NQYceu/gHZI8DxzCJBv4c9MxGYXBH8zDvHA1Ygpw3ZbGGs3eAA6E36Uqp
rJlXAuAv6/Tqz6/G1pHsyQaFLwpGgUtJd91i0JVhGP3FZZQtf0YX5MZAdb3HXjnehFMlnOcirnfg
i+0mLrNismuPnYwr4zjKEbZes1W8f4mgN4tP8Z1IR2T+/GJY46ySpNlMAaU5c4sQ79k32FoXGZay
zYrzVjzz9WKLW1R9yoxb0vSFclVXFaAVlgSlNUyYArvhHd33i8wQaHP8vOityUv8PXzpcPrQYNYP
rZb44omWQHIpBHrng5iCjHKU2sLPcSC2pGWZhYTDbf8ZdjKBrv9znuAEWSkE6M9HpnHr9OkWAYyg
c3zmOv+OAcn6F+yAewFwg+h/Toel9fySKzcQDGB+r8tB5Np21gnl0I/4spxr2JF/vCYlHzH6VEO1
7TyX3tA7IiEXfrafMQcKYVRD/7xVfAiK0M2wUKfKpXxKaKXYsIZCo07VKrayN89LoN/xFNtqV/ky
eRsQAtCfaMHUnI2nk+2zE0RWEACHJfV1fal5i8JZBfsJ1JLdWtlCUoCjJxBa+zk4xlA73As2SLIk
ic8gjIb93xK3jKR9Dr5O+XrUQU926yHBHBlG9MudEFcfj41nyrOZpMA72c9JBNhjJ18SPWBLHO5U
qm1vMDpWLA2LhLiw9xVzRRYtNQbxs7vYaPk4sJfLX4r690gz1CsnEaPUqK4ApwRzRFRk9AMBM4ae
DqcdyUqfnF9OCDdOKz52uIfyOEbbB9AkNIjo9H7aBuekZOChW5o6ujpFomR4ayc5x7BdkWRUjczi
aYBMTm66ysaMAjQZ0TO8moN1HWi0mnyO4T9lqusu/DjYxdaUtkuGYGoBQMJTndkan8pUj+RsGu+X
uQRnWjnbQB351FinFjB7coNic2KwyB1/z6EWRuT7G236KpdalTkTH/2X2KuXsWUwQ7//Qq09+9HB
t67f/LFj70uvVbv8hDPmK4V/C6XvJJ8vxYswFjkfYfIA9a57Tmd/NBcoNBGN4HradMIOwZGW3Uns
8wy5SqnY0fx7r/VcBaLtf1r0G+sp9B1xqiGpdLwCnkZiOuMtQp526vG8M/R4l/4B/Zb3KRakf07t
kitDVPYSy/+qwab5th0Psf4AFT9N+jKhMJHBXqX/03padIWVcBK50K2Whrl8PGEUllgQuONdYLDg
ouvp/4ONtRT9S/ciTQVGB5SzIF5qQ5d4RfaR0rdG1xvqV8lTmd8gorcXMF7dTA/eALKTMYKu4sG/
rHjcSmUWfchR0EzMuMRbYVMQC+cZ/OsIMMcyC+/VyFWQHnxDDr5PSob7mg47rDVUmsGDGvDf9xZX
SAZ1A+MyuZdlkrWppSC3bXJCEc3Wmj6SaA/cj1A3qOx4OFX0rNk/BhlskAEG9I6YJXPLR+hjA6/+
L8qY3ipTI2notL+lPlzCAaYEywtGugP+jYMY0HGFtQEYSZB4qnynElpRQRPxuTxV5KJxrbesGXNJ
sVxL7B3qUjC91pvRis4o9IFUC+y8yts4CYSYWAqDsZw+TPOGMa5cQTeSaX4obYFdssqv1+W8l6B9
ZeW2pBYkSXI26W91eqgXJO2kBBjFZjvXzqGOTyEsi3nmMfZ3EZPc4O5GuRZnnBzwQbeZMOwHZRGo
LbBgoJmC3UmfULVCV+n75ope5pRFGGm7txGolGOOcg4t+q7qlV84w0E9N1vq7hgAONTG/b9yhWjy
hGa0Bz3aItisDSA2Xr+O6QDH6HNk+U6ye4EkLm7EP4LQXCfSw+0YWjW972G4jCi/hl9td/Q2x/uK
dGrXyyNfAh0et6Qbvx7ssmXdHQowxdDleku6kaGxThIIgtAGdQDRa8rFTwnnaO9DFyBNNjeoN9AB
LQC/1dN7MVGS9sEArWQ6QAP6sMg3+w+vDho8ZpzQ/u0Qug/3ibzHqWiOq7lLF4zeh2Wycu4xA49n
OylPtJLsWFsdMd5Pvw76ve25cSi7lSSY8xapwFdAcR7V66Aw8mCToypzyHMwji2M4k9/kvhju0xD
1mHL3g5WQDksxL0IUYqx60nCyqOBwaKsJlhxrfDqNLq+uc0BN1qzP6/nwTYvFfBc4KWvX2p2yLcM
Xl0Y2n9ErPa9IR/hy6h6OO8L4qRDYjYMgPkKcPX4+21qkXFvaim7PPCwtCIB9Jlab1d+/eHvZtpp
/kJ6ntS6cgmKOKxh33DtCUg9046gzRwJ1ypeaIUjNEKpgMLpjN4ibrEIvE1rOQUtuvleV/1jWiJy
j0OcJ77gF4WiZWybol+qrVeUPvbrlkSDyBWi3TxHQNHnuGYLCX4YoxNO4soIuMt5E/AaSus37RKn
OI5BGoQAoCX0Qh+H0kvLSAkZet7gbPgeLhtR1p2tSXYoaVf3v5DHEzR5iOFOYZ4ZO3RGSTVyrRVg
YBIV8r5IJ1g/6QhiaXHNXmyeMIm+xvw7hsbgP/Yo23Vev9xQIMrXLOTvpO0nVpRgcPID+MKxgl2x
5EyZAUQ71DNlQRuT5R6ixQ3g2BcoAfwuibZ9AbNgIlXgToeVfE2Zv6t9Xu/cZFGurULXXU0jKNAM
h2ONK9l79QBAsYR10N/fJ3dcqoAepeF75pS+xoCrTFJBlGKfiLG4IRELsgw/Gy8ldxnTv+URX2YG
WTMxhC95BXlF8d7ygo99geuxLBriEbSWm91Er3Y/9/DVZP5yQJGGJ/4CJciaXTbuk4ZXWeSkM9OZ
+4Hs07T8epunD/6tYlXe6rKKTcYhZ1LbDBtd4VvC3gULOvYm8FA3G0bBAwAZS7Phpkp+dbgLLX2A
i+dNMbdo91ZGjA84eRc2a8YQlkk3zr0jT3Fh1FxyW+U80DBlTU6eF0s7vwPJnYFuyTzf2tyUj9Vx
S5/YmmhQSceszgzEFPATjLj5738ihIzr3UXNCcKUYmrRXn0MZSj2JcVr/vYbkNbOBKKoSfQ77p1C
CNAvrSkmUdI/HBcIKX0Tkc4eOBcc6U/13+eY8zlKcirVPNoNkAjZKcSA5WQOl6MNXkXihB0KM3PJ
Jsd2dHr26YD2Fm7T+nP2V6alPYPVMeX8/XLzkdg8OBICiAIf6BhMWSs8dx1442Ig3j3inHLeW3Io
ifiCKHR5ashHva0VTdVWv8Jtymsytt5BqdKwZdHlBnpU9T+JKx0e8PPiZ9sXPpsdWiDb4rmn+44I
DW/xKfoyqJh28HJGY37OCn88a3eoO605rMMYA6JcfqkPeAetJ61rIuQeVW/7FK3EyzMAJUw7K0L5
gHPdPPh/Tunx/O1KF80gfbPYBceGCKcG3DPaFteFk4P9DCWsRubh2VmZ+/vtIRhjz3Np6HoW+Ipr
EUnkLwa7wO96aB9XxybgM5c/9HSpNNAFqIa5wVQlHiKV5q9nZSvuPV0MBO8oKvwLuogkDK6ae2qv
YVkjGxboKdjW49ZSm5g4UI8i6b/+0KVrmr9Z4w9vh7kn3JeutJqNEtgRMwRYQ5xNYrk2cq4pK5nG
WOYTOC/4Xb96e8fvjulDv8ffGKuCTbAw7quizbcK/RZSR57WnGccgAq7PEycRL6sg18IPzkYks0R
iCFaIkRVH6iK6ZvOSHuS+gc/5HIjzSrlA5SU4eJmTr+qkzgz21ZHSguEGbjbh9Dfo2DZE37shgSF
yQEkhg8Pmd+6NaHCaUJcfXVW+vvRDllJjH6g9DhnkDCj9FKByvGyGyMKxSHw1fupWoYz1meD1MVL
f7HErUAWieQaD82p+6jWmK/dZ730PPkDSMoiBygzoZUGfVIT55KKD6uHcLPONkVm8ixCRgdKL1EO
ztxAADhMVyI2g5SFx170KWhsZgXiqmCzCSd3rSJRZrcGaWaob4m7CtL1gNwUU8sHAdvz/T/Oz4cj
4I+K7oThsUDd+BNSP1N5cvNfLyhyBsOBns0FJQL6Hw7CYZFWU6uz/DH2ap69HI+itRQA9QMjlLeO
eWZOAGq5lQQ3EJuyl7s2rbUkKQzzJKh7bfDOwuyNCYlhKwIgdr0oE68XgDVGgBDKMKsMfxx5cQZ+
OuJWPe4EjJNmthw8yQ5Pzn2H2E4MJ7zCgCxJ4WgPmCxWlfNywo2f+CVDYCmm/l/nTlbtVcQKyvqT
I2gncQT26TfTogDpBWHxUBeCQnh0gPLzvoUqR7n/MGzaEeEkI6netLX/srR10Cn/gDDAQoTi38+w
e+70V4NfrIrEAZ4oGN3sZ/flhtB/kTKNqxXRWWNvG9X1J/JCNcvcw1Q0Hd8JBzAmGIe/SbKP59T+
yAqV47MNYQV6nUzAsRlWE04swkUsnpWrRHA+/04m0bQV2HFlFoeX6ZliU1HrZFjIhbgwxlDEYepF
sIMXYbmSL7tKmiaJxb8AFgcPFmA807EwX/CLsGgDq3wGDczOcoxW4L7M9icq4nD3UwdyCf2aqJzz
Jpjt/wO4nimLSlYDfFe8qm+KdhF+V4t0qXoRKEdMfVukeOYmwELGQug2KvgG9+m3D3U5KViaKrso
Llen1KCaK7q7TJMSWIUZqhUaUK9shdmZ+hv2aiMFwbrawClFkY9LjDpFa5UvTKOXfMJjcyX8XpBF
2YJgjNCN20/8S5G3UXurRfRu8ZJHOYBeqn3ntJFnhCUujvk9oEYQWuq0SMUkCsw3kQxPPOJ5+t99
WOMlEj7AeHBNnO4hftHnfKvY8/o1U4yalQ2cTysyeTfT8nBgzEqk5ciyZvomRaeIc/rLMGJGNftw
BBUY4fPmGApCrmCXYoQ/Ze41X6avb08ZUa5UVOwXa/s3t5gzHNL8T/JvHVMBnhnSh2+/SCKv6a51
qiWDE4ldf7nsasitrj5oXTaV2C5br/smd6WTysI7X+pEhU2QRuc4Jea8mCMIQh9vBCOB7ClPgwIu
2+EJaAPug2M+36neOqpqPsSdOseaMNC/oN9oZa4jkm7aATiQ5BtBGOytLzEb74xXmeX9Vz2SACxm
zM1OO/Q/USZfKedLqNHR4CYJF1MU1oIa4PHlpxlTKYS+/KC4z6WLsfwHhxHW/voN3x1wE5S2LwAb
SfSs9DmEdCfUUN/4yPN6jt0wR9r6f6toO6dCULAMsgBEujsr6T5+A5fPQ4AFxTnl0MSk61wjOIqr
XLjmf/uOPShsvRArSwSiFf+ahrY9jOwQdPQfyZeEdaw1KTx8gQhHViX8uQWv3Yi2VxSGI+5UsXHj
U9KRbwdHycD0fo1EgTu8pfkzxCmQV2C04OCNjvopzIMvh9picyIIhHPbRGkUyp8WVhKVIujbExdv
KxW2bZ6yURmMtDPcDtkO31Y8uxqxIEc0IvFjpOqcK5zqj2zkoL5nJbnKXdiEvhnTnf3dqHJMWKGa
eXN+9BuXVdE+9k0gjLL1G9ych9gpF8qkLx7S9TLA+6B3oeo0pKB4czZsxanzGAIpN8RZIEMNCQaT
z8o533KK5JVv/RQFXkkjcKIAsA+Docc0sAaix4k6hRqwSnJVoHycbS0sw9W/b3Bfx90uesnabM1W
pZshOldTP47Kap8bnHZ/yrQJticVN1c5xKh9IkT+oxKssr+eTLl3/5i2nZFZcDFhOb7T0WYu+9bz
3Ig0Eb6qHX3VzHM193gn+M9gb2frKvNvFURbfXGhrusNpJ9g3849N6qYlow5GaYPO1dNfG9tBsOR
iu+mKTRkRvqTu9bL35tFFh5Xoueeh5VVXd6brB3blKosBwiL8pxoGMprCUJ+yHRzz4P9B7zO7If3
tP3bNvzPoxEX7BUD2JVdR1fgRM9pSrX4p8I+Syn7rO4GHJzZM/4xwsdw+ndeLjiREYvow47B5fPw
Ck+5QVUCNc4bJ36/ZG+7ygmFqDjTb6AU2mvIjoPsnTMafFHVhLrQtIc0roH2aN0InYFOBcXCvJyX
KyNfVru5oVCgm5peUAA8iX4B1DHG0P88fFcrwDjj2WkzyWFhXgpGEK5za0DNDaUvO/0Zi8b86EnJ
HKrInEcaP87zlkgFwCWozzC1KwcfJf9h1FzTplzmFMA05rdyHkZTyWAOx0Ce4TtcX/O8iI+cLFS+
jN3hjMipKD1sfjPNemGxt2T+n/diPmsV4DFa6CynTG9ULfxq0+A23JKl+0LEMJJx86V3+VAXejS/
uesewdIIxVLsicHUZFDgLquscvWL6J/O9U3BvzPJT0C/AdWMGWeAuMflB4wcwdn91hA51u0utM03
8nXnSxvHRWiJjObuEs7ULa0WVQDwt/0ix338BZgjowyvM8wMinNSYkYgc6SwquOgoXmeBPdr/PQJ
N3BTTqZInsxNFFnoCWZ4J0pLIZH942FfdNfgRuofgthmpUtAm5eEFe808oOBTSFiJALN86meJNtm
DRofjr2xKBUyA92cF/OoJNlY8dzdxvaUEypbeSRGBHDyi5Cd/EwZbqMGAdlHKUU7s2N/ykR9OMbB
vPa77Rr/FybGhGAkQdwJuXn+Nxn6Amq+81EL8jHz91JP5j1zHm4rqO+SCl1ILRW0VBZegQGMgKWn
hJJTh0JghfvRNnV6Fg4DTWYrf41eHgOihmZQbE8/YL9zHOybg1JwZEvYG25yuF/Busy+DiREyil1
M6aKK6+9QOzrP4XckZw1kR9Ab/T1q6pRhfxp1bW+mlCoIPzJv06Sfybb45rKIoFSy+H5rcCu2/ea
pUITJKl41Bbj5RjByHhKR2RkyqfpgRoWCHmBekT4zQps3GN+LbHxsSEziO7Ono1lBkCakBa2QeRE
WOXlKh4QfLIY/IcZImUEGRrMDtl7DER6fAnOkB3+HKsZvxDPOb9BRZ9Sc/i4EvUHFJXWKrKb8EXe
RSsO1Y4Ckso8WYC6fJYuMW2D+k51bHMjiaqjs6PS5Jh5qJhOLLrdAWnqRxi49sQxymi0fyT2VP2w
4Sk6yveWbPo82a6KuVFEL9E1hWeUChdnwXqnjOONtG7YFadYZAQhjSkeDN/Ao+6ZbkZOPMMIdfj0
FbBflj3G/xHS1w4AK9XurlRmBkhpofEwuConGfDUm55x4GJWw4gYdBfQ8ykZ1fA7XwHTVcdO2mlu
7h1Wp+HeTMtqj9Z3LH3vu1tzq4XOZvyV9iEbeWKTmnkQfcgqPL0ODSgKu28z+nzEyXQuVhvvW3TF
iW0nITjEEZ/PxeVktIjv+9nUSItDeXsSasgFzUkyS13ZtQpRNB5UzpoW49XifCOzwbw6EoCZJ77F
I3Ce/xAxoWXcxT0YoOKH+BX251WiVeaaNV20nVQ9wtJAG14m6NSBJ+nN7iP0bkr/2gC7TOjDPERq
/qX6evDYLKiRp8KqHq+EnoqSv0ohJaZNHGoM3Hr8jKrPfYnuloSircHlnMWH50sbhTldyMDqD0v5
vxrslitxQLQC56lv1U5EfDn0k7uc3w9Z+YWk0gnoiyzXZDS9ZLgKZGnRLzIDL8eQQZwaI7giiUwK
0tw74G5wR64ALLi8DoOFAtMzPH7Al61aT8mhjafZ0qRhbHbC3QA2Xjd3hlxU8MrDAMAJ4j4A8v2x
V7Swi4AoGf/auLvIEFgb31Ox17AtRESVllcoLZJ288nLvJLsSw72r7YyChzY7jYWAXZ2h6mdz/7u
hQPlL6ScjvTyOx0eVOGb9c9GhdS0SITbbp0ieqqqpdYwkYsCjoGb4f1KblDtttO+eSuY0wHEx3+a
ScloqNL9i/l0y+DnKU03nDPLAEJUT138RoGFPhTe9UajPhNnB978/CZ9J/2u61JdS5Q1ywqAQqWl
3BZuQhvJbPxkPsCbaHkhsOFyd9cxgN35IS32UAoDsmspuMcL4fs22MlfClC1AyKeT6Ir3jm97NcM
zywlR4dlFmraWCOo484qes8DRPckR6CeGMigJz1+Exop/xBcn0/OnzlM4px0M8ahWVdFyQINTu5w
WMVBkDBLD7zuyZ/4OF68c+6Nz6HLKzkbSiYrtK+HtwX+bFCNFu/KMONJUR2XIIPnQ2LChT48gJKk
zADixah2os8aswQmbhBPQ0j8ylXDjJUKlq47ZIfXpexWNEMq02FW2C8CqEWufZTRQXnPW0kVT3XH
qdks4ZH22h5cjU2OFmBKynjKTsPk9/SHlDtjTpAqEZgNv1x2fadMywbXGXaZGgmYxOuhmXhoeYfd
d8zPnxDtOmnserOPZ0U2KQYiCmoGtq0wcvC8VRlLvjtLTXbFjY4aZVaaseR5cC0UfzCx75hnWvei
06F0EPGyF28ZGxgcaSU4RXtZLEfPmOTeWceZa1U8CvHdVip4FOx/E/oKa/iyayxHakk6M2kYKXy2
u15NJ7GeptAxRxov8EoS7mFnWRqjyE+XzITVN6Sx1Loit4y0CWsyG87B6INFuWmiOSronssLCcrh
sYs0u7xwi+2nZkgGVJwt0vqwdO8XrvwNMwnKBLnw3ro+Fr/OG+KHAZObDnjwPm8i8pk8gY41DvEG
U6hGRQMgWxuuGSGBgJuwQczRtyIpeda3B5lIQNRLtb3mPGRudeN3Db4GpkKmTwZWu//cKHYFPxyg
yycn2j5mlCCj8+T5hootlZ0iBR4/q2ZzOmfk/6YXHRUmseXmkd1rWvj2DL/5xYheh9wFlpqPKFp8
rMkvXM/XFmW9+eh774dYLKtHV/c1ir7Aco8FvvAb0gb0oZz28ixM1Yb6ANQ5NAldLeGHGKVSIyu3
nSB+VdtIamzHeroyweTnY+1KtCJWEf32aS9daCHA0pNS9m5fw+MhVMTMeAtt2621FK1MrG+qTWCd
UQ9FERmEQBdIWYtzwEEoOgnLX1ICNNL4ckJpb8HKKV6in78SnM4tFL1qE6yNwdhgy5lmwymnvvp9
51ut/gTXTandHEG+SQgyEHX/F5DOTlpA6RJ/UWjMT4xLd2NIx2f/pefSliXIU5JfKI5SaV3YAZX9
CDJeVo/MBcJseuJddtREhDZnYj/XkSV4Xx0GGYxbzxPFjDJ/KtmdOrH8epC9yxuzCp65mfg6z1QQ
7MrLN/mfOQRiXKWmey2Maso5Ytng/4Hd/wyNePXinM/22NeOu7NXS+1hFW6Mwjw0dsRdj6m9ruV7
DcWFsT/a2Q1eWANOrs1PKyAgep5g8Uq3ayld/FMT5blJcdtcTNXns1KGYEmb54eYXXWYuiPBcuI6
agG8VCJvQv76e11zE9qOSZqGeCw/6a1gOmbe004OxoMDnlmQHQSPpoaEOrbfQmCK2nkEc5dBm774
8St6YBRQGo+6YzhBsNPbgM5tswNWETEqtSN79BiSx5MmMRdOAr5JUwP1ZG6vMtfZ2uoGUFWoPp+u
qzpPDJXNnKvzWUdLCT1Tl1mgKezXdF0R5ceF5nS6rE26o66urA+62ODManhIsqdXnXqGDxdGbEl4
XRM/7bshtFVPbRZC6mCK5RhcCitMA0e8Ase33ySMeWRb1op7F9xQIrei6eNWldaW+H+rRLocCrkZ
f+FK3+oDlRAqfyQjmgPcOH8q6kTQkmShcRxwtWfbRk43+EXFyimSY9avZ+V7uKzBStOIAAClyruA
/Bq3RuxhAA45JQ8q46beWTkleuGy8GmCmwHI+6FNdQKcaBAlg5kn8LztOHvUtAyeC8DIouJJJU0y
VKLYVx9eXeTo8KYvBtTJUM/LDEDXG2pUAR7v/xsw5BYEqGmhtkA7aacmxKcds9nElcXASxjx/doi
jaIBmjJLLpYPwGNIqvUruj7lFUqeX0I1LRZHRWPGvNoKDU2JCR7m4ivNTFM0JOw4MigrnV2IaNTi
7ZpdC6l2M995OMeM5jJ/vUoviSxJ4upiuvfsjxYfmWrX3B/Vkmq+leA3SGohgN5UA3K40ZM90uaR
l/PfMZSsqmoL+QqiVtsigI7B/EARsTiFcO953eCI+aVnt8IRscXZwr+/g3EyLQEN5DzfptWfJgUJ
BfVmwo9j7vtkjxFsf8yBih4LHut1HNhdpuOYMJUvgDhrXlQGMHavTzcNH4lC6rXHLc847GRhqHIw
C6tt+zfCR8lPPkp5Vis/7sA55HtHc6OxP55RWjUrnwfYBgvmIyKJo3R1l0doXLTYR9+6tqDoEMzm
D96+b+VPTh97cd3/sXY3/I9E1H763rCOeC7HUK68jRqHcX0Eddakhi/8gQTTTIFgRkYWaUl1+mRP
6x7FccE9ESi+Huw4Jh8TLFfWc2GGmILr4bO5SBLqAPJ6fr4+VQNL9A/AVeP5FaXyCYI43P8eHTIh
1A/5vQfGtFL1UG+dQInpyJi9OHLVcaOkGBO2aqllwzMb3+5aY3EjPlJ1E2/ctoyFyxA83ExBA8ZP
JGXvfj5waBjEUtQHf6xWWsR28j5ZpcrZS2cUFFrndmqKbszoRYFWw8cZgG/9neB1cTmCVOMwGK6C
Vfo3msDLS4SGL+Lj6Lnufpz02bo3JcpzhVOhZ123iXumGHSMYsRmDGo94Cy+zald8hmzBATH6yh3
Ix1dC5vnFf9wA/T/ZHuh3Vfs4JaJBsjM/qMIJpDA6Ieqz5Zgxeo3lbsvykLsdcecidcfgs0MUFK+
09kP9dNWLBx62kN7iFdSRd4elfzujFk2itHa74Qo4WLdff2gZWOM0tHiNTK18o9OFkV+Kymd3KKe
yoAmpCd3lPGEto6LyjQHfNQy5i2Ej/vaD5QMT86LG2vHRPdaE6IiWo62zeAg4c1ieH8ZEopMcE6f
Umq+FO2Qfqn5twzQqYgnVrenVXNg4xp5vnauwndV1Z2imE+cuXusM10FJGZMLa70aH4wQG4EkX3G
mVIz1WUeb89zAcfiTH/5gmXbU00wrxaAcvFcnO9TkSONGWeB8BXC/HqGB4A1PhALoY36fc0rGGzQ
eHjhyZbbImXIpKMLUDMlCLXjJZ314Uh6WfK/g48rHdjqkFmQfczNRa4lZgOkv6GEZltr4v2B87b8
Kqxf5Tte7DIQigZx1JGkO+hvUwTRI7HxgnKF+dOBm31UuvD4b0YH1aVpH/4NH/YOefFuV+uO0l2Y
/8dkN3vsl2XOar+rOYvAc0jqLycalNcI8s5UuB0uwO1QBsC9M6v1OatX5HKvVri3uTLP4tiiAovI
c3fqqku7GEaVQWnTxtY/g0yxW1wHm9W2FrD50kXt6WCLWVsnIhIaxlzncBbUnk9m7eU7GEhMPv6z
b364EgvBrk9/XoU/s5VLdMZA9hWLnd0eIQqNRNQXEzz6FTXG7WGMhntG6GfoLTMZKKyUW6d2Hfrq
EwwsaFc8DsfN0ak9w/6B5EEFdYtUSeo5kKi5NSVdP3S2m8iC240zg1BHkmrfGR8xDDoV5cRj82gN
2SEydXd84nRZtNpcZrJYZ8ukzHOJjcPwEoh4/KxUKDkcjKE1nKgKCuQUm5riT7QcIQBsZRCUBKQA
+PYcvSNuBzeFPPYk7F7GH6tXrV/1sedJOwqBmJj7NXCKpAg1+ZwVDU8fApOUc9ck2ZnnE/EulYxd
MRfAcV8n4jYa03wxpCCiHkREeMsB5svTcBm26P580ZISU1E+5TWa/rs+E/gTmcX0dqYXqTYvgP22
roIcGeQza7Z37dhGE/sYV6++nQ4k+qk45kbLMQBOccNhTzZBT3MIbCrWPWyBEVSmwF4eeqUAuFNX
oI0cjLJHThBMWRJye1Q+AyY1YRp0ptskChBzk6lOeURHBD8g7U1UJmSslHk6cXoX4JDuEP+6kyjP
PEqemzrHCE9ty+34U5mE/dDkElZGmYhJghVNNdYXyhl0Uo3f/J6yO3ceu/llyXbvIUUGylDvaDV3
yu3D+1Mv2jBM+bETOZ6Z5QhfdA/ybOQ+XugQHRbRIPFXzCfHstzFQp8T5m17TODdglV+ztwAS61J
UPEGj2gFEp84rlEwHP6ndW4AvOpcpdoiqW+wXcAmRc/4SgEW84BppAaL1QGmFgz8+1W2sisLvdCH
jSJy1CCYUJxX5F6PQNatfnW4xJZCcTDdns16/C52nAoUrpEHoxbmPFPdVwCpPps8wipvQNt7baNn
iIncTpfHkMzsOQkEndDTMbcBJ0v8if7rz0kmAjihDL6VV1+2kvW8JaFp2O0uk1Ywj61cV+xi24UE
08vqAZkJ1XgUGlb+TMpSGqgTTKGT1us/W5Zp7z6DMckRIt3258jPswqqp/1xI+3O5J94Hk6o4yI6
yRn8NQlS6LqzBFgjbzawj/k3NuKlkiRdGy6nF8ht9tSk7ZYzd3R4/OjjShG6MiYD1H/glnb/yQVe
hmcqODwYLSPFNBDtE/P6vEbZsQtKpo76O3MhgL5eJ7fvn0fiPJ4RNxB962uz+fBUIrhM7OYoRgiK
oJ9/No10slOL5brk/wapDcUa6GPGd6e7DvOlJ/iiQguekD6LqmkeGjZGUiVg6tSB1vvk2faFgqXi
bqWezx6Y92XYCyQ+RnpXNB+kqAbzTXooRnHVvKHWUPXPdKIGnJm0iA0ZcoG0lDaTq9t2IJ92TbTR
66qve/SGYArHzGd36VDp5XBfmOFALm2h3RXonoAKVB/6HbnbmHNqAZFdgptBXNlYFq+jWHkciHaz
posOg/sfu+l7oz4/U/1vI2a757VbIbsbB9zOnyZMKnTeMS8nIr26dQV0tsGvd0d+RhudiCDDw3km
4x03Zc7C0+xKv6tsDz3yRNuvdrNQsCTBV/wkB39/3ct0bp20flydk/NnSV9ovmyjpTrUUk5S7qPd
IAOjotpqpRWrKekRx7oZwhoAC8rmj5pTLQod1DcUIQ41gUtTqXzhUX5S3+FqRDLZ9UmOgUvoNgLy
bWHX9eWJMhMT505+0yNnJecal3KOR3t5fGHVYvo+IHPWdOaaNnwpDzS6SJQ3dKV47iRo5M9pafUI
Rf82m0datW+rN4t2YWFNKcqXN/Z3Ptkt+W7IlfZD/42ETWYCi6KC6C2NNI7v3ZPuqNTI0S/do5mg
2t9u4gTf7aO9y8p5BEaqdlsK/A9X/nM9HzO0lyobJLjNkBlGspbmu6FMkAmn8jSkictN3fnHEna0
xc3MvYcBuJipWMtIbN7bUbDsJtpf0ZzjEZ1OrAtDQK5QLec7gaLixb0Fckd0fZFOIiz6m2FOSqOV
fDUQvmD0dMswv7fuiHmUBQw587mcAnU3KUMfa1Khy4D69SwuQZY9BhJMRSeUuMLB3lfXE5jQMRyK
bHIZvjrWHrzeBalNYC1A1svdT9tqZZ1UWAwQQ/vupJa6TIektHmS+rRWICTK9OilsUYWK5mRe3Xr
7qrEAt6IfSIA8v9YRxhS5+G5Z9fQ+z6oZzCefBN3Cp32vLmJxZSVq/uzejNx6NnOc8ah68Q61LJM
+L0wWt1F2ey6Mcu/otiN7xHX6QrHjAYePXtRs70qNZmURs0f3UKDZalkaC8F2VoaqEmZ1/qpLiRk
WsjbmHrKdU3vVNp9/9MgUGQUBtSho8pQc8bMpwJqOkGxR/gC3vVYSNkcifs65Z15oRlxjp7mAbwX
aKdhgbY6OAtQfdbnBoRNMIkcmYYBdC1e3Mu+chbdL0HVboJ1f6kU0yed9qsi8ScJK6Qsc0wAyGOg
CGkhRdC6oVHbuOul0b4Lh3qq79YTBGtCDFTaMReONe90Np3kctMLhfbbmuGZarj8h3pkd8+7FISS
+vjIzqa6av3l3iRAb7O9gvv+o3mz/NFi79xML+13DLlGceNW/7ximmEy0jRHhythQVL+U8SNkmJ/
x8J28f4xnwLM7/eVpFd5Ayo8bcLnV7i3EQqNFG5SoWmgeNxLkZe05F3gQFH9k26jNGx4xO8hpDWT
WCf2KhqjELPH+uNaoKCyQBUq/h01W5vtZdUAZ9KQ7INUB26v3fhXLVyopSt+j6k6fYR5H19n2/w7
omvYuIfxjwEOdsGfwEnrYYd+WGg/vOABR1iz19BUujsdH8yrDfm96k8fdGPvdZ7c7sydimGqPfPR
2ZZ0UpRsrusaQL+A4htj/DG0HIsrhp0GYI8kV1nrDbjTB6B6PF3WMRrSIdolOpfLee0+Y7SDlyV1
VLtWXhCkCpyC6R0jeR9ahkrgsm7JdYBkl+5ZmzWVlJ7EndIaNRdWw0igDiYSH0S5ZiHrnJfypyk3
hN12qTem/Y9dq25hNR4MoKa5KYdr04xryWARm38Rx0jmrIqkw6AlUch9d8LjSn6Xs9houdg3k2Qj
c48DjdKGG8gBkWvv8zridlSbA2Qv/tzbNYn6Qx6ipOhCS6YkGHuHhbwEkq9Pb7kkvn58CiPSZZi2
EVVmVgDqpcrHZ0OQuK6Os+xnhGeo8+e5EPuzlHhrgQWzNpbFM8ioacH5+RfjUC9cZtnaUiZCxtEw
nFkM79Qm828a1TUu54rYHgoRD9A5gyEErOV+D/igtq/D2gmmpDs5GXI2gbkNw0aseWVr9VgOV51O
3OBO+itWM3RT59huAuPCCJM+EbTZt5RFesBoXQHfti1SYAhx6PNzDdugCckmd2yzGfO6mU8KZseR
OIdnbj+HXAW/LGEbRdcDq4vaayqlTcv26oI+TDRWwqdVRMEKYtH60I63UlPr2Fl1YXy5HpXB5MWP
uxnA4y4dBm5LhwcPINzi4Kn36jJg5lm6zwRGe+5Uwri4YEVdRPYMW3q3BmCQ4OQLk2Ytxty1EKdu
XSkAQJ+eyLZOywJSsSTW6Ckzvgrf22j9XLTHQnx9j0v83atVbNlxVy4P/TPMHo7ROR2C92QfZwIr
bMqDu2E26ctg4gmPfj/FP7ITwA0ec9QiYAd66ozPaJFBG4r7IVFvk2XfxH7AnKa7w8fIUYNFfd6P
II1LDn+XBSIiCVfFhth0QbszqwsJgUXlBKNPNR0UYZPrDpWGAeprzun3hYEiOxw2WJcAIwH25IAx
zyg2dBfWdbOS5jbxB+zKebXO1Rgqn26JX2lU3Xopg0J5xtqJ3SzPFd6rrOvt6+mwVZRbQ6Hhiv32
5KKg7MP26Mv/C9eM3bLD9+PPywm9Cffgi8V3vq6Qx47BHk1r+G9aN2NHhzv6C4YnQuyKtZDm2Ywb
5x0CdvCRdxRdPhGNw4UPeMRPQ8vthpun/KH/sSeYqgssqgW79qRUFegojeO0pTG87n1DA8c3EUB4
KdckzqTVsbZjqeD8i0KtMLKzj7bCWXxpsTtd9TCbE+bzx9/rrpSsBbaZzpv69VweoWw6VLAzVT5f
STB5khr6Pttwvi8oW0CbFkUuSlaDo704QOsUdICRGwq+dOhWmZdz7bb/ISHe0t1gzVB24np3K4HR
1SChzfVdSRWnmOprYbw8LqTrdfN9xPxMxZl/KVSPBocwG9tTZGSqkaeQd7uNTToF2Cqcl/CyFUUy
d7cgHxwp8gg2Epuh3oHYSRh0+Xf8ARTBHYBscl18GquOq98mDhf+hmWJch/hCmdS4sQLDDM/1ghj
DR+njLW87zjMPElpG024LRAzw+ehS5l4Z93eA7zCY1lqFFMnvE+slahHumi8RUZtJz8tNh8z+CNU
yHL2TF+VmT+iNqgUYzNo8iInV9uxOU/dKhdkqri2j/SG2IF4KKEPggMOdP1wSMavBEdlbmriMiEP
CwUAFjAilu3buv/GU3P+0L+L4TJVkKPgQDZlM75UQMD5EOtt1siOS3DO3OrHG3ijX+RW39FiMWRq
61Ywxte8TU5InEOTkNtbWikgif4tcvnZ6gYZsjHUcBJLfCNuBMApxcf6wml1nKgHQb9d79vuZelF
JSyVRnuq5/p1/Iqri3pQT+TnhWDvCMUoTRAx/ZQ+8oHrJh1chkV15qApUMg1y++OJowLzVSF09yW
du1MhC5CHQ7RI31rYAQCJLl7/HMcV0inrAgJdY3IV/zg0TMD7MKWyACQfOrHuoasTprvPK2fWgQ4
EF/EnnSWknaOjEBUVgpPOJFeTTpIMZvaO2z3yhUh8mF9tni7p586e01b2aFjVjriZ35Td/E72T16
kyFThKvBG1O774OKtV15827aIB9GKgZzplpSt7MR1m7GRJ1Vh3mwpP6nyrWfNo8P0bX0deu2wFnM
jIFAxJ5FLe/cDZKQHd3w+8tALP+4bmwa0dxBxziplqTbIXPfXUXUNvXAxwrlrnQdn6/TD31+PmYi
awuAHAuexKo6SHyRjbn7ouw8SmkXGRtBPG4PrJmsEHo4xmlbdTr0Ncgqe2VwoBAELfPsBLPG4Yrr
FE+WK5U4r3y8LrrqlfPy6Ny+/xN0/Ex04/us9Uf9JkXJ1zFbm4fqvIRiLScjrQKKI812uPwlqxQB
2pV89w0vUbuhSx5T6qeUcV5e7kdyxfg+y4WrshFAsmBMTd5+2kyxUKwq+U4NVSKOdoQ7ySRQjG/l
F1XKt4fsrYRgcHOfgMgVFAYj19SbOlJerrRhpv5fo4ArNkp7i496CkPv9Q0VRrtjxE7DzogEoLbj
UeoSEpKWYne+2ZrL15GxOj+wSPMccW+i6RNNmRarxOLL6WHS+0U5nQL8fKgZeeOltAGgX5epPJs1
/2CK7h38DnhTsO04eRXxmSxnm2KM8hnA/VrJrOXiIFOq/vjvFngGJCxxa0/utRfMSmN1JN0GGnf+
VQWEwLz6MfuGKvSP4Wjbc4S7ApwfFeU7FqjgeUrZphlMFgezn+Gs2hyaveeR0kMj0mOO54/CfAu5
asQR5yOEDwJUQ5IEIZvIBiq1ylIoWCHFNshTJRxdOoaJFHdCkJYBVKHahvfZ46OgLRC5npvSR+6N
7XUC/IeUFPsXrH/W/Q28rZ8Y/JOZzQHttdydAYjra076Ak0IolsT9zT4FY3IfjFPMxmw7FBmq6N0
voTdmeBIFCDorfoapXcv0J0e66c5lm5tjwIPzLwJsc/h2Sb+of/dF8j3Mm7DBdLOcfTxhC95VKE5
5zZmw3b+UL7ipzmA65ZZwT+QllmHEYTsEOpxP1s0/QUI/adT20rBuSJVZIxrVCw9p9fL/a3vwaAm
lE0hv60UB+EnPksl3PlYeFQcv5VJN5qvitGGlJdCbkvrSXLp6DGgLMdotw6XH4AcDoCSy6ORdlIa
nlv4+ZVMeFox+boMHaGsTF3aoyV2OdAeMgHZgzBzdyhq8t+we/WrdKVRwge+JjQgvrrv7Qwu9CnU
cVEnCtj/XRKNsZ+bV3fTt46NuMcdH1aWKI//YpxHJ9qsu+UECith13giVhI9ImffZbq4yYt9jxoV
XrVmO6YyN2BcbPaaOgHq2M3AG2FkFA0RHhliwxJebIce8+Ic/UVkNOsCZdYXPqPyAXxQfazO4Wgc
R0ZuRsj18zl9iwmU5cJvHtRPj0+rM+pE+IwdDwgMDEOSJMTOz/JZTPbF4hg2W9Y1w6xU2JQ+H/8K
S/yW/k9bAKN00M97qBKf3yIYMTDwkjEbzh1NhL6LQKyVgDVpURG0ktN+5Vup1xtLyXonqPw2Z6kU
ZfMSlpyylCkYi5nKkWWipBDBIVgsFmYASMS7n3PP/6ygTUUSki4MgoC6jV9GCL8PFt4PeEy2bdnK
5CFvnISRm+j1pQ+GdRvQ4kD32Pa5Ee9HWA6Iep0ZNAYOFLCema2v+W2ToYqplk8/tEjs8BW8FW7J
ltM4vYiSmV0eZ+nBB/2E1caSzhFaSDEts4Skkqyw63Lju51c0oCR4nn9ba/3juSflrhTG/fAPGfv
FXoMOUsJtHBdmWzxRpSGg79cOvTAqjsS/EJb4iO+Nb0QHqOjPwyeI79ENHEg9kg7l0ZfbAZOJGTy
egHSj1Ij8e5x8E9aA0Jfdl9fzJ7UskKtIswOcc2GihTj5EGVNUyG3DVfmp2mUMyu7H8sa3Nw3PXP
SMIB2AvTV9V7aj+X6J1aTGphz/2FzswDQL3t22j4Z/DB75Jevc7Ml7GdC7TfkutAVGF0E+BzI77k
KnngRgPuJ0v6WvUabYg3ckH0He3LoEuP7uObgREkcLn0Q2LDi/Bgnvh8zC8HswWY3TtjMRiQpUg7
OTrXg6viLdSNGB/QcfVcdhbQBgPBFoRjAVmD7WUro3BES7dB7hQgs/gC8EdL5ybo7p+/C1VTF68i
C/y5yHyh2Ak2pwtvIiO9Xq1DGfqZtR3lUIvEJ4wn8rB6KETuTiLCFqXryLTk4fpaLjdwQTW2Wxhi
oyean918DsgaJK7BQk4XTCQsM7+HSA8U9ss+u75dvBesjYhK8gmLjsohBM82zNTI3GVjOUyvppZo
79tigymgubc3lvZQ0rQ1h6HbXrn6HbujGL6rcGQyTYoFIkkcnM3SjNYfNJS5RRBcTywQY2KpbLmu
J5peAkA2N1g6nk4ZuAX0iWfUGM6Lmnn/D7VxOHtiXH9J+/4Jpkz0TYOYIH51F8ZGWKTkGlI835yM
YFVYHiR4PKQ4D5OVouni1YnSTPETYKKH/gt8JhNqCUNM3L3J7Yuc7L1SvpJDnGBDrVCvZzmJofnV
Lv/P77ZbfElp3rWBWwZMs/AffNIzTiJEc/7HlORJ2dl5kYIKkkS4ATrSN0SD8SsoEqls3gsnT8mc
KdcnnZA43mywHL00lwtZhrpxcfN1jP/YnauGY5rjOK/T45LO/kJeB2i2oyztVSUvWT9XGuLgCZMT
okyEr5Poas8OF+Tu0CVEgPzNMn+T/g653LVqqZQSJXVuFSklHNd9jCLoab6bAVxAtgaABjIQM5if
/+WKN+RDSoNsXNE2HGgYjXH08H5KGLZ9rWIyRusbhC0uMlsspZlFvdK/52n2wE1EHPoi0B8ctvq8
4CqYBnfdSy2DhdsWByoqZesbkVT9VJoRJmrzkz4p2yMKg4vcG8yogbMJyTIeSj98MwHGFwoSOdOU
DgRimpFJ4SgLLt5d5Dicw08XUtozwzKmNu5YO8B6mXn/18qjw8+mzq/17I1cDf5LCGlsu7VZPLzC
flcX6UYXEsSsYQ03ZftzPLkd21vZVnXJ8tOTwPpIP9686s5nL8ceI0+wn9SJi9Wjl1Gwz/2AE5yb
ZYAueD8y/fvtMmIQNQAwcZhHJeCOWmAYt5PfNWVAPlna7rGsAutIEJ2mfVaXWgNtc3rftDsVgd/u
E2VVsjJhT1QU/RJaa63D02QdXSYvIqC3JvYVrBj3MytXi7S4gULRdE95cWmGWKApq2Ezwna0TeFc
OevEi4MDNbi/dS7riE55+oQ3rDxXI5f8Dlq4D+voWaP7aYGHEatXpRzZEU8KBxRInJPon0zvNCGU
tP8Ei44ZSyohNGMNG3w+9Qz/VrnygGFwFne3kkqLdwBPdn7uh6Ukpt51b4kBSjkvP8wlisoBzwWh
nb5tOXr9mTpsBtlkUtiCLsdwPwdqUi3W2ulZ3Nyems+OXkLqyupyhJc0iG714gKJCpFE7fTJzcx+
JnNvJ1DEIUu1tSHhBU1fDqb8fAVjwBDB5pf20oqO2SdFib59gDgGksSxogdo/wo2yUo7hwjFhBfd
DbqS5AJQzj4UE/nz0QBPseDh0lKBTutpcjiQCvi0KkRHVSjoa0lB5qFXIsn9v/l3VQOs5KR80pjc
zJaNVxvH4pYCMtqY5kB5JQk8YkUEHqGybVgaCdujZy47MyNlXk3WPIY7pDjBho23EU4kPmFONsP1
T9qfAxw9wXBC/d6d9dScEhqAR2eZwkwRguddDw7qfys1VzobLKvS0l92YwGjMy5eJpHVQqWkMV5x
WeCRt85NfaMnIeCFi+XfSSp3tC4sN0t5KzC8PBI+F6eyjy7t+a7wdlQWYGVaA/tmNHyxKWsspt23
4ejgsD3DVUd+f6r7VjN/xNdLECBKWaIWESLZGB+xlITkdUVFOWmpfM1H6hnG0GjsDc//CArK9zaL
EmAvhAm9yDjYiamo+T+oWlrP6wkNDgkfhuYXkgSYrAvFBKYBGHDRs0L+RG22YwfvpVjW9ZBiVHLJ
u4oOxdvYvTDqONerpiM6BpAL91oGQrxlfS115eEHdo7cvOe3Z5/71mqoelaRoQ7v1Tjrmou8XSRQ
Ym9vfpkmriZPBmAwWThnUB2YnljbsQqOjuxRRlpucT59/w6dDxD0s9mfp/TK3dxwbgCI56QSmpUT
R5M0u450xPAX2ebNTxbcg81jpnvfO7kXWFKFj1798PA1g2pJZ0XUYCVRXiyebiiWq6huPKeWTpxJ
oAnL1WMFhXIKZvniApvffZK/iUpI1hTw3I66KHMDSQFZXSttoCGWDQUWnskAlBTbK+fJI6zlmzzJ
VCRtI8anNGSAPm9pSp3G/t2LX51hoGdm1T1OLCy/dFRUB83wEBAOV4emECWQuSbI9v/36AWW1bbf
dyQGPyTQaa8aY/bM4HeatPJhAiH7ovg3v3FDtQSlNzDNUUefitSjOs5xuV0BRYEdld8tbIN53Tsy
o1UJnuOD2o8gQen02bBCOhUuGyjcD99cD70x7JZl6v3hGbUdL6nCPc9YCc++aOP6mTKAUO5bLVA7
bdnr2uerDLMNWlqQSgjnPQkj98LI93SLF18XRWGv/DjErT8q71yadeXZQvXSBp2xNw9bN1f0FHyu
6dJoeX9erFtDNLozvi7F0nRiluu9nNNrmi6HQObzcAjoH1JYo/qs1mPb2VR6NghyHdOWTGVuT9pI
OTK0dUazC4MOCdzuzsF9ORnNQ2nLJ6Zws62fs0Rnsf1jRe/OZ3avlVaUphXnysKXzr4eFRQveeW1
OsWyRrY5u2pVfAaeijQMKgq7QQrdWCBvTfoypruwdquFd/6Ikk81lMmZXiqSRL+7F54ShD8qWqNl
/nGE05ZNxCxtqat3ZPqlc+tMpBoGztKNRg3KjQlOeyCJIRBQyGL1daehAqLqOWVD67foA0mXyP3g
nIVPjLdAJMtJeis5kPv2UICwAAdaItQYOr00LXi9YthLS3RgPggfSLeMkzkCMKLr6ap2OXYh/hTO
HjhVs9sAsiBfUkK1EO+9gpqY0E+7v7PvxsNrjsSejmE2CJJu5+X5rpykSPMzpWCkwxxQgZxo4XoA
Mef0D4cxqN7YXJe5Zq3DsTzqWvdqR4MWA+fadyupvZOeEL4FnxhywPAv1GJ3WS9Px7EsVgLh/VYd
DkHH1MoIhV0t8eyTH4ygr9LotRDXHwbbYNGD59w+3wHNaB5Lkn0UdScCbQAva9MadieGeZo60m0p
Cyi9CtYLE7D5D2UM/+Ad+4GA7i2wUgCvElX/C5qDg+M525GdFqMlR2rH3TW5G8HtJ5TzDtuuSTBO
F5FPAut/PK4+wt+fVGHpBFeuL2DjEpkzh+lx8TlW9KQQi18GdzhMTCJH9JQp7MTKo8k/7evKGBvP
IhDdKWrDkhF9ZWlcatanomban7JwSTKEogBhbHSh4H7KI9CVOiGRJLnzP/VpXEnhjoXK8DOyU8Is
0Ku9ifhUZ0XhXfdPDsPd1stOR4iJgRooOi0ltFJ/WEXGlenxL4cC3nedrDwQ5PCqRaumfGqXTQT/
Wvm/JGIlLB4Zie+9lqNzZ6kiYn71IKNXnuRFqP51vqw49T/XJvwraVcSStHG9C0u5c231u7cZBi7
NAvaAPoL+5M7IV17L+apuw7YRojDiv6FXuv/eqyfd5P7MMRHY4I4teNnvms9P+Wg/HKjjYniihz8
OqWrxeacZqR8RMfQfrTNmvkCggUgJJOB55/ahweJfhNkpkNjan1vtu7KI04dP/T6K2+9P6OyLJS0
HfmyLWatwQc+D1BHjCUxRsuk1Yaa67p2ads49nDl6sgikZzAzlcPlJ/3jtY7V/1AuPK2iedv60AU
iRTO1g6UnVXnxezcNiSH6lA7ZMgZnI5u6fC6pjD30B30h/AY0roPTFfXNLPKoUx2Q93L3TAMcKUk
CAlcRh5+UyqWwJBMzNG2sItupfu5u23b5tyM7FBhkPr+Wlno3SI5fNvJYv95XCLurLiZpOqHf4Z1
8+/Iyvm7LO3k5kjhR0gO0NsVlTif66+lPJcrj+nL/GZk7SlxCnY+ILoC5E10H2YkvrVgJwykwI7O
ieeSGOyc7yX9QPNzKrNvG/Eq8jCvIYTl2df6luddruuPR0p4Q+sjR3RC15BAqfdLkApdnFxq44T5
KsK8J3wS/mW9K7M4/pv0ULZbmgSVVEqDWC+DgcHihvwm4TQE4/VGpVxaml031e+iNQuiWV7IcCvS
QbH4EkP8+Rilpm6XOHfN4dlE054tWDXZwGcDn7bftEbo55oKS0+UPcvCz3z9drPmqsgQFsiPtb0z
JHh6XA6Fmu/t30kOAp8UDlPtwbQhOqTcUJojU1S8EJDlcTROW6Dx8Lz6Cn/vn5qouHJ7RFyVYcv6
OqURG7qPMScPbJhNn+G68NsTCn+GYxHQ9Jho21xYO8s+Jj1BInlcI+a+G52U4JvIdfQVYhdHfYAE
DgmO6XDpPHyfWml61iUS6cgHcMkP0hkOZZ2uh3AsFE8XV2cVkwPPAO9DyYL8UaLBwRtwOZiuctta
cM65hMWr6iOTkTsvTowRyc2dA1GsPr9MiVEDMDwGPHbr1VRIB5rDNSVBEOoJVetIACIOScOQB70X
6HqElGhKhXH5ywNwGY4DvzevZKy0qqzMq8323zOYbwTzTswRxLFSv3K5Wdr6A8z1Ve1Olk0VYRzG
/adffTJSxlLow9NaonDCJ0mqXpQdao5kKuDTGwOovHFm5J9oeNg1UcHve92DlCcNQLJ0VwE3uRHb
s5eU30ofx8/gFIenl/OhsBsYQ+JGOWMPSiTeU+fH+WNarBUWZkSyKBXsG2tnoYQ9xBmH0mW9rBxX
flAKgrcuZpo/JoH5UiNIQ3nnhLtMrS8M6IYDjsdR1+pyYuz4uzvNGhqq2+r9RBSizNArawJaty2D
8I/EPDh7haucXx4dUsAR7Xl6sJUbM9R1+jPPz/ZmCCptALUub8LQ6nPb3mY86/wCeasJ8v8VTVf9
YlQVrQncXBHhWohFkx0hoxioL+nold8Npqibo1vaCCslkrGBT5ZLLTefhnUd6qrySOythskFgAdJ
At0Snfzw9Ql2IYzdaWfXG+aP5FED5auRdpzdBZ2sWg+2sdShQ3Nlt6lVMVOCqVjeqLaPH0DFLXaI
3adNPQt5TZgfYyYyygnTtthmT8qOpnIcxJxkiBUM/3Rj6jC5adPBR6REDMI8gk62jkc/XCpakuuE
XRqAmTYyshNC+mCdyKkU9AwtJQnFVlg9nRikZx7774R4KiAiA7cSBTKvWM3yBjxLkYrJbneKYcLE
8YtxxvWpVVfzChc61Qzq6bW8lhv1Y+G1eQxc6F1XelFl20AYYKJHPOyN23rb0iAZTcumauScAabz
iZp5L7aS0SRgldt03xIyNPw9tRbHYJP4rX7FMr47b5qZQfWOD7uYkIxlL/97DpYVugvM5HAz30oL
64aQkh/j6cKIc+L1HeheZCowovTD/HtpK4npgSH7TpSnDfZ5ejroWOYT7by65jN2y07u/gBxO4ud
Z4Nhkv3gAqyXPxS7pggqFWo/S7O/e4xNPmFgXNbliaPfK0RqdVhTkOKycPPhRyhQg9A8w19vwi7m
7rG62vcUfNYHp4A6UHv2PiKDsFpQYCx9CouGZ6vdEoGBap5cMBo/JMGF2iy8+FbV7c63Q85kvM7N
875dgjjxIUMM0azh1I8m3J8NOYLcm1Oia1VfzrLZI7y4rG9syN2YJbArjokcSZd9EllpSteAVHhg
1ndPoa5KQp4jBuNITNFSvwcvLiPmAxu/b6hiRqdGeppIz/bvmcg3OMhG1HdCq1WSSIJHsMEf32x7
9EHyTMtDczBy2n+ZnCx+EZcAjhriyo91JwzTMwg+pZkrtS2MdKDDe84oTh0q6kzA5rhUMAikn1ZI
fku6mDbZ/k1wJIpVsBbvhZh0S9fTSDFaj83PZabiMFM+zH5ntPgvbY2JnUEQ3cl5m/RcjjFiHSjz
F+8bjY7JGMIQf1nXH4S4+saBWzj5UYmoII3fXYyi2oUOAzbB+OxaK3UJSQ7GbRrZ72qm2UJsqjeP
xNLlb0ySGeWO6FxrE8xSXrL+l+7ABsYYrQ9lvQTQH/Yr35r1xOeGvWTt/D0TlVcNOpKA87+PmdR2
faAz1PKUmjvwGIkmNOr+LZd93NyPRqhdMSlOcL2OlMijTRAKPeS2Nqp0FcH5eeRISllO6e5hbFAy
FXXfLQiJ8G2xoKxu1bhyRNMQ+AXcjXIH1hK7jyWcrbekIOwCnSjRmBsBWWfJUQ7Cnnfo+FxdgI6g
mFJIMA8nADztD1aXST/yv/uVQQJuOwMU60INKkI+WhNSdlA5RGJvh8ILToUiJ5dj1klwuzEKBKJQ
+9fVAjRgiSHLetdJS739ggO67pfsqcaypZjVqXT86mGPNbk1HJEOTLJ9RIBdE5WfhJKecRvJwoQZ
Lb5WpBdQoLpv+uvszz5eHQHKieBNth6/wRPakSRmEnnHNwkHK8B/CDXuq7XRtQerl+WtnYQqb7DU
PT1jz8LZ664DoMKhEu5/oy2mh54m2NYT88c9f5Intk7Roma11cCsLxUAMCXVLzMYKirtMlDPEW/o
9lDvOPOnBMm2E5pcQsxcW6T6X14xEyjL0YA54jazKbpVMbRxo7NaFvhwiaWTkSKX0cOq2LQjrDuv
mgT9MzJ5Xnky/H59OZNDN6AsxlIXsEpmPuSt9/MBZWS1C/IFPymydvE1A7YJ1ULlmmUV9bn15Tgi
vOdE/ymTzySE40ryVIP6ow2AFKiNRnlJsb6CzzTmS2Ept/tAUSL5pIg/RbUhmnmAJi71sFOxAnNL
531coDdzboRYq4bCkIpSlz/iyW1FhZ17IUXjREeKES7ijklLFtL7AldWE6gHDhnz+K9AgNveIEWd
0bM4ODwGLTYMIizvvSKLIMlC/9y2zeN0cKsl7DkInHJ8viiyBhKxBxoSOLiPr3q9l+SYSvSsFSje
srqm1fFo20RdoEz4SUnG5uBZAkgaCQZed2Kep7yi0S0JJfxqJevIzItrD09C5pSV0DtBfrPWcwv/
DM61oFT56/wikmebQKVxVbirw+/IoTQbjlcphurHOK4+P/M9O7rlmoquySzPVLHtmXIh4Gw1abXi
FaQg47NskaWgTAuFBclV10S7coJqkSFgPdIo2RKuDxj3E/gz5vSuMXbkjboGqdIpM8vg6l6uCeYl
ikZvAk2kiOIp0tlnqTcXMyj+7ZhC3U6Jskqa3hTDPgHwuZWLhMgL2DheNz5TDvM/33Dv5ow9oC54
202y0W0s/IDr2fIU/LUCXf4uqvHEdT+9H5rXZhe9Wv6z+1fQCiA4xBVK1K44gCGWd7Gvost68AVj
7ckk403+uLvQK4t83OX676If+FcLiAxnTKabkVzMR5qtST8LWeloPWxztf6HzgST8W02vykS7EP2
BlI/p5KwMEzpOiTjnjDc9IDuyRi0EN7CnuFONyaxDcAPJ9CUnPtX1eWFR1G07uwVk8Zz9uBKOzJ7
pZgXk9kk4KBPckHqvbHGbiPq5HOQhKUoVWuatMVITMpCr34PlksHLpomiYoH0onXGt7BtU/THSn0
DWg/rN/k1wJ0OPTnpZU2k7wOFZtdbrdz/hxuptY/vWIWeD7XvaYNrNfkz8w1MNJBl5OJNQHL6FMi
ytBCgawLFrdPjIyZfhg2wXCbq/SW0bL7Uc7lkR/N1EU3CvypWsbxOwgt+MsCy7rxzRxF0IgFtiGF
sZA+yPTtM1zch++j9IR24/iEB7QOtPM3MZA08BHFIT0e1Asw5ZHoOcii9zZb5or/GYlLCZs9HGaK
/iESsmEf0zXcpisKmaAaGV4hHvll17pMvJL5RSMTPw9s0ASt3L3xoMPMaW3zDJ/d/MetoKeaLWbz
a6NwCsgr6xA1P3EytY4ze5txuOkvbkEkfXPGTJ8IeBPjbdIn1XgsTq44u50c2EIhZTK8k9jrtanJ
ATFF5kbIocF3jnx61KPIHtmbWBODsIgxv5jZnd6i18p2gDywG2JRKOpphUUrQYqOdnPWg8slUR50
DmSGOBzuyuiG6wEgUWAhmNjQuG02asqzNlvBU9PqyNaZVa8gBN7Xj9T1mpQie1A73+xYx/O1OXfT
Ccvbngb8k+OFxfj2sGQl/zfLnJsIkAMeXoRQZRhCwJeLuLK1IOllzyKIgQDmMo8q9PXxxJYjS9yp
rdWU5I6tzhRPqSFBzNNtMZ3KVIJujUTFqlW079ba0lOhTXWy5ZHocj4gtHMwTfaDdPRt8D5O3bqw
svjigAnOltnzZ6vtNbl1sd87/IpnaD1VAaZN1t6tkLIUgDdIVCHQcRCM6+oyOSOBYtle6EV1cfMV
mWVFzW9Znh6tGjzT9DJYj46IeJlXXr+xvR/7dfFycgD2RIv4EHTUaJ2Su3sfNLFe/zxTvaqc/gtE
/qamSjo1FfYgY4FqZrrUEO/sw84Xz+5fAQFH6oAczZ0tKJZ4gEzWx/3f4WRCMMCiuPS0E9dB4smv
R2t3A5Kkks1vnPP9ZdNt2zXuTRY9MzBmPb3KXF5qZDYzH1tJ9gbhsD8prZu1NdVBo+MKiuNWcyeY
kye9iItqf+CxBmXhA39yetlTLtCNERPZoGfrabQsy84E5APCB8DQnnrEPi+vCSR+Znmtqx6enyE7
9Aeeuq0kkisnFdhwAy7dFmEv01Hw/cgr00Px+EX4qie8PADZA603ec80uOPmlsyOPeGuYCXTOxnF
+s3wvZYQRwEOzQ/g36pr9Ub++Fm1RrNU55fwCLvCA2FI81sugKjnnf7KUddrD02U/x5q9iRyNLg6
ubo4wXUQwEVsKPgoaFi0QMrTu7R/NaQGPi1Lbh5C/ZkiPQWvSAthlW5z8RT7SOtL0zE2GuNUbB6O
Rm/IR9hva65p9ULfT4WDjWVKq33GjYPS82Qgl5/7vgvPJAIE+FUQsBM1TlNG96Q+1ihJiktXYWr+
wextHbxw4sqbMRiiTk58AJbIIx8A9U+Jo0sIL2n6uCUwAY7jtPbZZafVFEqGVS4lGezPuk07l6OQ
pFFloofXmSlQeSgtFADEzX470ir2L67JyZ4prcaTGm25WhE92qj/mPJpJLumxh8f1dpmrj5udZUX
6LILoz80bhaWraTuZVqLbUgDhlA2fyFeWlVqUO/pHQCKjdH/YWsUdtPclGa3WPR3IWSHZTUXPLLR
tuurYG4Myza5dwCigLevNvKqCL3XgXNPMk71d3CvEoUQnhxL+5jr5fVrJ7mnveZVe1coiWWieQ1Z
ow2S8ccKziWeFgx2H5Q75+AnzroU5Tf+ptnH4OHgrKKG8YtEAhdFUmhNg/z8fhriFk0TAk4NIi8o
pDRa210EDchYPwc/rELWxhVkPBhhytI+DTyWETYMxeqOlogQkWy1Ap5HxfqNBPCbHaL+uxbqYu5z
VvotRc5ob/qKuIyalGdf5+ynSpBmLpaNiYZg/eyT9TY1zofUl3GNUbzaML5r30SpPXxCqh5r7Q/u
X3/6bBaW6eEbTKRzra2Y/++QdEBHNCwS8ihV2tS3Dxh3BSjJAszDGwG7a2WquCoeEhEO0KyVWa5m
MTqui44T36iKvmJkNtIJ1wnmU2d0GRbJWGh2jmECtdE7r7/Fwx2JKStB7gV/nunowG9uFfYRWZT6
MMsFoYPGjz5a6P5aQw8D4kgziqkR4peprKuYzxxxJOtKc9e1ZUugIVa4CCyZYGpeFb572kPQEHyJ
eeGCNzMW6+mja+b0AbA7nfMOVYxo/8AKH/hNe8ZH5m6r9dbcvk+19WVsB1nWQ19wXhoNogrrOpsg
ZtVMGg0dWI62F/ryh2gaq/CJBB3IxswgzbQupdH+iAWF2uxfghf35bgwLNuoLibKiehAHFvJDNLC
rKSWBo0cchoZtLQiRpVj5cTw/as1/cx/n6y5gb6O9l4ffMZIbdH5aGX39j4X6vKqQgdGhc7AxO2N
EmvR4W34E6gkxiZyF31xZLuscrZfRo5VtS58uV5w3zlLBYpT5/nZjj6L2JVBAApSpsP+aTKzKz00
uHAtfOSAEVqfCZtubddUu43uf9BydyDRkcqwE/nkhAT5TWHmvH+ydmqKb3s0mUq+Okp0enRQcxLp
ji4h46xDZtSd7/du7ZKSt4xVo+JbD/leyShignlLvhyKuU1F8nuF66nURO0fGKBViz1raKnXbfnX
auCU6FOxRUSrGggr3kdbQq5BffHyLnr4bLptqZraZu+p8HWT6q658C/RDJdCw+n8EjKxIdJXrUbX
A7ErnqdYLEW3vhJbz7u9m3jE3Fml66rLsNIqBQUo73k9aIEl9Y5o6rwigfmBW4MJQ6SWZR7YvP53
uHhqtCF6EIxIcQUmR3tvC/RGlPETFECsT7qiWujdLG8KhDy1dZRF/eP+hylnHX0KGrnrK/vUzW3j
cGid0sbzAeYBgfcX3wEYSl3J6lj/k8j5NE7pIBPPniz1qzoxmI3HAmVod1DzhLpncrI0w1jwhi7o
3ewHi/mAZkdK/2oVTHrba1qBJCAoG8O7nk9NK9xLy2CJHk4UcIT96rJXlFOL7Z6eHYdexC63m9/T
k4X5NB1xf1jXBUiPHHakidkJ0oHOFsAB8Vx3bOFa6+zox17UygM+T/9RNnka+TH0/5uRjJ8NnwaI
SipqNnja1VEbQoDmCzYUUKnGmwymOL7/GTMIuZ+oFoCSVJ+02sfGYWXngDA0+AMXlcOZIL2JcoZW
ZJsMPAUBGYkjkvfrwdiM/SJrSfP+MBj4oGe8pwkKMMbW4qZn32kYgra9d/vyh/Oh8FCAm3WPydsf
mEghv+zLXWwxOvIh5zUGyzxrDQ3Lwa9/NgXYmjpNkqdOudeeO1nHK8cdSIW376sFU6ldcnlldc+W
CdRPLuvKs/5/N6Y3CJUIgWiXMc+bD+cJBw6tVz5GX7bJZ9xMWMsD5kbBPzOsNSYaMW2au3TstTUh
hhaCImuWp6S5Buw6d+Fwur0zEIjXU6XsdLc1E317Oz1kQvHT5YXELBj87XMSNzfnGLLbNKkLgsYP
IiuusQH/JyrFVUUfauXZEFtVUyD05BYg8DZgG/HTB3TS5mFT+uK88ag4YZffjnZgw8O/QrZnyqX+
+8qRjl3NSf/XX/zysNGb10I6Neo5c5zDdgMbNfWvBw51R6CeGM6YThv0rQLOdpxZICp59FKem0sQ
9ErTBq/+aZCtLwaYQV64IbLfD6Dw8kOm9glnMfQtxdp3ZP4Qe6N5RgTpZaEwZOd6VzGAF3n4X9AV
Z0LoUsPWspiwLQZTTRScoLWxzaTqX6Uiaml261IJsRiRJbjWBp9GKHdqZUrPpgmloR2iQClwBBu3
UDFN9cnfEeMcgfyH1Dz6WYYEgqYbOnVPMYZowFPcfs9XrHuj9OZVzQ5TWIWZo54I75b9fLOMujHn
pSlhDdO87bbFcybrcs4dNtytbB36EJE/8lWL91FjRSE9fiBUgVFjCYYaoBsHp+fxK5AwqU+G7z8I
7UkkS8j4b0YgQk9L37e91DrbNhKUgL211HZcVsLDp8Sy5g7VSXGM3lVox4cr/ISn6TZLmhDhq2Ue
ZoyqlS5ZLqZN1lV5SOyU3blq6Qok1msyG5cfABflpDQeTIeVJ9xjM3bOk4aHojhQMiq6VEGIr25w
hGDJTo8wP+gBnIvz3O4SSaaHlffcA2mHxAp4sXL2CA4jTM7ZHYHl/WufBoxQOiiu1f4L7ckzmIHg
KiNXh5xFWr4eurK68HOo0/Pte0N/54N19cRnd+dN+c6+XQFXG45iHzgfrbP++j3msH4vFz89F79n
J+QlFBBO86X/w9AVXytuc0v084K8Ml36tTL6SMkac0GPU7bOOJUbvnodO/GIOgI6etHV9zQVhOWc
QkrneN0f/60FdxbbT+wIz1hzJlXuVrKR2dl93WpjdTjVOp081cijjFolmmH/4z7DWiaCytQel/Pg
+sVv0RffU3gywHLNvkZMB1xo3AbwTcvBUQSUCmfumH4yCR1Hw3wITFOHhfTVxJ/l+jDbuNiGjP9q
efKhksn3M+OL38VeomMENyYynr2lJacQENq98sx7MmvyQz1FOZoOfTdqwL9dpw3WaejDZ+Q0mXCT
BCp6Nmlh1akLzWd/kNTcczgtWJrzmbUlNA24NSgjPJCCwbY/CVYS1+cPdFVlpILgVZNTKWoWfPfl
ar0DChn1Jf75KAXr1kSOSzUjAkHTA+azuDYbBz6JEc7kb+7qUo/RIEmHUxUmOoAKscWEkQ4Yci89
N0sUEcMfAyvNIhlo8IAfEY4lLAX5UIV+r/xLwUHHV7Hf63NBKX5aMCV1Sc9m6rTE9jcErPDg31We
G/bZRs/M4YtJYFzWjEMDyRN0s995AGTrsEYA2dfl26OsE49pUCEm73Cf4kW3j0L5cbo4c+S4i4Dr
KpPUnsUJ5xECAvMIOvsPj+S0iFB0p/fqxRvx0014wle/c+Msu+V6xpWu2jQN8vffdaOArVjZTZBA
Z4z1wp/OZ6WyUzckKnRrBa+z9OqVtGrsebPom9xZOAefes+DYZKJqJnkPZ7Bw8nS9bI3/cyFYuuW
zBSZz5uG8Ecvhc4r+J+Zp/cFt8DL4qkxqFcJbbuuq/pkpEdDWSqRrOs13A5A+gE4nQBDT0e24vE5
Dr5Sz4iQ60Nh7j0FzqM/XIBZVqXS0W1emkGtRdXYmgSOiT+OoHbo6VoZt66AH/8b3kmnmRRpqxK8
TlN73OZZUVIh4jRWs+UAHhfWQBRvRe4qpWnaJ8ZKhvkA9O4T1OaR06GHHgl/OLRMrj/PY9pXwRWq
Hq7RmuKFm+Fre0YYLDxAP573QLiLiY1Co12hpaRV634HgtmOPaJkQGtMKhjeftFK1mTLAF1Z3oyB
apa4CaUy/sD6lXQbTF/IIXCprd8UA3MAJ0KznyjHhw3vzFahpdV9VQ+w4G/bmea+MzdCu+oFfs1P
aoqVCben7EmL3QhON8INWYYaS5Pr2lf7+gEgcl6yzAInt6/iA9Pn2Icy9hS70TtRJGfZdS5hcfCN
3JY8UUjtzkpCdCpQDjPqT7BSHvb0mbr2RsErlJ4wTE+ayUMsf5pIdEa39SKknSGZ1DwwZc4GNwvv
vEtri8GVm8zFeBiYghInWoHFfWzBCdaIjSMRacjWojoXgTeHBevtIvhfIBf5WiHLAXdB5dlhKNWQ
RZMYS16U1u615GyvjweXzkqpvn4SyREnFn1qT5CbFuIDRudcYIoS+RCgqqUl5nQL9yIgo7Nv0kjS
8vi2DFqGnB6Aif0M3Ld8/NaO/6Zh+C0uOe5qW1+T7dn2j/hxWoJZ+vloEHsb1NOTpwe7QQBsiv47
83b4WxGE2vaJFl1Ln5sNpzGYR2iov7vrQnHUfNTxGT0zPuoQFMIBO5OKFZROKoYfOsfKLUZbj9QP
L3vl1IKgl6+ctJ3p6zMdmZHZnq+BuwvNVISyAe784OGUVAHWZGfPDQjVmich9iuD8dz28OxNwLHS
3Up25uI39VHJkkDudEdqBx8uUqxBkXm3fNxEHNbdH3hISASv1YeoEJnwShuvm1aSdhROKboMkzDG
YDnkc8Vat/wUHjPcTn2M0m1jyv/cRGq7W6oaPdtUCL+PJWIb16FqYcIQJDlLb00Hu6umCSg+WAph
T9KOm3fs6WhdIjz4aY7heP6S+E1HdKI3Rs/1g9IXhD1SzCI0xEpCtAVaNQzCtehIRzM7Rtv2u/da
LVKtNQ4bjUSaYsT5f7nqcYN83co3RLw9/dsdWwG2jYqtBxHbvSYaZV5hInQBIbBapGZCuiAfIPT7
nb1y1EKezCg3Eo4b9EzZrdUIPpmInGVXLFaK2jN49rrN2lnpCSVeWw0YxbpkNif17FFFxHcmqnyw
2q0hQDIarPEzaR4lF0xb6A4m7QAT8PSpOJaW/lOwkoQFOlOyVgjbZh9CaIrQ8Kj2Hs9SS48e/ao2
bOOqA0MjC0vkliDHK0/Vzt6L6QB9wGAz4b4cC2UwuMVlC7SIoEADTMpMPiC4gEHsdVfsLiHYUBIF
QpJTt30ckan7f3bKC54EUv8OvBP8ukcjRIf9gryYqugnWVWgtHpPtCi/FJsPvPQYGsZD0qFVnNHi
2zR/hdguh0eH7L203M+IU1/vcew0dbRhzQo4KdTzA6+ojX+OhRq/YlEQDlV2SnSnpHh2k1fYrgUZ
qZYQQNyamamJiZoK/ehxMomLbppHB8HDOWiHpkxbCp+50APKZNrOlq0ZD7Uc/ksWuIdUsxQs7bpB
LDHBF89siDQovVbM7ENRwOZeNaHvQNYZB2x62gQVPxFBUfFqDcmNkaKeHvV9SJ7Vh6oHgQeAMLqH
vGTSCNYmv2BLoqIYCV/Amxcq7loF/BMfEdzLwwyjXw652bzJu2FbkNEkrYbeKKOltNUT+nxOe07X
drYnoEr+8qkAnmaX1KAlC+aeBW/0F2NmzkAQwXxHCPrFg+8YPGSqyE4sy04hDcQi3zKP2autXkt3
cuhBJYogYDsFRSdaibsv/l6DYkTwh3444rJVYPJyikZ39BetKEjB+gJXzZYl1iyyAq72KKre+Wrp
vI0+CvhrFlkKjtmRf5j5w6dXwn+MuUGAMxMfNid2eDd64ZZ6f9Y5d0rfHCOKqpSDjzNu9jGFLBKd
Uoa04orVExvFhzTScONkMruYaL93ccgSeC+u7F360kf/X6JAfPMwwx2I+kQTvEcZIb7V0U3ufOIK
Dz06GfLBI800ZDjD3+XBcw/F2mbfEeuZga319D1ZDxXlV5nqv0OF49mKPNJt0oLsCx4i6a0XPWgR
2a6s0lGvVEjRqLv1a59Jj7HIdNibmv10fRCjxAD11n+6hP4lpYm4XGCYPCBMCBzG9LOXZXkTGH9a
fVOsDiyofRwK0TjK9PImDrNyU7O8mlt+OR6F0RBBc+0B4q0irXpqgWxhEijLNsUeguAmJWV2GH6g
lvnbt9jKvDFsrCAMHh+SNGxaUXUYK9cFLXvHlhPOkJymYxKHiPYX4sWcnDqhUOZgFMPgPwFaxlmA
gaficiLIRwK0RXE3Tg/5xgKS3rRTcPdFtG0UoSlxiaVEX5qIBRdFSv9zax1tvbweUXyZUmwPXi5/
lbhBl/KcJukJRUzO4I+iWYBbBgq42RQ/P9u1r4Tf0OiqmyEVWTG7EXoQtNUYRBJOWCeI1ohEw3LM
x8olw4eIAq3Ys5qPe2NHZfODaj4ofBIlyFqOeGd9ugjEtMa0WnjAaeFpPgT3gzORjddkfvMfgOy8
+VLT9/LhFKwH/7msJBkbmRTpp0w7ASFy3aPZYY5ZIuk/treZBEQ5pjRg/qALA5/JqVU1i1PjvtrQ
K1wO5pRL7kBl95vJ5NJXbIonMQDpliIW74n2JmgDXVODuE6xxIPG4qzOtqyXFdV97DNLsijaZ05q
zVrjxcPY4tMqbVAmhLtG56rjcthMUbqZCjvORM5mMgoZe8zk3SwuS7bHPCfczqawFZlmRwatcljb
yy2Gcq43Rv2qQGkna52A/17LN355TfepqGT7QcZGM5VKxQ2UikSVBvqGQnp9Il4JNMXzXiu1zK+9
yl1ZgUuiFPpKslnusHBDT8KCSW9ONQDl2NLI7myflKmeOtFIPCg9FP4YkjetcOYnsM+7qH+97lDA
MJX1L0nn/P8uGXjNSWO9vkBiJ4lY3JsOshqaUY2LDvP/IiBpoHPNJ3+Kx05cL61Ggo1W/WymL0kp
kSFnSeEoX0FKl8dLVHCZIReqm3QqyQYc7FXLyqWVhhOCAe1R/B+yeXHxOClXmXB9w1qCzp2/4UKy
oCy/1sRJIpN/91hsO115IXwyfknlqKP33Xy18hCjS7GrJveguUhIxFBFzsDRu5hBvdrkfv7UnKgA
iFwbck8IMCVkNIaRnUzfT2gWwO811i1+OP1KFEq+6KK9o+XEJYzLMKgT+eSVn6mvsXTvY9qxFWWB
OOJvR9vOLaaKW5KeiH3gjc+vG/BGaXBDq5qbZySmp4ucsq0CJAxlTeFCrVG+bkX/vdQtBOyT5SY7
uKST6T/AUr3Bog8RTkHuUpJBvAcbqyRppKJcWBxSG2Cr8MYO01sXIMkHoFYJBkkIta2NizT3rnSH
1NoLWEzuWwKtDHuOeQhwBsKH36y7xryu6vnRYKgQjXmyiqut0gGzO+J3wTJ7gKeYv2lACVtHFAT2
x9cdbXXM56RaRJPSjQHx/Yy3/cB5H4jDwP4BYy16bvAS99L0cpcYh/D5yGjMIJZOcLk8GEYcN/CZ
44Zu+q5VRwJOJfPhqymLNn/I6imbi0pPX7VCMxGFdXM3fOHs9BdMjaazgo946MFxBe1/Uqy2I6nM
tQTc+0EAwG4cWw52p/GaolxSc/XWfWRv6cGQFSgv5D9c/JE5chr3Rve8GKt1up83YvbdldBbBlLo
nATRTaoiZl5DRDt+LB8nvAfxD6i98hg4mL9fib5md383Ng1wpPhfw7E7N58ldg4bxnRbPFTGlB2R
Fo128ix5McUUYx9FNXpNwi95r38OmxFQd3/fy0baj2KVbDINfCakZGqqt59NRaWp+TjzinH5ondl
u7dDPuYQn+dXiyqDBuzsmdWBtNPV5k+RLYIR5D8erwr6Ir7sJwK2BNM6OdPUr7OifFk1uQGm4Mx+
lC/3IGhlp8E6TYtMisp8p+Apyh9GRspCbb27tmHsmzbTZu5eBKmH7hXzZoppoIcNX+mSVDzMbq5j
heGshp8TxxC6CRWmYobVtuQ59qobJWtTUC6mV6mnB05hSahXN+M94qjZPzRblJNojew1DicjfnCe
S1QSUVQmEgMdcryCUFIruOGHwjIm+TDYTNyYwGesmY5V7HuCkBD90PElhOZ9sYY/dwpfaPeodlak
z2Jiqt87yoeLRk0Vr9XYUqdaD/LR68F4HozRqo/kDWjJinswTaaROcHiyjst8bLN8VmIDC9jwLBF
a98zaHHI6aDEKvLROvsgCXKTRZR35pQHyUvXho2jZUK9qsvSccI5FxvPixooIqx81o93yK15gFfk
e2ezqNLjqs++LdR3c15XZhMUfBApqQcnDdrmumlKMoknH/hFvdqqQb2cs7rQWu+Fa/HUwCPPEDlJ
GKTWvX/BAug6JifEFwUDrxZjuKaZYtutfCtylWGDMCUoG7//3KxqadmOwAOgZ+BTmnBJuFsopvHE
7FlHyue4MH5cQ5MRqFoJ+Qlsz5A/qjiR0c5myvnGEJ02DUeZpm5CP/sCv0Z/Qfy/wnr2noJx8r0Z
H4WN1VdMsgquwbLT/5AOX7reCEghPISei0BkNe3fe/1PpJdqibiDKZxhsjU2NSl2/ExKiJjHYGS6
EZjKZvscQdq0cAn5tIFMsSuk5lGS3YTIxCiIWaL6Gg+++TNFGTuUJT0cfCqMwcfLT0V29hY8B5rZ
7L8OuiT6bZDnRAW+RfQ2Do67Gf4cjNnv/ouuzTPN3Kj953cvH/wP2MGfahWpbPwttlidwHbDUBmo
kBnfE/8LeZwH1pDEWpS8QLa4ZBT4FKOjrJYno1A03fJF5l52ti9uvZB9W1Pqz34Fu+VS8aEFtFXR
fY35CodOpiHIDrXl95k2YUIa3DEGq5WRQdJkVXg+8+B9bWSxRe9yaK6rTnvBhyzvxSRX29VtHzkI
bjjOrih9wyGD9NP7Cq1AHyfGGIRXOdGBLrRxPlNBRpDbUb9MxBji716vWmvFrRMdMJKbI8C+nhFo
DGwdF33Mbav06QOQY8cy3hiaiAIcx0+ZWXMct9XJBzEG5jgSKkVVr6+mRAXgph4bEoVwodzh3yha
i/qE3pGocd6ZR4ZoMykhEJEeTzVfZPI6AQboNpgQxYnfafa9n6yQ8Ftoa0f9r1Rk9EiX9TlUk4zE
tWA28vWrwbdp2vHqWo7EK9hzhN2SyRnfGTSI/X/ltSMRwvKNc5/NDv80pG5NN04YOZxsQyyny+dM
HhsH8wZn89bZpU6qdFr53X50hUIRWXek6lWkZNj+MvPavpRg6kzL3EDxiME9NDRSlCBI+fAzM7Z7
k6Vze8LqzxmcokHegfxN8i9cOSc7CTh/ViIKelGl/yRpQTC9X53MrsSXPQ3MRzfScd2bRuTKTcUA
Q80yAjdxD4aFZx7PxqPN2bQFspyMPc3Qn84I3odWd9QB0+3YlT78F5cYmtTeewoyhRrnKhrU69Xp
Oezr2kxEFlO4/TuEcPiMubOIIh8SnZCN7XFPosYVDIqhJvyPsizT4tNtfPYHfgFsRUJ9GV5kSkVJ
U2cif1UVhAOcvT/GcKS2cT2mk2bc1l5/YbZGYFGXbs9QN86TcDG/bXkquK8cQhYmsZABS6vCh4iz
gJxjvauLHpuUjPCdEnr5kuTi9j0mSdDXtxuV3LR9jR6pcQIoD6FTcOGg5gB+HOF0Fmzx2TtXot9R
rn1/9KHgsc87hodJZsPdnJzvp81mItqdH0UMdhGaQozTfahvVIyYue7wwfiHh86Nh0zZSdcFg8r9
FQxvDhmfRns72l3OiVHSFNomLAOTkGBfZpk9cBdQvBExgZy3yLB9tttETK/WvPsJ4BJUvPIGOWc7
dmHx0QJkVNLAJj8Ur6sz9lEJxC7w49bJq0rLf7w/TNNMrVd0n+1jK7a2LNc/lX74EoH6++F7nuP/
lPYgeKOZp+IpoGx61wH45JpfhWbYvP8ikTz+iy/lfKVkWIPICN2HkJFC3Anc9I2XOnbOrDgdEKua
+XLJIZETMby7TQbM9li/SBygs5PWkSAbuY8ituu/Xj5OK/ZNyQXosCX+qjbJ5PeSt8dTsGBS8RUy
2CmaCfD6agYSZStpgg70JCiDCELKNue+yMQy7tvBkiaNZjjdt7LAMjpNBHx+Sb6i/E3xbznAfiCB
EKTodNguWGroEWbWEXYW2lep6xRN+M4rlHu74PQmUy2IMYpz+StHPB4sKthg9ZcS+RgU7sRpFUJd
ObLZrCltYo0Yx46TGzTkfg+nhGVZU7VJxK3FpHWxMW4UwNUzC+/uQOJfsRCXzJ2q+C8GdURJOOiA
mVDaHvhT/wVEdhUDZ2pWodNkXf83K540H6mVb+sTm2esCIrKLOXI0rYO3puLlpSoSV/OSc6KmWMe
cM6kh7V16w6cmf4KQwB+AhbdnniNU5YybLEsz1mVL0RuVPQtby6sJ4Cmfz6dy27ucOR7qCI0kpt9
EdPnFvBAq8Ngh80Ey8Tu9e8NxInlBPEJP5oYQ1WC6a4tLHTUWfOC2zWLTuqvWlwi2PGnKZ2ewsYU
vsZnXEAUV8anmyxEbrOVuMV1xZxmj8395z/Hssbc+IMfgL5CWOqkh6wZ6BvoiWc9te7/D8Q8FGGz
30MaDDnZaqm2Al0EjMJ/as60KxU8U8uuMTBiFQd9sDzn0BzvmfsEGMxw1pIMb90mlmzEUxXlzD0g
zT7lNnwxykS9z6fa6IFxXlz9VtCmBv2XpXtB3r+eWUYtPTpaDXGYxU8zFemPzqNQrI8i+KZ6LU+Y
6rv0+orgeYzlNk8w35LrsArFEvW56fqlpUIhdxCF1qkr+ndHvo5SNmiN2mMMAzHZro/FCL98ckLL
nuHsLXmrx6RCgki0SvZbACTmRgpdUFNywLpVFIj9EXwPvS9GilyWGR7jkeLuOqZJsY2TigIk8eu+
hg4nIgD+48vMy5rwT4RGAzSKILh8JgkWkiqdggnsS43xj/N8GqY9lNpMrqaqqGlDcvXDCS6YnoIb
4Q7eEOsuXC28fxjqCwbsg0cjr2VCvRqNZIQTUjjSY+zFkUuCigqhwnRJ8WBCWqNZDUtuz4ifwXWc
caWWInAbo3qRF/AntZtc+zkA9/AlpRnUxSat+/pm5RvyjAZHkoqKA/NQkdnV/rCvrOudBupKHdBv
5CfYlupOlahbgJ6YNd/4tL/pOuLw+LfFzEzJgsidi6lSg0BUrSede2T+t3UU02wdgQyg4Ic1V2Da
B78inHrrxtaMzhnHHASkICE5mEvhLWBagOQkjE9F0ddvZJwF024LfEWwwcMTK/4gNF201tJklTTY
c3vimHU3Ev025NhTudcN8fBtT4SLKVKAnYzzS2hKHq8wztiS6SlirYJBHFXhGt6hlwLPLAHd9yYy
kM1t3iFAYotjljPKd7/qiRQrXZGPvLoIw83JVH7rR12AK2ticTm0aR7dIREjxLsc1RA0n7T5jKAu
RdYeZtS7MYOCdLXUY9QJrrwpO/jUo6Xxy6DeS/AtLjemaMtCgWLS32ZCbYzhFzLmjxydIlhFzPNg
ILJ0+GkYL5MlM1LNvlRLUaVTfen4QwYpHaN41l+rgBjkh76Di7JTcMGYAmGhb3IRFjdO3B9n5oRZ
h7IlpFrPsG4WsKu1x8tvn/76GSdy2qw/P22LMSdMuQG2yDzhoeZxmilQZ/byNXZiy4XvNAZdInEx
HdPL7jsKr4wgaHvSD/BRzxTmgUKfZOavtHxQG+atcaxZPz9nnlI9u9yK6B4jCZ911ATK3DHl9KxI
td2LqKdnqsqoLo8x5t8vVvR5JLcZa5NEb+YVLTqQ8uf6yGgtwog0ZAoKMC8JHO7g+GAwd882JtEk
B53OTrQ/i60kUwlg9QEIbF9lkFlgWdOIkcCqXeIk4aWD/56NQABH2a6w0Rjl+vtDoIh0gf5pwt6j
MfPBEegGyqoApbM7q4Sh4ERQpkOckG7NQ6hIGr+4d99+nIIE0hoiLo+yODSQPXUrlf93Kln0MR+P
34wM8jCamNwmcbhjBZmhESFqxRHbMgbPsVjgadNovzD+TBEWw9zPnPtVgplpSRMQ/TIMhbtqC6F0
1cwJV3Mru1jmg8FKubA7ZtTOLrMwCobR7kqZB65ciAMLCYacgRMC8Fc0n6bzrM2jCs/UDQVrw682
GgjdKXgbsxjnyz8IhAu5epI9Vb6ahUpDt+Sv4WfOhouiD9uZNs8JeCyqhHNQqbBTzgszjNhIdF25
stQPVEWZ6AlKpuMFtsB8TnGxHBzSs8LT5865KSO/KKYaOGGwVKGN3D6WQDota00VdeFO3xoI47N8
TqofMWRGiGq3FFBw+gPN4WIBSiGI33QuP0W2/BEKpJksr/9HR2pUZp6ifE75rKJHaDFuCw6huZ16
LxTs05GcT+2/ZjcmbQCkbSZuPhJOVDOtEwDiakrvVkobaTsWWkn/iPPm76cxMluGpGBGMN6ul3Ju
qcU9ibyF6DplatiV+wRoe6UmEdhwd0XuspFCR3NttMdt6Cb9QzzUotvbvDSMdAP3O8gPSnPtRqJe
xGovf5VY+gkRTRXUHWQoNidlwo0CCN1YLBlPXLOcxMLmapHg5FFgxsSfNQNAKKvWuImsLx0mLTZg
Rpn0Wo6ysxU2ILNimDHVFcNzgd1hyQpV4LPiEEkYa+ubS1iy8Lp7eoMHS7q9hNckSl8TXxmBWBU1
Iv89odtyzhszqDKm+b35UAuu3Klwcxv+TFzwxVzAnzz2C6MGtpPvnYH8BQxzFyniJ275owecSwwe
T3LUT6J5WHACCxBf+HpRxQmCvSLVp1FaFRXvqhPSbA7PIBLbsR6ntbZmdsAdUVth1Xitz34fK0kY
ZnG6wjhlDuho9wp0Wo+HnjvUM94DidHreAUiUFVDxO2uNoIovKpDEWFNCLf1MG06sytPD4UfXZwa
hC44aQ/frW4jIi6/4paPcYhAxEIB1QnRnGwKsvU7lR7ffcn7S4HCGlDdasSJooFwbdCpKyud+xvM
rMt0zZwMhMlCR0jIDKM8Jt9Y+lXjOJFkf4DzRiWgWilbKyNzk6OZ9YQDK0X6RIp3Y88HBLV7uV54
c4hNN2JdkjjdEk3Jt5RSuqvlb96460zIkbCk6qMmtq8A+YM68i8U6MDyAPBtvJ0dlnHH2EaCdVqD
F3tS378Yv4PVRKBMLfsQ/ahH7b3HxQC603DS9OOY15D8o/6wDG2Z3CDhjqcl+EJB/dWoos97CsqZ
ChgTqRE94javnWBoqR/i9eeHLoxFedE9xlwBTZThBaXJLJwdVDlhaSVjtwXoalDXjdcKhHMa+KnC
ZaT8bmjT/2omuNZbTYi03ZeUJxeQKT5PbxwwoRp+JK/1eS2ry11sou2wYwKJO/FLVbcFZ/5qQitS
nP70IMqAMCaUDjNTQN0P5pqSibYGzVu6sNds9sZl0LEg1g6cwYFIXy2N4mQYzqfCGU0rQyOJgw3P
VA61xp/S9qX4MrOgIVsHQITfF5WVoc+KOsx/ko3F4v3NLpEW1R/Xdep3GHICOOPAX7MjeFQIAjQS
EMbvGMjBjXOD1ZyQbcwbYqGh5w6328GstufNLaB0c2YKx/bWjSl75XHFYM7WvX+3kafn3gwEbpaM
HnNgf3sZ6iWemgifNIXcyrv8XZw5QSJeYIJEWMIKe6mQa6GsCG4I6iZgQHuTsLftbTnUuXk2mNc8
7SFtri9JcFQrVsNBsL0Lp4lw06s0I/Zthq7QKuMpZkKZ+8NvLV4MjAq3llZBRqrPYGWcNRKYRewi
koqb8WOOi+vl83qDbGdqxYasiv47pAkNuhxdUgIv/xNsCoNpRqyj6zsuCzkCO6fuGZbkmOG2Pvmy
8RTUVHFo3rD1TxcpywZ485RKhorq3SGRo7v8GHTXsDJnRtbjAZwXOyiy5XkmlaJygHZ/RaDtk02c
btykY8EMCV5t61W0OTCJf2fhuyTZFPNoWJiPVUI3Qb3TlFouJazA1SiCdT6vl7m5zQysU6gdExwi
WD6rBOufnEyx23YG87AlKryvf8kf+PunvP8GAe0LB4iwBYUd5L+tXXMfz207+HNy39WhoBniwe0A
MmqQB5F1yDQq1bS1qq3nKPvDyn+ZG2FmqC8UCIVOXQvgbgV2l95sZNS18i5Be7qsEcXPce8+FBpU
rBzE3WQJBvv+IrOb4r5f8RiHxJTdqNU62GtFIgzaUqOYe1/56LT+DObeYb6zxN0muOn3sihRy5vT
0vMOTF2zloFHrbNzU66A6HHbl9d1YnJAJ5zXk8Bvg81fBHg4WUClHtad5HVwTTmKglAy0BlwfPNT
vXM/GTgkWFBcec62YOdO7LB2x3fq9O8UrwQbX+ncmDsf3RWosS/mdHwW9XwjeB78AUR7iMBSFxQo
5NwUfW5wR7Qh8bql9gXqx/gNbieiXl7BiKep5z2bs5t4+PTZHWY58OQ50rX5+iB3sgcNAkowZh1V
YRH2YTAanagKkcF6EoKUWWWk5FEgqFh/qKAVOHKI7fqmqPMZ8wIEsiW1vXRz6ZfOBe6Sic8C9xy6
FY99WBaoMiGV84lkcCKIw1oc1vg5wMWn/y8e6IiIkGT0Uuse9tbx6rz7sJaCflaKVsKNaSZFEnc5
1AeKqvzVguNIm+Uom5XD+yDkb90O0FSQVMii5uahIm3zp0T7Z2Kb9T91+oJSGwypxwvGpIbCHLll
oMM7TbBwi8IDfmLU64wpYP3CuhoV6yzYowkoLCsv96sKDRhFzSgsQqB29xFqeQ30lByT6SumPhWC
7pf19R/bF9z2Us5Ma/MzUltT9he/zSq1fhQI+cdLC2hIfZHfVDcraUzOlAxoF2I5ogDjFl14UQOq
0N575wNf2YFScZYjSxmxiUCmSFRE2nYzyu7pM8WRtmw1k5vOWWsjpRvI0dDPGTEMOYEJInFrw5vS
8wPpKjMXjqXmSvjATBS4YDhHYjgan+Hs7bwwEvAW/6sNBuKOrP/un22Q650m1H7VyFe5jK/6exhZ
alhlbMBGKKfxgw2H1rQdNzZxE9CufaWocCFdXIEdsUvnfsHuw0Wd+bGOmq5EAXpIbjYdPi/mdOrY
cgv97fecbJWFOHxx6ZZ/zQvSBirw1+RAiK49kPMoUdp7wPuVzkAVUWYPBFxKVb3I1/IB4pBbdbOI
7RT+YL2PSclZlBwyJxN3vWW4a1xZ1hcInQB7g1ZQ2o4qINfwEICU0fzSzApCYv+Kn4ycPpJyshtz
9boU8W4hTnhhSjaj1xT+yiJ8c54jv1xEzY5x4OMwm28afYCe0ecf+hbEQB0ESqX1hUvRBQtg8vDU
9YThonYClOp2Tlup6HTAl436KQU+/kcsMUPmD0RpuoocMNrCm9x+TZ7AHAq5yKZuuvR6VEBbc0iU
p+tsOAvDSOwPrdsFZ5HGBZ0OhkG+oWyDr47YHLIbJyotzJRhbVZcX8rpGEkc5yvIRSQbhsFuVGFF
+6HmLWfjcdzDNnSO9Y9oD8FvoibnMNKopea4tkBszpG3QW741ygMDdr5msjzXLYa/yZeZEUj0b67
/xi8F58pZjx/0ImfoYRVmNhU/r/rK0PYIYbnaB+nbk4SroflB/aoR/gs2hoDABCDFCLpiyoOepJ8
OS2wzH0zPlg1fJZgA6ysH5TzggV/xl2KjN+R6hKc4M38QvkGWiye9pzOHHBiImpRuU86mF1YzHUq
3eE3BY+LpyV+W1dNM5fjADRl/9xOdXowA4caoI1qkIUGU6e6nLXLrlHXTsnaZTbHN7mLfuy4iUDh
9isuLZ4u+NqjKfADLt7r7uRiEiZvdrnlg8LSRFo4d1e8/ShmrPaAVapD8pLjn4kB3F8X+5/46Oy9
uMxTaJLpikSJrGPwv9qzK6pdMqKJJHYCelb6dBaANyY18VCOHXu0O+K1zt3udH601jDlW34UkQE2
FxmefGikcJXKtluplg3UdpCDFY2OenB0BnRFFAPJhsqcnvjQREtjbD6dnaAQfWrAgOipgKA6lxyq
065TU2h7dpvbjAfTQ7DLW1LGfbSLYa0xyNlR6jukJZshJsNT2FXBBrWdmnvQzuMd0oO5/WZueYId
MJOS14F53FSdU4f7pw3iJ/x8ocM2NkWqsAg6i4ks5ZQLpTvXy9JDD069P1Cl1z3jG2OfxehPhKX/
JdonHSC4e/w9WP+GXwE6W6c2WKBhz9IwSYccV/Fo/qV+S32BmZSCW2dvAO7p5ViG9mZ3zX8ClwV4
ZBC3I92HBZG1FtaeS68kfSY5RUwRQJZb+b5+Bw6IgDqPl3u0n+DQeEQwRRm5WpsLOcRf2G7sl/JD
sG2Dl9234jB9KBFF406uSSLtbBGWQhGCk5azLuyQpo7n3gIJNL0ucATRxDnOIeBrZeHJfu7Yefni
W9fZNhnIS41MU+tjfgf7tBzg/JOJtxZ4XCgMK3HEjt1Pq5SryWp5r7bpRUdmeH8bL/10pjgf4v06
Hup36kmmmJT3qvh9dUVALc8WnLynAUlz8jVYhMmb1NxJqcaKiFV7U2HWfzKFXcX4G7sv8ze1Bny4
saU9ERaiDEEtBiIiAF4ybeWfNgrgM68gLn2s+0ZtLSKv6pYAIgNtLLuxgd+Gxy3jJR7+NcxwPPr5
dshrZgIxG+UTq4gARloqHFv3Y9vmG6K5nk4+75NDlkhtVVi3cuHQkYDOGFR7k0+m7N3mLuuDrnAg
QS1s66suXB6JT9iyb8/WOHGc8aDvZ3Jwu2Jl2tuB/3yisWodl6Hz6QEjURMMxnMi1JaS0QWLZqI1
piEmtPm8CQNt2KM/bq+xEzIjilhRm6dIO/Jghe9gyveEWlTYFSDw9Na/1G+GdEa/nTG3sWh9VqG9
RimRj0yxF0ZlftYXGMFrGzffAzHo96GaojkA/RzM+Wd8Lnlokh3Bh4HWLkrMxnc5/3nF9xy5BYDn
hIxNArK2MV7z2YvwNrW4SLl2CTjoTvkgGjmYEME+lh2qsrqydxb6YAWoIArkXnDXOCZUoLd0JosO
df3kBgMoq5iyLt33S2raiA3QGIngDQNF0ND22mUcKnSs3lrwaO0ko8TRSUdggxouYz+seqK1Ipu8
NHkd3+lNE/cxAvbDnWDtfiQvAFsqwQbN53qoqU1AHiGrv3BAFK7Oc55h41/aYe+DUnONeSwZxvgf
7TINqscWQbqFPiAciOHpv+mbOjW+aQ8YTUJKq6FaI+qMD3vQvtHbNEK8GqjMxjgqR5ap9qfUZ83A
EtY0FVz436sMVaP47ytuvDdexkQITyZ8CBXEzevMV8AByyHLUban/vGJK/dUlw9p8503XnwYK2he
nCGTNOUzjy3GexLS+LUkng7d5EkJElyYBJJc8lxf8xNnpQHVuP8kEvxRfU5lr8j6dsBbit0ngAt5
5cTeIUR5N4CbDQpYrFlDcvdy8F1VMuDVCwQEdxs4iI11s+IU4Te4mhXnusBuUT4ee54NXf3sjyfA
z9IWGNFigPANdtTMy52oP1OaT/VUi0+nOVyJ4ywUSAfXL29snFmS+81yJ9ssiMoFZJGcNxxZ9tOG
XVD9Y9qaWxAYBLbJt7cPlxiwniI2rXgOOZz0fqZcDWFbaC9C/AEPOojTawoSoTRA8CmAvM4uaK+n
xaCFxlmq9dAyuzbmC3VdYzq6cocC9daksPRz7kF2gpqwx49bB4HNnPtNbZsFB9YvnVSgZ80QqmLd
hkUNCPoYAy9iDZcqESCVX1KsDqsMM/N3yDfnMJg2ahIgrUtLmTOMV4AZQYelK5y+A/N10L0v+h5W
rDKLnMnm9T6nFDRCDpQQWb/JfdCj0QfT34L5SVoyZWCptUD1xENl6IMgCisOu/aSkeFuaqA94nEF
sH44VtWUaKrCFaqcl1n2jwnEabQyS/5wFJYTpNWJET5MXRyjhcswpQREdQtXObVN4UcLCQF6UTj/
kRSllytq66zWWK4aQIr24Knbwz4mZwdgHMW9KNrVvU3+o25TmLoHlVeM3K3QQQ0B+kEQuCi1cxGB
4dErsUZeonoyNhOa8E+MeoWfdW6kp9vQSbUwmEjsEKXk3AFu+NwE/Cq22uZH+AXJIUvYKKVAYSF/
LVxn7Hd31+9RcKlXtK2bEhcjtsG6QLl5YHdmcnnOQDJqbjDEddo/4IpmRo8urJHFuwlW/dc5g/YA
NNddg+d9VYDGq1HQXVi2/N4cJp5sJAjGUifZhU/jMXGlhLWZ2Ryz7KqaJbACDNQa2mOPQhRk1qoQ
ulpwBBJpGU5tofWYTOrT7QeGtY0zqQQ1y9zA0YTvhE6vOpJm+ADHd8UZvYHZeOlG6PFGcqn8sHv8
f8gv0Q3MnWS5oLLenSuHzTJjlCSocnkysb7T4LS4WkvgQibfBFVl74IGRJepgMod7xhQ+mzdBtzM
1Txl/plGv0wjEKyIYQs5IhvcoL70wNiE0JqXCTsMWgOZPbpfmybmVuj+9vUztUlqMoapVx9G4iGQ
jqxr4rnCoPaIlJavGXXVnkZX9kJXKqqkyXy6K3O/nuT/lFPTpc0zoOE6Wp0P0Me26BJNibaYAmjB
JHVTC+kLyPJOXZMPUyGVeLFNX9CYs9zOM51bFoH3hrZq0pymKmHIT9QgW1veJ9M2Y4d+kYQBYcU0
ds92JE+08qHkPjeL6AY5xL2Epe4UGpKkENbqvObnOvSuTLPo6idSNmHaVaJi6Gt3JHF3X1Mkf+s7
GTKRbQJZNzZjO383y4Eg/bwgRz59ne2wWrF9yuJv7s4GjdqOISHC8QUoBIpLLInt5v8/MJYC07R/
PMWY6TXMLe34CRQzanw/cwW93maYGWuwXOpDSlO8DQHNP8AsZcGC/D2ZwjU6ybDZWZTKup/GiOYc
0krqmxEEHkalxkIJudvAMa7wuNaqS73GZufZXcyItTvhyEF+qU7FHoMAPpc5BY28qruPkIbWh1qf
+kxT7zMXw9ZTSoCIL9W37qMQ8es1kyo3p5pHvS3bMDya9t4yi+T/fgQNUxqtcccJWT0TapR4Zb9K
bgeCks2fhCjiuG9C4YSo8+utasKz5bfxER17i+e/UKklnM5PrX28Bm4UntSH3PcIZndA/V35YAhe
+i4jGpSURt3ATsJUtvDp+ms6oq/fDUlp4ytB8ZCnpLUXRIGGBLm6D8mNvG+HNLdXTdBVvf/5qQey
ZmN9UYyd9v/TS8bD2AKDxCcf2dnD82dQCipPi5sH6P1F+7eLPo7cySsOY1eC4oMO1GVYnoz8hsRc
/OW7eeRr4aBkhRaQ0lukBNFEe3hfg86BGZziS8TnlA04ymPE2+756e1yiw5qW/v14Fz+KG1uJ4Xk
M7SbcfarI6ZiochjjqJX6nmR+ADiyWG5Yk5xs+mSuzRnWBwSzWD7GO7JbbBMYT71Fw0SC9pUtzAC
53aXQtz6Jq5QrWE6epcSRY7yGvDpzF1nCIbDixKkK9tXnR+3ICxFHvy3ytj6smnyBIclRI0+kq55
3QFVibaSUKtALJjZMAp/c+weLn5bZ9Q/GsBmR3C7ucQPJ1s6S7NcVpik6pWm4VUdu3L1F6A30ES1
9/jJwlsNEKaIpLQm5m5ch/4VEj1FYVxPSDW5/XLRXCohTEgXKhDuEVwvSRwN8TYzgUvjxyXHa29g
f9BJXhmqDhHSLiNgJ4SbXN174cbCtDsSyKTPIm2+DAgDfM+0IqZPU6joDBD4jh4Fh+OiAoJozVNL
n0AsfliYvKZkzOw1WaIAnyORS+wdpiDm+UCKGOnW8ngQ92EFsrz9J8BE07FuyQ50cPOVM4L/e+60
rv1NYQoaJv7bOJEdn3QDMjXCLcN69Cxh91LQ36GJAN2afhUhu7thcBm0pIURJXb2ZGiIRfZgPZTP
jU6AnylFiaLyd5UoZ4EGYUhB4wzujTFyjCaTSgHk9Ev9m6oic1VMkTIgBrw8/9Obuy1hK3mHuEbw
BL9shrQMHSeXobBg8SOZt1w9VePk/s7Dz0vUz3is9hp4CeUv+y9lg6cQNjAvmTJZ120KrexjDIyG
H5mCeffjJS2HIfnNmjf5W3LwaxL3YCiPo65bpsBokkLMSsCpNvaHYnlEiEY3ySgNKvJC5MRO2pg/
VE0GUx0EoSYUCKUl6SHLWKUSIHx5io/DdFg/lFLj8QB+QHnxYId0IMSfSDyJavuqhfS1HTipYHw0
AEvi0nwQ862LKzqoBDDp8p05EzBKRwQ5maQ+hEy0sqX/RfRFL5fJEMUytCapeKUl/LZDoQTU8HhE
UDOWJzZN2uwPZxkYPWovHiVnC+TIFDnRJtikE62uoNIUJW58rRc0sTcXSKtpalk//BaBmzo2+ifn
PGxabB9yFPJfhtJp6GKFNSzvf80lTc/O4sDhO+X1QuRqyyyz2tVclPmFulMqxYKIOdAbyV7aLLmp
pTa0/gTwJQHKW4CJbjmHM36CmgSC5n6bT1XvtIlKlKi9ZrUpKB8tvQ/WUTS7lE9JV+SlX2Eu4SPR
83e4aDEcHbu+TckILb+z3/PQE4JcTx+KbwzXh1QqM3sL4qX99ugYJ1HodAXoCbc44gXkoOH6Lf36
LSyWE936V4Rl7jsXV+f2qAiBTIQg1i3WOG98oYoX8WyYNdmijCSmPXLvmB7FIZUYUzn0ONWrFsOn
JKHsmkJpEzvLLAvPZWsa0Cr3wpQ0hIFCrwYrBUDFUgXSQdtZ8kqAVSyreBZiodqSyKnmEuNWhpjg
heg3VsUtoGzcjZHBIfQFbrFyZsMBxu99TNhJ4CHZGoCJeH30rdyEd4mzbteS58lveyhhg7w8wIDb
Pyi7I4FQ85Id5TbYDM0kHcgxQuG0AgcY0WoHZj41OPhCtuvE3LseeRVeB/rR6oF6tb8/ohfkevLD
4I0fzCksAsZBW+1WP46VkIzGwZE6x2qiSB5GYr4xH7Hy7x+7vdufM3qzzSrJAYBm238hv11wfRv3
X8WEpCkkc4Iacnr4SE0jF7CjUgk4C3f4CBpqD5F4rGkimHFMIjLWCA2wLM59uLxJa9xDXvhz77av
zySiKpoxwsjwip4drlGJmjhc+4AqQvCzhzF9N52DoK5r1Gxp0SaYAd/cVc5fu3/3oVHmGOWMz1vO
acDUj3pUJwzAD8HxrfZG/1ZSqFF5GLeuyhAojsNP+vAt6cGOhdcnMqlB6wsjDjCbS65IQ2f8Xxfy
T73nmbRn2/WPlRp8mQwUtHNftjsI2UXWZIeXxSWDonsODzoO36WsfOVG1f5wDDZ1jvYgbuctdl9F
wC0skMJxja0zmrzhbYIXwPZBjgLMbSfEbuad6xNpWSLqMdfzgfYduOsqIIiuuZ1SXJp5MEtV2pnv
BtSAqTX0Toy2ZETy3016rYbuHB0q8vEB6jhRuJZEDUqkNgjQfmJOeIv9K6/NRZSpaCpO3p1HmVGz
RZB/rhYoZHLTO513e9Pm98O7rszJDLy89ClNTGDXdhlSCJEVtmXV5Sr+KD+gjUc6yFZFR+f/uyrN
cSBmt/tTW7MnvcHQuUgslNfPynVYcDsA2SuclrPWM+/yKzLjB4pydi4mmV7zp0esjZlFEbAc6kQH
G8oA9APcf3ayYdn6fBewcyKUvh2sOtOMnMknyOlxZp4zN5j633b+YLd6EOrjjeOIG0eFCWF3Ed6Y
Nt85JCFj6Q24aqb3AmnSTGAZesev/sp+Um559ddjyiwJOyZa8QDF4NQgaz+8JEKPX8p9gJ3nDtw7
aI3uWyJ7v1dGGh3wefxHxndqI3z6fozApfSqxLkDhSFzyvCwbQbxmwJ1ohB6RYcxGB8dZdw0+RjQ
IMgr34cSxWax54QRRcdDantBVXwaHyCRJ96wz0iBjg6QzY49fX2SLErZDir9YcmiLTG77NC0vJH3
nhRHFQTBHusnQtgbifwTy86eVT5RqRJeexS9nJ3+zhqVN3ZDezc5VzZvlREmhvoZJnzw9WfDneXO
KDxxPgD4Rz34xyoPGQ34l3N0L2EkCon1x4aA2ALX0l6aXd8tpAfJX5ETIaADvJSmfrCkI99LSRjN
A5HiAe10NKGiLC6PiDOtE0pv9F5xcj4oi6Gak/MuYgdlJ8p2cXTr0tukDF/Xap0zQB1uGfnmJFUN
579wWOJpm/5MkXFrwGO4J8EPbMXUHnLPIBq5Qg8t91IipSyDTcq6Si4Od43RCNHNW/AHkw82bED6
3uSFt1XrdOe8iVcN6XKHZdvHLNMYE4XFFPfwMb73sNFq5n0V2a2QxUKkZE0tVkYinJjejA3ZwZfl
4nNcQTtY+DSlA0hrvZll2Tc4llZ5W0alWAJZdaCPtxBRZ/cBEbWCOKABtHoe+FU9hGgiLQLUR/92
YtQEDwwb2SZdDCWUZO2Rt0jCARNj7Uf8cSoHJlcL448d0Gi5aE45MbdWKjQNJtW0ZCqUs1MarLGa
dC7M1XgFrYjUxcHZfMQaCMV6Socyo3KbHp0rWOz76zRm0uuXkuJzTR9DF66/kf75mu67smEyWmEs
ZLhDIocCOWBYg9CehbpYFeiW8zZLT9s5s/6nQCHQpVJh7RnL7bARJM+NGHq3j2BcBqI/iIJr7E+B
TNpMulpqusE89FQvkDTl3B20/qefLrW5LbrKpbLkXgt6qUe9gEUsrV3Xmr2ir1YYn99DbfnaLG7w
HvU9ZNP2Y5JW5xOMRjiTB/ZJ6TlOa7f40ReTQ4c/rlk9E/r+x4yOGcO1CW/t+Z+3EqxS0bAGF0Px
22US8lkq+RTfu3eim3Mhb9idkB9QixqoMv/TDHhy64pocYPnE5eCNgoxJcYNXW/hmvNnh0Wfj2mp
4uLO8V2uiw1JFhfcnzSa6WXV40m5n1us2W50z9xkZyAUKhk1yaIU8HvVSlDiqqAVuq/xGQzX0daK
kBiH0fOEb+I05Q+k5l/+WToJViwRVqVrNoD4KDl8SJ9a0BPPobjf6fgZ6VDKjLd2D0XYNRTNJ23G
6nmIuoCivdRzk8iWm5OY0rcgJBJvSt1kepNcLPczvBHyRUvTx5Q+aRE/I68zwt3XoH3aO9A3xi+W
O8HqNSlgWi4BM/STkj+FuN5brjg9W5khuD/jaFeaXECUhgYt7iaEhO3YFGSnt6icpkAzA6OYUHPT
sCsQ31M52XSd+qTzWe0U052YvlKbkMokvfXPxHsRuxpT21za57IMs3TO4qDcxtUv8ADAr1+1pYr4
0cGK9+L0e+t3h5W8wz4q2bmiTPG74wDeMAZ8sIvR6qyNFUxpjJ1ftr9JIbYIzZuISBGLsTezBr0z
Qp0UmnQYkhq6KYSkjgDGC6D2ugkboGQsMQ+3euNFbvr8OLUftdg2GxOMN3qUiVg5z+uicSe6kDR+
bXgHGjh/oFWPQrRV3n7oDuXFcREuwUIcC6B51xCB7zOQHdfpXxh2Y2aPsF0rZjpPpn6HWd95DEBn
GMe4/TVFhb2RwNSIGJfgXx0QLtuVk30oS4dd9GlpEkYGxeonSQXgvbEQy0KpjyNbRvA/BZlJpOuL
k/wIus36+Q7Qbzp6AvDFcl1f0GJg2V3ldOO6rHiASlcQ+kNDA8AznQ3edMHTlUu1L+CMrjkS8q69
OTZivmFYgH399/rU4imRPd4EFm/xmkbfa02302S9FgDsTjgtBj6QjfoCxek7uWd5M0LSwBGdrnZD
Z4ddFggIUdG29ut/1mG9UoKsDGzoEzg655GbGFKC9RaO7FxJ0eSQBtq7hWMt2F+Lme4VOaxDSXvE
9/cfz/8bB6Y5KX+EhRMf6qZBuq6riyr5YXPcpDPj8p9jwnWJsiXLh0ClqvgXTdOw293sVc3cfOyZ
IndOtUmgxZ4hzsXCRHakP9BidCQGv6XzjtoW/N+Sx1l1s5gZM33BqBD6LlBudi3M2AT5PO0SSCVi
/9Cg3hGrFPAEXcepb6jbUNIHTbC9s2rmrvITjlTYrNP980VzjN2IIX7XE2GSZZjDULCU4Oa/KjsR
AE0qm8W1GZZ9i5Tp1Kg5yCBF/aSZ7J5YN7N4okfgKlApRxU2CKFQx7NUnfEr4OCpZ0WlOVK2qtcM
5NO7HmxGgZIv2zzyocU/E5B5BZ5ovtv6FhxsKawBzQ7EIX36Uk7Id3Is+mIOCz3Nt9QYX+lF+sGD
GJEJJD8t+p8bF7wXTX4por2Nso/MBtdaVAlytP/+NcG1PXSoWbuCP5YEQuWT3LJsI0v+ahKUc8OP
elJH7I6bn2cyfu0LYOoyKHmDPTKmgTIuDMH6unaR+PHpuYZi2rHQg0mp1bo3t7+8tMAcy5MhTMK/
PfU+AVFBlnc4fcC4+GUEHWZFvijgi39FXkDVI670j2iPgaX6ugVFTWRV74Ge8eGH9+2zbuXhNzFX
B764FLi5zICqiXGC3sy4KomolS4Nk0ZiyOuChSMkkIHDM49bR3CvZc9J0O73IudJZKOS95kHq0nX
z29z+xWjAs0+lYTimbhRuA8OMN9OTYPKeokedie+X57Iaza6Y8V3y7YLxmcnpIA/mkvqBudoZYaQ
H9UdSsVgnYH+/3RJeIyceFSitWueOhzmn9U7g7RWET0s7jMz2GpCNSA/kw6zSKKAUrmSHVWUASkw
9EuoAvKG1/fpujmxma3WGHHn+NxhQVfWRnQ9NFLm0Q5Vt/JLosgiZmqoapgnIjGLq7EoFDLB1q/5
3/R0T0Xhm/SJu49wQ+BEaJrA78exrUr6sNq/nLb23W10ysUDql6kMstT91tYcZhqEcOIgfkcT0AT
BiMEvp6h6NzGodVw3pd6M9chcMZxpdsWU+MOLokc+xdFrY4IBZVue1qh4zfqbT3x3TIfb+fyfwKl
KW4klrVAg8Dsio+FVnL8tJiFI8jhmOjemnfxPPXt6/fSsyaa6uVFvgRLYebn0BAX5msnzAZCeHbN
N18tgwVQGKx3BTae9S0YqSTgp2OfTRe0bBhWCDCt/EcrVYqWsa8tjsBOR2LAgFMa62gusXy4ey3b
I7UB5gsTM4oJCNtVUm8IEhKLZZslITQe+pkHlD+aGxiIdqUZXRYArnLdoWERiHmG2eTlYJYgD0tj
sl2jsBFizfvxK+LX/WiLenUSIb2Odf+iMDYGcS+iquDjW+6PqbCU5FOjaMEeSI8xpAFrYZMuVTy2
GCCYh2s5cWQ29Af+SUCFW/LMtqX+uI1FioYF4dOjGqfnDl7N8/lfaZ44pOuS+9bypW18vFy7N+aX
Yx++YwUv0xU2/xmn1g1EL6NdK4xE/iKc1tdbECn8Ma/R21YRkiFDbChlQa+9+9WPl4kysISS2ouW
zi/svbRK1CKvbV1Sffb2fH4a3MokMHDOGyrhM8AFAQ1DeC+uj3kxf+H+tfXMlUSVcffpGqO2Zfi8
+j5z9MVhVUyky+ffLrZukmyDZetQJBJOOpmrm8oEJGEChAIV0x/fObjkD6Y8oQ3j5XGGPAXfScvX
WWXAuUDac00L8XvYaf7h/J85xmyc+8iBbFoXU48lAuLZsRRQ+6AArq8rYU+zQ8ikcQWmDu8Q+v6R
+7WKJKrbVhtc/dEdn93eVe8RKRlADZ0XpoBGrcX9PKVwjYCl+nfwrqTKmLL4aTx63/+Ax6qefDKQ
AL1v7Pt30tp3pRRX8NvXm6RqjZKRbzU83xP7pIXHslk5Lqthara5q+jwBRLpvC6nqHaXikP5fOK/
q8iy1zazJOBPvru4I4TQiH9Bc+TZgbnzpY2kCKCX85wW3/s7ub1ovNjCsPX9mgfwIXuLUr6N6j/B
kxPdNwOpRrbsyG+gyvMSK7wG/LpKfq4zOPuwO6pokKJ2u4JB5AfIb3R+MubXy2zTmGhrcexcotCO
EpnTCxEDH1MWhlWY18gzzgpXr+BmefmKV/nUY4ADEP8FDScgcpujQmzL79tIzD2Z8CTL8FHsp2C7
0xj+2TQy6MTBdB9TTU47AfPJyFN+ETw7KwMygcJ6B8ft/srzAF0QKeM5Zfig7QfSbP3/Nt5/ivn0
K51LCF90PQsysa8hb8Lr6tb1Q3smOhAchOnVwdjXGrC67WvzkZGdzzqWuFv1fB+7rENkYTtZVwiB
4frFZpdI3N0JfcyVevDigAR0L8bLqMz3WRUlZ5XJ1UIMBssGn0YylOI7IyPB84K/sccfXLC/EjeM
flRD6OJ/3FRFMpBEnQQqVWdaJ/VwzUeWZRUOgciYdBeTDdkME+H/N9LwAUmdmJ2YyYOWKUaX4xOu
rKKJ8UBa2wb9wi9GvKTdt0/LjF+jiOQi338fDFf2oJXWtjcw0YAeZ6AfEL5G5l0xPnXIkFUXh1nW
P87FjEXxeuY48PAzOUJ8PWb6KIuId4Vr/PPG18poQVtq+saPX1NZOZgj1Vjlsv1jyBA2sBQic/sr
pGDXmvTxuWT4Ra8mMk4Bee7KdzA8lah74Qi7nGuZFA8sC/cIMV9WNiK6GuAhbVqmdj27o0ivzjUD
gtl56+d93epVN0hIOI+Hg+eOU0SYlrP2Z9qwVaei3L0JaktHDr1TpFJ0x/pvf2uon30DBGXwMaaO
XM/3Q1vJWNg/noxrvBO9dU5GzCMDSe0RDRVuTfB0sAWWwlH98QT6Gb846PlqDCRK0fVghGtet4+J
gkwwHHImFRr+g78QLMdQWEKL9FQ+Z1zqBr2hVm9h3DY4vXnay9lRlss4hX2B99hdbIdzwA1PP2D5
p3ezD4zZpkk1P4mQbJB+jTx7YS3I/himBj4vnjB/NXgJD5H4aaXrThsrufMcPjKOUum/gqXjiRz2
9Up6s1FDiBJGbn15k78xVLxIdQNM6U9PP9OIMlujV8/gk80D3PKuqUpQM0HjGvt607+DzGuhDT5c
ilTbjiBzcXnD5n1DSHALyr9rdCmUhC2P0CiQ5fQ2futDhJ8fkR99AfNWnKvoS0f1ukQTmHq96IzB
CHgI/p2KQ7IGAmSkDISBMG0c0j3VkS28+ucw0YmwIh7LwZH4sAnFQK/UkVDxBQSns+OuwWxDKMAo
Yly/NFKEad8jAYvOj7AEiCSXCheVHMGSnZru0Inq7ULRiHWFmr8C7rGGXyjP3iIkUvgaB0g9iWoV
m1sRKNfyqaHrHMV9TSHk0sa6YeCEmGNZqbZjwoxuGwmnHg1rtYJXqYsUs1gxuUvfpEAEhF7N0oCm
goL0ERmGRR4IqRJqqRgE+TUlZ6NjSk3wmKH0CfgdpsjHn3/oBtJlRzbUVKRsnKlkHojq8jyhRKaM
0vs/Ko2UOPpjD4CnUFlyBGO/ke5ptbNpbKPgV9y42M+xgukK5sNNpmrdNm7MKTKpXtHyCGlNXTn4
7Pqkv57e4/ugjNt266h+fqmAUHPQcqox0zZO5tBFZadA+MaadszF9f9QhPs9WAusumTWTWMY6E9O
Cc6LVaatnHf1nkER1Xp0q/FYbVMvgmUpMWPbtZiPAYTkDVCwmczq6WkfKsFU89O6lLWSQAwjU6/R
GE62yvIcIUup31es3ylzp+pqnhLXu4N3oqWydQ8T6uuhB0KkG7GgmUGSTmfwqcqSY0JnoeBAbFy6
UUBiJePOGvtTi0mb47zVa97GxXBoUou3/egzmn67O3QlsOJHh02LYm11UsYaeB5K/VVdfXXFpzpv
//jxuu+b/ik60kG36d60MInLtw5AeY+hvLLpP4ABIOjDnw9FWDMaon4nkMdrSvJELIHyKte8xxxK
Qxic155s2Nk9JA1wRE0Labu7mmefoxdOj13OYXi5LbRUIGjzvcVm+RBW8cvaiIOmhUbqX32DFV+E
QNBiPmmmJpDjcR8vjFCy3uspVWJVcKWG6K+0qLY18200QNo45cypaPTwQ1aulpEXAY0SGaTRypEQ
6H3Ayi7Ate7yteXf5sRKRiUaO+/N3a/zG8X5lPuVpi+Duf3FIEbiNDnFI/TOMKLzxXKtovwxTduf
CYDcscsNXhn+7WcFT/XiJBT/TZSqpY9NoXtjT7ej4+vfzewODhnNDF6fTkTyiF1HwVi4KbKPZDgO
jUl49DIdjnNJ4wf9wwaLv4BoAOvtegmkP9FissQhuq7w/9gdbVYuAIHqmxpvM9SZDY7ToUSM9cIn
/7N1YdAyqwQ5Wb9naX3K4oCHtlJJdJDbu3PPGhje6BIddVJBnf0p6EsAl7nEV+j3EDLG9GQGXrm2
y/cr7gP4wc1y5WjtaKbRJm650qwXJaxYEEe5Ypmb9SqOnBAOud6/GAi8J7u5Oq3eU2FEzJbJWfeD
zta3r33tzxFTmGrGa8EwqjQA5r4kfTi1j7kO0j3WxYxO0Xt8hK5sxTaCiFM8kGeO59ozbcLCcbBy
LWAZ+drsaW3GU+qp+VHA2hK4gV1GDN2Y0i9Nnd4QXJMWM0R10A9lGNBe1Te1lfogVmy+JpflzeFj
351LfzDEMBBJndxheDx8Gd3pPQZ8VIB9yADdo2Dl84kVvYrext/jIDCc/8n1WYlb6rM/tgFBc114
YLUdmTmTcwYsRgFW13qJM9csCzIFSedej87F+Nhsgp4lmXVImioDcfi9QlKYQvkETCNNCuclHx5U
Tn2AeAmPj4qIpyGgU+LoMmeN0NP0MU06RmHCbeDjIaLUuCFlTrx4dmmHT4agqVnHIIL4nw9b3WEj
bW1t4q1riteAFmOJNjFJ/gI/dJu6pfufVe3oQFsMpw+f2Z1EoEYh9ZJlfl525SssnAR2oJ5R64dM
mrmBEoiUqVJ0tc9mswIgDbHU81kcy75cag/irhn5GwrmkLfrt0JLqxtQu47fNl0O85Gr8uei5UF8
pUSCPpEU+KEqX7A00pfGikv8sWag6mHf+DfhCN3DHo1lkBZ3f6FMqRiHDLdm41gnfSwW3HQDLi35
QT78IMqpUIhKnHb7Orb52rjPU+4Ov53f5QtAfSuQRQpHnYEnMJCqMfd2bL7O1Gv1V4EbaMeQpnfu
iIIPBumEZgmp4PcI/lo+nhb6+VwNKJAimJiTPOJ3rRU5tTd5dyM7y+oK1ESjqbrD1vyt7QWC1gqR
eb7y6UPIVQpeL26UgVlF2nkoW5sgJVrp/jvfKz2NCQbJVdKhPFxX+S+fj46VqcMlT/7gjD1OGHDh
h55+JDdiGDkPpIjPYD/cQql5DAjheWJdIgDzhol0Y/ok1cNWb0Dc1hPVn5tm4VxJ0Ime+3Ag6A9u
sVGCLm/mRHJsK1OngHa4/mvkYsj2zcIMfD++yy93Hhwr+W7vWAJizd6w1PjDUpOAeYJWmwEgPBO6
/JCcUrpR0AShQJxY7IIMgq9cRXwSpI9e0lNMZ4rTUx6R8sViaHTKZu3aLs51auPfZGM7c1bQUZoH
6/LX0oIyu31cvlFkKRniRdmk/uqyMUszZcte0C0D3hXOAjUDRcRS9BT+aLWMHHkupM7DlDpCLn46
FV/QCmac83HdPzv+hxV7Yke4N1Gxyf6Ru7r7LBoG3XqybQlbP7A2lO4Or0AK/weT6F/cYk8Cbtle
fYfv6qIaRgyvJ/RkWMaO15M8GdpNTh+twq6LJFCuwSFKErqdyO/MFTGiKIaVK4seh6CI1ciaI/Jr
icAkKrQLnSK3IFdvQCyp5GFO5eaElRD7k2dcivL0jl2qg0hv2SAuYuTai/ZYgSQ/PIL/bMF/1mAM
CmXrQDjdCjHTc3DJ6IRQl8X5vd32KktjOnI59inVXO0mN+Lf1+z8jFkeU/aVstZ31DbVYJmbYUEA
/7R51wBFNOrGdavCM4RzgeZ9jo5XjTEXrAuPQEGuNNYLgqNaEbH71NC+ERP3Z++/uaTLNP8H6xN6
a6jZExlaz4Kku1VY0C5euMHuarHB9HzcnEEQuDCXZwtiCI1v8zqlfGXKy4Hb39j6/BDUA/mXeBsi
CO9LJ8EwojoOU3vCVN2zIoj1WJDBmSXtY0Y7cR4P2VuouIxluI+sMVEtfjbJwBceIg4oG86kcUFr
XWWnWIyYD4sIm4R8Dcn2uo+D33V5TQvbvEjhgSMmm05TzIu2YF1T7NWHFY9MBtAgC36gBMILua/D
UXDHBMDJsdqkNHVPC+HnkFACkFe6bNahpkWsdhPLEskUmiXMTYD15kgetYrZomEM0gwqEWXrl1Uu
SEb0uTBYG1spBgzLokpH7su8XkM9nqzzZGLxVa/KBvyhpMa+pzLixmeGWM7htDYMRnm9sSU5c87s
ATkfzQSUGRDwGKbrWtNhTG5zcgRPInI8+hEze6MqiDdzYbGzm5Hmf7RRnh5m/xTaxZfRLRG1IbJb
0VF/Cfpc6tVIMbdPeYCF/oMGp+nJp/bKZP/4Mw4W4UWzXYY+M2nDV+r0hrIH+3rirgJ087Ye3U3C
PSaFSmrL31+5pIvyrIK0rCYM+2J5ZRE+7YQCplYwL6tNR4pkeY2WerW847nyK7M6svbqfsIV0orY
5MDqQKIvBtr4cuLxwrD3ad9oXjkHROrS8Ao3PKtfVVylOQby4zSenMaKBJw0Bk9D9XYAXHllI+gv
05GdT3oKT0myy9GJm+4jcaipBaDYSvTl2td9MSmv2swkoOf+rl1v+OMMyP2ABe50GATfEAYUzlhZ
kww6lRUBAA54mu0WQ1WgfCE1bryqgOT13OMJ9qF36xfkyEs9Wfynl1frtkZUGP1uVbVZpogw4/ht
aDFPKoHswfsopxGu3YzlS5scjsZd5xSb8EOsUNMZM1dm+eL/lE6EUmuiaqvAMochFUAEYIVvdbhp
gBxt+b1O2k4tZiqm6XIijSl8EF1ZxsUVrln6P/640Lhut4oec4JO5wPOM858dReCY2YKHNUMoAZM
lh+nP3LZHfteMrJb9PlyYH4rwuMlv8nwvY8XwTys7H0w66aaSfheBWreSBzh8ZzADc12/d3+L1At
gnI+GJn7ASJJcOT+QdT94a+IEefZpon2PdTi+VQVa7J5HYoDkB/Jc05l+ZE2ESdhVRZF6U8EN49n
SqUbM2TA7sV3i81TmdqdIY2Uk5oGd1ZRLDMiEDMVAZI7F7gv+xkvQRpGsdWUCoLSpkpb/OasvHT+
Tv0lY0axNIxdSEuR6/2yO4eaGloUXB69b5B4WmhOWnop1WvOfzilad+dqhrdMGVrC+VMF5HRcxvA
pHpFABed0QWdwLV8jbDYGvmSR4KxOlNE9Upf+IdkrheVnZnn6VgbDrtFMWtTclRp3Vh4o0fFRumO
7GWlqY+Sh4OfM+dGuRBQZDHbw64Br3ZI3NOHrrVaCMiUIx1UoRxZaujuaZh3TvqAYtB/FXXs2LIx
a0P7jfh+to1yGXYcKS8HCOZYqSmxxFM7JBwWtkcsyhoqQ5OHHqNVZ7vbionnJDiMyqrWIQSz4KOy
LWjudEgDwUD1CKXFIKbfbflXy6ISmLoF7UeHDUy0BpbyV61kvf+Bb4FX5sVhDv3w//EFTcpdlKCh
ykDJ6nXG3Ib1wvGYUlFXyg9lX8cErDkTR30j4JdvxO8Ez452P85nqC+0AI1zGg97t/tqfqDtFv/6
5Fz3vzZBpDy8gB2/7zzFwVfPqvgVttdw9Gd+lwEdjSwgO2kFuyzyb6RXjfVjznTvbpVEP8JzluGT
rkySrKWwtBs7c2XtEEvEzjh9SU+dTb5Nu66askrlu2/CY9Nu8FRT0rqVnD0zLwgWfQAR4b4rN1yx
eGFNR6lDUHGWiFOih4vph5oapy+6+OfqFdqbGIwoGFzHTunKfjTU3hPlmXbXwrwiXtsNqLZWSeR1
xoUeqb4dPzbBPSpcfBJWQ4D0ajA9gQE2HbjIThCwCg8QA1jxkPCtT3ghO00euHJfbYImxNF1JKSD
Yedma9er/+F+S8yhXWIWDnYoDmBwmqjvxroP2cD6cOO8CUkcGXUCDWs3o4yXOt4BLLXGmWatDccM
LVgc12f0ia0xKLF1xCNNrcopQBxZOyvDEz48MCo/H/nyFNmGlZOxqjhGSLqYvdZl470ffeUVYE1z
RRxyz3cixVLu0FjIlZ2gpc5GLF5BIYv5XdcqdDKEppyIyh72w4OhsVuSgsaPuWa5HGuQdJbQDnj0
Q0vARULGywrfmd1fZk+2+CNK1HYlMWUmntqZf2sq4UrJtUOOzGJfm0ttLNdatex2k+SXhY+Vq+Ds
v2kG69XLMxjL2oDdb63h5zZKaB3bVaO4sUOGDCpzyQ7Pn/Q0zIoGMJV59UoOEFN5x0DZx/6/c8up
8K6Fi5p2X9uUagoQe9ikTiw+iCMmANoX/bIgqhlPoUCcgUJTjM7ew2tPsuqUsFZgk/QwjHOO/tXY
0WcEymJB8b5Omp3jvYJ+bKPqREURFReNFrjQW82nzKDFFfC2+dbuGvjuOn8w7C9m3l2ulxobdBQ8
19pUV709S0SLCBmTaxfKHYiu5Ip5SwYkktSfZAJIR0su8P9mHhgz7bWX6yBfQcSAUmKR/F0nyHqh
bt+vIwAKn1m/aVMzMkkJOj0cTv7+thneZSPbItT9o6eHSYjTInn4pdaBIU3GsmQJGpacuLMIBP7v
ooLATrqlTluA6Kb3uenHthNo3udW6nVEwrxI3nTz5GvriMWMpO3KByNfWwsZOCrgdwbLq5QQJnK5
9XqQVYzhjKlH+BnIL66AqtDVQvyWnC7qDK4LkE7kl2XH6weclNBuZkEgkws9CqpdzwaLCQa8VrpS
J7KqQto7ZPzqZNl+Jdt7hk0PBboanocK02OTjaTVp8N2J19X2Tvx2OMfGOG4YXR6ptSiYQwTymyE
7BDbWLgCV3j9p+nmQ1GpG90eTVsolSlBeF9AF5eq1w+PNtoUlHtMzFWIFE2NGsbMbdCbRLsBIPuh
o2+wdfSOypu2ctaehkenqLJbGK8jt38JNPr83G446h5sDkZ5CF50DuwJ9g299QE98Nd2VxnULy/E
YIuEyrwi3QqXCBq5kbLH14GCESWXo0l7fz2FcnZGBQaZxZGi0uRotHdKo/xBbd98UZ4lBhH0GWuD
O3NxhwoAjjUJaSegPallFnlD9a9df80ODLvJp0F2dkFISOK+PfdzAayoPigWZCN8vMtmXxerG2Qa
5RN06sanX6fZjAdjf+Q5khgskmpvLDpFcu5cBmTx3jrKokYUumoT0rrUK6nlGwKqWJT+KMCi4dCD
1GQpqNc3OlUTJabqeRcArz+b4Sgzqzz9ozGUeOBQeqyyEWdStBJnw39DXT4K+egwaSfFnkqVwrzF
KBEzASW4BUI5ZPRXAO6KE7/8YrTNpodefIXPWcPrcPPI0dOStgKIu/0wHYWGOQHTkeMVF8dS3/SU
6D9r1iYk37vNl9OOaoYt4tl599SA+hVltnZPujqvqkj/qpO6O8xmw5vVsDTEoK0AW1sqo5ExmEt7
ETRb+3ltNocCvvZD42Wq7r+fUTII42RLK+7NNtYnZ/dZMW1dVI1YUQPzuwCFHLzQ93auUGUBkDUk
NzWNmyLODSU3qpbOe9Y/zA4z1O1Zr0lrETQAITrJReUt6kb2Isp60z42hQpzRcv7BkYeV95zEwaC
VYAhJpQUFbdtKLywJAkoajR+KEXDUqdMgU2IbGiMlkJhoUWSw7mYT9nxcXYh+qXME2i4aURZkypt
gZGAwp+F7CoZDP8P2j1bgR3GIJvm30eEbnhWxgUU2noOljOLmpp2Xkwzi8JksgvJwrORJFnm05n1
FEo/PfezHD4nZ156qWLYxjUP/083ZXntgqlPwn2TVs0f74hftoO53lkciWXcKuiAF6YXm1mxKNn+
bbEdG/Mw+2Gsbo2S5UfHgbsYFYivaVl062bNLMIAtUXkDNCdC/cm7DFV4WD3q2z1U93Ehro3a4EG
6G+0XlfWLqOf026aNhdsLC2ZoJp2PlZAejeIZZ/blOiylMlsUOsrw9CFyNPJxiOCPKpxFm7fiudr
0t3KEQPO7+ATI2C6RgQ8pHSWOF2HmcgckD5YfswxSHYIXN2COm2N+jETOPYf/bCpCrZA2oG0Muco
COV22UbgL5y1p4ehL6Eo5Ci5RIIDDdy9mzawUARiMou6VGDtxQcwfSJTu4oLi+OCQ9/0Z9Hp3u4R
CLKy/AlRNOdFnIqSw3SC5jsHymjNL8TYVGOIuaOxBm6Rai88/C2wR5uHIh0H/yL7H71lM+ZjMYgS
jkO4SBUavXRTjxORIN4C2ZDz5wEY7NqAB36zi7GuOmHFFnRj2T7fM2Ii/f8uWGfudfKMGFWeT9Dq
50sRp6dNq307ChZqQxSwOcqCc8cxoxakRL+Y8aFH347ffS6K5I+Ldkb0zRFO9gq3TOG9ykjQi02a
UXcqIk9ffuWRKIYAkQP51jKgUMxAjaeK3sf8HcCeLAsAiwm6eL9LCm4KvsfeQ9/qVIc8dJKWCxEJ
o4jy3YMpIL/iZkQyHcnrIKyPJQjHra/0CGA0lOEQBogXVjRo4X9qcvyOUf2JnDDCFVjyIE2N/8SY
UUf7Ar+yYWlE9wzsOd0O11odaW1Gq1N+I9b1m+gVXkY8vTvAZNhg60hkHphoKpqrO5TUUacB8CSG
oRm4OHmoZM5Fbb6xeLsgdvhtE6UtpQEI4SI+XfaNX4qGkWJ+hYoniM/71Q3cNFjL5Xngud90FW15
o8lmQ5+oK9M0hMH4r5p+CuzQ4aPABmibTcu6cYRQFqDZ3B6FRS1RJaDV99V+LIRCZo/oLhsWWO+T
nWBl0k3clZBXQEEnz6IhpeIp2BVrN4toMmaHtVTHdtOOZ/lksi1DVnTZpK4QRg+t7Kh6oUaCnIrH
AW77B604EAPWbM4qbZxPG5HK2kKIAhL+kCVJcvVGSvPmqq5FF6H9hwIbiN8swA1TqxqkUIxSGBan
xUzr8H9FG1mpzvA7FMZMcqy9Gn1gerBJ02QDFBAS8Cf055YpPsWKWGzpX0bxE940W4hedBSgr1Mn
Sb1RjD+No+r0eAnnQWil9nEEbe31kB7OuiGUG8D/xFFepp8N3AkJ0iqcevRnQ7keO44ElUq3xll5
ZZ3+mUXX2fq6ioc2Rypp0NhQsCk4HdhOXYtlrpB1EGKqDtAmt/ODP2y30ejGQt2rV7N/QwB+e/+e
VwWgsjEk586Z4Wxj7eJtOuiPB6hmEMA0iaI0DtN1A0lbPGXSwPECIP5VZE5th49dH6CpigsJpGUn
/INuDzNGjbGOKu7NzSPVIp5WMQZuceosTlYQ/dvW4VFpw/Izur+cKzzMk4Q3OiJBDb7UBnzwAasP
9tW5jB5UC3vQB8j/LBesfJzMQgNf7ilQ++8wJnxcOjRZ0i9+LrIBoqglUGYluTZQHkx+XnqIeGtD
8eXgNdTeIPxdG6VRKLiqLHmomBRqk1SINggLZoy7SuWMR33UABFhkhM6aRuC27mJJ+qLHC1LQsMR
b0FrtFH53k3ixnPkmnVgU49KGN3/kyibG0AmOi8YYm3q+DoSiNdj/xpNMVdNcjkF681VYbjI8wZw
rOuwDKbYFWqSkr5sUPftDUPMt1UeiDCPzySQcK62RfZ1GDn85S0elN8HUj9Opoc9YQ7sd7+gtygh
Q1fm8cA6ddvas+ZZMBDy+Nk2CQSmE860UHRxwi36XnB00JqZ+cRDyS2WQZ1/+J+TSHnGUQzNVOPm
LF6H+Q7Q+MrGiKT7qL6kKm1UmOqPHcnlfwyWtUorDmxpX87EdMb5H4J7Nz5TW+t2I116Js8A0BUt
Kdg5wQ4/jFx7dYgUfnqkF8enOuTD7UjKCvl0DGAHabAxZfIElfQ1hJBgTdoSBw+RwUbd/noV35r8
cNponlFrG6JPBW7PIXP+X+vRXstK1NV2c2Qo3vCAXuhrYkr0RgGAkfHZlN94x1QyvYRxSqeeA6l8
+0yj9ffNzX7/GD05wkSsai8lJ5LyEeCfliEuhgU5C8ebV+h44/5H2exZFnz+9nDnYSxIyxRDlXpO
1Kg/HiEQSPXfirjpQnUKXPBSsvFEitruZIpaGdmrowvSEZl8/1PBsBNrV95/IPFuFILD/bw8unNC
S6L559vL+W1QftuOL/BDvChha3E22Z25tftt8YADIZktrpDNgP+2GfsZnS+Af/R7RekI8v+w0Uny
Ica7AypTuVSqT0EnBSNGwf3m/pTX7LxnmFLVLqhLNUx7/VkRpTfJcvw0dywic+qk5oVLe/4VUSgj
dUZ77cnEm3jmkhFwznkJQZ9Ag0gD5UR0k3qPq1xZdmOJA9kFA6u45ITV+Vv4Oiruq05LkD6CEFMM
MeWGuv93ck0RBt4Egp9Xz54orgQp+lDEQYqBFz8IzRiAup7IdPj15N1Ie4mPVDmoUetxkFmjUm30
Crkl3JHBgYcKCb+4zqLEmBow6/NMnmEwB1N/z7wo++XcI2c/iS6VcRq5HIdnV/Bch3m0tKmYdvkw
NmSVgqzKEZXRzK0cSSRXldNKuyT4gXs8aEbhZTZxfJrx5k7fw/sGYwXBlvHc7vZhLARK+bQT2YTW
K6pLZ6yH+qlGLMBtrbwV/sms+qvc5Ck/NeLUvRh0Y2QjFbPxB3HGI3r/vAnCPLjHhJ064+oacrUn
nywyDN6mxcfxOj5vwLTj4alU9g8KovYBokm3TR8MTdPrFHpZFUP/mU0smur3y+Wir/iDXj0N6qgO
rw7PeaMbh8wWum662dGLJnoKH2Ur/EAXXyay9con3C929+tMrTEgPEdWFSyH+VaEsiTxWJBcoqqn
wYSI7OBQ3PTw5U7Pg7oBzeueTQX5OnonnqSxmHhs8jA+1uimSxQDUzewOzGEBBJM9FktpVk+Y+gu
9T/WRGsl9RhdWZZcFdCck36EJNYqRjYBfFslWk9nJapKs0UJ0vw7qhmcXU0zNg0hE5K9tIMwbhfR
HERmZL+/h4KMKE/Gj096fWpoV4Z7Ong68xdB8pvmweyZ/IaX+WsGa2ULiwhRPYm7ZHQd/rpcy3+a
LKYtwaaC/VZATEFbxdOmUn3ibbNVEDYpmDuluBsPPZlctIUzi/LWctoG8yFBSnb6HdSidp0OZTg1
G6KX/1Mwh5hRvH2b4CXTScr//cQoBUp0yHNhw6JG3ZXROVIaj0/Q+B5W2THUcRzBArb6nQNGrqag
CCGrONe+437UOVMGPv4g2YhBDkiC/oIfSwMjw3MrM/EBZ3jgRbPu1Li1Td+FCE3/b/joIUv6eshn
RcSewBsPrLu4viFPJjFQtT5PRUyDkhBADr16s9GzhPmBIG197CVbvqVG5YrGyAnQ9sL2+DWFN6QH
aITwpTueq6fZbWBXlhw1wrtOMdceFV3vLr1ZNPQS2V7e3tSS4wr+UMEQXnQMIeXqikHdP9m+jLXH
D7lnQz1df7OcABnSaaadaDie1QNp+UBeLsxsM8caGtx90CPbS8SXiOGfY47EAuVC+SziIaeC55NY
JGAwVKw1PcH7MnWqM9KpAcw/hC0nwFXGIBgZcMbZrFwAnmDX4B1F6cAgKukKrHYASzV3oRq8RdT4
B123F4tjpo02NLHN9+3+ex6ZD8HuctxmoO1/sb/xI7sEyl87DK+49Ol+fT/X6w8J2RiGGrecTyh8
CZjAKtBArMdj1KT95Tk+Yuf8DtW6Dypkxg7O1bIhtHViyA9ySzozLklC1vqn5oO6yXfSw+WdOHan
xZ/AIb0hiQQKLZLFOG68HLGRLnB1+kY64BrKcqCAAmmYT8+O7soQ6/mK17RJ4AW2cwOx13eRPFci
R90cHbj00SeiDXBVYDTKcbisL94lqlG42rvwOM2YN4qvGQM/bR3VXewyDJYgfe9ajfDgjXMRfv0v
KnsnP32OZJ/O9U+RNZ7kWPCOHw5RineG1fhnDpt1jX4f3n9ruL+0s0Q7hDSD47Fijjxq4JPnmoiH
OyMEIkUOjM3DMMR+LtlJ8Y+gERZ43CDmN9kwYIJncqvC4pe7jQUD7OJe82GfT/2nHhe7icDc7drx
h857m1ATffS8tec3t2Z7T6tJFvVumexCeq/BB1amqhQ6o9ph/C6fZ3L70k5d+aMW504s+AqYxHyj
Hr8eKsN3lLEBK45Ka9OLS54ocQ/hof7m3jhEwtNkIoL1kuNuMddsikcncCPVKLIJ5IimHeMRSqMD
++Vdsw5MMWc9SPnEXiaiXR2Nf/o3pe8sTD+N7xgftFhj1DnX0epj0MSrJ0DX68JQZOvZirg/64xi
Uw3rnxYqSf3ux90IUU9kVaigmQxyluTA0BetViahU44rjsEd0TyvzEaXbeQWPVkVawBryGDMX4Ur
d9CmaBcfqbo1ZWfkjunpTZaco2B2fDZ6hMHOCp1l7RTCOCwlFq6o5VCBDhU2qhU93UEPleOPmb1c
eqNthv3N4oFeRo19t16yNOj5sjwl5xR4+VKOD1ykeV25NCu9KikWgWHs22YimmS3/4bQG9PS68zw
cn+QYgX7v6xD2StKnDgTfZdqo4SSeUnq2rWAhf7XMIEbj+nOJ/s44mO9twZy3X9wTL3S2TL0y18L
MnS0yTRpiBBZnwZJCD9KJd4O7D1i/FLyBdP5WbSa/BmG+3i3JJFvOk2hS7lpjyEgX/yBW5eoe0Nq
0D/gq2Ep1JhIZtknl0WKMbzNszK19BdB/O7nYM8OV6yHCaNMZVahPdlT0hFgMxUKrjye/EYc92q0
mA98P9391MDXIpo6rZfT38BW8wVuHNWmLhCcbT266506rEiLRQfl/rqQZZIWsE0uDy+1kqLG8dMl
FGex2T2tqa5rZirl3q5APnPFjneEFExmXOeI5RNmh3j805My1DRVV0+fVOsOZEjDV4eUh+l/peTD
U+F7Jyzv8QKVZW+ZXpnv+0k8xrAM92E0NbaYyW5jyqyvmlh5Lm5tK2k4Vu3NdcrAqWIXgZQbR16c
tHGKOYz3SpLdPnsmBZdlx9nQe3JmL0hKDS9YYrWZfgNxqhXkp08pjzRXQvnFojZyyEv60rQBQWqA
oNlhEPVJ37hXhkaLEwiqXfaaL/wzvb3EabLul0TQt46Id50Ybe98wVjCvqic29XJKjnG79wDEwce
l8IY+mlkawUoCBYj/5+lEAMR47/Giba4zPJRYNkMB2X6O8PEIt9t5N0vnTMydKRDmHcjPdXP2hEX
pPVgK+8LeOPiegPL+2GqYeD6A9XX3KxHPNfJxAxWkM8gbmrGbXVQVQb5Fqk/Hmu9Nh3XQGrCljC8
ix1gheHYBMfkgxZ5+wNry6kC7ankYt6OUy8ZMlFWcbBaGOWq7ks2n8OFQ8zQ/Ut++vZ5WBJGbph9
3nKypr2VUUIPqAFE1EQyoc+ldZrmY/vetoUU2QXIXBZicqac/GPvu+NcXSfdTV/3rhvzP802VxD1
a9VbxfUbKiAInhCaqmYLiSNBcIw4hzfnv3I59UcDsK7QtMrXZF8QHTuAIGcAq9caneyi8UyEmwr8
FsIlqpZ1J0TdZRIGOXx6b6KMBuazu0NPwNsHLzVbnCbzbgOfr4CM6mSL4334rI+j09DFbjOtf7B0
pPU2Kzyvk3WfueKWL7lSmk1DJcTdAatVGpCpLxKrDB6y/oUUz2vMX6mPhpKAv0K2+HPGKw6wxly7
AYv4cwGx6kzY/x7KI1cb6WL2xd/K2vK0Zib4CjVv30YywW5Ow5k8drl8ujSPdS5vbW3Apfjl4tnk
DcI9yZaCV3mvUF/PR+L3anOGw8cSwnsi2halz2GXnOBDx3R56Oxqduw33C/tR31cwJ36I9+74TGa
43jc1wr4PvIX6DsukcxEOWyBQLUynxlXqiDfCfEGBzhIeR2Z98K6Shw/hCjeOG9leOfoZtFpyfEU
/PJCTHORLoqmdAzjT+5VH7T9De7Y3e610My2XjlXUr4Y0h0wVxc/t5VFOL6XrJnPCVgo8OFV8zgO
BTsTyCdnhHrA4+KZLVlMjV3hemZq3nO5XrbVguNEf1//mdS+PLEtvIXjgpY/NVi7c025dXa+t7lo
0b9QtrbQV+mAb3Bpq9cwejdqn0tbnIQ4sD57u7N8KjuFqJT53p60kA7EkPOQR/Pf/pt7G2R1nYR0
5oxVmC5yZQmEZ59zprn8aZW3+iCWl8bMGnH+ql/tM/6P0mvYUjrMTlJBb2z+rASuRL3aMRoaQqFk
P96P3ykC3lOY2BdeZ3pIQkEhm0gCiyCraX7Js9MtOaNUaJHCMIN9d4LhEk3tiz5VNXk5UDHsUPYz
PjaPdH0214OIfofu6cLGaN2LXxkTVf87ebemZodZYppu86GpNRlzco8wt2VZM3DTwoqXl3NmRx4M
g0EmPvsZ/h85NlTXPy/5A8V+Qg0hir8Q2n2zPUeZIoYpamWs14bdkFW6OjMC1gxQaEyU6uk3Y1Fk
M6+DfAUOMeXxKQcm+37CXmhPhcwtANiwmlIxHd1zdciPX0NaHsyMt8xP3/ecVPEDpgRSn2PXGYhe
JDlGGNHQvDORCw95/B1aeiJJKMcoLU2RCaNbu4HcuJKrdrRWAz1ZV2OAPJFFpqUFvuSwvQxyANVv
U9qDHXaZVqAJofabSW9LWROxWBeU4SuJbq0ExkqtSzjEWlfNF779lnp6Xc/r9ClTKhPi+j662Fv1
4+kCHN2VczP7D8BABcD7Cm8V8Zd/v6UeCzoywlMqgKrY57yEMg7Wz6PylfjqKJluLV4zYWtRXKGC
viL12EGw2jy2Uz5vWwD29h3vJ0DxSQWXTs2G5w+Zplvnho5Ed+7BEJJ9eXE8CuSMIJ4BxzDE7uPw
CY3/saMa6g1MCwP3K/au2MXKmQ9FpBrFew7eq/uTievB7dys9T/zMNSLeJDA0xOzj4jrAxYymAK0
Wa4/nbcAfZArAdMpgv/zh0OroCLTF4ez9oNKqQF1ihx4BCyoZa30nVfOJ5OnvBqDIxn7jLvfqOam
BGIfwxWpsU88R5kP5jga7Ps4b8xSSpf9TYpkeRoiLYFoecf65/sKFLxukbpgwBkrbADSNsjzUauh
84krlLPoTOjntnTObSpviCsgM93aFiYhbhlFTlViiZSM5l3lzbiYKJFI+d150Y9lSlE843zfiFEX
4C8SPy50ol/sDZBGyVZXzIJ+jAJ38kYX48CIn/sX23KZLJJhBG+M7I9c2XigrLIOKw4Pr2tjtAi3
UbeW9aBYmtCCUIZTrFjvy5YC6BLlfLuJKvE9uNvgJiWU5ujnzgttOwoy5+qiuqaSxiXNpOI4YBpA
pv3rmQB+R2ojcc6gacR/SMiwqYd6mc2nc4uEAiis4wemm4MGSywce3hncvRbeVh/LsL9guHmPD3A
Qp7t8TIGQ6q5p8SvH/3UObAdwIEdS5AdFLcCywgtnNDIje2MxUOPXHflCEKEjBh6Bt39kcozC7hK
xFb7R6WOLHe0hoMYUDxLJfwzwsK3TakoHzUGWOeIRpF0B1tIlfnEZaHNACUBbQC9mnvN8xMjC0zf
sObYBwcl2evqHNX9P6G14nnimG8hV1wkSRbbRfvEzD46l2N6rp9Cse1rgxjAY6yw6g/KskdarWl3
kU5ss/6q7i1uL5X2DFMX3W6mennKItBMCYzYTF+hdE0R2y9KrAMDqUp+F1dL8lsCc6hK55qLPjMq
DMrtITpjUrQe8gkD8m+vi9+3du2isaAU1ws+eukjp68FmvlnUMLCCqXiYJ7Qnku3qwcEOgjDnTV2
+3VUMF/9A9K8Gj8EbP/4m+qXUUE42SMSFE+ug38VScQuI0bqxSzj3+O4YbrWnBWoyp10Ah/BvQCO
UBpGZEmvnjqsJWqoG7GO4Rm3AoqYR7CoRdiaR3BBPH8SEtXd8T9MCnn6xoPNwFiOIUXJHDBYC0kH
p6JPTfkvGviHb9buWlzgq8TwxFqooufju/Bw5P86QknPJDBlPSzMBKdrya1DIB2RpUD1KMjMk7ry
XWBnj7iNkmd+uwpSlBCKrFc6fD39cW3kEehykYmY9Q5Zq4SkXB4ctQpuacgYczEXVw6vT/s7iy9B
WCdpJrUBu6A9rhshnjZPMiBZGbGxvVdpPIIAxud3USerXwoagMdkCg5msRd67wzA4VVWa8POJoUH
NOOlwggznGqJLv6ESSoQr3Gl8X+Sgpc8HMLhyP4yw8dePAOhOUJ/L68UaxZqZk5Vs4/OC8SYmvCz
0H5165gBtHkhkRaIrsfSmhO+TQNKL62YZZYldMsCXuHK1Xar/ntxXU57EHdt9NPqi85BAq3hoOD9
KFqu4jwH7YmHZzJtVOwPV1MqYslbYKgozziAPBcD8F6+RvLtpEgzbzq4ib186zarhHE9L6VvnHb6
AMf7HP1CD3PWH3ejuuu0xeLWvS82KgICwld8AML52zixz6eb6XaYcHLbXNvCXdWy+gUn7lvfSY7a
9ow4Cd6Y0CdzRS8xCSgpOBQ2hhwhXzKCYzvybqYA5XFUQWefBLCWY+TEhHHyFN6AEiyYrv5szdLq
EQe0lPgv50CZk2VddR0B0TBnGquDD2cLVb2FIGf77pT2BdKJKs/RQ0aQTWNgYs7MZRuTqv/+k0E/
UZItdIPcM74dUvMKNx6r39EzT8sna9WgDfkwoy2bTd2APfUEs10Y+OY3RpAc95NM03RTc+4+JivE
DZmTqxeNqDy8Ln2rywGSxrVrvO/bKF6e0A5IGjx7irrN/Xz8bxPassOUO3vJFGRamANs4nDxGmfb
ZipSN78/uw/XG94+SkyhmPEiDx21xkzeWXt/aEPRFGtZ8EBL9dnGE9+FzMe+WrmAUg5E7ucAaP9O
+IBoaFivfEohN9jy0ZPo283AU0MCB2ZyblXPkHzx6ynOg3oEVkPQNnQcoNaUlkbDt103G7ydmNSp
Xy7UzWkRqd6TPCheD2HsNTEXc5W+QFmCQE4PQIWc9b2Qvt+yJzofSgBrT+8TcDXhNoH1Bz040UBs
W5jj9rD6ZySuzhTXMSnZx/Lcs9ILVJSrgCKaX9Kk1qbTE3NRuiiIgJlJClv+fQgDTBdamiE74Gn+
teMOrLUGb6lVpwwPU6Fu4YKMf6oG9peQiZIjokVmOJIOTESYbnZUkVUqQTaKhCTlqj1w9aBknNrW
MxeLl5BriAWQ+r9ZQSPWu2yQU83SBY7Vvb6rQEKgcj1kWeq9rp94KCQA4gjh79+eeYfHUplMyRxV
z+LGqF05Mz5CsORVd0uiyyktunI2izx2XZl24hdBXS8ISvxJvIiltA3U+tnDZbiKHQnzt656S6PK
8wqe4Raj0RSDw/y+HTz2n4OZy+Jxfj14dl5BpCnJWHqWcYwGpo/FBp9NbL8kkuXc9V5Rd+VwUFuR
Ot1UfQL6Ej76X5EnFYnxjWyjOoq7h7Q31KkqoHENsPd0GiIPcaXN5i8Kip519IweIznLNjvlVFNV
ydESPMmwSbGD+lsCZvUFoO9gkhvVH0+5PSOYqutp5vaIlP3+d6+Sl0SinykLsoIgQCdGN+Ma6xRE
sR1P3Pbl9VovFqIeZChbxhV7kx5e4Pz4ZvZP/fsk4KM1+2HUrcf6Co8xh6dPLj6/yiU8GeTYoqVm
E7Z7z35SXR2je0GnyzWypRSRtQWlHOFn2Zmo0aSURe+4I67SlW2aNUWxo4GTUkCGap3klM2QN5Vg
HjLkL4dyy5UswsnIOrp7ozOrTT3wGpvnjxV75+XbHq8tD0ymoIaldAOS4HKj1nFBwANMt5w2NAXk
Qfg4KDdmigD6qSEgADLykSmlugbtukEerLVl7hHBTK3jkIIpFQhC/4vmX1GcIQVDlo8toPnMqJ8y
r+LpMMtFa9s6LZvT1gZUBeQ3De3OibvsUb5cg63PEuvEFwYVp8727nn4E8x36aMLB2+V/A0p2qXO
ZdFSy6LafRYBlVDRG/XZHpyt2awEgw80Qw50jke7Br0iPdtPfdT3aEZW9lEdx4Nfa/Gb3q+RPJWZ
mFfU2UGSLmI3TYcdFLUgkQPvovhNqc/XLxNqTByz6RNCMBUSc6+97MUyOMNRUwx/iany3gcGNJb+
8V4EnMGzbx8diAp7vV+VQVJzaPJur3hFL2bnCW2ed7dD87bG+vkKydF9ag/O0fyUNm35DhNULQVd
R7cyIZDWXd9xLRAyZIaOb4MwcBWBFToeVnxtVAv3Cz+Yfs68qtgas7BQzY84Rb5GpH+XXJ9R4piu
eAY/qvP87uMw84KGqWUeY94OSaiF22wpsgpjT/hoRtTrlyeQ5Z/uSnyjXSa66ER8m3ABBHhYW9D/
SkGbHZHu+IkdMRTZsFg6PbDlH0CNZZHUKxzJh1SShIWR8BVbvIJrmFdRLZQl6n6bGYMKTQ7cU3g1
Y2/dMA3XMVLy58Hj1C2K0GcV7MYZj8+7sXg32bxcL570RDC06ABvPAoZlf/kBvbXqSQnk0NuVpZK
4oBzCqzLvLcqxR6UDgB5WNgwoOQemVngIHYmcZt7N5G8I2kXBLjn0msiImFwDGnVXt+PLNDfl+Zr
4kSHO+1vpgt2Ul/lxTHYmaLAuKlaiv3vKAqJGn4hgHOsQdtX5c8G6LZ5/NkoxOUEBtoypV2EMgLL
MFhPYIOJePJgwHY/U3v5GLJdrACY2QVr+OmX99n3UL1N0JqyY9RKT0HIGczkCFyGUhKBk3X3+O14
93qIDqixBjb+yATUNfUWkf1jaNARQLIEpvRXyukphqggQG4YhPGakOVBvP4DEc1XvVBLZ7nqsnp8
gpu5XSKlJf3uSvyy305qysiZW8Cap0US9LJerbbyIxTcuzO0SumLXi6MXIFwlZHTmmL8jq9U74XY
4fR5YToxSX7vsE03H3yx9t9n1hbb2uF2lmkGqTSvKUsNzKKuu6WHODkY32WlQYtUbkIsyMpdxypF
qY4vmuHhCetwRFy0Twp21bJfgvgy0v3sBY2ECthMMybyETLjXsaidKSsrstTM9gFUtKN6xWxhVCl
SqLSl5HRnW5eo6/y+0asVtw1G0XcVwDxygdaMBvOpDr0tYctnVCsTKOrVZ16h0y9FCMh1r+psZvt
JQLHzlGNhrJnv5MCMZX38Eo0llw7truFuuW3eHIpjq0cQ3gL6KaJjgJULJxA/jmJDtvhilZ4V0CA
lpHVr8eUmO1+daL9gYKJ+8rspAYnGjMf1fTFFvQkO2Ym0smX4/Rr1r+IUaVjcQ3v3ekB48rhPSj1
XRul0rEva17HBhuzDc4K6hN2v4eZwbrR5t1i/pjtjkN/cxdwJfjncue2zfAB359wmdeuHs1NtG/9
cO04XqKPbhtNSrB+cLyaTCBfSa3DtrLT7r4iYUrfDL4I8QaCEWecqM5SWUQjeCt7JGhgJXan3N27
vIcYvTOqWAD2OXbRKisFHrlACIQaoWUnHmPRnFDuivEzxNFjvrY9w2RJKzy5utVkF6Th+7unUd9U
B/FjvTSz4nu/g5vDaXfGjB/vHWI+c1dRZXpsh4KVv774r/f9f7eHh5Xwd0fVCXld+VV0Z29pJOR9
Qe0jSHMEShAG5bqox8giOXOb0OV6hWf7y7meYmpOgCWjhK7fs4lu3TaK7rk8flwdBGmcOJSfmJKL
CPBWxwNruETIH4WDinC/INmXaKeSrCd1zQ/r/Awm8G1nkxCpAj9LXAHVdqHeTK0E66AWupCr4HhN
U6RZHpX6CXuOS0VdeB+jTjvfr0yez0p6fVr1mvMrTIMk/k/cmafUw6ywISFwD/a01px5cqF7Uswg
SoNpnuhm6vh5fQG4cHi8oMEGpSM81VMmg6Rt18kQMMVceIXQ8a1A/KiOdNrdrsSjAZpSVCmuSgAX
OLU9X6h8V57djQSoA7x9ksmkLm8acOlEYJr+RkveIn2udZlIvIxquD9On2l1Z9J5LIU8vLnkZbVw
w3SulIFA1lo+KjpQko4TVXgYCEXA+4PFQUAdUO8PneoOzLoBSYmqBmNyvqvYTdF6GrhD5GHdCrxr
WgJalg6NayGJK9NwXjfjGKCYLtLzstHwaKhKH+V3Zxht96mNjrp7aTEdz1i3iOxuEdWAV2qcOg7f
Py3OxmXwuKVhqeAUOw+XcYeIbzRm7ZmvlFNp370tumyK2zwKi1U21Pm7ZQCbPKBHDTzY7s9UhBhY
lfNvCR/y9ACEbw/0ZHpmMO9Sa00uT433ZeBCnj+TkYuc1sRTI3JehnudD9/IBGZMGJ30oV2E8JcV
NKbWZvf2bw0K3o8c8FcJCIQs6wD+WrEyUO7Awgp34hc/ssYMVVaxHyXY7rRC6mjDt1vE4SW59tt/
NOfsJAN4PXBy4rKl+pzlxww7KvZh1qgSGd1Pb24QLbQHXNakYp1kl77jd4Zvi/BqraM/i69d7Eqt
WxQyUzRqlC/FY6oOlYJRimZgF3nGvz4i+jL7UECMIAVHwbisJENbck365NWWbrqUFcw+dn4YZSt6
BNbabFfwsITrYJdBv2FwP/iT7h+L1uB2CiHncDdFOTgpwyVZndPeSoDIuSocqVcajze8g4fpvvtI
JapMKMD059UOKidUYs7nR2zBpIF+6PqSyUrQqC1VvJrtDuQ7glCaB90prdLPL7h1NUYeq0Jzo1QV
9GJ+OUnPLMAyuJDFDK1JBWXR8E77yeKo6kLzlnSO3sxwewo9QIR7zSu0HLhjaJP0jxCkrGSGVxDf
OGdaUN5hOzaLasCmINqVb//YoblARXJ1IQNfCsLg3GVtZhXzx/bK4mrT9nftBFNBYq/ki8SxqdNs
IJ6slMJ7WyPpQgCWU1C7xtyUsACurXdGZCBWDPw1Yau7ATH7RHYFIxBLR7lClo+TVOLJY1sGm3GB
f2fuchq5EGwXK/8edzOjh/GsjMeLU70EY2GqJr6dtwg+vNvgdWz7sB0qyGQwBHkI8kbGpAIlyQkl
VDgluilhzuoSYXmymeHmGs56T8o/xfxb0fwWzOuqHf7RDAddHmelw5JCclAccgB5TNjTSPqz45B4
S/ajKEv3vxCqKqlFwbcScsB7R3L6h61UrjY+4hkprHQ1Y0bBq5YUCJRRyMu2DuVCUWf4D/A8dCuB
n4ZxLbUVVhKs8mcnCexprgraCo58otIwL8innu9tAloY9C97kv+9KpsuIk3EfN5grTSipYO3wy9/
VD/NDQd9Vv35uFyr62OQThaMSEQwYNUSs/TAK06Fx/7AGWoFUfPWT9SHB/CBvO/d9P/bXtDhcxDa
jPk+V3oAwH+tA8Zp/4YobTRf+4e518XOv0niLhO+sQyc+sj+LOfMNLmohKr0A2bXlkg7ZrQd1l+/
dJq60A/Bv7d01173jA+C2MS/+yTPwjn1F19qFA8Ucp0AWDpP5fHGWa6BvO9m670Jan9XYiOA2O7a
fwwIRtSZelNkZTbbHh5/0B+EVcUElnoR3LlRUZesxiibQKxLxyhs3albNup7XV59N7CPC2zsUuPB
Q6iS0vpWE3HeO1qcUtIzPFiiSt01+jtO0weOyVPtHY3aSMG3pRmQ05tbDu9Id7mQFb7J/8pw6rFU
C2Kc020zyrZjp5nZKibW4ZXagq3zkvvq6vR1985T38ykYRH1tPNdip5arh+Ga0VUzyxGirPUfQsh
/jj0Sq1Zh+w1O/1JsaFAFsLM5pXk+ZH2xd9PA5vcob74Qwony9h/QIIcKdVW0Gr4JUkh4uaJHo9j
8CsJw199d3F9phKzezBwgNKe3fzxAlgPtrOTugSzbyrdx1+qPh5qWDRVdZq9CC/+PdRhwQk1lzjN
rPU7sU14rcjYP4tZTbF5RzOrhHNEFeHFqHRI7Sx+tSyoKnGy/VOOO1tZqHgAdRZFX4NoA+kkqJwN
gYVE3b3Bv6dtgOOkypQJaep7UCWR5aYHAE4VcUzz56yYDhWV+4ac0hloOxmkVx+YaEzNt1omyqjk
tdfAyHftXzlUkwt+kMGUecgRuFofIIu5XJY5WaVhH0YFB8uC6tCo7LQPFoY3TK59kRk38gjap7C/
Cs8ywtz2r8DJZLLaor8kk/J8wnYM3WMkzD1+P5eGRV+yfD+Bk0ggQEnWtXEvA63zAJu/smGfOxDm
SwfK1avZj0LQ1K9ktui95HP/MIikSergGdzVIDo6ZKrXHvhPVA+4tDkD6m7tMn7MccXSyICmCn0L
I0hS+Awz2+fCU6i/Lsm3SDpwhIejX5XEaiRM0djxfJtVSKQC0oByeco2Av0L+6ePQNT9uSICYAK+
rnjw0dRtOh6kDYCgjp0VHLT0E4abrdrlIetKM9PnVMee1t4i38mvaYIEDBNruf/UcU+QgK9BhP6w
anJJ4PgamsJ0raF1aG0242GxYDPWh5QqXL/ot7YTgwQwk4rdLQPfPIPYiz7ig1rslmqd+M2TPH8T
TpmA0J3IjzsINRDpusOXe+8XyYKv4mWSSD1lbR34nNsQ+32mLPcBHj8bjWb1rbTMTwx52xvP1MEo
HVL2Kmd6uo/cJQbFB3twDporz62qR7vFGji579MgTFxDDPm78kP/zajDd2827+DHmGzbXfsQIfU7
1D/VRBPhDRNZKVHrglZysnj62ooJDm1WpNyR8rAS1Egy44z0VnjuQqAUKuP/vz5cA43HsDySJx+b
EGJd3cEDmFuVZQ7tkHn9XGZsvgi2vuUYjNCex/3hzYK7eKRSJbDAflwdz6BkIMogFzwnVwI3NjWA
yNYksBNcs78A/DMKzwerGM6bSoMBoi6IjOAg1cIak+5NGROdkg/F+Jm/mFn7tWI+eaVCCv643+Sf
fnhnh9FQLbI7BGH7wJnYLQnOK4Vc8/jslFMTycL5otl/3pRQKrT8zOYWjNA72Apq2A1p8TfFhX2Q
SJfE3UroayeUMTDrZ026qxTZ6Ob0vXbmUu9hljInpltYJAre4u/jtuQ3Z2wm8JE1GMwWSn5Ve+4B
kRmMkyT0O1g9ymHp8aqQsF4nfXGYMsH4lzMk4cNLL1QyZo1KSovUuK343JhgFco2CaaM5BW9b8iB
x5yRqRZFP9aE+tKZQE1SEuqxkt1vrwTYHHarvLe7NScW6pLvqVWYKpRNIZ5KRMWM65EbwATcsgXS
a6xnzqL7Fe/vle6Dc4sHJ0N1l6+ttQagvixgWYkMH+53P7QgaraXr/fLW+OD+Wg2dEENsQ7PO2x9
uWBAghRr6van9uTsn1OJQebe4XamxdLO3hAn8JEgxzPXfeicPY9vbbJo75VJVbt52X9wSDatQNK7
e4WZzIYWcws4y3q67yrJbE9FgIRhc6H/kzrzOIaZ/LG79ximOu+gTMmFhFhJXBUY0iquwEEgapXE
vKbyNRbxtLuQud4DzP5+opVZxhtxS3L6bM+Gsc+eP4U2Ch/u6Xf0oFdf7IEzRn8PahSogNkJ2RT4
mXb8dvg7yRdOQbFdx8eRHdZg7KmelE0apZuxapRb0XhEDijrnGdY5jFmO/7pmzjWw3utUR1IxQRH
KAxlJZc45g8WqRfC2RPpv7Vw/ARA86PCF68kCabDhjKFJ7NL+gq7kClyrheTl1T3gxX4eE/fjo2E
36e8y/ngIkETUnFxxZ0znsUefxNv/oJKLQuoNn8NbQPg8vZgntITJzpILDYiPE5du8a9CgW8U/ud
f7qKXVl79HpxXhjs7H6kpnGMOZnERTdVqsFu/JcejMjpRg3ziNrV63ZH89KiCRrVWQBKubma2y3D
v6nydIcNRkG4WDHPx17E6IHG5AwPeTcA9/QkBh99juMfFAg2gp3jOaeDvRRCwInTYWiVoFEMo4cg
EPygOsyeE/Lt6CGrUtcGifr0iA27YOZvmtXpiU14O7UPEfAj615EzJ53zexO6Wgwl8u+KhpJs86q
+qNv2zcTWLHpB+20TrvjSmusW2Is/b1ED/Gzl1ESm3rMOymsPtKvoSp4/02KA69Z+4Xiqesks7Rr
vG7xdU09Qp0xu+105fFjdEG8bU4u9VXSaQerHYas9WJ0ZeWv/AodwTal1Jk+2nxvrnO9CMqJ6jGa
dgPIJ6BRMm50hzCU9Vdbjqb2vuy/QESSmVraRdYq+UjB0g8LXZm/a/2GB2BR5V19HYhW6sybWHQm
Diwrvl3t6fxDr4yHB25XTTxFA+DmPj7oDi8fEIGkxONdBO9/bhyQ92z0mHlbVffash25heU5GD+8
ftUiTBEeULolD4HwoST5ZFKuzm2fpGwfeBuorQ/TiEmNyyz1CgzKQBbPMZa6VGn40J7rOi8nLCax
baj7bhI6adoWUnWd9B1IUZz8yhaepDfHUOQTgi6so3h/WJclinD6/i3krBIp/4EfcVZ3vNVgmFVs
hSocrBzduqARb6Id2CypXVyso/nW6y5rjq9FKQ0HU1UtK6gPhVxMwuoWXgGUe8mmfxSYWhBgnHyn
+bAb6nuRqG5Juk8CThx5v29Ke8ryUnRRnOgvYxqJymfmx1KmNJQGyRi+jq5qvCZ80GsTsjeHUSqN
67N+lJPcCkU/+3EvIz3rLnI4fE4x26/1/9MxSpSbFIkFl0Vu/pxmWMzLPjEwMEkxFPZf32DQpdNH
2dCa7cxsCYji2Kv+QuqKBC2+UzhSTNtPqk92shx6CnhHtvxJk4fuqPC03jVQYEmrtSfPYNTDRaeM
AlVksHpivjxVSaRFIoLPKXkP1vIO38njL6jIGDPB+wJ8Z8P6Mm/35KH3bT6guuE1/49eQVbF0Eqb
gdn3UJzlP1UjvnOG/8js1xSd/WiXnD5C4uBHKDKi4YL7VKOIff9OmKKEH62krDYOYRUbIjFhfR5L
1/HpQ7HnCBUEmCJxlOc/lD9+GO3kB+MT5In6ZHzPekneWYpc1pFJmiHPBM26Wqf5qp/fZHz3tbGT
b0AJoDy5AFgF/ixe4hrjJEHMpNOFa5VFxdSzb0UJL7CAfLBhfSUMQ0TEDjorSXej+aTgZll9Jwi5
h77t4Q73Mkv05YWLQEvMMhIO5hrjR6VPMEKARdauLzwm44YBYBoIOUIlSD4Naar9W806HRXpoA5L
REOh3H5u94KlSt1Et6uAzBSDc/5SFBw43c0moJm4VroREOFDlOF6XCI1uGwNgK2r9gueU99qqH2p
mq34jm5hSpY8g8add/7mTXubLw/lEbsB9DS8sxG5zuM8WqcUX4DlU1yWi7KcELTkXFAotSsk92vC
BfP+s3+cxANiXHxqR6gdjhz0xirTJWrepDZy8JPqHsCe6CuY+OJg4Ye55DxSrhYU3BwOSn7LjcRB
JnKjc8MkG+incclgbTm9wkjg+Dva0FNdnMTAPr3YVzOcCkjtHhpKZlr3l6Mn8wqEIyLA3w5KN4en
8txSFtj2RpIaoK582+sAJLLLm1DirWk3ObZfQf59ZaYCIVGKON3N2RSLgkeueEk2h/+ZP0BDOhL9
lZv9vmKz7R1GyoKZUZRP94iWzkwUd1FufMYxmdrsiqoitEx0IxTV/nEF02nGOjlCJeEVYTm+sYJo
xaGnj1LW+VFJzz3yQJsDZWveFs05Ww654ekBHs5QJyLXSEhlKvS0npAkGLxQF2EUbw2zplEHLezr
rIH49XeAaP4LocXgmqyxeCDAKa53Ij2MUGZitrYM5HDpl/bM9F6BRRCQiyXyTteOJc78PhVgACiA
AiltbhCFULgpqX0Yy+10rUpdd05HOzLoCsZlyZ5RGkRhb5BdK8DPFzHQZBZuafyKXbtqk4gyNHLW
wN8q0KjZ+wzjhmqQZYg1Xt2piAkaJY/QX8QZU1+ds3vbp0oAiiUM9penPj2M9PzkHoREhDp9Ax8G
wjw9BNh/M6r4aeqiV4IkLUS7FEq8XpUFF8KfZJjYNe6rnvYtMKTVoDNj3d5mXvW3US/RsrmJna9c
uskJPSXodvx1oztuoOVQjOJA5/S8d+I7yMNXP/wjIQEeSpLeQOnzxfZe0oq3H1bUxJIOy8SR90xC
OXXdiQgYguzcuaJ+8himBsrESygpO+QKCS76DJfiXFI0YrzIbYkuYJH/oMbcVZwSGvkUy7Ywxt9B
/m1fjAeijc8Onba3EsK+mbErf+W8IM/sR+tceTWzoZwnsOVmiKeJyM7X0degmJjYvCwtvlWsRG+W
ZZuB6/PBOXY7cf3Ilac4KHQrW/N/kfdJjXdQQqpy9p0FIKrXJG9wzUhYdyh6j2C4jeogMt78XM/c
BDjqW4nrA+dDLty1lRN5UfjYb04yJrZ8A3ACT9Ai4KeE1pqAjzeywNv7Me/Zel+ToEsdyt1Zi2KS
CLGkbxNPjJz9tl2yXdZdsy7ib7hYBiE+QI1Q4Nbiwjs3IHWQDj27A1YRI1WYk7V9D6chw2CuaE7F
qA1r8XdNj0gwbQG0C5jnZHOr9SWIxGlkqAKWq+/fiFzegyCaCaHuxQK13KwJlCad3a3WWEJBp2MC
evRF25Wu7PZYEszxUMdDSGTngfIUjCLazcQS6udHNlGQIRWpaCmvl6SBsxEQSuUx2X6UqJAmyxpe
0JHMypwL22VDQqz9f4CYABSlOofcgMz/QG+L2v4+JAmhtfrF9JdcBoJdMvD3M81yAMkEEal6SCzt
8pnIK8EyJSvlHTKqUKSUClnCRIMq11PpSCIh4e/0/M3n3FkAB5CLsiuoOy5x7OvqNcEqZUCkMHE8
Kh8zmtOpDkNyGubM03BnDN6BpPgFR4Y/kc0La/SAhkNyp3k21ePbwTlrXw1IsG/bcz2q9mfkAVz1
iSkd5qyguIlPezWM9ny7sCXvuOsJCqCuxkdzv/FMldVfSey48D8xQ6C6OV43QqLIFF5hhnfvK2oR
sWRbHcxOySa45ihB4OOc3JAF1yz7Wt2lOs/yH9GxGk5N5BTou2szAkZQEh2bRweKy5eb/WNDUdv2
ZB/5j3ukSqvqIydIpvOagl+ii45TusGg3WIpUSpNV8EAQsF9vat9N7tGvdQwJRcg+rNHdfO3wHc/
YmlMBJpxSdc3woFrt+lE0d8id1BL64LCrpeIJ+eLGNl2TQui5KFwQ4ojlvk4EbY7iz3Lo/wvqWHv
pnyKLoM1p+1MWfKplwswaDkKe28HcylFZ9Woph8PPlsWx5W9kr28xpspXv07I7T198y8tw8V2682
9CXJWaL35GPSeiVbzjE53ju7dkP4ojS46XSpIhEF/1SBxQXXY6DhDGQ1Fkv/onwsK67LEN0pEUvn
R2Im2v0BlHJaZuZvOzDviuMwkiXhiebdVWjolS2+uNw1cMVZSsYwt9ZimKvxmMKHV/7LFCamSnif
Te8cJhbFulmeZyuMoHtIb0o3cikGyiB9/SAsz2Oua/5awH2ZZTvNacKagEZjxszkNBneAoDAtnZP
PG5dyeA//Var7NHTC6MdVSg0yq/YOlIOZ9wQxiYJZSj/I8Z6jgTgGs0a/Q4G4gCo8lgPijkt5ONa
/6KnAVFFr6t4VhlNrRoUMv491lP0KcJ+GPVusIR7dct2twm6mc+l64qdAcUDhsQLS5Hr65gTUMBN
SXMUb0HtO9ghHoe/Ex42Cs9SfzrQhtfj6oM/tVFBH45FsZ9uIjxBofQXqU9yNqHTPTyDrL43qfof
Jsf8mtqK9urHTq12KnlhoDVwCbW3Jwu39v5oR+2Mup9xOpQpOW8EPwpA2wxnbgoAy/RTaGEsgCAX
wNC9SVEobTJgGHXusiBIy1eifWPawEfadxcUkYRNiMY3j+bfo304z2cTGMdkDr633cleR2E91xwb
iuZXSzzIa8oaLpU6z0JP3Lk2F7KThw5rXcD/BHUNNxggvXtCfWSHs1hEt3aR43zH7AEA1moSOIdT
3HIb63JdyNAYcGufnoNmqHSjA5+pZiVZu9UA7Yh4WgawXtL7KPtL4DjInEl43vsMCKZ8+qFk0TIP
fdF3TltxqB8nH/yS3whyR60NxtXY0KzJCF/LuG59ETz+v2HjxogcEwNz3vUsiVysYTPkwM4it/oL
P+vagvL96+/IccDqkWzKc4STHVn3Syktb3D+cRrlhYt09u2YzxrrxI2TkElmri+61EJyhRWkGwvh
qGIGcZq5gGzOyy99MNLyTHICnHWSWldMW2NGI0zqxr5KvE7peIMdNgGVCVnl5TfoIHcSutrjFwN8
0BYCkD6lQ0fPgMjPM2bIXGZy3HLb9VEkWXDae4QagfuKE/7H4z6PrFl4nmNYrOLmjgamUrpavjEP
RDCc39yKdfoBZrVSsvpCc2HL+R9W6DiNtkPlwln56W7QkI2CpPk298sexrTPuMSeglTEkcdt6Q+G
OoPFVdhb4eIN+Ekl73S/6d/2Gb7W+0HLb+zSz949XA715wzvaohlKRwFejn1JkQbOGzN0U93gkOj
OlrTfGrzHY6GmcPaQq9CEAzibAPM1RiuiZOC52lnNSp0u/DN5z/2tcLB8VL/2j+dPEglz3YMvfiS
LG1nqlhJdtEpXMmZ90UU9E8qsH8EpWXerFVtdiu3nEQIMhufkOWZFrXrFHYtgIF4gIAbmdlI9bvs
SbuYehXo160iJtJJArjYyhXWmqIcdbwrU0D/SQuCVBRDPNyl06ERbqL/PA66nE46eTh+aP/WHjJb
VYDWd9AWte883f6pUhJQHESvN7P54X5s0dAb5OvEUjuhGzEEH7KWe83E4L32SvVHk5ueWyjSN+gi
VydpdNmrJahi+J7jG5haz8ESmCKtbV0PcbkhU9Rx9LMoOqNREZVe7E/qZFLILq5d/NEM6MDmGv/K
eynWoC7GcbeQToh01PHlUeOD7kxWu2u1hYrkuScxF9o+Y7dYEROqeiUXImSnvs+okcpt8HOuLYf/
4B/FmNclzpB2VGBDRfLgmkor5PlnaIDl8SXnPTNxzeCkfKFNntzKfO0bR3FSP64GEc49UnkQhkTQ
Zp7eWotYYSbV6pMcrM+6Qj9KZ8WrQ8y+nnKNuQ+myMejDrKLqbKl9Za9o9K4+a9n+Os9m2/zkC7i
ksgiItHof0m8/HePNyKS3YkIiomvbRkMWOMZNr3g6Rb5MzlBW815Bc22shUliBCT2PFh+FVeROyz
fPFliYYY0BbMsiCs/MXSUCmcSBfa1hBHMmNYnuhOz25thl8pHwKn6urg55YCuwXo5ERrVc83mOOb
2asDa7S8EKU6LjngBEcxSv+l2iLOvVj3YHa1Q8titkdj8WTPzzuDI51bPI7WK/D8BjzEQ3W6CJCQ
LvosoXrpR5wQHu9Nzf32chDo3sf2zUHBcH3wldVjJmN4oId3QtFXSPILsJ1d3j2VNPNauzt9ezgT
L4ty/0PNJtFEAFT0UQ2ZdCq3hA8MurtCEHcvuuC8lW2rooxckDuLSsKRcY/pZMjZ7DFdeJF7AYT1
bXbSgMAbCUbbEls5gCIBY34HJHTfGfrv49uIvx+HiPE6bcUWzUvJ/EqFCRVXKlm2vjePSdfU/d9b
jsJl7kGuuZ3a/EF3PXRZzz/kvk+9GRtfmIV5oGLGKc8m4R8pugdsGOIfYeOquRRMoat/zQGOw15N
4TQK1EFiCr5LgTGyWTVgSLNviKxjhYr9mgacbjlTgjjhdIRNg/ainc/gFYkmruZba/3kyrqMOrue
ia7nzX2WAlY1ojaARUX6NB6g0d9LXJajblulpqiEq5JrMsOxjIR+zb7CMAz0vFANRLxX2CLNpkWg
6c8BsoDQIxUNxlIQKuJUKWciIn2eBeaJjiPA7p3ziFNU4WsdBfMvWC0Qdf9fLeo6U8/tzZBTHGhd
9da8LvUKXGa0oW7ZbH4DFkgeGsIxxLTNOzy/9TCrjLyh47OrD1RimrLdOHqdRk+eIWU7UuO5yuu5
f2BYwH31ep564Bvq6VXHi6y6qFr+MdRs+UXgFOIAm61uAF7mODCvJnRnewl+iSatCisV8jO3RYus
VC/HaxG4eeI/D5gQywavPp7Z8u5Z2m/FhAQujwqTIZM8xd5Z1nSLeMOqi4kLdVdPh1932pDeXohY
/oY2HR3skSuXSLNBZ1VCxSQgQLbcrj4/9VndGppuSxweJys6EKPigeyeXdPhDGYv6zNneczPbWur
oxC//FJ3ZGklwxD3f5CGRFijGUisbMJ06Z+wYcgUr7p8OYSwrVtc6ws96dXu+8Rbiuq7FZ/feSBN
Cb2wkcbXZnqRjBnPj/XQmaJA480fq6nY5hB1bQ4lHcI8EU7qJ9t4O4jh2wyBvsbssCqh4O+9waad
rWXaBxSAorXkrKTQrYmYB+EiiesExFMiL+WT8dFfvtPpWu+TXAwGa080MvO5Rxl9dUa+f8LuUtw+
grVhvBbTzVcIL0Xkf+eyayQW0uhpWZvylJn26F56toYI+9ZBH+SiRgcH4Th6PL7wXsm+CD4/HoXT
cK727/B68bbAkeN2cdxuTTcB/pdPhxFHyeqz/vjx1+Jw6a1sJFQNG16vhCVdt7CvAEPwwdOS5PZe
NOTLAdXsMKKlv1drefVS9pR0gibJcl/GvwFzV78mRtk7OlszQCmxxdstYaqxaI4sZJWlpvQo1yQ7
d5+46Fe8ZxOkXt0kZY4AZCZ4NU6LsmPkGQ4utNcd8r9biQ3tky2FYAnh9E5cnMnSM2KLZWI/Pi8b
YyIatfnAWLGB9SfHjo+Gl+0+sQPgNvlhbp8jjrvrabA8dlztDGWdbAgE/2aQZ4KEXR4QdxnnJGmh
MJbKSgTxVv40Q0jVWJIvFj1cY6Ro2x0k4v+AA2Jq8u9pOk1qtcYDIBNFIlw0I+EK+ybH8PKVbkfe
hpj/3JNEDIMtgLHRcie1f4j/+r7b8E4xqObXwliRlh0Px6klKfRR0wn9r7E090SmYjDCzYwA7D3M
ujVqIIzW01emAzBciMJIJaV6xvdu6pJCw5wF6oV20XYT6jyazlLWJnoL1LwoWB/Y13lTgbxSp6hK
0YsY4Cwasa+kW6hD9m+GfuOXVSTewvHAIuZHiZJqibeXWtU7kP9qmMf1uu9nwfnBaHM72xbuHZlb
HGc4PcgaC/8Qwe/Bjn5ljNzLofJ8azdz4xI6rU2W81FrZDfYm6TP8G90hXQ57PnR8R9vatQfVUcz
pnrOVpJJUxppjMj6YgpgFruUah94e0ouoREKGhwyaCZmQBLSdk+k6h7zTjC5jkGanPBsu0M27thi
YRrYE33wWIUE4lOTJygAjV7FZbDwQn6f2x+VLwMlVQWF3IqypQk/7fnoRQm6Nry6NSpByYI3Q4rm
ahX9zRMV5qEFx/OBxykVoJSwFCSSxZM26cP0y/P1oJFB+XCiJcy9KgeeSN/81OgtduKsby3cZAiB
idqlcsA9cremMhmPfbtrgJMoVw8AbbZtX+N5U8/KVN5xj7dFTchnsePhFScAY04JgrSgSw7cgonw
keKxYgrPqwFIlUOc390ZooJp7B2HmLpboG8ht9e7WMaMBRCb49QC/L+VI2eLu3sEa5TtAoMqTcvx
r4AEg8I+HYANAnL4k0eB+CWuB/uEoNim1UGgYgyLLRSYGgmkY6EVzn3Ye0jG9ShZyILWcI1XTpC7
9BI08ZcaKpkmOxFl/sPm/k0MLGlhqMvxSu8owhY7G9ChNveo7nfn76GESx4ejJHEpnqfYDCuARjY
mexZmBp+IrFUwT+NwG1IbLNGvHtjZUIOKdXsWrgOWhYgTXKrEBVeMxIJRn/EyZ9Vy5ksSTfwT0tu
7pWKgm/Vw+2LjHAlRWPamg4K+hvqFknFnQ6ZzhfQiTOkSlktmlXC25wZ37NWcQ+E8e88+YkmpCKV
w8BO0Bv5lS6BEUGNkq//K6qVBzxPKEw7EXjgzFZcZDU96Dq0WtvKiRzysKL+rNeaNYm8L4s5rofF
xS7SC4x9XWf3TCM2n6XvyHWRuNRQUqP8Ze7rDJ0CXpeXngsRoTvN6/A4s8W4eKwlKmcndz5gUcl0
H5ZztNLlFBTUxNuT7ZxbJjSaviUrkIjv1ee2poQGl+gsNhXwWM38lyO0V1a6EvgFACDfgcXT84G4
YYxlEWEmplETwoyXt411am2IFpw9pXbH6YwOyGiGHaMHDrrXHO070mrLn33FZJVG1Ii0I76IJlvh
ozoJ5/8eww3q/KM4Etv+UDLseDr2ZZ/8zv0xB/LTsKR51SsgzYCGD6ItsmDXUfc8Fsesa86+UYmS
hnHyDbah+3/vnTPG/X8vPYDwTtFqf9rAusXLnDUwtU2cKpT/UFk+W9O14nU/XrX+XIIv5Fsyq7Hd
La1mfJDLtl49hcDBbD+XCvF9bkYK/3CeGOpuu1mIueA5H9XCOLDqNI6z4ZJExAbMA9GISYNIkIil
/W+6yPbxJE4AUgJXxThE6VQF60v4CMa/0Ko7n/MsL7M8f0Zw49FxsJYooZF3xnHf4Lw1SUZPZ8RR
33lu8JE0DmarH4Lw9jFxD1j/7FH4OmACJ46UOTc0e9THnpGhVc4qwQ9PLQKD+V7XwzjAH6qbstPE
AV1KNUzYKi/nRwEDskzM4Eai3hrU7EQ4t4XaVDUSHsXpKTlf1Fi1xyK4EUDoT8R4npGL39HE3xN/
VCVzqZ+OX/PGRUnEm9+jJu6TpNGPMsdUGnLQuN113JSl1EfR4+XfXZNjNe50N2zWVrTCDRIdJScH
VG+45j38nipCy9IezoRFwoDJjIPwF29HPtWOo07VU7//f2i1yPU6SXSIxaHPdKODnJ5fdB5z1IUF
W1eezlq2FAmY+KZRu0iqwE2tTr2mRDHdXekmRvr/l1EbydqQDuEASmYN2yrUEc4fkUzoJKtENHXw
G22ui5gEtb9JgFM3EI2VNUW8WK2/SULvZmDskO3v2ii22ldWzTRgPSc4SeuO2r/jyXwd+tQjMp2n
uq3blfUQe/AxQJ2WsuQTmVvmCkN87YCT2ayzKXiZoeVgNwNmGUHRdnmAMe6PY5W5aCKS3NTfUmGC
Fwh2NuyXCPPrG+aprtrGLvCAwdVXKfRWyvWWRgKP2+XrJvkT0sOWx9Iv0/a/cDcxlF4tKMwf5FUF
7prB2e2jwSD7R5stSZNedkcKNII/flrpiYwF3dHOC+RHJTyXI26AmXop3A4cf/H+SVjWxnO7C0lx
HpgBmgBIlk25Lp28x3wt50EGyujTPGAIa57wOwR33YtS/rYowH7x7Q8VYsQiE2/zC+3iCGWeQna7
Nj54U5HEksCC/GeTOQHrp7/WN+lT9ItACdJb2GLKfiUVZcJxhKhZuFegGESiaI07Iv7F34/obeHW
4z/hg/xftan3fAZ8jSlgsryfGY4Nf17XDjYj3S11wwV2rZ2XjgLtux+cLgMiwuLrPl5jxjXNTTCG
FLsCbBLbeuyBSfwKkbu8KcLZkQ+umYehXfdv5pfApmH4wx7FPiarX++ndbmAuZiMS0Nq/rZY2s2w
RNoZbZNHC2bsC91pMSTIGJVv/l8dEp8oWwHUWgycMDOnw2ut1+ohsVpq0ph6nZ5VzI3bgSUQj/sj
2SNn6RqW+ObFVc/S1v65Wzd/nMoB7Gla1/SyBF5p53jGMJE4HIAqKVshlRg1sWBCH5PN78dL6cej
PUdKZwzW+Aq7fM91fRWVi2s72SLECKdYNqSLS4sNYA/picBPG9hOUP+hPonE9RqiCI5GZ4LSDhRQ
CaK+AsBZG81coyXu7lVAoJCo3reyFnEb6hYjabblNKZozQnIBuQvENrlJUUNfQpU8NLnA6hDIR3S
i9U1m5P0FgY1nscmglNEr88Cc9vp+1KRKS2YgNVadT2Ebllkk5AbsnZJNmqO/4iTt8RoPVMh0DE5
AVXiV78JpxGdQhQz2hY3ahQPzt5crVPknuqBsSFZwGaPljGuipjkmE6TUVpzwKj2ppdEmOPG+HCX
Jg62T9h3PwTz1gXJGKOaUgj3P/BTn9qKiGrPK7tKR6XHwqkRfKkK/jp7WoEU0b33j8uQCqkeW/6Q
Mb1lLEma4BWZBbbYrTsk0j2NKiOt83Rpecrn0KLCzDn0Folvx/EtI4/qty+iqZcbtjY3CM6vLTLt
T3KbhMJCpTtTMT8IkoZ8qa5qbPQPdu89FzoYvq4aqKCAepVHsnBvNs6AF0GD0KOF9Lw6a8hwF6JG
EHTKoLN3HUvBmsjjrdJAI4wKKhoG811cmZXRZmXeD8GQ0syU/9RyuHGwxEAnEV6fHYwU3S41zl4T
srOv9R+O1Iq+OUUthYHZ0uNzHsF+XwGcA9cvKTckk2X0VABSluwvK8qRNKaqSd1FtR7KZ/RigsV2
oXY8YcdxX9yAfHPD1Nj8lHlPYmdKrHlv6TIYE/SWOojv45edtKKjTH6Nm7th0hFdFexch1oHOAxT
VMiGjXQSt0SMdUCU7wr/BqtWn5otnkSZ2o04F1AKxdkVmA4t1TRVc206S3CPosg02rv+hqLQwoRi
Sq+IAuMQ2aZ5NO80enGTmiqaBNPWGU241av9FQYhTLERa8UigkaAGSbkCouPneLcCem+SDP8jx1M
5WNbesDKmITlTEf075M75HOxhrINcMf9H9mxVivZuGCI36Qq3cBRtpT4Pp6jTZLEL5VZxtK219Vs
0Cibj7QvUZJMfwZBwsC2p6CKDTohdCmESjhYlnFtb2D4t4Bsik40UyX+dv2c3k044kiML8qbqG6P
U2rYX5wo7eGhEWXy8r0mes8HDCTqcKYLi8UqE37ruPHMnNWnl+22PlyGa3YB6PsqLYIsjg7F590m
gDk/SbfpM/bqJK4RmjaSGIs2xCdZXRvNQC84r91XJp3yKk8+d2951aK4TX9sYz5YDhYumOvrU8EC
17eJRKjWy7oNeEFTez4VqDXtN2214NSzIYurSmGCRKL06RkIuyOEA6KyLiVDC+JutEvOMUVJeOMl
zK+5q0+20/2hSNHxpPacJd8qMbJ5J9tgComZFxzy/E6PIV/bcOOfroRz8RcANiceX0b2SMsVRJR9
7OfGLgtDA6EWFtBQciJ2/1zsMyN2GH6JDr2e7I3IXdviXtBiYCetxnmH2Ylz6iUQzzh75fYoUsyV
YZ7yqzYjXCLUCQsTJbKJoQ/ydN9Q2aFhfHpPJqEcCLaqPjGhrfZ0cwTBaga4rH98VPs4HlshHBS5
/TOsliramE3+0kfullw0Dt4k6U5c1WpMgg3sELhbj/Q2YrNPMtRFbEY7ZvdcWg5xYz8K7MMSSYUW
RczB4+6E8fBW/VE2mozAIcQhW59T4wGnUtlo8W8Pj3EGlwy1oqr8+10uTWu4GEz7Gj8pbh4w5nAr
z/pwd0+lDCf46L4GpvefvETT4G5hXIixUF0DB2220CNu2XjnN0LRzSdvkT9TrPak032aMfTnivK3
yLrI93pZhAwj8W6OKrflfTzVp3pIBLn0a07AfqCR5TQzbQW/xSbsLJ54EvrlIgaTJJTOKi25EhnO
IYRNdpOg1iM0ssjtmnIDLyilcl17gxrpZuA+/WjvNBSj8c7EeZZwBMWkznuMtLADpzkaR13OEPS5
QFokgIiGbYeMYYsywy9qYq76poISJRvo1SBTE4rElHYT3jDiT9wAGW8u6PP2EJxmGZdGu/vNUY7q
0Goy7az0Zn7ktCIrT7Cdxs6NSRpePui3HRV+aAi1GpbGJJKt/G1YssbbtHjpSmQF4/GM31xbJv0f
vPY3DmIMz2ci6EbF99goe54FqSUkKzJVeOadIBkjBNyjeAl254DDesSkwJklE0aISUjW6r1jTROm
c/m2aYM6aEZ+NCrzQD4ZWgg6Y9RttTveSQDgV64naApisMVk6MKHk+qVmf5Ym1UG/J1V/3n/qtd4
sEq1DqSEp7AOFnk15hI7aJ3FMv/Ux0qrb7gZcN5if+qE6bTh65LOTq3bT9i7mS2lbH03XPe1UIaO
lNjwqNch3ZXMBZwqJUZm/pCo1jJwt20O1A5hto1zFgtrfLgJR6m8TX++2fdb1f5Je/nH9HZXkeaM
dnwe/LujqsXUD9gpap1NeStNc9QBNvJJ7V5cuGkhfywSmLed8iM2E7EFuJVarDCb5QIMpsXz5tSB
GHkpjK0kVzyVT1G2ST5+aImVvIRg+/CZCSCtPjuBMEkt+a83cwFujKeqWPjNu3+tPy1J2zY+KQU7
LeawhNOqjYPyOJ0f31CD5OQoPheLG8Eg3o41dfdPEd9vYpoeORQMouryaqKxooRDUh+gk5hWZzL9
FGbEZ6CMf+jmIit5ipfMdwuyWPiXnjcDPxViiJHiM7iIlyERB9I+bCaZhaMSQZyHoaT+pFZ7+Iju
fMGaeYa5Ulgg2+J0p8ZVrBaKE0LFDVNvksf9habNzCBMtxJ91rPbBRjBuglhk4ZEZm5ni+OrJkMf
MV+5OV6QoE6R7i1AtEBY9muJriZY3O1N3eetJceDWXOSA/113ZVEaMICO3qqO7RmyoPQFjBsKF5P
FV3sT7M2E/+DHrJBJ4LwtXcs9h5beNahbvJFCkLcrVCIMev3ICx3wLYQVpX9q6KcaxOjh9Pvzk5z
gudW0sV79SPGo7VEYzB11bnfaVkAKUbC29pryrRDw5NwtyYLRMM2txq9ny1CBoDcU9HsRiHJGS0f
+5066p9OHRQudFdnEpGZOooSXhr+spqjd3qEbXb/LjPPFXRD4ybgQ+Az0DO8ZmA3icZDxDzZAuIw
eta/KW4GxYobDxRoiMvoYsYnnByHWawI1/lY2uiEiqEHLOJFh+EEXCZW+tHKYl4FAdjBBjxVtwX4
MwGxv71kCVGg4McSTf7xg45qTCVgLEwuXkKSO9jSqb21SdmcTzo5ulGwzFgrYS+Zx3YArMwxcMCE
unxK1p9hPxd7XaAA22nvXCXIYOlys4Ju+HEkD0EEeB6iTU53t6fmj66YnWVTTMR4LKu/IPuyXCzI
XM5KK6LHsHeAg/nKnwnrHboxaj/lYTM/OAhCjOnB2Xg7wjePjHh9qSHwaBiOl0qm46xYNtQOsciX
0Fe+AC3esyk2DXL+gkG9J1orhNlx/HdpnwLQe2ZAMDe7qFJp82/mNQlb9vIpmf2LrAyCsztaYZJI
TrhbDpLh0r3x1l4F/b7xZyC9H5OxrW7FIDtzIo1mpDHJvmF1RL2ArUvP0IGkvICYPgmxHLahFSR8
wIIt+XggIu3jFBHOT8bujnKepi+1yTjNJISWgOR+vgy7A/sMWpUWJ2D747335Y1HZQuBHGZAEeoE
jtdm+W/Wd5Udz9QwVCUccvU8xQaaxMGSPrk+JWKErys1YGZBskW5yhHuoY9DlBlht10gZ7wzF463
IVnHeog+0e/9ugPTfMyTjg1GbIjHt4/8BDZcDFvYIPwCNfN9t65JOikPLC5pd63wow3smoSh1d2L
fDZp7KXRrDzJ/Gzoli5wEluMdB6doYJVgsCvlFfNDWRXLVNgkqOFRsloxfKddWkEV4EyTQF2iAsI
xUYiKCOkBaOL8cq19gM7rVMLPoPYMa4yx5NsAas/8aOJ9w3sNzxM19myHtV5pieWc1p0Zz420ivs
9HLwYd+KXu/LdR8Oo0YIfi6DyTl7/9jyMLAuXipgZuRKCoR1sIw07QOY0crpEiizKIK/zixkw+Er
OntCVLf5APrzyFjF0DM+6DPTy+1A0S7wgoNN8aX0id9NuvNJkGPlImM21VtQc9k9Q4ZFFaeJknJc
YIqgsXAJHsx7CUcKSOrS7/30nw38m1gI5Maj4xIP08iAnBHUJUERTj1XvcwafulmOCav+L5e39/+
2dXZwUWfYj0PPZfwkjlMQ2rdeIq8tgv/UR1O8jtK/t5YapetsMlydblsS9mWwBHngLQW537Ialty
sf8sZmvVis2KDZpDW2vmJ/7VuRcAfD+hUmkEIFUWdtrQIfZtUn5A4dYebTvOYlg+pJjkugwl7ulF
xO0kIuBRAvili6KlJg92tNAY767SZnmPm5Sy+4frFMze31nknthfP1JlAiPbewYcLxjgbCKBmieg
BzuaTDnK39OFZ1NVXsgQf+Lt3uOoDqY55HAogxqz0PQjMuDAPpRcQD94tpM8AWJauO1FQwQXIXy/
vEUtl2UXBuT5UeCFzjMyyR38q4fU7nrHZ5+qq098klQK+39VR8r6ep4hyU/BDp1D+/2WprYnlSxi
M1egWsjyPl46Qt2SD+0MM+OE+8O4OfXFcKQrnx5bWmvRPCcqQL9JHTLAEVK0f81STMatxTtIBibY
kptD1wW4pNK0NCdPNxdvANeWxU22GXasV0H5ZdflcfALeh/D8ihIoH3yzmaWl/Dy6bjM7oWvDdlg
9d+Z2chNtTxFOIZH8+SKRtvLHNW+O/leC3uap/LB9qewJRl8hrqgc24mVh93R1dplTAov6xeR67r
ym8o41Ex9TKPXgbio4LUAEzekxiul7qMgaLIey6aKAyi6KJIoE2wSQVEtSjZcdubkfhw8E+r3A1O
+7WfZr5GBjV6HpFpCHajS5DXt1QTkLWzbV6awDJJX2rd1P42ThSe/XVzhCKGiyyGYE8qUJwamLZZ
x98/0+s1FEavT6i1VaBeZLttXH/XQV9qLobFkEXqgT+KrYg/lOkoVm6a39S6avIBipuDg9weKMoj
s9YzmPSfD3HpZLI6hNjICZvpp788RM+I87XwuVTfhWexl5Q/QBQTg5k8LWPJiUuxoMZXrl4pFEk7
Q1llsnoVfS52yDSIoRDusdxc51iWqox2anvX7K2zfC17PRDXjunim3ofKh8ET1osfVCnBM8HKKdJ
ftelPkYQ8SJa4DNveR0Eehm1ZZkrA1RmgCsWbeHo/ULiH4zuIct9Gc+aB1bUBqZSLYHG8x6NA79g
cDDoOTUGiE6+nuWc7bbmrOBhGEkG8Bd5rMC+kEKSGz4QD0Vk0uG9sk2T1krR7CGhDyfndFGFB4I6
7JzJrZzG+8ujY38WbCnlQnCvSsGQEdm5kbdh8hFOGo/UBattRlqljvGN4rnHjN8mbmHXwNtrNtCJ
s4sd077JjpqD9FwY99eCxtZ1nkbs4LUC8n3GEp8lq/E+4bYTunCew+9OO38PsBGmtfKqNCmRkEwY
c5+nvE8kbokKGI7ZRw1wUJrG0obBatlGCMNPStigGp2H/lyptWoUeLyg7bAR7CGTNvk7QwTgy1VZ
oLw0ga7Vm9hCTqAH/jl92CK2V3Ggpyw7ClZg6LcM76F8l/ri/7Nl9R8ZcMduvbB+eZehIXf8prFr
dbD5AYLswsxrVX5DOjpZsve55D4LSk+M9lPSR/JeoL735XHkWx3rJ7JjZDQcJXa+fWV3hrlctC1A
qiWfTjqiT+iDQ2oc4+TijUmv0LVYxkbJEn/drtr6yDVtHbHRSVJQrhJ2TClEzNzORNix2e/somoN
IhVji3xYV/xefqt+j4C9kPJ8jAI93og/s6AeoU59YmUDdeVEoDSC/WXFptT0W0ownCcb+C+u+kbT
rG42q3WPf2l7S0cXSWDETKf7enX/eMsv/a3HXPRJ+dZmsNItybQTZfDpvHTVB+ebetMST5l3xoFo
BC6fD4R6vwjTlVPPTopKXgIDqU5ND8ILXqSl4E4vpE0an1VbGhjFhLkxxIGfGUeZyEBxjYMfFgWU
QXlQLkZziDA/xXUawYv5BhX+OvEjk+3z6BBENE+LjsWUZ+Ql27chB9Nmp2kttF3KIKtuhrCOtDM6
QY9KnnBSuN74hAuChR/fdmwoCGxBL/NSbr6T2czSh7m1CUvpl3UUZnpWKYTZ+xCk0JrKoobN2v1f
5g+F06O0t2g9xBTiGmogPQ/nsVpiveBxNwbV+0ZZFosxzGB7aWnbhf97fKx9v8EguBAqybRgcBsZ
zmSo6CWWqd36iTfvGDZKzy9JJn+bWQwTXSaduoLPPAi6LRffFHUTlX1qFWl4iGCKnxX75usnpwwU
MspXt2WCAFW6vegVMeAu2RGHZjI1HxA8OILwK4yv23h7y5A5XuXTsje9gaSbXK385rWsBlCsJwp6
y6DsLPs4KRVq90wmMM3SLvYZWjnavNc/sl+PxMaTa6PgMoJF436scTOA2QkJ6ouBseKkV1al9RcO
Y3nLV4U8mtwuhPXgJperbShsfTcgY9T4MbqQJvDDSKj+kEmai7gW9ImSjAV+titCz/3MQo76oo4C
YuAx62MxByOPilIdukP8bnmW4AQY8ycNPRRyF5JanCbQzxuiD/iyzmkaaeujoUJgQs+9AC5Yqj6Q
qMXDnfztp3SmM+Dym4DsYuKR2krbiajtsWcctUnkjyiePEC/G3F933Bk5iAo8CI9JJHxLfitKXm4
S1Q2FfSD8GJPLlAQDhSNBggkQ6NL9mDXMz+1nx0UbgvhZQkCl63GTtsm+F5SGzra9mZAsYiTc5f3
hJWIHVOuHT/20WnXK56DLdEWrInguh8Du5f3D57m1wPLTu3xzndcwIxWJgG+zzgo9bQE60+HkyL1
fxjNSK8bljCOJapnlVxhPn3F8JMtQmp45VnNC/700lVhCqKglxIuyqd1AsS8O2iVfS2S63NbYjNG
TPVHvctazpdGlCRzVC7szdkDM4xYy6dx7ZVqjE4blxCP2zefsQSIssflPx0d+7i/XIwUjFwJb0QZ
qUQRlMVf+mW8r+0NyynUnLzmKv/ebYWyn0WVJoL5AQokYtUbZ/XdQZNCZCe2um6Fem7ouaQG1dN6
uPIuFiaIjGsFWYf2ObTDk3rPDEUWALIjH1agbcghsebQxsff55O9j6XVwrz/22RRGczCX7FGM2Fo
mQEv9CJch7Ns6PEPdubD0oys2jR7IQ2MCu5u1IVTinxdVK4EgR+TBezYPJ04iUZe+EGfrHMhbQG+
3xKTVp6BnYG8XAWEBFlwXvFCGyhJnlqTPc+s5Clg+Jp649FEKUuwOrRv3pjJVCd67lSIISWrwbnG
vM+7E6XAURsCjhd5hrotYX+wSUr5DyrU6drt3tjCR5tDzWtd19ZJBsFZnotzjRynxOrQEkjaKz8E
rG67ere+h1/Go0d5gV89YoyRiuw3AGADNDuAW/Y5nzQ/tX0pHrPwYbftTO0Qm3t2AnOyezXZrmpF
yLsjqmE1Tu0UUT44rKnqV2mM5nvCtTANBu+u4yC0ggd+bNK+RFANrjwNpJo1BaPa+D5iO+Ch0pyr
8xAcc07J76nZFmllh3UAJujxcmky+KP5nqlgWoEFwvA1mL9H43x1Vlw7BsRMTO9+vupfAqiy/hv6
tb3m6goT1PI6ljdv5/akx2i+uYgujJP0iHpvkO6VqN/JP7AkYCptiCpHO5iV2RvKFbtWUkbMUvcS
5ENZ2ZiRyQbbdrr24K3bakmhH8l35F+V88LHlPeHx8p6/D2QkI4Na7XIrOomlhZCCl8fZD7dy9Ae
OL7OhjdhQV/dZRnvqAXQSsGE8i0gWUck/Tld0ABUjEfXpz5ee6W91100CYIWrCNeqH56nh2rSZt1
A1zm5zV5NK9fDkQXYCMKLG20s4+Xpn6Cd4M0dKrqyhZVZ9RE3O0r0Qk6svrxlIlttH3kQr1Os9CN
xLXLZW7QsUolmwpObJcaOj7iLGgqr4jdGnzvwnpke5gvhbYxBrAtnZhUbg7PNnk1xSncn1erTRU4
hfKPNU1I39LCp5ASksf8xyDGQD/QU6CGErtpfGCA3pmMrx45ShqNxHvKhzSg5Wo299CAr9dxayzf
q8grXQbZV1VwMAzJoRdHTZavqnRD5qWLK2fG9Y4m8BeRglGqaF5e7LRlSZvuKtIIZF2OIzt3vnNV
3K9P7SXeCa/8gGiZZ7QWslB1H7nMpJgAo+KH8DzweGHHapo3/mPle26cbF6QTaY930rZMS7Ho5U7
4K9N2eUTDSnV44G/44gHcmZiH8v0KLqptf3NbmV37hoMcuccH4xD6kj4RxYzSs2igcTD5KdD6d3j
nVrKlleyi2NKY9bxaf5MxLNemLUz78uSfBZKD2RIpecoXojJWoL5CM5amPvuKv+AdoxFEhB7U1Yb
eT9dIviIBMjZqVHc8QdA2nofgSKza/YY6H33pZfzMIwt/1JWUlsEyZsmY0NqaWHHg+ojxpV8aOvg
uCcvKQaRfIRjOnDN0cl7xFRypM15IPcE/julGSytr3WxYhFo89oJfe3bW9uxe/p3mW74QXrsmaCd
ybZT4eCmMrURCnCCeEijnZ43zLervkX2jjUCltthCph3+hQ0uOJHsQ35kHYYVg+5X5JGYoo7w6yL
Omx1FQqHa+4ddIf9R7crPS2HnaPR1haO1ckwPaCSox6ALNvMXvaJab5cYBqrDPimA9L0mG8DTNPw
Lwv3TNVJXRn2sT22YwtPG6i1wk3+QCBUoSLneXEMY5wGgThvU00AIPspQcMRqPZrkjlSjuHfliew
AEPO70cVFUEEojz0C1ywHyIlvFyI6d19mVZdRg+jZKWb9oqq7QQf7SQT3tgNvoSuIYIZbRrjAh+i
WNmP5PJVFzdVQuilMVIkdQnr3ZwhSwyTHcWbnGHx5jC6P2K6WTgu+hDDulykrpjdH5u+VoiW3lvg
7+YwP8XIUZE/xk8XMhHjG4e9Z4pRnnHruVUnEz08P1tiF/wzBP55MMfPMR9J3iaByfrO77X28OM5
jJX/p3TiBA1tDkLEUrmDPSELvxcqILvvS8cwFribn5P3tDrI3ZkTA9btRDIwKOrFQQVn+ZwElE0/
C3NlZW2OyWwf4xnw6mwsDXtdQl1Iy6C34dPViX5FllQvzXglvT+tPNITXlaWH9+QQ6YAlzkLxnMV
mwD2g2ir02YPi6Gykq0Lqun8sLZFZhpr5VPvm8xsK45/DG4yQob+P+fjYPMhVkPhyOvjNz3A7adL
ZyHoS6vgOPv3nRX7PnphXMpXPIrPCLsZKuj4Ewq9t+eNbeK64FszuzONeDFMqiwEHL+dyQJEQ/FS
bT/Q0BkEK16KMF5PolDI6znUPDzVQcLkFVN2azGUn+keo1PIS218gTCCBPyDwhw158l9L9lppqKH
sGAExUslO75D3qzJMFwLmPeIZrDwy7sITwqgvtYZLxt5wJjMlzTHb7Taz8DHWravkNqHw+HzVybI
UPCb8+BM7EWaxwrtAyklYhbZDsmhp4KL6WYU2O4DDWsp0V6CvzEUPbjFGJ7tRljCdtE9jAisgnx1
aRsQAbfg30wmISmpomoX1j2PqQKyYA3XPHNGiOlQT/vfCI2xnh8CGIT2ZOrsBBkyrCr4rjMGqj0N
t2XBrK3Do4Qlnxd93BF71tiTFXFBH2KHr54mnpCUoAEXmzqQMqFNvGJng+3DoSo8afznaSBYeI1E
09sNHwT3+/7VBOJuxavzVURiJbw8SGJ3MH5QEl5HBtrFxANqOcyvomkRzzavpv6lEyulCoG3hbXx
m6FydDp73bgTMd9cFsNvxQx6nUOF0/bbW9bMK9eh7tdv688zKA/Xzr+LUoJnyAVcc+I2agw9CxZ3
R6aQKaFrotpd/6sQ0DphpDOujohYDKaxyBefU2g9gQ2Peo5VnJgoKEL0fuo/7VvRX7h8/TZXGlra
/eTU3keYx7Kl794wGWt3VJftTYOYWL4VYpl70BW3UD+b/NgMPH+h5U/nX4W7xxRDZtvsWE3+Gw67
72+Y2mdpPzSqVRLLepx8hQm1lgaA3cqlwCgOE0cWC1ri9MV28srK3LpssLiWsbuH7okS8T1OClTT
BZSg7eKZBlVl4AEmiF+4/mRBTc/mQxHS1asbOEjK1ogsgWpYZ0rO9VgVo+/Dwm6+5dXoc8SuV+HF
96Wg0vW/BP4T14nqHwDSHkiyp3wM7NcJadBtT4tqkMqZgSQVOReHBq6VZ7s67vos47ZAVnBlCgn6
kJ91vlPn9ozYJMKuq3vt3flYXdNmFZwcKQl8kCybsF8PLQoXZPyOeplG/GmOjrpo2kGUMDBUcqNA
8rMH3q4AZMlY2PkMpdAPtNERAD9asPOPdmVPMgA9rmPqPpXDQn7BNza9eBtsYZs5IwvGOVKg1YmJ
4KDjjHU2VuCsEY/kbyNdT6melTEQkHZaWnRPfVi+GnVBd8LUH7AnZJWeA9ElcPjSBtr8g4gZQdIE
XvgXTnNYpPIuu41cRsaumdqMrwvpMNxyI2/qO8c/dxEwJ3xi5914Zt37/eAsaTLhzqMEobMvRoMn
fjVLalIrf0v1Uc32fe+dwz8GiEwWlczLEy/vW9TA9LKv+Zs1RC09txUaeEKSqtmhhcr3hXVohCoA
JDtqd38J/T5iW7pUtfSdOWtOz25j5E2l7Yyn0qKplTj4hs7iROP563x7rkFgBfZPbXA2nTj7ZXZk
cbvGXVbcSoyOcTrxRrCKdJd07NPEI0dpQ3Fw2VNh3u8nm0PCr9Ly3HNZNNQCg5o1oXWOPUg3xmvX
Bb0ahE/PYpCgHffsxUTuwv2DMj6GnExdpjDkMBktOvd6ZltyYSxv5x1ZxhGD0N/SufRLn16QjS8v
5mrLBBPZ3fgjwF4Ve6MOF23oNbCpiHmFSAKmT+zwH+IvcefxSzhVQhSw11OLg9mjOz4qQjY6rvKE
c7kgkyD8Mi2OV7h6ZaqNRXgylBfJacBwV9wz9lhw0HwCJ7/QKxXqTWlu8qYyxpylbjpkMmJbTI1J
quYHY3s71M87gUyO/mFcDLrklgd6swpFNf0F+7fXn1KWysiBCXjjUKK2LLlXaJiQZMD09YGPZQoB
0uvHYJaFFjVSYQosHF23LzxE1E2+i3eM1vIL6GyCLazgI4nuymyGHiN2HdXvm68yoO+2x16NxlZq
ZWoxUWGDdlPiJi7cPMKrCBMOjiRtDOXPYE5N7KjG1K0L0YrbQ4fbc/ZbFlnsTBohyfQb7p1nwOyq
omhB1NVpY7uHkj7Hy1g9ZKXwJMc7tUk+yL58g+9bC6Dw5r+79c+4oGS6bYitVZt5i77n/EmPzY3p
d+bKo2KhN/cz+QEB/cGcKt/CSKHhnlSdWg8r8fAYJqgtxE9Vscy17DFlB5dz5MXZ/cAXhgrILFBS
wRYIKn0yuS7z183IfMT7IbXuGS9QhwUMa+TL5gWYdWoeUd25BMY0n5PPi00zxugPOhw+turxOBBS
h53mHULoAtKJF96e5bYVFW1CpumxBMba4QjGHQeboUsq5azeTNgM9s+kET2nU20hqvLCUThrrM7L
fhskGgXMrYmlhXm7RA5g2dhkuP8DU67AIxgDy1btexVGLWY8OcO1QJaF3+EBK42Z8KWbgob3ypn9
1567MN2M6Sdgi3Ml5q2i36bmsRzDjER/jjnpbESTx8iJv61cYEWMPGFC3fwi1WnXyoYk9PJlz8TM
DTeQ7thukGR7E7yDBDJBuCo/Uc+rAYz0LE4kyHHgrXI20BzhD8n7fhfzkw1qGXW3YAZyMrDe8iGS
zV10Aeu0zfObQHMj1GCV6nH0dmDrgNDelCrKrIDz8OWp2RF65ktj3BbwWEXo9WfPRm+x4ryRc1Jt
oNOWB7KaIln2SyrVkcM9pyGVgHf8JcDRiXgIAbIJPQKtwQKosZVYo8kv8EU+mjk6kO8o+7jbrA82
tlpLn1i7PJI9MgKhJEWYiiL5VUgvY1+2+gptYmuwAl+czNjFKYAnjywAHSUs9D3ZcpytryD4A5v+
2kZEL9EHEuAUiZLZoojInzWpJz9K6ZvpZIoeoVg2vf3DMSrHBqW3+xfweKioED3lBd2Fry1H3DW8
SqQB8QRVQe2Xh8Zb1W3xxsmPC7m0i+pBt1sga9sPrqYpbxy7Nn0sC3TZqqBYAvHxdVaNFn9TrtkU
Ta+BWxoWu5rj/hM9+k7bXF9TmhOvpV2fYFjWNz9DrPmZ5sXQL7lwxz9wJCxln6kuKz6dzqGVKgPZ
2Kg3uB+PkzedsF/wE2OPFYurvrQIGMyqrjTuyROg3fynvpaAA88S8UWuUPQeU5vBtH7Ip6j+5Nrw
nomnp82LizYxbXwGv3vE4e/wDx7EjX8tIDAaWI6ayJmAlypRyVse1p3boWVZmYfe9TAq9q6qxnbP
qI3KWJkzBsL3WLQBLDnMv2ZBYRG+6R60jjTTamYkoW6+H94v9fOms0+Zgb7ZDn/HRpRTYdzgew6W
VvFweFS39khiSGZuf3p2NKsi7VDXrMTT270Z4wxe0/cCHWlzmVzpBbpnLHAP9IvtX8873QWdWc6E
NSS33nm2JD9OxwPiwgD61cZBu5WsCEkbEcke3vWp9jwdlo9cNf1l74BkO7L9tmlx0huCEbwMDts7
oCOi+KEUo2CzC1lEMoadstsd/ElELhNwgVUGv0k/MT7bZXd98toSbcJQThfr9Yd8RhZYgstJeHqh
r+Y038WAcmraiw+siZIntqQH/MZkZgx/xobpdCCmx4xjlkYevK2zHs2JRDbSX6P8ARYIVWNR4jkE
WId7ahXDNixJWpYlZfKCdJEmXZUhpd33jdAoEvLfMBnX4tUdMHdW2Tk1XpgHm9dFHYsDxNX4/Tzk
0WVI0XzhoA+n+hRc7CMC7/OmcojKiOtFTc5OCjEuFKif6Coc5/jK0nB27y8QE6cdNUroEtwvM1os
HIsYkXaFSLPHCjeOGP57oNEwm45sX9ZrN8iu+mhpZQrNsE/sTRt37f/1DdAzMiWtOuN+lwVNTmyd
0V9Qrwo9KGjBKo4dcu+S3wJrC5UBKvsXQCXhKj5N3QfLiGkoKRdT7Vymq/umxvQ0BIbCAEgbjSs/
uONuU60T9RC410c5dBGDQxU0DGgZxj89cAPENQuwnNczgzgswWDWAysyjwOtlywcvv4U5l7nxM3C
CicwIxRIrcm0Vp5RSLu2SMWTNKQOe9I+nEJfh/F9Mtf83HDN4f5B8yWUy85PKlqwFpjS9Nrdsos3
zfBOtGCJjEqkSBdkQNizIiR7KnTpAGBWcPG1nHGQ6nYz/cb5VCOLUO8uRyO9+ljVCAcLJp2mEj2Q
9U+L94H7tExnwj0S82tLqnlVjGwQKNpC4hJDhi5EofHjEWABC5dLJnpMuHUW7z34kt4nGkoVmMlD
9YymW1vMTIRUU2JAdlo/5MoqA6MSSAnI70Uo1zQVf/3yk1wXFXfz5ATOiZNyJYwyP2o/lV0Fkm4a
s8hZpMB9W0sJaqafEwAUsK2rmfoTWiOU3Yxq42LOvqqJi/7EfLMcYaoLWdewPbEgnVXp1klow2xy
QWCdbcouFy4fJWUWoDzcJsQKL6kDyibopqZbk4ieODo65OeNIbcAwAwngrSEGyvTvxmwkG4LaDaq
87HF+Lwuj8hi87dHppFyvK6bJXcrOTxBgU8SCl52BsNjHpk5s2ew5aZGUn3XxekhcsoSyiypvG/r
UuMjpYxHmS+lkG2evsc2A6JkjbdcmmMwZdHMXF+WtJIyClr4ICASPzVOzT2qKPAy91DM4sum1G8x
PiEc/OW8Et4f9MeS9p4oHbZA1NaiSfDXYMY3vuM6ZtoCWz9FBE5iSXgQg+rmw5eG/xrwmkgnhRF3
9SCG7dVx1JVtyrGdOreJpXZ9TbWlArRf/focUoba9H+NQgY5BBl2MmOcM2QWVjQl32YZ5dKiQOX9
YTvANdaV+cxZbMtcjYZstJSbHDglZGEVYZzsIRMA/yfQZf6S1EN9wdMkJCTzT/bKbHZIEuP0kzAO
LGoc+qfvG4UnD65e3mBbp4bhpeor+lqROT/YxUxvtkHiBtUZ7w/PCgWRZWbb6eSogOvAFhJRkxGg
BGsXKxUzwEu6+BnrXgvG9NCA68FuP2oNjFxIiwM2uMSRbCTtbbGNsfXCPCLTlfhHFrCubQge6oQz
TU0yQHbYZfLyXj/Q/GlsT1ybQNW8j3vWIfPk8AXqwUWffNA1oUgBtMR882xQCNH5KO/jtHfKUol9
HkO1ltxk75qjSYG2icNjBwS7JUt5mwPzGQU7tj1swWUl4KJ5MFuAyjPvDuiRqMGUpKi+OW04/5qZ
WGoZsnXX0YVFUU7r5ya5zak5ahlrlhD1nQrULvg4nVJbUaJb9lZyosFmCSe3EjyDnZRKP2vG4eK9
DaH81qmZFkJqT0QNT8rO1AyUPiBpWgQzPC8qfpR9+PX2ZT+RHNERjkNHiNJgHzMlBG9hQWqeeICS
FHCAnO7HWxy4OjAdsPBUuOGfLqMwwX1yEl/Eue0q4g4Rer4aFpzQHgofIy9+lAam+yltVC5Q5o7o
1Yq2TiKUo7vjfRL5h42I5GcyXHUgzNZYlruW+u2SCZ7j+5BhujHF19zvjmYOn4DhY36BmG09dESB
/4r8n8KKzrnBs2ssQwenc06zOAMJt0Ro7vRfvfxM2/121/EqVZWt23IpXcYeyVw/GL1I63d6i7fF
tuMDrSgYeyVMuSdSMEQDa/moOGk7AvWWC21c4lZ5OmaW1lA6kjvyyjA3ByLJydeTchgO0xwEbwAV
qzYgVKLdluW/NqMr+RnHW62OFoqZ8pFaTRKeJ6EhHVCexuNQZGctdUbt5Cln8v4yPJK5KdSd46Ye
V5q8B9EWhViZ064s5UNJDvdWui9udxLEUCSrAFBq7yMHZ8BGD4PRjT4WAPq6bQ8cacoElY0dOBq2
1Ribt3urrymGgZy1pAmeJ8hnI857dAE42nVVHTYo0qhyWSNVY8NZhuzVADGHhgAZ+DX7Ta2Oif9j
LDKJmltQ77uedHpEwIFNYo0JC0ktGYmzYYO/uBbjVcZIaUOapLxG/x6BK5ms7XpqNLQqumf0lA8E
zixBQXDTnw0eXCOtxnvrqn6R1ZcoQZYjyku+EkSj3tTyJ5lGSBXNDfzydYWD0CI8xgbUZazdXpJx
TTkwDir+dCQ16r50o/2I/byopX8Ei2AG7yDtyWJ1Ek3yBwNuGWRs8izx189T25nUW7I8qTOrRX/i
J8tOUUWK8sS8jH5WWb/BPwe1gWIctyl9i/QxOwQmvvoczuPjQv9MLUTUs5m48PJyAPkCQRKY8nC4
/jMdMu4Naj+FOcQaJF6lc7uNWvDyUb1UxTXUP4ClZ/gGuqyk69mVX4hzNkhv+a2GVctzOeD5HoVp
7wKEZm4knbTN3Cyqkow+FHE11Bn8FgJkWtt9HMLJFQE5FAcbaim4VVWQC0MGFIMUh0MYxB1fgmCB
ZO5npc+vKr1S27+tKT3AIjycaBS8zQ0prh2ZXm3dvF55HIN6vLYTq/q1IXmS9Dkwgv3uG1RGA6ck
ut9BjHPsR7o8kpnRe2/csIzeezYL4BBSJT2wx6iLX0bS3KrIrA7WK0WlN3SsbH1PPZKPChmRPcS7
bXiDSYowo0pbYLlmBSIWQ9ylidVoZ0vfYgi8sIxvC5PsdMADrqs2GDLompDqz4ZEiU2ZK3CTJ0JV
tJnM9NXaQSgnQ6rEluvbe/2JO2RYMUK3O5KrXTvUGkSpYOkzIg3MMZrbzq3mRjrb+wuaqA3TsAZW
S9yW3UxQQndXOVh8yyA9wXotQk9QVDxszpiElNRt2jCOM7263wv1XNiQPsBoBn0tLBQP1b51xCyq
NDBqUn9qpnxuJ4Qe61JvzaAB1ehh6Im3a/NQofo921CYNzlAoWO/zkMlNNdeteNIi8mCsJ+35fxj
yl6bOBfcXP7/sHtPDVJar1HdTz8cgwbEtP6epvmpqpRrxA1y9USL9QohnajnY1pWnH5TslE2/QwX
Dmm4HAPJD6OrGDeUV+iv6Coy5bwsEak+9v1X91cgvOudB5/p7UuuylfraGUalgmAcNwrBr6jTC/D
hPEbyKPyopKR/UPyOvNniBdQCTXMd1ON52+AXqIl1Jkx8Y3o9UnvPSua/HgMGm8D9cWsFCQgemWN
htlc5iAiChCMIWpAvbZkLDo/5NJYurocF9Io/buBVWQkRZzjoM4vz32LrZQoP0Gny2yJU3Y+qmcr
Ye1uPp7mXy9rh6gWZ4j3FV+w7T5lFEHvbIfEWQe4/CmnqVpKF2gWM/njgQE7NNzdRRMAnxL0eT1K
Fs9zMe6L1XwYSvDrtGdsIO2t1GtxOlUp4GLB60qJrURtvFnLw5/yUCiQg1gYgiwr+GXzC4s5Q7NE
AkeKOZ3Br2mUX8/nkZzMDa0f3mtdV6P0fOb9QRjcTcDkQ5AjuOIewm+RFUi1jMjCDUQkLYyb6GAO
j+tCyxy2d9YB9gea/P1b0H22W2yXyXFRSO802XnYaDNHYyBaAlMM/lsY97DuIGDvXMLZKo10/ZD5
LMsgg5fZ9bl8HsGpfj5Jqtly//oUZUj1d3KCIncsu3hJg9rKS9HMRD8W/+KCd++a8qzwdMGWlzfU
dhFdvPSexs72DuLUlXDmUnlvy6mvzsJTuK5r5A5np0MN/+S6oU1TzHOzXz0x/2N5N8V4SlDRL7r2
OC4ctm9BrFDkv/j+iZCk1MhGnl5PiOs7bnz8RhFfCM4ky64SlI9i+Oh+kCEFTs1UvAAmss3D2VOy
iW9n8GnkZjrYRrU8EFA/AVmMgCcrtbLkOIRcl0dE0WE8ZWDeEYXdl5h+0FLxmtOA+fvgm4gH13Iz
KAzQmws04D6YYwwl1xEDfyq8QSLQ1WE9rUQ5YD1eNk+U1h9vpDPJjEbsbmF1Jbg/gN+9inOofoiE
+dQCH7kp5a35C5vlWmd+Cy446yuG8n59UMhgFQAH2283B8/nuirAfqyJHjNZktbnyRX5glKMCtDe
QwRD2lhDNT8tJ8pRKdIXB1Kra0R04YKauEarZ87b+rGWpWE3LMYW/NI/TNhiU6bsCqPTs//dy+Sk
6SQdtuBvOi6cfL5i82hAxbCgciCA/VpcQqvjGdIfWBaCOp+x74Nev1q0cRKdOWtGO6aZjSHZVn8n
8etRMhrIwd36ctIhwZKGx0oO8/mY95Pt11KlbDKtaeIyKtIgxW7SP34HtDKqxtp50awTeEb5QI5J
4zv4o7MPje9WRL6x6G9Zev2xsIEccmyPYhYGzcE2Iyg16Lfm+AwlK8ebYnqNKyM5Ss4M+zzO0iqR
gTF7DG7XhZONESypMnBRCMAd3Jft0zMYgTxAZcevCXH83lQky2EFaLu/lSPyCzlcYL7c+DruucoD
D7UsObMargxFrKOsyhTNCqWzac4dLB8ZE5PuYNm6aO6r0AXr1jqvi3ZrvbNRqYjEjFBjXUFdyH3r
e/MdB5B/jfgQ1LWyA/kiKnGxd4Bp0uGRNtiGwbptVueJpPJAIcr+uFxPU/tkO2FSbYDa8fMDO+TM
gGubZhrv+t6ULBZdJ5XbWvXBVNjukL23xJHV7eE22s+VX8VAte5esj30N2hyKldZxn2GRLh4FNvz
j5s0cXKZZBJTf7DczF71OaC+8/Y6m1y7CP4SGYmB/facTEp3HxGtkAqgHrMW+HaBWdzvJDH5IjTw
rQAU9Ih49gcQWXiHLKtB9tS8Za1EPjVq7GpSGUJG+SrviEkla2aYv6QS5RvrRrxFGVInDLWB9pcH
Nle9QlKI7XZHVWE67vN2w2iHw++UibFUv220v5dJKCF0XEQ8KbZq/1QvJoeWozETKXHvQvBEleXG
my9tQqbLj8BDuBf1H3kh885uAHsiNe7LN+YfGRUFLdNAtTzfZ/DcgiLqeLUeTDthVVuKc5BzHhTv
NI1nbyXtbpLLROgqmJt79CgBKfRE9IJHHyo9rBBl2ABApDLIWws7gOZ8NMd4IpN2zX2UG40DyryA
C62ACY1wERY31m66Fk5Rw04F6avXLMloYaoKmOlKeOER5Gdj3/LGoGdWiDhw/0/ltCqBtgnAU/8J
6Ak73jTKEZ96/3WeRtZLTA0qa35tzrxmT7NR9dHfX6t9Xlz0Zu2gE240W+8phoKxxfglrP8+Mq4h
F2DOgkkyeVkGpLO4xve9ukFIOqykitoiqUTzyuguOm54tZvh4k6gpOxsQRfX975DyN1r0xKi7L/S
I1u/z/CU9e+qOVnm88tVz+gnE5+avzyoNJcC8nLIB1QJOBZhqeWJYDT3xUKnwx6zUpjG3X/gplq9
i46A1TyhNYhS+rv5QJxLk41iiETsdME49s27dvZgbPZN3/CgAMQQOVvA9TPd9posRklesOxpE6E9
sURz/+jkv+2OUZJG0QNb9JMR22dy1DxEgNUFMU7/shiPayqBqbAD69EIMeWduQFauQoBDh3zf8FY
fpaoiKmK/49PVPl7wwYFlKNlju0J573TptnmGJSrFQ9/Wyl+a4WunGmuy8G8PUPANGMmPGwjw7H+
nu90CP3Jz9EsHxNMhMXRL892xWNevhkN7G9wuc3ZOjSF6FPRHJigjMxexLJb2Hd7HnAY8oB4NKpA
YPdcZnCcMs7SSsL6dvkHrlevnvyfxV3PGUDNZ0W/Ekm/kHCbJjD/uxHMxtpXt2YmvQY/anLI6HC7
Sn6/J2tQTwebuQT/+tvf1lqgiOHcfPeAHc1m6/SLgVxATqgrpWkHaB/SYDyMjimmEvl/xCqpDrOB
I4vTdh/P7yc9uB/4qvMRPhSB1XDfz8y+2rplzZf2w3do9z7f+1TzJ8T0x1WF61tZxgN3XmFsYKA4
/V1/7Y2s2Ls37pZOIvkf48bY3XYRDtWc3G5qiY4YlLSfXlJpbEZHXJ8ChFEAkNU0f5xz/LMEl6By
9P6jF5/BscKVR3F/MCpBzITrZcWlKFKjoXedvwhpJtrg3cbdZU+Vi1pM9t7X6SYoJyhodH/50Jxs
0ZqZY97GW6IsyGOGqT/hvlWxFNVT61hC0rJD3wTcUF9ZroZfEbiBNw+eKBi3Zgo1wkbRRv/AEo6h
lQak9MrqgYpkQhiu5at7QvXXbc6JBUnSxJaUAiBVy11l8P0iYssYUKBD2DffuxCfJVnVgQlcJjn8
PtnnZKSa7llLcSssZ8BfHTeqJDPNunxLzjBwwlRWS8ZSjSd0rroSkxmRRSEjmLKxmUzAVV0RsnCV
Ei+M+d0ZkqAmlT4nhtlMsLFVJB3cKY38J8/cYxVEGMyaX0j4jmKqKbQtfIGYXWJ91EqxKFSRo/k0
Jz9YP0eux6Etu0dzbMBKlEYI7tW3MtgrzGiyIqWXVK4H8jxaYV2PE1tk+rr+ktmwhlOV9L8xqVyu
Yrja0TWDy+YRiCPUBV9dKciqaVlg3L9MLG/EwueWJVdYSZs1UENfUR4/diLgqac+qnpgHozqpsHz
3n21nWG/ZhwHPtJ6AYoGF556HmRnlMDaYWTPLJpDVoXRKjWvbCxpbw7AIcPg3Hstb9cxK+P83Up7
ytIOxjCpY4QKLgpbCn4dxpBKm/VwXlLdEG6F57yml5LomMnNQc1gZYwhRJbUV+zN7R1M1D1Np7yl
19NqctihTtlCongxqMfbXDwsW2URGHCWFx3/vFxLonj8HTexA/mDCvopad2/bc4ndG52Eqg42780
HZJeoP5JyxGscNBQjzr9XjjkPt8ZK8ghwCUEl/WftJWLCNX8J0Sj5kQdjyTLa5vAhttPzvYvJbiq
SA7oKpwfJRnVMBTdDYpecN3B/cTWwYEF7BakEyZfKDjI3kKag4qVdVtL22gYw5Zbhx7S/uOnACmI
btaveno339+HweGJNajXWILUe/wwkIazjXOLKNVi/RBKZWPUz1FMnI+MBmnu8gxfOkRB9naUn+BO
bJxedwdr53nuB9oK/jp+m4ur7H1qnkpoWpqVb+qV7gAJk8y9XhqDG7JzCNY7MH9R5KsoxAyQ0tKG
GFnPCOEAf7FVSvIFl9Pl8N3SO8r0Kxr6mBYeLJpYlc3UJngbNllv2FvNM6//Epq8Pge5zxPQjK4g
ADWHDVayHsnpbXzROURqF98/XKQALIYE+1QQLGemZ1MJrjvs5spsWCLaPeWDQZ7Dacz/l7eoUzSP
uE8IGF2swmcsiaHLOFolF6dvvZqdp+Pm6phcp2en8YRAdOOEGcQB844I51nn0xggAVftigl0sEtP
p1JSuto4+oVJKUuiT662sb6Q5m1aMLbjAlse+KQd7duTPflQxDQ4gAf/rV63CWBY8zKuU2oAnJzs
QrpxLWYnEHVnWxt43zOemVXHFjHzK+Ppy+Mw6xk5PFEvMMlxr5tNaEiOQkRGAwBPhNJjLLJ3VjPt
MTcbRKM0BxvCms3FS87HAxOV+lVTSzhNjaiytiUgFbPhnsuxV+FMUNsl+8XOMP73f490J3uPUOy7
i7HCOK5DDoss5sV32u4L5nXjLWZeEC5hTlHUBaxR+siDZF2SwBNb8Mm7uVtsPVXh8PwOkO6qtY1k
bE+00xPLM7/4Rf2BvBNcDPD5RyvxZfcQjagzEajArL6dx9fOEvC5NDNI5mW7tRS2lI+LPspfG9Rz
x5dRkC2kKGqWH7Zs9JMa9pfVBXB1UltwSFaFFKhnocOwJkwN+FNSklzj/UML1zRpLwQLItA/ID2H
ehDxSsn6yc375y5AN+3sSMeE42I5eUM9qkPshd5xatGQZaanOol50kp2dBzwuYyACd6+pFfWb/d5
5lrfDBKjhgeMMb93HiGbEx1vMLscgvcOupKtUvqJ3TTDVyLNb+SSo4lV6iRtKirgW9Adwc9GfiF/
VKZ2/tdZtbfxXEr+K6SCJwXnVl11lOfFUZJiU6w7vbydz8mnyIxKlGUTjGdM1Zt9Po/kww9NOgQC
jFfgrcZDgbIZ90Te+53hBb+ikw7ijoSE25sBOkugcYcKiDHha+vLlFcWmtIQmvXcCI/C864geIRw
TxJzdI+F+qNX6i7jligGYFSU7rlYJ8GwUl2LCGTgRQiQRsG0MKkgBTAlwW4AYJCdg+CrS0Td1qzq
+7oIhkcbQ5XBGmRTTXQW5V2/XxGvXzR2rDVUOlAP5ukKVHD+IuwkH8X58jKK97ESIOTIuRxBbCwE
Ku8UgzK41Tfnr0edz9rEelrCtYA4QwBPI9F2mT+GktI/gNIi5VGOkDOa98lEIVZB9zMxrko5aGTZ
bS6BxexKIqe6SZlW/o36G2TEfoIAm3XKHjSUmgMcMigV4ZB4axsKPLKPQJVZc0XAb26NXxkr4r6H
X3zQChLxRALNvAkf3rZw4SmEuostNcG6lBu2b4iHIy0pP5FdkvonxVmxGKq8EDipQqaOpQjwRRrU
j4vZwKIxL3nMzWXmFBZlP1TE52+RWBDG0NBux6P+Fv3NdQyG4CjpwHlwaadp2l8PE1S1akAxO7vV
D2sw6e3B8W5xu37XRPmO5ZA8oZ8ot3s1+3NUrSyQ8OVSsf00QESoF3Ykj33y5wi4/rDY0ddHD+ES
fXbDERuSGGF7FqNb1ZYjpin3ZnA20qysqjUju7IzQ1Lyz2fsTxSTGLtYrrsckyx+ePar7/O7hclx
mS53bwT8K7/Ajnm6JwbrY++bppqBnkV+VYj+42CT44RgAscAbR1Ko2Tqm1aQonaI0qdtLEus4G/o
ylKD0qniItSHLur7EQPn/JiCKAJ/5XkN/7z5FHIPmBPWu4hd2O1SaKH5iZrvn1nwTMGVznzGHP0j
J7jCeeExZmqNeuoZ82yxUHswKyqsLjaf/wf1E4tCYz2VU/c6bYZLBSb03TffjkqETqZwL6u5YOBO
9FnzuxA1vQzAmfSF+e94cE+FIR49jYPZ3977AdPdifUjtWHdgd60yHXFLd8fciA9oAFmv8kbyNHs
Rmx1DgjK0Dqo8YK0f0g0xt2VFhdSHYi/A/DexL0PSCAKSEXkgOJ2Lkj/AjLm3CshHTBn3I5wa/hv
M52yi73EDUhfnaVCt0PAuSchv0X++HQf8BLg9+WWXCBjVh3r7uhwHAsMsqP2ehzea8nU4Rm58g6U
TjDlSGBTLziXOo0Uid3Sf19Nt+17tlurCHPJOwJzED2h88QyQcTZKMd8zFV2BbQYzb8rU9X/Ng8B
YSvPausYh6I/Gis8PwYXScANUbjpCUZgiALGHPH8R8Fyfd5xArPDKL3QKK33JU/nV3FIt1vFPM+y
LBC1MpDyYlT1mDsFlHPKCbRY/mEPgXVFvHHvwVCROFBcm3qgxIdaz8J21d9qmGu5xNcMcYIsNTeF
XKqXA7W0vAfblSxJnK90Ar36kS9OPfxhvRTWo35BKEuzefINAOmbkQ+/G0cVVPTu1H0CCT5z9HD2
Z8qM4iASw7JnYBhrRn1Ej1CllW/XrN1J+1Z3ONRk6PoOGV/E4slP7UroVR2hOqSNw1gbhAdtI9Vp
XrQ0P068sm6FFPXJ1kdRBSLBwIWByb2mDUsyid7ii2uKe6VGjeC5n/lOcpybDxMBIfhHg3Ioui9d
Xiv3l03SpHVprKRyQkC0PmuXCntELu/F/1TsWdwmVm0dD7ZAe5QdFFVKqK1pGPT8ZNEz0WxGTmZU
EesLLDjm9p3KLUGyPKMU/6YTDM+2P5kt0wT5qrv/Ue8t53EzwtYdrnEUXkPJsie+1F7z4POt047V
NCSfFA1pFhUy51yUqQjGcNAmR7PQJuXHdst+LRbHub0rOz1xeRUzZsdAETOmEoj2FCFH6aMe89WR
ueT9ZBlI1M3ZpMHu6BIn5BglF+OhVdiGsfnw+Fya47gWSRlc181zlSQHR1M5TfTajYrhOfWvGtgx
g1tQ/rEj+GKBXo/oKODt/b/9zlAIpIsJgyufUHo2pwWkCQaa7ew5KPzQ0UKprJfn73TwHZrzR8O/
uEvvhRWkLUZ2qZfvmKOhy4tKGIxUezZAppa1yhNheByatJwvkpHzAb2w5u3byipQHT6c2EPKSBjH
olivAgb3JcEuu/e3scBrSoJCm7SEiymCNRjNUGpz/vqS/sU2SMssTmD+cuVdpuDv7DqS12VwnT5m
Y8l1lvF0wSfjRz957aCh/afe6hC9d5nmNdCwQrmHGhLo/icHj+B3m7Kih+p/cnakcArM+NsZJeBr
KUHgeYc0O7QDY78Bvnvkz8cFMg+FLvlQ+KSyTpu6h8v8wKmUCt4izqBeA+jYMPL8vSj3xuO5+DXQ
vlvM17OtNjXryNQ61p4ruziBLWm3zFsLqEJRCJcEvtu1BYWeg4bie04vb5kvxbAdJMjq8qKnLZMT
a6sSzM7c6/B+n3QHAGwBl3DqARvsAIebz7RdsjoSTwtBFWOdyuaCPJir2Ylgs7ICJs9RkU4RiKYA
sriOm7HYbnBtavs2gQaVA3dYltSN2O2DGXwPaw0wUY15pp8z2zOB1q045125NtDzAJdpia+BC+8W
Ut0DxkoGXoDIdOASWxj+RYY4gB+JMCLMshWIOaER+HuZfYMHYd9+lChx+5gLRuhkqAyg7yQtjFk6
f8rswNJzjThiw9nh1dPhHElpUXqt9qGs/MICdWVNAg45+bAZyncc/XViSxiUw/x8ULp6ybrsVUmL
1/coh6ejdRX/9JvU1eBpGwMoKsFJF2Mj9AF8lNkRvukkVkZUzguE7a1I/VuiruuDpEAkeZub07W+
DuorfmXZbRgjui40MksBJGwgvPfryJ8c3qpp3CfAw61DUvoGeD3MhTbIiRFGKg7n+ZAsTYMxmOXx
PnuI+fizixqeBvRhjYO6B7FZDePi3eQzjga4jKuJoEg4d9VT443GpVOmKsBAomz8vXrKMqEbcmvE
CQ+kRTzjtdDpQBpkPRzCFUpneBIR/jXEmx+LT4fuse3gBtqaRj1avFOyIGPaL92ds/4MujiTETWP
vliwpAPfN5DgAPSG9UMjkEtqA1a/UgFkoV+phsMLDHzx4Z34Iy/iSfKh9/Y7UJAP7nKQctHbjDzy
CdfHey0oDZeMY47z14Fkf6/4oYwWCkLCL/fcJtExzHKgQ3Cf8mjVsnCHGKINoMptjJWVN+VaC/0Q
jNDZZ9l2xrrl/jrRejzAi2BMnSMz1ixwnjcQWjykkowHeyBYQvYRrmZIZG03ZE/z/V0IB0gaPxvv
jsyAlBXvJLDKtcG1XLYc2G6905zd5YuNkF+63WyLJHme+ATczXX9LKfEB8FxkLW/XstdJDMwKIIN
4ZyDzsGK73skgUH37z5f8yreyZkGmWDWSaAwY/nbSyWzijcu4ntYxmGhhL8EUh+JUzKQdhoQH+j3
gi1ghTV0OuMIddpkpJosK+7Gflo97TwV2NUGD//x91+YAgexbwl8A/Wa4x117fWofHpokApoduv2
+MgASXmlFaEUyURAXwlpGJ83wzRKABi/Y9j2MD1V1nmUyzSpwHGybF/orn18e0YEB/TqStUIpmMo
5jLZ4MW41osPfVTMV8iXtKxapzzZ6aKxyvg3K5IkU2fCtDhCJ4HQIMeyfq+1HHi2dQHO0i2ABPOY
OVWS34kZlU+nNwx7TUcpNPOjTPdPs6fK7d910jnQ+JEoHrTlj0GZpFOQycj2dSazPd6BOhEtuTaj
3Y12ZD6sxlCGne5kEAUJH8YSnLk7H72RZVZPT14VGtAap2o6rQ9xBq/RpbHQ0t6AyHP9cp5SIPBx
MgJDezQmuSJsbWboFmKMp1ru1Z1WFHiuQowb1XFpPKY0wUENnwuhuyL5LxMvQWB2tt7mNOXDbMQ3
B0oaa/af5YMtTqPcnyGVUdNjg/qFS1KPaE62Sk3Qd3qtNz6algFHKPdsHuhjnUqwx4DxEfT/+7bg
toSE/hbkDq5aw5sj1+7pRmKBiqCBKWA1rNzrYIz0GQQ9IrGELJPQzmSK+sjBOvZyYVxnKlIQ1rXq
G8akQGAj+yw7Fd5gFDax4FDY9OoE/Bo09eXVnqFRlN0kYq8HJXvyqTMazvHTW5Uqs3BI7cK75I2Q
4HTZl25NEmDC7whJaMniUN4jmXrx+X3SalcjL/skkCdsWIeEujmbDWf1vLVCqrF0bZRWcZHHa1R+
g4ic9tsXlNkBY3Al1oNw8uoi8HjsILuWvqZV7twqdPjm928ltBU8rvwsEatIKaMYACfaIANJ1ZJb
f9QHCflQCy5GdkAtfQGY+93cCj8obXpQwyInm3+BQTSoPagkAsde+RDVjcpuysyxOFwLjbNkAABf
atwY/KSBQmYaYBBJFbXf4sUqLsKb4Fxd+L9gkh93Om+DesyVh8xTtmBqTgluyYDuQXmbUtaqzk2j
+7Xp4L+XEg4UgoglrKtGp/jzET7tIc26nTuh5uYX36vMDetU4Hpclx+xhRt2r+HplSz9Jjarvvgw
QY3nNj5lH5FGdACKs8HxQv5q5ZZRL7aC0Ym9kDIL5340MY64m26WEv1g3DSlZMbK+ZJ+uY2kPbe8
1RrI7Hvy0TqUtqZcybkGrfKQh6oJtRP+8cTXzQkBQIJvVUiH5Q1kbhQfFXd/FFfcftT7DydwYGS9
goimFo7tit0K92H272tMqVJsnBU3pzFrKS0eUcWtXwQLEyGusRtaFqoGx2ny+1qPqTuYXDxfqgH7
TUvAfgoQqBLzpqwv/A4M2BV+UDOS8xAZgpnTMKvSbt35jM8ZXG2C1Idt4S1gIptZcItpGstX8qLr
GWE+u6cZijA4C3fPDycJU096PAGazKyT14u5QCZJ/Vwr+FcaUq/s6IxVHWao9vGAw9s8pVB8RUji
nTdIi+nEf5iBw2tn92tl3j5URIwCTBgjEc5jP8Dnnd+We2VpDDPgElHUHGqZX00+FlrY2KSdMduV
esSGd/aNR6wm7/ZesLxoEw3a04bay17rdBjVRJgOV2VVqwCowi19BXJngvD88RmfslC6JFuDpbXJ
EFDSlfQGCQ6TQYLRRDNeMnouzynhHIaznJnmFSJpvWIV/j9T78gAZI+OIr7uVXTM2q4p/wD8rpn8
mO6Aqvb7PDDXr6+FzpdTU2EFIiZ8SvcooPZVDIgk1FYC+VKpIAmEDJFqBfUf1+sWI/eBX3fQizOd
wJF5p1gCw4iUKagS8uSgbcIKltsv3CTMwz1UVnAxHmrPJ9c++bwY6ymq09EfGKVMjqhxSKmgnxdf
y8YCCYPyCkOnA9lDZ5SprFuLmWuZVUxnRfQJt8G4PweoycoyIVG2zSOWF3pXrLFgUXOX5d+6Y6Mw
dBGxhxJ/wZ00Krxz8TvNm5obAABf56cTf+lhQy++l4J9D8HaQlC6JnizTjv5w2BkhN7r8g9U65ul
tg+HusLQtKoCdwA1KqpWc+fvlMKfI5iIgjT/GzPSzyETJNSTe8ALegPTnMQTN6XtzMmisbSAjKgF
xp3Gaq7naNtlRrz5AZQWQjbE/RtPn1lbBx1lNRRkBlvF1MfFN0f1t4NB5rc+76QNijnjF6t94NVT
Be8ryHOQVY8UVWwO0qPsWkHZy7Gk8QJ9m/lWPSxsBNd632emsD82slQGk3RqKXO1mbCfKY3vgd9l
uT7QvEP6cGn5Hin5++bU3IeacIZY4T9V8BvGGBEES9hrE25Kdnv2oqjpJE26MYNK7gXe28nU2vlN
L9gK5aSxaADFCDNO93WnsLHXrQMFpK69mHzcH6lXzfYWWm83nvQvtzsl0giL+cwe/nQxeed8Nsza
MIN17qBYO+RiGISkUdsaMoWjZ8NAHFmfih/lr8fWFdwFwwK2HJOdqKVcl0Elkai03A1DHyvplU0s
OD/+iMhwBLhgmwkWokeNTS6hZ4a7YvIqGJqUQBa46Mkkw1ufDoy95qzd8gpxqGLqgC1AhS8R+9P8
6lZENFlYu0jT3hb0GDJKet1pspNiyTnP3JRIls8wBOSrU98YRdWyASRy3W4Y/SiQAD5+P7NbhWgB
N59dOrJRDOsXq3Dv6xsbDa28Jq+Iyex7P2R02Vj0PPmxJ2mB0sNDE3ivUB56taZ/6yUX5Vaj6LwJ
6l4NaOyOtIIjs/eWEsGBRGqYhojlwN90JhT4xvjV4THUrdKjzHdN+io3xGxA41GA/oy3sZY6TGEk
lqMUkPWAOBWgtd4/sxjFr5DhVlT61B+B+Tew5Ewrs5XT+l/lr0pSZ9pGwMNkUDUJ8oFggj5cK0iT
sHPSyApb6tvl1b6aZ78FczwboW9hm6dnu9ssbr/O0/1F1xFQ7bU6AlW9IfTnSlADKz+TLBrcxWBV
2tkKFkHjWqEQHSI64OSNEPR4/5s9JpOQykXcHhmafmHzrbfMtHby6aS19Wed6qVb+pxf40Lrm8QP
JvX4JtVlLBkueqaCvFen5LNJIOHilkoqWdcmEVKjjSNGzsaIuI6QLQeoRUiO1Wksf4Q4WJe9ErXh
fd5x12jd09gVr6LXOZnatJlv99OT4u0D8IxcdF2rM7RtApx8aZ7TUlT0tu9LKNlEeA4qLN4FgOlM
gIRvqXdbjDheTGXaDbaokCNcLs/zcRto5u1NrasDS6E/gpE6If2TW4Y1B8uMGaeRL4Ix+baVtO8e
qpBEKAa+d7h6tJ417EBwycQu28opI7TYDVoMYVIK9vWOvim87QHauYtaMYhl5WNl8/GTvAmRVjeG
wipYcBL5Cg5Xwazw9SBvX0qk+bBe2mY8cAbHqZmPsjlbl0FIYAt7aQHqeiBtPqHOqQn2ZeIgYSlY
MNedpqJTo14L+7bO1PELux2wrxCzn03rD+LgbPrTzJ3a3Np+hpCOY39EiOX3wXGUMZ2L1Uxi7Gf+
c+kHmSmtq+xaFFsQDJyQdLb5PcFe6rKFi5124Onzfdp97OLi7lrxPzkawmVL8lM7uvCioot4wYaJ
DoD4yqTBMt8NImT16BrN4nxOAJGiyIV6ut0y9Kv3EpGmyn1TPBj9fKnvtL0140onvY0IHkQMxjMl
lXB9w+o3w9/FXsYQyKcWJjLVAO8gAK6gRPckHhCDDrSIw+7bcVZGQIEG0+6vR4faIbs/hcmfgmqm
9Iw3JkCoQUbV9HmBs7I+f2dXh90I2vASoqkETfZ0lxRNGr7du/NOE6gRCl4zgw1YxtWtfYgh5zd/
e+kPuz59BUnwpI7c41uExT7RHYid3HXLcAM1YOJpg9XJDEBtel4pwjcvuorxMmTE9wDbhNRcd8uM
ZAU0y7JXArCSJnwLe9rGysTqNH8Zg0UEcSD29R/o7g7D4IBOcJEvwEqchQidI6ycWmbpWX8zWHMe
fESqMOO11X0vF4ksTa7F8H4BX7TeCvVvxAu1OOTl9pWTE7FF8UDdTP2HMFmQFWl+i5IFPnvRA+hS
DyFcTmL7CNeit0c+vnpxLzcv/pf0lFIHr2YRHu3I5RNasP5R/ytmEQ/1gnHkJX8Djq8tY7+cRD8U
2KZIV7F1GJovovbhURTFhFyTaeaNIKYHcHwfmgfkgZfspBEyT1ZRsZqld1cqNK7JNW/aAd1Ze0KK
8qrni8GP9Fn7rcLh/Om+S8F8uD2oqclSq0WmkHtaO8zfr3PF9TvbQfSl6YqqjJcNdAn8B0JEvl12
5vefPow2mAwShcrxc7DKryTzLEqGru2OZbITx7ekh92B3IxQ12oSQCP1Kj+d7W7IzRNErXx+Q7Fn
AufTaYyR0lqIf+RPpwMHepJfSPeD9qYmSe3SLLbsesIGoGzLuPwjDLRh54Kg1dOSHcQnGnGjkXJ2
7QPFUNtYx0Jf+OOScYKH2AES+PAQFqNyPa0PKi8I/faNnMuw/188G5YTMNp8ernnRbxfOZzED2Vs
2lvgpf7PoktuJN/Je0FAJYQzDAFYflANLyZcKaR2h5J4QbIQyImH9yHkmYH+BjR96aMDuXQbWCHX
pWXRuATRD4V2281/LCGRpjkY7jUBm8MXRB1TolW0u+4nFxad1nxISpe3hF65OEzMr75uYx3QvqFO
44LquNZS3sKyx5xNa0mGcnbz9qPtffZQ83o69cfqIqevvc5zmCNjscjdqk8hOVMV5Dir/oSB6tCe
S8n61zK1P6sGKtwMr5kprjeR97sjuFtiHmxvqUF5Bo3aFsujUKOlazAzI4JEb29M2DbxJfsciZNx
YDPFSVmgxqk0VrBAT2MiQ1wt6nQxrmV12v363ONBFl0zweq2ZatUoIOzgNvcGRWPb4JhfypfeIWi
IliZ9SWthg6GH2bxQN8tHaiFWJQCo/pa3tvBvNJ2wS+O3dAx9wXDTh4P9jpMDEvtXT/0BzfSFGvN
4btPfUnNP4CDA3dSmrvJLLVpXWv82Ib7pdKr7ZHDX6u3ordBuXRmdADrVcRA/NiWy/IfU4A5oEwj
YNOyF1bS1z9wxmxxQ5v4MueRoGNVFOpMwenuPifp6srioR3lzVxpOetBmcWrT/uLRmaCaBjNX4bG
hG/2mOhZ6eN8MagHPj5BRV/CtJTJ4xOBBfntJyi8gwBbSTFcrD73s1VnZJwr+GMg1/HVPaDEKjnk
oi/lbVplsAcNlIdDBUXXT2XWFVxDs8i9hOb2sRUxUpYJaCwJgmzA7J4l9VyN2zyKpUQ6qJfPiMWc
AEJoiUNjX3wQYyc+NqWEXDk2mDE9SzpBsTSOm47Jtks4N0MQpAiGGKAN7W/4U/ElXIfdlcoeqcjy
GzvzpOw6eJM/sWv3TUGqSYTONWOVKIoyA91qyYF0ipQlTFmko1XkU7EAvbCqJ/lGw0b+4f2ojzTW
hblZSUz91zZkbC+9rH5Y5qfiZuYLV+2Zuv/4H+UFSTykvqo/M8qq+z1UFZb0fjfFcfNXfR+17E5Y
dlh/1AfP85ZmKMRJ/4/tk9JelnwvEEBAzPIufuyN8sKYVbXYuNvLmZ/DYMSHJo38oddVrH1Oa6KP
7r4/WGLB5PQ+tUUJy6sQped56jlyJwKKaRWAb63zBmDm9ilN0BLbF8Vn78xoTwIj3HxpTAclSFMC
FiITHY/4u9efEPMvHOoE2sx6ogrX4uFJRgkMWI1xW+bGYy2hgnGwKznoIIG6BfAId7VIMd6QrprX
e5TU5zd0pnWGdV45AhBZrOeB2BwzRNWDKiyd7KNDx8Eo7B/eSudCYmt1G+an//JpFUNW3xM8iPtu
udIKXgKwB9DRBDN1Y/jpyyP84U0BkLSyH0ZXgOHM12xrvkH1T+ictgQN59gyb0ntejZGwi39w/Sr
e+Of5TXWGSWdMzE9bzbv2uHZEfp9O3FGftOjWf6LdxfG++VhAQBfHJhbSu5hNvWojZqKv59M5t+q
d2A/UrhvADi8QDI6O9caLKxEoChdfRfN85wU2PUVXvuJO3FyRCe5zBjKhOdpRf+KnNVcLscLsRpO
N9OqdaWvyeeXLazfUqELS/qoIm1IR+6DEzlh7qZdYstLxNlAUm6N3ZMuxKOjPG0SnlVL5mKMADI+
Ah9PihH5xgpnE7O2JQPeMejFZoVg7GuePxuJeEx/WUb2dTibLSejSWNdZMN9wXvEA771W2y0+pX/
QsmOceL+MSOG74xSYB9pUF/IKXXD6bup5TZM37ZOFOBStQJg8U9RomSLvOuspaaaRuwIdOwTIJl5
6LwQM3DyCOQEk/ss9cV8EgqaygROo8W6nFe7hvEQOiUf4w+7PhYjv7NAWfWq81OZVawRw3KfT1ql
PRkHEEgBjtvHW2Ebe3d4SFI7+xdCrLaskNPslEprvUzZLCoy4SGsMm4fpV1NxVfWr2WTE0U+O2in
bI+ljlTsIJS3G7L2PPwFjBAgiJ3FOIpbhjnCpB1JrgULOjlU5S6cnXUf8v+MwA171rYZIw7r2yI3
JFHN987j9nnlfxZMEItfUdzvHDC0m/SgQbfqm0zhwyWeZU+jajWNT5znI+cH/kg9b3lwXVnWQiYe
vwcw9WG2xAkBVBa3JdEdBLzG+VwTgA5KD/NQVBPpVCJU9W8LerX+yJXUc0G9UmChSRhygds3AVgc
xZZKCmTiRNdMWSPX4SMnq85JXPUfOs+o+CuCP2Vv4shu7UNO4nfbR6eaQ2abjh4/wB8pN8F2SMoV
8mOycOivjmDhe+f7V2ILR7rSZHl1+bmGhSDTxLBy/9dYtwBlFswy58tvZdt8x4tZhDzkakQpLftJ
D0g+7NWiGqVSl6m5IOvQbS9OFu3lMWYC6psSDwPrHS4kR9cxTh23r8cFRhcoaOkNZ7tX9mpW4/PH
/pMaoC+aye7PRiSXdP/8HHRVN/ehSShjWWCApAVLkUhFKx18WVKIzXHzkYyK29WOZYB/uyJVnfYE
cLiDUvtmjEj+H61HpTBtHCtwjrlsCGsLlKE7pIG83y0UfL4nCXT0VDIXMeStC7KgomT/o3PMauZJ
SUJhjcp6w4qKnEMjMX9XC6M4tRbsAAquhXLPmj3p1fGuMKBO1GKT5Q6TLo9c5kPk6WECsBxkSSxP
oFm1eBKlLpmPpEMqNeDcqgGc3LG0CoTR6V4841McyTnDBupvZF+IGOBlOwJgSI8VQe2sXTElHtVM
wBgaQ3cnjz4fHLbnWp7VX7ilBmXRYoFziPCWbXYlY8WG/ujDwquvALQspTLabc4Q5214e5nCwxVM
gsPhWezZzItn4c0wk0Je4qPCmrrj2vsNXqdRNbN8t13vIoDjwLaqvtqgAMgwNla4f/rbp+NjntBF
L7oWs85flBLES2M2AaVCroIkVePD4KYsRNlrQrMGUO+1Z7m+bTNJJVwtHwPTz+/Bo/ROgmHNpQ7O
1BAigzw+shFxy6sALJDvFRe+QQR4PEypGvWOUMcQhZ84hBgOsaV/yfnASG1zTBDOYyIWJke2/7Ex
aBTMidqNkAr5Z2ogQ2cMsBRwz1Lz3b3vSH/HggnkSH8L8gzCZFIZIEcV2Mk816Rxf0d2/WPkJcD5
sD5yP/8ME9F4rplR1IGxLWlpfX63cys5Zrk2i3wSx3wJJfjyD13qbvm4nt+q3QuAciSKp7lHXFHW
XIOnWA20TcTIIvf4Rduxad8MaauM5pIQqRJJ8+vglHVSy2oPWx6ZIoKq9+JdTN1gndVZhP4jfEro
30DQGLJ6z2TNmqTBeEW5NVoRILMFKPzKyCwPCWnU43K58Alw9rd5dIY0ATWYUXiLPmzhCllJN1AG
g+zahdoV5+6ulRZt4D5IwZgRUhIUYhq7sNr/w86Yy33SswaQYGJgOtP2pcBdmTD4GhdNUpCuPT+t
+dGw5OmD/k8TxA/hxh2KcDyRGdpg5GIqqHNQIGfhzKV9CdTL/ojnfKkJy1BqWBJhz981frMEe3Vz
cu6y27Jrqb3AEn7/z8q7AthzQC1Q47RIxVUU6z77gcvCynyvve+DUDD90T0AuQd6mtsWCtFxjLpk
I0v3PV6UjVQAvJam85pQYEa0F5MKu52jGZfATkHf0cFlLOpGqB/f0kOn+2qn/R8jAT73QFcEPXQV
JXnPZhTQsYcFKY0HwGa2MKNAMDFKy4sJMa+Y0rmOI/sZRWhwqoGUZIfJ/dGD0XPJFb1mOl2U7pEX
B/ow28pFMpzRhWiDsEOEX3Kzs6GBfcxVtSTzFQOAxZjnEl49JQkwuye7RX7FPgCgJ61C/5ZafNf4
XjoXBYdHUihEuIj5jAszc/imv/769DzDEpXh9dc8NYKlexf35T9mcZUyhhdV9dGoB+mNf1dm8lWV
cm4Pf1dqOfPEe6KWGUKbnLpxCYfH+xZz8PA5ZwjB1Oc5yak7iuTf+UyPc1ABsciry8PY+Y0sHmwH
tHcoBnB13prPmT4tju9ulJELCq5eSZJBq4aUybUXyFK7ibetSgjJC/eIoYPuN4lRF7XVedAOoqhv
1rtTqHzBdCr9Bu5wd9jwdajl2sc6taUTPsa7sfL81Sd6XMb0Zz0lF41uJXweW33oOyi74EcNm5Ij
DShp3LsRIHKzbCTu4vNBsJ+6jgDib4M7P971sjMNw6y0IjT6RLrUK0kxnAJBKwVFxQJj4XumTZFB
ikyp0U7DSoliTeftoLnMozD7kpu0l7j8DaV+dbjy/xvkSFM1QWGml+Uhp+wxccC28IPtvr/K5ZBW
ScU3RuBy51ccy9qXtixHdzbntCRDTSOtvYlhv3wsoJMNt2mZHX/uCX+rJQxSRcnjSSfhm8oJaCMD
sTEbCQe5+CO71KqJlEoGOoU5J6b8x8QfkoyB14T1kLMmCPhT3xxLIJj2TIIKLIrz8ZyMUaSd1pg8
PVvEt6VtgFPyVgn1yL2JFIORCT/tLkrIuQxBrZhfOufpRvieha0ybPll8IWMq0iSizOi4iw+Aglr
MngY0F/TC+seFeQ+fJaAoc/VU68bChvpGobjDHkiAqe++4aFW+2Ai21jG7QkwP4a6IMud0iBg2Hk
fgapMaAadSHQpXvg0MAf45HazNe9cS+28ff5qOfGFEu14wmw3Rv1jEm2a2on2W4XKG4mUF1rMoU/
2BpyIP8JKwEFVfSAWuH+UxlccJePYpLVbzoP1uNb6Urxfo+FguKSkn1t9yTn5DZSNtMzdr2CG2eX
DE+lO2fopkeTYAdcJes98SO0omkJeeqs6Nj1RJgcvJDSOrMfRlZOmjoPPZZqnnmApmcB1U+LUUv6
ndqcoV5VwlcLqtZdKR8mJUtDLyj5TntYZ8QZLQWBROtamymbzBgZUnDnjqm+SaKvhKfaz9UP5K+Y
Fqm3bFuGZS3RPP4H3IvijF7QqzCt+iy1JmrmQgaqOTItNLg1rhRV0BCpgreZCpCk7ZC+RAUgOObg
Hf+pkBU8QxUl0I5NR8Q1XVt6F/Z43gaO9aVeISzQUflq91ojQ2htrbnuufcBz4/+oQrKl3PU4yz+
kga8OYWnBuGjp3grYviiIIld3cBy4D86VszOXyTzEdlZk6y8U1LG+kICJtCgvQ4rtvy9KtHL656g
iy9b2guBY685CJpHgXj0Pc1ezqPOrA/H4ZWNij74IUJ9YrF71JTLx5rJhfEVST6nch3sMO1kkF1D
K78W8nxtBMfdB3bbIa7zlb2ql3gh72Ld+9sc0/vL9t3/qplb74S0aIpp+hasu1hIXYWD8vxxMPUT
BvXRtzxaXczvxn3H3ZPauJl6K0z8gI+ed/hnb5AS69EIFGMP+ujZpb8RaHpMc7pWucFM3EPwl4y7
ieJd1iPX9SXBo4vHqGQ5g9pkGS/ziMJmpNQYfET4j3VIZarY7qFwKw4Pk+DEKeSEUmkBJRHoJHTN
4tU9KFfRi68ccHcNP5IzPZmCSCjpgXCoqlZMlnkXq0T/783Ns71m8j+Vj2esUnjjT50Sos/L8cr7
T2Va36d0wdu9Ucf1buu9qFxM5PbZLcsfT18CrB/WT+bc7CgT80jMBqO3iUQA2OLpwyqXoHrNEGYr
GUMp8M0Fm7uPlYNnHXNGw1NHAn1rybl6ehOu23eVMyNiW4fwCmMYdISp1ajTOI/QRegFgprxL9Kw
JaUEc0eo+ubpMdGbdJHmwyGKr3XbDpx7XVmzfaa252gFvCGC4rllNdxcLAFOBO0Yo2aRCwm8D+oB
Zi60IP6T2ACSDTG6mqK3t0Nsxm+ycMitGf0sKrSApY6jxW8oNuy0quQW35FaCYCsUtwDyo3CkOoe
dKB0DcnU3KeIF/KEp84nG6SJf1rkGlTIAOeJxPSessdBTdLfbq4jqZOVacMvy60MlZvDcUnp19Pu
qaxHtHy8HqZ8QfcjymIz1V0abVOELRogSPRC32+vpYkhpIA/vw7+M6NrJodzZOeKnXnngkcJIL7p
wAj1H7VI84l07ttPwPERpzO7RofcupQro02sUdqFjoEc09ZIVolFGdexXnH6n3BlyuLSELpGw8QR
upJONc1qDihrypBmQPnoGL1Yd2+oqVZra7yYueD9w7BjeL9rc6VtQYzE3jowRJ+MwI53gDs4kh7b
zIwK+iSvpzNkj9ECkmrVtCpwkY/0DOlb+U40lsFbozm+0CHnBH+XmZCOG9AS36rUP/yxmodOaxqC
YWXq1O9cRtdVaDe6cYnpgTUvB98ftwIsQVr2md5NzY5yo2WdZKHiWrOSGuWewWinyNjjVblT6l4U
jKEhtmcAEsBKRm1uP0q7ODexgM8HzVm2Dor1ivuzWI4oIw6c463+BSV2Thz0mjSaeQJ4KUU8rtBW
Ae+OSbktvZIkRSP+uCSWHx2THFr5aWnhIVBe6K30jd6tvNu4RrvBSwRI/0gHR5BtGlwQyylX2Lbz
/tMKzXp4fv4YxtBDRTBD0EKH1C7hlRhEyNGISeTXR8uIlQi1oscFF73LRqfiDYULSiNdDJnAO7Rg
L0Z2quXYjLUTxu8MiZjyvo9aZ6dNeP+tqX0KIh4SipKt3xVmU4Z+J4NKmHwHHPg75C/ovUbmEi55
FKeYcYh7bajnmzTIPmtP4DtZvNa9nzYiAt7ycGqJY16RMXoTzIk5srwlxF/bufzxv0K33yWhYZJO
RsFucVKgHkxHbjZo5dEUPZ5Us0xHXg/66T8pbzx3EZznRGPjJ9x1tsMz9hhbVlZMPOL4rBwYXPfw
PODaiF2fSdJKD5IiaQgqEw3SPyFH0OCzuJEjgM4IrmAyDWxtNiav1832FvaLgmoqazWwciqYpuGc
8Jr7E2eR2ak4HK7zcpLffzDn+f4b2yQ+aZ4Oizqy25AYUVRq9cRvD+FX5K1GJ9yr/fF1YNRVNyZO
5v1/POVxstN9lhbStWt0t7wbnSM9oh0D+XR9O4Hmo4Ki9LKO6e2RUe1CLClT5/8oZXGBVO5xmcb3
DR/oin5/tQLEg6bRPPZacTmDbKRHbCV+ee1/Td+MRB2BtXD9xyXZSXonNtY8Fjei6cdL75QIHLDZ
PPWRcH8NlQDUMsh/WAnT41eT5pamesDEeUMO4hfoGpmq1K0mdcgRmHNEQAkN3ByiLUsakgWmEasl
QQgAz7jjVmhiIDc6J4/YsZ3lIbe8rYPwK0s7k8txhuZQxXsIqSKrn8dq3qbPYTkJJDgwKGoSXNsv
GpGTSTnkGssNrEDlt9yDdfYixhYpui9vefBlSgoYz6vWu6sGkAvmriXAFcI/4HUuno/czLWSmDH4
GfCJVAYdS3kOGiASx6Qfr7/svklRoXfNGBzpKpLM5Cg98TX9rWrpAd/AMS8Pn0V0Lf6PhJ3JtfEw
oJWrAc+w3yvgP2HcCnwc/POZrYBY3YuxFg1ZJJIQh4jf/DXauKO+hkcnIll6erizuTGWdOx8stIQ
K/lA88nr4SjG+wCznVObN8zhWfuFgd5mnjV3cSHiOKyBoO0q7p0lRfUwgKhfFtg2zd999i9ydNon
xpwBwKxVqIk4bxkAzEapCwTNov7LIzKeV0+jHK3OxaprQnHxmuOK9oEacR+HsTh/iJAWRJoQCKbG
cd35pJNhDvr2TASp1z1hM5wahwz2QX8+ITYie8VtuEmPNZsb8sI7fPXqKAwYjFvYyudQpuwaSEZV
zC9dWTwatwtGy973D85QIzaH2yCnXSGDCPKAE0g+ZbrN3717mXBgiwSe2s+gvyQultLBXiElNVnh
6sj55geNixpY1OZbzVX+Dy8XuX591pEGygDtG7fgxkc/95cUmeXIYvctQi8u/AIs0zT/Fhf7qTF+
nYJPn+aWVulkqWEIceeUoVDDr2HI3fazbFPay7Gr6wmjGT1WzxQuGj5CEGDPLEPBxN+5EBoHd6Sn
Uph/PvttHLuj7bpJNNAYMPR3ceChxKSbsdT/81ImP5T7M+BRbyg/xHUxoAnioJ3oux2e9+yvWMbH
thDRdGbXs3F3JNIsq/6nApRUGg7QpMuF+oAU5OzlfhlxDfbFmXpanUeZ3HEs/q6ZzO8H1lqEP4xS
7qoUYFgB8H3SkQhGoJEKlhWv9x3F2iPUuRMKHIA+Dp22EQNbiC7rGnH/iSvUbFAHall9L809ZQbH
WFYyVAq7yPgNIseZ3Sy15k7oU2Zr+KzWX+bIGzhtjcpVJr4MRePbYnY1BoxKcanhGIotaVPVTGEP
bkDSF12Z9BjtOy6rCVHxuXuuZ6aXcDNg71+L+HhzdTEGOyuLgeDeCiY8jvvri2Mroa9YiHIKOeft
xEdIC6pI47b8d7nhW88rMaa1quhAiwBTKAA7E8MUNSyRp8VIxVGVgKWOgKKXfMLFUG2zO/5SIsVB
sOBvRyjQi+35DgPdRtnOW6TnQDknkqcDcBFANP6Ebz/HKK0KtLcivXmY5fp9m4IUtuAHwtqwGZ51
zLBTGMW8EF1uWINe7+ytFWLDEZOHJgGjaxHxZOPJjACvLNVb3wt7eWgjButy8GKLmL1n/e5ba4MU
8wdvORKQLY3m6pZNdDnC8dvATw8sWJedO+YrG4CbZpyukZl5OUR+rSSwULwzE1ygAfjyb7wYRIQN
cz0KQoyAmXK+sSxwa1BtJoOay+tSQfikouP1ZX+UaaxP8ZzCs1XpY8PPHuyT0GUtQ6IxpkuQnk4I
OV0fqD+FFOeS+regmfCaIv+ltL7gRHXTGDwdxWs/REqM+6DjjtPGm3E42UAHprUmtKW82Mc102BN
ljNlgqEs1rsvw1yNgwM5e776CHA0gtrdBFZTbTtmr/DmN30/4iP8vY4/Iwu3e8oNAtfdPk/Uz91L
oVXuQZeJEUgu+kPq5/XJfp0wisCjm4TEVPAg7++bm7ChciB+Cs8WdUIBom/g2aetG+5M7ImEumxo
54UxJVcJywL7wKmOWGoUhjOcY0cjPNlayVguCOt4pgAsql1ucN7WL1rhvmZDUSgXDn9iiB7Px9s4
q71ig5E2EZYKvian4aIKoBibUfS/78EGCod2sXQePGGzWSP9tToj4Ga8Pjwt+P2sQ7mtmk1kE6Cv
eJuynuYQK+hUlmzeS4BVYYefINiptZS/8pfwKbFjZAlvLggOhNu0ssWiU1oxRneFVJ0++BHntV88
MziKPMNoi7fyg/niftnxpqyzb/Q9Zx3CW1PtAqNKEIj6z7/xBE2bprQoNZ4c+XKYoQjL6Kh79KJW
y6kEx1yeb/jJF9ALU1lLP8dsTBTXdwG6tuEO4rSKdJUFloFdKHI16j5DVIb1poScNmK6ExIY7WlD
GJsKnCifpz4VBFm1+4mvSpft8caVdMzlqP9IL4ghHnkqpGamixnIpjRE69DBmHZwViUMY8UFo5gv
5rRRTkHdMnxb8IamMmQVj/JdRrfIiqiZpnWEBvgX+xYNPax/DMytXs4WZ54YSdnUWuovcxxI+fai
SgMXHyJ6pshzxYVpVy+nsQ+AqOqliZ4h3h3SRJpjebcj45Ed0ft3DtfFI1af8eClXvoIH2WTG0W1
q59dvkn4dOajahO4wy+3tb6JlSwsoO6TpmWZFOjblEifGBxftdJljH3MvdtUqY3lXSu3ySWzEZln
K0b1FC2fS2UYZMT3JPrGubQS46qf8eKUCXLtn7+onx0Y/zZmN8Zgd4NiWGRZlDaXl0Q/cSXlY/g1
057Amiwp6+5vMaaX/x4IRuprmSmgBwCOcCJevUl/J5FHfoDgOyppqQdT/pKjVg4LEa/YeJqLqFp1
d17R+IoyXfE5oi0+dKybUZ3rumJcWBW8yxpczsKu2dBURlFNxU92Eq0xxAkpLezNX4G0BSEo1rCt
9Tlz4rdiFM4W6c06DwHf+ilLlUuxhBmafGZS1aGdgTkpdqdn1bycuLA618fApv2IPPYLAWvMwO08
/ECdntAyvWVsRC9GpqYDuZNQ3YoZQebprnKew/GibS5DflkKChDLPIdi/TSyTWh8q6t8rHjhPTcO
C7xtaHTtVcV/xNu0Z3EMi4xJVIVKJT0XUQsVyD+eJO47tX5AdsN//fkW09pKrk0bgJPArW01IpmI
bVbI2rUgSGKVtmLd8Zl/lQppfK3xz7eILCGNVd1TDNv5Xo9Cwax9HvdUJ1zil28Hcf2dWPjveol1
LWEWQIOj8rGLPpLg81SVS37+VFZGpap1uHQYFfJysvwUX1FTqk2eZTnq4OIgYJQoWQHp99AEqPHR
ywta2v0qX8OIrWjsWKoowgPCUbAVGeZTTfig5lERNKVI7pr1dhP1WOkqp23KuRqoz5dG71ommJyd
M91Z/+g9Y+FWIl33sktG6hT40zxQLY+TkuG5Bhcs4ExVcxdMqkR3bhf9sYII/18tK7K71NPAINh4
67grgOfkDg6ZrYWL3/03fdnM/l2dIP7sV+wFtU6ijYVOkGw7mqG/6a4jEz8+TYPhIeus2obKpfNi
/dUlILgc9nPHTQDDQjAFLu9w9K4AYiyXCh8n7bsHf8lxzihjGbSZohG0qIpXPTukm6buqHO9vskj
RfdRAYV9TxSywU2TgK23RK5tRZVh8NooH0ERewwk4HeU0nze05P9a1l5RJkS//5gHkdh+Vns/5ID
GFXdJQcrcq4FxUu56g6GnGEg0D80a5f/KPdVL3zw1bnpji+2zWdjw5757mamD8spP8qlMUX5JI6c
uXwqCveVvMpttijuBNJAqLRPbhiyVWZVTD9B8xeyncGOXbYeJzVqv9Rx2ZhrMULgOtX01+tBoBVX
tKNV/k3P0rnhUm1N/waMMryloEqpPXru5FHFFOCX/ABnMICx24G6/TBlwFgRc0I6IkhVUEuZu0z7
SIZNENHwN9QmZFwLoRDUe/1/B0udjEmp12nI/roWVVF7wSTuqrFI7/T5SgBYw6TRoKo5vAWGYQGR
Qyduj1+taIAcQBs/ojF7YgKzCFJPmzzINT8QrL3czjZA2XK96RYNa0VZgnrEr2EMiU94QiKgYLhT
moRnO+nxh06Uq+uAicd8T/EFq3+b6xFhfzLoPaqwtZEWEpSnjIs62rqS6SSd7OdQBRbSF5NAsByG
Em9WPQ9MiQQ1vJXd+2Icmkq1fi5Yq/4OFfLNtcdlspueKEMgj0WmVYbj/kPLtKFf5yZHaqfJAUVt
H4KFuX21HT1p4qKNqANdM2cFi0c4ffu9n/FxJDLLJlHGHlpqFcdbDcWRjlPrKoOTprCE704K80Vb
duz2Vosqh+H+Yy7HClIAlPQ3xurvyFnOPL3yMJLYD7RoX+UOGnwq1bHadmTutFT+vTVaUa1HuaIY
S2B0ZeKFwNvtaY7v+quix8tdI8BueOfX9yi6jHU9eMGC1+wzQhYmNV/X01mf456IJHLHtIOHL4IR
WQaz2pxixqziyE3qvbnzPqXMjzClv/tRNs6tZlFVzzjYK9Z6mlBO1jptIlOZ8OECnUVmEWIg9itH
k2tx+x63hoLV3+bf6PbUZbwnqi7Vkw4Jxq8XlK52/x0qZUzsso5EjjjL++6vMKhNtIP8mjStPiST
AxYFNhobteQT1DHKFoU2ViZT2+3NN3LybqRnhMrbNajjELewoVAiBAnrfRekinNWJTA4TbHsm4aH
SdVBAd+ep6I52RjlqAa6AD4zi7S0K0G/BwKJENfXCYn/C11k+cNfaBChjf2lOE49xarDxq13v4s6
Y+NtlTaDfKqbBtgqHJounMbt743Vm5MZx969xIsJx80CaTVulQtWrTtJC0HjErLSUfd6x1zrODal
h5yIRmiE8ItSZhELucAbKIUmkXggVNRUUikzl1GpbkzuGMYNWiIKJgk16uqEu5iUv0bSfcESUF8V
UFH+stLNBkHnqrSnZSfq181788JaLbkP/JdYpIaknMZdXBXuuu4NyNgW4aOBWd/uw2hvqXmEE413
9bzIopnBMUYEAnrL4LP3oHsjcGSRa47EpgorWoCRjpQMfjJfaavtCWQLQ6Is8P2k02XgSCETzUrd
tAfuHfXH3Z7VXtBJ3AMLvnDx+X2OJv6c0AN9djJCLQoIOGaevkzMMqVnvhhqkPk943EfsrTKD3ox
fBcgDCPmCpAzTKCWaGYUVMiX5+87cHTRvPs0Y3rUPLcoFQ5OZlGBt/aKV7v211GgKwbqnyk4njZL
mlbP+XWftq7GD4rhN4aUcUayKjQS+2561V/pGDzYyJvfxmQdoV2TI+R+i0FTrXlWltWhOnNLFv7t
P7Mu/bWF9TUQ1yJ1Wf+qidE2BQ0J37bYHW2GobWdBxGdx8YpfgeECun0bRsfs332Ujlu9HIy/dO7
j8i7zHVnvPFfn/5BMYtM4+kBVhe/GBwkAwJU8cz8kdOtVmgKNm0W7jXwIrmc45ZD8u9c/jMfoEzu
Rb06dKXMkDVimRttHCievdBebcUw7ibcVQ6ZBgB13I4ruir5m3/Qt7RFfkQkHXmrrVDBHKgFG4Ez
VN+mPz2QVVWVJHmfdivB4w+cBzUHun6MUhLDY2o0ReFKTluoPbPHfAIXGshKcRFR620tQhIQv/OE
j9FRW+aaejD0llNa5GKM8HATvuSGA2iIXAVaedAPDYfS9RoqR2QAWCJoMLAEi997omJUewYsnFMG
TjB5JcdcvBb8PMeXrYrbWyd2H1De+ka7KzbI0le6d0v3Pzx5LSbOaxSqk1qvPxuyq0fqmKQTNqVc
yVDMWsnIPWU6VF3a6TMdXdPpy/3NUK9BokFn5i3RXmi+3lLvFmgP6UFfxEhwBVNrr6zt/6QMRf6u
UtbvR4mLPWkUvTlWMbpgLhqwTk+h3G1ORe0b7YmdMRcLxDb4WrzraExFQbZKe/1IO3uTPWuh96x8
/x6kMV2aeRBg43Z1lMlYVwImsMG8I1hA05oaeCHXaOcd9ijYZMAChlFvekNWhecL1G+RvCfzsrGO
JSje+FnfdCnBleS5xoxqIv10UL2Y4jiiJdERVaA4VzmlItA+jjMImrOo8mYeQnWRCyqhYOaHPDkb
N+JzvjSbvef/s3QdzR+kEQG7DDgTFuaU49y6dc9dt4r4O0WGryZTeFvyfRwn4Vtl8RlSek45cy7q
iTwq/KFLOh1nbDG/Ik3MPtuTxLCnGPH7Olh9noUKcMNpxrTWHX5Dh1Xws1vaO2gc0cqGmhKu8kH4
sT9WQMCijfw1bqLlC5WKWPj8yjbGuoMQkPwH5fi6j/YaS1WR6aTfi0HiqkpYGdae0QdRcq5o17ix
n1GNmmyuAfBFX5GhL82n9ISFOjZeqp58R0d/TvevxcFtHvaMIhJUP8MjNH/58NFDC3whLIojxokU
N0WI6jB4VY4Txl2ldCtS9fhax6Ac1Oi9x9xKJnAnYWp8Mb8kjvZRlwcrB3C07tPtfb7kF3njRWCU
eXggc69qfIzlN0TCMGCaSik/dlJnm7yv2+vp8fAHERupdYJKaxxy8hTGSTNDLkZa4Xtksc8PQehG
UtuZG36ETEVqjlRgsJHV+5YhGFP1tsHbzGDGRcYNlFS5/PVhmY4e8pN13oxSsvD1dASC46B3vLtc
Stt2QtysdfHfY+inpRdFtQkcVRZ31S88nCRgnv4/Eri9THZS3CqHBerezPsgmtEDiGoP2uwJZ9dM
KFbb3YWTWaYXplh+t6DW94COUWk9YHJgMO8mIWmDy4ZtQ5GL/Gux9gIaMJ9gWG82K3Rq6GBT4eXO
dou6eEmVQgZmEszxCG0R2XbqzKdfwX+BWbSFu71D5+8AGsarHq874c/m9spsnG8E+bUdB7XryROW
LUQfWlPcrKO7hzyfC0e6Cm/Ysx9Z09r2RebkNigcnVk6tuuQf/exdhL0zkqcT+w6ucJ+IBkcGAYe
343uhnhzwGEcG4pUdJynimeJvLexTl40K2J9lkQNNabcVMLnAfXSm3OTrw64562sB9CX7pr9GUYS
zAZhgTeRszj5sdtY9M+YK02llqYpoFX5s0My92pAkRbV7l/6IhIQyVbmmodhgQRLIv/mt6WwFxFb
xoFsRT2xs8Qs0BmPSS8fl7HK+y5A+mpqarQnRRSVr72qVIB8Mi4NIwlzGya/31hd0mPSdRN+ozgY
N/NUVqx+iOmR9LhR7wFcCMo3ZoEO7IsF6xcvw9srHYaeCzj89+TxaEIpzQ0Nu/b0crX8uKCDfkhk
8wv7tgegr6KLWmt2uFzZfLtUg1EZa5TMOZuSVR9oLxeR3piYRLY3mtcWxJYADR2YyxmjGsV3hf6g
Sdya/JgNm1BaEuOxqH6+VmPvyAFbJBaAIqNHBHGKT9GWSIk48Zga5/IaLgHaFM0cavAxqLtB1RLE
QYtNFKLoVO/F6i7rkC1csuSO9GZ7ucXID4sZUGVfcUR31uplsJPLleAC1yQmlcM9sEI4kpnmwnrs
2gvVBWjCpd/Aa/Nvurwq1+l/d7ECpSggI+7HXJHgjRARIBbZwen3KvD30tP4wde1B+H8jJ13i+IE
3n3TcnArcgjgg3spXmG+CM2xjXfdgTfGhVWmheBsBfi/1+p1bn/ykxTXijEXJ9VumI2BuAJgekcr
3KNxQyFBHGDqQWA5AQRrzBA+plbXugudI4oh+EAN9doBulrCv/2A5v2URaBsCWIePDSLI3BF8ZfI
oHvQ1yO9BqAqft2x5hXYlAGCuymaC5aGwc2Afolp8HWRoSAexVWLOffah126a1wGdQfIYS8UzLth
MM66BQatc+tUfkaUXn1jrH6Ff7D4ByvYRTX6ir+eJIHrywW1JadjE34qBmMkWjF3PzvNOqexLImG
5k85Wh81THko67MzaH45BjSeeJul/mUv+4DUdyUQtGsvFt1HGUR1mjSfggbsih1w25Me5tK2M1nI
CvunKvfSmj3bazqMzGWE1i8/kBAJUNLE552e3ts8JR2SJtGhu0wFeVia4eZDpYc4HdGIkEjP0bde
nzcAlV9Yyc6x7dD6LmszqJwl/SBK2lRWTcVwivXhYAYg2NplPyc4E7Z94yNDItvBd9pLHN4hMsr4
z/Uq65IFJgqcQq8IMHB9cJxEVifcAJd58NRlaO5jAqBeQg9qaccjAe/nrtwiNifGzfmidGIaPLyV
z9ScusOJbdo41KLfNxgYm0/iBvqt6agqRw2x4+fWUJZ2zmstiQCkeUWzkJIFh62sVikUtDsSPKwR
0N9aSjj4DoU57z1EFHdPh8WP/MCt8Rx5mDKB1fVidKdlPkPPBt5NZGsNs0keuGdXBtLGNGbd+WBS
1jBjuYeUMFdV0GkH6dxj2N0MxQ6i7THcQkj0OVIKExVbpNTOd/l/wrrEqY90Ki3yPxdY4yJ63hIX
t+VAFHLKqddo3+0dApu+ny/mUSNYt1+bpWwntH9qyVkX91ZPjR/3KWnF5y5w5WY5wgKgpRQRcPjX
BifkzXS39D8qZGKO1AM8sFEjjtaYlxPkSXPgOFz4kus4/vNzGEBTesHhlvNbjeDzCNk0AwsXsQ5C
Ks64XDAHK/3UCG3TN3aBR1dSSiOag4xzCISGDrJlyZOmHYRFMM52kU1h5fAOwu3UNDfneqPEd6KV
CYxxDy8nhv1chx06YPCKOAGFTta73GD+yfwuJ64OfflO9lm30YiXCpFw92oKVRnkIXIFQxAYR2dy
bq0ozB56YGE9F8S/I8tIrIZ9U140k3A9a2PVWbhcs4eU0vngmD5n9hUOoEWcI9EhNuP7iCHqyCpe
UfS7OqL1rI7x7IzPKOQDxed++AxwcZcYwC7JgkcQDCZYSVklpR70LZKegPN9vCpkJjVdRHH1EDwC
TQlF4uZsIpOE/FdUKanWbaP2AErn1y9oYnr19K/HeF9TQKx05W701ImlKWf/1NleIIhRKxNP7+Tl
3jmq2Qp/8tSyBqLKlASKr5x8gCcDOxVKk2hRDskfeh/I9DgpcDeKLRzQAN0TDg8KEnEcg7ZJ5wY0
brJpWoWM6fJo7Qr5olgsVIErS/I6s7JsRnl2PBdbANcz+CLcCuVCB/ARSiFl8r7et+nmRYHWuURM
ja4DlV0+cp97rl1qo4nr69N6sbchhAOmYgtX1fV8Gg4QyfeUjJJIJpO9L1ytlum4K3foKj5K12+N
afq/mVNOkRn59OzE2yV82S0j6A9h8WRN92QXoDkOaNaKWwhgYQ7KKFFzE1qABJsGQdOFsH91mYLm
hmiFPHn7E70IRCjQX5YDa3w8MRm5ObHelXMMfffmfebtRvoEslgXv+iU8tbvM7r/rOgjSnFdBz6n
Ttas5Tyrab0t4Z9R1Xtzlc617vgfnIwVcBY3/kte/2m0UESCGIX1FPskOPWTcUkDipGh5eFWzdMb
adM+dAsMKnlTsKMxuKEOzVW1YFuA6PUCPfJ+/BeCeKX2zftY2EkDXrsY0dKuxfX7c9Fpyj6WBVnI
3CQQ9F6WnZRdt3qLbmq83runuZBkqM0/SPTKwuE6c1P6TQorbFWWSQH/ZnXuFk+7DKEGgyCb+R0i
dAi6Wkb7TjHijB+wdaAyNh4Ti/2LL4U/Q+VuLxtC1n3BOzQEyuDZNTy/FyMuejqVBWRJh3TPItF3
+KSP6BS4FE0g1ob2wEepnC3izv2uzSVvUvyjJGeiMcIn8vT7z/AhM44iZFDIy2CPX0cT7SfN7kbG
3o9AruvnjXmHA2q7GDozbqYt2mc0jug3ani/3XANQc+1SouBJ30kFsIN1hnVVuDNkRotZhep13L7
eUuGIcWH+p4oAhd1+0VZ1q/JOG0i0ibGYu8s9IhEGr2I69xIFvsq4ZEc2YzhakIqWaa7bBfi+kjX
sBI1RAqQgfTu2d8BMsvYoH1awQhGybX4aqe06/Ib9p2kOEi1DfGH1Mh7n+PdWjNdmmNkBzU9dRZU
eOt8XRwpLzrqzfxfzDasJM8a9N4T/67JbmFvJcJPCFO9xmi9fjElKPKFEkp4eXD/CtubZKpCbVnz
tH6opjsgpRmYVs/vHrw212t4CF827wJ5lTdyBeUxxOLBycsZN6Y7YIEpTnmUKYWCGm8T2EFiJoIB
Q3diANfobQBaoClXvkohFAyp9o3Hh0wp80JmGjnBvqcBwuRUyNH99NIIY6kUZIpU2IDoq9L8sP6t
W8bFkOZaRs37scMTFHAjKchzRf11RObFFl8ItSZf8n3Xl8MEg2lgNOpTGk8hFfb8grOE7TBmdhdQ
if3fpiKsp8kokV0jUtlJXA9OKDBSPndxlzXvNghiXgWWMYGRCt0j67nOsWRH2kZyHtfYEJ8La/w8
QSfQhasOMa7XtjTBKoK/w9n8NLrqSoz8NIYM6alqeIyAZnT1l4BBCINKmDTRBsVFoU74VQP/sTYt
zwidzazlK4wQXuaSAHulMmpF6NO4035hzdRey4wdY2wqPi16j/fi5hcQ17zAR2jSb0T2nQlZec5S
PoUyukD3oNg34oQUVyxtI0kWbXpl3UY37DerVznvik/zrISFD4+2cupnXZIsmeiQdin2sa/+9I7h
UT2DQ8rZYtovOdEL7H+DgncmEkEGwye9piFTTr+0TlIgsblVbsuTgNmkWUIsNKsKRLHgZir3wsSG
VdblJPFP662lwJeNYI+7pjJ2q4eGXgDM4/6A/F4aU3d/Q/wEJUXqg1vBHkJL3ilH1viC9LgbmBKq
N7fkve3DDNty7zAVazMf8AFDrbtdEo2gFnbWk5Emqu0weM/bGRE0bZWXLPwJ1pjYgFqxJgKEAjiS
adht92etpMTVVPM/7F9plLtTNyeCvFlpi2hIouPrRr5O6MQCMCZu324wVFyJbf3djZwr7SXjgxR4
GzAz0xkJcim4JH2z4gOmoOCzKcHBA5+8P7Dr0NvUwqpDYX6Y/Lij9yCsspIZeFiz3GMhIKzM8IjZ
QtPA6rpLYoY2Sgwn2PQqfn3hzYjku5aCwK4acGqmOWUZBwzc/Yjd/IKeHqWvFFPOZ/0sw36EjTwQ
3wka5Cjx4SCR2w2H0ZGBCkG1MACLAw+r9KkDC00ER73krLzWLPZvI3RR2CyoQIpUYiHchcbeEzKQ
5EsSA/44DGg46J9Ru2MLcRpgJcg8rMr3CUh7AM+53dnK8wipNv6fTLtQKFn1CEdO03esIbaMLegr
oUhlPW414emO8aATRKqCCq8TLryo1z4tkhLqijL3kstC4F3XICX3ehFUNuNTdWLmlKDfIWnrlkzf
5GFB3Ok7vMuf9VUofxpuLkyg9sjDxkz/i7DNj62rgSrUUgtXUCs8DWufQq+7h9nMsZdDJIVoSVsf
x1r6nTrPuh+IfavwXQI53FzhoeOgXoZYyrA+leUmH/YV+GEnw6aKnPFZwgrEsnVtiFyTPTQEwWZT
4/Y9LxhhnOtO48u3mBKL9r5zkkUHKOWHYQ+FRiWyaQzSTzNN14qvwwCQnRUtgAmvPLX2InLUpC7I
bVKJrpC+r7hkwCEJxG0UUtdrWdcEloZPzQpkymz1U+yAlp6SciPdrdaq1qfkRHz6uHPF+q/8PgC0
nS6GJLTMozTO7agkNSOad+xAoT3MPNUiZndkBjv4RE6WwLMHEcaDxKOQMaxWwLRT/q5L777zPAUr
GX1Tn6Ur7yhOrFbX8jKthehPGylPb0Po9BuRS6Tv3RDFDEInMD7OdiGusQLQd1oMpORK/3qF2LpV
P57XGtFhohHm0GmosZmcow0c84g3w6LNOz27cX8uBTe0fsKueV+2eMcEy6xE3UhSDhMZfv0Zslxv
c52bMc/9cptN2zN2ToUvkftIbnE/wch4UH665mZOMKEA/J9ItY/zzU4LG59ZW6gZhtbCgKUESUpg
qbOV/bl9DiTlUQg9UYyix5ulqmo2xb8I5FlQKGK/qnS678FBnaC2gG0LEU5R0+qlczkwGsbb+QfX
lIzLwT944gWrMtoI8qOX7oKxdNFswD/sJVNyMJbhdGxHXp7ItTyf8VxQ6+xRcGy70Q+i6JY5yhfB
dx9qQpvMW3LRmwzRndq/5PxsnENjEjQVRvPlyWn8N34oFQzAof2I9Gl6nbE0rVchLzIyyaY826sJ
10Mz28EOrun7w9g/RruCgcMXeOUBPi7vfperLtUaMeA4bXNX6WecJzs2uVqxfO4ER72W8LZC0iv7
ekyn7oCRbo8ZEIP7L1S/UOyfV4j4YvPXXgJs6wPZVBazMWsLOCDgEPJF2D+cVkf/qQcoOky3raIk
tNu8vo/ntMPlEAbxIK1EPZ9b8EvRi3jg4ngEzgDs84pOyRmp5izEyTsDOniWnQiwmoMchxyzrj0k
3MgI9yx2UgR192wL2rKpBOKQh3qfMUCLEyf2xyJn2/XJCjeSavHIkk0lW9++8qWnppfHnIID2MBH
kxD1iMKjCBxudEykyb4GWIMCRDIJFL09qu34eMzZd1FDWoeHSa+H6O0QA+xQNtn5pKcjpYPn7DTe
+f6rUhmY4fp7oKCWVDfK/eYgYQ7PogsXgOHxYX6IiN+pPPoVSJa1F6FOd46tw6D49H0Bbhd1ANxK
DWvADVT6kfR1CYTa/n8aKjJhxe91Pl/hygE2n2uo3DooYmsndxgmD89Jo0yKlblz86i6DgePhwyA
4q0xv8p792g4nuvzoezIPF/oASkXmI20yeJgB/xT4Yl4jmm77zbvjXK4B4jHeQqu5saCq8ffKltd
NSYTEhZ/GlJE2asmVvkHt0cXY2Bv38bjlhRKZCfTAmqGGOOZer7T7ujFLjksIx8cCh8zoM+mtfOd
ygimLRiGZHP9mv0OkVpGfE+sOCDWr5XaYczJZquSJtmKPnuGhzzY/b5XgIONyGntZY4ViwLj0hVv
XdtcjFpL6/voq5EyYhbWcdcuZuMotD4QzHmSSm39aaF/uNa5Kz+H7Y5FOpdXOm92/Rd+PyOYoCn5
EPVyDQ02P/tcjIJZcQm1SUU2YS/vOSCypmJicc4ESyxbpMUv5fVfXymfOonbRFr/oFZwfLi1H07t
OtQHQQwMyKII9cVeMRvZVI8B9a7LheMu9/yiJ+kfv2TicEs1IL0dvAqlJX36r9Y/YVUFNhJDSkN1
SAWHbLmOIJJLTJq9gKEMdoNKFl3oZRq2yHsFvDtqIdRI/Sg+FA3DtEXYk9V/rl3FyaQIGFXef9nH
rIe4+fQbq+AAp0/R/MKDAXrK91L5FOWkd0qiPp7U77KcpSTnui2vvCjSt+IraFCh0MOlrtnvldzi
YzBwdGd4LpthV18dkGfjGAHuMp31o1sTmcA9rvF3RCGMXdQoS5DxAWPeukDuDmdMxw/475+oUEFu
R8fIiscM1mL3wdCklHunpvqpJrqrQNW2hT5CFkmiN9zj5Gu3OHVBkfZsKpl4fikBC++CvpwQ43Qa
g3f0Wo9copy2qDpo4uXnH1f/YcxrR9jQYIJV6ExwstfbgA9vuEF8yqp6NJx6zPhxNjVVlaQx7f0L
fJvwDRQVoR+mKfJKvogSV7UhJN/GLoesrxeMa86hGplESRE5f2GD5kWqjUzep9FRnBg/lgIV5i8L
tAQ44X6uyYiBntYD61xN0TsZAefF8nciBOoHz+9MGMNCP6v1lBhGu9Ryq/kWKSZHbNyVjV0G2VdD
aDrStGAwg85KQfuRg3owNe0NqdcVs4XPasMf9DBX7e0UAZ2KZCPQh0/dquGIpKMGgP2qMXfekdkn
RkkxgqM5hy4GM6X8wzeOqVKWOhhpL1ds9DFa9OddN3bno0xj0oGmksPPDkKXqmkP0t7zFKwLJjkD
vOsh45gdPLimA4X5s1VUF6NcZ+wdoZ1teMIIysBdGOmNbMB4wuCIcdaNLglydKgdbMRepbPlRHzT
MJ/bGKVRUfFabKCrNVW+v71nMp4Z8CspJrb/X31NaSX06ONNhNjqahbjJjDW+Zm9wC3FnBTMAOrZ
ZH5hsPMCnlFxZrv42Hm2rr3gshKVpFG6fJZntl9idf8WlrgR38Ehf6eGezQrp0szPsRVdQeE/pf2
fJJFr/WS2p8p2yvfCn2Ru/mTWXHuzX5I/DQ+jkKmlOC+TMt8pttKdGIJBIxx2fN3UHPOnLHoRJ29
+mqp5CZDQtx8g9o/qbaCq0eu3xiMlO+kgsSDiSvndf1lnOFmg9C7iP5e4S6O2aArPebapwtQcv+B
SS8DUWFZMHv3Fe/VlVYO+206lke7ebvepMaM7bN6b2w5SOQd3Q+NFR1kh3YwLqZwXHRUzRR9Zz91
qN6Gwz0ENba49Lb5jE3fIi7VpPXdv2jZlUyZL4msDD3cfI59Q5gELnxZwBCWABoApqt6hnESbzJf
12rgSq5FROYbPpTit2wcbpMw1V3NpyjRbIfUrPSRU8af7/2tih+8Sud26JxywWN72kizjthq4fvT
utmHHUjMIbPXpN1FEurBQW7p/LPE94YJlsPfPKs0Srw4XRCaYqsqkrztQ96Su67cy51LP+DE5sYC
yCJjqHA0522vYj1EPEOoHxgZzt4NBjxTJHnXrVUCly7QE2pcW57EwsbGYx093qEiufC/W51C3t+u
SBuvWeJh/LKR5p01tKVfw2OqzKE+N2F9Ee/Qz4vUItn9R3OaacxrX6v1TcYvUYx53mCPNiAslcvp
6NiYnXwq3gR7WHSEvnZ9ZjH0xTsFs5rTGWwbdhU8ypHJ060gGiJQ8aejUOwflBEv6LBRi1hhbDW2
kzodeh8D9NmAxiRScJnmkYUC8X7qKKRm8ZrkmmEraQvd/nvfv5tsLejQ3WtyJrq6MfREJF58onTO
JrlcGOMsGpoaWios7rg5AkzKOLSH5pEu12ZLVh4qQtoAJMAUICSu3ecus66gF0elFWy6L3OizulG
lfbINZwjQYz6UfMOpoVOawl0Mvjghiv+d6/wG4iWgg2Y9nEz3Iw7P6HHoiXzgnebHp6vMoWWD1SP
b18CsgYzbPVXy9ukS5utMmSePlaJdQQJ2Jwr59vxQEBQD6Z0R8fDMogh9QtA+hKm5svlAHGm8Q4Q
H5abcWyv8i7EnJiAz4ma19wH33EU0KZEKllouz6GJYcmstChQkR9EqeNU0sGer4xzeLF3V9Bnm6i
F/rC7bjqoZl2aBYvi5Mml7TLW/nXYBsj/7UONURbO0yh83DXuH+R65vJsqq4/1F29AFvu5PPwpD+
igQxDfgfrMVq4whsHoz3Er12JxbWULbCEMFppzYAQF1tMx/zkqQfvMuBjCWid9+8ejp6t7VLpkMU
7qUbcufU5Bq+vvA+AIEFy/KXWg+UohuIgZYB4QUZwvvLAYYOUL841lOFk+OLJUdzfIzoOiJMe4q9
I0DvpTBE5FjHLvOFllIZrA7moYGMUpsTIxRD0q2TaABAywa7RQsDYjbIm73ZsY4NQJBUY/qmFB82
xbp6KkJOGSqrviHv3xKr+wmqbjVGLP1gPc53qzkmpKBfSrO4MaQxFSuNiCnbMBq+hoag8n87c4kZ
TAosJ3XBg0wWdTkiHF8i0gWuY9I8LVPNUrkzxf8+hzViA8KK+CGnGUvagJUG79lux3b6ckyTBeo+
CNCNb0LDmWbrdN+kBym1bGpIqVu9Bi1Z217aPrqEzqI/ODqGkLr/P2+ldYnKnmI9kpsfLyrjscsp
2vJC1HQtp3OUmJmXfmjwI1q+7YtjmYVXQGt8ZzdF7fSxTBRHAxjJNbz7uvr1uO+a66xxvj31WLLn
kq9b+7vUtAgyUdnvhVan1yOFo3gbZ1rnB1OG46xCMma+kjASCjkUUhtLKgFfEvTnJdla0T7VrvLp
DcDKclZzT90gFcLRG4a5my+sYGBHNtAm5fI3l6vv4mWtOwYO1ta4IZraUZ4DWRfRr5C0lG4qg50O
B7k3Nbo7n+6/Ak9Ef54VI6rIXwNtLrIQFIllpE65D9HIWkiXR7WRJQk2Ijn0IA+HDjuTFv/S8GcR
bfVxanKcZnyeCNME6qcFKcmtTVAiYnJ5ogVxpEYUVQHqKc0ZYEq4TyY37K7vTLszvayBdOMEkkZy
lFhsA6V3Se/SMw+cMgHI7lrrYRL5e5aWsBiPypEZ+L4sfYhD5h5UphuhBktNVIge40ZrNxBJHD8B
wdHSd34JwjzmBSvji3BKRk/4sdIN4r93nGPjwV+N9sjVb0JYfgqq4X2iW//nSAvjRYEsToJN/KYf
9Jw9qAJPKBuXIIDci/2JbrbIT+lW+gGTYfJKVoFKk6+hRfusqgCThvPN8Iz6ipU+x/afHj5HdZTP
thY0Fqt7Qob9/UfG/Q84bId2ThpYbdxSu8ktU+rpLDDo1ON7+SXZrD+50M+97/QZpSfBm8lI7oYq
Q4vokD7PI4mnbbySaR1I2S8yyby3lbfKJ5O0o3IyBVRyISytN33YKeOXg5ZHASvy/dV2BotXNOEt
e9fW/1tCPyxfz+MHWzDhgmhuXcXcK3ZVC35nMwWppMytnYex1A5WaJBRBkM+1xEd+Av68EkY9/BB
BAwZ1CHySVFuOxUyblikT38O/FUFUyzSwx43gP9IhzcTdCWEQR6B4/AcYdtoNoFKiTwwlEKL/omD
qK7deoTZwlJfy5iVGkjRjy1ev7MyT3igrgm84Ri7ZT9DGQ70zpqtXmhpJqDaVXzobzuHf8yN57m7
m26HkG3s7W8kQFmUruluCywy8L70rXH94cr3Xa9Y8PsHdsySjWG4EsNlnxEnqyDGy5YDK5Icc798
qCjBLds4sT90wHyragnVB4sYlV5u5QSCkHjeBRXlBZ1H7g7mp+JzFlIHQVAcBDI2EVl5BL+wqobg
ij1LKlLt/gNDI2qWOsgHeiIeiwYMvxL9d9U2NHB/W54yk3Gh7UE5zEOJqBXT/lSqiIRJdPegHrNj
2AErO1cHIPK2CoTuEyqOFjuoRXWexPvzZ8q6gz7zXF+sfsjvxvuhdbgD4/4Cq+GRp+bO6cwgxM+7
d5GA55B9pI7tZ2CIJIKf2pA5IJz5kaDoyxYrMfNSOvtUdqyyBAV+Z9jJR+ZQL6eD/lYYXF5zaEBz
+KB5acETE7hstF+i96nWRYhZGS4OojxTzKiHcfWMbYd8CvWfXCcAnSSQGiWtgFIxLzSjoF0/2g1k
p9zHcyagqBLiZ80d5nj0BbkL/uIDsecsZDkGU+eOi6I6R4OoEgMucow+c4+m4tdGjPvlY/9+Gn2+
yFHA4aepbUv3DlGFLMvKJbkbNDXKRQkQyaLtH5rLRNvxXE6SwgA94YQAOjwlJRYep9vdJr+mxsV5
v/9z8ic0C9swBQA0QwM8BD5SULmKIWKfg8yy+vCVwcpNYOl0j7ewpisHVsdBcjc7ytmLB01bzuIa
Pn9rXTFtqNOfq1xaXzUKSikO50BVxOmWl71kzo1JoJRp9eQvLoSdlIce7Pd2lFavmj8hjvJlX0TW
oNfN0q/1HQ49qexCpSfL7AitXJaazxIfdg260nfpanAs36vV94/BslY8L/73fhPP+PQGrYdHSNkn
J4NZXT7tmGWeMxuVdmJYQaejZcEoVxP/teI5mfJLgLs18pRPMSrhjTNQ5MOCItoKCfAx26XDxEVK
bvf+F9gLXzhHwRCH45JLpiWh327QEEsVEaUV8N8Ipl/ghty4BC8kilTCd8TQ0KekDG+9+ggAMYFl
1Nq4do6x8YbnFYvb+7sj1OKkmcI9rd/f+Am0qaxoD4XaRoBBtjH5RvyNkE2kT69RnWyaFj0ZJre8
ZRGTsWCL7DQGJaBrETiZL4XSoxeoXDUSZGAXzG9bekilH0KF5bcR/Xd+NjREnr/3v9Y+KjtFViM2
MIibjedKFD1ILUGL3w+H3dxSKU8uBrNeDPIq7Ld52nGoeeOfYXWCHVgv0MRwnDvDIxZ+1q+DStjM
jlcV15F19Hs4YK094S1uGcvKNyeE9sVueNqBNqmqKjYaAgRGk1ntQA7LRMl/dAem603iECgb3x/6
F/A55K2oEFgtRGwy05ZZ0Dglq/fNZ3rA9g+mBt+/F2fB66ZuDhfcAUoY2AAg3L0MlDhFbQQCxv8k
3K22Wp5ZWI36CnUnYvjBeh1ZyeRebINw1kQKNgrjUJj3zcjbRz6IRYF/uB41bvn1lLBYXlPXvGj/
3XdfIb4wA1VUIY+d5J9zdItnb8i2bNaBE7vr9nboiCXPXOf9UfZtAgXaaPnLLpSnBVxZGr1vQW0O
K5DNkSvGKbOR3epFqHxi3fWZfxcV1rNsK+MuZtKSuIuR0imjeOBLbg+RSP/FLe1vHqIBxEdOeLFS
sUSZaIH331TKC8TIxRTat1J6kYRJg/GZTp70NYxfxKsPcqcY34b5DlEmco6CoEH7TWz7hrv2rTLD
9FK3XBb8qyvQuEmbxlVgjhECAZezfmfJW1iubj/B6IxmIPjxaFI9SVTot9j+DpW0NIo7kko3yhYe
1W8xiwTdzKNOyMYJe5LpwnGxVJFt2M5/LRTdhb1ig+w/xr4FhOTumHIuW/pR4HKyB8xz2PnP4AHk
E5XXYrFAEB4ofid6hW/dgde1Fue7oB96FAIcGBCfIOVoAcX3ko+2dpohRyGf8qVaUEhwoDO3196F
wVxI9A69t1SBvCisl8Tw5HZp0cGhqO/tm+lVOJdMCoutEiiYpuFwdOcKBVXpbscWBJaFJHoTlluj
0/X9CVRD/pAHNfsNvyWMNCwPThpcR34yPvx7QhYdoKDlul/gLFRiCkgmiKaO5i/+QwvfaBR7QQPb
iMuIYdWcGlYbR34ptrCtA+jOSqbpwVgRu1b5DGk+4t8zAHIX3NusIsTk7HwtikpESM+jj68anFf3
CNSe+CRNYOzIi0VD8RrdmVtmUiL/dKnSr5rh0nbiq7/Y1g3uL7nOQMx29Al/PPcvsv3aBNzEfoeX
0mrCHQiBetn9yEqtySZ/ZaVn8CyplT0IPxu8niTMWm7EHP+PPdO7QLmP+wqYG0NSAmWgT6e3zO9d
bXo40mvfg4wkTheC2I115/ElX5UwA5OAJJnNlRnNjAurMqT4EYr4Kzpbku+gpEWIiQhynfe6FMHy
jPsThk1nregYk9lm+AMT64WZ8ja4e7fL6u6AQ89Swh/tOy/z6TFAALKTDs4m32gzJWXt4vR2U43V
FxnDTFNyLK8TQuotLS0JCHp7noWHP0lS3JvvuwZie4kaUeWGuXSOGdpYKkwEWvos6JNXmdcxkWrY
qMzxDlN/fWvrOEJTEWExfjrCtUzugg1DTBwa5eJTMgv6p2YMD7x+elc777lbnrkAwPbuNXUkHHax
woBvhx/hyZemTwTDWLj32M54AVIb9vzp51q2zs9cZWqNqQR8XwBcOATwjqvHQb3TRqoilrr6Edxq
iyuXrP/UPDZrRYKlH1v8tFNB8toDgyOmYiDAiYm6x2j5dhPRerO1DG14V0GDvpHB+ZNLEr70I8dM
KRXzbtm6hQW8zbwdFWsm+6Al1zsA5tVadoWwh4nQTds1di1Iq6OTvoKl4p4yZoyokDO5JIC/ONUb
nycSy0dheh73Y8vF6kG13C2pi3FoAEqj4fdojVX72YJ8WgKsm9NVwwloHsGNE/bRdUHCZjXxcG8y
SSaMk8zUwBP3heF5XlWEPWTIQO1EKcZ/FpCg9K+K960gt+mRFQ/h15DrP+cPTI43NdTL0dCTrKLZ
upcmsWDC21J/UM4xa4m26UEvbeEuzktPOuGUk+0rRV9w4Uo8AVLVGyabwLrUXJ/GQUxahGhx0ESe
k3tRGvtEZ29l9KZuYSFsQ7kx/SHsW0bnEpUQ/z4t+ZEkuEKGuD1/oAXwhg8HGBa08Z+Ur10i3w7a
WPabW1yu6eOZubvnV4lbCi83ElryJt1Fm8xDN3lorsGfT1Yql6czSzsxUdfiRdKaUVHnNSAaHECA
+u1wBzVy6ze081f6k6FFER/h7AbTfWSY9WNgC5sBlj9eAX2N4ZcGvmTNLymH9DmYH1wpzBKf8P/F
1b1wDYnD/I+hVGceh0jgqkthmGaBpxJjGMgJgtKlWTjXKKDR/61vTUd/PKLBWHWDFZBMtsHAyM4Y
aV27w0WvtEZjNWjmyJmWX8WN5minNldnOCpa3qrZt1gcaW3zcjtwK/sbUkWrqfByqSflxFAe9A2y
B2rZuOkz06Gw+tpvTXij2BnvpQQkuMvnBc23Tnyb5AKZL0xuBtoi0CtLRrvjOLVYEG5F30e1pdNq
1d2wLAq9OO9dSvDa+vUj2Ttfa4FTWige9SPA93zQPPJtpJlREto9Ng8Nvo/kbnadZqPCOwrIRRZw
ok/2a2JUCP4MAZw4Tc2aIqcbVLe9d4k8AJb6jFhvM5bYCJ5vQaRQqQ0GH+Vp6S84QfikWVNSttqZ
tgoOJK8XiLD3s/iAui1IsYQiUhZacdwWuO/OK96Hm5GZtO/eGkdxD9yLlvkyHr/Pi/UGwZTD0ANi
AhndqKGbEE6K5DAsjCFHJQA63v4H1IoN7oux2ABc4CJHLiU9Pez01UNkYlSmxlnWq8T7wBRHb5Mn
K4ObJSFuSU9q38GzKI3W7jfAGg0YoTPJGirsx2CtdhaaBHDpD4LDRoqywDmPwRQiiNgc2jIJFo+9
dzudLmICYBaxxDSgNdxMsVd8ZOgk45tmmxk+TPWl0MXd3Cz9zog7QclFxvRfgd2Uhv9hkTFzAUJu
3WnAV45sv6hR/gi76QZ/pJ3x5y225VCBF/PXcpVcxc2wg9+fAAuG6FU65nkBiCLPrGO590z0ml5X
zwX8tg9zdYqkfiVQEdbcvKRbFzYvpR4jGQqrMvqzIXrfAJQ66TrygCq0UjZRr4XrBiNrL9rBxQfi
oFH14NDVXYHzKa3W74Tm85lqEAYOlGfF/oz1AmEI0eL04JpxBpLEAfmiTVjHmhy2djhU/9WaSDq8
9HdMZKxjx2br4um5nE3NmjqF+pJnNqUAtTl6vkfXG/zMVPjxMeQvC/1wiEOV03zlv65oHcB25oJi
M2SmZ8Mmr5GbzYHtLWAm2dXDnrnix/RQ+YxDaWORwbJsMJ5UDSX9PFLo3fnYdR3FT1Vyzkk5iJvG
9m6v3Vdh84Kp305CaIEcYy1DA9/Dm9yNabewi0HRhMx1eTpZm/2kkfYrEK+UVrarGUB5Iqmb7+0B
KWT5zcPylnOHi7CrhZ3DaUyT1NwmHHGyAWVqWMYqqXWNRUdoO6QPveWRDIiws4Ew6gqSmqddbu4d
QqNXEVl5dT8ItRJ0dfsl2+a1N67RjFVAX0W4iVBcvSrS5ZEscL/WfiAa8+0wDCnGBPBidfPlj7Zk
oSez6eoiMAaaq0F2ti9W8a4bvhQg7zAZKeAjlXhzT5bOV82rzJpyk525jat2M04kyF2dsfoJsSYm
+SutUUW4ds2IuPbotE8UUW71hKvqQ9+XG2nvXKFrJAtotBpTCsolAlCH2jCguMhkrNk3dUor3AYm
CcAlpjsedORWXA/VWXMTP9X9fkzXS+H/xIVR25EBvKD4a9LRQnTDre8vFqkGKRfOW/yB9oxl5dyI
6dDiOgFQTqTVBfTxctDPVlT94IrxSlgOQTblpvlkvtPZIxGJowvmQC4PivduV6V+ScFnjy3ckA+k
7hAp967iT6DUuDMZAQgVDG9ouKTjHBRKLE/5KbXlT168Szqh1eW9MbtBLJVR2sGWzoqfaPvnHZ0Q
77HkU9qeLN4HorqNho1P3xbFvQCWodVQ38RFStrblNtjIfteRd7I8sv/1umlccyeml57P2g8jljU
VYn8n9QCBerQkKh22EDuCOwdjPcfYMBThFcbzQZ8FiMnBNrBS+VGXwegU6NB0c85Uog4RKGAKnny
6EvmvBkrv+3YyNL/RumHFqKiKeGdl47tirhI1FRxbxr0QvwpVvBc53KI+Ma4R4RFp9ZknO4XRNtd
RwCQKgwrJ7IHgvbyGlLeRbEDnqTZzmEacIzgvrwTrJ3AryYXdkIDJipfXpH6/BEZeQLKk3Bf3y3f
Qhz4dOiDjBuYtsX4szKxLEtBSIUqYTNy0yWLPEy0anVUshmjrCawzkjRw9qjkWg9uIHsrexp3LPK
ATe69pVE1fsFgeB63T8cWudotHG6HrQFmemx2Im/YsLXLP1SAnnKS1buVlkUJPoNNF9Fh5lUWQmZ
92d6gwGP5D14C2tVbmXp+UMG6tnBoeRh7oUKir1oEg7EoDD5q6Ks75cPe+VVNZS3n4TktSjRaFw5
nR3GLs86wmI0Ea9SHE4+/qomU53II6UO+ruiaZ8iHmdE4JT/ko69R7Ju2mo2AYrOvQKTZ6cvhZTk
qHxKjftJbIna1olTsXig5BnmUec/7kHE82x86ClctDr4YEyAK7fRRL+wjRCfuk18S8vcxQdlyl+o
xy5/2wNFkUShayaOSJzF/nOEs6QsAD/CtBXVC7lS3F1GT2YC+aVusVybq5g6dIt+Ov5/ur0UXyaw
7LYRtGqT6tY+5dgrJ40A5L65T6kj3RJEA2IG05VPqL/uoj+tq60EUJH0imvoTysqvxeWXP7iZ7IY
+nCEBmx+sGmaJGKPUTxAODQikOrFHUAKuanqNSpZmgZEljWtaQE2Q918b7zdZnnlMlcimRCus2Fp
UQml9mlKNauNjK2XavTqKA2yb6LzYjBS+fBldFeuiwEaqP32eOPYcsMvqAibZVAXMBXR+fgKhEzt
0yFQXMTkFQf1ArEZCn1CeUTb+Pxr4ONPstjH+D2ugw73tZW+sP7GiJAMIBWIHtwrEVHEDgHr3UFL
2CNwH1L16L3FSSjSZFEuZW99qMnJVyZfGSCYTa/tdVMSVtNqDwOqT2lP/yXxc/eaLnSvxYFobwfS
7+wk57o1ocryQS4bDFMIrAwirl0WPuCdevk3tpKygXQNf0oB2K0buo6jj7XyluzQCouPMgWE5+EA
vl26ItF6i1/rlKEHixDkTrixPR7j6mUDpHJbipjUxPR5jBCt808zwOhImaDWE6ydjeVKlKMP7xWs
PadLm9u3SUNztlY8T/aPvkzx1yauzgWD6ZkiJU3QmMFEvw7evsiOMPScIn5LOu2M/hEPj89ck/Jh
Ce9RYeLF2llGoISEZ0inbXNytUWvOkLE2rPWQfI+KW/hBHQeWW8vP/4iNF9uwZDrVB5vH/25dlxC
wi4bVj2rgsTPwQH6sJO/9lkdMvd5zef9ow8G+LMNSyXoyE5gO/3MdPfwo97VzuwE+HEpU+32pgfW
qsmEcdpEBR/6IvYx9Z4w2nYdu/Q9bDOWnCNcYhkSvv+LC1ouA+CFqfUvmVLKnp5qWrS8z46rzNH+
LOvNDustr1Fnx1MF3guH97H46tbLWeGvjcB17tSIPUe/zmJGUo1BP/UfE0X4A8eQvXlqSgrGi/oJ
Ad7+qA0sQnrwf2Bo5XSAYzphcHfk23Bn77PYD+hJaKAOJQ/1E+bACfkT25WaYdFfm5PpiT3+Wk8V
7rBkssBVM7xJvHEERvQyftnnq356h66B7Hbpk3htxeVHC0JbYoYpFsOjM3/fT5VNcS18etBX1OIj
j+NAIatTFlsnVbdU9GEiYOvM22wEaUJ8uocWt7y5xHkTjqIG7l6ewKP5LSB4TQfztGsNmZG0zDVU
7YqjcVTJeNNdfLusZtrDrOJqfrwtOgntH4pI85Heiqu4SwVKmKIiRdsmfoCqJSQAWhYHZPtzeQyk
MFFG67otRNRcD4G3Op4tcNTEBo7mejMeSrD5+OZBNlntFjuQ1N8ZztxpBONVgGL2ce0ejTjEvGs6
1yvZBEkwiyJVe5cK48iboVmd4YWat+uVjcgncJxQNnnGW47VPJHCGD+9c6r0lqN8wQP96B4ELcvk
DWvngh05V/BcwtgDAMfyZrAGeWRR6vLD2vJEbAOymcu2b5mmPsffCL3tcFFdUJet4q6N2s6X69Iv
nRGzaso6Dxi5WJ0t7r4p540IVWdfOv9w+/eBgFC5NHKkGfJa4GOvvEKXsUnBC36HNLNrxIxGa/YS
elvZse+KY6Y5zcvkB9AOoHhlMn6zGg7+9b50afqsmJ2LXx6YotgrerJ6lPjXWgGlEKZuWdy7znjA
+Ak8OUMIB1ZHXRt/v3B3RIhrQFomVlPuu/DfBvXqvNmgnSFY3vggBzGFVeAhkZyLs86rmh59zXQs
ikmJhrFwoRh/G5/qLlcrjeHDfeSdbRzDrNShlalWVoEwhCkmS8kADZ1w6pmgiHf9GZOXpd4dK6hP
RmGhfgcPZGZgQ+LdTgXqYkzAaddhpz20HupC9YflPnaeBRnyqogl7orsCyuZBnKcAKEoT0zkl3Dm
GFe+DCi4XRe1D7T9ENrTLvLJUioHQuatRBe4gg+Rkj9L3SVKcBr4WfZ9WR3dp1Ydcj5JeGYhSqE3
IgeHPlgcmyyNUpSGsxsJWS0jaWDVj1XKOyv45WBJ/i5ACwK744mGFgzODJ29f2GBljRUz0pqdoDE
macXLFFmJC8dg3w0u+/gpOaSz83lAFSOgUrTDmm4nS2DtkkV/ZABtX24sno57h6J0QXiAx4F+MrH
UStEFVf7PnnG0Ri11rBtMIDdqWZCzVvYZJd14uOr0H6+lJXTr3lr41XBjw4g8viTWhAMh4KMBlUE
CL2HlCTru7QhiqkVLHZTXJITG/HI6LqX/a+/TA9ME713cVr6vWwpVCXiPZcr2+sI/kVWBY/6zNPe
OnDj5G09n+KeFXd37uGT18Oj+ncjYAmye1dXLFNB5bQMnMgNpfeULMf3LOC3Px6L/OZxFPy7dpym
iVmeE0zIxdXARsJIqqOAJrqKGhNF+m+E3ZvI4rnAhBGLRm7Grrrd3xPxu5MIZdntOvA4cppf98a5
G8DM7rgifK9/yRE/T2Ar5AismjyADTx6y4LoM4bIG8zDHKo8raRRCcG8P9V3w5tgCc7ZoElaEyZw
b0MpS8NMYbZka2J+51gp3I5v1jzTrbH7r0SOiFT68kFs43Q6z/lGqdzcAURHpDD6oefrd9+fsXUm
6ObMNnFXdP0R0krXwhTXT6UylTDpo5SpPnZ22qTPr5h44mGGIWEMy9r2AJbFmEIB1hoTIoUnANgL
AJzDZmitYkpLhMKTmfr3lF1kleV+/ZeC/8aqFUNrZbYV4XNMfn0YCFJnk3hWJWxIpSPFTgTNQJ+O
/h5P1CzwD4gKxvpYknQvS9xu0A+w3xiao2Z9aGtI9aFUHR1wlohWB1BXiikws++Uo7OUTKW+5SuV
9UPAgUPOcfnfjRDkfMcvlH7B+sS+rRrCPEGm2PGOENfrI9tDH5tdntZwLooZrnguUwffyq2ILJyu
vRUu9koEdGdbEs/uK9xPO/jyLh7kJskV6wNkM+RWEoaQww/rPKStydpLZnARa/RyPOkqWl6WKhCD
Ii87F5Fg616fL0/Hgpw3vWYS8B/TUX+OjdpT42HS8fJfqh6fTKdQtQjAHkFLOcPUuRiz9XG2widH
QyI94ScvDNtOc/lk/KcjB/5zsqRVoI3Y9zgaIQ5d6a+nAT7Kn1FApPuieQGqIv9v7bALrqP5yLIO
of9KuZrbp70xeFyLPCT5Hw0a1aI0Vd+AgYE8cX7WBesGT1xyRYcl0KmcqHUJKi+qvkhuT0o0fatf
LAsdpi9T8ztQGn8adAkV52FIzPPXqKKmi8NsuEZ9eXhMrln57xA0/aI5einqLWYytxUgLiPSkhVM
+d20GBFPnk4UMknEtRRBsUxbDZypjbEfU0CuEoG7NwfM64ndh7wBwpi3Pb7brGjfpOtCw4z8kWly
6U1nBW58cWl2j96GzKjee7ONQYiEJM4O6jipPN5ujf602LTa/sl5usXF3kI+EG3aSlNFVLkFmNO9
OrTcvwi9mU/FhqHk/KMcxjIfqyXql9Rc263EsYx8UnB2B1rsYX2BZsjAXy9T8VD5rQ5xSoLkzhoD
/PYHmL/KuW8xvEH/NmC8D6D4aMRc8ERr2b4tXXdDiVmpLiOXBatqSe5Z4q9Hz3rLoJeAutRnnwf+
D5+Pw/c70vlRVKE7A7gIQm/krVNMTVmOpfr4z+jO+myuV+brr6GZ14J5cRJV9zkGvQnlp84Pfz0U
7k5OJAsKNtkrskqg/QiK8WYg60GxE+wiRyqHE7jVW99kHDkiJ6qpjM5bGizrjoGAg7OiDRHpQMwO
oz8vkMHP5BBZztWsN7bRNOepgprtKXXrMlQ7eoSZx0T4S+sVrKmYUu4njrcBAmb9f4UArTGNfHmu
0+0nqhBrz33Dr7QRLhqZvGlgJpuI8b+kR7vtbzAsVJMgqetBDitp1a4D7xyRekcEVaQqVdbBn2h/
dJmDCyK8EUMfcQY4bt9cnnAknTCM6HbtnYx6pE6c8SB+JyDLXsH3GTL6/1nnUf1b0k8Hz4JtEtg6
0EUlT8oTtdw9Ldde4jIl/Of5vNKCP7rOujgxCCOJbKZnXkycLF54ZEmzkc/reWLdCvMfkttkV9MX
yprgj3OxVIWobbF9dSWus/+jI5UL2Xp7NvAv+ZVMJRK3blVlEuiiiHM4B0zctC8+RjdJ27uZCOdH
PAj+/90RfRzVbB343iE7Xu91hC3L5I9yidViJqyuXxi/DtLBFjRH7UDVQEe9Z7Xf1C+lDwcgE49U
JeRxqcpdcy4RfBqekTu/x/VAnvI8LyJpF2GQ6Ue15xlyeygOexdtGFSE8SobPxq26NkERSTF4MC7
LdsSOFxH9FIpKgVkWAldHJVuwj7gFv7Ir9IHYSRCIrvNDzYz5RzThZTVqgZlRLD+zyi1GXmEMKE5
HzNpabAFJ6/j5nKE39yv3ClR0QOnXV0ipnz40xUn0kjAVJFKEW0kVBdwBsCrO/WjqYcLdi4YvJcu
YKwugiJOYR7+M2pKgCjfZLM2TlqbDCv6bcSf661o4tWlOpXZSHNtCTRIuTqS/ldG80rBxC2nRnnC
Llu2A9vS8O0tP4fJkkDphSHTKHvwkMWoV6VgzuynIwdPi4yzthbPpFrZKWluFinxDMcdW63j7QEn
EI/TULgun6ZaOUCjbLkSE+aAFYSf5ofUa7oesALoIuzRwvFAXFXk1SSC8Qnda07ed+zxaXhaBlbY
3soo3G9icObH+Ow+3I5eAhtdEfUJbRwQTgFN/RrLnkwdj2ftrX9RKHf4zSMr6TOQoqqztxMuipDK
o7iM0ewiDAUmGppSzcjiwlySrh4gVhBDtcL901l7AEgKiOtBfraL4zrd9AENvwHGWfpquD9VRe/Y
4M7C9tv6Z12RpKsiTkwR9DkyeXUBEJhsP+4jT7kD5bLq6f27PAWOIB4/VV0Yeh+ZSgomLdAI4MxH
2TM4d9CG97tc9e/KMssszEF47JA58lUk6aC+ZmfxsvbJyo2eV4K4zs4q5QSSaU1Ld9ogW/SOfZfB
qMVB6/Y8tLuY4/UBwzuPT9eWti8KkveN5qIKG7BnNAmz0Y5QJZHsZv9RNCq3DPITrSM7gLjpe1FT
kQdtAIKnhuk8qx21DTEixEXHt0wumQMAcCU90c0Mt5YLi2IB7ycuGt1xzJPoknx1O74jTGOcW0gS
yR129iPDsJiu7p1GYKkdG+ZXpwRqK70aqmdYm5vnzTQJCjUSDZwDwH+uNBUl6CeoE6zbkDrrK/Kq
A/3A474ef97EELYIO953WtIfU73TwZAt1w9+kVpBPAQaYkCESi0dOBykKd/uYyGe7oJWAo3R2vYN
AEl2v8thsL2sh1xgmEwnO9p354v9SCOQ60VXehD00hR6zA+LHa03PclNOU7unIqTMA5a4cHYCDDv
kGPi1bKCcLG8ZjEKliyMHl1RkFM76eKk46pUgf+tIkkFXFpgZGtqLPUKzieoRdOQin5puEbNXLzU
9BonWFllRQ9j9wl7SS6vTJ2fys0cP/DoAkAk/he6mdNH5KNfpWgSZwTpmsXbhfUxNzCtcEJldyem
iKpJolKtqjGgrgv0o8xhiTFGWfz0snQPHfP0tnqTrKGubZJPTffAqpejEhAm790+hn99izZ9XaQO
nca9qNBn6BziiHsX06jm4pJl82pYqbz3CncteioaZFcl/LOmk33cRQnxi8Bpy5epzIiaWVBxwLz2
TT23wDZT5P+oCyAIeGGwEniqicaaiirwcMmq146RuociGFaBtxoZJ38aicFx202Td9nlGNlZoUT7
vpoxPYA7VjdVExNZSgJ8oDJpWSDQglBqAm9chbvDcIfJ0lWA50pKhqjRuB108cPpM/o2x6vFEu9r
fGhQ9vinr8QL11kIuPdcXX8e3S9V5XIG3C+hTNT0O6LxR5b9xk33BGCqPrLCZkwVwK0B6ZZzJ5p3
O8IFpzIcMmHaCYk9zwuK9ptJ8MYl1oGgBDw2EsY6F8mFCpgkqC1R9ayFwjcG39Cd7lAz3avlcirg
xZx/RMU8bW6KGOI6YOYe7J5yfGvcjLa/VHWg21FOXf75UN3pFJZvlKrmaZUQSgH9Iv8jLofQ4v5f
JQzTPUId3cBHDkIcqzZcLMhkdt4H5bfSopzVniu3kVhJBQOznsRAYAAoWYP5C2B7aSykK/Q5PqTL
q3qi7cy80zxpCQOWYHr0TEXHwg4jTMtqLuGCGQ4bDSxVw/9zRiPMqM5seLfa7mdMcJ6859eddvtg
u7SrQMlu283pbtnDy9qO9X+WOdw+M4EzR2mQjrxqwMNwx63fu85Ycgm0lnDui27U7DqYWBpbdxJm
4pcsz4b3nvhrlRmxUQva7e6rNIjtb0Zwgh9OPkPyT5/M8WbxO6lQY6lGogaKIZQmPvmRBwCm9KIU
HeIyWnQEPT9mhrKxmc2Ero0HUxWo+fkjc6+rt7OTQdoH60KwTpluZjRYPm7NEN0fHvU0BXgyYCKp
sKj1h0kYU+JLFUMHCPt8EAEcxZIKAx57I3cRUr9JLn6VReZaTAR3C/JAZTS397lfauhsBRdP8OGy
C67Gufq8aGny2VMcTL/6XkT3K6eB31py1uc2sCyJuDMA8Tc8Nc68OaSf3NLobClYUv3fZjrps6Es
OvjCOCHZUEJaltJEc1uieI/wilepYcohEHusfSFdrYphMNAOWaYoPI+ymZ7Cj5QDLrd0nV3sHBDy
ROZhhAZIaIDL5qt/xOBLjXBInme7Izci0mc1J0Fq2RajNiFIV5rgI9YH5B1MWAdU6pzPcmZBKV69
2PhOVvN4jyNma2i3MfHvQ4te/ITdL/0uoDuNc+0HDmHd1GavT4/Kuu9FTpSZk/FcM/mege5gvB/8
hdKw8vEbu7bAgXq07XgpWBmgow4yaP1gVLOqg8IfAr5uhYK00G1NAS2bJyxFV1/wKKtW47JC8f1X
1tHsZ9R/9IPdV/AOd6BM8iDM9wRnnI3WkYRFuysvQKm1HkpAGxrKIEC5wW5TYZfsNw6Q9hzov9Mq
FLaY1yZk3fydmIFYqDfDh0hNoQxfHjut332MBToFz9qbLPEEw7ZXTNdaQsluKXPz5b038qMYHhj7
Gu4j/WuI5UUaszyksfcmZ8kWQm/FvrcwnQNnVoGOpjpVtoJiNtf8UPahPf/Xk6cBbV34fc6xQKlX
knCSj29M/XtP1ZKBVfiXm3KItB0cxfSebjux8EpmEWNO8NU8q7xviKTzxH+zFoc1RRMVaDS6nHoG
si8qNmk+x56sa+5wHy8S5a7E1qORWhnOvCTp6tQN3tg7DbbZhiUQWlJESmXYyx2TAjYKsJZv98Rf
bW6uRAKXtm2AETWOPHVJDVFMjuWk/FOYCvGhkf9Xfb302GqDR8tHBeIgCoWBMKUwUK4xW/5wGaeY
VsTPHqMRqSlYs75XGmbA4CV/LZEnvZHs7H1eFozzixrJdo+I2XLuy2oPowIE8L3gMh1AmX0io9I8
glyC6pWd+dkZDi7A53KCzawVcOIhVWdxHh4j6gjoVPonsU6fXcZ+FqjvScu4TUtioncYRymc/yq1
paOK/2Yb/CjjS7PzrQUBh+w2dzB1V3D3DS28kRvXpfq4yEPVtoamyhP2mUPuFguW9HwPd1KDKXDu
yU3MnVFxQHvrjntuWoQxCsoglhsYQX+ai4A7HvZyiJV6VdePu0onS9A6QsN2fnQdn/Fg4Rs50x5n
B9L37seZ8XYD4ywwThzqygeW6yHyOuPqOzmS1y4V3ix4oBy0XqiS7OwTWLSMWdcZsJi1pVhQvFsz
429u61+n+lW0WMDvkAsDh8VX36e7TNUAExoZL0vTlSFTSDpahSi5URQ1vQq9S3pB3PkgOkIITUEg
cnouxdtfLNsA3CJA8+Xu1E6tbUQlMPpVJL95GpygUo01g2/xzeevY44NLRCnARtymLlQEhsaNhAJ
QSQwiZf13Jtn5bOprHImv/3uqXEyG0gZTQF9aefRPJG/iAKLt45xAuEb2FL01cWYiWgwYokxzmob
pj2BQCxN41K24x9JHUUEZ6dT/2Q/cFAczTrgZyuBxLwN7Wfb7U9k4I/08ZonlpYcUIC6yATw0jyv
O6/E9RnSe0tXUXhUmpNWrPwkep5RP4kAUHz3wwoQneunkFnfPR8jGI8PTV2CArCmQnEbb3XBILA1
mFWkeOhB3l15ep/SsOlho9aPvYzzTy4Vbm44Rp7EyUH9Ge1ASDWHT5Xkr7Bx46LI/vx33hfPi0fL
4UhEaH5h4zyIbfdissOi+eAlmv91PLkGMLnMXVtOqKJTihuh43Vzg+6MH8O72v6lLWQarF2e+fIY
WXzw8U+dtrnT73hPUKNRO5O0Is4jo+egtuCpBA9kccawH04+J5F99MpXNl9y0Ne3nT76KuULfhDZ
reZY3mF3vHDEgAKLVxhOJXZKsV3LD444XqJ2y7ebQ4DSJPsnVS1/RBKPHsoCb6kVuYZdSPC7tMsh
INPDQluHk/X4cobsAU0s3g1hUFrkMfImUxDXnr5nxf+5siId9E+uKgBKvqBSiwOvMaM67tlTwG7Q
mn7yPWgnmiPw13lfsJvSXEQuOJ6qX/6y2k/fMecySKN10CPjaKv52jt6OLJ/F5uhaNY9Ty1MnpUJ
ez0sHsPfE+WCRk8jeDjPuWrtlyBsui1OY2QmVpq2h/IoywBX5Qtn7Gckv++O8HSQKnCQ5PyYZYc4
qGN+fj9hjJfIz3Ny6xMJaj7CyYFvTA1pRCS3SxT6rO+p5XXlhfyQI2Vt60eCuQZ5m7PupZ6Z06xP
QSKiBSFfJ7DQauCFBHr4JB8J4dj3R//tBFVRlWsiK2A8NTzTIRCw3jl6FV75HI1HiwaMPHwYWB4r
cBTmECTHlqPzq7wDr0IFe+ecwK4+hxOd2QZBvirzuu37B8RwudJ0hD4RJCnbnvsaPHbeq/Kyq2HM
EauCQ7nmNcKe2gL1A1dIjJTMzdB80Y115/3A2taRhkZ45AZ0Kf/mdJmEUutczbOckUVICKw9fW27
zLCNPbcFgVZaP+SHZJb5OskAO217uirWyzRXdLDxHc3odB+XPE9rsiaHFIgrvnwKVwQoa42PzmQ9
WdiVnaHcM8MNqWOLoluNXx45P1kaqCd1taSWiOVZvkXntyHNtm1lOqQ47Flb0rcXQsleVZt5r9F3
l8quyZohMwRASol5wNJS9oDZRl/lAzIFhN9vrL1MNTHGPf8fwFmgDL5NfjYYmbxDqAKmWV49YAPw
P/8uoIITN56XcbaELYZ2fp5LPoEyHhn5XfxtbnUwqx8YIZ/vIarGRLIEQBIXabIWIDlnmZEAKmw5
gHU7sxzUMicQWaN3DryePYUjp+qjPKSthWaKmb+c+FJctHMlzQ7WS0YUSpoNjG5fpsmaqBvnXkeT
+nVnyMjjrs87fq/SdzvHNwekA4CJ5Ew9ilOV2b45kVxOOJBQkso1PYNrX5PxnbDd2Qt9ALMddkj0
xI5Cf8wOM6Qe9nt7mogAVi96622CS9ROO6WS4TBSmRsypFtTIZZlxI0BodFBsHnQ4VXoGR9/P4fo
EyC4bQziedDp7qhhiyQ6E3tk6j1tFTPPoFnOdB04WhQ+7PiSN+Fj0r0WwXHo/m8iJ//rH2fnUs4V
g9Ghq5z/7VB8Dl4/yn91JG9Zoc3MzizsPGLGIN4n8f89+qrbpQrlJXyaBD1OVhAM5RSSWXcVdLSn
0veyWe++o1EIqMRO5sLVJtr5TtVpImXVdyT73NzogdvgCyIHt6wEQicmourK8y89BVGyeklMxsT/
4cRaL5uAHfHxCKwh8w49iZZYWT9Mpw6rPbFZrU1FJYVolmrRHQ2qn5tetkXAjv23jhIzN8Ex69KE
0ZRQPWcgTfssgfHW2fdUfO3VwHZfQ/OyTh1Txv06w2//BRUpjHfsnUkbROOzcUfZR+1tWAujb9ux
RqjXMJPxQym1YM1DMfStW8x3BKsO8hM0zeS4rJEbSxBA9Rt7V5kHEKCkmzwaPlgf6iTufxQzCSa3
IXgzpW338YWggLLOcXNTF/bVY0yOzewouDoxkfuZBBeCRQNeHIBpT+Yfzh8XLn/shgVBAx0nflMQ
2lbEhngI2HRj455vy47aeT38OrDCeJ1nnVTSspT5SS9C9pEtFgPle4xYxwaWxU3h3oW/xmVq3fE3
GxStaKUUqrTuFKfcuzi6KGcM/yDo4zK9a7TPEufbKhAdwMBMXZOtNxiybDYhpRCIRfj6coEiWcb9
JYIhYi8YaF7T+Y8yJXvkEfY/Kl9zqL0Wd2oDSo6Myv/x6LP19o3934hdfPqaFdqGnc2sNCsT0LC7
kGitFhkTax52LH4vYFCjSzWEZBVKipzQemHb2BzzCGfgpB4bdsxOfWGWN6sDsn9doA8Bfz51w5tX
TbqJvtm5Kh/U9fT1vyye4qsmslfI/SKu40CVGmHjUu4hlmOODsO2hl/MBOAKwiAg5bOZUjnrWELH
knIdHkMibPxo9+T8Ft5HQ3A9+A4TweAqJQLimyXmUYhicb38hiyz6PgDSY7tgcyQ0ipq5o5KktrE
e0kHw7SdrNqGbxJM3BXjkl/n+bjgU/cm3YNXPSIblwmCebHZFCaH7q0wezMDNK/c45Sot3cZHkqP
kOALy41E8R/e8dBBezQKLiCrPMSYIjfUYvdmKx5ImLJ5mlrCzuY/Gl0V6C9zEgvjir5IECAA2ocR
qNQg1Bj9FM7EReuwuVUSebNd02LEdp+inKi0egYGFunFLRBV8lOz6vbCyYKzId4hTLAo5ZcBdZC/
a+fXpISZ4u+RELKVm8rVetZWvmf9RZ1Nt8RQlzPIRSfXt8Cc2QMsIORG4dSnKxtyGWTlR+BUKUMV
+bPEbosUfynUG2keI4zoVya9nBJFie9M2PBzTv0zsv0Xzaza+If+WeQSvMjD1WAw1n7HiYmo1x7x
XWkMEn7/cAvA4/WT7FOoYcH7mO33lBAVH9mYpJfVe3tushsQ903AAsF0snkPzruy+J7TJ3W4LzoG
e9Y5472DtBOO8G960PxXmAH5iBJwvPv/1KYr2SfFSdO+Al2Ratk3yFXIPQ9fbIpn1BjzlSnF2Gk/
olcDnSMcgb4GyI+A5eRgI2ea+20lrYhs4436V6dzsVIziqoknDYLSFLO4yHR17chIFVZ+YDViZaS
SOVPcnSU6Y2M80qBly2YAgZYmbNxdSWiS5giRyX/FA4mXEMeFY5mdE95BgXpPOkRq99xoIymZwfQ
wA9rpcHrIgrncnUCDR98bsn65COlWL1GZEGZKKBYE/eL4OQNaF24eKlNjsbwNUhDFtxDPrFG2kb4
b61Yp/jhEZTCnWlBWkzWts3go96Mf9dK7dHeUsaHM3yzOXbtnOIOlfjaVIVnRYsnIbAOe+jPJsBu
bDYIe3JbRvA1FGchGHW+PM6TF+4bMEdGdcRvdin0hL2ejf6bcVvE/mZ0ttP9YGmFzFbS0bw47WcS
o7a9hRozljV19k4ANnlRkwdiRkp2RrtiDIO1zGsngi07EgqwocBS2EPt+BNiR2oHFadlIsA+gsJj
SMKct+SBXfMrVIirhj5VNZN4mFc2BV3OtWJMETm+XXV/8kMeTU+9c5uVTRVvUQUvlJrd5TxGzWKi
Oa0FXVJ+OAcBdJEj23QjhDyZBPqbTwrVXRBklqz1Zx9S3UCLZub16gF+dbU79eh+uFrp0i7zsnNo
O7P2+LIOB/szOfd332W92DGDWa4L0dvCT4QuJWZmUlL90MAp8X1jyBkQ9S9tmH4gq1agAvYelj/D
pETk3Ddf/wSZNMtCd2390E+8PDZCqXPLq6kiIEMngQjSBeXy4pJySoB2UQZSzD09ZXnfwJ/cyJ+C
84cmxeiOnc1EdtbdFaIlFfwHKJ4FI1fknaFd+I06xRJ3mcIYK1ONilxHXEfJppn0ZAhqA58X3cJl
OTwbNigfBJlMdDAvmZfkJ8ccqEfs8AzQH+KFQrPDbv7AIfZUPFQ5sfgSJojor8lSvQhCCqGNcQLn
JkPoQObWwz/iwBdE54tslJvW+cCb1xshYR8sWFKcSvyN+On/QG0qa/1RtijTlBk8f47o0h7OJoR6
XeS9f6CfOzkb6uxCaR2euUMFHdLQZW/VjO1SBkleQ/AT5EjJB6DK+YGA3kJV14dF9okluC+0PlVp
BH0mAsH0IYhVxqPsOenqcNUDM0tSqZ1NO8oNLeJq8qkJ9TwNrX46+Mf2r25ZsOM+0y1DKIFCFBcL
H6b94IzO3+WXT6/5oZfvsgeU5KcK1ChA7IRtRvEVfxymMLUepms430ykPwnemdMA4Ozw6AOeM49J
1f+NTqSkoOpUjaplgTIRIQAIw6BUKAHSiR8FoVlKf8eEpWGndd7D54aZ+fqi7x0TUKUTpcV40HeE
Wq+H+GsSsDYhcRy3vQg1KZgGs3BcqBD9M8dNHTx5KRIiQqsGR94UGL6vH6tFRIAyGsh3JT+k+RoC
mr1Sm3UH2WHx/pJpIRQ8B73/rkCpMeADAUmTUkVsjbKl+mxGCBteVJcO3+Sq+mGqDIjo9PNSzRlf
BSouShmxyRe9uoFLQm8a5ZhZM6+H9Cxl3KDe/4qpA5oLtKhGxHHp8Ik+1m4NAHKkggHY+W/3St3g
4zPH0VJfpZk+DwkT3px1vS23/+b9WcD6WciV2DQamJDOcEVBze/Lla8BbKGoWgPeGeugHBYJ5QQ1
DElqyvc5nNR1EtiU3fVE4+SY0omt562I+ikOMf1pFDvFPy8ccIqABQ/pmSwKkH+86D9XVr/vnSi0
pVndrxCh6L7FAfbz62/VnVRklfh93yhXSzstEdFF8KnLO0/t6yXDty74Q4oHqQBHvZWzBM0+7qoa
D7WyBzZ7qdmzzx4+NTxwdJZrLb+pNBmM3f+Y4blUwkoPojrWPXq8Dj60a8NC68kFfPEOHmkXRs2I
WL4FEs/3GPjKnyUciCk0jwOEBTSNLnRDFuzRef2TsEphk5YOJj4fWKY4AGRgVH9bthk/puMDU//0
KJPoAbVnBMSHd9BA6sRsakc254rte52H5dhXE/llw2NNKP9Xf1VG005yiW1UfjBlwuIebK1TLwbZ
MlOcQtzXzsE004vUo1kY3mG/x3A7ClbH2smwcc3B+D0XbPYK+7ir5zGPpPBuxBtGFGBmdXkzYXV5
UN0N4OfS4S0TLu7KDKITdoTpKkQr9/ZOezTpWRfWEoeTo7HFmo6LukqVpnvxEB+bUJ+LxJbRO01W
8QC+6q02d5ghpgslC5IO4shhFELm1ZPkOjTxarwjPxsE0cihqi6euCQqTZKUDHWWZZ+TGNmd1+n1
pzJt6Lq5OK4nB0gbuBvgeBvwnV0tt2xZb5dXZ273A4vj/vRxWJAan5BaLEyOH7hk7OtykfXbfTDD
m7EU85lDwpf9qJoVSPnp/xFuQhsslkuJp9LKOTrqGdDl1NRYxOJVpry0SkMpCYb2ZG0nycbjIQqD
uqxZ+rSP4aWmZax+cHEbhM0EfLmRpQ9dTPuQOUuEjrWZnaAl4NFR8FmKfcmP6nzB9mp1r+a4ne+/
1UFzTYz7krIj/Zv3jYeAZ5w+vasEyJWMGYuCoNZvd6h0+Yp2MZCXNKubc0+nVY4PpRdgq1lwGXze
6ldDdChIiy8VWSMO/ZN72vIx5YepzZysxBAEfs71TVRY8AZEvoIOMcnHhpz8jp+V6YWjCrWjHUj1
GE2ZiIXvgIyLWjaUc5AFE7Py1FQxGtYNdR/pxPFkIKxGXxndSyby/k2VJxxZGYcLY7Hch76XAd4Z
9fD9xIL5zDyCJvVS1ZDNRz1qhQwOfXJZ70cvF4qJD9K6IiKNx9VePQYon+AFk4gsZr+uYTtNzamD
V3wTc/7q0IMQ/Vy1gOScm/NdUDLIqCyY/x9bhOo3jD2z+lFUkBxr1SitvrDzYfXOaCiXaaa06Yko
hfyYibdjDvmDr52/gB5CMlNAS/6YjCLO0OqO5zohJjw5dCq34wf5N1q0qtaegcg+6VNj7oVOfiC+
IQ+S4PjdnPa/IB8HTMQLYpYnta8E2k3rqkUsYTNEC1I6hTamimHzjL2t2Yq24V1vTjQzL9ZCmF/I
5WiqSXdFbbo/TbvLt5vW4hdx2zJtPh1S3B6tyrKLtXOtnPcuDXkSvRBL74pZ84ry6Tf8ORIY0mgY
NuNGu+mhGTSQeGCmudzJXJpBEdeg5qzk2/uLGgg6PYYX/UwC97VAST64VGkdMm8XBsv5E7TXvzn7
G2CCzV7I/b5VkTywccl7YYqgzc1A+EcYSHn/g2dsHUpIzDzdWafs7MJek2o37kez+a4utfTEr08x
TGEnxTIXQRgcLspJ8JGsfCj8dnwxQsmpVYD2eFQpAWz5yFFmP6HDThJmV8hZmcwdsbR+V5Hw42Th
FtlS5Cp0UZQ0JNyu1QKYc789DbjcI4gm4DIX/TnWeDjArU9UjFCxKJ7NTaySTOzKpNcxXyBqd7LO
BRg2qa7iWCs2qb+5Qm4rh4+1ZBarnhCriYd9Hsnd2fE706+w7dcqPj7rqu/JdodBCo2Ef/YznYt6
HXRWTZSIVEEkwBQnAArGoDYFVTtev3aTikiI1yXqRv2lIWcnpQwuMqVcdgWQOcKk1wDFoEwPzCzz
heJDBYHEunFbRJSi01sXmKt7aeJEycr8FaLKNLlWFDr7qAnySEODa6IV2WfjIuG1tQIXqwy2LnOk
R2OI7A4sh89+b0aQ/DmMdhPHSElBYul0VqSPDUi/RPwL46P+97DvEFcZsQ9IeZat66GZomYyB1im
mV/wfOkcsviIEyzEBTcocv5DG3OlSsl646qMm3pHmG8e4YZVjc/RfB4iTZm4fb24joCH9TFMkRyR
DpJ0GlZW82eyy2r14wrth0gMK8ejbGo9jVURoCl3l9alIM5HJu9iJ/m8v4XvF3+KkngwRrvkJj+w
U5y7MuzSA2aJ21fcHFyPd0wOPY24P6soIwgR2ssY7ljWA24OO2qgSjRVEvpTriEXlg4n412zYO+F
TEabsJkT0M+JAkK+MQBSOyWPdkbwlkJoG/DjaCtHn80SFR0fH39Iyx3tb79BVHN18vyVQwo61X6P
R0z5Ev+FkfQEJNfBNelPNqpIkeQ1ixzrPZuEvvrunMI/8CdJzYcfZKrGcNIDlUR6v2T40X82ZQGm
wodKKY4YVS+q+QLkuoVQAqAf9GtFLZiuXsP3aKhMwFj/Qptzc8rcC9+QJqLhhH0qvOukPdi6u9WY
dchnRAhIZOhwAnHALsKXe038CEGpWeBJeLp98Dmrg/uYbzb2jxdNVMHE6EW6gc7Mkknel1lBV/LL
I2B+ZA2tWA+0ev0O08e6bL/erM7sgSa8uGl8UfkqpWGvgKyevlAUh9bLJQwpmYWGD80co696xnkM
YXOY2SzlaJDpHreCmU8sgdSkaP6XbPcz8DexW5t+91KedUPhrqo8PyP8S37YE0DI5Bv+A17wMV01
rsojl7tCZWwXZBXB2f3k8dG1lz4a4YC2PDlgKkHlgRy2+d28y+T4vQZi6aNm7QNaT0szMDjVwf/Q
eYw+qw/3tfMguouN2DriWpw5it5K7Je6eteJfKE4OQcS1kdV7aVyeEE//8TjVv1nnmnt1tAxj8/o
oDJmRMG0WeYVcwD9NjX7wD/Jqxt2U/agI6VnIp8itCUyCOgJKajnZW1q0iAOq1n7b3a0KD9/2eXJ
63f+v8eHFxP/SytfbyHuyfgUxvfkSz7qk2x8xiV5BgZkze6Ik2QmSSqmMuVWcseOT9l7iM3mH3F6
d/YUE41HOFXG6al/t527XWIr0g08c/wqNIpNe9168No0vTAVaz+YmFmhFovPKHgIcWXZ8nAcBlCM
hKfonfOWJOKRhyJdnoz7M4exvyxcPPj6jn2nK6Wa2DpZKo05NAv6OsHrUbj3v+/HmIWRl8qDD3IC
AF8irnVDjGI3ILPa9rU+YS248Y7iqEuLz5TPL3ssizkLdaXwVXGWuAHUt1QZDyt6exvyW9cPIhJG
G4RpbNUpIo9wQnk3qPh0I+OBIqyEtmwzz3JTjo2USeP8XeY3OzfZaiGcqM0mHiNfj8VuKXBSt6Dn
5VIFdfHsegwpYGy8fH2EQJWOuMnU1N7LD3y6BRdzlAs1RKKK5UAlewBeM+lwPa9nMP+a0xhN5NKd
TUNwhzmfCxR2U22aR9llMghgU2GCVE/iHIW8tI/MV7xeHhbSPpqI0AQKNqRhr0mLgq8dVSzC9KTL
aeTxfykXGCWkQbLueI4qkevNuZKbSo4qGNDi1QBPS1kW5IIl2Ph+KXSwfGI48ZbfRddetuqNKUNs
j8m8ArXk3P7/t8dVHI/5k1lhUDNmHx2im5DMAbCuGCR0Q1zHHV9d2JG6xGoTsuBA/KbaYBP+/RLa
4jjKUBF47V+cFmkjITfCHu1i/9qIbYuPtcb3z+aXQ3RkjtoNm5BRIKOdVl9HyUhmd37OxsuKML/G
WYC4J/DybB37qQDMjtKX/suRL2I7fh+z7njYp3JrgJkU2tu7VT+1s30T9O24Ish6L1aAAkipdFvV
UXyPn+dFc+B57D+/i1go7VCODPLAhkH3MIhZJusxXedfqqgVn0Rhlgxu49NkZ3P1Ag1k0dIPnZJ2
v0X+qYRYPDHDnoG4PGcpgOkisxMJhfMGCZg1xCfUwyjg6yljtu4qIh45Yq/MXiCw5jnavMHU0d52
Ypv3dELzeF0d2kON7UQGHqIknZQdibLS3+IOC9wXr/Nw6+IJc5O8RcH3iLu/beTZWJn53gpivYN7
U5rz4QUzTQzmz6SzbJgATx/RIzEpM2XmpxEP1pUm0PLh5CxRzhVrgLPtEavj1JGKEeaoFVnqB3rO
ANXFAlXTygY2GE00LjLYlFmurk748FhAWUkzu/BNykUAJCWKssosit+UfomPIhdSUMnAUf0m5qdu
7o0pshXXwOqkY6UaS7Szg79BLUyjs9Vfeo1qYUA0sQ7zNx0IP3w3tnyge9XZ/wmspok3JWfv54qm
noUP/9YhGaeoH3cPaYyrDrbIU7XUWI0xHrY+KC8/jA3fYPzOY895++KQpS4G0IdJ8iKuNTbFtt6a
OxMv69HAsfbeo1HDUdD/8jlR6/j0xQ2gktqx/jFUzCDvbtrc/Bhgm46yjA0T5H3MTH/0/G0KhIAx
YhOptpvClk4V5rq9skkUocT66imFvmH/4556zSEVLWGmWdjtEPuZUGso97EnQpvFenRi8ZQgXGin
k/NBUzHlPvjJx+9zEebO9gstzZEd09C98S0SHRamvXslPGZ2Bj7G8MTgDBxfi302B8PyvApSPS92
XxZeJZwJv82J7d4oc03RyHX4moogcEuNVMT0HKexXuSzmjNvGkW+M4qJvKnykt9I4P9KRh4ZMTKd
z7FaCAgSxAhky7l5US9CfxGZwYqXQsSTs9O2sj2vVgrVsGbw/Ix3R5OzWnTU8DCbNAgyRqvfsYjh
hu7ByvprjdGN2SDGzd2K8GPNV4r/0qDqtwME6R1lyd2PsaZ8gKIsosCn2USSG33Dy9tLl12Nkxp9
rBXmadfZcW0sKVkqxYTdsjv8QCv5GR4J11Zj+0oI+C3lhXfW6QjhYuMj7OMPYnOGUl4V0FqZTAXo
or6jYLk75G+3pkTr2Xl5pQwVznI0hQMYAf0gfhPFjIzLKD2SajpuxrmHJzU3QZap0M/mTDJIWFJI
bxkSyqAKet5v6V0WpuIsoSpJVmoS5hNwh4T6A//Eouu7Fv7Hj1tXd9hrDtmok6XqigUJzfOe8ieE
ZFeZP5m90VN/NA5pAcskuldDlaaCAG7P05ekfazXlj3M7rd4yPKIrdn9H8/PlvNqv61csTIZySU7
QaEv5quyhXTuUop3RJD5X4B/yhRvxdniNhDq2n36i+CYbuFW6C9vLswXGIG0O7B8tIoTVUhOgqt1
dsNx322xyblWOHDtwlr6hcT3tn06UxPWJLrYaqzHBrQ3xmgH/OHPX3Ee3tLoDD+mvNjHR8e3KGq3
kfCA0BYJDjP0mxRlrfBIlaXXNVA2toDE+X+t6aKmT4p6adEalQ1yT2EoK6P+cGYRyBXvVldX7AVW
rNUnGDoRrq3Ca1ozHqqvGfwxIDkYuVOYup1vH80bokGf5vbG+uF6gDnGGZHe74G0MRRgBbd5S9cp
ls03D6duEEq8ME/jUu23Ksywga4BqttD7PoeeMrzjuFMRrOCzOxOJe72N3lFmG2xzV/izoAbF9Hz
mz7HvDLHpIHBh1jeQ5yeLntarUM4xfmjxFHhKu7j0dPxCnQ5XllPoHsH2DfryvFwNw8rxI3Oe7hx
6Ne3i/nY33x4TYoTPvBTWFVyx/2lksEoM7e4CgKuWh+8rrY01YgU2NjeiBTf9/IoKeCqLVS7Muo4
KUkk0nThMsc2ACePiFpo/S4FDIopPYXQXWsKluErTGctELomlDrFkNLrco+CvmUzS8HxN1uFTYJF
iRZ+8hspQvXS9VPnf48RRTE3mpOjGHnsSYBz9EQh7lzrTSUs6Ce9PHzbG52/hZEJfUpFqgqDh2Ko
1t7JFApaAqdkFDZlUp/WSWiqyRByp60dL44pNcTdWdhFqtUlQLXlY/I5OrNj3xi6ypRTIxLjbBbn
upnnkuUJ1DKSnMYgqsWN0usAMovsrTAGYrSxbFtquMtzgVyz8mTvMhK35+ZbihptIJd6eEhBaJWB
+P10lQXJd3zjFUrKBVQhQ6QMwAc9yFEIC/jKW5oCsZHdp3ArWOvtgSUA44x2esIoK5LXGFMNAvxM
EDQc4ILr26dI9Xi33kE0DHBd+RuO7kIsKigACe68H/VR0FLnqhYn49kMukBKEu+hZtyw2iw809YR
DB1KYFx8D6w7FruEq6o54oXqkfR+bXMCZjapX4jipPi8qkFAQETiWoSgmSfgfZIKzV49TOc7cjHG
hd/6RgNxOhPg2ypPqE6ceyeP0cBUisfgYCHHeMDjgp0btO+1dhxCHCzmaMHNr1iZi1jy4H01n9cf
XCFi4venqGThk361YVTSBArBBG4LHXAjQJNQV7nB5tPFlUtzp6EL61YkWkQetb9revOSFSVSJxWn
5H0//Xl7S0nh7M9uVmoDJQkiZKt663CCiJ0KmryuYnimJO1v5gmOQFjq58x3xhp+NarKKPSSjHgM
2l761QdJMrPjxXiHe+NH6n1KkdXkgut0T0MmjLhO6ILNP9WLtcyG5/6dd+hQrlTmsujTBDLK60ZP
7FH9l/YgcSJj63es4LKH7bOL/HykmBFw4t59SST6ynYA6giDs5IlcQZAHhyKhp5HImMe0wWx2/QD
fcT/wVuC1gwH5wlsjhIX0rspxvFSYaUdxsgqAJn+PwZPss48iP8fh8Qflygc2WzgdULtdXitxpVL
FbP/58UbpBngOvgHs+P+8fZIJDT1RO2yl8BlHa8pAXniyz59IjianT2HA0fOKhp1m5RgfmSNfkuB
IOifsO5CGvv7XZcJQvtW07hBNrXepYAd3EXi1uA29y+jQBjXkfUHcVkVkQmbi/rt6XClNmL8u20O
knQsR58wEMs91YHwmmZFzzxWxQgLEeHVFS5jsTjqQ/U4z4wI0luBE5mVyjTj1rjElRmF9+l4NHrO
bEnlJu8MjUm1D+XAE9T2O5w3cHHyJNY6/tJkcO+Ptjeb6UIIofTnHVr9IppnpRskcJJX4ZHkGp/V
zHdHhCFvQnvNlj+QuS067y1gc/Fy1s/vkDXuFth1/jComQVJ9G25JFK9/mPpBBQDyUx4VeLpDkeU
mN5X0Q8pOWbc9vcFjM9DawvFARgVg9HNeDyv8IHzEsqCqpm+GtrVqvcSjsOiOKD3q9irdrIGng7X
1EkTdNpnUU/Bv/0vpF7iNbNv3cqxBumZr25NZrOjrklnijcm4fMt7dfvpOSDaJEMAErSrJ6qlnof
uYzm+83Tecwzj38kbEZ5L4uRSRba8cPh7gXGYxslFjZhfjhYtDz2MnDZT4SJRIYNG489/9B0a189
PpLdB2tQBIDfmHPwPujRaBz3Iy+16LOBenMb+hP+vFyKJZ+IodL+5ILrz6ahpk0xMpyqVo83MnCC
3AWR0nVFnW3xBRZblvZAoRmTFrZnTDAIsDXbGRYrd7l4id9UiEzi9IH2ESn48aux6yPbnOukNhYk
+hnqiWEo4ektvC58k852DYVatp1bMx+/wbYWDoZr5wDI0TmT8jH3kYjmVKn0FNTCf4jOTa67FEvW
Kd33SkPPByFwCvvWHx7Red9C46nDh1JawBQc+7V4RCazGFFcvxby2mqdIGTin8zLIioQK4Kjpo3b
wEfTFDoYKTEwlcV643a6B1s3Dpy1cKIfRijsRv2koQEmPIogLG94GH2LgMKmgnLrFIhaUMiSSL1X
s69o0yuuCwbevxrn9lYymuK27T5qNMg8NbQFaPZEbjEXK9ZADqA/clTHXQ/E8knxK5PWMpJZvsfY
Ymay4G1/XncsIxcd3mqYG3utdQ+RCGMS5IZ3JjPMRpcA7CPo0kyAQKmaMI5l5jRO75Wkl0eo8KXD
+RNbFoGokJnuAQF4VMR4FEKaLBenGOSkbqs8j0UneV8Mf3fAyRWeRJmp5e79oZrwopqzVySKCjnK
G2nbw2zJWTuRR7qShqabN6F9/nkJje9n5e9BlsOolGWFxLgwDBx42Id1pjfy9czMBwE9aqHLpvu1
IVLmJM9UXNG+S0+3h5fBHV9zaDboWor7Dt77BtI5m8oGC0MsfMSWCqByl6Adzk9GWAEf8ZJ6Mbim
mpgpDP8RlEUHIo9HJ/kJ4u6bUZCh1kdtzgzfISrkyqhaHc9Uy0qXA4we9Oy2NZOPdluSHF/2ip07
i/2nP6D8+XZc6HJnOnDFiY8RpRz0VwJ2kBEtZFWgJ0xvnwcoYoXZ7w/kKc+CwBWWpri5meHkAylk
6z4WVUvUZr4/pjJBSrv05SZS3/LMory2+WYOZsnScWsQXeiG4WVib6BPlSk670W+lMcGKCZmToj6
XNMW/PPpAF7jTNz7WzLfBSFZZCmmKQEa9hGU1Ex3jIKbifqf7Mw4mp8jSlPMvMwG9SK2lBcEg24H
GdngUIVG0dYb8FOjGu3UJcdBlFb6F8L+TVfzafFd/TiDVLvgbj+U3ASOfObvea0GrRwdnC3mm3r9
77eQX2GndUFxGnAMc+pda89bBsAvT8b5XjL6A7hXsta77P/DA3Isuo29Nd9BAXkjognn4UJtQrNO
TSFMwNsJw5jp1G1Nt1QQqXbXzod2UshqoBdFFizoH/wOWlSEefiJ6vXhmDeSa2D0jCMWtuP1b2DT
vAP4hbV/d5MQdD4x3Cd33vM3t9w8iIGz3ILXQndg9LPlgzRYmq8173NwYghO3eJ2wkywnHM3UK1a
U5AhfOF8ia6Tf/HIMFlw2f/S8k8z0PMOXjqIw3gb+SnJBqQCe8qLgAKQi5kY/Wmci9ygEPPpNMa/
Og1kLBSjYbnwnDmJzWVZL6fbGC2Pqw8pgWlDPpY716B4uKD+Fjwe4m4ebZE4QRlsNbnd2sFIwJAO
qIqDsCCwB3pv7u5MFPYWwOuZXMT/Am1vCTK2rjdjqdspqqtA82BQKldtbB6op/KP0YqecoY9zRQN
GAD+AfMP9NOsO7mCTvOXv9RpmFcxaxKhWfv+uPgR0XPM4oxj06G0Ka7HFpdUvKA4au456iYPDK9n
VCsghdh5hCqjEobqQ05Ya67JdNG1at1+K9V9obptNaDWwbuTsbrNRIjLnoz7Xgi1AtW4nIRY4tp8
IlGWfd2Ou7TTEuoIjG+3rvtyTUPonELQzk5qVL5Tmfi72/KgHXxIiAbTZ87KN8NTIyXAlkF9T0cL
EJffoosSTej8AKLG248gh8kIwFdfe/5r6rwK3z2MEQC6onje0YLYBmBvNO0BUTtwzHSOwGXyXJs8
LFFQU3y7YYi5b3ukzTAziKqSc7m++xJ6c4mIYJfq1cEn1a0hCXpq+9PctOLbWAsp3o3TrVUnrBlW
IcH7BrqC26TpAtnoIJubE2o75CiOpi6bep6zlKFkQmT5hLdgI9Or8bL037oBRX0ruM0rWleUA3bu
oRJZB7BOhKoWp6Kh1tYEndcjfQgB+9jquhzXSjAgkz4ghjOL2HYFa5QFMePx0VBUWxGfJ1YOvSyP
+a3T2d3/RuZJq0OSPLYT7XpwYCDoFzeEIV3yAlnOIV6EmHFhl4On5oomrxKZeKmb+N+2NFvvCc9u
I5gDsvwoW0Vbar0d76q7qb0Yjxk8d6bxtPdaFTBEp1SpFwh2ukPAutRWT12GQeHaUsL6VztJy6L8
mUOn80JIPDKzkjugon64l7YWLVhkJLgKV6iF8j6+h9/eufHu5ZNg+FtD1VrFANWc6QHmBmRBSt/P
McNTVyT4ToPa+QnK40vn5bTumuL5+wTBvAPQsLMMTdJSqs3R+r4XTgtsWgKM7fsZ3AM+BshXcDFF
fHY8IX/+k3aJEz1dilenUhPKC3gvCvXQnRPwmZkQP1JvGgT6gaBLX3GHzYGI34PXDJ2LnmMCEZRb
c6gltoEKK1B1bKYYnh8iHaPVFdYkHw5XN4NLhN7rskIF0ej0/RXfHkZ6A0TIR86eHdwsJPLEkh0k
1hsfwYr1pA2oH5zYI1bGBqk2Ghatj21GnZzJW/7xHPZUoHrfjs8fzUH67yrbqPNn8j/3TnnYHBIZ
72TDS43j62Zp8FRXW3FzBLqlVAzIEJQmbY3vJbSQVrXGbbfFpusfYqDTC9FTr2YNum6NDo6LigjQ
p+A2LVreQ2pDxbzcOOk3PSVVB2dMoUPvpqTSOa/YfkwIEXb2X/jkFpYwr6tGDqJnpc5DzBiet7Vx
ytVTIK+RvrY7+cYBYC3cvnO9pwWP/FQc+C6jRkbQcI6NMuPvlrJXABvtIfnvGFh3uxbWKWs91Qeu
mZBUA0gu0CIAuD25PRnMktZ8cd4EoPYo+b9gswg8UgZ3SnQkSKqsRA8JcMicdJSDS5XhLDLueTdP
tNpIN7XQZAhAL2rYuOqDLACZYnkf4cqktnnD2cx6W4Wd6uevLVkCnOBg5Ovm7v6mly030Gh5a4Sp
c251iGPobJF4eTEe9yhpJ/QFb3g6Xx0gxYNIxN4kiycmNcrNySYLBj22tnbt7uT0TvXKYnILvxFM
VCGgtIULZejFRCIltgLNnUDapEm4MvpbpyCxrPyKhoDXG297k0/mAT5HGd2dtOKGD2VRjCZjSx7K
5mtiQOD33rPjwb4VL9QPV6YcEEE8ETo8ySQqzxdne+t680ROLPYAclSm4ztromtUIWa5dpl1u8Rr
MpS/+GERPc8Bup3zqH9QERuJ9keMZOqJ+dVJ7FLs/c1Wus+jhBjzghbqiq2IiiVaeuIF+J5eZFK6
zAvz2rq1ZYwO2heo0AAKMEUygQKKzFY63BqOudJEXKEy+qh1IYqZVCSr6eiIP2gPi1PuiXiTwkl5
wp6KnFeo00L6hQo7+YrrpZd2dQqoqaEOSuV6DCunU4zu0sgN+MivA0lptGwPswP51pec7XyWHmXs
loKH8Auee/yWslBF5rQKWfmoiV7QHs329ktwDQdf2YA4EWM1CG4EDdYvL/IfUEWUWZKxTnFlol5x
ppJPcNGPQBuAIc7IwfZbp1p8WeLpkUtCkzX3t1GqTqJfGbGv+5riLjrgLC6n7UqnsV/+JVTag2t4
osnU2nMn2LfB9Q3+HWGHrFfO/aZAOPCtQENQb8ySkDo++q0wagX/uJebS4P/kGOEeq0Ge0nk5leY
KbtEnYNKcQE2wAkaASpK1qVXqMG1gl2mfuKbpuzQrYXMhU6tk/IvkKRYH/zx1lMlm98CHOa1FgK3
W/T9e4w144+12cta+sdmbWQBrfBPueRRta9VbwPrQI8qawkA3sznQr6QYJcGIKGg1vsEBYLYGB7a
hW9QzqSKLFAa3uU6zXDgGtzYMTZkEnjuUEGYuyBNbC339DQYt8lKiE4LNe7E5DIpH45BVOPOKxm9
08/1Tr1Ouj1qJupvmLthpcm2FOk050l8FU24CZ4yz8zevin7zgxvvKgDWOeXu6rZPMhHtJxARwXg
OkKp0sS3huUUe3Id9u/swko9POhIwon0d0990FyEMlBpVSnaQF5sKvqm2nNlhDEIywLRT4L9dwUQ
JZjjYv+3kYKEcfQnDI7z0enj8c8nHUqYw4cThyAY2zaTGs/5qDFQIni2EY8wcptNuE993qaKCaWQ
PxQbno9x5dIKlM/atj49kSN569JpKuSYF1g8H8gKBMrTbg8s8yQ+gBWpMpb1U45hyrJeIURc0tZT
W+msuoQkjWB8Y8ivj0f/PrmpE740boejqlU9ydBRpnR9VDIhlhoRwPRUqR5eH14a669CpA/GSZA5
e9/gkWHG2jYLATSp7EvE6I1uQxH9+wBLQjPTiRhEQzOvxwfwRI3F1slDinJFe/jjwDY77h/AkAvU
IYWPIBfC2+nEt0oXV7uRjEw5uw46ldBRIxxsk1F/DNWbVYa482mQriQlSSu5JPE673WL/z7Pnjni
fmG2Y5P8Y/fktnsXKeDfARpJ4xmP8Qj+qRPFzdJYH1bnx22S4ltW1nTjDxDA4dr7i/keY4k2sub3
nfYe4uwAdbYYv8xGFiyJj6PsUN2LAwPhztiP+UpTnWTo+S5vJDEppNYFTH18S+0B/RPfQTyX4xbX
RWIQM6XfgCNQ8NkbLTJqZtJj1cQf3kxg1bgwAfzJjXB9bxh05P+QKeh0wguXVvZwicSMNEUw4WEs
DzFqQ2XdqsaHJMK58ZBmZBbmClWJgt6f559LNATn2lg7a+GIPaRS3lsQSxEzlfjTDtL57TfUemfU
Wk9W1vtNm2NSTN/a/U1VvpvoUdNsaYKkC517tVLfgl9ez5wjjgAv7g47//1JmbppXQnRuxUknYM1
57fwSJIZ3yvGMbl5kluAk5g6dO1CWlA+FLFba5ro9OIoZRWmD3750dKaWVzSCfvvYFXCBNyLEM76
rSopOW4viLxM237eMF9Fk3DKYw3JTeg9omBfd05LeuLO4/deexed/6Md6UIj8NOTbK7pBp3kNUQq
ULDKDsjWC3osks/TXdjmkVkbEIuBJVVbp2/Zg+fTlbrvCVxZcIXAPL4gCD9Zd+3RIuOgpswtOncu
ZOYWdhTHLNhdgr3CVxnYjvd39/Ot/f8bqYREmC5I503tNEj6DJ/5Eifu/AzH3bEH8C3YOrrel201
P/3DIAAaMYijGo+2cDuiZYja4pX9ZylSoAUmxtGUvh3AgGDtlo0T1HC1ptHkgXYTaLY9ABJ/NRhE
OuDaVU+06PI6HTx9WMFsV/rpYrwMcr1PYSF0ECcskP0N+5pwYJAuqyRcvUe2Tf3FHv3FriX5vpx7
ocnOCkuGGWjCQx6XCN5VrCs4lPJKiXDcm7RKCKc3FcV6d1HWf4tku0OU1EGrXc7IaAOICP8Wtn6W
RdIee8dBrYF2OMnDSb4BVPVqZ0p+pb8o3/V4GnOGKzUg466d9zqiI9pDVGsJx68CNrkjUsl878YP
gZs+VwMTMl9hnatuClUgk3epJbZetz944viaLnPynfCtS4rdqeYirl0IgP9qMRoXymutDWblPBOn
q2B2Ek7MpLPQ7tBEahgQNV8tHNPt/I3A1VgXsPxN7MUA4TSd0SWd6G6eeMy4/NMvjKE2wq/Z4cVD
YvzC2c8YiR/YKG18ISNwx1GlNtS//b+jY4/NgJdeGxfzxcq32FAdzuMl3HJQymXGS7jBKzDCB98L
3ThQ+ShIgqVDsrpeVTtVtzymSdZ81/wbL7usOIa6RLmJesQTHEDvMphe1QlDGTbPsCJ/sztOCHEU
ds8BLr7o86EcppbGlZ1AMg0ZFnYQhk8/lzjy73GB6j/Lp7VWEKwEniS0+12x686g2NLd8+pwXESB
26eTuYRfEcopI0U1oXQwwx8al4KJLqMiJClrVN8zaCvq+4Y/Vf3qrBxXwF8tRuRSWaXD6zdFbcw5
Qmw1x2lM08L/hEdjEZtBnxIfc2D4g0LZ6FhMmnQYWqru0EvueVWct7C6/ZMCWXFajeeEwvJ5mPFE
Q9Yw9mDG+AT99phJIAPHrKPVX6cQ9P1mfGP4vLg/1K9QCi3bnpY+rq1a+0makvwhC23FYXMyOG9Z
8gZb3j3dL/7drcIAltQffFOPHzygq2q5UjkSA9Wlcrd631PmkswMjIlhqDnTTSkBdhSiyCd7XKF+
p2T5h+pqKE3cax4zYscdsvRZFx9o4ljk5VZChxABN7tcMTD9PheQQGUalSVzdkbdRknF2iH3ICzp
QUoxnOmnbqJdjNtiZ0k8WwHxBigh1SWH3AlfKG9KKMvTL0s19TL73Lp5SmTzs2EiVGmgNBFVxmrV
YemTBugAe4BW7Gik7IfdK0MaraR1FnWMr7tl9gIrKzzIA3pU6RVMZ6YJeL8xDRIa9QPQbGTs+CuF
d2RFJ+KMRV29pujAXyo+/IBvHAR7a0zDMGtfHfqwuNmBBJTOw0J4/pCxYcaBtf3ZkK808UBqzxch
gKEYPOSTJJV7ADfgXihBMh6Rb1SoFhr+9Oc4lT3v7il+JWtj1CMn4bA9OgvYSaDWfT+fXIKWwlrL
tk8/G5ooM9/Z5vz7cEXXFJpF+BWzbrKSK7G+zas7luh2wC3Iw1xkT6mbozePSf+KY0VyumV385Qc
TNUWS2FzNKwWIj2ergb/4lJApgimI+GHrZibdyWC1EbD+CQ7rphDRBQeWZyYPEbfhRxHaYvLdTaV
rRn5ajFitX0qUQ+qptmG8D6A01s48jRXqziJRNRz8MbDIe4Mbsk7OcScs8AwAitgZ0TMeCwUZLRq
wDS9OgCM8/oFnwQajQ4W4lUEmUkd/MRJrcVxIFnQ/dO6wxh6nTvslpOe0RSMLbNyJDnTJwJANOnZ
i2uJwdNMpTzdtvyRXd91UvW5E8/q/CZGj3PC2WjbbQ+AKQaReQ30rw1UL2Gb0MHtShFRsfU/nAjB
ydTFTX+52hP05pCFWcGSXm7NjyoAa00iiKlPoCCFDgD9/pf1k5N0CVrBdtpCgOLiFvyc85sphrSj
uU2zHGxC6AosgJ47E8CTi942fyAjkkh+BlcWsXPxVQham1kvIQnNbjCGaJNQoKaiA1CCRhFm2vJx
hzVt/ZsPO4hwhW4fkOwF2jNLdXybjUizl8c30PF5uvKWtpXRc/uwBr7FlbrEUnVbGTKG25DBDGXy
6lEP+3K9BZnNS6lE5deIXCmGvWWSJIuFIEs+jeQmqR6I8DfaZgvkY4dhilHuVwXFrFPxdm50GWpQ
8J9NKlw1VL5RLECbtqlbzQbZjRBBRblZMCxXl18g8uI6Qmh7kbgOFQOlTQmyRrPGfgmDqiTwsoz/
PhqHDxt1YgD3qquvrzknRPofOoBn+aSTxZlSzva5i8lCjLy/+BG1EvICiaXC55wpGLtV7akotWw0
0YiUaxUH/dHmlTznvkguoEKBaF6YK0dNUtmeNlSQ3jjzNr+RrtZ1Iw0YLV1/MELoK3KWzN4hwk4c
pwsJKQrQkkUpqbTjPpTusJsR6JH6p7ey1iweYqOxIDZ/F2K2wJ5voJnivlIvH8wi37BaliECh15U
KZFQ4T1XoqxRqxTTtpgLm0EDmmXw7YmSV3AAo+i+9DMFEL77Cje8gXWJtDcuOK7pikXVP2yYoQHX
WbSUdW79yhVSOWGf7TwiWK6Q3ifJIxldLfc/2D/UMILBl5O3OY11PlDzVxD7vVBx65IvWPm1j3fY
zHo1KuSY17R+wbw9dg/4usBqQrsbi8V5Qgq+c97vJR4btP0qb5ZIuuv/lykl0z9tkNfhdGO/r4Vo
guTELCASETxdyH+ChcvU0G7kFhvwv4rLhMtGluvz3sVuC9tTr5qjwCORFaNvOnlQyISC9ctKe3LQ
23GDfEgNDPKmG2EWivtZxEDQOGjlgxyNCmEklzHXQyZJbcakJdiOxHb7u31koZwI4+f6E54gKw41
Cc2uc5Ub/MnKoGTn8pvQcRuwnouShXBH/KwSPuitUDLANrU9kxpFLNonPpFlDZztShSPTswxWPSp
L84ApkhjHmNfVyKyrBPhjfZ/Z1LiBgdK/OvxHBIHCfKOptgp8LSg7dgfSWpC9GifmTf1es25C1Ns
l5TwKMRD80lwbhjnob0OZpOaFfBs1l+7RDJ4U+dBcIkhGqBUDC04ccAnY3BcYfLpy9lFpEFUBnuO
MJg0hc239hCAyF15/rBJFfe5dDnxfmBJCF5CkwIKGw+Ykn3DX7CqxN25e4dmRt8+b+2JKQFe1XL6
hpdIP6/8l4iyWQY8OLEhphQcAb5ZTydIlLIENHnDsGjDDR1uojwwzB8oZoirEOMiYdFguHJpc7Wl
qcOjjd9354wqF/pvMnz8VsKhxZ9FImDo9nVlz9PeXZxH34gxVVq1CjjACN1oQVu/O5fpOyu2Ig4J
5lX6Sw2vK7qlEa7ZuwzgHLjYOxF2o1NvwsiUUO5nG9SBCbDuyR4H9CvHVnR38Wt6P3mfMa+gT8jc
AI9VHhJCB6eTSHUj5yw2rm3NFnsD5DWIN5L1uRZ2griHcYrOSBdEXMpbakMWynIbR67Ps17nNabu
i3CsQEul5NvrbcjxhK/spGzWIGRoHE0siVUjiyHLTeJNC4+f/ueAqldsMSssqISqSMD7CQhAStEH
HULKSjZLclL4bUL02QSdMW2A88jXfCs4Mj4vm7QB+lTRjpfek2semt1GJHpP42+510VSEja8+R7Y
khMhuwW6mJMQ9o1pdKvRp9bUpCvi2HCI5J3AaWGZaQAlqxRor1fbX8aFroWmT+C0FABcDbYdNj49
xtlNUppVemcK/zwH0wrec5TidrJ26csFA/gZs5FZD+cMY5IogMaD3kt+nQIX5RneLeXE4qc6Zlbi
MjT8BS9N5hVJQlNP1xyMnQ16GKAwyr0bypDgvqNKafjoYsPPX/rQlVICJzWNrykFtlV7xwL03GEx
5/iJT/XEBYirySHSYhwsoTftFIKyGyxAFtGlOlfbUVYt1dEPM0kbPbpV4aN/JfBrwPvE+yk+yOuo
yn4yQa1A+2aw+ELxen3bXEu08HPD5N/eheGmP54Vf7iiOG0TedO1srIsGRgGSlWgGn1UOKIF8JbG
SQqrlW9fAS/oHfY9M25dMxaxeF/KZtKGQ4WM4ScjZfArRtn6aqwVIIVYoglJvQk1th/DnQ4uLugb
3U46TIEtVARQP3iZ0wga2xV/tmk664cstMS48Gx+JBj3sJu9PeDnqKnt+hWi0SveDQkbJ4gpLZ8B
PmG2VV2RPomkxXP/+Yyxwe5IoXeCmFGUnB4TkAkhc7uKvGr0+SIALGFQGvxecTDJdrASW3cabf3X
RGnK6zZdnrLDX0AlQj1vLVbu0tBa32Uh5cfH4r7IzR/Ff2lTLVnxiDan+MCQmAWG7z3JIk1L7PcG
CO5fEdy6mvZ9fPvIsvJRLBv8sVlku36mtTY+WUKJZ9EuIq3YY/sHhOqbkFKjdNJdak6I37PmDzC0
xp4m8kDP3AVNWiQc/CtL2PQ8h/Bjwz6pkZe8Eprq2acFwh9vpK5GLYT+d7xwj/ZLg7VXI+ti2sYp
60ecGWWH2vECAqxXzgXtkzmFxDogrosOXKTXwk+mMPoxcUnxRFpNe1CN8J7ZkUTRUX0WZlAQp8Yv
ZnxUioAbIkgdO2XHO4Z41Cfex/Ouf9SMW07OzKCOSI0ti28Ah/ZntvD+9luLAufppDH4QJPhwHbW
HbFWLVBu/svsmnsapf0uquGC9eRHPIsUmImpCsuXNoMa6YmxAxvYwdadqZ5bC0Q72U/APpFzqMCn
gQt70TOzF9dnIvavd2gIMuyII3AVLZv0L9VGfkhTTdQ4rJnpiUVBP96ySrQLY5UqlfJHY9D0ZHFQ
Ol+gDbWW3G7GklgdLWYa/NlX4P/Bsb9xEkoU2BtKgIDN6HT1x3gfHi7my8dU0o7u7BShda/7wVrm
ip5K+RSFcwdkuPn5FlYHqdieoQGWrcSXPkXOpus6oSAHjzMRyFyiIMLN5kJS/K2KIsRkP27yrXY+
wazG6F4yXX0W3sRTVftoW8fVmu0U4lB7ipTMOZLrabBlPc/72zr9iCTNQdlYMp/tC3RzsP0C8vTt
nGCSpQ5OR2f7IOoSuNz/moz51FOyVlOyWNLJipw0YaZGNddqpCH3Diq9DcmC8fhjPk2+EQktPU1C
ytJSd9NgbVzrnc8Q/3h/DQ3LG82A4fIfGSAWu79ZzZEo9Ew+RCv/mlZJeL21vhjnA8fj2skN1XKu
CG9fTMeHDqgxrv/x1gRu46iqz198kn2vd+gNNU9sO08gxykZtDylQISgemNoPTYacXMcrihKh3Vz
MT1reigPfFdXv9WmgAEG+Xa/oiWPYQ+z8Vtztl7vBfyWIfdY1Wu7YdyZkYsZFRfUXtd7MB4F5Ova
Biw3mfJFW/+lJ6DnFJ01Hv0+w4LKyevFPXHXQGiH6YJZbKdoE0kqRl6rUzTcWCTfUP+u9sRp1n7m
bPRRsFPDokTcgI45XonQklV6oHV+eKVPohGjlcPl8ALuoK8N2m2Qvwl46B1m+3kfrsPIK2/wHBKA
yTKDtwWgu9KciOR0bgoI19IuGUQSA3WHy2LBkLniQyl+nb2Q3oRSTLx31sypVuVtumGmi4wdw5g8
mx5XpmmebNwcc39XyfO9rs/GlCCl/0fYvH0Pqam7RA7CnRZ4vkgs0wH7hFKbNzfy7TiQvCs/URZZ
Umvr/N1KnacHibGlwHeT0Qz5OTWEqm8sAqjySWHqiTJ8+cNgW1q/P/AKig12X1xHhXUpr+1x7m/H
sGvOwYnmLyCGyyl4UoNHeFpYa7pOzTKoF1IAxbxPd0j0BmTq86QeP6mGhw+wQSe946lV80TzZPbS
C8UqdOJVkLKQkHYw63WCTHP+Bf/T4LfaEImpAWnJ41p0cFhAp+r2bpxWeCHjbLAfktEZowZ5ay1U
EDK0ckHEt7INd3UDoVNo3O3TsSIBqwStTTIWx8mVOHq7i3dTDIeK9XWnQcP12soOYtF7hkcs9Cy1
7c3PRNvpC5Fq6oZeaTXOIYvQNu+efYqjv9LXeC2E6F83m9TqspsUAU8GoGIXbp5qnZ9x8jjqgCeP
TuCxRCKKpstsLlMFyx3cTCVuiArkydYMl0fwjXvvHKsnFArvt6uqRdFso8tXv5IZI4jHV7DxSKxe
/C0NokNNq2eu10iY1KNEH6jWcHM2iExhRH7ccId3IkQfx9IkQ+pdYbZOYYZS3CLIAqAfqBN39QBK
hAHa147D8nZoDQqSxyjLpcb92hhEIityWIcIu0GMKW5brXuT6Rjtezc2iW48Z+WLLEzSNoECULmc
/Vk6i+dZ0LqmV5YMYnK92i/gA8vg7ZpU6hIFBbMz0LzJJpFEe/SaVG3ac1+yKqtJ8LPlvqoO3udd
DXRuMXIeQW0maKJGc+RW1FzPE8Zn4ZSnkSoQOBAR9vNE6Myp+5MdnTmd1vTXZCVIjIRYK6jwqPLv
9rfLgZAxDhN0UCJ+ik8GHEXa/0dz8CfAE1diipNJDFb5Ek9GokP3JEv5sKbcXYMmOiH9N3LI8S/6
T1zZpDfFf0U3pHU3nZkke+DRCydXvKHXQhL51FdiiKRxoQbomphjp+3mOUrhhVFT1u0gHafcgO8h
CI9fAQI6gVDAB2O3Ir+/zuouZuhn17bXPcCZZfsZ0VoBa6T6AweurMhSPus1JA1idby0o91yMWK9
YN52lYY2mvJlMTg2Pl8V+sC3ECactmruBnMI5tEwmitWsQP6b8hDF0kDgbpfwawK35p+0+KhWx2Q
ZcPVbJ2y2YJErXVHMUpx/GJX2es4R/ZSTr7JMUMlNrDWUv67ku38dlV8kL9t/PnqR3W2gW4sLB36
ga4hZiPRNXthX3uCiRVXHQbpmdfGfzhD23tnmII7g+6jJQphVaBxMV8XAhNber9pzvWrzO/YPvyn
wkUK2xga/EiBdMN/UJoRBDwQWKyKS1vveEefuZNX25mIViCZO3UmKL4R08uUQNo9H2+Mc3jSfW6r
YhkaT2ZaHZoxDBElx2dFqmhobPvkuXcBEMyvuktWYADm2ntH6fpW9w3GGLlpFsInNdDL8I7aLcak
MnWHYk+ops5bg3o0oCsfXkBGdh7aI9+ZDITnoaNNJj2KI8gozAMSP6QZntctWLqPaE9KfuMRHqHV
5BW5ij+cXzpAmDxwF3yGbVdHCI2P5bor5VblVVD2ubBZXjv/1GiHwsd3dCGJEeAZX2FQpuHXP3/Z
ls+fOqavYUzhtrSjW7il0rndkenrbCP/BfkMee1sPNVV5H0oLuJHl1rQn0PscmbueayXqxNXv9zr
6c6pVIYD9TjX/jxZHpwDtpi3Y7eGItTSZTaR6dTy+6dSk9nKZXVSI/BS1HR4zWPXI5VSFNoW6ZAa
GLNYQoSaHxqk/X/rSyBJJXWDp0e31cLJF7ZuY/iVqSyI4mRjr195/ccF0TSyoEGMBBNA6AqQmS+6
RWRIBo5Ha1ryGSo32kNvKHTubsPR36tAuJ/G+pjXyx9EdPxZ8X/F/waI5tIPLckvbel5z3i90Y2N
uVAEcGvJw1QIcs1IWJ7YcWIRaIi2bgWbo3pNZJuRdrDbpBwQOiy/Wfo6j6sB5A73uNH/c1USJs2/
oluMoVosrLpfzDaDCbsj89VuSF7SDKa7kL1ELWyxRJkkhWzGVmBikUKHCkoyLFBsHtpCJ7UgK33c
BYW4MooiR4BASzNObDYXdsyRdnmJHBCDewk7YZesvCPWOkYyYLnorZGEPkYbmiy9FUclflTs+Ikh
ihOpD2tAyTpWoJk9nwGD7AqKjl0ntd6Dvjluy3MpMA3TqBZmv9+QTEEAd5wTD8HB2hMA8qEJVp3U
sZGZB1MY5S4p9VY1kt1HMG9IOdJ14t9/KAJDLPk5Xhti5+Rn/LslxqOnspeM2gjCsC169AyMOB6a
wqjIGwfBgStl9BvdBeZDofkFC+dhpOkWB8P3aCG03hrav+lAZCmExEQS+n/Ib4Nhhwa30P5KUahc
o6CwiwE3t2/7s/4WSK81uBJ4B/YYcNpxB7SfkEB3dY4FeoL9v5v8LXNZrclXn6qbHazhi2p5mQOo
7pZLzAPmI+47Y01cW1JRDoSRaPTOIqeyaRQYcAfwK2lb/MNauPYI9SPHbzNUs3ik/WQymQWMKWge
/G55r/Ml9HhId1wW3DfIQqepCEgmjIhLckJFSmaoz52GCX6C5MJH9lk/IaKmWzugLNqlinf/rmvp
GnX1N4oLTKdSSUc4/FZDlsqy7wXY+yWQucPv+jiL5cuAkknY3HGKh0dAOuquka7Y9x4Qe9ytLvRY
c5HAegDM5hYatjXD+lIepOhjh3VbXg19Kg3xvHZW7aRA+oEm9MhHKRgOq5Jm5wrQeUmTwkAp9ixP
3XmBb4DEtrPB1vZN8rUVi7Pc3VhvdqKAKwH8ibLwH6y0tmRj9s15fOhRd/5u9iuqN6lvUNIsa0V9
vEQd9OvJ+h0Oe0H7yhShM09VQrShC25GdI4Tv3ryv7nQ2q5WytKNX3MrEEiaEntlgeB+3S444hhj
4AO+uqKkXHv47HhhscSOSbHanidefCH34CYeN6ouWA3zUh173LqoPCHFXvlle/tdj1nMyPhFjJ0x
8O79BLWa3mDEf35MU7ziFX/yBNBZHz/GBacnVyEuDZM5uFYd35S+lSdx15YMnKw5hyWNr7VYM/ud
VL3xIKKsgXvccZ1LhFEI3MaubiPGzXwIYSbnVV6VsiG7rvlINv/9j7yiLKbJzKa29u0PPgOKSqcp
FBFc1gCNzANcfDmFBbLg6eilnFv+XYTnItNOusRCefIR4PomwqO0D0tY8L7xXACmSSjkrKZ2wESS
+WFk5/W66fPoxFhMvh3MdO9WF8T6kpeum/lgl/6Eu/q/0tnjpW1i5qIEa668KlPqWYjwvObWzJmH
763iITkCATpsNKm9mVVo3bzvRvj0Uocb7Ef0SpFd4Lq0XOSPAFajgPD1DXbpMsUZ/qHtNJQjdm1U
iR0EU+HHoiJUp94sO5RMV2zRFZ6R7DGGf9qFjTVMmac3PEbn1fHaeG8FM2WVpJra9FcONGawkI/i
RKLrPgMZXqkoHCyxumlenkxbqNPiEzBup+bkMdNcutpVaMNkg+A4rwoPJ7+94pSyC1NnIvWgvajz
4UX0FbGurjW+/wu8SOwsn0cQO0C4ilE6BWmyPK8ChByHJmkMhbo9JU49oSmD4oE8HKWw0Ar9qTHC
LTWXLJ5q7C/5dK1qagI/oY/D+yokXPTJCkCA4vkbZrcGMBywboEbIZoSfO/KWDl9BS2VLVT77Y1y
WQ7/A3wqB+KrwTZogwWqvufiPYuZX3MbFPFGj/EoRXzgt5xZsh4CjIjXyYlzcF5U7H7sxcGwNNQv
Ef7Rs4rKQ72Pbp41J3fVAqkLo715+Cw6avmQYbduRoZ6IMMsTOHVZ7mZtv3S9HWCRXeWj6l39XUl
g/hV0EII0Jfx2tU4BB/HNB6nWkjMqNSk1ZJI6ipxuUhHnWX40kUednBbPtMZtHgRTQiajYzq0Vd+
AKVsPrVoZy6hVDuEIIVfzlNXkFmOw1ufLWOx6FiQnVzZtOfgpyRrlVC35BMcgajPeUdKegD8wrB8
YRf5GD9OX8G41xn1saytY1oSkEGYBgm5p9j8mItaL9YTOBL5ngtFq1MlsUIMxS1YWBPEhhk+NR/K
WKSCvkFSWGt838/dOxCLDBCV2oQi1cuihZmdcnhgCTtpzXjFlTe0TbLwn+hH5IxXlH+Ll09GiFvN
ZNS467IhF0Ijty8kt+O9SOTD/DZMpbBZpIvUDeARTzPbDNsjk9O2g4qbhbCXQjn3qG542WD6rCZm
f458Zhn7OJbO5WCrL93cw40uAXF/FAfQjg0ItWkvbxdq4O49xUcqKLhlHEEdQBY3cBYiHWgZlBl+
AIOkty0vLPrCBbOIuL8JXoNLZ1EMnat19Eypxw61GuTyR28L1+o3imFoHIIZAJhDxfiGYWZb0zEO
1unAzREft6oMgOWA3TebjHU50BV+WkdZ/r+s0DY0wc8sgj4L6pF13ZLyxgiC1dfDqgIf5tQrdyx8
DZ47N0IXvKVDfaret3Yc4sOPjfn9iX9mJroTgq/NcTfO0nHelGRxFbdotPtcbgYmX2QqaFdptp04
CQmO6MLdIgQq/1FTu0nfk2VHcXsEZOzHGoyLM5/zVRI0sSxdbQGAuh3hAdq3fUE7NEFhAo3VA7kA
/A4ttZ/xVAFZxJHXCMeg6h43tJJtj8uCbsdFelBA2Vud7gi6vyrNfCkz+ZQIIrng8jMwCS1qC0oh
2DYBwzk1m0LJtvFb0ImLI/iFMsKTWOOKZ/91qwOeZUuPCGJYlpchNVq86gMr/jfhZ5/kp7otGJtB
rVSfIfk2hIgdUvNUJB0GZJOQbRHPvUzifalsgDuEzt8VziAndUMGlCJwzPRwZHWJ2AZVVHAawybb
JB3SGlfQU7vOV09BJPaEnCeoLBIFPcWbHVlMPigdcOJb3t6Im4chiqeRn8ZhSTfJSo0BE7MzR/Hl
ChFWgH43VjRJVqB5aYsx57BkVqxBd9LzN3BkdvY3x7pWd4xBZNErC5WTI71RzYyHHun4fhHujBTA
coPYHvr36vWpG1WST/Ph5D4uVH+G9QHJXHWnJapxvjjlh76iSgPaVgUZhnQePmcCfd1lZrXbKBIU
keQsELb+NgmPtnFtxre5gApCKju9iSzfHJAJpQhwm8EF4l9MDd9XL23EdVoJEd9ZwRxDtoUf5LzB
JDNPeco+abp610ZZqdWlUzxFNqFQDCb/gcdEbbVZ62qeS33CU6+UUoV8qXg8s9H8PzOfkXPSaoNk
an6ebj9DDbo/uNvzEW8PWGN1xpfsmaGkef+qQNAVeViXx05j/tM2RbDP0Kh9g9D2Ud3rsVv9D8+g
wX1oPO5vsx8RHE7xzy6Sz0ZVnfZxgID5crnxbCF+wWt6EGwzA8szFrV6o995S5Nl/Gt0VX6vRf4k
A2neivdHb4FtLgLK8+5mdcI/D2qYKdPoGCRHL70lh51+dGhuz1h7n9wBWxu2c84WQwR6wg4sLwXR
Fw1X+bUu8WGxwO5CzP9D0VFgKZlUEPeAoIE7kMFmXXpZLrd/L825/+OCmf2PSRpqZiE77SzJRHAG
dUUZZiYrg+Alt/oC6XrMn+A37I5CmHqdo/zZrUtyJrA9XuGt/BaQCQ2uApRJo34tZXBVG8WZ2L7Z
A+QUr1h90VjaeR55uKZ5SGKR9JOBt9oZfNXoeQ8iKk2bN3+/W0zejioAxN1asoFM1Nih86biNpfD
udVenjo6FTgXR7z5f4lWKp9U3G1byeHNQqO7fKFr0pB4sCNKvicrUkH+VoTBxbAzf17Gg0kF/VVW
jWK7dYKfrll6XyH2hKAEsN2Ik9r0uWHXR3WPj/5pn9Z8sulh/W+c6iHdFf5Z/PA6SQhfw+Z/kL05
boGAFo8swfbStM2faysOOy/Goq2Cg/SESzJKjPfvCPATrNE1NdqmGSH2LkB171GHr9VAgommaHIZ
+RwGqzjYpCeIFxrfQdbu6W0Xxf5qlzq8hc92T6lO+Zl41tl12u3+HPx/l4gjghatc+eNLFedew8j
rFM2xPXbVjsT6N0FNoSpMHfBg/SJ5hU1DkS0v0FwsvYzuThT+aa2+5Y1BX8Rww6k6My7VM4N6Xh8
sw4wZhXtqmT5LIILSmpahfeeXbsaeORzcbSU1cM7kJedgLeEYf+7naRS/Gt+oMX+Nwtfm3iwCtMZ
V3BgArUnaK1oXtqV0QBj1ZlDMLn9Y0CjdTm2pP0xagK0Sbee7WoGIBxl+QobU65NwlG63H8J5mEE
AIMAYWdUnYT9Om9THFrj53Bwkq/a8IH8fvvzmJHWQ44Sko/83xr2dbSw9uRBbQCdh9Zin1C0J4L1
kue+AeWYZsgPitcxeMI+bLGZrI+xxddQhHJY9K3DDNMUKn/tpYl90ktegOEmtSny6V48TofmPesl
2dO4zGi+wRCMpqYtO7/QKPdCgtAn7nRq1rmWptrx+FO0OJBDC2VujmgHQjvXOwc1pgMVQ8H2igoX
v6BF/for/TSirqd6N1/XDT3slWiOYtoCbag74SrfNMX5TVacHnZM2+okItoJ3V+g9YZmee/oqLnl
HtMYRIuR0Bp+jAi2eYrlJEqAmrL945d8CC3rAOe/GUZmrqLJMn2Ezk/0hb7t6vulxsJETAot1MUn
EhOpJ814jw72KURoo1wnCYmQ+X3Wv2bjlfPitBmU/GbDVKDQI6o/Cc+AUwqIDUKrwectK3zazu54
FfWQFG8PJDlIevbRZ0aUNS1Wzg3jZ9wOihNA6o+LZFRnf+GEign2bAAVS1AtcnECge0ul8hNvYG/
/YCevHkg+bRtP+vTrdcOpAyO0lSFT/BettBWvdJzAUNFskLa0od1w7y08WxByzNcPz7ZiK7jYS/9
P8NeP8Lx+GFszD4yReiEbFFWNgea6EJx1TQ7kp+GaPywXCyPskEIc/3a5EDrojs8zX5wwbo6HCz1
/BqwY0DsUClNLGi90N2vB1PfrhQLZ5Q3Ks8tBnwRIzAg2UzTOveSkWJKS7iVZxe5NArIJAXOOcPR
WwZMBBKoDeVoY3Map/5tz0NeLu3IRJqUTn7f69sMvcC3evwGaypvJc5JXC1M7PAcF8TTGCPqO7tc
kBTqKQ9nS0ph8gpjb0PGbp98qesEIowBELcs2dULDgIy+0QuNz94PatAdUhKXSDkdW8uE+rOVQOn
Sn9978P5t3L0aWB9v/4xfX3cTPWiRjjdbQ5FPFahzJ7V3YGL7J5UZ5oLm95/Szb4odaKAeXusPp5
mf8RBBja8IpCPfevmPWVuKyRuUdvPi407fDTpFKhTvc1CDz5FlaoyEArxzHwJp3NhdPotmSiMaqR
0CqjrfFIvmX9F+i8Zs30iGmeJITkkgNQa5SAjz871JqdouC5qH1tkf7E2RTEv02VYYnoHz5vyq5Q
d21wuyJyiWg6shC5PpERMU6AL5JHwMCspOOyekD7qqZcOkR3gr919v1n7coLh+AV2ssK5yxud52d
mP1hoTw1qx4IgdI6kUkF4gQNqbNgGoto1WC6zsFL6UUU0GZC3Klc/U+5unlowwlBz/PFftm3Onw0
c/+W1Bi1GDO3ste6BqSias67VRXvHFoZssEAyRTmmCbj7wFAYoDGfj5aVT39lH622ildyLCKyKeV
x7l3A/cxDxK0kIC+tNJWClUd2G0+qkyS+0UTM7PfGvxkxVioa39hVA8nqXWtJNgimkb20w9+s9BW
ujtkah3JAGrzYHGF0CtQuuDZv8HcCFcFFtFWANk1PBg3JGXO9nvmKWhnCYNqDX8mgjq2XTTbOi0q
KAm2uCP6NsL39Lif6AwXzozVumoOgZoVMmiVedSdiHfYjQLRczvvsh7nW4EDgwZmf29UpVDQDCz5
wh8gepLE93tZRNHnu+siCpVzQOHccDoiXifiNkx/OmrKcBPvuKT/7+y4hEc4ohlPRpmt79lrOxA1
2cXuySb65SbcOI6c/dl8VKDgMgJ6XjHOWORvs+v30suTMeuxTw8E8v9e4ygUMwgxa0DUho8QJH1e
dfD6y/KjQaNdOxCGmx74qXXsEUtK3/gVSr9LR9FytDRBDIO8z4MsrrEHKUCVRdApywQv2FXK9Xsn
QcX7cBG3lHSgZDax2LGNZ+G85QAh4Iy94mpFPMlqycj35u6M8HlVGS1vKa21Sx/gScayOTmBh8nf
THoS8vbnz7sdSMEMQHTeeVXcItzd3kSyrPvp4LiPsf1DnwQXl88Yns4LKBgQPw8sfviQ+6JyeXq1
HzwpLYMM8DrgyEIUU/AYnDsP5dS3WWZG6sFG7yOiPtWGhiaZ0rLTvgeNJ46VGMbluW6zN/6i2eOp
l+4A00KWTnX3MdtYE1T3B376INluBUfHCrIAOIUXTwzUTt1iO52bOtt5G15MlC4a9vWktk7N6E9D
Wzb4lW7hhc6lF6j4Vd1qNGLYx4lih9ctdBQcjWZTo8GD4u9upYVpHkVF+L5uSIbUXyiKFFqvwVnB
40giuQ2NznvN2JUPdWwHharkM8j/17graoYzr70ox3r0we8zAA8d5sdeYpMVRBOdNVMouh49AIhb
7gwB/Bqcwku+mQWD3FpIVytnVxbVYialHMLYKndMZFhB+1+kcTh5Vnr0vTrEqTM0mSzsdT/XDkEf
ExUHnwA3JyVhTdba7ESRC2tmx54lcpCJL49/sGmhzWheB99+5SUv2HKuMypIPg8l2SrUIMX5Qntz
JlfmupmLzx3MtPzakoytWgE5dQXLMIzXJ7iewglltV0JlYSCeCrZSRefAj9vcUBCpy9Bs/fCm6BH
P6hGpx5bHKa9z6MU6q/qkx2iwEtaDgnvUosgmiiAU/pqxFBNEAi5gFtILofcTa6UucxdB5OXpMbw
P4/KK9JDsRUB4S7cIKPLbX1hBDF0I6MWYV+1BEDB/lpE8q0WecL7CMxZnzQIK8SfSw3O1+atkVtG
EgqC8xihsHz2LpGa2vQouInV8OF8CAM2yLqekBWq9uhSHjEgxvXNNUqJRQXQitcV6Wrd6BgBlSRI
YC4Y1wTuLbuzi3Apj8Tpkul/anQ47xlAzdXhdQGIbwPc9DDLuhO6xj54WUHhoplzJYp9PcFIAQnl
3KsKQbLBmUq+QbNb8i+F5wqNTk4Sqf7tRFJ5d+jwxRS4IFIE12ewjvvdmbm++yc1/ZxcJmrtcvmC
QCO0B+m6obPDBo1snJyJPH/bsCROtEp5kCxSj5eiqmv5uFNbNWq4UBPGVUvcMA2fHLGggz4WrIxW
Tfr+A4dxpvn56crowMVCk0dBimd04CmkwlFM6eAYL5MwYvyWKWQyO+yr4rQiqB7cu63IQVVDM5Bz
0sa/SUIRPsGnRUDztDDDmdpE2ohCw4jajcyOkKbrF6cZ1u6hARFO+VdlvSPtdJ7GzV1m0q3RZa+G
EYft3SfGTUt+TVJHyBqcNT01xroiWpiUK1umd6jtLOK78RDpWkGZ01CW3Dm8Uu3d5X9b77UIAWTv
4vPC7Gbk1F9mkssmh/5MCrzPSZxnTLfK41TMM2UUS0AoKoSJanbSVHxMqPFsO9YWdj98UFD/C/bG
PinhyMseZ59HOCtoG/M1YJatWyYPpc49H48n62XVmmmFbu6C3ybhPXo7sehm3cNdNYXWUlFscLYU
Foc8VR5z1a+Bwh2lrH9G0s/NB4biJJqoTW2SMKqZRgKjPUiU9eRLM6eQriQesUmadoQCzVLtvON6
wGV+rn+hYmuCoJvhuBnaHdFHS+uhHyohFiy5HlWdpkd/Daf/ZRUSeY7mOMrr8BYSJ2ryCnVoG9an
Mk0bhMMyop1y2ddfbJC4OuMnU4X1UAcqP/Rt7Oykv3ToZqaEETlR9JdixFyhWT48ZGwmsavYPkpF
xmoZrwp1vZ24TtvdIa2ikfYKdkiJVLXiEZZ1nuv8Q5rFprS4L6a6uEKrJcmVYSYbcKsZph8smUXR
ZQiZc5emVeE7d7qQJHQfS6BbJS0qwPelHrA85aP9zun2iu/uQusleQ0RcGsKwVbkOrdjPf3TyhJX
IqrzvEIKhr5WMOpc8vR8dYLpWnIYLhcXP03rxdaqFp7hKJUbw8WkRr9lr2lzIYvM920I4kRqcaXL
mzA16MBM6WjnYV8z4v9f9HgiqnNN37TMUnbgQyiwfJ6Th3u9aOst6G16UmZUnaTKBxDI2hE/t9MT
QygjHTd/c0CftOUs0r0QdbincAmIPMS2XeCRoJ541nM5sYYqqE5bCMdrB9TALyaAzBllYX0fHjmi
rkcufVWAfE+dVNyHwAMCHBul9jlOjJ8gL0DU+9k5XF09dSft8bOA/yKJP0oLCXCuNo5VT10h6c9u
k8d0KYtzcdVsLQ7Tr8HfqrOvxbeEr0AufDwEHOYIZTbc6oKxL4UpG25KAhuZA3mxV5tF94TtA6KH
8TM2wmeG77D3gsqssTFeoA1OWDcDEbRXb84pdVIXEik+8ns2wHffBOg1ZwE1IPdMQrVuwPqIiQbq
+0yb7Tloqo27/OBaKsNIrtR/w9NqOEzfV6msNaMJuUITOXniNCOWmQ0c2H1mhQETgmbHT7hK2p3z
36Vd2PDPS1nzDZy5Sms940p5DXfhjeK0zps82ZaUf2EyK8eC1JlvjiO0YOTYuNXgP71bysSf+US8
b8/S8aegt983/5sv6PygIdkAd/dJUPiykQz/JOlrCB7LRnKi78UA6ebsaSL6x9d0mKg5iA/6Y+bJ
IkQYeRZEe8PlAfrRzf+YEYFn7JjTtE+ALvdXN9EsAwPsJTi+n4Viyw/M7H+pznrtKZL4VDQYYdKB
FKj+BKgcGpJKrUX79VGsAiKZyxwfqR9vCb1m4BtJXdoK195XR2PrzvN5tkcMHxYS9P4bCS38Zww2
qtk9GOc7KshYNs3GkXFTNqUyoA6zMjP6dHvBgz8F5dQ269U703Z2adg8Jw5LkyUiy5aNXj7eiwjs
Liu19W8k3Euj4PqYMCB8NCRL2K1tHNfk7RtHny/OExu8vLzqJovsutPz/UPo1Y3Y0tPRziFvEBlU
k2nJWdvrJQzFTFNmjwQN0w9EZ3fap6mrf5PoqRv7tWgDDFVdrXq53f8dXAIkMpHvxKwzS5x7a0mq
pEGEd5Cjfai65MdPJkO0O7KMt/Cqm1TJMm4GasIzPHDjCokHAQ1WReWT7ggeigHm/Ba8YrM/bieo
gfRqsAZm+xUzsN8htt7+6LQ6Y4vGgfTF3qWG+8G33qu4o0pAtdayw9t96F6WU7MojVOQC2Cj/zwx
WQ2iDvoBSffCaEwEFQnhoTAc+G9UxuVN8bj8zTZfcaKCkMUHI88o6w/0o23WuWMDqhccVxdT1nHN
/QT0fvpDbmUBALaw2VG9kck+tBsQVgJAca8/iaSAOKu8fo1GSFD/IW4qd9gdrt1311aEkTSWxCBw
SMkxTH+bk5nUwJ2uswRiQD1WMaAR3weznEkAnPSYUFqmbNO1vLLDrmWmFigHn1k1xytSbyKXlr2t
JJ5VMjtbODJm1exncRxdpOU0GkiCSfyCjsa86w02LCnUXVz+Kthjgi6ePHwAhNXV/N0T6FfeNf96
lj3RVXGbEnoOLg1RBbhsz7UyRY+yFV4QMncEUdNniCCWtCakUN6bzgquc3UsZzkTJOoeJ42foEnr
N5JE3VZcCDOlpP72O+/sPOUfr33LpZffyzaHL+ZPoxWpL3TBfa+Ae5FMH0wMU9ubAD1rxOE6gzpg
OwaA2rxKxYZJO98KU406WhsVEUx5KD2BKO7tM96Xt6uVTKcFgYQR74posJKfUyFbW/GQsiV/eH32
FMe6JRLsG7p10fUiN4ytGBisc5R0dD6zfoi7HhtAP8mZSkcGBcqmXhQdDmNAWmYM+RVKfi9yGYzg
1yqTA5xzWS/kRpfhxrsKrnf/6UEtglNxiqcQzQRcUZ0UuOPQhn3pCnWD4xnKdfiCUxGaayrxgzVu
HFQbBQApfna8IPYJh8gsZL3iubsNH08VGiJjlSN/KBkqJQS003nMVo22HxdekCTLc38uUVOSuu2e
B3yYmj5nSg63I6z4jFbrNmsK5A05Qd+d61AO8vR8uo9NANzA2zGvhTxXZOQtTdpHQPNL2tMvYyVf
1BejPV/ePq+j30pgXIHn/hIB3p7x0z6t01x22uEXkkUpVmWEfFA9GD+NOEoVnVeKusts21Ktyf5c
zOjKPkgcMx1MnsRtUvGJr5CGXe5y+PARwRX57vo65B3NJhD5cSDVLnkyIWXsNxhU0771YzgAkrVT
2MclddiYXVpnE7M3nyS2Wd29Widx02TvZR6Fd7a1HaK6gs1NgnoAWiO3EA3Ko1QQoXTxm6yoxwDI
gNDiuvP3RZfT6y69x8nTQK5mvJz3Wo5mxXZxKWTRpAhdZwYc3rGW4M2LdfGDPzmQST+8fNvZPmyt
dlvtbOr7oa716x4ZU07S/jqKCQJcP1Vgo5Amw2szBNW0q6Nu5kcQRdpwVVCRwd/JidELj0pY7feH
ZdKrRPRoHoIwt8K6MyPsJlYiYvNOlXwMyTfOiMNbKs0BpvtpOjp8/Z52QovooSnVKxsPPKLtvYPb
xtsLhpqc7CSzl7fGwvYrNxWtvVH6HTDLm5x561XrgHpDTGYtDayrRFKqglod8nypq9qI0X7IFAj2
m1LVMB9EpzI+yVc98W3hn2HmIeuybbeH3ZGGhe8PHyENq3upxYyEjMj5OwnfJ07IxSIpP1EWDtp7
KRZKvEj+87Dj/7rbDfdnSnMrtxiBWMqCrXLWj602h5w8hakvkv0VbxdRc1sE05yVxS1XOEW/YuZm
JkjKgCLs7COX67wy3ekSPMxiBMjvNCJfX/mCYEyVpo+d0DGHIvBTFYL6rERcjTuT/uFMoSjPZzHR
LvH7Mh8cJpy5DaZf1uY3ZNqChl+JuOipx+lUbItbQPzESGwhQJ1whS8AkLjTXjj9pIUSswUM7eMR
Z5u1k3MzwFSh8T1+whJYIaZgc1gCM0duSVSvuXcmpdI5HzeGmf2IbLNGgnIKujMAKdCB0L0z4UP7
L4q6syvmKEyStgXFB9NJmelnhj+uuo2ogiiactn/69RIC5qJvTFBNhOKVEONVqrimRkWdksAZZFy
8gKDx1n8cA03bY/hARN4rC+3FuNEXbb/e5/DK3QcKD7fu43em4TDTttfEm7GwnGWSH34sOKtUpbs
GouZa/PI6G6fjUX9kjc9X3/FijZWTqkuRAlQFhBXahaLbyqxs4d3nNjYmlS5HUcUjO7Lb/s0eipR
yt+yuQoNJtszMMXvEbvVWv3V+RZR/dI8WkGASa7qz9Fn2/5/fWDjseLSU9xq4ORy92khHA+K2ink
xACworFDCwu2Qcb2Q28HJoxoE15qWwrhIrj1WY/XYYg+NBen81qEUM12JWeoyUmLeSDBPr5lVXeb
HN+xl00svA8uIpFnKbFqkVrdqBnW1bXMWfJwJTigO3u4qzOTqUD+VO3tl+L/qGBFqWoIZ/rMYYF4
bW7a3maig2uQoMVnFFulNiO4kkAgqgwuF0faLapZDq/AymVR7rpqZHXspPIUimqdkNO1SLefZlW4
KJyy8INzhEa1+VuFMqRJ1XymqfoTI1upX3DEQDSF4XCTvwgP0XTxQBpZ0PMgOJlFBFNnWC1EuzYd
GCalY8+vIICJBGUFBacNzPDw2ptcOci5UlywlNgMeXIdGJS1ajNjqebNfZKGc7BsIpktgC6U3RXr
hcFCbHOSRhgoT90LZHfEzXhE/koSic0x67DwvUgNIcH0T/6SZOr4k3kKNm1k1tJeZHcqBTUktgNq
z4dbuJu6Qx/OlUe0xamge0w+n2sh77GcJdYA6yn07LLFXKKZynx9crY0slvBhVo0oTdO9cHKrMnb
vm+Iz5EhzO9uanNVK4NAhDh+wMsPrpkNuMAUG73YM/82Z0F2w4kNdVPRJUREFEMLmLlpPgTgYG9D
FSgEkaQGkdHP/xZkqcozI8/GlFOqTRWy1UYLTeI+Uu1qoY+BOhrNwJlOyfNzWRBo7YKqjf320aFy
XDT196edWxt3QnmAg4oO39IpAzsV9oovSd5QETzQXBz2926pEdgzfiHouFaFS88XVZf7wOY3O/3r
qIFwelBatvqsqNMWdRL6J6AoTcMoi9Uss4csSUV4Yp6PZJmn/YSuBhIpezsNprx2G7uabzUrjbSA
aTPma//0Xqk8Ch6KnDQVmzXd23xOggefZSrefgXBbN8SYMXcR5FEbW4lg9GqrKkMYWyfp6MpaTmU
jOJ+A66U4zF5iOK+usPYXw2MwMCCUNQjnwdJody8k1otOWgqOc86zt2Qtlb6diaMs1U6cgMkNuLB
IRZnOkYI8YNC7O7b+lMlmTad4I9S2A6y7yvQDm6jxGSWbPOlfaJMK5rQpC3ytwBX+wLP+L3y/7aD
LCVWD5+BlmkCYl+VFo80hEwDKFlN/eB3lkZTCIaUUNGS47qHo6kNKof3mevzjTNoj3G8EiIoTBZ8
6GpctkAJaDUjHAdMv4tYVkRv13heQBFIeJOYKxs3lSydmwbCTd3Ix0RMTgzbnrP/soxYjxOC7AIZ
WkMu8yWhucWTTpCbuhKlMHbT9c1V+5mnEs6P3NBfackR2X+ePfBFyTOR7puiyeU6IjJTYSBUN3Uo
ylGTg4VfJgGGcFUdo0PUAIlrZhUVFQefSR8EtzTAziThvYtIKNaAu5vcoou7kYnP67P6KKCNjMnz
Mv+pFuJChYWLIHFqrwW/+kyYfwB4VP0vr8ibuwqwhmvqhnXsSu848lSk3+f2OLyxpw5OgRww7jqz
L3bM8HI9UFvikO1VdpwS7nPpOZzhaHXUoCqhSE/ZJNfi/iGG4ypGTdNQf9t2mVq4UuaroDAUZt/I
Qb31LfNGJ9+bo6tx11ZPfx/3AXfPFI5x6XSCLrCog1g1AuFocQ4mcPx5Sp+TV40RBqWvil0W2KeM
KD5vIhZr7kzQIvmDHF5kDYmsdkVJymGQJHSmowp46CoSIrshndXqDV3fKUv/M8Fgz4QJjG42zl+e
ihzKWC5bIHlJo8Tkph/ZFaKanfI+eyi1XdF2uKFBBDt6UVOurdlDDjVPmg3t25Mz8789Pzg2Jxr9
xlGPywf+N59j57wxTZb18UEzVFgHgZwJ8xQX3T3xzGY5h/fXvvxa5fTQQdA4Pxk4rHhuFVbehm45
Y441LVWvCJL/7hfADhJwKydvNoUHE3Oro0RthVvvrF9nWrccG02MIq1eAUXERbpl6oH8bXDif7qA
ZIidEShEKKcQcquiuxTJaSTwtc8b0g04uXJpLF9M0Do/B9+ML1StzTho6nkzn7gqSSczw0SBSCyD
TDxr3WS1QqtqOC8jNSyqgYepPkiV/NBJf3xNyvyKT7AvB+WDmiLPheUTNr8bH8ZJcYJeRna5hVol
f9joFLlHHq4sJmLpmcHdGQqhd5Hq3tk8y53ZTE0OOniOveIIMVhoBjv9TNBaJIzCkfoKvSg2zy75
/wtfmub/zZ/eJulH4WKGG5rHuQZAJhN1u9mH4nQAyeggfTWMmjWndj3dCC6/9sMQkGKPgp8wxyZH
cNpjpw22bH7bKAGLExs8fpoxAOjxTMM0AJx3hX1lbmscWZhgrzOnwNLNijbDYiTEuG5oZ6H9V7HH
oB6UA/9upFhzeCg9d6ddsP9gLuDJv+y46yZXYvoUS2U3kc2wkvS5ZKFYoU1eFVB++dnH0YqgOxvQ
m8yZ6biLpKyCQhiszPjyzzGkL4tuQTH1Foefr2TrPBJZh5iGicH/OZP1cYZjvqBhxkKxD8NLDqUc
ZFiLFlUMPiosxyHx94kIQVvjuMVF/uOE+/y5HYgypyzpnQSrcqzPHmX2MzRqGUWAFnJU8oxWRsdC
qNiiBnLYAy5YJUfLKspwBfM412GTV361XPG2Al427VflY/MMgz+Fu3SceI+lHx+JYilT4SryftMc
b0nD4PYV3V4rmUfHJziTO64le8naVQ+aS1DJp+y/QHd5WpPO0uy9KH9L1kqm8C+M/8r9yG2Lbjmi
eZecdbRcoRY5theqQHqbDMeQv2orGdP2CaoegkJyQv5xhSfuRq4B84mOjmaHTvbjkAW7BG+i+OJS
ngjs7ZzwbR5Gwi2AiPuwomOSCuaWVd1MX7qnQa8fk4viEGS6keRAeeJGtqQTba7f8izrUPHmewU8
DBfOrHpbjrox1xWrn98j904npel8gQe+6W0EU1EZpVoDnURqhjRQsJtlzySDoz6/uvmGZL7ZWO5Q
EvJnqCTVS1+HUrNML/WWjsJ2LXbAEKheGTp25jKEXp6WtLLajYFMd+vcEEO4TfpVq83V3IZA/+WL
iEihhg+/4GGM/cOGelra/hOGKmVXxMKTm6ng2jaCL05F1im4j0jt85yPWrKtGpC0MtIn49kF4iFw
PLE13q2fy/aORbcRYW0PhG4mGNM1oaKsehH/4BYv1miVH7ZJUdKpyUIPafQrbj76FxG0RtgmB4+2
kVQ0OSvp/m9UZt72FT9pglq9IZnanzBfdRctlxS4EQGaeLhlhf7sbrRAGNZL3ToZQTr7owDZ8gXC
rNBhPAPysdxRUbYgmTG0ZH6mtJs0JKuZ7DUTk/ft2toc/Qego0ZPYXqyAQEoKdG70HHCwtPOzAzO
TMfNetaf+DRODfyWvgBp9CG4q1bENKgaJROih5zeatXGB4CJBFoz840Qrburj81mrp4m94/REo9C
guPlOUWbK2N30gT9b28gTVa0P6blfRaLEN0p4cRS2F0V4uuvMrtNTsEokfO5GV0CQSlhfVRklP+C
OK3H2an0iY5aJw7gyun5pZ+vQUOQGntopmesGg/p5B+5yt1smWixMFpehId1GvkBxECrw1atjQvO
lcoYNdXVxlRh75yJRYE7feb9hv1A9JpKp3C3v1zK4vLdNe12dzqrnfpcAoYav9aRYhWe9Qop7Pfz
WnU3mXZXHWLIRfgLP9Ztpk4OPMBDx/COYEavajRf+cKTh7PT35pMTLVRfEzKuOHfWDaDXof8g4iY
EnPPzsEjDqxvyWfdXu0XemnSVgSFULtYjkMd4GWjBVFYdhLbyLKEnOA4JDJJbBf+0/aubqOmHz8+
IzOmrYeZvhlFPvng9jRwhzdamdeuCxrl3cXuoGFP4v3MGOAwi8qMia6exuT5qCLh8ByM2uJUr1Jo
hsCOux8pbVNKZPrZo+grypLYg0xbd/HzuHTMX3EoKe/Xp9wAJVXcx2+q5FTuNxUV74TxYAPsdVF+
UlCh5RFa8FbZOSSRtGE98TPnWbCV0ehu8Mj6OdQOdXRakGzsvmspO6tG8O/sKQa37HM6//c+bLm3
2J/26amjWrw463cHkwq5Xkocwd8cE86Bn35SYOfk6qeacK56kNm2hIB/o93ysI4ZGyIpzIAObTXI
N/Csi/SuqqXzX231Y7o6lmXQsNpSz0A6I75aDTV9q8q+355mqSX2KDmv6whvcCZ+s63uEvPdkzW9
cbaI1qZaTXsEkL79ODpUE+pm4W+b65HECZy+J6w2m2C9zN7HQPwgDKy52nIK2oQnHWXq+9a/KBvw
3boh3wLqtpp3CC60ohYcjyE14He/3vvwnnU0x6FJ9rL8Hfnhsk/oaHP8vUqWYnEl3FrC1yNGFanc
nfshkZGrV6/9iWo8pvm0cBrM8CWiUuHThHnJrm2R6my3g43JvLAj492URBCXuEed9SGvr5hIGEFE
EC0ovEbMs9aIsA8RrhWYpgAfP9QCjMAlv468DJayRkzWFVFl4EB0y0In/GVMO+NVGPH24nB0O21g
mkVp8zk6m1tyq+pTebTu0y8IWLWP9EVovczpt4ERJS/nna6MtI1zkStGiQ1he6swFDvf7dUDP8hH
JValwKt1nItHbDfNIV6JUbS59Lmn+uKSr/Oaqnx+VaRsEB8ZUzAcrxxWbp8wH6Hw86j/LH8Q2nCo
TdCk7tuVw4e4A2H2QKYk1p9eqnOVfjYpeFd1ErrYPNqvXkDx5YCg7DQAQiI9kIXa9m6i88rsR4VW
U5tVzitvRml0pAPIbgaW39OoGk9EII4CBnASmPhgzMZaBHzhqjFiVViwghgml71mRAyXbsEIh5jT
yadtGPN10y0hSmtfun6Dd62pzWYWxPqzGNYdMbWU5X4/VBJEq4YspWp4/jRAqdNq6yWKUaj9OljW
yV0QZVVUhOl3sYzrV1677FWY+Q7QqvxoX1VDMsDNC7uWE7AL6Mf9DD+wnh5fnd1e8+W8/ZZ3HQqC
0pscCi/54oF3bhM3p47n1IBStx7F9o3FDQQMNjIbS/84sxOttkQes85SIHbLaUyrS0FvmvqkoXWG
CsSLMFn1AFmx+CGPxVP5jb9FDls89vIw0CZUGmOm4a8AI9rGcqdr+8WuKYVGPl2X4DBqQmjrauTQ
VHQ1CkkcSGaK37bNAfJz08HeR1guJLRMwGsWkNDf7v9qSrkaQsZcTAQMVlfxwM2w9er4Bw8fYI4n
fLj7v4rp9BqNvCsL6n99ik6X7cZ0HBf8FDbCISdJKU5+EeU9CdJdfgie/pTpSowPs3FESQaGnJOl
0WbsqLcqsmBPxhkXL/GAqiz/lCJtJLn6IbyLClPYTEWWcRAlXY9OWSGDL+YLtO49POPIkYUJAqU8
tRtw1D0Oa08pUoGh5NwNcm0nhXFajzCYkjHjEq2uNn50paqByf7V0PQeyMmIebNOjKtGAZLd5GTk
kFWHZXn2nPGCxy+Tg/yVaE4dI1J1YW4eMzBiHz2wiCUWqvO1ezSz1MHansxj008ghDvhTWdq0UOQ
so9L6dn37/TS7SE7Ufebe+rcjugnkR3ZlSxOrvctkyLuSMtWQ/G7m1EJzdLOmlt4ekwxvBZ+fxc1
AMdVszRbAbvODwDKWG9XairvOlYBh6Y7TSEHJfUjfW6FDV8QCjL2RIqkDbGZPvxDV6CxVv4b84jA
UGEwYP3fjsayzzEU3iSh8KyPED91p5KFWYJD9x1rEEbi4lcUd0jtuy5DGbwUX8P9Pjh8Th7w2tOI
/K7zf2oWQzoMvKdZwl+dCK1nSqzL+WcnzZLgcQZhw6hxeo3h5JSnPUQ9cH/RNxuRMkmobZyHGGly
sKqrgYT2umNXXfGBOfSWre5WbQCraG/X2AQbcy/jpp5+EiVaDGnn/vyP8abwDMWCeCSw1He0/ZSc
T5Tj+w+MCInrFyclHj73q7aaUZlPYBNxUKUbOnYiw7tcWQf5ytOh2NK/iR1LH4sBCMAifZmIb605
Qpx/EHL6CSVyXotMTLvYWiOtk5DcXyv9pvKBxfMKqwBU2LDSN5Sz0EAGBJW34i77O/+5N3xn9mOW
Rrqt1k2Tv00A6PPkN8AXjjOZMHxtyMC9iKFrT9RTBSc18eeq3+OgshJd16TrvVoRPxn6BWfRhr3N
i+BE8kHBM5TUe52kZUWSlo+FiPWOg6D5GvYrGONhcP2w7VnvcZ+ZAo8yyRUNUL19Y3ohKi3fu1YV
SfWb3TjkPYagPs7NjJLYNxVjWxV2GkLSzIUF+d74LMsL2LesljXH2umqYBEfuD8a8q79ZdzwWhLF
DKrV5CS6QuDbP88bf7ZJDxWk0CTSrhGV9TR0kbtzpvZJjVBpIhH309KTwDmBE3+N58Lzq2D2gMzk
4b/EnkmZ++jqcxLc0llqTNW2x5bjAR7R1qO3/juteWwdifDOGYkICUo92iiwBRrabYY+LXNTdKEO
dDaNnlKgrOGZkzRv6IzS7EaCOK+LXkmAz7/Y16duEziOJO7Ttunl8qNyIg/zTkrWJ1JQoqBlwd0M
I2gGhYx3ZKs8G83PF+SFNsmQSvznkv1zvga4p+N2ZyrG9rIblMoSiCSmBeh5BSVWAcp/GuBs8RXl
SPzboszFdv+6VrURFmHkdA0QLyowhgRdJq1QmuRDmT1sXSIj0mrcnG+zwKHFgKkIsHTjk2QpwHLE
acs++mwVtfvL4o9RYa2PbHHKmRBMm0c86Wma3XSYINgfQcdFgPKvpbRJcfu0rKlp4TgUX4O5Y2YG
r0DUw7LI/NtwKQx3LcLVbNG3cH1T+jk28pIAZlJNIZdVqEiHgTHHOYOzWtwI9/AyPonBD+TG/Ny1
xLabiVDnqYVQsxfr5xxHWzoCwBprTJiGsLx6D3crA1cbGJuC7iVx/kr7S/4/m1ECa6nKbLE0UoE5
rXxfACBeQBBnAs0t4WqEeSF4MSBL6Fp4BK6djPJU74HgwTdrPX6LWNbgNt7vOK17YZMueXRTD1Y1
V+/pug53nrhEZRKhiusEXd9gS9PFVUXp7zPp6GGwdBK3jzrXo+7yupc0elSLgK/xY7VvIRQSeHUR
aI0iWNUTNMI/7Sg9Xa+RZHhtxoXFzdHAY6ZXWFwc1BTKN6eSf59gefhtHoEhgrIGvvTLs7UtB9na
isLHVGeSIHgXyNft5BgU81sGCrMmr0+Acbm9Aq7NCt6xrj2xVN8TQisd4TW4xtH0AWuYzyM3BEZc
CJegHy4x3Igj8lxyxdd5VuDTAVc5QB/SCYyu6/iNTNPd7vSmaU+s9sK4SfdIXdpUv2ktYXs40/+7
/9NXcKxP7Xc3HcOsbrzVhyql47Sr5DtNiohtYYELWY/SropH190HxBi2qabu3CcHZhw6oDGQDZSg
w+Fq4dDAhrl2IkShGYMZ5JYo04Vhgg6yLu3Y4YBsFPg6Vht08kwgSWKTOYiposBJ6rOhwhbVoJOm
1bfO3qPMU2sVcNgihC17gjUfZ25qxxBa8KRTUyUOpca/ccBRUcVru99I7GUYznhMRkh/s8orj1iW
bTtNbbkwS14cW3rexuA/P/ZSLeeAqip+1LSF1t4Tc0YwKOt4CqeynMnwDFcR4vR/157WYIUVwSxl
Bfkw8x2WyjFiwQH9GAZSAFrzduOxOP4wP80cMaOeXrM6XC6F2HgHX8frBxpdqtLvVROXLhMPHkhm
JjysOSZTgcB+J3FgShoCFs7wlARSzkeIPJu3VJOJqlKJ2WUurOquUr5lnZahGd5avcTQ7C8BmIGf
XH8wD//hm+YwrluIEpC80LQPImIdyOwf8Ew6mSm9ZobYxR/BdlutoXFn7Ufi8+uYkL+2K1J8+lZQ
bv5Rjx4W2xGpqyJpvTJKH/LmI/hXwKQE13ZYHBNDRhgioxqSaOif3gm4nkNAgDzSCjBNxUSnfHqE
aYvdTeeFJejlvzWGJaSdUySzda7Vno5dePyCRoMaILwv6uSvHwJYk7q8piQHR1i8zUisQrY/DaaU
yNEK07LluEvnWrquWmC5WL1amrHBvSAYp3PI4qzndMYuGim1i5OOIdH24gE9sXfwe6CSLEudLcsI
R6B07h2MSwTsUw854sBTpTv5OAEzU6jDnHJ3KEYKOfMHsOJdLQxXKUMeIiYPa9/jE0NbAsD0xtkc
SR7O0a9JqQ2s1kcExTK9cGd18kEGOORjUJeEvhn/4vQ24SJ/WhhhXhtT2p+oaILmcnACAyM13ro+
BJLJrnuYabSZK/EmCGo2PiGycn9D/QY+2LWByWyxh7myYJ4a37LHBnI+EPeVIMGfxTLG6X/qZtQe
/88DtIy3dTwGUqpc7eKo9n8vtLPvWWPWjbhWCcghusp6DUBh1s7JlDGEp5nKn6PUkevjXLTeCWld
F+zwL54G09FKo5o0NjHr4YfuMFX1qqwDcULpIg9EOmJoO9DPNGddq9NbIebufzAfun9/QN5A4E/F
y6bB/Sue/0re0YJwN07nwIVncviqUTvcrY1c6xzvAlTitdAPKY7pifwPpxJOlOnQmSTdsAmJufWf
Xwey9lPuRa6zvSLDjQYwFIObvLr3jHWA3sKHBBWqnuKlF2FZ6xZsMrPrYjfS6rPVYFXeLHv9XtvG
CMyi6OpFmo8xWVy2ZEGduxh7cToZ1xAByuT3kMw3Ehj8X5zvqjn6T1ObhQS1J3L5luiVPFjO62pl
q0OPmDzupj4GQmo5669gTN3KGsouy9ctBT2KkeOW58Q41Vd0eFt8k7ISZrNAfybvWAlbZsBT22zK
nGGnxsa6mxoHeQA3cLraWc9HGsV1hBKQfeC0WNQbZjpNphYnUXd7PQoOIo8vatD4iM8+hOuVeV+o
d0GtuudhDLtOhgRBRATGS9gn+bxNqq/o/tHLtE9ZVwua0t97dUKR+YFtqulMJ+GuDAfoWa16NyPQ
jwklAo4vVL//G3h1qGuYnnFq6P9LvJYDOdGrKG9jxqLjuiTIpzjwdcQc8LqcbXoLxz+VqIqVQvnC
Dy7pZfio6SG+Ft7v2fbcYeukoXcM2qtEC37J0CKO1Hc5KjwUlvLfKG3mBNUzCMaacF8EpALHzuzk
U1/WYUNrbVOvXExVfC+bB/TiYRXvv63UT2rfuwp0j//GsPsxr2McaI7GjOrJS6mi8yXnq8qsrmQ8
mQq4PbaKaCrj+wzW0zuratuhk/8kv2NC24w47alPfmAPUuLo9UsAaDJZ9Y8nizay9CQt4o262XCx
qU/fXTP1t3awJOwewSb8Y1y7L2N2kAKGPHxyQ+0NreMBQZyKixXjXipKGUGKhyXCc0h4HuoxrpKJ
t/H1x1HzpUS3IMH9a6Ow/nUrW5XQDeUtKi/qUcuCzl1MErLnevW4jR36ZgKjXePEeq6v94hbT69i
j5fEJPPj/urex+8OX7dZrKQKmqBjCEC0kNzxzu7AQOZnKnEdkvnFdL5S9a1i+OERREL70y0XmLkx
VJivF94xOD7McnJID0EzniteqMI6Vii2hdd4rYfENl6zWto/2PkDjUgyU6Y1gW64zN57bbaXgpfW
K/ybm9/1K2pfN18MhDwRLj13FPXtiCaGOCQR/9t+Xu3q7LsHTVjAAlNPJOeUsIiV1lSTZWdY7MqB
RUIXF0wEnbfjBBnB3V9/di/kFsl5OzXmf/FP0yPvhQEGmT7jtpFbCvhAHMWwP6JSxfiF1h1oIdMe
l/14eg4F9DBv92L05h3y3EN73qHWmV3VBM4iICQRc/S37mlXUmx9SxZ0ltISC9Xmitcxt+gJtfBz
68TG+FMJd2TfgtYMM27bRbL8B0dMezNfU0f7vRZQ+rmH7QkRwazy09YIvDH09ufxGEpQTNG4IeEi
77xbyCuk+Xn6V1A7WkzUG8vrAzNZ9xtSxBf2a8BcwVlSXNSCgy7MLwPl3W5vhPr99wor+TWg7ooD
XsaDo1F8lo4d/LqzBAhdnxlu4NPMcHcNZBpCuISFyfpIENq2LQ68Ppc+14qtMSaE1oCrJif1vU+G
0A+7vMhkbn9M/6IYFkY8uLy7AOYFNuc++gGUsWsFpJzFpXF6gaEXg7FpP7QYB4b3Z6HMyZWQvYcc
u31ovk2vkljMJpY0zGCoBacvmiKmL0NymNypDntthY8FDG+75bPN/RKlTEfhmlgRpXwcJx7mGlwf
WFerkMfpVDOWiPzV5zyr0BVHbGQw4LGA+MUjtpH0Uvqe1ku4f7PWrEnbVgs8AFMfisPfkk3Lw5H7
rDoV8dQpr8kGEjXUXT2tiLVQcFyp1zqyvb2C0CF9+hsVQWd+EiVk6VuFqWpJpLzzkgT51cDO7zye
reuRKp4bwX1F9t2vtXzzwcbFobwQopjdLILTy2QeapOW/T0bY3Cpxjp8CJMxW1w5jTY2NfWWtFb9
H61K+/61J5Zy5sLzFVd1Jvf1wFOeq4GxsjbGbvH3YJk4Iv/9Z1ORsGnjEz3A5mWCzFcbfCgsDcEu
I84XAgLyUuo891sKpLmY4bfDIRKHkJJcawBDYhic+B8YzYn/xhNaKIjCiIx/RaQ29UqR+jIBgZz9
dG3PqJL/O2jVuYC7yhzVD0d4T4SSNtfdIi+gL0xBKTt+CLvkdg+1IYErvjlBKk0j0L1cWrWHIfvO
1i26h6Y4luTXIyfMBzeUvuTjxTqmT6ZdA7fldwYn17A4N4oJKTT3SMD/2qYQxYfwYGKIWyHec9l6
8h7Oo/EqplLwU8Tr5O7og3RW4UiAqdB8+3rFCLRNyn6sYRxfSKRc5SWrxqUMwp+jBk6T/NsIsxnP
1cpELXa0P1o1u8Dq9/Wp54hCMfsgNVj9LkGgmsmS0RkprBsB70/e0gpIiCBlZnW0RxGK1l4Sk0tY
ijsSXIsj2fySclusDEP3UqYwPbpzlA4IE+Jb3f6wQLGI8YugsaGnGoAAgqL/3otIiOtkYPJV8jY9
qS49IKKGhIuzQlq/36Ua1pb7x4GBWSX7r8a/TxrHk33BLBF034FXU2ShAZ6OUuT82erQRuZLeghL
ZE/uBK4PyyAqpHpd/NEbqkarqHP/8ay3A873O//ec8vS/fr9sd1afba0TDnQDf2XlUirypzRYGq5
pa6A/9tBDv9V+3m2lFPTcpoPCEiH8VYW5Nxa1UxYmgMN3h+uhc6WPAQLw7j4HJAMMFZDk004eVPU
+GOMBi8SsQbfIW0b6KD45JL1obhXbGKNGGIIfqzx31s3Fj+ESurHLuY/kP9+Lg8xLZuL2v/PDcxz
oKYqWQVR1TqYnBarqtYnoieiY3t63ORFU4RSviWto5sSDGvm7OPew6nWN0wvmdFCaW6vOlQNg5A7
CVHZEjzdzBMWuiF58YgKAeRydgzfA2T/HtFxVe6S8G1r/lmRSDpic5ODCWnqBJIMCtx/DDq4W9Sx
8s8uuQAuFANtrAysY9cW4ecXzxjPl8V+M3oMZ4Kc4yjyTTX7pFk4HEN64eZOxAvBhnQp+5s4Fx6i
ECDGmjsKtbRHD6GD2YE/ZF6mCcnxAhZMNSJ8SO/duJmk0X+TQng+GuB/1D/Zcw9+siWhqjEL4qO9
ZsYv35qKWThQ1VO6IPQXtgKv5TX/vDy5L3QlqaLUukts9ukf68APUWqpu8DgFUD4TQutjgJ2LXKo
+Snbyd7btrzKaED8QPkT+IsXPcvPfd11GK/3insTE4xkklQigf/S/rb1p33dbznD1t/dXyWQr6QW
2v6Gx05ow3DIYGEsKa6NPNhwZguEzPZhjTspaC0pL/YnWH8x9UcKXfx+Z5eFPmYCYRAk0XZnVcyF
CqgXRW/QtW7ckFcpDxT6l/Hb5YBXroxg0XB9hkE9Oxs7t5PtF3LylmbY4u3YwfZd0HEsPAa1Yq5j
NW3y0scGmKhyILOlldRi3jqFFzYxWkZnLQkqyTArLM7wylJqlXpz4tQBbDGD3WEMgm8/LMKGcskl
3us1pGLMW8BaJ+ySTqDkw44DkNBVsyNUSmOYTbVelTlm9Mi4r43NdRE3chJRBCd1citBwNfkIwt2
av5JrA1972uKb++ES1/XdwS8YrMfxbzhSqrCA/KRqUJwucw2F6hda6gNpUJVLtPrU3zbZ5paXSSa
LXIL3Kr7bVDCOCHQJM5gbrGwin3qSONjOj+xVC6bzaA3KWmJ4GStsDe618pa4BTH5EZEtKzGVfU3
yBFsSSwghBkYWWSmEUUpgjbOFRps4vKLbsTquXclSUegWFA+4qG56AjNo3WFdCVmgU3WZStNcxah
h+TIRPEFvgVU+EM6yyTd0qWK+eYLEEK44DSYiGI9qJdQMoYnwjOqQpRxsb/YTdHGXXcC7hKSrvdX
iweUKaM4Ko4idSOb8ntCOd/gRH6M3XoEyJ/mXxnR2na1WhMpJL576nuRFe1BqGiNPt+9OF/3BqYQ
H/ogxcCjxK+eSaKWvtRJIi7ChlRoDJJrB+Wvjr/nxG6neK59oTtcm7zSjuhk+WTsqOYT9WiMuin4
ZF6fZ9Uo2gD9Mw+ivXCyXHptrO5x1zirjYDBHJvB52pFKeeluKVU0ZtOZspGtWrwfRSAbirZ300u
/w1ZOEJnPCn4C3Gx6i9y6vQo+9Q6HEt/X21FicI8u0M5ntoEDctd2WGna/ZYuy9/Qq/BRLKf459t
C2MlMZM/Jx09I12KpWgpu6ZWWK0CB/8jDH+XA6KFi3uYDTuyD7SbfFDzypgbL7v+V7BX8wJaM2RU
e3LUdKbbLSsT9FfadCqFnhZNhL6yVfwJEXTN194ZlE1CY8Tvqd5uq0oiLalsbe4hagzi62A7fuew
FIGhZcIMnu3oqYxgWJRDLKOl99KCaTxv0JI/S0kpjH7RxSWkaTVllqoAL+pEov9IPk6D/6srC7SP
6SW3VixpPLH6y54s3KfVV4ZkiNMdsELO74tZx4J/kUAP7dgpgFvJHmtHAhGYHkhbr/Z96VBMjxjB
WxHDCDBVMAh7B9VQCwfXHKgHBdZfUmR2lJERJDgyjBmXBar7Y3PRU0oxvfuwB+m2UIJIVebpgDII
7CT8h5QKc3iPgDgl3IqrliwJJC9OQ0PdCFPF9/n14rVe4gNUpVeG6SFq0Afx0gES1SaLtX3F4dgb
4argZq4scW+0KrZIf4L4+Go+uLWoXoMokKyyFgWO9zdXACrWwd04QQCApicjvkDv45+MowLcYKsf
DPyNKoORX1n5ROpDhHXfc1sV3VP2JU5+kDJYvlrD38Ingt9JFxhqRRpZ02O8TAlNxLU8IDfZ+ayX
uSUY60Ef1kE8MHD9g2l/hzL3UApttwVQbzVfzXrVU1a7cj7KIwaksOtEpvZdEyPPyg2ruUFC2pjs
rq8B6oxIxYZTWr2/e0htX6X1+873bfv/dln6I/D0cnxBEb5q++s3fu8t7CO1YQrPzhnPhbGx5ASt
KkmcCNetK00sLaBsz2TqP1Qyu/3QyIEKRSsUTa73J69wZNSbDJpIX5rRkrearfZJ4yDlglVUVFhf
0G07qSnClRXZy6nY9JUtjPyhSp3hf9HS3qEJbgA+uhztG7MjvBlhHwdS3uJLFow/4dF5SmZpmq9O
Em8kxxjT41RmeFYvBTZ+d25NmSSH6Pil0822T78hKZ9CAAvSLM1VHlSw2w40+AyteyEcRAWotcBt
r9yVxDt4qdVGci7IyIOS9bP8S5ESSDVkcoPEj3JZ7dUEleW2lTU8/QSsSKsdr20LFiWAs5omydTn
wpRL5ML/s84NE2zUzttSB1Fg5XSFiauNHxGk8rps6FT+GjbUC7K3+8SpIXNOtvedejftt5tMhqYG
Y31B0CJYYQ7tN/SHxjG5pTNRQlfFLHbysu0ESIUuYVYgqpe6JQR3kQbeQefkcKEce9pvNzMFE3b5
ySaf9u/I86wS3boT60dbYkQyAcUzenMA0LnbqLTKD4H+mIcJiV04OaXPr5Aup9Wp0hSrKnGQXTwW
VyY8OfJ9yCamdCsA/QN5loth6GMEyPFH8wdGDsuZXEVet/+MzzTCeoWPF5vgROAjkri6tOYO3TBx
kmmpmgFmG+dTKvi93oWtAU0XPKrC5p56UBWKcQRgMxNLYNcVASjb03rWhBRw8be7EWjv0Zhpg1My
Im0n0T/Y3FDeYL4y9u/0okKgoZBCyYIQeIzxcDDZGkxs9Xgo9iX4q0Fmms5IF3Cgfx1ve9plg7aB
brpmp4oj472IR/u36GSgqNgH3SFGE4IRUbPX0R87cVFblHkBZMiAgJV8m6Dbij71VnIEBMByL0VB
iiyqoKKhp7gHf2RJwEISEzq8kY0HbzrEy5AwC9lfsmgHeNRwi1TnQV1Lge/HoJIy+O/Aidmb1ZkN
T5DslZyLDDYQCTKJVuONZetp5wpwKfHAU/9QK6qv5YXRVW09eYq5R+8lc8EByUEsFoliwaY/FK/P
0hXcKFqvboLiCDGoDCxv8h+DMU0SA661eZfmznza/8EA21P9oHdtqQw/Vyq1PT1FCvbr7Q01p1vh
TUwJ0v4oSJsfL8iDaO6vavvv3LIn1pMtnjGD3kYBl3dIwj7KWlHRvK6d+Gb62Ljr0F1cYsyuKGvB
SVjh3Ilc/QOUZfixQTRIwEs9X2+Fn28K+CkaLDfwxHXV4Y1tRlC34LzPqcX7iqJUvhKziuso2isB
rgdZkDmdrq0Z43cbZALkvrGaSOPE1V9GtgWvcRywmGzp8fA1xGGoPWnCaxsBWgKkY1wWZ6Ksgb/d
rsb/a2SG3va1cIX9N+38n/C1EjoaYYX7OqN5+az9e3+OiSx9iBRYzevTcyfTcFZd384zDRzWAewL
YTm46+ZV/PZiDc09ulpluBF0a6Vyk/0nCsWc6W9nDNG5KZV/DH+i/C+hjka/zJZMC3rmAqvp+Luy
ZtqA6NnDi5b8RtlGaGHCIMh6j3kmlvmCgpggT8Okxj/so4T5bNxPRfCryhwKFX9CiCVD7zNvuWbW
75lLjzmFfBR+bBe3LcRbbzSZjrd+8rurqADiJ52ZUIQ+hZqjuWIrksfCmouvDIVLqlY4t8KnVCfl
4OkLdaXJTIYOjUdI1P9jnkdqXvNPfsYvAllcpCyZWgi6IfRFiqj/MT0tZ0OPPCJbAhE3Bi6CEf8P
R4+4OmnWdVksYi2qYhZV0ajbBN2S8xw3Y6IIpE0P/4P3wcp1ANx2hUjgKRZoyTccH5/ZWxXMcUKD
KYxK9oNOdMHuESDMh7B0RbxXt2vF0t46BpQoPm8Vk+Ws4TXMXm7VHUPnLTsMmKSefwYhUl4QzRfu
aLTK4EOFxe3H1e2sTFufhYwOu+6m8CYvEqBhJSEi8KCaSEutY9I41ME72En7n1ggWi/cbImTAz1F
Vlgazt/3dbEk2Ee+ZCLv3UpfiD7PkZZrbRqANG8Xq9ul8x1JvkFcstWAKDzadvHQel0hnI96bxJn
eEuavXyUgFdlZr3uVGEHpyItvbhWo3TkjldHm+3KNBQwabAH2a+heIneu+ABzR29ndnbKAeiF76Z
8ifnIV9/xbIUooD1ooBioCJt00i/vMRQEORYspm/5OjZvC4P8dBox0iayJfVWMrJf5RWJKooxNpB
hiGCmbhm0IQsMecOFpf6fy4x97V/wJUDL+AZ9UMVeBMlcEzVzio5zqLau1Y6NMZEpc0w/DfGETqs
3T+ZGH+xPX7qQGa4gN1z3OC1quHUPeuyn7PD4CaokieiUQ72gClBlvPVySHyzSNWRe6sxLPKjAhH
uC16C0utfsakXOlRBp7q50fnRqUa9F3m2zvkAMG6SIGJt0r9h+HOaWXSL6ZbtIsUswLs43pFpbqq
CtVRK1npnFdh8mPZfWrFxHyOR7ziLpattUGt3JqwX9o4m9W0G4/QZ7w/2NfxjdHd2sSCa6vXLD8b
hXYGOk3CAIgaouReYEQAA1/V6xUy67bjNbIWcW/cBaeCUjTiLhZ4ogJLyUuFG7JtzxmX6Q79S9vq
lSvi1fb/5eC6WAKkeDK57mhpD9fEOihCT8ZOoTv95eppbtL6Tgx0CEsyoZ7DLusXRkQ4F1xxCIrU
duQbYtK61AHmmX3SrqkfxBFcQmCtF9CbX3794xAqoelVNXk2DfAzoM0bT8BtcFOsjldOambfKv2/
jaJhubSAYPR1PaRapWsq0Yc72bVbG5vNFuA1g4wLSge/yqnklBkGH9hzPJuSSZH8RVAiPeUpCAud
FmQnvJDUQFhldeOTq2NFZkYSV/mXjcJ7GrWBqqQArIq3UalfNnUVcIY6+ZWEsp74D6FoyC/5+LFv
4thN9QElyKy6WFwAMaRo8OkBnxIkkykmD5xqdHHdD1i+ZL56Mrdx3XT4iGiNr5xs76csLhRpcpjs
wyVH/ARJz1PREYP3EeM7pShwYG01xfB9ZP29u1YIXrtghUrMsb6BjjLojZ9sp+R9FT/VmLk+6qeu
uRofrVUQXyxW4qMkCQEfQj0BdV4WDv6DCbCdp+8djgTQKhg6aFgRSilpNXpPtTjm+q4Wii8lZObp
+r9jqD8+VkTW7soeMSDu5nkq2PNWmlBxHtuubViuLCCmRXZ9dlNYkcM6BvSbC28rsMCHA5y96iMN
mPmBztnsY0v2O/bUqMRVH1GfRlZ2QW78oG+IlPWRN675a6kWis5j4likAFkxBYBrkSnmck9pzO5n
J9Ya1NboHa9e2f9x45PodYFtWRd3NZ+gmssQyraCUMFcb+QU+6GKPLi6wvNHYtMq+x8P/3JSvWXO
LJVF3zozw9pv8RtdHu85Qdp9WeXzw23koofKI2c6wX+acbGLIqzJRSFae14pCA8b/ODc+fFbIbmn
bp2Ry3MXqDT0wFA/xYZZtorXv/VHM1Ssd66PZd5u2MeecbapjMes36IJoNgk0Y7ZegvpDHboHkE2
osmHJfkYkqSQKufZy5Ml9jqX+oVm2E4nNi+zppopUzzcbUHa3GbFwcSo+u0dKhfX2v0MFO+PlXOP
AOeS0xjk7kciPOhEt4BVoTEpy2Hy2J1Xu7P2ZGe3EDWFZ4V1jmYlBuxxXTa2VsJIwCrZ8VBbySsL
3ZVfBkaSCfaYw87BuC7NMWilXgSYaq04a0I+6TE6kSzG9zUoOWITRgkAySBH7xauaqGmooIUwQo8
yuh3bHrqX+TlZFRDC/8IwyckNLt28AJMTgihIxpBUWLs6IUNuwSek3kskMpY6nBDVr7yA7aP8gFb
rLu0uMKiVcqjwHmcWaRn/Sh1BbUMVAlSE+Y0IU7jV5CaEOtzqauKOHriuEHkstLWgjiJ5hTBd1P9
/Or06O6KOZYuOaDFc35DIZ9aP3g9JRc/m42HZuK4/WjyWJwhTeGH2NT4jhkrgFdyTsraEI0k86om
PnH24rDQIyauOSazNQ0Nj6A767/qZKvFoiXc54fWJ5ILgzGMOQiSEXz9vWO1j6cwcgONcFmGwB2J
F4sNOWJaMZU2bZNd2Q5Kd0I1kqkJEro4uMupp8jSyX95Hiu6s1y+dmlYb/h64DGRTMBcrfQYoIDG
iuH0muEdUwMc9NVM+ghkV+W1I7ZrAVSC6UovP3ND80LQcPFxTF9H7XERJaQtQWwJYoXUnO668IhJ
IAPYP8+f+FqOmG9abNNh3G59NLAxr4YG+J7cajgVkIbQGK1ANu8qiLUlXnyI9GRTjZWe2R91zVnC
ciYzbFjsMcXV+FZLB4Y8x87YZUPdUvgdM1U5HreFEY8IoVKlN0XdT2GJ9aSTtzTPplNMmzVZXEQM
5GoEOCxXR6ncW3GIjTRDGXZ8+Dne6GsXmwEtRV1sz6eDYGrzZz9ET4PvkcglmCRZae/+CL0zA9dU
JXs6wwHIishT/ndD+3zUBeHpRhcID1mslYUep0FaHAENNolygBQBnTYXv2mIGziPeejikYdXnwUb
Zzmolr3df7vES0GF1yhtdCfigVSXCLd0n9p7qiAyLbgYLXsr2lqqemAhEq/CfVCKJTM0ZgwPK24t
WRb/22v93rJ1eTr/5itCFyfzMqdOfnzEw5HX+yUGgDPvLnuInw3MboWRS9WIuTtgto6QNMBIpgAl
NmcXxryYXju3IAO73QxQ9GLTnVWvXRk7Q8CC6jvxXWK9R1foJiXc9xb7DFSj+zSnEiKLz9tBq9A3
LEfSc4r4wpkhhRf/1FNkWTT6OGkiTynvtbxFFETkiEXYjB3Hw4tXUTT9cSYI7A1IBVwXvjoLB62q
Fhjk1p+KnXcsupGxuPHsbPq4js57zxGm5XpRCrCN2j6CalGAg65yTWJ/E7jyCUGwIwaCIovMzpUs
mswqARDsdaTv0yHA9TrWJIOFCdb/kBdDrpIUzeT8Y2vpKFfVgMKkcCJeIHHVZWcyd+YF4o4eBfic
gSlt/jSeIkGTxCGomnkcStGDg3bNirueIdnC533Nvh0eLIq59T9uM+PthCt9L8C2Sc8uX2KAJbkG
CacCmDvy3/tB7zqPoxMyHe14aVJH5HE1BcbzcCtvbffMmnaTNgIX25LiV3PaTjF2GegDm47XZY/Q
+jwZc9rpNDbcd/gx4BRmF2nz/QMsBOh5nFDRn9fp1boUwuvYSMlkWPvIE3a58h4/e1LCjWWU0N5D
xmRInTPkPGqxzHsDxGpBeqD50h1fW6d04sl9td1+rVozRrhkJ4P+A1kxAwiZxZEncKgQ/C+VyaLp
Du21OE/t3EOXwzoKluNuLeokyucnU6D3qFg9/cxPN4V0XZcU2cg+OemAue8ot+TaDA7ha/rFWdcX
1gXn19itInbN6B6kDY6uSuKfrJ8edcxFAfHp0iW9VfBbNVPDgUB3iRVx6vaOkpeFEZqOi5P2sq3a
WZCXCr6SX7FmxJCJfArgwvBu/UNiiFHo1Num9MzeHMHVELBPLWEDEg7UhSSf/Ch0q3o5PMeltB7D
Clwl1CaUfjsSWXSUkKaPJ9dh+Q7xS1cX1WXKCbj0+FpMn9wU5zCrwH75pYkuzSjQ1B2oibNVRWOt
iWT249kmde1ZWluQv95EZFHhgFMX9faAK/zAgduU2z3UBf4M/h7xab+75fWj1eeffqQ9uZBOaaEC
9+MsDrI7UaJ+1xxUKh6U/DglgiEZ9VZeNkzeaKpxO0WZNc2ND3zbwTPKMr7wyRwz7nTZL6w4h2Ca
+//vxbt2BXZvOIPcyraWkvlwIMoRBoOoNCGltWXamMo4c9YyTS0kWQML4Edh+YbM4FdGn31i8UcM
ooxhFe2vT/eoknKROrhhmO+vFVG9Yqvjh74t0F0sCiTPej1H4G179k/gJ8ajLJDak9q20Q5966oZ
19yWD0etXtOHGbkVDcaJm8mCxPGb+TeeBXO4nmis7V5C/VBO0mJrLEmf1bDMGoDP8eECwufdWVy3
lo0vCkB/y7fuZyW35Ea/ZCzR6/smZpLxinWo5uXYWOwD3+4ZAT8qJ2wRyyntnD3JLWVjk2yx7OWY
UT4kNFrJNHJJIsD6WnP38rEcbz02HKfzXi4hc6U0p/qRkzVS55cnbAGSYDeE4umdKY+iliIv9a9F
ySFR3ybzPyB7WqM75k1uSq/lWAtNX3LaxgLuA+V3D8c3NtF9XDLWtmjCX6BkFK/9P3I8bxDEFzbO
GzRyL16dxCZcoYJvm7AqreqPdLQ9DUHeKxuZ6HMQ0wgHnIAc4YfTYRpu3QXiAf6b4wK4av7dV3/I
NIxAmat/1bGk6vtj43a9NBKhY5VWZ26wCCWGbJ7Ls5gHBSpnOjLNWuIM7xxR1NrFlGr6/HwhoEmr
snWtsCGnUmZ9C32z3FXTXyo63jUavSv3om/5GAyBJR8AyX+2MYqVUyc9dphqVdnjjlHgrVd9LAGz
+8P2at6ZsIhgqx89F4P+tU3/DGVW2sEWtnMwZ/mCAdHRApnyiaPt3F3mPq3amlNIPgsjQ9ZaCny7
HfPh+6thCGXTi6De42uT5Q4J7UbtQmkmB0b8/69LiF/IGnXG0Wv8QgADYIAH4SVEq2xgyuBo6N4M
/a3jFU5ORchtR6BxR/pmlo0F2FTEVwKmAFumP0nI2ZgLaW7alDfziH+l3tMW3Zr/CTerQlwvI9Wd
r4Zmo8qQbkY/ggqk0zprpuo9UnFQbEVFy7M5SrRTvD0oHd4jobA5Tmr86ajbkys7A7STIo3tik8L
Dt3h36a+BJUnlqWvPxgJD+hjh+D7bHYOjLjqfqqcEBCUSJu/PAeVdkLHGIYnN1ZSiSno68yXpWdy
kN/OAJzkzUJ34n9xhx55qOrIKMMWaB6cJHyHiXySQfvYEkxPVnHHs1N27JdHyW4F0pVTt7Y4A4V0
zIzYj0nkH/vB18jzIfPrdEx4MZhq5bNGWoQsD5QXvM7sdKdHQaogBkBz14D0KAei9+uTqZp8JroU
DB8U0xT6z++eFtUXi6kbNgrPioWl4ei7gfBjfR31+/mUE4Jm5j7q0bckCm1SF0K254l44tPXNEiE
tvdTACbvAO6Gtb8453sSIkX0i8gzhvfl986CxxKVd/oKvFTxncRN5ygRpyXeSbgKCdn4xYIUK0Gr
RKHcg1sLnpwsaDZ5cmNik/ex2IhBcqi6JWH1VDiwShc0nTXsffiZhq25H4GEbYYmCulqXXPR7vWW
+yG0BeRuSFag9JfkDH9NgckdqDvCCG6cH2wscmpgjfAv5OWb3qOhoV88igqnoHtT8iPIuGHPBLT9
sGEG996ZDEmbcEZCvvq7ULbk0Icfk+7hhnWNTVO3RvyeXHnt4CrdjiiFX1kSafJTWOf5kQsKUa3D
DPEt1N5G9Ud1ryzsxBTICzG3A6hTsAw3+smED2pC9bZ++E71BOqHGW83+lHEcYahUNW5wwgPs8ex
HGDld37BgheD8H/+TaxJPsRP2pjvfmAk3Khzt5shh/IGziDmnX1xrbZofvw6RQmvvEvD1L9tCHSB
DH9/8fmNOLrNocwwSQfMqNCiMa+dZSjNl/GhJCKeVv36dzR/4uX/U3VeKKj+/1qqG9o2ube+w0jN
J1qDPUpyCObeHrvwaQy4/qeTqJg9HExCwjpH4zjkT9W8gVlhtzEbVg52ejB3SKbGh1gU/zDr4n8+
DHO4tNABshXdff7mTQelR0fQQTkLeUXhKF7wXrGlVJ9B0w5itbtmczu+T7sOGMBAMXt3PvM243Hi
hyWKuKBOYQmmf0S1pcnX0yAxgIIHH2hyG/ET8AfP0bfhl9esCFsAxgVQFixZa/4BMyoobtGN8NPd
VAZl8g97hZYgep578u4dNuDwlzc8ub/TxUxBKSgc2tXd0PyWF3kloCBkt9cHKS54QsDiUVFTWic7
NpjIpPkmeyOoQI4gJzXmKoj2Bngu0dnHFxgaB/Pbz7r774bGOYEEoVUgTXF7zdP7wqS7dNSGuLGl
ls31z+KhDerKJocY8VeGnsGoWxpC0rh5KjdLv0mmlGvYsCfSI2U22MPOGlcbjeSMPhlHVmFRuHmL
u+mbQf7whi+RFXMe+UHDbjA5RWxpM8e9DoZaT0j31XAx2GLHa1//n1SVF82DhRtJrwhedjSlyKCf
91QWPLTRyPXTeLou7KLhbxc+nFZhK3vV9VzSjqMlUyfyjBdnzQAcD1mbzr3knP/peCk4Zmk3lRcy
kR0zp6VChyIP3YJPCpZUOWaz+ToMIyM+Li+3xcIgHIkwNcnSRyE1CTDIItL4G4VJQ1KoHTq/sXC0
fM/5Vfndyf+0Un2tssCdrLiTO7Ydr6Ilp1vlMrQnISjeB4VqkDxvMp7KvVMmWezyNzuOHJ0OcPNR
XDJydeiWHFKPQIBln62yfVBnwju84QXeP7zotjV1J50vq2TlSDKTPLZIKNTyeh7Xkfiwa51CekYn
3T90SBGByLhu/oiXixRVrVN8Rfa+kZQx008HT9fltMSv0Li4k/hIeo4f+qQv3xkoo4nRNu6VQ3WG
eM9SvFhJAuc73z0i20hb3d//a3Ao2hluc7jzD3T9xNPBQ2u/hbO9q9irSgSyT+IUJWMlYoo7TGmP
D1sZJOgvd3rY0UHDpACYoAgEEkWniG6N+dHnyU4BEvyI9llXExbNhPcWx7yUo3qAEb5zG937OwsX
gEzHZDr3RUl762rY1mIpgaVwKAFQd8LJizFFUTvqT/G2i4d++FSr2hUflqFWdQooaASQI5fON3Lt
f2HGoWZTD0VDJyjMUp8mI8i7Yq+/c/rIMaaIYYtrvkw6B9S/q4MK/ez6gz6waGHbU1iLy4C4lMID
IBJb+x3XtQRBGKByKXNsYTGFJx/3tbYV3sKFjNRMn7pRdL8PudCuZFpvyfR9ghUHhS6P4UYXHT7S
muB+yowB4Edo17c1LtAcHWBxBa6C3ALN946eyjuJf4HMHAbhjsfbhRuP8Ijy5MXxJ9aubVx5d9mJ
zYYnngaRbkVhHzlNS8zpkO+W2n/s/+GI7CIXLV921jyD5tspxTpO90TWXvvI7unyTXXfNNF7x82h
vOT92WAV2/mmmaRJgmpNyu6acT0iGHIj5DgirERoM/mL/XHJ8/eqHB0J3lVO1ciDoFEhfu3TQG9Z
5vxO3qeqA5XX5AD1h9zcvDXjGyIW+hSieps/xOnJ5MgQJFZRM14wwpiqmdnD7pDMFrNy2PIRvZaE
IHk3A2LiZFDoq4vCLOJYTLgbXwJzRW4KYorlWmWyQgDWOWdaEeocWj5yR9rqmhoNRdnrQFCDwcPz
q2+jGR/D1S0sUhWO5NTZpeqIZ822rTSuwWbYuFg11Ma5+Yez4H8POYuFHCyZjH/NQDadqTH28wkg
VzYzUkpOWbesi/11XAoB6JEPhD7ke8bqsD9EfFen9ibpD3nV8rIyq4cCfrpGcrbY0+033AP2Tcj1
F90roRCAaltGAUXguw43MPr/eqk+4PW0YrJ6UK2nJT8ML0M5iTcAX/LS+XkdR9IiW5kUfzEeWR+L
I/K9de8WIH+gigXLY6m3W3b0hOEKCkByxsm62XnkTXZoO9Ut9kOdn77ELg24VjZBmHp/VB4xxB0F
2jfI2TDyj4YSjQO1Tr6MiqSa6LjGNWm5vEf43VOA8vP3NCTPpTQ4x857a0UH1oMV/1CE0X/BRVh8
YZAcTniQ9jKfvkIDqnyrO2wU/QmKktUpRWhuxCgHCzDwaYcu7uXQJ88ns1WP6n6ULeNwP94vdgVn
8SlxN3nFONjTyDjn0+/dJi7r1P2XDGAMhhwfZucbfkdVuHazae791IsWVVsCILqwp7cMyShIVZmn
PWFZslk8d9J66Lw+55p5XIz0E1g2cuv1x9cfMw77G5IA9NhmxuyopfmCr3CtSSKRAelu8B81zVMY
CkfY1JhLbBYnIH3w6EuFQB8oBaxThjzeD7fAiodnTPGUjtSi/pkOKOfHVqgyHR2TAiZd3WHqNFnQ
tKruVPgNhdOKWeuWHm4c3wTPRgDQd0ddWf0Wbp+f4ISx8aJQBn9kXdulsIcFyoI2RVMosIw1xhSw
1TthWvGeDRneOR3VIQIoYP9KoV48qrSS5whBvG6faOYZdQTP/C0hgwkkwMxYMcVq9lvnjuF1N/ho
U+v0v4bX1GlwhclwIuMY9Yvhi0uInIF4aq5posn62I/3nz7I5OlMc+HKjOWTtU/cvLl0zJ9pjduS
FMPaB0rP5cPq8nQRepf7+AxPHw8Rncno5FxPQdA//sDStU0GKSmEBPfMzlsfpO/h8ZBfc/fFBtZI
7O+OGSkJdikyh4ZNeIV7YJH8kZ2TykpbBp/sGLygsvwnYomJTibJZ1rtLL05SEB/MObmzL1Hf8hu
GheH0x6MmUa5RSYCMVPIDWyMAZN/XAoZFdRq0mzuaRrYXyNW6Bk2qSi7L4V/8N2QSwbXPWJDP09z
uKIs6RxqHLgxVYJGXK1pF8eqFnpSrk+BpN20qj4i8EO3KDyZg9PLhzN4sLTfnONmcZIBZnsmL+Tt
esa/2nirbyhnPCrNwAyNXh2HS0PCHHrDT0dPN/HWM/SH2P0Nva9n+TNb+6aIAUkOEZ87aE1SO9DT
c0BC/tnDJA2LyJluAccRuBKMEhB02OJfVMH6H7wx0QOGpRYi3hs5R2gNySA2ZLrdCSDwymdj8uTZ
rUkCIq2BWjwDu1QctjXmbrfiGeFEsTPP0OuY6w1n6hrLoTo9MdKlJhU7ka3qTN7vDDSvxfuqQePa
HtYDGfnPBVeVrwoR50/idU4HVaXTEOYC5s8ML5ybvCqdUbdTUTXY+Tkad3IW5gZj8+dAfCm83+9N
z9ydQP6jMiyueaHM19sS0noqdKHew1sAiRYPwA3c/WIIjN9m3O+hmHtD7RoOzElDGmI3G/InblgA
4yaBQhlhdit0oq9WH4wJJ/KAytO+w51SGsE+18CGy+nKtmjuVYAd/CMF7yZViCxYsEPrYv0wtf3Y
oa0NynVrBWow0jKYhossKR925n6SnXYelcpO2dL+Vb52j6Zp70iulbBacEqpBAHAOyOw19I/jko2
BF0Yrs/q6PzRuPfdsWp2HQ/DO1oyasT5mXS6/9XKn6AvXgcGHM9f0P1DqyHENBdVGl35aMVEplM0
cOHq18t40SmaUxYtA/EA6WAOmnuFaugTItrRyyMmT1pa6S9zJ0LiJwfEe8jT7VqcebXy9NWRur0d
/c31VJa4fqSP999tGjO2W1SffEnr7yiOFTE3GqS7L+Nt5BEvReMUbJ6HHe1G55g6Pb8n3welk6aE
SdnFe2lPcVfJbXw73ygvH+0orMK+YbEPw71teq9n6nJeAi00ANKyZzaMoqhBkrgMZBNTukimabhv
l168kFyymrjXE8MQO5kQNpthVUVdlm9xAoPEp9na8CWDXKmkmvkZHfocF9pLOIDwTJaHPAMawmr9
thIEhho2xjtgyu8C/KO6heRk983C2n/0h+GXg7xruGS210jKwU5GmgrMp3fjsyT59scGFk25I9CT
N0PYnxf1h4ZPuc8DP/vTKrDYjaauk3L1KpXKTOtfOaY/hYkpJ9ylVILTMC1aMUF0soOXvlCaid1g
rCIVKaYIdDxPSOsOAQ0NblXKbaXWVc4h7gVDyrhY85ZzZp4nTrgC05zjVNicgubyvS/UU5FdSZiy
/XUvRXIFzDWYu6/X2VB2nupZYOl7PwhyQNMSuCrCdg+kphVS3YjTXwvBbm2s+J8CNrZg081xnkoH
qMLlFNsjzpDCkuJTzaLjrmXdaEMfjHwUfgAGVsLoGN2FDfbf6Zm6oosTnZJvMdbEBon7AhTLaRu2
As4zR+f1PZ5H/i49d9vttKlsrT3/vsNDTXqF/0UGQwHX6xr4HULVTjExRGV7+LxfVf/rV7vcDeTU
zPy63JW3aHoxvOcsO6ubf1GRXYmnpL11HwAVcxRP5YrJDsV4o5xHoYR33RvOzL91nLetUlfFm3gb
6bgNeW/EAf1YyJFMvPWSkfziDA9M9aKkThLitImXwZEkucksAAdQ+Bzru9LopTZbeE7RFWf5yXU5
BCPHZyJ5PPCfRtq7FhH8RfNOFAtv++uKjj+ZiU7PimxcluxZxtumG/eraxnf+doWoyk3xO1yIodT
EUn2Nhjtq5p597P5vD8e/Mv1I/OP4aKUQ86MJcN146NUxHH0rmzwsPG9hE0NR2mll+o4kvO/AqB6
CbQAgGQ1sMdtV4l7UhRPOkIELVHzlUDaQa6zQTqdZvc/kVUOViz67bCxrSxracVfIFf962O1w/wp
DO8Uq0YT+j0eljzwkvgdpQ2UdJsKpwG02dVGkzR6h5b7pbO9Z9Nl01pl5x/BpSAdlaM7ZhLjOfXA
+oe1ZUVTY0e7nzDAwSQF/9izJYsql2xKCp4b5JY/uNU2WkwibVgY8iP7oNaOh7T1b+F2/nMCApjW
ZBud9PdjgdDuUzSCKLLacMMF8Bry6POalBjrGQXQG9lBvKPoC6qXDzmsUHgGtjO8T7QMAyo0UGPg
nWpv4rTgg+A4fU/S0+NoeIWVvO0+/palI8kasNHUgusTrD7ENLrUhmirVbm1RML6BzWGMn1iH0wX
qbG/IJy1WBStOOWuHmqLl8lHfsMW6YVU7G/l7DgFAUgv2GU42BYf2uKXgQDB8wIkLwNtK7bJyUZM
As/7wBn3wNQQYPgqqkiZQwH/v83Ybqhq9IWHtB662vAVMovhZoZP/RHTKcA1JdyuxJ2e32hx4T28
fIIkIjxUzrnUE0HFQEtjNADzot1CHw0a4pV6Ah0MA0c290Ij9n2W/JBqHgqnV0o87WIiyx3/XdVf
qbsFR98f0puvtp8B1WGntdn9W9rd7KQm4P4t4DXKQr4JFmzrl8EtI3dLVSqV8TCukSterxxwASkU
1NmoV1NHOQzrNcBzJEp3Rn/CaAo0jfN8begn2/RjRwxvpPWkdYmRHPOtevi/tKNiCuosIpAyugjv
UfGjyF6BQqL4cMO2MmyIEkszbqQvAn6NbrxgY42xaqBmviW0P5Z2gQLpw1QyHqHs0/TGZoc7D+Yt
s76uD+ClhValNe6jThsezaQq9odtgeWqGQTNs/F9pmkqHW2vEnyLVo/2YCOGMkYesHLQ64+2WMkc
nPlgQ8d6pOf/X/i0GRofyz3OU8WSX9ByA5fbkzh2DMKW2AQ9l1bifq4cSFwCdyFp5rsbWM4qEKUr
FAWCo7pck6EMoG8s/6Fc6C3WEsclrQmQTP1OpewQXTDbSzLrjivqktLShNbwh5aDrmIKNXki+tfY
Met6sNzl5l8qI91we66FjsjhfqvZuotO/98WIixguKJW6Y8sRmeZZSd8I3/ICTTtOsRFTN/WLvDF
d4nUdu/OwIe5NeL7niFZY8XbxmIo/AGJp20R8mYEpD6VIvCZMxdPxy2Lj/wpDlPBRjzNZP1cwl7X
L6xNtuidmqUFYSLJ6igzV2gGoVXViiV6u2/38o20nBsr9V3rT5ofvqZy/pHK0UJEpGpIyYRgUWjw
Nz8E1jPnOrXmLCSCqdug9Q/MNUgBQxPshb11Hd46ONnU27Vc8p33f0J+nE8feE8pSgFBFj2WaH2S
PYH/ghkqHTNjTKbuCqoDv2i6tQmhJ0L0BDCNklJXa13crdUH6ZzlM8H0ZZjgO39tRcJyx8qxX5Cp
s02hoGfqnCJrbZSGbYSbFLvLG85EBpgPAOpCLg9pUerFIDg8TYc925tgBddhxnApmt4lYHAocCpl
y9R9Ne45SSyDooMHn13dc6ieY+xxCshitKSoIjEOrwotStR+jr/JX4GfB3Olewyev3ezvyS/WKPJ
5I+4LkK1F5NhSKeOQKc6IJ/FiMXWN+KvJ8s+X6cfH8DzA69TXndFaDGYrCdLkauGPWUqLx+Lrj18
P4ugeEtcMexOPuVKkgE3ykjzhhj8HSBkLfTriTp+LNlUWVsCWVnE9goUZCnvUH8jdfXccoFxX8U9
bzRjq3ToZnF2qpTKeiZaxeYG4sb8FMfUD/XGLSeGgOlCTZ/h+tWxT2CcrGGO+G5NQryvlQGvSPII
ixTWhVaiEghubUQlmGxNteOKhYm5hQemKZTJUuEdxq/PfVje/JOKoxid5U3uiURa2K7T5ynxOhg5
QJdctHyFBfmVnnuWJeHFgik+VDqN71mRi33b0GRI+8X00aICCIIiI5tfZMOk6LoCBmAU5bXdk4hE
1CidEtV1PlVx87gAdMi613+7niZOFWwr0AsHPmEld//kfj0JqHkzt4+W2CJTDLGuQL3MCDs5BW5B
cE3t6p5VoP6eK9R3XT4/J8NIEYNUAZ61ET0MMgBnX/tWOUhts46B96GTzH21DG3gw8XPVz+obDj0
a8ffXJejgNPZHPE29IM6ErsFeC/ywNqK3fd3cM/DU/UMMrvk4FKWNBQIeypA32aWtDfZ0RwSRBQF
jRRuPffn6ARGWshobhiIsitVARDL9uQgxqOJ2hhDPoF6PelToORvFtl12A5gsz0RppVoH0LUDUVg
1eJYnDUA6Jhopn0ERvtdUUu50ilFpfVFo2HHkVO6XN8hx3gH0gjBB+OUB8RKmdEtBqszS+yqedRN
+hoyfmyJp5y9b6eUJGeiswpfR4JFMEH9IWnhNyttlGOPpwDUmOUVmt9ItTf6yee8qMnogK0oHyjP
3LZ91htWX7q31GgiWT0vlkVIlNADQA5DT5FX8h5UHpK3z9OANH4Qk/uaLAsem1cbaxRL9ZBcEB8g
DflRs2MbqwYI2ZmChxb8wHNgJHQbHCZHciIYI6wuC242ol0LeoE7bGHpxkjcTX40EU7EobeLcqty
q1NbmMfp5AnX4PYxFYq2/DhQN0JeuDEBDqC3YmYjz2UV2GLj3u0TLBjWeL5wBwdC8udLNfCqzbv+
HXXlv2g6p34ZzozigNJHSxL1+yuie++oiCGv5OhGnqJDWmjVzeaRfnrX9k6b/K7DzfFPGhrn2fea
TcPKpAV/iUGdx/gM8sv8vh1S6lB7MF5pqe8rmIqKqB75elS/P7HiX7vd+IOA44z4dXKt+nw6S33A
TuQ8KlaSpClLSvtB5rUYx7kKYuQ7K3VyFwBcZ7lW/1WNRrZCmLD6tcd0lwEhFNGPYhCvzjiJoKf8
IicBWTw0AzgbcSlMgHuTpBkiSJ13f9OsUJ8V2v9ce5XGEgqsGQop8JdKHBtDMnF2pWGFGR38LDQ9
MtzKjggMS+XpFVTU4k3uQk8yziK+dccpdMmT6uc+5lo74ix2n1vmEk1hacqohPA1QNGMVwVBXc3P
K/1j1WNjkj3drcBmuViv4kGNH0ELcu9ZVwFAqBCpp1vwEynRG3oMFdKKAV56BJtq//bBYNyncgvF
0MMattrJdBFavHzA5oUtT3L+Zi6IG4w1ul4klpLlllsUoH/I8mLdQObK/vX7rfFyNfNB8vjmJln1
cfbuEstAYBy95rq+EICd8nFlwNmXrSKleG8o2ldZ9t2eHkJ6JgGYQA3yt2isXKjdbsqR78YLQjix
zhwpm4c+ScEvZK/bStPTpL3RlaC3z/0wlJZqJo472yYpQddcRn/RrEjxHyZgonymsIwUVWk1ormZ
0xjN+Sv9wkpWf62hXVAY04WzYbFqI8NQ9qx+1afGcJ/U5YPQwo3I90P7RO4Ooi6ieqKtzZfUEDkb
k2BLoi0siamwynCDpXZx46K163dU41XESComRj6d9W9fsiQIlJhg/IoIi31cYe9kCy0e+3yVOBuB
rQFpbRMWhfPEx4eXFr/a/Z2/7eONjh6B/scfJJXcoMNVWvH27lLeWKMPwWuUcH8CLyeF/zz8jeRg
pwbmcXX9WeZKpjwOrK8y2VyTYe+ETkNkHcFFrSnRRCEt4NncCtQw4rFSD9nUMYuu1VFwqAS7wJAs
w6cWA+4rBBdv+Es5S07rXJx4Lv14iAsGG05xcU++Bl8bsKiPBONmp+UGnSlDNVJLSygwZlAnL1cE
h4ya8yaXVVwJiUTwF8uFwd/XQenrRC/eHuBA9GtRWMofGeIKd3MX41XfLeIWEswZgsX4oiNoXvpG
bKo2R9Jvn+E47HqI03vUorpTvK3NT/zlmHjy0sZCEOB6PZTlXJwIpkxqE3VknCRwvZtwL1y+BuVu
MmLEdvyjBpxVq/syrBHAmaajVqTxNsfn7tsL5BreSkuIqOI/ffA3qPMmAIryt4N3naq+174SZbA0
OaG6jmdT6u7AKMwJRZFJ/M5BZbpeXvO3i/pQNnbK5lqo5G+elWEukoLQ7F6p6iQQCjkIankFjofp
6LyClC+bzVtzVzwmuJZpAL9pOtbK8Ll7IMvU9EWtgTvilZPUGJO51PZniU5mBbGIzPnuaSS1EW82
5UjRLusVCLuSUNnJr1ji/JPOh9M88dq6xV82JR7Tscbff/LxG8+PL+VCaTPmh+ysbIw6HdzFgkB0
e2ezzTyXH+m29A8HEazVKcyjMNbzlx2IhVYgtG6Ws6c82JTV2wEvum9TA8VRENj7sgb3ip/1CzRx
kilt7T1vsuYupEpl8H5bLdHwBwt/2Pf1giytWM1UpnRlt7BTCeNinRpzuQ0rFbgyQM+3b8RP51Yg
sDTEycUKoPs8OizWO/0cNi+X9b0FwnBo7WKJRlOwwgvwK/lrCJRhFbtSg0Dl77IK4kd9D/hO26pD
zGYNrzxUrgD5UFHYm1DJbPyB98AVAOhj7RSFOEZMK2jsgKT8twyGiphOPPlNSAPUBSGOrjl+DFaT
hRr46EqY/mwv7PoIV25CzM4U6t+FmgxC7VeotMUAW06u7iFE5MY50me/q+2i7bpmbhAKptXSWSik
ROgC8YnWpzVUsdSvVyjQVcSWckPqimw+GmJsUfq7YzrAyQFTq5dTM5rGjRUGebF+GflrjtwCvg6E
jJ5HDwwJjmwryYvTe05vvePGvdh4+8Ela8akgGWEYI0TssMCGs+wI2S9qNMo2t7KuBjeNTyoGRf1
2xjGEH7PQAc8v3SAJMIf7gp0KpUSzAFnyIGyXrAnx19NpJp/HlNZLmOaPRRjutgj+rwyQIl6+unH
yHi3XBlTxHpG86dxFKNXcPsVRnKBLdtjjYdix/o8bWZkH3JbYszjyLK9iiYIctt/5Sl6s/n6lqT6
B/gbA3kz5zZYglvWg+D6ge1BlCcmwnDkA4uAySk+13ba4irS8X8zrSPNqhs/QZJXuUTAhA1qQpli
hgvTyNCiIZmQlNpNgRqmKcWct3tTyPy2Md+Q/hWZIRoI8W5yyA8r7LqbpVKncKCVG4FmPCa6iTIT
7wyU7XEsY8ClzaOYALDsThZYkDdi8AhIJXndFNtCS23+WQ6UUn8wPBdp43c/KZoQC42ZBFqpmZH8
iUUGuTkzOA0pMe6BFV8GnPGK15eIbSophoY2pEtVMocbsezMHrmMmdB0RQEUtvW1TIZCrONhc3lN
H/ffaF9gIKtHGUmDV3H/PCrP/0Sf2QZyVNKM3a/d1Kb4xzKyZfxe9J/TBXIHoy/ftp8PzMUK9Vj0
1gcwj8sQRqI7r45lVGDhO46uxiU26Cd+mgBvyOhsi81vbi8Yu0PIAiKmdtrp5XHtJTU9MvE0dOwZ
nRHoETpgiZIa++ycVqggfelwGx6ruulYnhe7qWe4gQGakIo0I2D9ZhyfsCzhDrWZrZCbsobMGtk5
y0vvAio1/ucmzjkd8+XJrc14pCVmXw+ZfaMrlZSV80kURXWvQp+ePJxYV10ewvrwQo6q6b0oMkik
co0oeDIWfI7vdtNJxmR2V3/F+ANlydpwq8R+JvHpWXhjdAi46qoFyQv7v2wTssiYlWKN/BPG3cFX
XOhr5tiwIAgQpRwYKSubrw4guuzJNNgyYvwdBnCJ6Jai8liDeom4HqQmyaPGFKf35+DufDe+/LqK
pf9FeG0Ag+kQegzBJD2hYzbrdX5lg/6dYQ3DWr2smUaOmkbkleZTvlSF0ARaADBqTbFvBzGTfr5A
9fFY8HZFANSiezZ5VyUCLDZXwWEtuTmrmYXXj2MHSV3AJkZ9WIFbXqr77Co70qUDtevZPMpW/khT
+LXYv+dfSxZxYVs2Gy8o+B0SPS0EyDKGOPjkWC+qrULBTG4DuA8ruhhwAJ0Up910Ba99GO2p7fLz
L4AZk7fXood2Z5WeT6bTl6jn+ivFgMxHjBU+greZNg05algX2envKNgZsHyZKJj+HCSctnG1rdvd
bxIxUcWfPesxCAdwPJ/3ZfBqi3sVT3bei/KokfuoxLDM+wpsOK7vYtoO838dWcSoupv+V0jAzLO5
rOv4pnRSBCtlyAlyl5gOEmc7pDlUtzNtGLJZlDQwNUIOgMih7+J8VBpUnq0EneVdVenbYWZTB9j7
qWRztWgSBXjeuBo2HgxzuoDmcGt2GdeYDpyHooSLg9ESpovB4cHJ0h24CBneiR8Ve0xfEEV3aurA
Laqab+eah/cqpFWQTViV7O/werk1iU6Lfx7qMU8KCzWgNg+3QYWuQQRX+oBbY+9XZbozXRUKvJB0
H7wdhcvj79zLxr48uI15fzHYA290Swbf/HLNO8o68l2ULLxGBojUKBFOT0vCurGO7tO83RqxlKd5
EpgkfMN9fNboPJvCXnZa5j/DlI1j9VmOz/giUkSulOqBGTMywfXD7JUxOxu/QuE17/eA0ZT7Jdci
CcOOYQylnGTgFxORnCGSXUEYcyle3dkKKkoPe6B6KFx+S/Rt1OlFRzlTR4MN/zB4eHXjAQ/HZi7I
e4yTglzvxUhgRTdjNG+0KPUJdID0+OOLeHOl8PbXC2I7lGOLNgTf9QLEfIYMgKmTAGKq9EX30JUN
9fVELDoEEXi8fqyi+fdOMsV92DcQJzQWUeQm5oYglKMjCOZ1xBtoNotUw2iU87+wa/I2FT8alBI7
VoNjdZOhF8Y9msmX/uo6jbX4lnZD28EJpauJjz0K++kVkPDWaBOTPiQjyl3VGi88FLYU1UzJiAvn
MhZRCI0JdJojef1PcwhHzqgw1YheXL34f6p7LdiZLie1hsC73jbvU+l2tl3h2QqjMG3oYCzm8hzG
0y6EW5/olNJA6HrMQLOe0uEn7b8PI6f8qi3IjL+ouV1E3eUr4qax90hURAvle+WkXJb4BSqkybaD
gLeybeS1EoIDBxnRd8tDxz4BstqB3M/e0x9Fs0Iw9R4roiGhBR9oryyNeLq7XGb+j/V1uVqweksv
X6c6r23mkJVmsobMhEWKO4/igJdbEyDo92EzXbJhBA1KNK3P2uKVRoUwyXWSubfvk+5IJrcUqlgE
MKcG0nBsyOQa9upiaWJun9getI6ME1Co1vCHTFO3lHYkBjuv5YcrYEn1ewyuePyU16zkonlAQ2Xt
z6v3hjEQmu0DJahDzS96oYMY/+0jYX9lkKtvGbl+8F8+o+aBHSGUUwRC9SPstIif8j2YDK6SmDJx
QnB5VPg80vZcW7xu3fFJlGnmaTO//hnnWTbOOVutjljO4Rp3JNMwbp439cq6aBzd1KDXSvJhXcgv
zH42Y4ybWBs/kDCRCXHrTxva9n5v+mrSm/iJxICaM9oxQ8ojIbN3bNaekb5FGasV1P+iNtGF+xkG
64CHYQdovpFMNW8PDKyGcddQEgTUu84ZUy7CaKNI7KTpUhFj8VUS9RxAkg5JvCz6EyhV1ivc2zsJ
KqH310bTJV2hwbacwJjejKQeSqIuWb2Uo7vdcj1SGoIxIFpwILZMD8YonpohT6uZkzPcCT6/QHO8
5d7HBMcoK3s03FJmk67qvuyqYW/huXrVxq19BKWnWt1i+3fiSkAX56f0qPspzTiaVdWHTbbZgew/
0QA/jWf7x9Z/HCGxCV/f2Y1bNdXEKYM/i9DM9j3REodwuX+Sv3Q1mQUnfn4H5Xrvjz4P5jin2HUB
Uoy1C6QsCuHLmOGCjjbSnXSCpJMJXqgatcCxA+CeiS4em/QmOqReD6lAd/DUlEj9BiFyWJrXueI0
mXVzsuhD/6J+7IzzV7JJXXWWzk37pkwtmVbAPJ8AuNGTJ+eMsd/2gi5ryruCd5YG0GILtQcp8Okq
patOXgBIOsTAHco4dCcHxDnmRu5/04gMpCJF2UUK//FW2l0DWJZ38fXdqP6P98bA+R7Bg1emnAg9
xJSMTNBpad+GwRifvTj2KNNp5C0qJ+Z2B90ihtPFmp/vGzytjW4gLT2Gu0LLCg9jT8bc4Z7nReGN
Tcx0JD1w7cWCwFBGisjcASi2ZLSA8XPUXznV8qqSe0RT9sZI7pnofujZa4TIdYg4xPW9VQR6987n
JplnZ04rwpSGKFo9GztJ4Rs/nQXUQmPCtXO08HJHKH0iPseBpk16OdPYeEJhNqnzjsqfNvqex/FJ
0ZLFRrlXqUToAAYh9yBBzU9bRPfwT9jRUNgmZOgK0eTsswhAkJrMTX+dz//yKGAfaNCK64jkuaYS
/9idEiRo+ttJ8KOkoTKbZ8d6fHZxOo49/EV1l2vGhMzM0aJvoIQDKnrviYhWeqsZIt+EG7COJ513
VDg6l4Q26zufS8D0Jqr2NW/Jsh25RX//t8WuWVm8RTnaB4lOECsNcMTjjy2rDQMa9xk1Ssxlbr6x
B4exqu+qr/pvOT1bYHTDamXzObtj8XtJ1L0x5Amm9m5vj5aJuCNlJBi+GBocYsys+5/MzgK+/L78
/2FtC1D25ccDVAOUAGo3/6vlgjOTknN3BGvfl+rjMu3PCqAY1wb40Ucc1mZGU3RsBBnNk4yhPmWO
Rq72oLxfwB96rI4mbzrJo77+eEEAoIw6+XCGFHF2liitCOjiMPeMVt+Z4xMQ+ItwJK3yljKpDzHd
oOxz6v3EfrJO8waNj9LnA44APaIc4vN7vZi+ehMjtFKFESUpGSmq/KPLwdf3ZhXSaaShRPHeK6wa
xeFAPgkGQZS1d5nWHegOKnsCOxZ6SwWgGL5X0yUp4JdjZRN6plHFkmwePXBp+JqA+AgMkA+hNGiV
QhICmKkj2WYVhJUsRtpPgDQMcTYPdQTdSpzlUEkaLM8fzzafT9Z2fp87PWQ5TAKRIyVREGlcJLxS
YKUp6M9D0jEC3v6/rVAfhczhc6qUL/KYh5Pa3EL2hVCNhvczZg0+Py6eO0lFTxRNZOhA7pHD2GM/
eorKp2ldhBYRS0kp0OWfK2TOp4BbHmXtStzB7IHzpWVx8F7y+l0E0C0uKATZUjoNYILelem0NcKb
M3XFexg1xjqs/FTXlA3lk320JdaDj/rWw9wubIm+vLmN+au9HyZPF2lYYNsf2IOgDm2NH8bICAqJ
ds+V/uWB9BauhR7nbmVQ7W/m1Uj7GRkm154wiJ5+hf7ik8a+saswTKWE4ksUCwKhzaPDCVor+25u
aUSMyWJ1JMTIG68+bJEAgC4ssitXdDA49QeK1q9LhzOAI5NtVXhtWJ75AvutJbsfRYxt7bg/OXgc
ymMULNIvpwIvvb8w5Y0qJ6JaTvfiiByT5IT6vACbHfLfboDCQ8zwDjxdlYocLdqFRajBQykGUash
rfQRqtQKLLDhjbzmKaHLAojWwmtqRP6DbcMuTgelkF4lqkpbwNzdt9EB/0eCxvd2WoB30y7pXXkh
AoBBZo9XV3eX4mqn+rULh2+7OK7UcFlC/bRIrC+gTPn9WdCB8cYLpd3/zr8vCVNgbGEat8y1pBu7
IsPJfuURO4CPAr6td8LHoly1s0g2txMkOlYS/O09n4dGdV1VX+lQ0ieGweZfASYzRi3SQC4ylTJs
uYPmTGXyTnxjBlsKS5+jKfNJMSpAWuStbM/b1NqxNd4S4pIij/4BA9k/zgli3rGxY3LfgKl+W245
19ZJVHNw6HeYbqcR3ajaVWNJsqjwJ6BNt0G17fZMc1ZLLTOGjWrMAN8FSvPSObU//MP8bSxircYj
V9u4yGVO7RuAn/9EAmlZpVUjULkSJ1/6PSUJBfXYTrNkh073PDBuIiFyTjOMwqm8liP8fKBIg0kN
t8yLWjg/d77HzlrNnVhJqncuVC22T++AVZnutsduHqMu1jrmF6MfjLh7YLtl8tw/Y1zmVgmG4lM7
RRsjkPCnHQlm4hPYnNhBqK+9+ExhkOzOZ8Yjnn3+lIPWERy4uyJdlmfmXPPFfCSxIt/SPo24Tcr6
0Ps6DVczka4RQcMTT09p++7nnOD7vYAw43Km8Y9/MrRD0fr4oxUTPLCq9YcRBg5Oo0xR1OAPraav
OrnHldU/WHnD216uVeuHpq1C2ic2d4eSOwKeksxDBf1tVyfY+Gul2H2CKgOTP+EUObV301gYfM17
CoQDq7P+Sh6cnOaaDGDMJiTOqX2gq8H0kEA5FXzDLDrZG8Fgv9WT6/Lk0eyLhDieVuF+kabzgPbC
YgwC/SRFB4i5c3nlD1O6yicWXU7qN7m5OQHKFpb1v2/eV/ft53tSdGgjU/MbMDk3gITyXMCSYwyd
PWvF8hUvpC9EnSU2RQDlLzXZXUaq2T+lrymBxtPDZ9gaLTvRA8wKLYzMPVYkVziVtLqIg4qKlZgt
JMuP1WHxXGk8ybtqEzLm+cgJOTwobxcmMtiZ5e37IB56Dwblv4s2lWr9Y+k6g0htwPXH8SYtSn+9
2bogLToyChi7o4oIv0+5MksMPmXXMX7i6ecVOIJc1WyFmaIW6luAhillrMr3/nUbMvChIfgT2uXe
M4DNARABRgFifIEBMvrvhWm4exsgBe674ndB4JI0yitUzbU49upQaNxU1bGIOinh+eDAzmZYUIp8
pb9MJZbb8jOv3nohKYsYgulrEAX6aT0E14D4jXDT/daGD8R10i2nzaVa6pNhioB6fOBaM/1WsaBZ
WfJwN7dehBbvD2RhqpAwq7TxxNPAcSjmIBhlSdL6g0XuDbVwHx2WJmvDKgMf0TEfFO1BD3kP+b9N
vKKG2nqKjqsT6z/tDYPtCRdfMyKkxZUDQiEpQf2Msm6o9j6jtVlDfNqBE1RykQm5igbA+dI5tLy2
ZvgBmrKWbwA93h6Tw2voEdMmHV9O5PcwXF2+RzRnd6IkdeV1E8FRXQCKVsOmTekJYXnp9yNGScp9
35CGXGH42cYbgzARekUj4B76WEHcqYX2IzriAqJOCkRXnao58LGTGFSqFP9H0hn/yv+mAIoRN/Bg
9gdZd0fUwc+tNow6XTUU1KdCrLz5xASBEOEzKia4dtn8njcIUHkV7lqjAVAyyjesaP9SOS44bD74
fRppD6tyAt0qSjaRjkQxiVdfH2EjhLRJMMfriYZYMKV4zqKe2HRoaZN+ro2ulijWj7/+U8o0YreU
SIrZIvvOwHMwzx5DiHupmEAFa++I8aLXGAIcfOo4+L1aRgnxsm9foM4wfMYmyg3b5N/k86q+jBH6
0bihmBNBSj7X6Hx3vXyH7HOfX6Dat5F5zS6Nt4negU9iKHzBNJ0P6M7M0NbwyoRjmSd7PM04Ovmk
MIrTQwovcOgHglzzUAUjYK85laOB3+ELHGyFuMlOmId1Z6M3Bk76BNymTeZ56001blWjUYhzc23e
10uyRld+us2d7L6cBNRqVWQ5JdoSvYmaBwI+UYKQo3BKdsLU/e4sSzz86t95IAScuCYjSa5ZcTc+
KIG7NHwtca/hhyxfF6XIBjRRZY803fIezyFk+SUL42fcIxFe9u5U5yuX+N10DnFy9Q7Ep/6nVSqn
Qc0BEYT7Ipf2s9UmurxZmfBc/Ps821n30Ig9jtWB7/mro5EVETdNINaTOwOf7VpHzayBPlnCAk4E
VA6qihRraJl/u69kIt63MMKv3Qgl9lsV27pIsVlbCyQAB4cZMx3W/32d7oqvkssRgO6tA9b5T3WN
31Om4obBB6z8Dpb6Zmb6HxVDc7Y+CRUAkkaRZ2HOt0M99JeP4B9sI9YgfabsJIhhNKrgeK782RPn
FQu9ShNAwrsUhbVCJUug7MnX2bWaEfaFIG/s1A771+YtEmqhC3zXmwv1m+2wr54J+jzRKOUkdIiy
eNVjgd7iCnpegp5gaaxlGK36SbDXXMZt2eRIwNOSFiTt6K+xkHtXfNO9i0UxmOUbJVeoZVvBHlTa
DJvsNLAH4LiFw56xxzqp8/VbQ1s0mYId4H/HOul4KK1PjlooI/AmBlDr1jVZsKsC87HsxykfMCSa
oj4v0XuCQlcmkeNVhH3iEjRwzCYv/a/wgoIg34wTemxEdoejvhtrEIvboiwgQNJUcSn3Y4L6q4Wj
+9Jkij8UDLMMZDgd702DXJlVU890x513aC1vVye1Ng7a8eH2aAbsxKe/xMeHhkRj8PkH4Fgk+RcO
cMGw9cWEHLI0ug/5iDZHQpeGAc18/d+DVEuuPuVbyubLpACE3ZJoYTMJxbmu1WbjnOh7lNmUSbDp
r9zdFYnYTSxtJYmZVS0qU4SKoIPTd7ofQVOfGY7i5isS/XfVq8qai8P9ZnIKhybZMsmADboezgWq
Pl30u1HicrPerXS6gqNXdX3mUN4iAvxcJeKoVjsThhV7ZO+AthFmM8v6WeS2a3vxhnEeain/noQA
TW97v6pWjSCzOkulwTm9u2Qq1TxdM/+CV5hbGEhIOEJaALiV9FAwF01wNcgK7f+Hlwi7C/OZ3HLM
iZBgmJLjyBCAr/aln/ttuy8/+M+LyQkpTpgT+vVG+dcyaYvurstWVZ3kpf4N03POHBc8b8ZkJJBw
UCvrQ/N0/QJmYtdjsLuFrp6lZeCkc1XWvqGlS+Vb1/M1ysiLIyyxbJ791s0mwE2DmP3wi0efOuzU
qdklDDde7mIHn/ZEYH3DrKjTpkKComAN/3I04qkXXmFdH7s1YooU7CGF0l1Xkymr6x9CdGR21cdg
T0HdcxlHdS4RqPfUDjy0LptQbsftmShmFEaQczHa170yqISLl6JKNIfk3YCmyOqXpqAyFs83OM1Q
ofo5fa6lkxzMzPc28IB2sIhzHWGdZ4MG3NwoXFsrpMrm9uY/Hws1V47o38PhcTWlEv9u/B99d30B
Kh1lECDEXXP1uSfDNJvdzflyXiK6HiE/YV6vJQRt/lf5IQuL5wzuHUNfZKsaAzmabxvmT3hdF6KQ
udRwS9+diyeSGImQkBBfmk2IUQ2JPqjN7YLL8Bv4ZbyMUlLSBUHxzEK+mSiuU5MEDVDFrIiekBoo
4b8t0nH2hhNIJm8NEWz8xbFPnebCmjtz/+DKWe2WJMg3Y5u93s8Xdf9/PYUmQ0gATCLEssCitmIL
cbECZNmVhFcYP+0KC19vyJQalGpqIeICgSvpM5GUy833hyjZWvmv6yWNocQJshvww0Sz38C0kbLl
K1MPJHa2mjG1QZYtW8yCjLZyKcTGbfPIyDszUQkzkSM96J+ocBLgv7w/oeBfgpY0oxCogWO3RwR8
wSdVjfWgg7McIKByaDFw4Pt29k6n2vOotyrYPMLTAAtA8orbUWiUsphr6uZGs8Hxd6EkDfPOAxIO
Xic5WvutieLKH5ElyxK4dWxkn2VbpKCq/hmPnid38Ll1TVXCbV2hJ8HWJul3h9oFcz18qKw9MHIs
1WqfT5oYdnznCx6CAZyZPtaE9jWhVvN03oTyKbhqXjT27R8YCGbt9at69KzHxxM3FyLalKiJIMgt
xwZ4tDn8fvgZh/N0aSkY8oz6cS9p7dr6x/K/IFw7v8nAcnWf8l1qohoAYEWJfecJ7V1Vh+BInhBf
Db+F/J5wFMliDOTTJ3RSTIkBBFdhUzut9PfumBPQWC8iGwpR40y4OsjTEkM7wxpg5TFEZhF8G8za
9Tu8YDqF7EwwhibrEsLy6HMH2HLUA9hUFjam1TTSdcNm0HoWjoCCIOGiYOSgaDxEPzBB6PV00/wp
qDRXa3m4xbj77mRBXFsupEzdtp5XRca5oQ7Obr2Ezf6nsJdiWzu9PXJqsV73jDecXHMZyZyS4aQR
q8PVAcQ54liYfXtLaZ5lYhJphbvRIjRqCvOixKzDP5Vz1katHjICTk25zZnKTZ1mqAMHocrSXZ2x
X3TMLc58snivKdeagUsJgivAkLECa8lXl5F1Qg8H2/TMGjmPk+Nm23ASgo8lzhMZqnwqIy1wezke
2Kv+fugBrFqdV/wGsSpOWdEEQCcYLol4SjcpE6P7uW70WAmO+C686tsUPnXPaaf9TJFumMq0HydW
WdjoY/HLQKdxUKYzn1FX6LKbWqGO0lM3AOpFH84kC7WRSq3DsUf7FQ56qS5yOWTc19ac9PXW5gh9
JhBSO8iSsGVCd/5uf1PP02zuBYNPR64j+/NgyjEnTa/bouFEv4QDh2p2akkoVBaQBobILy7WaDrV
NiZXFrbaiOPUXovUp0SPdfzr+/GoXQ2hioBrRGORdRATONMCIbdpGsmMK4zdUlOT7nu0Yi/VT8qh
gaZ3/OGIQE0FJF1+kTZQKAOh0iv8O9CJN0JxUvCfF53nH65/eees+ARPiuWLg66TYeV6r3Yjd52S
UUykCnSpDpJekBfZ3/iWeOj+k+HK3Zonf5jIITDi859u2nVHBF3se2yXP5KlPOD1lT5tsrdtvjBY
tcvoG9V1gP3ylpMSl+Rtb3DaWxd335Hq3OdPOurF1D5ISfCToS2qF73LcRNo/uyNecWNjStsZpay
CRwiIs4CVS5MCpOCAZGpA+X76FqTo1teIoEz3LsRVxDv74RKU8XVB2bMQ/LHrxqfZjqT1BXDPTVN
guBFCurs9YrB45oXdIxt2ei36Mll0fu1M74eGwRoCff3QPdLias5nTyboTNoyLBR9xI9PkHl9hVB
bAxpPp+T36gUSH0oG7ktKbldR13Wzy2ROmgXMtrY9VhcSXABkyuGDiG7yuyxaIVHJahyH/Fx1K3c
jliL93TCizqZipvknUIjvvzsM7VJfSxaxdxkuPZOqKJu5JqqsYxRt2j9kpRDDF09/JqnT5t0fqPv
TT0++hcb0t8pCDHdRyZO3EcBU9ZqyjRNDTWWX5sbo0iWD3O5oADn/VM0wx7gTu1DgUeICyei235E
xIgMZGI7KzIUrJPegLBFBfuZbN/8CwJ/rhxStehm55h36Qp3ortLlNwWi6bQ5ZFyoSE+2XGKHbmE
o7ehnt9rcUigxaPuX8HD1RDIeffsgh4vxqFKQ4oJlPzJClYS0fgzAREJTZe3RbWvq9w54jQbobN9
CfJgw4kjD/p5LnXaRM1j/FeAYpC1gFcr+vKdOnLZTrLtCymKqnPUZmP+ghq7/5ucvsnWzpA1Q0aN
OZx9CFL22ph/rLw9R5fHiHDu/it9gVUbCrdM52EeFAQ1sEXSWXGOoThY+slS3BxhmHsDPYZuMwpH
WHVQe11IdFehEJbASe7c0Ngok4iksakHMSqVlG12UghrbE+LB6T6LdJfwv2GlWqKmD6+jPPOEegr
rooW2DsWgQQjc6ysFdKRr5djfjb4oVZEmWGEJiZnTfTasnAWtqU12ZIbJsw0YHsjlTHh6R3qYDY4
Mfi+xmk43fLZNiOBi8agdcjR2mK+xnFino1r768uDn+hlEDUVY26y1wWr+CC6ItxDd5b/ZmVlYOJ
pTQnIAsuULWjFNFs0cCzNpRJd2Acq+cJ7aa/ChN57lhcOEgzQpnJNBqa58aiVhx8KhzZs7AYQPdf
ssS7cIzpYAUGJ69EsbpDu+8zJ1PNCm111i806JkLvRh8Bw/QMN9dgNzdO4XuJZUdFTbq4b4TIWQ0
8DzZQbhleTPFkJ/6Du1Fvxg8lrjGcgvgJjyvVICgB5BB1xpQOrT3PQc2uETJ26DkShmOEE5UY4WT
XRNty4P/VJH19q9yX2UFgtVK3TsqND9xb6Kc1Wtzs2Boix9R8w51UbUh1x0dULnZmOVCdvmnSspz
Mtwa3sLUvo6em7J+wkjpjc8U+HPfV8cvTYThHY6qcXj8f3IHEEnElff+m5uU5QhsAx8aE/sINic+
RerrYp9d/cLzUGdYatN5u19pgI7jWV/+xwGWpZe53d00nuOHQcEcosdf0hxgZ0iJ/OXu1B0pFSGB
4hRfnWCRO0TSGBVpBTWBqC+vsWOtS7nPSubFTCevc7aBaxVbXkoNR2Oe4DEw4UVRGacmshfqnIFr
qg1R9okV41GPlibHokC7GE913UaJe5V3PothYrvGQygOFwFs7gtWibSoMBMm0Ung73gOSz1W8Vrk
IL+crQ+rTb9+Feothox1aUR9XwaUmJ8eGGM/c+sAwnOJkhlXNesP94VKWe8BKbb5ljRea+Agpgyx
LEAW+st14i8e6zg1lMx7K1/SIzJ5lorPd4EpTEBhBbQjdaelwiM+ccLPyDEDkX5mXYPgjoTFXhFz
ieYMqxvafhFRfXP2cR1x6hiNAQH38iofvJjxIUph1wrQUV7sIrg/OKeh568kFXRX1WsibRx67tFQ
7HGVvzKlCCxC+IKiEZY05qCJOeCH+KOVQN9N3sXuU0Q80MxT+loQnnN/EYcJ2bd2i68Q74hga93D
IVmVc0E0Rfmv+WDDn5B3kl/IN6EMFzS23XMA8WUjEoT5GhNv2da/fFEwW3TsA93AhQSsWqInRwDH
vLfmC9U3rQK5bOHei9+Ako8neI3fbTbdmzO8/9jFFdqC+I/GQMdvvEFqZORUzguvOu2EVaG+/0PV
eX/pfXSbOYhDu/gFhpGsFn1SH6v4f7HggWquXr4iSS/adG8ZJQkKilK6yZx5hgu2AOQGLWbq/5wc
boWSFxr4r/xC2SX24sU0guNAe6h+SX2fWOaGrymANTfEyasOiQn977U8Ugxy3YvEsmFMfPyvIOJA
rNK/zqJqTSJboUEYieN/eAwyqMLK+HxYUgddaw4m4MYoHZ91ZPuDuCEN6cpQbgbpJkqvW22jK6p+
TN6zCzDv0wY73iWp3bVpYWSmDWomveZCQRDaqXQiq4lqI5iYU9Ba65IsloMV3HbNa2QkmPi7Uead
9c92voGrsVXgPHsEzS03kMISG1ntwZOT51Y07BpSt62MUUNq5PQ/7LBrEJmCpL5H1fo7/gN01rCP
wDUWW0zwqWD4Een9wy7X0xzH796EGvR22oz4MH4gUMHvBfvWY/Ngn5firho1G/8Hx79yxyvntWM/
OiOgV2l+wOJyg+07inlmv6jfUjwELaPhY+1hjRYfonYI17eQl89F/Bk3Wr470B2sbh1vHZ3XS6yi
PTVJj39HFmgl4STdkWEJsNgBqsLByooVdAnWJ2/C0w/Z78goBkilKlfL+JQTX3ZXIy6CL8KRrM3Q
faUhVF8ae8FytvmoSTML2y9UAuEdI5hH5/mOK7DLeD63GNtBtoBIA2mtrj9V5uq78snReWJVfdWS
jl6sNWvb21N8W1W258+P6WuE+zHrsXL3pday0pZSkTxAThXmNLbaErs3tcFFolPqvA6SIOnaGvzE
00ayFgOTu0zVjNAY/fUbwGSxMWUCMUBvJlBGA88rrWOk+FQE2+F0SMSONxjGV/n7+Vae5rc724ie
/IObceblEzWr4KB4G3hv/53aOKPfPNWYszaumoket5s1yCJg7IpSACp4JEsZgl/xL72hqQ1OZUMX
LxTjmiZceuMvGzcMbIHOdVL9Op5Vily+fcYivFNsQp5q7riVuLgC+Q1PMI1sF2N8ohxHY0WQ+dgw
CApCEdnmmdO4Q0OO5XcWilzJXkD4kiNRKub4nvfBKlkrK75abI5OP6Nr6MVfSXB2gynU3hOrfr8j
Cgzx4A40sNXb/GTK7wwVn6nVPDqouXmPdnjAY9pxtkleQC6fXlIr8I/FIoDlwto7qE/+0McXfk7c
T6L3sFhdSSWN9fWDQ7jKd1WHyhgbPo5nI2DJ13KFn+/N3SDuiz6bAtNYYe8QTYBJAW+roNinCf9J
NWT4TCS0JQ5W3SWioW6AL0TVBUbClHctMgrJ32WZz//Qzl34BGX2O+aTTJiwRXHawnJVC9oCZ5kM
wgtspPFPyjbETO0JyRfE4ilsGG7UOqZ7C6lVx/oUeSPpuHT7NWPG/HMZtE+9WHjQZVpDnQ1aHxYS
WpzZC2pKw2FOy55Jfx476XEasjVbtyEOeXbqs6aCMs/g4Y9xjsX9lL5LCk/TQyYqXEOk1wigB7EA
cufN+v6yYZWRhnz69b7PgD0clRxtYbKZOe2kCGbU7V2rRwXf/OacgpJS1hLNUcerBKfYB94zOp+e
mYYmhxfYbAbxlMeZwNq2p8vvbovlN1K+qeXjvkzsXWdtSQteOBRvio1bK/tZeJWa/YePCmUyWzYW
Mm0MntxspA97QE96k3pXH3/YLJJdrY7pS4Vv3z2Jknl4xP1PU50YxOJi7Rw/E7B5EkfBqMFxnyF5
soXOfLV8eyUhSWCaTsw+tV2U1Yh/aBq4RH1xnlwIj/4osiNd6OsyyoNuQ6wv0ldQrm0OMTB0iYaD
rTuMzJimT2SqB19bFI7TqDbdSmJyBB8TDE8RgQVu81yC1DDW77BFF0iqfbJhtJ8U+WKbc94rG1up
EK0CPsjq5efMM6HI27dtRQip7YhT2Q5bchpmGJ0KiZ1Y9dKliwT2jGsVaU0sihThUDab7zHuCtrH
NkbPj1JymEARo9qlBDc/3mCk9anq3DksHnFDPTmugRWHl7mwpxj4iLnFrZ9kWmuIdljD55452uP6
VqDMLYVBdvwrQ0uraL5OuKWOvRtuzFH/+BE7bzwFJQevXywus6KuLNuFNgqqAx6QbGYkqPi0zf99
elORanvza7VP0LM03jknwDKB63IqGpXcXnBcbU6yqmkRvyaoTlCkoG/nidclZJzlqNry7e3MvAKE
X6V8b4NjgaSMm50T5aIKuwQZhqyc+OIMzsdu8RHUSY8+xRyjzwjQRFhEql6qNoNSih7vbtwco5c2
oPsSzgEqeoJpstcE8lgnTHE5HXaA6/Y44ONfNdH2xxYzLOVH77lSA+DeoNOx25qBQmWOBRpoTnO3
sslHncYWBPBiCsAM92KvFH21u6LL14GL0ToMfp2yVOM9nao+jhMCWHKCmYNdo+aGZNAxQf7izNDP
VfnWpB7iDv19x76gbtTwgWu959qp2Ii6DLkmIVVLQlFqigQWImHw+X1o2+i667MXn1fCXAf699E6
mTmJnW7crUbxjDUfX7eFBXBcl5HLaZXgnWvxJE/Y4VWFRPbrBoElsAn2NgrPCmh2DqFP0ktMXooJ
QO6irknJv1qjqBZUeDbxTMTz+BFCyNaGBq5JyZ04M/bQ941PPL46qge46FvSfVPnP81dsP5qvyGb
iXn+/x0XPyW6/dqRCwxlE6VeJ8hsc44odDwFrE5+/LbetUgD193Qwm0tVYMynQ91o7E3Zo//oFl7
F42iPUjoxV4fJPa4Yo583nK6UmTAV+C7ZMDPKBg+V30W5uzoBB62inskVKkLCOSV1p/ATJ3Q9opV
xSjTAGNX0U3kOZUi1RzdT6IeITPvsRtYVPmcVHNC7cdwKF6YUEwzNh4HUbKlyedjoHW9c6yzb3Va
4Uc23aeksjeJt0HuPOMEruBmNFpwCyleHrFhB+bIHDqyZxZHLIX2II3EUUAi8E8j+IFaOyC/C0zi
w4sI7gR9Ud54DmAO+y9a+hGhdPNUnuKULPAJVjvuy3EIX8dsbVqVTryPkFY/L4jsX5vFVVSOuLUJ
Fci8Vnp9F6e4VIpHkevZMvuM3wrrb6HUKJ2bmFtQPSmOkVhBxZ449jN2tM3Q4/qNJH/osEv9JX5r
KaODxDd4vqeNWDim++CGcbqmWndEsGxe8v3iRzMF6BVGNVUhGfV8fwWRebjw/KTD5mp1xU2NAe92
GIfE45+DggM5tqkF5bV3mzCpnRjHiV1o/aRb8H9M4r4haKg0JbygELAaFw/V/spKbqIsiXlrdGax
bCai2w/rfl/K5lepbkqPU16N9jfmVbwXms4erEsnsDkca6eMyK9DLlMgyNmSVD6Lxe+Qh99TYhmt
sG6MTWa8Veq42/uVdE3vamcYLjRKVE2i9E2ofb6xIFYWWE15CDZRoccl54kZuYiAj/A5LiV35V40
oYjFlCnxYDDOqkHrtALW+KVrXZ55qo6oneDu30OeqxquAYMGf9oCL8fbQxKvvHqLsCmFvYKTGrBN
FFEdcJG3n0GW89MgiQbOSX4w9+J3spUg0YSRJmbQQi3sMQJsg4mBxVTxEUiflOreV2hMrMTmbShm
9loQXe+bwcsi09cPYfHs2+LE+N0M1iy2JZFKzp+57L5KmjKiAPccg/YaEfINZDKsrdzRw4FcDjMr
NJ25jKswf+TCjD9NefluyfdIyTBhrk/osk/y914xflq5fXwidne6McgFXyo0kH4FUUmLFXDfWplK
eL0KQ8MiOK9lHawPowXi7J5rc3cWjFqgqeyZ+RAxrfTPRcj65CtG9zULOwcx1wOKJIGz0MwpVUYh
HdehlBxnJJMRowrs+MnpfFIPxuSJOuhmvsGv3lLdyMjo+hUpzxfHv+1FLvEJgZ1lPiTlVLr8euOP
2QaKHC47QVYH6iF3V2W0l6y5kpkW5Qr5rp9WTvKAugsZdYfVjYaKvc9I/rJGTeqrMzotcP4oyZyO
+TR0m+jYiFuBOIsZeEPq/PQDwN5z7KugfZRKn0vj5QQ0gxsw3vy+BUgMvGZTg5NIulCgCl4YE3q3
t5HJlraEqxhm0zs4I85DNpE7VHpifpsC6wZ316eX48jThoIvc0zTN4zlMM3x0xEeI49n1dn+gmAz
Wcb3kWDXR28uMuKjpofYg9qh82iynsbFsbTOgdTxEc5hmVTdFp0drwW+MaQKnkT6YRTeORBL+hin
QKZrjtuT7sBdnMXjF90Hije0hgWFwrOXSTHPH9xef/OPFs9imch1OkEL2rklL/sLt/kvWF/oFSjW
LMdic/8+W9TIMX0IFaiCnu/7zsTbNVpDoYfAJN5+VyhxgNxqfUGSrW2Z9Ay7r96dnjzQ3r2hQBVh
leM5tnN4G2bPRNBr/jj+/O6sMKw/MMKvmOw3md65oLCXaBkGzFOwsY7zwzTcJhkMkj259Wk3TiNS
jSx8o9td5dd95APq24EJ9IC4nA84JrLaVh7zQLZSi7pgmwKgQxb+aZkhopyhwv5ugNSlc9KzOMoc
d15Qz6GjzXRGNleTxaCq19eTaR/kNkxJMCHM+dCSynz9YwK21ucmxuLA7K5eKBG6HcS8rHC8LRqY
Su+lXcbqC3sxYArSLHaLTZP3xif3wN5utqnTUVDMPu+QXpISzbU7oaSSBTRcdjouAe6WAUv/Z8TC
y0xj3F/xuVv3fHzD3ALeNeUAEsAL9tfuqdzwzK4xwnWgBADNuQzcjRROAjCzr9stHGuVraq4R4kt
C0WFekZSlXgI2SaPObJHX+IKTfQnbqTGk7iyDxgeGm3Ci2rhPgRRKbML0qyd5dlnfmDQBP8UowvU
ZotJ2M0snMaKQGWOOKzlie6hsNcUvEFASMNJRekMIzI+JhLODOXn6nAaj7wfgFg35MFKOVfFrgam
Dy8oIN41VpizqcgSx4jMXdcuWPMinSTtgGkIIuApY3agCnjXk4uT09YodPmYrA4FHWRwcOEvIVCf
H7NGIFmTDsOwv0BNjOKL28q623cZkEOGofoxq7ZI5UHxRuM88C8T3k8z8jSOQI/Z1nWSqRSurwvE
RxhJVjoA3nIRzbT9F1eJwLGFDu46AqeMQJ+QVMSQhSIpsdeOAz+dvoB3xcJ00TwfUCPRaJP1jbvp
w4518ppBpk8D7BLVS3Ifo8Xyot9ATprrjF+l9vW971RFUufHw6Moxm7IjtGN1L23Sg/TyEaeR0QN
KBDdburpnUTwLCE2E1VOWvJTnWG/r6AgQ+hXGdn9TxXkgvRZn+SgOjOw/ENMZIuzjwG65dK+HgQH
lANCfEvdiMfTvcNMAllN7BuAFEIeJ+1tE0fJgPELkNcy3tAMIZw3uiIFrvRriU3DWcrce2wWCOlb
1EWk5Yexl2U5SdxcqPCbh829vfvHMSsL9/T/eglZH6RkSUdECWel0wUuozgO2u3ot44D7raTnrbz
b6ta+YC6qBvkGBy/yUmrtNFoBRt2tB5t56fD4TngqFUwslOH8QGEbqAY8v9nCedAY833j3jzoQqu
BvNccOwSgL81DdVpDR9vwzWsXjs7gvJ4KYpo2kItDuQ6nti9XW1MOPAE++aRFC5bMZsn/1PePnUD
wHDCJyKTM6mipcXKfm4oCdBlLOBzZX0Y1pU3oNZUjcWqpOc0OsrqUyqFN2Jn7YKAtDPuPdC/Tlb2
IHWf9T3VasoB0hBgeU6K/fRYFEBQbOPVR5uEWN7WMvKR0TV6X3LhIucngglN8mefzkR2XMQMG9kX
lBRih465IppCB9tfFF8qvS1v/q842IKeAERL1XpfYtauz5IONqRapiKmFFI8hHG3aOf+n9n2cXsr
tfN4MeYkTxHXOTgPi10vAHfSo2Nu3tN0zOvwX3nUfgg7FTbIj61YJMQ7EuEDlfDixhpwsulP7sWr
X4O4XIb+jyxsIrDNYw6HFU3lEFxyz2Wdoi/Z7UMl8Ws67HefiQzY0QUS8crA6sFXSAxS8w2b7+Vb
92mkytxn7dRr/OM2B6POno+8E9y6uc2D8vbyqhks5y/yB4RyMggoJ7x5SfzZrksgTjRXR6PgFmeU
vkvDtifW59d1o8JMnhC4ULwQlP89j3GUlinhA4gISRkU9puV48x2VROgChqZE9UM/Dvrc+HJCa4U
JFE1AEwvDL3I6SK1pomJpilG2310k4jVSVBD4Qf71MVBbpXqTmS1bhCmn4k8cd/ohtuLBg2xj4AB
xuQJcpcEX7Sk58GtHCSWbHHohLEFhDkQstFUstBDjs8PW3adlSGeqhlnm/E2TB6HJR/axbupLTcj
EDXOgg1TXIaekx8ntW90SNHVwCHTWV48JS0ckfqqcJbs0XhrtixyNL6WcFgesRqdiAUBu88So9Fn
MEjX+BmVdF0VtGPzRvaCxf1L5imjYXI3GfFwV7FRTArVxX570x9RwyR9iP3fc5/dgG/EX+PGnckU
CH3nQT56NBicUu14AF4nj5CzaP8SRnfox9+e7/vplrQ/19X/LWpu+mz5i+7ZEKfn/WKi4oLbeM2j
LJPJ4jlRfSKzCrKXyI6xIXYq5g8leb3dC2UgoWGPERo4YldBUugpz3zzJBgCoX0Fx4MF5+kkE6Z0
BU/3mOEy1gBCoGGEoxH4938oSYlYHTPKIAteTjX/8Qu7R5A550eI+kijaRFwe/Vg6SfBGw/qa0uk
mQP4muJaPi67gXTsWW6HJ/hdYTGxIs04D9YqB+97ArML5VklM18iILi2Ci+34KLzU97+cOBIWhiK
D8+0IAXlv24WWj8yhiQe8ZcGJmva96Zlp3HCB4LK8F5XxCzCu+vYTmQfSLRiwB9O0K2v1QMWdAha
QYGRDaMqdGZE3UJZvr8+Bin5A4hyF56SFIuowq8lgv+6qVg2rKQjrAY30kK7QkS5MoeUwz4s0Qyx
cTq8k61yZ4PipL3iDlEwWhXSDvcD9YlPyBW+Wt/iBWrrvrXgk+IUgOhgDFjtTVxEVX/1S9moJox4
Llz6Vs8ZEn03cZJC/DGl657PjBWSplvR51t8eMBPxH7rnvbz/kGFtLM40s44Z3SedJS+QqccGWQr
KKVyR25JFe3ZOyhjWede0n1qheZdUSY7hbtyhmjQNOV3VWCwOnykKuV91jg9b9zk2R3UNko5uFsd
NhaITsZ4mHDYK2ID/b8V3MK2LSx9WiNWKxl2RmdOwpYVc05YNrVLC33ydnFkRy2kQGmyd2ckxU5v
zgi58p8URe2igyYMcpCDrGQObtynImQbQaChsdybc4uSgFt2C86g47Re4oRht1UpCMq9aQwd1kUl
17SXW2MRt965y9flfce/vF4ag2BC4m3pQkKEJs9sNkJo0MCACiqy7WkoBd8FueGFq14lp7CziTqE
tQGBIFwI+DwCluYZvxZIo6lfGKTN/MtvTMQHmFXSXQ2WC7RANNxOg6hm33DPyN2/iS8VdEEL0v+6
mK7ssc3u/uhq7WBNy/Gb2I4VjlQVnbWYT9um24lGY9cGLnahEEq0dSYSWlbzdFNBValOaJlZObfq
BJYeunZFIMh/vLyCWdub6ZTyJaTdWbkqr+xPJHMEB8jqzg/gRm6+yeOt791gmY0mT5jiHFUJoZSN
tQF+vc8af+BGFx7ULp2ld1ypdZg9x7CqfYkUIsJ/Ub6FX8ccUt9CmEjvEeyK1LJB4peaF4JOTo/m
yQ0jV/pa0YN3g1DjJsYj/0ne5YpXyiEsmMV//C7u5KP/lmX9bhvd0fsPrsW/9k/KjbTh25FDgHoe
xj/ygOff71VOw5Ctk+0SMRlLoxZSZ9016ixdTfpRQxYIR83yj8z9rrzxISWN+ozi/kJOwSehDZ0/
QJP6IZGcySB2uWqs9kjD9hmYMwXoRGQJS3z8nVTHwarPWKXBNax8EyNRnIfT332z6utgh/PJ+PuC
hTzRzARqgKHX90ePWwjydSi3YJX/+20kXGn/N3l8VU/WYxCE29qVm3l/2tIw4KHg4TaDleWib5rB
b/SNrXCZE39aonoKHCPOEUF4Ct/O9NrXJ2RtlFrXvcIBg74ZBigVvpmkRzwNVUCFqtSKA+y/TMjT
V3KzPJUSi/nU4gljQ0egXa97vtqo4kHWKnQp3EzuIPjaOXcfC8mwXveFVB6OnQdQYe5jZO+zDiOe
aALOJuqyfqiEeOU1Bsxj80LOO/TwAUCszVgEBAu+OXakWGcuVVgoz8rCb3cayOAl0R/zKxyeJfFZ
kdv+1ctdnRegDjVyJFUwYqGXu7B0GI7cExBTHsZ2fofvKFjTRj6y2TaYs1EYYxShxBtnFE8lbP2g
9w8c4Xgcv0HmF8TBq6hvyEVnipDX9hqktWCnOJxAbADzA2KEIVNmREV/ugPzWKdHGsUMhPwIUYQK
VQGCL01bvJMPQt/eT7UrTR4ANarSZI43Uo8jX0aLioFnKrOaAhR2kNptz6hCjBpiYMCq/SIkPdcI
Ab1LIcjE/V8Pl4yRlVmCxDkbh9mWmao2lPjxG8YS+0jtowFAGIxhFVyYEwXcdac0Uh7GrPNXbvkt
5GdKtGwwGuWH5SkNW0vWlbq2w2yZgCD/G592bPUwq9lljjT9Vs/R4fKqPKjmp6br3WjR2JQl+gP/
n++Q1kvoFOJAhuaLdJ9IjvWIP8mXjS5JfDXbfaeVffAZ5gjGjvXK/1GsYxHDAz96ZEk96pY+9C7r
mD5s/t4yVdciaiYzghh2HLp2DRwgMUGZkJxo8zxTiuQMLekV3wt06jR6zyA1HdtnRCv0kWiUZSaO
d07kqicMxhGVvj1JUlcOTIBKxSrZ/qNi0rwSP0EHIgUR3hkuJ3bqMNbKCjNZwk7XQx0QyDmWWqW/
+oFHEjILeqVbQCRdxZ2P+bwUj9Hb/vDqWIBuiLYmucctttifu+37KyDz7NQM6sXFZfBNxaGCFp6j
68IB75lOPDgvfVmRGk7vNmtmysyopbkYr3ZOtajr6L1Z15S1p7N1YnvOJ0/7ey/+pT5CubDQsPkG
uVwm863gLoJkGyuJSefKewaZQMAsvH1HTAAiLfYyrer8elhswHO6OSDHgT102qofydDGhjybyWsS
CTbGIazRIKV7Ye1AFyQuTH7nq94ABIsvWSPK2MgSPPT3w5lJ5D7ISW1g5ag3uY7Vov1+O1o1b0bx
5vccocjLwVJ9CuhFbQrjUEbGa/jkPDaHV4jS07PaoWFn2tPK6p6vCJSJjSHpWFn/7N/fIDVndVUe
EmtrbCsMw1a9q1TV1py24ayA3gijJPAteCKCiQ1whaE+MA93hQMtNmj8dmH/gI/x0ROqSb0DJhLh
ObiaDkZpAnhamYUMH4bRmb1afnV5TstiLW4PjqiwiJ10iUCAGYkHs00Q75PtOqosPkffGOidIURA
bCvqbG2aO0Y+bBb+xUCEBJbRvuk9CCsJeIeydATKVjlNUuILUaHgVfIAOkTpJ9spzTyzFG2VPKsH
lgy6fxt4PJd6AE0KHQ55OgyH5dKC1WAi/3zdxceiDHbXCx9tptp5ZDJKA/aZ0sxbF8Eg2ZJyfMA9
hbhUvg9RoSudtE++q3B75JUgPZgWQLLWi8nWmRmJJXW6IVIcWf21xytIzpezzhea4ZlGEVUHNPhV
KV25Cj0uTYRMqgA8etRV7r+eT0hmJGxtbgex02pt1R4bKCCeM+1BYiTSIu+KFktOEKUm5sqi6xSU
hO80vaZAe3ziykyigYb84Oszze1dyqRzw/svWxKsunBCEr0bRIXW6/ms273mnMjPumUGqa3sColZ
+QaRhJdNLjt+Y5bY2GKPiBS6rRCU0v32t82+Mi2m2NuY/a11fSMR4Ur2UWziW6y6LbR1BjxT8GkH
bAnyBDUH2FlRnPr3X1B1203tPkMbqwAtTWclq27TYf4zFJdfoJ1+3FsUtt+UzBbOPjm7ePIQhzxS
8rJZbMYGY/6o3mCLjJ2y5JJpNoyY0vN9N/sfY3VXRce/gWGQQ7qOT72a7RjWc3SobaNU7ypJSWdw
VXa+fTIyqskPw5o4pjBRk/z1ojZcF6cMg+2AtkLIRXPDyftfKDJ0oFzrKZiadk80KrXjjhvhikxo
++8vZIP7OPY3HBPUvpU5xr4zN0k2rq32mRE/QgVVT33NgF+8JJn+/Pgb4K4qM4q0v8dGDths301o
fk8OrmXGQ65VntCHlxe3IBlKmD64rfrzIrEWvNUCzdKnImTKkza9DLOo42ZKbBtcZoanYAbsoBtE
pcPJiXl8p1P9Ijqj/wnKWUeUt9QxJVAuDKVhqrsPbisrn6ShXXJF/jnFdEkIpFLeakWCsnBnUOxT
bs8N8PnhgXshMIK9ErUFYhr1JJelB5FstlCzEcDBYJ0u4Ryi9UuoE76UMa+rlZ2irWCLVRULFoXe
03/6ONyx2mIq20pUm8fv+0YSxLT093OynA5ZH/6a13TtgOSOgVqlrLCtkXs4TsF7DITeki1uQkfV
h+pmhHVStrUOmxZDK57cYFQ4jg90+woRaonNnWbAg8mAutHlPcBqpTJOW7lxQQmc9fa5c5GKId3P
/t/550+4rU8EWjpZwLD33MCWPjnr4h7eKL+JFEjE69ESv80B51bK+uk9Qj1t4IFEUFp7KWsIGIiY
JM3yYHkoPCd16cpgorVy4dbbhwjVc3f+KA9YkqUdfpmT+Ad+b89CxWve5+EPrWOdLtmJOLTsRB4Z
CpITK3nlOesYfdiMAcXcX3jjBKPPR9BJiZa9eyJV0PePBTEpHUYJRqTgSwWudQ5ZpuoPsLCbDg4l
w1F2M0yl76pnAZ/rtr73/UXfLLb9ifUXqXA8scGBa2gpYreZ01eIarEh53b/h9SbImFPJwprvzOK
35NllADpVEB9gYGmYB8qpY/w8nsGjVvlHfdPE+eo0Y/uByCyV4l+5JzwTJNsRWST0fn5pbr3c9jU
UYir7mivouSTvj0CS2suegukNLkoT80UX1JsCriQvVi/jI/eb62wuq3xsoE7Dna3rDF7g38286mz
ymsKyxKzzC0JXK9OENltqyG9GuTvZBaa+TQInTHz/9FBuZNK0vN52xIU0uy0xUDIXCKyRtOUUbeM
gqclMOzP4MU2X/Kv5puol3o0VCgbwhMgCWbEMIPNKtQtG9YJ+FU/e2Y0cHunrn1Mz3661fw2FCGI
gLAJQHLmGXVBm9cW46Yq1aU47pOdsyRZvwRlBKBpi48b/fbLM1prfDbJkkCjwZ5FG+UYbrue3Jp2
xORq34VoS8zrMqmbr6fVL6RjqCKTa5uxB0hreztPF+UE3eWoX+Yq7Z9YpiwQiAB64N9k25I+/ioX
uiddDUw1JoCknOxyqU5yv8zPjwnXaGKIPZSJkxqf3sTtJ4hW6JYv88/Jt57TCa/7Fw8e6jI3gmBd
MK0hdhDaPllcRSmNv3gvPRqlWyCLSEO0U1O1iqFTUjIl3zaKsTfLE9fZ2c+vJhurNX7HEAxE1KQZ
RapOrogLgbFbVWylltPxuW1NnGA/rZyBl1/hK/SkEkyNONdlafdUYFuejnCLjsurR1Ls7WCB9Q1E
Jf9EveMlsoR/jeVdXW2DnVLP2KkKfudsktdcm7etf0oRcVdvK1kybJnQ6WdLAykwiWMqEV1gdZjr
gNQG/wjBDdvfLSm9iBhRHtmkbotFtJpjHD99FgfKlMOrgUL35/o1QO4gMWV0Aky+IzjPpKEHcX1w
ARcq97u0oXlPNWFCa5FMm7qeAnR/zpMMLMU37Wd9JprQRjEiJNJXoxXuIjZY7rc+6nJpS2BGRBOx
sMsSGxXgRnEqsofFo540zJA2pVC93D7eqgUJJZq/DQxpO5BlYwNsZd6VgHW5/sBu0iLxKao+Lw93
Oq56d4fV/DKGv7qyfGqRk00zuPJA4JeKYGNB8Si5HgUU6tV+vU7RN0ETUcyXQ4HYwS7edltLAraQ
fkGjQ5DnnxDZPUMMsLwHoC9MVcdldGHcvOZcRrhLPZQUZN7ZVz69/ayXnE99sZzD6YFpfedyD93h
PqEwaZnxHQQCS5LvY2Dg87sYXL9BmAdlMLZ1LtUoirpkBHbeSugnv9UIy6QNb7rWVFJ2UtNPlPI9
ryX413mLMJYZwVqGBpdmHg1JS7tkfwSc4A7+XzuFgZ/9012xBK4madjUsye9oSYulvySu4K8RVnQ
R481S9WeQkz5gziYQsF4wLhA4+DXHIT28yqsIXaaq7My6VqiaCtLem33GdOfjecGARCW+UKIMs+J
k+/GNtFERwucCTCUs8fzisU4Ehdxa/RKvrvqX2DA3uh6IugyJhBvh66yAhCmadtSbKsjW4P22c+R
FML27qBRAyoFSogC0fbdQUnZYvZhgw/TB/p4yejjX6Aat7N7aF+tNj3EjVULybf7mtF/h1P6ja6n
fdtCHENl4yy0TxDEcT2ln/lsKZThKhBBpJfBkt4mkvLGAGHUWInlvrKMfj/esOwuxibagK4LE6ms
3plTZj92/cCpcPTfXKyxxdSN5/rZAhS1tDuvZczgQZr/W7qSbEHEuN7aNybbI4w67LVFv1PQrn1b
tnb0z9iXxkXr7FD34SFNb52uo80G11qIrhFXeQ/TB8zDa0ax2iBkHuq/HVbN1HCPZHIiGutxhvr+
0yhHVkobRsnfvcc75bBDUiAWK3l5EkvhtGDdBkUItev5BXGX3WMjlvOOohEtoPXczdP/UIT/RzVs
cFJw8GoUChEWGspMI1lufuTm4bZ1E5kiJ5CKcOUXhyL6mklYly0xWAXVQp7bal2WhWHMTpaoifB7
Q/KGvqrN94bwC7e4rl652mbPUayhWvfx1tYrbT++ZKHtTIqD20vZcIUAV1CrRsPREGwHzCXQFaGZ
Kz6vEYMTwn3YVkfp1AzJg7Mzb6ADwxQfj3qcD5NA8Wp6MH7DuOyTwZhHgiD07GOXZjKVLs2rfPnN
IdsMVkyrTkrOElca2vQGcVssYzJVSljL0sw4E9VpDLHrboEnk4hKPQj24TjQaK7+0TYOQ3iSu4RK
uSHRmKi2HuNPcFOV7VS1CXeixWHcZ3JQ8E7uyDzu6oUVeaApVE+KYO+HKtPjyWTnUzx1gTbAhVk4
td4RfoPTJtLQFCqb5nsQI823GY/zMI9k3RcuRucrbpuYOufbnembT3JxJxKh48B+vGeZXNnlIemo
A4OvPtai3pAPlRW1mdJTMf/jOT4sgIsWdMxaOfQpgZI5ONSqRAyRCc4UKG8O7Ei/UUBT3Vv4bHDW
7B8Qlu/5er7GvW6YWifzWGaqB+MAocGsK7wwGRpAD78KrfWZtkXmlmSftbrItDKYIryf8LE3+VzD
O75jTdiYb8gJ0XGpgc/8EZ3RBqrRhQ7lsTt3jwpAOJonE58tQl/6qinz4NyMXnwHStFi/oiBBHDT
gUnYlcS/Qd+w3ixNxxLQcFYCPljwCCrOL76v+pmbzuYD5CpLvLf1KsBuIelp8rIKzesAG8kruvy8
dowVS9aKLDy+0MRKoBiZJqNLN3M6xdjINCqgMv1LD+DP5rZAz/fH9MhoiPJCueaTESOM10WBOSi9
OzzGtYAOPQ+224lLXqQNyl5w3/PhpEowmmfpygbclR22xi3ORj2szzb0Hqv4wBopKzyPNTlAf7d2
oZqKvqQW3sx2rsEJNwf+lFo9lpuTXPNrnxSNEtpQsCMP8qSEyecmIgCCPjjjEpTB9N7L1ibQ/YXN
CgeLpCvOObLeWE6uQlTqmuGhMeiXtGwKDqMh4jel7aJ7OfaRcZg5utjlOxC5sDJ1MOoB/z1IVTkv
6G1glDqgcQDIv3ACsYb75oPU5ae5b0O1YqSeJdfb0RpMphxcdW/dn4nSw5BqbXpabWyqZ8lbFLrH
w0KVp35KXJ4jOktxIO79on5KAP9mWTywnCZFvwZVPhVwChqQjrfYx/cZT677FdNyFkZSQ4HTwtks
+P2RCwnfU7qkg8hqHGfsCd+SBrY5W1YG3Ox2AthZK/qPDiHVZpgYkLJ/Z/p4pzrHQBURoH9JsrH5
mM+JNgwTgTGm4FqGpC/dpkgii1/xr9008RFTrSUQBy4xmqL/XFuD1pjdlrCz/wYMsGTBIWHa50ed
mC+eWJmydo37LxwvKcUzPD7nZjuL2RSEcspDgQDFB1H1i/OZMDouyrKWoUSYCgtt9vayPBxhn6mB
n6H/4inbREMFktCpY5aMfDBnJrz1Wi8Tl/fRqX5wH/kiDKbcj9FgredFQCP2rMDjIOrBB11Nkxts
hgw9ECizPFW+rGNVcX8euBo4KXduoaVu/7hSVxLfmM4cDoKjtNg7ds9J2OSFeOi3nVETmb5E5/Rp
/xUyRiiJCHNuDXUmqsbzuubCnODUpgeQ5h+2JbUsARbhekllIZw7zbs+nQkY5Vp7yulF0/Y9CiFG
07gvoLED9wt4D+xIuyk3R5IcD6IpexmpfVxbV4hYo9ceFrjjHQR90JulLS86lcA3NaaUwxU2OyRt
vTAl8nbtBqwygZtItPzZpkCN3MKXtQMZABdHRgYVprUPN3NedkfZ5Mwe39gEex8niiwxDu7rmAWO
vEQJkx7Gq2axj7RZMFrn/UZAokldnBWFWQ6r+NSxQ+uRLNyaIWWBl8AVOngNK3J5zmKLKYbwDPs0
05lUSY/T97NuN+oOnWPb35TZD2eQfkgqT+EfTX5LxzFfTfG+peh7FjLwcIvcyvRDD7k8qZEeKT4E
61gtIiAmU7B7k+uaUUh+cxAPvp4KVOlw9f9BRJPjCVZYcjMyzbC4iUQQY2F9oPGy3E/yIqVOwYgT
K/RrraJEMhtdMhiJa7Z/hEp8OhFD4nnOCOOyWyba/HYKS0hhhqJJQb3gaty4LTKdVNqYl0qm04/Z
HwtFzj7/lwzSMOTo5LhsyBuy5QJHYABr207B3ONI0qb2GVXXG2HRZYN8wAgYeicKH78CorRgd2ec
75XJJ+RhCuYKtFSP5RcyzQbHNQyBHEMLiaHrwTI+3qOrxKoznjT61uuRAREICTSL+s6C2bnAeKdI
5ZRLmu28ShTys576mWwkm0u+7LrFyJ9cWzoDYBXLEZgQ2uGoP/gEPJ1TLeVIki1WhQMiNCMXnNLk
Ii8DgoawveSi9dCES2x+U7EabTDR+lEj8xcvFXpsY43zkMd35dVre/vxXjktcf5CniFpzvSyPMd4
0z/AgCK5whTu68uq8jOPy539tuwxcPzsdE6DE1zWNVoyX4/8K11i3r6DVmtDOZTNfIz0ogWjeLHk
DzRIZFb/sarwkRTlQsxHdPGUn2/d9/Mgcr8xK+V4k0cy+GJCJLHyqBnuzCDx9zmyBUXx6cJXEBXd
p8ABWi8BSblaKsNzfpI8+c95G7fovDfTEF4TGOgSsZ8XDuprrPMobCqn+ebV8D5OF7Tzw8h8D29A
KQpPGsjuiK0tdjNTqbewklxfhB1IAkMhXNA02CEWaKDZw4rjCH1piEej703LK6eRV56/7SGGRfy7
yCtdwP+KDOsCMevqjqN31rSwLtsjYkiSrX2hz47EuroGKRqmF3um1C75YcI+yfDFDu3j3CHMhtAA
3tgTDwazch74dVYpXq+hFGDEmrVTY4qF7BVKdOFR6jvjQzZoempwEIoONh1xotwuKleb5rkN2PfU
vwf1hG8NOYkIzQA9IsSHNgiU0Q0KuRbOQyeX0GsVZvbHIvE3IsVoIdcuc79QpQsi87/7iqMnGj7Z
TGLdhIVh80n/Yi10lGZtKlZZcxteYexgKYAx+XwI/lQ4GFXNddrNdhC2Pr7852FYxN9DhICcJtY1
w2idzgcz5apC/ZBrnCG8QRaElq7BkUh20gw6cf1xfoJCyZN6USOUVWqdZznuJ4H+HFhjpVB6BHiS
/d9SxS16cw18A9RbV/XBEx5g3otEc/m0myVw3Aq3nkytLSnNq54CrzR5B5L61GZekzoWnB0gtNTA
NP47dSnVJjzwDvfwNDhv1qnNs9ydQmHNUkDTBptJ5tZfCEaWjnc4IG8ZpjjNT4yIZ+CyEGKsXr0/
ZaUM56l15l6FkLVy4zHkwwKEUSW+MS+DCSNnIhEKPCXXtVb4NV6oVmTU9CSRPE+7GUcipNvezbx4
WovzYpgsq5JFRrEUQDAnuLTqWAXaAuQulVplebOrrzniDH9Q9EsrFvGEQeP9/Uw1d6WbZdpkoM/W
KL4Ydr4JPZydNQL0I4I4+n34iRNBDhnmu+rsVLj3XpDfooEre+NkBnZjuU/dm90jGw9g5KUSBEwT
SX7C7NF3XWZ4GxWCu22leDpSai1/95UE/hjsUwuQUK4YjXSp4J8dcIF0qPdeZKZ8TgYjj0s/7kZ8
aMvraJa1d+U3O0Kpccfe/WD0Zo6GEZEUIEUbmGLF1TVORMfPoIZtif+ZyA34vv9UEBDSf36Rr5nf
AZbrN3yIUsvOGVoiKvmfvBgvoe6Mzrgz3i7XtL2Uq7N4YENCifkdFbItOqUieUAV0wCBmxGDhGne
gTMIxmJqR/IhJccnl4e+0zPK4DdJnTVNQZJfhKYlzRJHRzein6I5GFIdPHPxBFDvdDhMW8mvbTkf
tpQsip7pRQNSLL0nOqe8JdBE5xJ+XWrHJUPw9YhOSffFx4qGlm5l8xGGWJkPSfW1sUd3mkGCf5oU
yxjTJK+S6rpkfquRJ53U9R0yOUchw8oXK4Uya3oziLh/FIdUQ1SfHvgVP4vnCmIXpH+1mmRpR4p9
lZtIsQomCFPtFXNxYlddv9Yd7zomuH6wWFFPrGW4cZkYUB3YDwBEPsW3SkYCIPOP+prPREL9FebU
974f2BuJH1NFj5KYQ5/kSCLjpqpmvttyf9ts2YOKm1WD7ISqGnTrYqpijZXosWzYUBm/NNfjd/PM
Xx4aUw6Y3OG/Lo/pAmUSHyjB5OdpXAVZ8uPxDH2E/AcWoRBhus52CgDg4UgOKyVBnZnoGzkauvmv
+69VORsBcESi3CK5JlbKwjwPGTt3BXr9maxV0VkW+vZnd0awpo8ZFxow/KV1rGMmHeNJ2WIS8enJ
wJuJ/068bSUswQCcANVfkHJgzpH1Llt2y6efzjIvMxhSMNc7skttZaoMoP9nYzgbbxTJWfxVkr61
82RonUhRrY0Bu3N4GfQ/G/0hATHLIahK2qW7B7A4v4i2r43uHJ7dbKNzCuXXzDoQxoll3RtmYgHt
kc6OId+kBolcM8NeHM4kdjKxfafJx22hdpZ0Hs5PsPuv8sa6nYVfwSvXcsbJHHC9Z7bEMzLxce8V
KVGXni2hqSqfCV8ulMeXV4LAgUpJkYjLiLnLJQglh1ZBZ9olznaNMo6Sb0YNj7gwmbOwT7Wvsv/s
6CW+Z/qoN7Cog5RplzL+BraEHX5WEDsNZfoZDJuHAK/qfc/ckpAeNWm9WGLA2XqJrNZhTr1yGIqR
+0rfO/LhlvtqZYNTJxHsXg1ZoHM73QfTliSKYU7I8L5vxAXMpC7dLlC39KCCtDxKSIYn+W4p43PH
Noxq2TllojcewkpjnBruCvFf8yvQleTCKofpyFQH0Rc2BULJLDVfOK6QyEeqZRCXfyYTpmqCAfi4
w5fKtWmSYTuUMiikosFWJ92E9MhlVfM9NaF4kceZuT3OSZJe1aXJnWmaCU/GsOnR5gjDrDZA26Xf
pwRDPwMowP8OHsRLx1kJQuTSPU8krgpueFnjxJntu5g+Rs7+x+C+ctK5mm74MJbIWLgJ1NR6oFbC
mQJ3EefqTKarrYiJIMIsBMM3wKoBXfhP5Hy8kQuFqJMQC2pKo/YVYEqI8rYKyg9f9IiTbJNaa7hc
o8TFz7ktxDdOFbOdKwWs1ezyZ50QS2FkAsd6OLelGEjFXAmVcQq/YSZMogK5nxrgp6lPmLYBi3T7
v2ae6StvCXY+882Cm14hTACBbcGKfi3fhh5C33EZhjSR7u/U07Jym/kVW4np5w9prtv+n/UC1ELx
3Xw61KeHoBT+nVQZGi7tAJQo5TWdF7t/Pvgev09kcKZCWVZkzOSQKZdU1VSn8MACVvSHs0kpGnhe
lJKMmd1/fVLZ4bXly0AJwTHpL4NsHZVceJ2HQv8Xzndc/92IrMKIA1JCKUGxD/5X+3OsPQNSVxTC
bYH0KAijP5SrXQtk/7YKdLVZMqUSEEUrSoHeBphg9cgEqQyhvephdew6fp7ZebW19RvGOzFV0We2
h2aK2F5v5IfbtmZXE7lmIBapI37ikf87rx56qf3029fVzxuuNU30Ltu9JmjTDEEAx5jLMSBj4lxg
QQvmfWG0WS1swZmKcPYW7RVRoPPUPb6kH7V4giRQVi/azae39k9Q2P1kGiy0upJK2IR+mn/YNljb
syb98tcfMlVz2a2wIn52hMzJOGvl/PGLrWZqlRQkVY3NxHmEJDQzfYy9YlFeKT/17jNc6xN4W3Tm
1DLxjkaKbrs4AgoOFLON6NKA7ZJC/sHlHIbT0AReykHCCInDBcy7MDjvReNPfFB41X10L98Xvxa2
z+Gmwqy03VBbN8OQKe3YeuByqTITt2n7c3gRShmIMiwWhe53Ho2rv96LLBJoOGtoEU41xb15Jf+D
dKFukitO/7Fy7waXQWpaTztOVL7qAMxDXH2IinxKs++yR8RbXzekKqS6+dOh68JUTRFdulQbSr6F
DMrWXnd8biE2Oq2q7CxqSaobUvyz9/UHBvbcwZlJ7gjNaOP2hmrbeIGy43+JoaXQnRSGt2vvQ481
IiX+eLPbQw8dknvrAGe+0CA307elgbHzV4R5UCOB9KSyojHvdYi+L/fN66uk7w0Z9zfjtQcc9wAP
qO44RPHlVLFMISPV6IGAQvBwfdjAjXOc49VkDGbyaBeAf189wcLfoVbwbvc1lyG3HNmiokCxg+pQ
n3fc0DCQtR9NLrSwi82G4V71a+dOZrOp7cJBzT3fb2kYx7um3XKkqhKa+Lds10tE08FRa3o7J7sd
sdWSwBQzxtV5FAum7B1GLuuDkoaVTApKDQTQJqoW/WAFADEwZ2mFtWKdtHVHcqBci2gpOGnZSIw4
mp4EjlIG2wvkdxWr1wQ8Tg/2Zt7DeWT0ZR3njcItmkHMXvYa/ODnclosL2KTDrq3sO/Cgon9bApr
wc3nE9hs05LBJ0uD+J9OKzR/CBpKbNBBlqe4dvPejVei0e1PHqpwuOKHl7xAGHz/kH3Yz3hc8Vep
L4aLpVEOzifhYHsH9SrG0PFROBDgGgveD0S/rTURB05J6TYoHAUgAiVyVqLY1oRIbhXXOo4OyyDa
S88eNRFxZDU1LmkiGC8YyZu8njWO0mXjIhBYGF8IdoJ4KPBdXuhT3srBfD9H8qifap1capuzDZJ1
ta+wouRdVVRSsbylCs/GjbmvFHpcjq5pHz8cQw9kna8WB6+GRqGFzzp+8OKLzo1ExjgoCOoKSJL9
nKFdOv6tqd+6e1hmFh/vMAhWWmKDpSbdSSr9Cqd0ZINbKxPCYJEM4o9w82uOly5zS/zuNM0bpSrS
3g8YzOnSOYGlNpWmViuHTxloB4KDNKm61qTo/fPNtMDr0ar5erW10qrzwZVnj7LiTQb85QEycasI
/40eTOlyaMVBbFn4CRGV0wBTx9L14TDzZob1dMBhF1GePCAFbmrMvpLmxkIcGs3lUc9s2drrylgC
VLkiLV1pn53S0Oe4ieJAwXED1hMQr9Qqg5IH5b+4/U3wrt2p3g0OZXC/n3UFsr53haql2XRaZX5u
bRWcuLdCT8KTgZYQvM9Ibatq7oovadCWv11JbOUgnwuGEoZci+3L0pyXtRhYG8iZ4kpdRsyt+U2p
3yWWtdhSJI+SWqEUHnvOYlx39U+kPaZxquSiaBWqr5nGDwYm9Uc9s45aQpl2ruRuMH2PQFLZosIL
AYS4tl/A6ex0NuSZi7qmFfAoNo/PIJ1LjVug+xQ0Xeq9+g1N2wGvYJ3qUsl+fN8wAHkD96vya7GT
USHAz4T0HXD7LyUBMuQSib0Fw2wVf/ppiX7jwzC3ZXtyPUMI/Cf6EmiZ9/0tv4m7Tshe9mI1Q27C
7kdMobh8+unJ1Opjifg/SRSvX259n3p4Vg31ko4lLVid71KbB01I5hNlnTownxpyZe9ygiuQenL9
3Cpr55n+GoLcuOJl14rUOs++ghP3Lp4N9IGvASLtNEfA45CHQ9McQJybisbxYJdyemAdw6kR7T8m
uwjCy3YDmYueKmf78DPln2z7nGKmWQmyq3ZkneD2y2P6ACyAGHkqcnvTboFojWns06MDIi3Jt5tJ
S21Vyk4/Q/f+itrBWVkEtFIe5wW+2jJ2Q61e3t070lu6DzWo6dUed+2j3OtxPEdeW8F4HehQ4MuU
M02LU4vpfalmJjDT2Uwz7b0sRKc+p6z4EshNv8OxK7OXIisEFMVLnno4HgsHIGZcJhZzX/4OTke4
/eZ6ibXZnjpLsUhTMrByXxVubXWFFFSfd9V+PZmQbabgDLKPBxe9cU9Cl7cuNT9DjNajFa+lJ/mc
2KPhJ+sWl+STdEB0UvPhm6t8V+RXDDwJ3z51H9f2jkuVnwXo5F6cLyJqvds32Wk1DrB2iHTLuBSV
iuPt/CRmaS1+iynaWoVOcCQnFOGCeUj5Xtnp8gkMSil2ujv5lr9NRgaueTtWLh1coRUwudEy816d
QBQIatU20wOlRf4ruN+rTYmpFuB8CCyoaudNT4vwYPvv86JguznbIHBZ15+ThXEDBHys+Se+pzvq
icTwxLUBRht4Vs6YwKtvu5G4oOCaUMuAeBlnENnyhOBKY6X4Ui0+NoQVY6IGRXRGEeVtuaUVd5a1
saoLtmt7ODkkybppozYlutiyDiKktcW95QgLDvTz5nkSvlK+QdQmOYgAqmDYVbojfkyqJh13ngBl
HufiwqOa37As9jxUrwmXHMImRaWR73ZE/OtG0qab3Y0XqVMlrdeqpGGobH6vYw26R1j2yB1PzLqv
veulsm3KfNcwZ+KeN8GZQFdRkJ/8KbqAiMPhRHFxaI2TRLg1SScA0kgmzmCtge1RRoVTt9GXXypY
SYTHfk8d//gylRV9DuE+hURGALP1h0HSNAucuUrJR/WBFYCDkUib6UJtPMyG85AI+5uJrCuBLIm3
QPkSj0/GRTszeaatINUUJThLS09uw7Ujrp1bZ6kSk35l6hlKZfAZgJtTgo6mPArL+LsN4yu+9un9
fYeFepDBhsQN/E4iLsoSO5b07N9v6BqGemVlebIItglZ6qfKG6S85lyevi8YcNGtEo/YSteNfwLy
YtDoSp+pipkeVHhZrZ05eY5+H3W1CX2CSK22nEO5t1dY88NMoNXeB2RZLoWAYCTEfCCbFN/EDIse
H6R5GUqRYEf4pB/0RthXr5NEHb/Avbw8965f+a1TzNe3a14snqf5LhpqYnAx9q8ytgIjASjY0brI
v8Zz4EK3iI34q1bBvZ3j0VOJc4SspgP2Ud/oV1k89PE2mdJeNX9bWC1tAz+bYtzE1gcsX8u1WalE
wD+GtybtoxTUdGrhufcNyo9it0MOlCOJttP21sO8UA/l+T8p19+qWDi5lbQgSxWfF833lvCVRq06
mRyNLn3A5Cpp+Gom5zdZ4VbT1Dav3Ym1OEmtIAMdb6klI2BRMmxWg0XfXqlfQDi9E0khf7RN2w+5
x3zKyZxbIp8RivIilEhnnpaI/AHvUPNulBrNLG1xL4ktLhEO9/fA4WwUiaatcgBM24MaPgLRZGNC
HVKuSnjzfgNoj71iFBH/FYkbzOHIVuUOeHyhEAvxe3nmFzYjs2nRWorWzaY6yYIvA9hjvYrPlIO6
LEIymOtN66VTvmAE6FvMpK+uEM7uzT8HTKATwIntTrftOXwQPJlznJVxZpdSXjxjznRUWkIMbp0l
UkGuDjHcX312derIcgRS8dePR5awxhbEh/7wZP3S3I2wkfGBfLlLcOW3yo1nGI2qtnVXoIhsOdQj
5U/bWIbJig1gmjETuKkK7nHkGSYp0sW6vcHD8MDGMHglCm2PoKt/IM98p5VDnPLtXjUnl2HKYsYw
j21x/QeOjiI1KEk6zRzK38dimBypqUyItabR/sRHuhayqHKPWCAmdXKkwDbyV6ATaKtdDctSxQlp
JDJKvlrHGBVoxXo9KsIpL/TQhPFi5wfCrzFmMbxf+FD7fxPi6Xj/bME8JhRIIRiB04WpyCKW7vyJ
SuceamaD4ml14k4yD48pnsTPS9RemHFLmSr992PxcYNHtZ+JvXP+wNVpuV/lFvHzThr+Hhh7MxEx
g4NfXG8Suu1f9OAKnNGIhVrd08+X8sbhJjPzpOWE+yJ1QN4ZLpqhQkPP0g3CVJ+XPDmGMYhBiZjB
4m/2Jc42JyLxF4Shqb6tyaUO5ktihUpetz13PzyD0zpKrI7l8g6xYlSX/vu5hvT2X0QFpmbupxyq
AC6ZZLCohnR8NIW9uEE4fDW88yZie1OIN3CQfo5hIJ0FTxl8VrO2b6pWoTfPyqTaWYW+iDgzKwkU
d4lJjooEMwThU4ScNwaMt7m+0L+e6uOQ2ie8JiBfb+GNwOi/DHTuL8AaZ3qRHIiP6IVeqr4ot/qg
KdpsgC3M/O2yphcrUnQWpjkWjld5G6ObYpGdk2A6rure3kucyfG0HuFwKMpJ6exRvDSgmnNo/+9k
7mmkTVyqRKWf8nRiqR5loZG7knXyqVqJKZC9lHlP+MDQiUKNqa/ZFrjiYwFoXtTuk5L5EqFFm0tj
0JHngjHtUei6f1SoSRMLl7Hsew7pPzXAWpvRu/NltuHkVT/6eA37251ENCEH+UG9kAi61ZvNhfbb
t0mZ+xkKzoe1oDAwAvIJnP31JojL1eZe4F3bOFHmCJrjVIIu9gynO7/7tgpr9cWQ4xBQ6p1WlDHP
ufUGb0DdTkyPub3xb+VZVFeRJ2kPeEim4msa3GdJRYL+u3rxpouLeqzXLHGdQ45gri733/4rBAMz
FqgpZdPSeVSTj0dyuf0Cjcbs1pujNmbq+xUYMQI7uJJf0d+4V93zXDF6sRNU7XX3r+/tLQNYvg5H
sN7BnCq91fSVBzFn2X+0TP04TTjFY9EOsQwJZcVwh1p8OBSi1hmtT9gCqHowmoJYu57hnW+SSp65
c/Li7OFeuTCL7+1nbZCu0ScwqKvuy/koBGWbiKgudotPHW1hMt/f9VdlQJfM/UYR98lKSC2PLeaK
06M5MdjGVulw3PZ3HXVeBluPDFlwHLDevDncHMSSCz/n1gG0Da550NJI14XlGue9uG5DtRJd31Rb
2tdDFRI387OZ8GjpDN4V//Zj5ySFRiro4D56ID0CSywVSy4UmT+9QMSNzUzWuJgV+Vl6yiqeRBfR
CFaIgJkWuPlgUgqZyqPe5zHkVOQkpu8u87V0tSy10+hAcNKirIAh66Ce47TgTiEpcajsb9mcFtaV
pRKWsJOClbx0v5neEumb0BGMpRQuiwsJS21SsLBYXbnTITdJgBIrMC/ZRDx7ACnyhymc8uoCbjem
IYuiczPMkUjnVU5B7UQlBOg3ZXunpV4m3V2/0za7fUZ/dPjmL8LOcaNeQ+2wjrJpcYEuwWFJfDyF
x15HTDMUdW++MK7vHp42CiZFKUYFUBdssN9Ngg5RfJpYxmzrCQPV0hcfEmbfbKRGBwHyE2Hd2fAW
IUpRi0x/jeADLagZCpHeiGNLaG94BLjVxkfksDoWXtWcAoDiSeC8+Yv7eu6bGi0p7knNanahxgXZ
DG+jizd/eU/I8aESrv85sBn7Ld+hcv/p8DXFfigDgbR0h30NsIvhj/T3gmfuzLHzJKN3NJBBnOEp
D8TqhfTfhf2O7Y0KfOH2Kus4uBb4I7RhP/Got50KaVbbM+DCrc8eAcvihtIr1XvuYnvxVYHaXRY2
7IvorX7t/529qxn16BEZid5D2JIGe0ECAfCDu8T2ncaTPW3//XDx3hZo7NVXGHaoTbvyowi7uaaN
dhn0HCyIOZoX1rJgD/z2Eq5Va46xlYJjkTEwmQMPHWUuHGPLlID5fUp95vwMOR/oFcdWb3rPSD2h
Mg5wsSrALrJa1FDO7jOj3LXymV6LoH0RsEN2PP366VAEpA39VuT7nPupRnw2uF0ysz+0hZSG4YHZ
FWjg/dwkmXbhZvbGEBPnkmbuB0n6vse8oULv7syNt+YcT1ZYLC9tGvSFHD4B3Atr6wB/ycrb4d1N
rroOxehPLQ8tc1jJOqNGqTHr0qe7olKJeTiDFVVcsAtwYBt4+eZkVw+w88HOfw9/IRpJaoee/jvg
r+LM9+B5xPSGGrIuw3M9ZjsUZflERCFcgnKPzYXJW3bMFRQh5TMQ9gjyEs5TV3l7ngmgfOfICkr1
uUf/49Lv62CR6azswAt/510mHif1k2sKnqG2i/dICFkbEp0S/Y1Rt4hpqtGOCp7L0yuSjRBnr72y
DrTkndZs+Hblxd6eWMpMx/O8JL3cwLqFujXlzLZfDZ1rE8vHgw/YM8KNwX/w/E8e16XjcgYU9Gi9
DlUlV2D2+7y8rU7GBQP2x09ibimlLN+qvQNfUF1/PKlhzvQjZAWrMq71ZE+8jOxbhv07b2i7GnR2
UP/d4piQsqk/jUlj4Bril/IIT/v43C8GRjior6PKqa74iuAkfAmciAc8PRbibeC8ZtP8VyfpwyAd
0uRKlF8npENOxMZ62muWcrdemqP2WrzIg7u3v5np6IWA/8aw2JJCIh+fjVQE8u4rn8N4OFSMbYlx
XNSc33734KCz9RD+U0Fkvaqe3ersOjHhcfvVZ+xQHX6oYgrBpaBMPAfRUw1YqyUJN6fcyVzZ96v5
brb7ZVJoJE/gmDXauqdsBX5iKOolV4nrXAzkKPBNyOsy5IYaGsNuU8WUTNv47Tflq/cDPT/qiG+5
fB++0Ntl+FW5vn6WVQXj/EOocO3+46nJyfBeQkRaKNcEpltUFlEU5/Z8mOUtLTrjOYOls517SNlZ
p1mTPixwLwfPeXO7hinRTUkrp77GPUk4nl64/8MPCtqDHAUfWGQStpSHur0OkpdwRx1zpetZ/8dk
iJuT4Zgjn2DfD4h/gQFmTsVsN/k9F/T7rGAB+vrlEGVnlyUzaaWyGM+WQ4YaHuFfIwc+TEMD9VHb
trtrWP9wJOLhacPNqcw6CV9E5E0tPrsYnUZbzOXlgnu8l/4HaVKIOwbKLXd7AXukmRqilPmUanTN
Q/Jz1MTTzY49mNQUQBO1oyeOyarA6goDb8eEw4OBqP8VHyAVmQhlhcQx/EDxU8RpM2xnEO2AxmWP
NogmoW6c/RYWElrQ8V/6RNrthqKcrX2AmBfMkzTG9dAcm56bTbb02xvKLZZ7sAYtOgnSMHT0bnZF
xdQYgZUhcKox6irFJIdTZiakPnJgXKM8cahbmnpHJ4RZn4Y4CFO7atN/d1+qZIzfM7FKeztz/snE
3P/kx4TKe1Ze9NAaI1nW3R75E9g7Jvmf6pVwlAqR42h6Jqb01YFII2GGTIFv3WaZD2LgGFOWP1+5
CYzrY7VgMlm+312jxp8ccNdXEdDXYJACMhYI1PEV3+M597SnMsPvaT9q3q6/iUrOnBLzJqgAcbrM
PKGZT1Uz+uizK4TrDdzs4ofCERQA3y2whmiyoWfX15lJVM9ddh6AGjmksfsIeP+1fpDr5xu0UlYR
bCoz0uSkfV7HnE7IDAlrCj3174wXZ8A8VtsGhNM/7BZLHztH0hWcoYnPlRA984tvaQc1SIZuiUi6
7DzleX0fDMTPO6dfVoolfg6pkmGoGeL4qSkpOIvffReczxCKR10xU+DcRmHZcr8hAcIzjSGhDtZn
2Kkp1VjfTRPTLYcbbTR04KPCQ4Trq82HSNRDy6yx7mBtgy+vpyMBYfX3IJ51OSqlzkPtQwpori8l
jsx0ylwN7yY/OImGFGBnScAAWegAfk7arwluLp4wvzShztcDGCRWi59rMaAf4FHIR83NWvVq1XUJ
cNWaKx13X4cfu7ps37GRsk0Xl/mEsdpBBteoS7iX06ql6POSvef8hM2zPig+Eust70I+kaXO8Stu
xvp9g9oOMRo7iImsmWRFEpK2psc3KToPcY9gkrquqBivUYqgaKikM5dpD5lyRCB+E/SILT8hM7We
2E8b3ZBuGr8ivRwpT7rz25QMegsCQAhm4VVfDUPJXZll0HHD4lThFAmbTGDQShkArUfQBG6rPcfs
iLVzb4Dqthw+9ok5vqmuqj1arPztvFHMtfeF/k/J96w3sSfCzeoCxOnZW709+MmcIeV/FB15Xp+p
p0PA9pq1phYquCGXMzl+AI8k3cyvvKqisz65bz9fDE7/wyMt+3vrpiDfjyrmvHTm96VTticiKX6b
oZ5uU/08Eu7/j4f63peL6Dg1ZOBjRV9uaOe5+btr3aZmHuG4itSSCJal6CV59fnumsIdpztdeI78
MYXtxMjLLRWRS4iE5We7Xri/dRBfU60ekOPPdAhN8gB903KwX8jqkrV/fNYhjENkmU3i4lOHG6KZ
K3KUar92qwLq3o3+3KkF5h+c1fLjSEiQ137Sm+PRxa4PCKOre1eHthxMjTCZSHxYE0Q1ZZQkn/4v
u0pNc9pdnXriCwGU01Ytjk7XNKmQgYPy65ZW+em3pmsoygRiENepMcKQBwkUExkA/ACwcwGEJTCc
lLwAWvZtpmAdJUFFilkRufWdpMx49UIA1DYAUWA6XmQzGL2qcwpMtYcQYMgZEbblgZttIhy5cjnE
t0t3zoPdczJmPSlG8th9nhIu1eixe82h0c7kn2bInwmQIVTw4H0QNxf6vHyRovVY4FbqU90yM3km
Vdo4QMX+6TxQZ2JEkG+jCR2UVSbHnWXmXvwBr3I5NRGoIBG7HIyIPRcJ8PH5Wjf7ZqRIz9vkTQNE
y/mbnojji4l+SHJzABEMteE6eGFXsnWSA3LK/VDt6pUTU4MRMOfEyg5sWx7zap/3kv83NBW6mNrt
f55yQXMEPWhqRHK1zLqH6zecKzmCdltrqw2gR0AfdX18+2qyhGXTDIhqOPzA+z1FhJmrLE4OsvJq
NlFc/oyL0M07i0ZsUgtBe5P8H20H+FtzWrY4VWuz5DtYyRt5d1gYafMEifi7eFHsXBUyQFj46LOA
1qgGEzMM8yQXvTwLI/EILgWhBl2crrlGFB09PwbNaQuFDIPzbkX8pjjLhXO65U88Ybff8VdLc+cH
0XYXRMTh4HCzIFDJVRruMdFmHJ9T7Jg7zAgQnTDMgmAMVSv0oAEI/Uj/Mqb9PYvHjAm3IJpg4vIp
hgaQxKrkaORUv3MUHmvsL2Ir6NiCeWcAOK2VaD4zQT9N3GYT2L5PQphQezuUqSB607mGB1M4YOJU
AzDb/THW5FhVvsch1cZ4csZ81azAwRYJd3wto/suMrQ2eqaJRNN7Z6yY8RB7fhVqRW3B22jvilFd
rkq7LwSAKZQ5rQ6J9VJBW+w9vN4zL9jD6u8Uc7cO6NQExY6nn/Ox3CgJb9OWXwBWII1Nv/pE7Y93
+QRr1euJ2TapWn28EXsuG19KAlCvxWTooRQP69lmbfz+w1iwqK/44DHjHJZ2Yb6Z6mq8kyXciFCN
KW2w5wndZCLRKjq/aMvYUL6AN8a3QcLcK8OnD9CPATobZBZgGLNQyKt8E7lSBIB9PRNquAecPrjg
rcXYdcIzN7HqY5orArPg1qoN8YwwheP4BM7c+JHnBJIoHoEK9XTHsnMHtt7WobQaq7qHAz+LVRsH
MMhFhhKvwbPHMAPO/ZVJ/heXl91ShizR1hU+euH0PCy/AWXeNfzLViInp7Y+DIURKT45uIJYXmK5
ahsAOSfvqqyjK8hlQ1AWdRguG4ApJNFAuetK9/sqGb5p7TqWhNS8vlG5ejPraA/XW59cirN7AFQR
KFANjL7PnXq9yQs/ygFN4g7/V/fSBxbLopf05T5i6YxIM08+xpU4c5Yl3J+1RxRzcThewMDMj56w
OfkY8PKdt0zBjy9KTsOvHPOdVJGEIquD1P5R7hRw1DxN46UWHf/wXu1EoK8/H6AMlAzZkfmlMtXl
GpxR+4ylhXQPCbC5aFhJmT9CW39a60/OqjAGxy3bZux6aU+NTRWh1TezLhh2lfogFyy5TO4btGft
G+C3A9vpzoRdViTnev0TZVDhfArDVR97N7lcZCR4pwgOfGaB1Vzj2vqv0VxLQgd+uyFWNOIcIeHS
H+hWxQE5IzcoJ7Lg8ppbM+lvrnQXe6rMVoT++NshyxGrGLCWVDg4kjUXS7gneow5pHanUxPMSTzP
ee/Vk8vvWwdSWs3K4abnyWZaspnPpgxbene8WQzbnh1b5K0QbnllenmKtOCmCTuu+Zd+GRhj4EK9
eaAiPeHHXk7AF7XDcNkV4vi+La0WG6gIVsTSQ0QLkE4N9Cp94YbUD0Ettm8pfApTQXgx8zjbeC9g
gF/rJCUYQj5u19z+E+b0wrFesjPC6voEd5icE7yTUPuOEhZYv7eKl6pMG93Kc18cx7NNsYQ3LI5q
34kq69xJlOeNLQxu7ANUL/G5Te0XibRpof4X/YDzn2p7PrUnlj2unjiiIY6Y3XJLvX9uV3Zffglb
mevhaseUI1okHh2xj3QREAlFVuULcUPwzFdaGA+qJrYp277xbcS5KsCco9Wk/Abg4PFfab6arwpM
9hAMjOZQbVG4ZRtWcvAEJ3Vj9eRbcthVStP0lMWc6qwZPzXdHXW5NSVANKBnCAuhqel9prUQro/a
aMskglBH4HDXJQhwJ1GfAg4jSYYkQbpv7M2csAdE8An72PdzXo3h+ka+C6xoZ52nXEyAmkZI798U
YI5VXlUPnmJdJH9LbE+dmAxLvmT9WFdHT1wsjA+0CWpFp2i+HlFlRVy115dGaDhjFWzahFZnAC0i
Z3++sdTRQ6pqHUIitddJmv3D1HmZvIEkysGU1ZoBS9GsCzpGl6tzyCsGFKcwg1KOBQRGqWEcBFAi
msGB7N2en+iBfq7HTnkLv6P9Ooj4wXo9pHrJq4fbR6fWvgrW2lSqtSGECQw+d+CnBRwvfBQ+hjIb
1Vww39BWDSioqZ+igUtgWjFY4nB1DPYz8I+t5oAsdjlXJIllImsl09aCpNlXlRbc5XIax0dbTIk4
qD/VZZruXv3LbUShZ7LOxX51o9h4MpGHyPBUkum+RSbt0RnA54sjNKoB8YpUKtCIMXye/lvdKkEu
U3GokdVtCOMVG3I7qtUnTj4rWzbWUlIuVZTLLF0DDCeZ91XnYfUqUvsYo5TlHDsadPP3JhHApIDX
XCAL6R7szHLAM6UJlWJcCzKainPdJ/hDThhLgCui7NSFy8e5LHkTTwEcWTHmEGHEsAn/1Xkmqdcs
zIS9bAKydQamnX4+8hSM7tmvLSQ6lGweQV0Qa/CzRJKStPzAhfYIGborzc+WKXNWfgyiZqLocPTH
qyjoIVBFwLr5e37kw/4TnmRAJ3wYB8Czog2XfUBjJkEIpY8yX4QSnoHziYu+6ifAcNbha03ZtznL
dE7XNlhvsFSA4D072DmTLG/S0qFDsaY6EqcDAYdfSuldwtmc8CXqMLE0YRg7p7g8+nx0DYRAD/7O
PHA/xeQF3ckPRgQwqkIw0tjstu507LsfH8MsS8l4Gd1MhRFPHrUyGrPawVucBbHV8QHyHlkAY94x
D9M1wyxgcDX8pdf2eUFaNzdNm3Wau+oTDG+Og0Zga2T8fCn1GSmYaOpeGyQxZOXwzaljk6CJMmNg
Z7U2zfS8RB+gyXVqlel9MXdioD7jZGAQJgh1loJYidkHBsx8qZDue5PRHma87prKa24DQVWg4uWZ
NsebmW50u2VRy6UcxI+sZtbYuCsYm147tNuHDNcYBE1ePH9EMW/pLDiRxMPdM2zm9safx5b1GgC3
eQeIUaGyIux19xbmFRFJMzv6DwVtGid4JpcpBki/8bed0/HDIaqNI22luVHidHkAweHupaBPmwjk
D1VGXmv5zcXIV6Fwm9NG8QzbSKcU++9u2oWoQRZHPQP04ZOKLcxOw3TZY69yhES9gTZ+B6UBi6dG
ptPxJjV1rC/jgtG1hdH4XAjJf5jguzuFdCNIkn5mh/ZoSK+rINPTIKq+/A2s7ZdMffz37Lu+7mrl
w60ROu7dN2t7+y5XGkHzaS9n7wsM+I0v/3RBox7mXcVn2xyG0wsPqkqRBqOJ/aVBRn/wGbOUvUbL
aIJuyuqkgMCOlmCw8ZZ19z9eaAzIttls5R6I43AVacrKkVAi8TSJ1GjhF9QavnJ5f79ONalf8kH6
vP5guVpnFBbSRLlLsXYopDabMdnBj8wkQY37w10agN4YORolEy0NCDeecaZ7lA2cSg+iDtN4PMa9
PANd4LmMwrvuesZIb5jlNTz4dN6cURgz4PqQ6ltlt0m0r9dQfmBUydhbpRM8MKud/FlzA3lKy7vI
/ODghsCePYYFGxr4toz84ThCUCSLAVDZGb0BeZ3HAcIoPcZdaZD8xBN4YXZGIZM3JSIibkiT1flo
ibhZVB3j5aaDuEzmHcZ1hL0vb+8M5Qb6RHoosg36Cp/ymAXawjdVd/X778ZIcykApsHaW8x+pT9D
rt7dL0k3I6YVU1FytcFv2LH3b0BcA9o675jAeZ+ZdKznh+kkE7f4xenyRv3Jf0y8gSCw/LDVGgcX
2e8fcBLrN7vmfOpdZf5ZLYTkPzS6Op3OoPS8UF3Hvzs/Pb0sWP8ZWF40J1U0Zd18ApOpZIfOb/7o
jxkYeyxByIK+6V6SyqKxwqWmeOwLcSzqvTAM3JyyQpBSJx23SDyE5xra83hyBMM25fg1lKx0O11q
tiQiCj81X0ooqSSLZVgOvRAtLP/7DrClM346KhLBrS1PPtw5FAq1DDMLNQ9Z/PtpTenTUNqb+t3T
f3JGm8qIKVNtfi1Y+A9+OqRkIf38QthzRpD5FjtuBCa4sculcuNkH2rROqQZ25BbG7FAez3h3s+M
VsO8u0kH0vaVlUmN8509+n2eFc/SSkfkZALYVrPRUlxkZGerT2Zf8TxQKNjYoxm+OA7fY0CN0kfn
XEZToaH4VF+8puzsXgIvxEmoy/o1IlWfLNb4VLBy71LYermgI+KbPghaZzOoiDiE7FRU9SYJgDt1
VMjuBjSNIrqQK94HE3q7jQTt9iY6BdCpDWgFTzzQ+boBuR7RzEIpVUrvw4chRFX7Abpxe4qem45Z
WFgjYq5Vd2fdX60P/E147JHyz3gxuTNpyFkgH5Cfiegvo9Ynku9bd8abKiF76MDdn6yYMxGTit8L
CDKvOBEkD4WUCjWUw5Z6f2+tezLiL8aWmz09k6jm4g0O8UL7r1JKPqcyws3uatCucEUH1s/ocZG2
sVkiNxSgNBKD5Ixov2SgZNpY+hNabunqjUFTbkWqrXJ3AbRGEudGIRjx0zEuQRIuHUN7aJjnjvV7
WuPl1rrRGbGjREI79+hhdz+aeBsk7mbN7tv4xmMXJb2B0QcwBOTX0I8fkfR1Rx8B6w1+GRomderk
9YbJWpg/y+hIzNR2eyQA0UrLCAaiodi7WSDPQjXx75RNDFtJVJHN51PZEIPogw/Htmq3UmsNxOpC
QUmoyewFxvofMuWRWYMmCoAdMFCUF2iBdI8/diq3EeNeL582c+Xy0l/wu46aL1jaE7DFuZd6WcMP
yKi6nz/T1LVZeT9DbwaTa3MUbxka67BzNFD2820bnwUgdbmz+QeVQVUZfoU+Wz7/atNy6a3rFzOO
N5Dy3gvGaqhnmdDrDZr8+OevWj6l+fDAT3YT5KSAq4LrPCG0wjbMooriGeuyH5RjMAk6KtL3FS/j
rWHId41hOXzTemk0OHwfGHYsExYxjCvMbITw6prOHLwuBe2LWw8xRAKiDD2zG4h6Lcq0bYmkGZzZ
K8ZLYM8QgB168vJTtVs9t7MvoDDO2AzFogZTUDBnqhrxq3QE+FDONeyQ0lKAj6yYKUg1ht2h2u+Y
ZaYyHQARxOAQonGtMjzJhNQWp1rtYcghT0ib1Lk5u093Py/j+SRcqrDjS9atLlp5XGVrUNg3buYh
BDwVZQfdk0/K/PrzLgNHAE+8D9Y4h2v5FHg+8Y5+3z608B/vqdbeiJ4RA/avfCpvywkqKejT0obl
3skkwaLacDasonyV4W/+qYzCLSv+gIQKqxUw15AE50448eHHfLMBl7Sk8padAfXuPOBIuSlilZMk
DeBeObcRTAJiBjohGGad/86XPpPlmfvK+JCU5++Bfsvk6oWMP7NyLKR08rnyqV2POiWSkejm+ij+
0kMwaPK4bZxqwi1F+C4GfLcHqILwbGLpMj5SP2S3C051hoP18HqI/s796BPB1O9T/geqW29I/CKX
rjbxeQNYYLHjyYjm0tHyqqNj73g4cUnAMUHqs+MwQ/orRcFgRClQdDfKOxJMn35TtVm5vDb5zHx/
eerdMaNB+K9up0dkLTVClbuzguOa/pm4zaxiExsyJEu7OGT6RLjks/BRWc74PXBFDcluuAJpy03H
yO7B+KxRFpzT48ZvtqIBbGQiCA3IOncNz4py1jUC/QvEi+/Dg2Co49LXJU/Z96D2HA/L5IKSIfvu
4vkAw/B1eb1CYmUGhAiQ01uC/AeIjAqfaUbUJtlEi22sq8na4Iyh+De+R4iPl1st8HBjBpOjEPpC
6ct8s1tpT0O2KYsegenzsOIEuJXqSZJfrR/jOtxC1yokgcL32rq2ZWpUC9G57r5VXJbQAOlFXoB0
td2woXNvkSBZXavbGDplgMAhPk1byGLdg5vYtln+0Oa1pV2JQX/NAbLNHc5XoW+qYhRJhVh5tsTo
c8EXEO6ylcoKGgBCTadCxhxi2dpurc6IuQdLTG9DEUt9XBI9+9MJObFLBYBA/aB1IFUSpztLYme/
2teOLmJlOSdnRzejQPZExmjYSp0ZKrDTMc0Pxn4X5Cv2PNA1qAGivZDLp4AMaV0kGhHJX+ZEXdpY
4wRszo1ifz2Rq1COCmue7aGPsJn+5ZErTdjY+Z7PbhBSSf/jcH/8s2OYd/sopLW4COUIX6rDcSQU
9gn6K0eSI3L+bCokM1zzLSyP1EVJWxcBHuKTHimDD85Fgbh3V2Y/P/R0vRcLldLo3oHIYasmqQnR
g16WZOVKcJzwrQnwn7yGxqjMkxTDMVtuZwAAtlB7hwFE3WQqKpbWYWNRPmRJjwM3482cOuIqmCba
dTyWsNDI5dhmgaoG2Prm3GnvdsN3Ok33ZIdhfCdeurg3q3F9uvvtQokmPcoMn7vaEY1IQb3g+pER
5hM65LVckLam2lu4Z0INBjzAckhC47ngFe3tf/srzxVGSMUyLe4S6ye1gsJGxXTpDJtO8TQm8Uf5
d5UHzgkQJd5ZrcSIwx9QIkRfiilMzfFJs58PVzfhY5RV42oY/fupoS0tv80XnDBqDsieouu8hHSV
+RxZi+UrD0BtAV0VhFIIMXdJL7UnfHCEg2x3CK6+Yea3kglBFRfipgW+B36kslvFFnbiKJj+rrp3
xJA0xzb97sjaWWACqg/2ZqVe+7268KbhluraHpuPLDVgxwBgytRLVZiqe0hMeR0nwhfz8R4IeqS5
vVH528Pis91eyS5nmUC+uSrKL15ofnCKPXyWSb79ZQ1ebuNYDlmvG2LWW8xOTgQNQhalwbqV4CBj
RPkns6/0KOzF3S0DSeB9NmS4YZLPh3YflMHrE9/BSw5kFiCqxduqvfBg0+Cm6h7pLQFZ+Qt8lO1E
c5YEQaZ5JW+i+WWJTKT76ww89uc0EDq2Xdfp3u44xeisI4OXqWyRs38yKSWTAkFejOLfhKhW7Buk
EwYCi5FrOST4tdI1e2QbgVzGMbTQDG5CkLTI0A2PR13rCXj2HqO2jet6q6GGCnQaT5cw+PNr9h1D
BaI/T6bqbiJrytEVV5X4Vsh6ruLUlp242AN260yV22N3i3Fgys7aR2JtBq0qbGc4Z2grE7QZECIZ
XYDzym33QqrBKozZGsAtBg718M2dyziPQuUcMUklQBCyvu6RtuDf9eucDUkvWXTBiY8Qt99u0lP7
t1EPyP2AT/KY+twZeW3Sfz50y3MgQvETWPLZVCnmwHc8K3sdsaxRM7rt0Xhqwn2ScXVtDVutXmGU
C4DHNeU4OjSCMLqSG/VqrZVPTWVUU0Bt5blmfCCHweOxU9GoqK9J6vYTueN7MA4IeMHV+RVYLKP2
ZtzhdkyW7i+8njovk4l3BZ2pHmycJwEqxFywsjng3WI0o3bkALPjiZegYOHGqgQvH0lxJRHCiKDa
/Ayii1QcTR0wpAn5qCxOuzl5HfFnO8sWr3Q6rl89JGifBJOdsWGD1oWLjkTIUO1hxIk16+VADMHy
M64pwBnLl3nNLYpFt1t3LkJX8yPYdr14Cb1v+wLjtqF/Nu/Zg2Jb7xscm90aUSCBG0Vy7tYBIYaq
v0Y0KACb+LRdQ6gxQOMQtM4Kf14XOOu/UET6aQtJ4Gy7voHLXybBMdTg6ePqXP4PfLuzCqG0NtPd
IkysDAl2sEkxKaQKyttAwoH7rJ4GnIDV2iwlHDzVt/ZtsP4Jrmr3Nr5OaLqRYxiyxnWQ9/8KyuSN
AV8AOlqDN//IAhpG6b7fMMVtgzQUdeeNCI9VqbAm1RbFjJHaziDHhr3cLBPrnbkAmXjDuEye+6g3
jprz2fTONIO3T6PmarUStAACqpXMhGMcEUWMaWmpBjEZwiZCYKzXzUevOsAeIN61UOAfC9SPXimi
JjZd3ygHDHxNxok2SyWjA5Xrv23FHP7mAfTFYUhrzZzzUQo5brlNxszpqroBM1iunGvmF+Ib0mXG
5qoyqOwhZhqTlviKznfvKRCwH54gLaFVsjCqNuGkQ1xCdaqByatBb9ApoSTtenyiOutMYjeTlX2h
yASsv7sS8ugeUs3RJr+YSBNiPKcvN90ATy4PCLMb+JfNP9u5FeFxa09KxR9E09erogEdElblfumG
O9jXVl3Rh7VUpSh4xQHNT8/VqBtNuSk2YpBIj5EG1UDGDbQjRfazmRTZIMnStFC3cMunTWMXNIPC
AWW87nfszq/MG3nYcMcZLV8lH8GWe2RTYgByzwha5kCd0Fuw2KuZeYIRkYQWxuW8jxdcyUpHOgxx
CqYvtIcjCjHqNzRL1B4H1ueMRIm9I41BOim/XXkMGSTbTKXIvRsfZq0j+FZIIwFR07ZAhNKATxvi
sSebNDVIdDk41CsOA0ocMTi3LmIABImr/5FuC081HyXYeyY3mEphVlPseJXfkml8iFtXKXatZzbd
hfE1EDElaukUmpKJ5nbkJuK+bBTPrN7y1uwb0kGss6GyTjRZ0eiQZCykokRHNith6DjU7QSVJi7z
ESoMN0HgyuqW+zz5r6j5TnCXA0vx99x2K73m0tqogLAbFMXkt94n2iTqyNxqxsFL2NP0+0jUv14K
RqvjEgplt2fZqThuRh7m4DSmIRrGEzeHgs7MrEc4Dd9SSTopt4adiP2aRhEJxwgdLxYbRkceQ2ow
EZsdXsUFKWsoC/lBEmEcPIfQ7YEVeO7TEoApq2UGO785so+RztgR1f6zS0VRZKlMY9rWV/Nw84xX
s2skqVcwZaYM/+JXgm7EhLe2hbxw5EG7wLEV2ooJQqi4dakr7UhyVuiUzPZII7LSSdnCEJM6wEw2
lwmgjVJOO/ceiRTERKXiLexMeChPhx+F3qQ2uNYI0hoVDSUh4MmzEuDSYF7A4+7BPeyoDRcMOGag
FFnb/UPc5RmNaN/bwkEPQFvM1gd3358vkFRWTgg0EH6lbPsGYRmhpf48tqTLocQl2g2V7+DX68jt
nkEFteiGPsoUyRb5gRXE6k+IbRiU3skl//2t62Ssgsvyr12fGAIC1d8ZTho7jod34puN8XfPrcm+
2ToUg02XcGWq8OHZ4jcDv/Y8kIvAq/0ncbLolPkPcs2B9glv6UaveghN6rKpPGMEqP6rvjrOzKbl
aI7S1t2dNQmw/GRhFGlXFTpv7GeILpg3NytzbXmfo03ok7DTXkAy6CnaPC9y94w9UKISXD/ZCW32
JFwS0lB5qrxgotpjbapZjDo74i7cuw1I0W6ZUnvhdF/NxmGmfziz19McgZ36cvvhxrbUMANKPT6k
wYW+cQUnbhDGhSHejy6RD9QIY0SuKMU3Za/Z8LJ8asONHrfDLadpcQxCpv/AzJ0VzYyHlW0E3h06
TkfagCgqH0++xikJpNCBumsY4+bko9YOsd7ovENkWBvoCzcKTo6sOyCbJ3hxnivuB1WvZPQDA0rI
Exe3y2wjeB+xFMl7/kLzsGqhO1eter+m6E6im3Q7FIchHLuyytsq6d9Yhe+wX/JEPmfMNi9dhIcR
rYvuM3wKBmCaI06s6leAh1o+I2HGZ/T6n1hiroVOk1ZZ03qSVibA7xDarYXt7MOB01DS67iU8cuO
JvEej7r5ZHsmUZEmegrn0padAOKsflOJ5aOVKU25gOCSfsEgVeSILXlK6z9yCeNFqwpwUpsQRxSt
7YMdvoZNLyRtMsC/7KvLGiBAJMZMmK0lw90p1noq4Gn8njSzrQlaKfFiPhlx8hoeC4kTsIcM9nhg
kAEhG+1bFT6ExbtaoPcKaXofenerSw1EuByX1+XNClyukgyM4w/FqLnDr0DMLf1ykYKv6JRQrabM
5pRukQCuq8LlwK+d5hYvsK2tWrpzy1YdT1N9M0OMWTiIi6P/pcyQXvYuMt+vVWsdxRwPZMKuWC7o
xvSn4juJZ+k3jizJQtrs+afDienISuijqHqX2+o8QVvXXw907LkBQEKbV6fWBPfyOuZ4eiLvVOD5
yFOvIzc/CXB7HGbz6bqSkUlsQWJLfdNPtXQn1/5U7h+a1PSilyAqcYmUDbviwmYUhbDzQSNyIGbH
Ye6eTyY93JJsFD43J2Z3HTAEIJ0EWxJ+3KABLGABej6X3PW6pgVwmxJ2tpxImRpqfv1KW2iyMpQo
Xdl+iN39bzuHzevf1GiXdqxPxR+JqXPnKwGOQs2WzveE94J849nrvykJEePhR2m8AeYYMgu5mbEB
ta2S7HT8E/uYsHZptlvYRxh+ao3CTLBGNBTaGLWSxWx06ndhI12rnEwgjbbjLaNAWRSx+2yqtxdo
tmItQs1OlWp3+dNfXnldsTtyKdkmtn3FNprQ9GwxhQUbl+kKz41qg6VO1pBGAsnKK94ZDMxOB/a3
1CyeV6DVSCjn6gwk9hfLarMFDRSzuKv3utFBQ7MDsLkM7REmZWfBMhpSF3T1UWc1uFi+VdRG/R/P
VN1f7kIvPqT712abTIpym6hoVyTJ2fkvxGG/Q5lOW+Z6OsFeoymzvUsaGrj7k6vfZCZAP8jvJGS7
HSHSo6+S+nOKOpYkCbQeNzBpyyeLsA1Mi5huZDWG2JrbD7qeeefVenFwC7ZkU3rCA+AOvnnuHsvL
zgeKVIN5UcqkG979Zobhr6KIGq4DPDFUYEfT5WjKYtEZRXmLp1gQ7g3b8iNcvskDJ14KmQS1pw5r
DqbYAQtw3t03W6TgJl0ceDuGS99X+5bYxdAAedSyoG67jNR7UFv8Y1SUSCM+iHv5hEc0PvH30XcA
J65SEYmfpJDGZM84vQWiH3RHFrfT1+mc1uMiEbhmjDx6xtRSUruQhGXMVoKUgClGr2F7zPBB8uS5
J2YGiYWIq9N9gv7h2Py3q5aIIzFYjv+UE6DDMy0kto/Rz3Dk2zhGb0ea2uFc9G5xoZ6ob0lTFW/0
yJKyZv//Ck3gmkMze/65UiI2+8gNAB/7orS9TUPkUP4uIblpXEbr9ZNWfin73CNx5kX4o5/3+5kL
9E1TZ8aiisvq/1UqmQHN/IAOmltmkDz9opad4bF+hVHlepn3XNXrc/Tp9l7fUKzsSQOK0ia1T79V
vbYtEWcDx++tDjha79iYNUeD8HkOFqSAiEzs8j0QaSEGGDqqRF1e8ewNTtbO4/pmKJvcCG+GXZj7
khlvcPALN0n3hhmRN+m2+M4kWjZ9PvFV/kRtM5FQjNnpVigj6xTsWjlIWkb5Eurw7tE9tUqvepZC
Y2saJXGkMLc2uY6J1WIK+Z36kT/4IvpNNG8tHWbxbHR1x3YzLBG06Y/igL11Hv8erUhvPznllFet
WOC6t3ah7lE3IbgiJyNt2gMN1l31rCe/PR3wORH24I0K2dSc6zSc0rzttaIk9Gy9YEFHaKhn8ZJt
umkPbogOozccps7/WVC6Vq5tbLXuIoA6PLKlHy0nBkNM9omUbtDhQcLFmTfxWZ4dHl0sOTyZGhLp
EeBZZTBsenp9drbTNYURoefomJmC6bD/VMcd3GxxN7/1jL5l51gwRrE9LVYF41/bmaQhRb2s8Jev
q0v0lfneNwU06uDh28FuNDLQw6ApZJyG+RlvpOIyJkXO7tpCRXTaHgTnT1TfVIVJ56JPEGoKO1t+
cRzfsV+FBDF+mlRA4ks3ZMKWRVGAZhU1Ph4ONT0L/IHqPB1HHPEoWHV1jlb6Rg3IGKx5I0UJTrHy
tCLu0ygjTQ6eZyXQAXonGxJs38GRFzLY/+Q2LogaHYbchGvgJVJjtgDa/9VZFTrpvrvgPBDwnf+6
wT47q8z+buJFoLgee5fh10h4gtTbraoJMSp9sfSgxLWLbSPRgtUbf6RfR3r3XXUcbUoKCbPoJm8U
tnNnk0KAGL4aZqOwe/gX9t+y0FP2Z+SDyvGpjD0GpD3lK56E/yM4Osu9LKFCDv33vDUtqJ/2Wxlk
htJViSYI1VblyuHdBe4/YLX1Wmg+4KmZEel4FR0WAjNkb6u1W5RpY2nNugZ6EJ5Rsx3YEAMTxDy3
m6aTvYshr+cC5RILL1LjX0c5WRB51uyUzIOAIbawWGxCq8NcngWyv0lxY++wnl2dFqEKZAgvsbvm
zOXmNq2lY3qbZ/70XEfT8NZZ4XgPddsVh/IhoD8nWIjxxWJoA+ccaou5OY/cDBoMXb2pDf8df1b4
yKbYISWYO/nAWVpHdROJf9LnJcyy/mqBq/7ZvzNg2LfSfn4aVNUCMR2aJ27F3JQ0kORngcMTqlBD
2gOjx9IhHfpETqouZfTSjzBP9o6525VXb4QOvRUPXKW8PA7pv1tWrhFMSI04QTtY+e5rg7IeoeM+
QizBJGN7/bHhgl64l0/tnD8Pdyfkx+Hbo1FpWpu3vqel+rGE9uPmYi7Rv3fRMRtIbCH37aGI7OW2
fPa00ZW3tTnl+/GSMdQ1PTfVy0yByaU9ZTL3fgCVbvu7Gwv9ow37ELxw/a0UbClQDOpTpqoytbLi
QW117RAL704kXSSK1ge0q0QwiLx5h4Hqn+SUEUDX3x/tOpczU1kTXE6FYroHzl4fGL1Q6ONGXl/K
5cuVCBwpfb7dhQtvhUaKoMH6v/JO0/WO0FXIhvVuLX0BScUrPz4o4wbYFoL9Kl5Qvg9LGhVS0d3n
MkrWc2WdZys00HP/sY/FbrFmng7rWoNC0AW47Z9iRpRNhxsDy12wz/O3xHFbXK7GLuY1I+m6RYbn
5KLaAI4FSbl+4lxwNKY+QsuuOIC2GN/IDyhZkWf0YMrC1CzpXvbolBjnrph/juAW6QtFQzVEDoW4
7UHfp7UDAVgGuXxHtDxxRQJBzmFEa0HUM3qYjXM6E30kBNy4Vxj2rWVyavDxi0JtmxCr7XxKSJY6
Vre+yOBIX2dpmhRiHZCc2YQa9kZ5SAVeOA0CiSNsf7IN2L5couaYfIisA66RwmL5JutONP9N8RvF
hUYr7LQEW38nj48XLD7ktvecNXuZMTc+oLlro7fL/XMukebHzj8LX9b4GNlERYGtaZNcTuRErNKD
vZRvfuZ9/zVqEI6t/arC8gOcU9fz3NQxyUUz378o8OudJofJR9Jw3oIDjWr+pDAhs3io83PgMS9m
JEa8d0U7iyHntF1hs9h7e+wSxtK6xtkRLAmrv4bZjS31tjqYf1qFr12VN7nALxLjqmV8Tdc2cvEp
745YFBvZbpUIlXeenGVkGqQ+Z9IISX3Yhbt57cmA8kZt4YGeFTmKjcuu5J05JOQ5CAZF+4RfDzEb
SG3ID0DkpgZrAkAU+bKvw83kaZj7AK0RmuTU0mWur26SaZmsbAsj1WpBUBtiN76iuQRYwzw/yqSb
IoXfd/X57xgz7JhvW1YiIwEn1JrS/vXHLOTW2/QfE1KM1PbNmK1ytoSrUocxgTaePOocAJv8OFxa
hbkWkXXroVGtcBEVIKIypRL3Vhb6tR1pWDsr3fWQh1oq8QWra2/GJY7GlwVYzArhX66H7Yt3JTFf
z48q1XS9RPQdraO6cjJ6w8dc1bboG/1GnRSK0rI7GplpSo01rBhELsMNHJ8N8S3Rv0Z0nnxhbt0a
3BsWiGfxsK/QqyCYSFzknGAdBcI6qUG/776+FQyVf9DvWHsjCH8juRG+BZFPop99kLzDtHhEYoLO
bf/E++f/ZCJJBb8YdTQ3JktcXU0xTwN/gYHwSIjt7/wfipALIPAkH0HapxRt5ikwzpoyTUB35G/j
orNCYorb/UioBYFHCZTVYuoDyiDxchtd/q71G9FZ9bNJhJXIrfedFC1H14411hTbN67ZEN9a01js
uPp23zSd7X0yskugFkyiAPARlbuGrunAO7Av8+YLaMRfBsEm4V1rNt7TZU7gJRBEgIT3m/plapyw
O/eYAisQGTuiNBHwKxoMQBeP5SO6JQ5QL+qPVo6ogbqkKDlmtXCC71+1b626If1GfOwFrrH2c8NX
1MkPECOT5/17Wkx5gj6HZTvJ0ZOPQlqJfc197wPTsfbTv0AtGn4ibFV/Hw0fnep0fvHi2m0+JJY2
S/s/TOqIZ0HHM7wUnmn2Zpd/0uzNp7Z9WwwtkCw/fGKOLSvcJPS5+OrhBbiBXqcvEnXQd+vG3Ts3
uby+0IirwDbFDNcNANT/QZko+FVVAZZpScUN0uFMVAo1chy618zUL+ZV+i3KoBk4itv/aYQj6Xwl
7AywFUx+n3D6rgsb8qLGNbdhdfGgXYoddtGuoYR2zmetn8ZdHF66rEqs/8sFP2O9QCZEu0bVV+iU
/m5KMjFoaE3yIXwa+7R5abdrSRrh3MTJtQL4bEzE2hMOdL99Csi/FOk2hV/0Z1k4QSITC0a8S53B
yBX0vsF+Pqd95GfLpHbHxVZRcwN1uxl1S1QSiepNUcbyYKiY3Ek9gky2Jnnh+GaJIl9TIyvdyhgd
zfbTMEeYZDiSoAWKZk3UjVRJo/1APALKKB81c7CJ0Xt9wd93sNXM2iYPbrqLoU5vGGJFqswDApIC
yn2NyQxOe9i7z+SN+mSRRZ/qcDzMNBobimC0fkgUWJhTSdmyL7bdSuRxvOQQHogRyVZBQ6rsjikL
hNHx4nYfcgf7fBdj7QSIxYRNNOB+X5baTUAYk4kXiiE05NId2FxgFaSFfnrSi8MTV3+YNKixd5zQ
cOVRhtXp4m57kfVctDk7KVM/nN/jEIDBZvC2PZwuws5EF9TRQq4ngJBbX7gw04yX7o9zgh+936Ow
h7Hfv9ZInaslX/JV0KdYh5iUqG71sNuC0r83SuxRS/wBnwzpaTvZiBzRRA4YjMxyXhFHHfIt6UA7
kJIZbX/RJqoY7+n4TbXLHawaYo5o9+cKE2zOjUTSp6Zuy2WqIHZyjhGTfHheYtF9wtrFOhtTh5nf
ou7e8K6MoB5WQFPwZBf2WQ+mOeJYbY6QhANXB4GQPOR7WKHnneaaT8aOZBZ8CSmn9n1SfCbaVuUh
aMMXutOuoGGbFKM13nUZS996MAowBWJ1QEsD4KhjvmTtc7/pkohESKcqxyOhZcetSbWfCnCthXuf
JnXyE2og33xci7j9Zs/dN5taOLn2AxxKAF3O1cRxTbeKfAoeeAfHVPRHGDD/AwPdVJJOJiOSfZpI
6tUFGR3R7OWlrzVLjACg3x1K8Of5iAms5cWlcESNPCTCsu6LaUdhjscY4S5hW/Qq8inao/Y3JcYD
xMt+VOafeHonOXOi0UOXzVB5FhdUYAuFyWbckCt5pF5KatLVVAxIfcBD40NWNV6dxavflg4VENd5
0ynbwpKeijSGvMMU7U4oY3Mqg1zexTOkUfPGxGVnL7a/DrlQic8fukVq90WOFrVGgfa27cdAoXx2
5s370gUYM28d/MkF5gmJ7Ig29dO+5lP5p7eN74GvOPAWI0aHO0WaWpGyhrZf7S+sf4cPs2q8ksEA
DuI6JU2eKJW+WN+dMPPqRMO59Pcob9RuC2u/lCjX2ehjxvsd4PM2Tr0fXfHhKVzO9x2Y6Q2nljmM
nTR3M/Sv6lOMf4TBZfOcnVE+SM+hFI8dI7RIc3RQhf9twVLF5CBWWMIZyYrf11WpES2X6lgtBJdG
shhNZiv0mTIoDcJnVOOyK+QRF7JuO9E9eaXBzyOp+NqvhhwEoY4TKw1iMld1RrcPPDzPhyK9NlV0
e6mMeVkxWR1kgoLuXfiBaFyZnT+fRshpIk16sQdLWDgSh6QwnV383q2YCpwn/JrDQ/QF4inogNGy
937k+SJRNpd+Qn2z7NJBFPZPgHtozAigg+NcgRBfvhQpPXJwYHdFUYiC2G/rfhgpXFLFgmf8rYlZ
voROka8HMCGZIjH8tNzBB7d2hqre7245/JzbeoYu82T5FE0Ym7UyzdznQ6Ir4zxygo4DuV96zmz3
RG846ZcglICOjaZi/rAgEJNO8CW5+9tM3F8IdtBtHv+sWhOg74q7MSgew8sXAToH/8ng5AqXcRAw
Vm0j/ddBhY9hRmqkhWl4LMS2NTcTUNOUXTbVYQEJClEobGPaoagzN2KPQNKnExVeAofwMB77VVwZ
sbBhAiHPOZVjmXqxCsBi6Az/lPkxOwJh7Sim/4r26nuWddx1qFKeP23dQvLP6xkWEqiDtkchNPLX
5DQC//ND3FIZDmiTW40AquCQPTACLEvGvn81RIGkC/ClM923AvyQ1x9dkDQGyV2hEYNJkgK4DAOA
N/nw14MNUzcAe+kaOKRBtQE9dF8U4zjTGkSe+1T6fh8Oqvm7xXwJmDlH1s3euo5mGrf4EL2vHRb6
rlSDmadbWWqyZLU8wvGyZMWbd3tZfQneszJMDzgrqw8xnmbwttrj/VI63Xppp7oXEuVMbDsayN5g
/BrNd7OrflpBKFA+dY5CD4r0d6qNSbEBIBBXcmy7maur0tGoPBgsDlPHUsTlftFWScXtiC2MmZ8y
l4U6uOHIMxHlBS8y9isreOyUBkKLAIIX4rFKPKBCCKlVFKv4La2qwCBoCe2uZZn/poxxZUTgcvnO
nfSStc7V3xE75aMLfT4Jcu5F3tYHxVJUd8TzgRrXZKOpz8Wr34VysYnOaa0WgZFmr3qte26IY8Co
PAwP6OEWOFyLO1vviSylE1gqhVA1UyiE6b5q91IdXnsD6B+mEp3YoMnEnG8e5HNFK3nR+EZCjlXY
k1KRNk24mJhCuNTIMyqcFUIdbZVnf3e8AhFlM5HOEUi/EfxkGVRdD1eJBhlSbXpQDZlcnJWHvkop
fqcQOZl2tBrvSgvXJFMFZqjcCFAnJ36T+5AWTm1P/mo1PXBa84I5P+2vZnx2cENzIx6KtkI/NWC1
YMY/Dd8VGUc4nZ9C6Vvc8ZsOvNSgwLjf19UVqw91pZUu8yfEm7O01Ta5gj43DkcYTeKjwCk58pKN
kw05fNsE7gxc4pbGzQgdazAnoUYU9B49G9OPc3e/DaoVBBC0xwDGzDUZEk8ZAecDuWw+9p7vEz3n
hUG79AFRTQyR8QC0zoQtLy0898ZTfsf1JPW918XafOdyE2d2xP1e7bgfEjVC83BTmtnarfi7zVBq
t4a5mN+bhpkZZmTrzFeWjvdiGSo5z4LpQWcbONvvZSwKBzQXwDI5VxdaBQYF5Tq+z/U7qYtvFocD
YmzAw30FRansV+rQxTZR1DQ3bko3OngQ6JvEsg9FqCxCuaPY6hSqix55sZwHUu+LalcQntxTMOMX
z2HYMsDIIBB0y/xz3YYc/+HTSLHggHawdEvm+sC8tl27QOyNrDNj1c7JmDDEcMZjfecdGC/+5tVs
+BntoRE3jCAJzTuVEnBI8Z6MhAn5bOD1di+C1VjxNVJjYQswdHqNYtDK6vNs8oKOJoonknNLCgC4
JPMdUhvhv0fVr21TppkRWnjLuYPkdarqPiRugj0JuobgJ81utvS9OVWHqAAczswERsd0BxYAtxoT
Jr5vGWY7NcnDkWF55sBtjck05Ko3E8fVlPtMdlo3lto3NT+kG5PLAcHVAdBchYTWS//hMowGe1js
H5KAMCvVrod5jbNYK/ZuCRPkQMU/nfE2jFtiZsfjc/WIFpUgUsEgIEQvxgpK/q9tm6qkg5ghv33T
Q7nY96hRi71hLXVaPdFgj3Hp5pZbj1kKQhRz1j1WBeN3Qe+Ke5QqaB2w3r37fNHB9juaCvipuaXJ
b2smM/MFlKo4U8A/j90mjYLCWIuX6kFLvthN5WtH/EpjrgUrMivOLGJiAzFqSeUXSsAXpGi+qHVU
I30SRcqfAexHoQRb35MR8i9xPNXU3+zRLZ1dhNVvKAmhALufosD28IAduWe09AvfgQDCz+Gsf4Zy
dK2yz/IZ7M2JZzVLU+NnftIshL812u6DSQMIBUWUfT6z7mpJNGMd3BHbGWGKJL4X3redfNe+9X6f
WugWf5nvld2ofLBYqVV7teQspnO1xJq0+Jh38sj2L4947AOMZx/IpHYB6Z650jF9qwY8E9iZLnHU
waSqG9mF9DrHNJOG19iPc/fpVAf2vWKcQDQLoG4mtxTdaaeAFRmIU/Juqq36id2QcGO96o0UW6Yw
bzOWa1zRPQuVos41KTV/GCJutGyS0D8/qTIIHUU9dm0Uiu8jNCdZCDYRm8sdtJmYpEJ/oxweLZgh
iqWo6ioUZrCqHcYpHK3gcXeoRzwNI9ZaGlYpjv5f+i/qzXQaxeJxybuSLT3DfOiilDteH6eP03bW
YJeJHy3+sCz5RztMN8iRs4p3FDz2sBDRzXebx5Lq9Su1JOtkk7UiIsITfw9tOxQ2K52qi3uYBtOl
SGyJd7oK7JBsZ4i6QLCNYr4pO+hScGdB+7c4W1/oVEj9uATGLjumtUBvvsoG68oAs0chcw6OSJxZ
8Fl7Y3MtXc4iJHxtHAqNvpqj83p1yxzcVMkNQr7medFY7Sik+bXoaq1LILxj/tidoxkVHkalC6iY
Uanx32E9Pgh9bmI2nsZKXVvnLkmQZi9tJs6ylKZJBSdQbhqn+Q6fyfAzX/NuXC382basPyEdtiJa
t0imsbiFQXl76jKt2HI+orqqKRDtsG50W/3YmYBhCISCa1tsBJvurImP/rntm568vD+ZQuPeS9+m
S0Y3+5mXj49CabEi34XQdWYt6LtgRDPNkq35w9NutG0xCBUP4HYJdu/wH9VOqFRVGJM4+chqFeYE
2OcplROpJ3XWKhjbthGXk0y4ufnwp29ZJdpzY/jNnknBiTwwHQ+RctgN6RTyEf1cYWdZwKuyoumL
BzuoQharcvuaFtKtpcKGU3wq/uPmjPO+f1RMEymvkcFRsdIFYLVx236FNeEplp7A+co9+NK5tJMC
oBJIYtDcMXKmAz726o81l5kYtdOInUmCQUE/a1Z/JR4tuGeo9zMynUuTmn6ao7tITmfB9qn56VgU
Y1dxTsaFwbz+ITxHKy2tj3SM1czIiadjw5avDi3O36kL0y8wgyxI2TtAQtEbq+1NXwYKBXxSRu7Z
PdP65Kcb0Km5jxi+m19qzwpuSnJR7VPuSqwFl67SVkEHAS9PBaN8AcI8hCfjXgYT9E3PSCr6hRva
eGG4aVfiSrGZ5Jn7t6kvvHj6ZF2Sz2BTFjYPHs4RRXMjrRSIlEo4mj4ljNleGux2Sdxr9dJrioRj
RBrX2vTcf4M+f93/YZtpAivtmqufsUHLWRTNNR1ysWyCQIB1efj9xCKNa38+1/EIwR7z5mGZZf2F
dBS8XMlq1kPQR2h1ZoSlHK7AUYjZQ2FgGF9JEddUHU/CI7Y76Jy0bEind9vH1S3sscuBK5jsLLtv
MqKU0PH8Uua67OlMkQ4uu+PIIbsUWWqizafz7r2B0267tJYx1dacaWMtX4JlkaZj8xfYXZeqm/yt
IANIl0VZwYNKoOjOeYjhlmYUjAgtb8I5Qp5oSBQLQyrrVMdOOiuzT9MWF9pjiueDj/Jinrz1i4PT
rKiO6an3FhU9uthmogw4ll8aPkTcRi6RzixY/S8yBjSl4Ii25K4oJcIOhtIVbt5kaBjCVCG9wYAg
rhW3Xb2hPAmcc8hhvuXV5Ov5v4DA/lB1Tc4Xd+uDn7FGqqv5EjGB48CtJyZ4DWpI3/nsuv/HX0l+
LBbS1prlicSuO0Rt65Y0aQW0T0d590tN9g5zIs6cwQkv5hdQE+sgvNG0lbZg4RXCKLOfhdtKsWA8
Q0P3ls5mMeLU7BqRQaGQn1iVVNvFjljRXoLNPprZE9ZIRNBk7FVgKkzqvohq10lWzXL+LUQWPKYx
ptrZj5xUp4nnsHiYA4MeyjyJbsu2Z9Jo6AbrnHevpgFe8raPtokmK/kpfUDuS3BBjaTCDuFQh7hB
0at30evYzMowQ3piT7ljnm+OR823XApmMvUJYfBWuI5bjhorWPMayrqLryUYSuLhWFOEZ0xkbVMZ
d2JP9jvLIoWUwcMQVE7Lnz1iihaWsx0a9Ogq/rF4e32RRWj38jNzh5xTVrW0CGIUpDwe/9/D4yam
TSA8C7wsgW/sxpOZqF4UCuoYWqGW7pwCeSSbP+ob7jQLrJhwpB9LQtCkXkutCeKZcfUtD/Cen/Xg
cdxtOpjMzH44B/vG6+hHpJDN3Bjv8tvkeT67zd0fY9XjoV1kC9SspTWd7HxdUhu7VXuHpHymSYQo
RnWMNVj4UkFhyGf9/A1Al5sEsFNBDqSwi89B/qdAtIFQrwcHV04jO4kjkVfWrigkGXnVGrNIwO2/
kd2tWkYc4B8sb2rCsIlUlUfliyEuo0quFjymO0pH7nyulQUiaTiF0z0a57VmSK+2NjUk34pg8hOo
tFn5P+JuZStWL6KUTIiIxrCpCPUSEZjwdL52LH8+6LrJm4ZTKvX+3IzAjyejBl4ne8MrUnizFgU7
ebJ0smHYEVswuqjJk6QFrtrq+vDZRVf0L/EsqUrQYAxT/Bkpnue8rBw8ko5rzQhoURVa1ueUDqkX
mGYwkMUe7eIfBhuitBF63TC6d1sS421OlW7nyRIGucOVesrCtvCRoV6T13NQLvHiWgqtJ7Oyq/eu
ja7sCubKED1nlyIvoEoxa6QDc9rkfLA8hYRmjtHo93ABJgHu8FSHbU0SsXSBH/ei6zdod3xkp6Vz
JdNjq5Ulg4f6Qwi2S6fZZdhfYAQJC+ZhHaSQRRNlmf2zpc8oWrdykZg410yjjJsgYVb4yrlbgNVb
n0AS676qO2kqafMTIKY0yWSyhnOnFrAd0rybcHmPgN/sDVlw4XLfWKDc+chdxhxxe/q/jbvRy89k
hCHHwq5HJu6SZ9hiTAIS9Q0ZGQW8H2MY/fAdbAfTdfJzoRhAS8idvA+lzS7pPZXDqaq+L6FxqA5v
G8D7ZCryBxjAsId122olfX7b582IIiAvIm6aYRfbghGpl5mY29K7aeA9Rm5mv5hbxcIC+N+51X+F
YRAFdola56zpPdrIpXZUDTi8kgcKBjVGTL7upTLkITF+q7c+tu6xOaz2fLonDQzwHRE6kdc0xn9D
cnf3u2YbOVdOj+wTc/zANy2EmBxP19s4tKurudPRVIIOeMZM0uWgQkfWgQcfG2RgqsZ8r2ke1IfX
sXUybyOAj0RWvjDgGuVmoieo9mN1E09Z4q1nIjL17BUaApyNS9F7ddP8RsQJnyUDGahFYj9mzPXA
Ax0Z7CV3LmxAg214euNgt6O4fQzOg0g5F0hpyxPvAum5WOl3I9/utDPcGvc26adhNinQvc/wwISa
buD8YNo6ioI5oB5F2W7E4S5zl4jhXU4Z7RMGHO3TpiQ/g0Bcc/YAXV07dNwArvqbQ69Y8v3Qk4Lt
9rKJSSMUWrr/jO34D5/Deck0u4FSBt+OsJSQ5wuSPRJk+6e7FmjjQ32znnlA0lWCPyuK4Unn3+Oo
D0JJ6EfJxICvRY3byCthSx70pFu4Usy1xuS6Q8MYxNzwqG6eapWAYaQzCE8UHFYl77bfRfNPu1NR
bMlCx9U4yTbdaNSCFiDWYI886T+u8pbKW7ERy+K2LIAG9WRu0vqX+KyvRyU5iOMXjsHqWqklyNse
MFo8ZvU7K0ILq49LXBAKbrUiIYYriUQtIlqlF+Abzn6/T8nxI4LC1h5TEz6wsq6JiX26iE8CunCv
+5BfDeYy05/9X8OS5KZ19IJY9SmqCeY3EFJiTCxWfCxPuBPDv40iidkzSZAX5SGcV6i4RlQIHLGL
tewUWTMSin82IQkIJlXSqeqzRU2CspTXXuJtA9G7e52+GPsQszJNB9/+ol8uYgX5HixK3ljO1Ax7
SfOHW77aGTx7A9sfYKb9GSw7lT5QqtmFrqOe4qXxLSSCWnlOD2JoYbr0d/tkmwCVPcChv9EZ1Fif
/hZJ+9E53/xXgD0q6NbvfvbvJ0Sw6j8Cg8raOj/DndzH/9kWmNaihX9JLaVvgpcRGGlZj0OR4wue
6Uc3rMJrGLfOLhwPkudfZAGSpeGwMlIUr8gQWKMgwK1n/L3OzlVkiijQFhR81aRP+m1kce9bKXlt
MBAM3uAwrSMCKraj42wT4clVVKhzkRLw1+gY8OAX+fd+190FUDuGP4CBi+SiClov4ezBVMBuaB3g
SfCQK6Nlg8Q3Eht+lQDelIDfed+TqJmQW3G0yuE5GvirsBwvt0R5Xb5ftfvlYOMfF8DD1rqzspBj
2GsRy0PmS0X3BrpV7cct/S7FTaCRPSpGDa+UfUeRNDmR2JqbhAVdmYZbHUc6O2EYG6mmcwZoImxs
0XiRaaBB1UNmuWvShxIvFRgBKZKamXo0Z2cclRn2mPzSCYvQYCJELorNGEhOld/NzH7by+UjUxEA
DT9z9niTxA5fToxs3WLsZljos8/SrBJS4VSK7k7pHuu7VmRkuHRUGCE0Ecjt/FlaYjZYAXm2yiKV
hItttTr+Q/EU5acSXTBiiZ761xLxXhrEKGFgTNq9Ym7+uTU/xUu7RiENo2WSH87zpIOehbon+jHU
fb5Np1SJm1WgeBtOUVI3i2ZwWFHgqNheGsCx1RSRAi3g/AQzxC3MJ1lkJuK0gA+e00USLZJzrBxl
GKVykPoX+Dpbwm6TaO8R1SLm/4FT0eUIepgFANBk8650kZBEDwgRX3aNEfGUCm4idSSRCe+RmFQm
3/vIz7j3inqxwDKv3Qlih36bt4ABUo8pujlvqCK5NyN0t2ss2In/J8cKiOoQOyqgQbFQ9VUvhWsw
AsweFGhP/RwhHVQJkAFaxMJvUbClMEdDk3kFL1InMlYUPDolRTIGwtaV7IGRmT9oMw7WIuTwxInx
lg2gkG9aldBYNWICzb97lktfZ5+P2qltXbjwLh4RAyJIcDqcw8hmLwJFUza99tV6h3xOXBpevtPV
K6m54nGmJGJt/V5F25IeKCgZEZYawYODXyjGXuE+EFscdAScqYIagnbnughlDJ5UsSFo4DN+y3sz
Av0MLYkzFrowXmO+nAUMnzk9+bR25My96CXiD4K+seWJwU/mx92sHlo205GlpdN8lkbicX+F9LaT
vJwn1mKDwur2mUzJpaLdQrm1Egmpl/QOd4lkFCR/PhDD6bBRc2BxpN8N3wa3GmCzR/DRyJnHKy+8
gYwAgaexcqyfFkaobyKKPWXjREBfPeooBHz8t2SmMQr9mXw5Lr4yNyepk8x+2fln/Q7q2/pk9QXX
CKNxjAV8tOGRxiDXT3Qi5aEmse8UEd6ntbXVFHDRa4ay34uGkzoM1/6kS0KNuM0POqucmUW8edw5
WMXJKX8oYMrrFmFUvLEmH20JSG9X5UoK83NaYf4heTeQIRBA1BQNYGCJ4530sAzyWTaB2vfMtjX0
PRANfL2ezQimYu1OP73dzubub/Tkg0YDmbfFfM6r7dg8xxfoCBvn6O4j1uIIBNnVkqHtzNi7vwa1
1pj1CvMHciYm8na5Zkl59VT+MFQgucE6D9nIEGbnvX87Jg+cKNPsC5eS3uUe0ABVRvgOvWix0Db7
jjBBqAzxNleCFtCcxkngJwgGxnxf635uGcnI20h0Vh1TVO5tyiyoNc1kieS6n+Kgh4Wo4jU5yoXf
7yiwS3Zz5TXACqf96n/fkxmbCPrV62L0JYYOzTsSHq+m3xeMLRULgG2RIhWZk2znYvb3aBJ1QFGg
IunDZqh+NlLx5+qjwHLgJ6U8LmNk8bVUMAUfXJ7vsgYc4Sn4+J5tLmOrRxM0hHDt5v/hVEHxGmx1
Ok2hAzNrhQT3Hv2uVK4eCktOLtZRQ8g3wSHaKkzluG/4iUaE1oHdbK2H62uTFN11VKQrY/Ym3D8W
dg5E05HJD9KpqNoidWQWKrYzII3P4EhKT5qPdycQn0QhYgMhz3WSdViRyOUt3z4k8SRxoAbH19Ss
G3U2X8SrHXeQbLeyU9Wq1+xH9mFYpYMJycUAC42Mw52yzM91Cp7HUhg2brCIvhLYmY2+/N/7a4m5
cIVNB/ZoQ+ao+HHXgfR50cWfPjGw/udjmDQwMkKHG4xLDTNm9L6wSKFYl3ak/13iqEoI5TRDmzV5
PsxWGVec/fgZLwmbqt8qFflkLi6GesQe30PdJRyWvHKRAfFB3cNLhoCPaymzwR6O4h0i7eFcvnc0
75ZbUutVP167oKpX22Bk+AdWYSfEwZIhcpELxdgximghbXh7I2gKJAoUD/qJqlOyrEDS2b+7/O9W
G2dVfI6Ka2YMGeznui2w2Akkbj2C8ZxCQjf4Bba/Ep5lRsFSvh3xc+y+BBPXfw5UlHd6oqaPzvNW
9rqESCog/++Q2qg/ymOtdWV9WYRRseq5q1RZf0uNbjjLvXkCIrZVljk2GaxyID81Sf1KZvcRE1w6
E47XddPCRtqIDubutItrr5n8MJJOob54eDJuLYZjX3/tlTp+oLGJKyKfB/EM5pSMM5CRV/457tzJ
j81JjYZvzp763v6qytPVQvgez853WzHRLA8RqvbqWsF1yhTu/ZncAPVO/jk2xo+NTEazXfVDVxbm
vwpg6h2rOVkcolgBvZuVUC2ypfQNxXnn9HOslsLrsZf33OuUCzp1b185wGjGg7RWjDBjqiS1D/7A
yvq34R7b9FJvqAWkwAmYPkX3YmF6DmiLPDk7xx60CqyxRz9zR1efAScmn2TQcqHGajxeqqk18aBR
eQAVrwRmu4iv7HSMMU68/3iXf56CxB3rTZv99Pzahamh8qZzvcIzN61kOnRqP0PXs9qhQtc6uOQF
ajjI6EluM1L7KS1Rlzm1PU3oFcqjfbKCvO1GYEifN+SUU0+dNEkxhg0BlufxAYsPew22eZ6Oeq50
6zLH41w7nqNwfePDX8iy2CNBMta1JLdx1ptVQhhStWnRxevDq5QjqX2X8q2XQZwS8y98/akDqEMG
+pz5FRcoRVXgCm1uA8Pe4CSfkMpG1YiJxeNWKeT+TFGw3cDpQ7eK/MgcMqco6yrGPds5DjrFk+A1
arO+vkRPLtFPFdxYy55ZyyfzzUnJ7OSrHeQ6p0VscByZmBTH2u3HJL8JJ1kLfRM64BOxPMK9Glk8
8EiieC4LFEGw1Ea/3X0yayqLHmrdZwHp+o0Mz5RfiI/SJnZZ55N9YEeIQjQCsi2EkgO7zcXw4nqB
muVx52K2K3P0/3m0PivEzITnxe+ZOqWmhxsbzGvAo0CTGcnYcnZbDxRCLCQag6yCH6/rY2pfoPdk
5qG77O7hgfRjBBZYYKzlFg8xtSUawSOtF2WgI14qPq+xkg0PwIrW3pUl+cHEkxHI9K0LB0HpA9e7
Ozbvc9iQUKcdVwbi1R5795BXCmZ6RtibsvIsvdYV0Yr9FDuJd0FdlcLq9tbpJ37dRVu2F7J9bKpE
Ahl7+03YjNoeptNBU9U2JEvbmxhSjPfyCXzqg0dt/nYISxESMwIrJOZcqG3Ohzwv8MpmjNhbkmOi
JIQjKPQ1aYoO1EnBckvpWRo29xf9ruGFfBIhbpFazWDn8EpEyW9yk6zYDCHEexpGVnxdXZnsxDeL
carZbu9oG5/GjdmS/U4z/OMTBuGP3Xb9h1JxX6MgAzs2z+ljz/3gBHKE3Xi6sNTxs74iybdzg4Pn
c038qr1QYJz/CHR4tkSENCLMQOhDEq4IgBlPfxpRMbl/bsetEeSo8GH/H/veIiElwwW3JiyRFx5Y
BOBn84Up5j4LYc51A+exxj1jQJ8lYb7EGb/TSZjnRuavb+PPynZopvaVOb4OTyNy9aGvua2bFbqC
ioQs14fUwd4oEjhRGzSoJNYgy4qhRGfrQk6zwZfCREx4RtZmSZVtEiF7zFQ9faemq3aIhFZRxacI
ZIkIyeEAlSzJvle4FGCh0FX/03YbZ++ETl22AhzweQvq2f1/7JuUEhOAM9YzMyiV2K+YF6E/f9Gc
WP9hQyx3JR1ZiwKu0Es1wbI0E7ZO4Q52tfkKPiuPa1Tbt6E38xHNv9kSdeRZBiBtjKm/x/m4tNQR
I40oFC96TRXgP8HQso2SmqlPkkRgpd8YL6d48Ay7lPGXxv+FuPU7fPUhtCkxAvCfWsfCV7MrBWKO
RsRTT3u53cUO3uzbKlWHgbKBFnIe7AICFnlieFUOJggcj0T28d1AolVQmqebE3hHwqHeMCYgW1ro
UkhEJ/NJ57yQpFCDmvs/++7eZ/kjPjyPyBYWboj6lTgmqUP/rIhS6es/jjCqYK80bs6UFp/G971N
fMTY0VRv29GJntFsW1cO3NZkSABwycYsJ5DtCjyvUHc77PGbcs19ySl+csM9Bx0YdbNjADwdKz6K
Y00vuBnOA8XFQWDROESzqdBrAvmjgp0Qzh43utEroNTdfOmBfSB/1wK/N3hTMP7d9aAIy6eqgiiH
ZDpyTH0hetSjMvQjyqUUcRSi/ToKmLlhl6YSWPbaJeNu8oneU95uK6YQby0FkPtuiUTOVepMV0+9
i3LnEZbXBH3LxoEJCKsng45bIWRxqlryE8kipbZG/AMEK4hmnRxY+Cez/67fQ5AXGiqUwBQesiIJ
m7Df/Af6DDzBXIHVf08VcRcrtO5pCusWi2piDs3mUZSSuRdBgnNqkuUi+SDXbTwl+vSdji7qsZ9p
C0eQJ30PJjgY5o4nAglSkYCb29PAMx6/pb064OIgY1bm6FOyh/dDsQ27ssV4pIEdpnbO8bP7JUUD
PbNaZqGPbvqljyK8l9AkEcg94tm3GoziZOTFgApgZDTrsKcjMvMgm3BFCTNzfdghkgPTw5R9HHzW
vT2M0hGkgmkwAswa7i4bI2JI4+ZZEmXb74zoI8ODsTjr/C76tr/6fDrNoaZI/89oZzQAPNnWmG34
xBRee8NAGwX4N0gVuZJj7zxenqkSG5ifJ39MfqyylFeUDIDTqkTSl6oKSV25wMglWZNzowaHehBY
231LBo7Rtrqva49Ownc8IDX3JM5THaoZSgqfJuFCt/UolTFn2bpoT0A5jxsgSVfLKgboW/R5zNAJ
p9OrBkoNjHxvef0llAY8gPdeP5DqNz35xG//j1NTFoTkviyDbbbc8jkSqQnES2vg1EZ9bwv3STXw
uxQcLUOub9ATbY/pZBOQnwPf0q/NSp2SCxIaj81GT7U9ekj2o8GH/bM8aIRVe7jPCFQcaLugZH+U
PAoHzT2WASwQqfT66xL6J4ZIJ7peoqVoQsbfJIYnyEkiyycAkxXqi5hctmu0cMtVBx9F3skKThOl
ZUfaGCCZrankdO8X352FsqfdxSinKwuMalrNlSk1p9dgdYZJ7zCAB/MPlW4Z1rOaVzz5fbkc43ln
mPKguIjk6e5wS5wjm3pbgixyi4N6sMoc53XIpIm9XUYwY4yxAOz0+iYoG2jiSTerg0FSt6H7pgO5
w6552ApJuBOvPMW+TPPuDGIjUjHC3KXu08R+1jTCAd7QsFMdsluuRcJKAZ/BYaavKmsejvr7mrIo
8iwNEsFsFUPtbCCB2hDg33+QbfPIspYk1kKfjsAW0X4tTBukeys7hpCDEoJNmjua24o0oA7ZVnAe
NOXQGgO0jom6OY7KO60gbsietXGpwxs4bgG2sod9oP0/ozHNbZQJWM15fBUvCmxG8PbeyttdX5N+
c0h0yJ8r8BoPheI8AZxNo0QRZpr3zhdhZWKjmvCYSrGuOsxeWJMeHjDkg+aV+/zif+k0nJO6BF0Q
YahghVKFBJbcZ0AXSAJJyMOH2zFyPhr13ytVY85RfpgoSn2t1aTqZeMsX69KopQ97YxHnyXsMypS
TleSIJsBYsTf0F1pzpaALdPD5iA4RnWElDLk8/2guRxsIGe7BKS0sLxd95yUyKoOMKvMhJI5USs0
l18oJ7sceNXn4RIQfKDMaj43Gb5c86vkgRVBW1H160l47eCZFivRD0YO2lA4aaiE7CTIrvgMH7oP
H1SsX3DirpttwYS+akx5ji4krxUOzr8xa/z79BHhlKesDa1Uyg3lRbSkIEb6BravFMlwe+rnN/SB
iIIkM3Cl6WuJYMHUGDIzvieKnSKUjRk8PixOiRIE0IZpcweOhqPhwQ2KaYXVA3RGxlJbr7zDW6Zv
GePZted5lLZWVKWSNbYZomuXgI3gS/O6WnHjo7ff42np5/UW4BLwOLDPvv764oC0j85xtudwof3P
7IWSkKJ4Dvk0kt5tU/ZNARJtcf2XOFZhtTZhSuoYsAulm+38HTm0iZjVVQnBBADNAqtyu+ThxrKO
Jb+jbzcyfzqKNOiJdb/uFPxb54vNDWMUej4sZMvMjGb6ZNloQIvOk6MESUxFk7G7t6u7azXC//Sw
X3dvOEBXb2uKNISyBF/zYpjAeAwjlpPQLCJ2H4sMlJL1xGO5+qqTNwezyAV279qsBiDXEBVJQwGs
W6EB8KYY3bHOYvbpOm6UpEPua5zvBhUdJVfY7F082LsYNLAQ5vXxHiDToQIVxz6CBf4Sxrg9Fq+D
IbES01a/Wad6BCqg4c1mrX5l+SfojVJazYNzsufTr6lBO4oKPSzu9N2B5DALnmK3C3XbAqMst99b
wIC+KsAcy4F9TYEe8Dgo33UOzw5iTQTmZSeXQeEeX7eKXiOIWvsoKxDyplWrA+psLFBx2y5C/zqw
Eq+4OV4S/lDo2emc6MypL6+hJ+L1hoAjnJpM5R580q4sNyuAVR0Jr45+0dxLlpNE6t6GzA9iSAHF
WNfZa/Fym9dzCI3mNbuIt43OOH95n01T6Dt2tbHMHLKabiAIxXzBaYjbjpHIpxrEi9wctATcvnUh
xusCq8ZdkyQdbFgHemDJk17fX+Sb8fJS6HEVHI77k9Pjo3Y47IjqVjCVNsOKfOuSm5mwsQYEJHZ+
WSl0iwfSxhbgn2xSE1MQbuWWJBR78Ng6zaQbu8BJ6OUQmOX40f72zVdW5o9gfcraVAPdO+Z/W35b
HZgQIk+jajb8RUgqeGeH8jgld9iMg0LLgWxU5nJJNfVVyNc0ar0ivRXv8ccf80BKUH8+jIzK2whk
0Gcl+/tQFF1h3q3XmrfJ0n/pJL2Oj1B3t4YHnipKgIU/LNTUHhtlSwBLMJzZUYBv7hNnhn/yEuqe
vjLeQczhEgXCXHSvbW2rOXYh2beJTOp4W1XaOLOmckX3alTHXpUjM4tPcVo5a6UZm1YEXOlKseyB
yWGlVKTvvSZaWXW/eOhwLSUCVMsE/t/dpgFLNCbe1z/pPryZS+cKqDNu5EoGG2OOE6Y9ZxtufHQi
JYn8F/rtl7b8RCPmPatdKU1cgW1Elbn90hDQL/3PMVJT4sWrYWlFZ07fom1tfKanLdRF5r70bZff
zxizeiRwHm5mWaVih5HG/fHjHyMZ65dHCcGK0zSwNidimIdAzvg7j7zmQXXkQl98Zfu4961zsK2a
DK51dj2/+vpl77t1Hymv/5lZzVjSE4tWZTmhCea+SzPQOvVs7peOW+E27j0oNmw6NxOnJDsH01SI
WnmiC9NrqnHh8N+4H9TG0+pLXS1vQ1kITUkAPA/xhR88zwXEaUNndicXK5WwItWXTBBlxFkN7LXN
ux6rn1tm6vCg5TjhWVsNdl+Iqv5s23oTu3q88/tpLcJfaZH7wkK2ZEbZuaHAAoJteyaonW5LNaIV
RvRQGD9SMRpivqn+2FtOmCmVLCFRCJAXmG2LpnVfTmAyAy3yCfQ2K2wx7DfT3IbXYxTHUiJ8EqCI
t0idGI33BqUlu53iDbLhAuiHncI6UqUDaOf1lVpYauHiypjxVQ3zFnTWYuq5ovK7gkfRzBK4Fp71
DAJ1djorhT7q1IBuWDt5V6lpm+7ZUgR2aCuBqibjCfX075RSZzTfXNhkauY7iI9nIz8rxsEQe9aQ
H0MTL94KZON7uymJUfwaCTa2FLylQRONigBytDUOozoLpd5A03rEUYRINbkmr8/QZRGfB6zx/JRU
ZMmUAg25EAYAC3CwTywTOyoTYnMYpAEH0Fh49vvNW2hr8BC46QoFarE8RdEiEyjqZbRkFZrYdpXy
LpfnE0fZTpT+4dnwSLOpGlrBZ0kXS3dFYxkbst0QseSkoXkI5hdpDPnu/L/SuuC8wkrgatXHS86S
LWJR8oOJdRKrxBHJAD98Wc/Qu0RYKQVqYfj+BoI6QDxdOv3CTCzdlfN0FtKybqJNAo/4AKImwogb
ROsOG6gVkFSv1TzRU4Ijxz5FVJVyHAkVQN/xmJ1eYkUYHz1EyjPimWKee7ecfbiIM89jR1LO/isr
In3y811R76EicLzuflaDUrRR6x/y5gSjoBhpyfDEp4eG3tCu030uPevoHdljhbQCXiPPM55gsOft
eoiIMmco3Fg17hjFNUPH61D09ixlKNzk0yILC9DgQKFrIx0gyNaxna717D2XjWi+2AhFPDHYGX+3
5g4TSCPHUPvf5Me/Z4PxZ2d1FietQL1ke3Ywl0ZqzJAnrZpPtlgh8lgzpGHUO/MLNuFncpVgP875
i2aYN6wtGeXyrVGzst67xbacY6sE1J/RZXqyrjZFUqa4o4a+qloID0XfAG2cGJCsG/fknSUkpyg9
mQuUPN+6T0bawzNkRtiAbBD8ZbWNGRlxdc/gIExmlG1LqLnEtxvn4rh8CQYM/dJU9dTqRls7ZYPb
OPKlf+z2M0bkLqKReSxJRe4cM5byBk4flGxfknEoqiNZxtR7qFxW7mAzlrRd1dK3zPEzru72f+i5
IRoUL0N+aLvbRGjG2U+SJURdTbI0nbrIvUrs1JxKgTb4rs/UwJimLoPLaFYNiBEc8UWxcNxayUSO
Br5/m5k2TxgP+/2qmJd4oPDvgSE7+vzqwECqOvNS6Lsuk/aYKFqV/lGj08P8TdomKdgRjPrFQBBN
GGuYVmqVt/HHL97tksd836uCCOx0pagPUWwGcVcf2xWmXyM9fWqXMuu8EUDWfDBRRCKAE+X0BV7m
58EWO2raIvqFjcQPHpMFCZ/0ZdpWk8s875TwVg2KLeFIkemzPn4+rzjsHVi1f6IaTtb8GF+8kj97
h7o747RbB3/7stlxEDdDZEGcDFYJ0MGnYQyG+5ZU2fpYIQcDTl2LGVJ9t09+LlWYqSxAg8N7zST0
68ETAiuzOCA35y/i/q5p0k0puRZAjoP9bTqXPWK/fyh8SrJHlU2unH9p1KvzvP8MBuRsr1UF/GB/
woo6nWQGgD1fA5CDX6jJdLZKT1dt2YDdcHS65kvzxA2cWP/Dk2+am5DQrx0Q7cRQ1DAvQ/rH5O2b
tGHc+f6FXKH4maLwZvtL1kmh/WT1jUZP6iyaZHSv5rzBBza+8uH7epyIIJaUNagG/B5MJ/NVxbQb
nqceJJw2WJx0BSYOQ23DupYqDhFPkYK7+UYtp/SLwaoJbrkteT7LeBGPc0zpc6SCRzJHFv+1Q/wI
sNduHubDSh4pna/owSbm7xDZm3JPIDkx8TUrFixlsqc+zybhCof/2bvNOiXKlflTVxMcR57k0QgE
iDL1stdAj9axrxRgPJSfzYY8MyESHz06zhbov7zwD7pfZ2tra7esz99JasnnZyQVgDy6IxoOlm4L
ta8yWAwqCK1PLsQ0y6SzpQfSHjzfawfkJJjiZGCvfvndNIpp0eVGJCOuxQNNJyxzZacmEf2IkoBg
sPoJLnZwnunF3JZccKX+z28lM4tkVosccsn9CJRPhBmKXlbdyqpZf8RoqQGSiHX0y7vDJumbFmbp
Wfi70EK/3sNnP9pyRal2pPZFzsHt/G5SfxbbQVgMKuhFa3L1Xb8v2m85+f+l/hqsqwGl/CateqT3
jR2lu+P/DXbEDRz9vHCflMZkGkptU7cQD5nd1pN2HLitGRNmkewlMeoN98Hh74di/xe0w4nhygLo
aabk9JEyjVSoiXovDp44bW4L2Fy7bKYRl9Ni/f9asD6YTpY5dcjvFtVWMTFAK1yXJ7FlpxXPH5Rz
nru2+N6NPbKT3UnOsKSb4Ka0Y0e1weeH7dGpI1wDY3ZyKfuNgLHl/0xeQNA9Kc8Tt2qOGTyc2cAc
mNb/UraFWPDaKrOpCO7GQ92hE/vKJ07Dh4lF3q4SXuBZIEJC4u5KAEQq2lXtVsCfkLi8h5UT/exB
NI+wl1C5mqzoaz6ow7RMZA+t9O0stfgjz2YI+cuJD2mgR5NjUIL0Lcb4wmA1D4YmpfLOgU2NpMKV
GxDdRg5hyfymc57+2CQnlCglWzpD3OCG+Ba0Lyo3NUnCdDn+83H5uN6xz0OHOuZD3y8vAbuGUeMS
wJUmH5q4WpMgehABzQdVOKexoIB0lhymeNYu+o/XMMjcOEAKJqSUEq2lxrrpnhlzbeTi8OUFEir7
nNs2DK42RAmH/oK5te8dOD+x+72Ilj176e86wQf0T+NLM6bRteJB4av+HxjHxzNnA6so0n++k7LM
A+En4EcA8pwkbXR7MMpoKjuf08+IuLQNutGGy8i7lQGccDLiHk9x21BfIOs9QEWOEKGQvypRnDQJ
di/BD8OTvFUS6zCCEgThxFpxSVzZWdoZ6HZ5wAX0r5mGN4dpD81k2cKVDctrq/gzF1CF06VHXhzy
0vbOUt7Crz+cAX3T4dcO7x9pH0NtVrIXSb5voXGksqf6kad7nD/azRuFxj8JBRKt7hRWhB335WPB
bwO/rthDmChrzbO9gi53OsVLfKt4ps7P7xGyAbKBLejYuveC9G37BxJ5y8W2VbwJ+fwUr47HqUz3
rzs9rWkJgwSK2rnJ/atmZPZyzp5kWVVyEyat2cEgaSYUbpnZLLdJIb8HIMI2EEC/8AIZ653riCEA
Y4lG+r75KSAClRuGTdTT5/ujXdtJi9Rmx2n1zxFqHRwouaPqBvzijnsV0PuwCQB8tzPMfb3Yqao+
xAB5g3jVqB46/WWQEuEj7SMBdgIwCCAHvC1mhXX5i+Ui5NPNhWJeWwl8xEcQRuDbd9w6uoYAkbet
WlGc/0MjhO/biNnjCDogkipGNF61Hoq55y/x59HmRGfQsnONRhOlubvRDmk2JV/BYMXOYZAPu5Eb
TznkE6Z5W7hWoMz2SX6edo2Kq5c6Rt8Lbv9hFihkYSABx0YEagg7/CnQlLfkFe5adQma6nMVGdVH
ZJkJC+hnaiVjVWgJKGwIGgkJno+TiUZGNv3Y2oXKzCJg1p5UvooQSXIbQgl5rgngfe8b6pvpU1oB
9DElJ0OhTbH6tB1fbj8OdJQcDrwRvwwrEMk5ya0kbNalDyY/Fi0emJxOGXRHW4mpGEocjSGfPGbz
di1iMbQIjNGDZuJELL+LGWr+puQpeXq+tSSPfzh9bIW0SDExgG1kR5G2fl41drHPZgzX6I6xraKA
4nNYJMVXd4OS7IhjgasRYTCpSB2s6ACX2wY/H8tk2b6/cflDabEwykvIx5tShvCvLTS24rWK0BJ/
ny+K7wkV0iy/t79AtEM+j4qiV9M9RzYqc++lHYyNbHeoPfT0I7w5LaqeswtAXPlCkdr/xogIm6wm
VPyz5u05vR7HrftYNORkZjKdNFBaCJomH8MZxaRYxwumSVd+f9hGoqKoYIl++/XLDZ/c4kRNffwh
8mU37peTafIVOVuhMU6Kc8ibdYCky/N8aXeYJXXkw+VQN5Ne3+ycWKXVnxcOIU9t4K7WwBHbVxK2
zZYvAWkKD64EDH8P4EjNogwN4aZ/5TeXVYJEO1FDAAfbCQR2uKXvGDxiabIGwrZ1vgAKHMYjxJaO
kgi2BOezsv8Q3VzaXBy4NW8l1jPC7mImgL31NCdoDH4pj/lVpD2ZltFjDoKwtZco31mUkUzTyb3L
K8OuGfCCcUWDsCwe6zqGiv2wEIRv4OMrNMaiqNpoTm6gkQVw7mJSbW08C6eYoIffTRl7R1DuRhB0
J/QeCA/x5DghZw0ZPV05tCOH7S8FXK2ZAwqyllDJodys7NPUS5PzjcivVsYa5DdiBXE9r7RPVmGI
Qh3ekhh/9tzFSTZ4PYcju9vJTXIze1It0c6fX0ZGMYE2525/d9ZkkhZiAnHoNXulCi0YfotLJn4J
WxdowoE3HtXXC5yu6IfHu1nhW4TiFg90+UZPCWAa1pL3URcGcHUpdKCxQdqa/3dqjbOhZoWLnvrY
vJWoXVxQvXFKun3NVrEuu3RimWlE1F9hAANaz0QYGVpi80F2ohJFfwkup0WCdtwjqJmViBBKqdkH
iDJdf++MdtH0aifKaWEKGFgaww817dILThn0A93KmhYEKLbU8FNzvTu1XamXSZvpWmJK7dEul+GE
NCnMcwfSXJ1yyKnHDGsYtElAp/WTacp899vVMMs+JXZVU5NcerM2izvIoHvhrb2o6iivzaLYStoV
QQFLRiWSlRTAN7PiRbHWlnOYX69SzVWjqA6qkWe6vNkWVKJhe7qA/bLDNyJvuhlxycxX8ePKwKW3
TnT30jovN3UOiU1Z5scQYzXQCCcg2sSrBe/tqSJ9UlwTSN74iK+SgnnHGx92VAW+mtTI1hAH9rA8
P1M6vb6gCNjWts0GKl844RS59KGxmR/mPt94bEnE1qaNEzePWaGIkeOSmq0FMxaR8ehWC2bOv0e7
RK2ZHcViGRJQFinb9PDKAV7ImegfNEzq56TgnHLbb8h6xu0lbfgw+uddAz3pAojp8EoPxSGtI1Yb
t4ZxjmL4lnDhqN7UG4/SjdDD1yPLU5wqEG88+LiuWPOZ4iD9Tz4vC55XiAoT7L4sPef8c8Akv3cJ
PJX3rbdYhkq4wC2Axn3DTN7yyMttWwDfGcktP4ccsQpfun+1EUxM+zmRevEP+NtujNDBxqP80D0O
G4Yl4iivA2qf08EyJgylVk/iK1unbZ9hXBLv8kXpW/8h3aangz0WU+0k8bzhrr+B4NmLFMtEv91F
7iquLM0VG2xgOZ3iTOCP/OaGlT8ee2+Ssw27V7LEM8I4Q5TAh24p1Oq2bxvQC4b+eaRnrfQOucEN
j+p4Eq7einhQxLGCFN8eR1c4hWyPNaXC36Lxs5JDwYvjgr8rPmz2PdZMM7p00e0M51Ie9yHXnPnh
Q6gKFmqazpMZRHG6V5SY4bAZQYto0yRpG3qEbRF8NI2W1gVU1TmC8SUEaReblR4Rzi3zZ5NyzPXy
RDlqLYwMM8ky728mwcFtM3zA1ti+lY8n52DOl/KxJ6AVJzD439uEHlsTHH6xXrwesvXPZLB+vVDm
3a2VSSpcXnnrh1wEa14DqBZF1pDAwBi6mDDFkf0ST9iTYgmzdzVlmvoDmXpKFwxWRTHkNCxLOXmX
MRaRt/ilyXsxU1kkfH7eBftrz4S0YM0EQCkkZw17DeqEetG9dtnD81JG7eShrstTywRDyYEuyGCp
znOwX6i8Z4UZICgoI5s1IrKwSN3jAAVMxmhgdfDimq054rm/DAXVk2Q3iGEQvuCF+FXZ3VSrQRbZ
ERPVMDdJwPcf5/GYtpDUFeWgDHEdN/v+MwruqgJITHV2U0FFvVv9KSLS99snlYvdxjUTjrHxgqpb
Q18y3ZXqGYF4DBCHbytNNmmpSEUjiLxVEmCX3V47Z8U+QBo8HxtVSUwJ330CVWknu4IYJhqX0E+i
NJp4TnsO5UO2KKq08BUNlWX50uoQUulUoYTvkctO7CZZsrfSRUNEcK0X0mdrFp8q/TiyQ4WK+SOb
O9p38vpd9DF7/nPHmiT2HnAt0o3XN33u+VE5RrpwhfSiFVRFgwUX/QFLBnrFpxMmV1hSoQftPWj6
3DxzxjdORlBjQDEiQNbadL/g28k+zfQX4BcrnzjIaslXIIV4q9JElWqeusJb+PeT3xRYymECd2oW
QpJ5rL8clpJ9cdrVCnVu74Klzn8OY6HHmjfvWWQ5zNPlKa+lHxvyCJ45a7rh7VXuqEhkkhWymN68
Z08LYBRt9RQ2+3w2WinX6f4c39DlcoAlz6XQRdMVKltoOUa6H6JcjMYCaQ5daNkINQsy0QDCkyOS
rAVQYig8HAFfnlWMwADDXORZSuUdfz+Fw5uvEos6kTbk4Tb4iwdBlHYdakAlCbltNOYSkNE4AFn1
dPXAnzJH34xYmznkz+EO3pKGNxcEtXFQsSPOCCmem+C4KEEBnkkJITV5X4UHxbb+0YTbIaMStjgX
wg6TQLlRveRZUzX2Zzm39VPcLfzyzrgq8JBtrLPDynLAZAPtyHJx3dNcD2QQJXntuP85iVAea/nL
EOGDqsUAoGQgBa/Xko/gVu/u1a91lrdFPN0BCO52zA0mK77V6o4NG801dospS2ZVJn8tnDRXXvXA
Mi4bmsXsOPmdZihEI57cgQqRZ+dzVY3Qc1lb1dbVWQzVuIgIATUF8uMlTmdDNb7YYJ2nadknqtKO
dHyc9BgPKOvIiJrt2vCDHxQ2wX2DrmL0Ya/o68g7IW+r/h121bLKXoloYCpLXVP4hOlbFOxC7GpO
JX3H7XnGsgCpYGAtOngwwScK9fze4EPxUHFhuRBTxm282RL2agenQgnfFSGf527bfI9I3Gr6erQw
E2yhY4cvXhHVI2btnhuBtfPh6cBuh3bwItecTAp/d5TZwMXJRa8hm+U0BxhvjlMRkSIoHE8TkCUy
k4zusbf8Jn0xQVEV4G5SI+ZxlyzfppHj7gewUhBR1NneJWRp8q9NhsV7weE7Ofzmvl4J1qSLJuXJ
vxV5NrQgPS06k3abWNahwjbapk1+dCX9A2NXgfAg/T0p7X8fx0RCnidvocyF26gCxRsabqRhecj0
D4yLsl97bxdHEAjnRiJpHQxbPy95pSzLMUj8K/zG2Y57Mmj/rTjNIJVdf3eLleBPCNZBiSIrzXpv
48Pim3eVEXP5ntDEM0ws5xrJfOMdTsk2bGOV6JJf6LDKhAlf6FyW6SLLZvD/Vt3B49L5rWrAt0Lv
qPKy4p62jmq6nvvkDfBZvv5/CuNXx1Qyr57zaIpUbq/P5sxEzXaAYw5qAskg9q1DtIDKtlZCx3Rm
Tg8iY4LC28S23bUIM5VJ8Rfyu+GezsvKfhHQ2p+7zCrnbSc8u0BRr5x4jcHLN5yIwtOxdzGxXf6P
fpGWvKUvidpaK8IUehkahrwrPmKQBQQBPXKoN8I99c+TZsb7VCTBidLePARv7UC+5gSSM+c/XcOg
6DhBqofn0drVnc8/G5iZ71vbSOyEAxdiYswBiVDkXjmlsGLt90Hzwe7mGeKZvQxG/luf9ZAdDWIq
jUcunu+jYF0ILLEUJss44Go19PgNXHEAO+dX/hfwQUp6/FY2/RZLrTLNUoPYNoga5jECkqJyw0Nt
W9scR6fODaKp2UULMSALl5atENo6s9jxiWc89A64jC4vafu/8P4CLtEAixI/0yKCip4BGtSgL0BD
G767ztr83IxIVx8Y00x5iC0naD+5kFVb+NXDmqVtTVbatvw3byjzovyc7Mn+Jkf6k2WGnfksguzQ
wzicivE0PoI2ZOm8+ruoDxZKJUB2i9Pk0LI4Q3TFj9dCAADShbF7kkUBwEF2XrocAQiuNW/Bj9a8
9qkWJABaM8MtfMjkNOoGF3WrqHwg5/GwDlUpPXaEFJ/V/lJhpRwzETLv4va38emWM47yBiOVUhs+
t/tHgvqmdALuRxYl8zgEaggx+fpaIG+s1B0mcQSyqWidCeS2WD2VM3lA09SnVnffwZDADYONV9oN
oYGolAimfJEqzgUxgPkqVXg6SBr27V7UpfrEj56wwbkyuVFtUV9duWnTccf/jUeR7n2VU2zgIYj8
2Z6RFH+r+ilO420XTbOZPtTD43h+fYihuo63x0/cli0N7wC5ZEvpVGcMS6CGQZYgD4wc1Y3cAZsQ
GKQ1WgYNR24BgE3eJNInsHm7RuvMtgwnsHrbKcTtkZH1fUaAO/RBwkanFI6S21RDXAB3wJf2BHvH
5uwEkN0KFRVjQOIW+0IT8ubCOHh8ljbs26cOzZT+lA0U2/S38wNgXoqUW7RrAdvLQDF+yOYEyfO5
jIhHhRlM5Mh+ExBdJktK6oOQE5cZQJe7ZbKNeAYoPsZATltbHtuJCy1LKI0tM9Us5AUv8yMLG0w7
8E0uqD3xTb7GZp0siR37iwthPr5R6D5nQDZzjk8aE49ZKPgJzmC9k3yV7XViswtm85untmEVhsoE
9aKGKg35C3vwzKdoLz8t1rrTzk3XXO3HJFj+Ah+ZBPdcMqpey8kLRvaw2dr0GBIIQEV/dMBb++uS
0kdfUNG78byRt8IYdB3XmDnQ8/ArjOztz3tDluvBJIlwCfiQhDIM3peJK+3WKwUphossLJG2dfHI
PcyCx+fmHB6rVQslVK+x/VkRn4n5MbhblcohL10fYithEmMSTvkRuILycGGYmCBO93AAK/DJ82H4
iOkiEBMvbwsoYFgGFCuWU4oEB1lvqRb/b2FDrqH3uqJVxkmNb3HfWoD+huRgwHBufMCSfooLOEZG
21SGxzkXsTFQEZjzfpGmO6XZo+ucM8OlyL5Oa0IkfO7w+PSlo+2WyotiUioIfJU6XPEJHJws950x
fhPbeFuWRoQQcO0ICQmQkhcLfLirCu+gBZE5Esb9OJiBk2KTeU1W1AbmuiFC6u+Xu/RLB0kSBZY2
KWFlr1QWObZq8ttKFgAHlO9eLHvk15L31BZ7b8FpqaR51vaxysZOUnEwGJc5mt5HYdIDjp1/ZYr7
p3GeCOcITUnq95WWowZyBryRzzj2vR1bmjd2dCog+mtnoOR+VqSrC8cJyHJ4FbLhqvzsmeZyLAJI
kcXS6nBz37XHrQmD1yDXfWmzT7lAF8jA5lFO0YSyXTsRyY3jCwcvCRdUenAAUNjbphiK5Ha7fz6Z
MpnbsUlHuqpq1dhbcuFJNpW/wwMWNSu0BnTwS1uqQfLxFJRPxzN/pQjJ3YMjGlQM6fAnOiSaOH01
df6vauBGQsPKuBwx5TAQOaM3jylNSU7LMv5R/apHh1DC0OT4OupW1nLMH7jI4Kbw/omH4P94sFva
p31HMxcLMUsjp80tOQ6YVCjRSgzosW4RxuLbVeqJVVtH26W5f3LaXkyaSoc3plsLMAbHJh+De1TO
CdUVlag6e7kRwP3XOb0dWr/7opKMP2CW5N7JRGnF3fwLnG2kxvqiHls4WTvbjN5HtZpHsI8JlmZo
Yjj1bM7ydknM56EDEvqb0nzNloUgg9rsNFKmuFQ7u89BehmbEGruZP5S0BB6cHLkcdIFo6s8WXBf
hpHk0RCncBf6f43j9o61DKKaCQ33VzK1Dly3BJHG2g0XPk1S60Ap0ihAhYAJsWATOEMi75cMln3p
omQiJ0XIg1qH6Pp8c7mysoZquB8t3tnJDKj2RkWvJrYXvl3dLA7eiieGlv2hrloSyGDXrJKVLq/Q
EMa/yWbMoKgDL35N0KH8TC3cGfXyQVc94SrkyguW7lEgT+eav5paJHDQtjCsgBzVQktBHbWXdLn+
XL52nn6n0a2u3E/sleZuZzpB++JBC0P0zYq0Mxc9R4E0tqXbZVXk++KRqF7sSxXJR3e7/7Q79ENU
JFMC+o9rBOGf3DfA46tmTiUzS3DQ+JmPMKZecrUug15QHeAG50b3eUOGTupAEQ6THqy7SQvrJiMJ
HEob2qqgae/267aArAD223QyH5HLrBKbg8wA3A7ZpLw7TxmwQaCABVrmIOaIMj2l4tYq2tv6nYU+
hlNzCIa9bcbNPHc7UkSJ3ox0tIq9lfnhy9eIcQLiagBDJbNsfRnLikWtXnOEOaAHgRLBm7gX9ZBk
gAntqPhegL+7F1ZsebbWR4OmgStBYt/yyMj3YWL+SeDdlr74uUhR0pgYKLDjgyYp8O7NHG8SyUAP
KtYt9w6Ss5PGyiaJ2/r7ZkO8Ax+vV2V4fAJ39hELy1cCyr3g8YUwkUAiPy84DoPQdzd7WRVRvk6a
U2guN1ujQnbLfyQQOaXrd6EuPU6+vv/Cf/eBLIQxOT4qIQ1u365GzMu4+E1vbrAk4J4hKMaeaRnn
Kgzfm6CRV3XpJ1AtM4IxTAHMzXT1of99rzPw+n0rZnCae7T462ujFJrhGlnAx8zrwurqGK2Vty3E
QzCJ/wMXvMt6MUuooSQwvbzrna81XbCskqkvDG8sbXQ2SnNI9g+0pg7aK/FjGhypgw0KGQ4mttYf
mFNIjlnCRKgbsloo1vgZqS9L6KfyCQFwalXypqLtQ4y0UQtr5oje+5OlQlTnGHfO71T3Sd0b9gEW
lnOYg51rBWO0jGyVIJnxJ4CijGbkt1y96nnkPKIJLKMzXPdSVf7GEVzdM3f2qGqDn35iQZMwjYYW
CEf936V5u8I3VxZLY3P6dkZ8zzA8mS4zozswj/90Bx4lUF9wiSqQPO2QGH0AoMcZb5lRTRkr5cQz
UTr1xbOctF/hautMVdEJLP4uAjf702EgjqeAB7LyP/RrK4NX36TWBm8VOiBNYVp7mYzsnhXAyn+3
SMML3h4kyHMrBqp0b2MemFnGMYXIMMb/t3cRc4iplj1mDLuweyxwUoeiIagBiKpAmNKCWZRyosDX
bOZoLD5Xjf+SI7SPcel0fKFTQiE1F892yI7QPPeHOpp+VWK9loI+7f9qqdi9EfbHBN6DlNSuEP2P
zwtAYKN2xtzi/fA8+99eUAjddmvzQEsw7uhXiJM2iDwKszArJh+8Sy81tIzfvfusjwwJ8Nx82+C0
NcChIFeWs3q2vmzXfb5dbiv6bIJ7Rl0rf2tqUw4HjQ7c3OpICTEwZs8wZSw4BWC+U3gwCuKzlNQ4
QyFAQ2Pz7Y4SKIoowhSulNINqVivp2ZRWDZXjHkQJaQR1IePbX3RFnkcrlLK0ypsalV/jCdprN1Z
ep/A/ZDezKpwVEmabJcVeIuynXpB5gGBAtkNJEzK7WCLl/AyBmnBA+/YajwqkYxSAK3shwVfRqMj
JCiw30Qg7BdGZXXzQeUbQoPvomYRZyrXwbTZ+eus0gMHiqfDjtptBaYBYc6qZStg86dTDhggtPzL
0tQOWFEdRqlg2V0PZCAZNd41K94CMeG4NGxhqP+t7Lv9+XXPlMlNUfi3xrrK/H2Jqo2woWH2HJcf
owFUOE8xBiK3gzCUAN0wxB8UQdaP/yEuaegDFx8SRGufog94/HOvplp7cxU7uC/2TqGXociRdPP9
EkSXfLjAxB4RAdppoAXG+175ZLzwZUPUSSucgKzeBAia4INQgo5exEVhD72EyM4uT4V49A/ne6UO
yEiU4V8RbhMxC3mjUnIwHCTCrO9c9CN9u7NxMxA7+vs2upZY6iB+drmGTLWiqFs7IVlDzs9iXzM6
Grf4b5YVBuCkAlkkCye7w0kfu7UHqCoZ1Hb6q2F7Lga1kPBUI/Q/az6TQUoITOwxVQBnMS0gv8fK
QExkuqSbIHrIRpUn0+i6OlM9ISpRJtGJQkMpVT178en9Q5N1XKvHcB7Pf+OxG/rrh1c1SzwvQmI+
yg2M4AfNNT7AiCBJI75aHpv6YThrFRiYCIVCoK0CKkbMeTvpeBbvs+Jp1nH6yYW5ie1r/khNKy/W
+1jPVYm1J2a+eaDTrDlx0SzNG7v4OZhTv3NAKCi3uIxhP5fGGeFKJq4huIF1u9eYAs97kd1a0A7+
LHGs2r+9I4wM6Uw30hu9otLh5Z7V7bH5LafCcEPBDCnb/0X9eVb3sQgbkOl+5YZiVcP/JnYB8ECj
FZHRSrgzDp/d3x+ikZHFrYqB2J0RvcbvSfjfxlwnftiAS8W4OfsYZvrsN/XMsmTnZ7P1DZvBc5rP
2QzryQMfuhccqdb0JwCmD2Amguq7vIgQNMRjpi6G6NSB9gzMUasY//rilY6rCQmupaS3dp7A5MfJ
R3T6lhshanTKzT38CWT7MAjbUrSCkfbYwwiHnj+YfinHrzof+dHmeUlgUy+I/CWTZPDqxO/kOFMk
287UAyOdQCAHdTwsOm+sVTKqeVpfo5dHRuejVWMT3LiTXrn0NAYXEOAljuYHKdFK2dIt/t2pVH1U
9iDwuDabJnXH2ayZkcPN93eKaqdjM6lGBQiTTus5t4O7yL3Id8mhC7t/eYKDVOWlRwdMz4ai+OID
JkPVq7BmIKDCdcXmd2IkAeKJklv1boihF6Vgb0so1l3aE8mJISTXkutuxlp/Uu0Aiky/Bz55CJdJ
W2Q2kG3cvI/n0N2gb+qwpUZyLnlpfm4JC/YiLlO4w3wdSVom0xns1q7U9TD4AzPNxoxmAM3/0nVK
P73Q8GGsaBZZ8wcd0i9WCJnLShNp0OC+tSIaNLH2AUEnUQCebGEuZ9x37eZxGmJUWW+UymBEsaUF
BR6keU4T1THdXSVZv1TusZb9SEIEvh2h2CnTnu5jX6SUC18O7YF71f28QHbT/pQ2bMlLECO3Hyjc
+6xc2IBQhstU55QTTAZmCNbQKJ0Y6LgLE90R3dXS25WtTi+sIQBxNIYpbwHsPXALEY/noHwN6qxp
3ltQQmDe2DvL/L/4sIOohUJ8yOUpsoJ2JkpcTqbUBWJNsn9RgGr31bjaKJ0UNLlVCEMgbK9duzSS
aRw9oi3PxjKlnZ38UO50YPDM4hoEsmJZgI8FdeRB2yiivoVcikf6qTYBZKWE/TzJK7UOp6TaFHCW
NB3zA8hMvyJDei192kAdT1ymgpVBQwSPDGXBC/7+dk4J5/zYdOxGF9DFfejtWjVpJwm470YSqn6A
P5txHZDFDkEZ+p9XR6JfJJZJtMS4tc9nnI53mSH67xex18DTdXcu6rEC9JRt0pDov9Kq7hgZXW7q
UK3OpVOT0KwjNF6E/evz6PD04psqyA7NDZZr60eJs/nSkqkccMxsmoEqJ21YzGJhhrsqPJAnBo5L
I4xY7GMOl0EBgTz3Eq1RXBLYdsNIuzFuZ8uknrDR8naf0J2MkayFG9+yX7YF61f/n7wocFoBjwHh
JiTofZWXy7PGSjS1dSuA1iLlAl7hl5T6lDmpnDLX1BmTe7iJcna9fj0WqKlofB+XtIVb3RCPa+9R
0LYB0zGYia40uoc7JjiurgV/2SMzE+5+uHKVQ2w8CIVNMThEazeZqLwwjz2+aUkgXB6PXDXO7R4S
hNMFnCnUNAk0btTBTf381J+y9I/2F5WdFBsv45zXlNGnQaPneGPv0k73Dt6ZkdM97a9u2h0bJKFq
h8ayq0mEF+FlQ96l0zRnIgacFSAxuoFGZ2tUIEteTqCtOFCuyxbooomdu+o5IGvtxXFo+zuLpFvD
WsAPXJfXsdZIs+1PtvJ6t1GjnfYc6KY4nTayXyqL4ucDmSJJVkpHvvz61bzpFHMuBJnN0vP27y98
5W6RQgL0n7UvVFo4eOzMSUh28Pl7wozm22VLZOh/T0McSH5s+MXS51Cx9889ZvPTp+RFEjAa9wKb
nkIs2LEv/D+qtof/xTejo+DaRLG1T5vd/xysr76w9gJ63a+F63P276ImaFPGRyrHZDJNAcjBBLm7
TmwcH1S2CjEc69wWUrCoQdned/VMgqb9eet7tfvOZCZE137AzvKhudKt6Xoqpny0iT7uGDZDAJGb
MIS6vMIVoiDmAKA2MxtDJpjsq8mEDN21kXD3QcfVLUzoZwgyzBajGQgYxW7zJHImdh2SmC3PPCB3
Xd4zI++LGyBuvWGRWdJnUun2pPCxExI1la+nrd291yjesFz36QcKnBqHdMb2KBxJOsNy8SHBaByv
MfhyT8IU+pDRfrErlpXlESdykWD9pmlySDa9V23ndPl/lsJzw33LRmxJJQreb6EC2ym+/bCqMwHM
Eli83DtVVqGyp1zt0m+e2P6zOlzx/yi81D5nqGLgLPudlLhmPdpgG7457oT3+sEGGToQ/a9aEqf0
sXnyCCx0yDEGET//uXQjiNtt6oBR4qyeLUaZ6e8vYzsZyp9NQcZ6OFme9cKqRoEzqA8BP6KCUBgV
p6t3JLfgx1lQht53dZ4CZZzl5OLR+fh8fpXptbbtEvkncnSn5BE3A7KnxkmUu5kZ8iETOqgM5K2n
q7VpfWY9WPZGZtg+91rcQewR4sz45gXMesJ4hS8k6upzZR9FoiOhw2opS+QuRY/LX4OLN6qcg3Yy
+tCNHI5I5cNwjsxfSj0COQmmUWqXvLMIaFwZdYMA4jya7zj9l8gkktGjWj4B9ReqGG88RmAKEGFc
V/TUT4lyZFAIzJ257k6NYsI7bmMk0Of/eTqa+ci8PHdA9yxhCqVlHuNXxPbA8XEC3/huY5LlCboy
VuGjhKXqbZXiYbxG75LIrZESyXkh/6j58HrIMidLF9A2aW0MpOK25B/3sz/x4updRoBSYQxXxQ5u
Ky90WHMCuF0l+f8oZDJz4iEk00VZkwg0eVdh3QNBqtKOCyD1iZqb2IiGavKjSkLxaoo3hJi8hb7m
aUpi4FYcvuKTKhfytKsfwClug/fUMlaVYoc71gHyoarIsf0YXXldHHK5SDbM3cazubRgXk00ftx4
wqn7D97iz05yWfR6ohYNbHLkYFaqaNqpb15+IIYkjirkWY89pcLIaualUhvsLYpSMNblOYNVxR63
ssG+YIfeaDbcEKQiY6hoQTazjDWBD7R8e/OOvp5kbC444GX4sCUQUkGSgj4YZqNwLuUNXEyN2/MX
8y5LbmNa/YtnfNGIz6v2fW0w0uXaCH4Y1wrkwmdJ+LSLqCu4m90WKXj9FNcTxi04i/5TjC4C7kyU
3LRhXZKBCQbvZHKXbiK8L9KjhEk5omehQZ8JsV1VaLwvXOWrG8mgfoCkZB6Vs4Wg/p+7en2v6QP0
c9FNDS7RUkd8RgqCmWqlBTEKEmKBBnsbzY4Qkk0ZQxknsryTuetwkK0wP8NY4OmVjcR/OvnXqUVy
i4c6nh/eqnEWFKWb4VUWdsp65CG1wJDtFPb9SUx0bOtlmp1s3zGj1IlE3cZ7MeJr7F6kMZmbzOtX
srep9WSn1EvB+jhKU8YIrzje/93yEpNTbpcI6UCuHZZVJ27hn89ODg6GIErFpyrjt2Gn3aSZRf3D
7Br7ZX4XpfgaJbc8EBDxYYosjZsUcN4jG9pG55V+1TBFd+wnQe9ltWnNc8Xzs++LGQ75oOBlzhd6
Ele2pJxIzxvrRs0aSQK4TlcB66nxmktvyP6AqyxmzcN+TWXEEtSvAxYYaZuwcoKHEbwLNk/2X8NB
Rei8+8bEmGhNes9JAzSBcJp2ZnniardwgKUL3AJWtvY12d1gZBS9w2u77/PvC0Pwwc6sfB9a4/An
0U6HoQoHBjftUfsgnmBslPQikVetLmspxphL/CUW4/7HXonEvWRr4hJh/gFzJa0qVpv7PWnkXTHS
f5SP8z2jrHGTq8a9Cr2BuJ7keEm+4Kdw1j52noGpGTOyAFc7jERguaiOmDTTLdaBu14mx/P/WbCN
WryFSU19KrNrzK2J6Yzx5YHLxbUMfqj3XgDye6V88MNKasEBdsZkAgEd0OyDKQhKctsCsrPgMLs9
6GL9TyZ2rRTmoOCWgZQ3W56cS3/oAyHbjeaQkDMM3CBVQzJkB/kpgEsGK0ggOcBmdsS8LZoP+oco
Ji3mSBS9Hach//eK5ipBdrkSQi9PeSdYeyYVP2GNIqZqelRrrP6PDX5cW4WRGhs5A5VycmViD2G3
WWPt3oZJNBe0Vtfi4bb/xkYEHyY3JFCqn6BpsA8rXdheiW1L2BOQ38fX3lFzFJpcy/LAahehu18n
KkN05/7IppWM76d1xLG5bwMqR5XNIkOL8p3W8cXDmkct4TGvikTSjP1N9I434aUdajqkkZQvzMyn
myW1KneHKalpR8AcahA7MSKtWcGGe7WIeGMKqdEyXgl+knOFPsXkx+owIeCPGmzqNNjytegBu/ay
4Io02pRiSUN5kyD1LDnT17Q8RjTS5lsTJW3rgcTMHzh0KRB4kntk8TqNbzWaC3RUVqGq70p9QdWq
vAe8cRh3rqH+0MiyMhvu3UwF2sN+TXLp60qdRqD9jxqy8zUxQ5V7hVSPgDJdYjyuAq7Lo7GV07NZ
WCk5BuBBZJXvDNdtQa2Ve7B+WgIlR9QUs4Lhteyc8HYvwywlD3lL/vF4r/BU+ao270jadXXbRK8M
5qciR5Z8Hh78lzlOTVtfvaiZDjKPjdvECuNrC/mv7nhymPSx7BOIevH/aYEL6J4YAl4rV3ADCNlT
GlYa4Bitu3iIHa94zZ41fp1Yrks9xYMKAPlyssQ1JA1gd+oKABMjX95GeFizs9v0X9JRUuElAWlI
5q/0HfA7ZelEdObVHl6XHZvgsUuLd1oOISVNeR5SwU0EJks7Y2YLL+2DSSHC3sL2KbpNxzv3Ph1c
pp8MeuKiGVe4gZIlv38b9JE/kw63YAg+LS0CpewT+DxGIjkFdfxPjgXEp/bkqLcDgScPPo0VI1CJ
1VB+S/WUHImTrg7uCo/hbHMwLZbdFctwPWWyhfocl3m73cbxS3ilgXW1qGFALFNkGffj1J+kS4f0
IEuTy4p6NpnYCgI1IEL4SHMdSlQCHuXWduaOsP6Q3LPmif91dEOMLgOcH2bkIoMrcK3Dc3ulZVrP
wtDAeGkCLkXRo+u4SNIA+nbVzdZkIx3W2iLKkYT+V7eYOPZ/NTW5gxGfFgBy0nx2sL7bDNjuvhfo
QgHZypw8hSbxqqlczD+mV0tPIzVLxCX9KQwKUPkGa1PN0f9+uLEsSYuEpNeRazSVebMFabYOquTC
MVQoAAiD+jdj8wgTUJrm42UqvSrUz390+IbRET6d6H3JKu0S89cDME7is5NdU4VCDkw+9eqTgcOA
1/vMqruPlq2kVFfyfLVwS9TA6qg84640l+syQQXUNGPpDNK6sBCoDK7caT7Jd6oRip6CedJuhA3T
mr9EgBqXHZet9I+5D9iUmTC19YnTOKmbS8ctY9L+u4+OR3p4AQV5npKOS9ZQo+Cgm9tVq/ZZD5Qg
Z/1WkB6bPjlJ2RuuEDAp0wxNhcFp3J0xFOIROmdcwDNYBIuNImi2IfrOZM0fqMLG/5JYAR/lkPHz
hRiVPS9pYpk0PXE0LOF4YRZhpMCUyU3wAE9xqp+ab0HW/hjNPBjLyz+ZEU1F8tFMcp+bZgeMsLWF
1zSZVb652oIH5fxnE8K834d5EIQBR+fv7W6XmZj+8UQ0ew3+XXqWsdUqF46sTualUh0HmDk1caMP
CxDgxnbcEh2hWjKw4QiKMRKdLn5sI/Q+Nx+SSIkv6IrgxYAKzdmtX2MkbrZVAGPEZCjDykIknmr5
VhU5ginRxK4yH4FxC8E7hD6/7wZbGZYdrOw4brGUOI27iPNfPFJtFDpFoFg5sIAj3tWLEphcRmcL
RZdP3N6h3RkiP2croLlZiKORdKWYjLwofWDBZrUizRAQVFhiaMiTVjHR2o+vVZs8LevlsH+/VgcI
gRMyPn0j/P5r/cDOZphWlq5NGLCi9pmaxpVfaIFI8tegskBujNZhnfXiOijQMpIhtC0OP3hFF41J
PwTrnV08s8mElprAkYWEKuaMxBgrMAP3mfr71amWb/o1+2OZmnkGuBH+bcKsALUzZDTpBnNLpkp7
Vl1gDAnFQYC5F9PmMIHXXo0m4r2UFYx7Te94pz5jNwLEIVahQmpIKyTaLtf33PHzppk3beCDDMff
PUpQwVtD35HLzwlUqJg0m4Pk65QCvnZZLNDh8ekj8dCK246Kj9sSNb0ztEZ8Fe2ymapwMDAxWnPs
JgA96AG31bA5hqXN3sEx18IvLtbrs3VD/ByxAI0QnglB81vcs1pFcsW4gM68RTQmseZ/mJAjwtIa
TQS6DuK+Iu5ncMtG8SEPnCNW5iLpdhArpdOEAkVPXSusNW6DfsJzcFlp3xZy5QVLscpG2pYz7qHs
sGHz/nz8l8ZmeHapUwjGCDgH/VMDPZQPj2QJlU1kIyaEfB+fVr26z/hKGrs+CH1tF69Jjcb8h8lv
KGyMNzd8pc+/PWqqrKNSXAE1zc0N5x6C30O4Q1vbM3ttCZtwejp6RUNTszZ2NyZuGKkQgA0CCu+W
HbKh3fU5cNWv7edDH9rJUqBGV4jinNSwf1N6sTj/Ce/tYev5QH3NY7NfrfHNBlrGeYkjqQx6znkY
W4rD1q0AjwBHcf2Nilj0Tl3AdY2AnILePZaOMo8a2Cx9C7P/gDBOQ2DFqIvH6rEyoWIXNZVF4wYk
cVQsH4L8a36dXgaIrJ4y1UplCsxP2m7UibJhcqI2Q1QPHbfA/bJ2c9VbTzdZnz4nwAgWR61MX78g
YwJ83RGrNSnNYyno3hYNee1ApI6gUJHw8tqkfXcgc88lYetGIM/l+jgJFUjWBO23HMTo1OMo+WkN
6ZsCEyX5GrvTU3TdhMjF7vdVLmAj++y+Xpr/VX3fFoWLCz1xgYtQeR1GSQdub+LvodHbRF/P+MsM
FG7yMETZyjOb8DVu+A7ttZWr+4Z7r/TUHgO/XM1q+aArFil7zwOzikSWO6Dxakm3hekLkfVojZ4/
/EbZbk9Zarz1IXsSw9tZtz1+pFwf5gDNSXAgnEz40Ymx7epwiNlHx4HVH0q0tuXkEaVOQfrsy+xX
pVX+fmEMY3/0YT8haoVjOratvLzFbzKzIXZpIuVWKbz8GWKqO/FLHmHaeuurzTNIfh8LvzoV95SX
/FxdcF0R/0c8wVzC0fkEBWYPJ0eaFSI7ZDCcE+de2KAY0r9M9l0p//IFgqSHYWKfM8GNQeO+i+Hw
x0saj4iA3L7XHHUzqMaq7nRHiD0h0eazDRsFduCpozKxXbUkKJk4mUUUO5lLohOlWDPU97AZRvY2
JxP2h5xyNBwfJArAOIWrMco6iNR6s6F5oWqUZQU8WESN7aSyp/sWG5bPfcYsQ6FxJxTeLkaIVdfi
Y3Q4THGJ+af5TnYZiBEkBqvF9xhSJzE/L1K9zdF9pCQPoJqHyMfd0ZimaUZpd1ODF8/9SHxFq9o8
uv9N0RXkB2L/SVYNDFE4JVjlrZUwmM/ZaoedR0hJsthlBvMD77GEjc3nlzDIq/k6fHO64YzoeMpA
bNIWQwDrpx/C57VtZBRqDcmHsmxW49RFipoVgvWf5W0fj8WFdVl2MpAA3tyL7/mkC161JbmJ06Lq
5bTGIiamgjOA/HrAb+eSgPFkYQRyXcklm/5BSTskIk69ezjuTRE5Xra9Q3Z44BqX8jpPhbXYJ8U3
itXnO4FlQRx7mk0PPkT1YqDiteebd8SEIwdakuJf53WXxf7U5kW72e/Tx352EQcRsLWlcqKtnLTQ
GOIwXJ7NWaeNEAkaga0k2TcHY4Y0F/tazHJ1NU43Ig6E+DlqzUrAnlgarbRDOTRk8ldITAVbVKQ7
TVzOR0SH78L9VM0FfiUXg85RVatlIksDVCP6DuYWD0NZtYfXFcmqaGeMtKw9xaEKGlrNDHkvsA+f
yWaH11+ioiFj2tUzDaGXj8yOxjWjxlti/9PFae1L7U4bEZofy/saeSn2VpRNfYRql/xPpEZKYy+Y
+1WmyNSv7KSxvS59QQqcaCiiU7MORa4BzliNBFMTVLH3Dbe5zIVvBDN4mw0qti/uudtkcEYWzgLv
G4tP6RNfDiY/DQQhE4j5oA4Azwp21lKCBcQDvagoNOOwsmi2z+35OaPgomlj9PbcSnTrp4X9xhwW
HsAdFYLBm0rcc7pmjsVWJgT9leJVxYjxTwEO/WbtU3znl/OlP1OxHL+n6vTisLrhTO2rlNfuZoRQ
n+DjglU7ANqhngpxPheJsh7yt6rE4H+p7ImEcN0ZaARQ+vgyNg3d8omMfAZaJb6mP9ewINWhHx+D
sFe1fEN6hdsgL6cT89g/Ay3IN9565uQTQAKgW2jdw9ElfVDtWUkqYXMb3pC8v3iA96Z/PqDZYSiD
GoSQds1abt493K0fPKc/ahc9JiUcfABkao37x0XoehUMwmPvlabbpvs0xe6gu/V+D2Cx7DxqKWq8
/UJXwJ2Wo6CSDVyEkVfJqIWa7vtt38m0bDrRZyd3Gy41ZKvFw3AXX4G+d+DDTplLhzwGr35AA1RL
lKem3XwBJMpaRFd3fReOnmvIbGaODadOiiGm8bsycFQBlZ05S6jK7RHUUI+q3xDzo+a1oaWx6cS8
Xs9YBdM6qXRlrn6VfeK8GSoBES67SvbkkRXZwSneAwbbzwuD+svKjJVO2Z5DuKn/RGD3ttnpD7/k
oN+Vqc3pgIdr3gmGVs07taVZTt+RnQIPi0IcBS9cT+e15PSr5OYFniliXDoxkIBd1q3aHW+v0CNF
+fz6Qp9SGq/aUEAewKrWlt4mvFg+YmyFD3m1wftiXBBKtAkSrVw+YJC5TEJVACTBTCwiMXuywnHJ
IaHp7eineypTv+y7PzK/PpB0+8In5Up38Hr8pynQ5QZXiPcEYgz9Kvzk2Si878rYtqCvTzCkZ1DC
J7CHc1zIUTGAbBbsfeLWlp+rGa5o+qjl+offDSVV/EopxLOwo4KCu+9LtOBJwPTCwV5iz79KGzpr
9CTEUhQ25nllKRKWvINgh5UZvQpq6CsX6SJjADEhmU/KZFPb7cCIJlH71FZ6lUE8+gUIIeIzWuQH
nTNM3cYoP2A5rW85P7xnqoimipGbDwEVMZm7l7ZDbagEj7TqtXKahbCHRbFhYtY4UnDmjcI8hbg6
B9whYin6f+PnQ2SAVYmulxhjMbiaIVWfMHNIxiS68ST+ePI9gbL0cgNgSDqn9VyVWHBSMddqwoyB
RqXjnuTc1NyNxyM/jguG/tPJmWDIpRgFUNEDazbOd7UlqSprhLraB1AzE+enLCKYw1l8ZIsoT6rF
/bXUNjoKrxoBsdhUSIuX3jF8YRe6J5WqLKNnHDo39ltvpWraXvbZ/BQ9kXJcwTAri2XqTRbf8o7b
+v6SmFy62a27Cw7v7XEBY5Mt1qfQsBYI1oRTCkr3RZ63JY73T13C3JU977vxiOO96gYTd0XrpVrD
Juc6pPebc1Cf5ToTHyoKkC1+LwyuuQnTt6S/KnTKU9OPxTTwDL8m0JS2k7pxt4qshTRt1lbHE4KH
Li9vK1IXA/KWTGVhHZPvNYubgCalsDYJxxrgwCsXV5B9hPKrr2ReBt77PXR2lqRuH+TJCdF4rPHm
wmJABJXIcMCMtl7DaJSNNXAxYHvmYHnxZUjb5sBfqWuIMMK70jIOIPlgsIdFXE1AhLxytY3hCxUm
1SrwanlgXVgPuvAP2i0ZHBbqIQsqH50kad6juVPF//jR+8GjTxI1Pl9nT6SmYPPjsN+jnbm7q25u
ULrnHa8Uisw8F/G8IF+AGT7svccq/tznOP23igdCNelv4EGDaPWhn0u3wnJcDZ9+kXQSeVil4Xkh
KZl7Pwi/4el+zeLKd8i0mHh2/JMNC9y5qxJtGIViDu0l5e2p2utwNVWVLX1STMt0IX3fA9GWUvbg
aO+ieDptpTaTNZ0kJbZJ8OPdwiPhkTRNY/OxE9fv9haqyvjvQv3bZnz5VOeeuJmK6BvuK5AVgWqU
TVRIhDYaLbNyulx4Gth9WFqVg/tT1WktGWwU1f+SrwG2xlF3RPJ3vI2WkV4jJ3Pu++OHtrDM0q8h
Q13suCfqk15XznaEuITkcBqSLt7zi5fgNW48EnYCumXnJ1vXpwS0MSf0q6w4cOD2vpXddX+OvHW4
iUP0LLja+mW5g8vFRoOw2lb+WDhe3mfoGnpdsBuSEGFpuWK6tRF0oKBnoC9SgPi4W5D4D52cNsIV
VSbTpIQuK8qIRUYjI11XEpy24e/DHU/5ir2LenPSbhriZJxsvytXO17SR6fbSQsK1HFkUTOs3ZPK
iEhflnvfnZ/Ds+YgdkHH5SNX9L1pZz/vKPJQ/IwCi9bz6CDb9qfJgCm5ahSNkr3YZieU1h3IHBWn
+J7rmEIr981L0XG+tCVym2Af3IJxLp9K7ijoNHfYgPO2sDTDVAf4DCe3NE0+AuQwtvwMtPfvFRjF
iggenZ2aVSmuBCpyCLB2p9aaAZYcPZXDDtp/kwW4d2ON5jJvFgX6KbyhdYhR7Bx6bCJu9xZLqRId
1BsKN3NYhJRPiaO+mikaKbREveM+/QvF6kDdVMde0GHTr0p0SyR3GtRvLh6Lb/Jo630ZimOz1Opx
bW9SioSh21pNyDpv1T6yK57TXE5pgf65y0D8s1Rsk6MSGQV8OMa1IMYgxB0bWJCH+ajTxrX2kZug
v9oWINaRfV3RwHvrrOS37KWIOuxjqO5GnduPM5m+f8kC9eH6rGEbc8h0PMJ2nNvhYd0m8vBaRxlG
60tE9XxL8n4zUBUPkfsbkSeJCZ1+B3J2ufT86snogNYRFiaYzNLhOV4LZ0VRv3KlmfDxmtz/oc8Q
IWNTLKT+lml+AagQB2HBIHfMSd8v9SnW1AUaS6gKV5tFbTH4AzAj9yTyUdtafjNqai9mmsJ9Xugg
3axVBLlBwf/BwppN6WxZKGEswwk+S0xUm81LiVloKDXhuYD1LDV6y06974qM+HSyTkGA1qtTJHAq
Ag8bPI3hKyfZNfwiB+/qIKLHN5JiRDw2OXWf/8r5oSGIuuWQtluHoOVPuw2Vwwo7eMk9yXiERPnK
FJVYcix7b5hhCc7bze/qVMbftJODqF8UH0pl1K5g9Aomf7GcWbxzlg5WHGIrQDUwze4daLGDX+kh
ptUnSfVBWij11m0KTwx8UK1uiXEReQZ2OhlngfzOz3OAIcd/RPsfswtg6zFvhPAbXIJQqg5gnF3B
Pd0b4MAUGsgX7sAbBnRifLmZmHHbBdcuew5EYnJ9DiptGa6KsfaSB/GAE7pS98/NQ7M0PfvyHoaa
DJaLQvD2LpA9MGviNQZFOse5O/88qNOceVrLqeWlawHvxoGa/hTcybisupuTOERILA4FGKMKMuzq
RFsjULVy9fcwX9gFvUVOLYu+ujO87uylqQzHUHn0lYVkJfE53SiYPJ0UGe/0TfpUoRE4ZE8SmvsJ
G+xiQ3INjSxFrIxQgZS247x1ARyNxW8rlNI6AxYpwfuP01EpDeP1nlbMCuP9G4eNCraD6VSOrjBZ
QVH4aH5SAHGLPfj/91jV0Adv3pwWbnmREGqGF5P3BHWumxDH8KTUVZApJaeNvHjfbidECw1frLvr
jxcbMyX6Vqv3Zsvlmfso5IBCteLGAjxh6kttW8tDFzAPK/byvS66sBvDypTzAZOk/Nc0N+KELcir
i4nmhMnhAjKJIOY8zaNglZnKtjJxvH2udkBBtv5sU3v9BVqUzdey6s1Oy8jHAqpmFmDdyeRu+snG
QR7rPTwW3nWHbIv0ChBbxzuiqqAcGV9v01g/F7mquFWJ3Yc5IiIb5Pg3CEEGE1bEjaUPhJewNKrP
JP8kCq+jvnFv+3SUEI2D0eoizLFV6JzAFUaK7Dbu+AVm0lZZ4WX3QwRR86fYhFckvE07TX2y52rh
gQEILFEcoM5LH+emk6IyV5bd+rluMTX/2B5rn86J1AQs2bHXHtcuRS7oNP14WqnV6JSU0OVyG+uG
/ZJgePhNcbc60ALG4HY6Fvrjj5dv2GnVE81ptZavn792Ldv41JC3Zbgp+B02lRFvb77zV0sO+Uaq
3zG9Lgc6c4M0rENwvm0eU3bzjuPyuJ9NLu7VPYA1wOpcygOSAk1vDaL0Q9a4JtNKJsfX0XWUqd69
8/VrvFWJ3Nxmqt5LseEYpm2HoMPKWevp14ZEJo1nJqH0mZvYCTnFUXJBFpfyo83PFAwMgqTbZDb+
L+cFs4124hNn3BhJ7PvzT+BnjWbWJSjMxi3Sk6Pzh4SsLTyvjrUjT9gRJCpQg6fk3ynnhbA4oaoS
SxdFGjgJwTASyy1Ih5MQwoyNXzxWNeLRYV0a4R+duVOz0ui3AY1U3s83hxwb/Mue+XihOmJtt0Nq
9nWOOX9jMh2m2Lg4KhuOMW3NayRV7w7JOi3pvWPHK9w+Dp0uv7ILk8wQo51qWU9uK2oTIb8t0avU
dysQ7I7lQ+PqdMhUFyXvQwLDPDWxGL88AZxjc4Hj89FboDJEUG7UtB1GKMg6fI/O7Fz/QNMdKj0T
aRWcIVoN/H0IRLvUvs2nDpcadJKw/ctIKm+gPtpMamxsQ70PSd8BOCuTujDwCO/qoM5w0ztGDqqS
3zkf1iWguSyBu7szodPVcJHnHUUycGRPdktKROBjLgqxquMQgjMAiNx3tuzLn47F6V4BjmqwEq7w
oOWSkfbd5sOYmDGPTXILyEuHb4atCDZ5t+9AU78UU1/V+/xdEUcYBlmyjdBjNEHLiyI9XB+OqmRv
15MALe2dUqBH3DsAgBDOCJlV0NhrVGKngJpFykMS+9eXJGN7fn6yz5OSHF6sS9xrh+8SkjX7p6ft
J1JJv2JjQWyE+sjr/HnJ5COjsNcSZ10ipdaivq6LfUmT9fz6vinsP4k16d8YWx15WWdFcWEbh81I
PZLjNL69KYvPZX9gZDiB2ZsthueslowtMb59kSwxOr/jbw5UH6CnRxFlA3CLel7otipkmHdkmXXq
lzYvFQyKoj0pT61gQqj13t0QRqwBNbgnTq+MV7Unid6iezYstG7114A8/17MCpYSsWDhUuTBWCae
vRNvw6UE+x3gPACyNMqEwEMBBhgz6g9HvqWEc1YRRwfNMRYDOFaiWKOP+TFJMtvpK3FfIyYLUd26
0o/BeDqWRQMdpn2jp1iqAba1YO/se76XLs3QRyqy/uvvUyVM9Y9qp0YwTFH5dylZaoLy3Pvo4vU6
xw6PY20jVuqbbhuF4JCv2cN7T/N0ipMQ++yVP/dqcMhX6ED4Qw4M8jgM29akuB61na5xbD7jRmZG
vREnT0ZLFa/HDO3BX4fdIk60bwBUrHjr8S+0jK2E//QnPU00aMbJuZ3J5jCOvFRhwAiK6mEt02c9
qjZpJywEue3uac0zbbKVbzpF6wJ7lrwXa9L7I4X3KAzKJo32XSeijYVT4lfmwP4FlQ2QDopEqRGo
QwWYMgqRbUP4lCzdxmvpHvJf1zjcO9F1ERpKQud+0Gxf58JDpc8aW1zJy0bg0iW4MBDlaQBkpteF
o0qQlU2FJFmGVZZA5qAHzgte1lTWFr1aCn54xJclJggY08tTG5QDZuWn49K+CEw61JMc01tm4WWx
gRXobh23ow/ySwboTCbC/JlsiM32kE2NY3xXmafirRoq3X5aMreFjfMSMcR6il1KGjhIRD392yID
kz8IZuPa01ek61Pm2A/qsNzEwjr1Rjw/pSBnTMP8zW6uVnOOlvB5w045Geeu3wR3+RzUe6SZr8hs
bAcQNk3nGmlaMqkvnj2v3yeIoEkGCws8p7yRLNOBFla49Q+G3RbB35E5VU1ymJcR/PcAfdw+UQJf
aaAOn+5M80M2rWXaNY4DC2wloA4G64fSvQ5shMKkSbR4GhnL2q9vyXJXv4iOs4WB4jalljAwljUB
Hjz3cQ4o5djx2OzrxmK1X/Ae3zAM28Ig7/yLMYCmPHqTFDt+nOrPQ2WDDrWVjc5BFMiMFKppFpBM
KV4NCXLoLi8Jcaq30EHT3vjBgBXvsQn8JScY9sbkek3Dk18TTf5pnKjABvZ6vRm3FFpkitMir+Wf
eJAMO92KzPHQSKMRwnXr8MkKsQH10gL02SD6C0BiJ8jDj3+s+LQEIVJwUrpNMK6LCi/XZru4TfPh
DAaKUrpuNiCvHHVoIWCKU4PgUuAi7vaCmESeRQL+cjRLpjqPF0NfHpwXscFeKjd6x3ozt1JVaFCI
2I9PFuO5lYYmMkyM1m2rv5ULsv5CebkhnTHm59AmX/7nd9erPeYvSNkp0o0XjfTsJ4RfJ4j3aQ01
IpbVnhD4cpiA48hMlNL1k+ThUk+epSEVu+juzjbDYHRyOcpmLa8P876k1OZAN+GXsaMmZ3w3KGZI
P3lJbJeJVsnKcZ6tBhSm8jZv7Xz/A21zw+dWn+U1TyGvjbjeBfQxi5snCYAyHWYOKXtYmUopkiLI
HXHeS8YmeKSYZMoxwA3JvNl0seq9iCxQEvBN5ZKAW1zTW9dVrfVemtN3pRwnILBahQU4bhca/ncf
dbQOox0NuneR6+N7cYo3zC+57V8V65naXkpeZCTAUD/Pg9PIJOT0vdy3wZOl7Y5Y01nJVJpaWo8i
h5qS2Z/J528X9X4fP+AFr9bae83m+kTrvTPT0tP/GviMp6GNUY+9S9lqXmOJEXA8j0FNRbGMncoz
VTkmKcfR29R6yXQ4gloxZ8vc/iWx5g3etQIT4Z4Tq3q6TXl4a09akvoYmiqXko6syq3uFTCGfMrj
8/TGNr6fVB/HmIaxCso+NtT1SqdGNnH/I0H9t/Cdo+32RIVGImmuapA7cpCqRed1afF3GEInELMM
8Ql5bVc0zuDTCOkcky5RSdGoBv/zBvCLNCtBNbXlkA3gFNLbt2GJbl3/xfoFG9nWRq7Ywk1jULxB
1rFkr+zrUljito6AAmstWEeRa/wAhj73xDLdiWwepNK96vQKSqqiXAg/8zJj2auCLsCFptSOqyWV
NXjbl/zaamRDN0lG0pC66ALHBNaoKII8WEoTHn+PBh/j64qO2V6KUIWtYuDHcO/IGdi8NIFdFTJ3
8OFHhOh5UXVtGSAi9d2oin8uJPPghbO0xghEVWazucO35LDUiAj1IzA4LcLl71VmRsoSm0c/28sJ
Na5xOrcxmlTufSYVQHh9EOFUKbUKe+X1zJVPm0xGWVgzyQihcyLNLV1qxY0UjGAxdGbkhozRLNXg
4Ug8ASjzAXKWJcstOjKqcF6+rVkBIrnkqUop9GvPqrEmrAcVMp9iYi2h3eMAP9v1sEzrKbfocbFQ
E5nV9HkhYhfl/oKDPm+EcC2NF6sY8zSbtps1sF1ZDUgiYQHmmrDR4wAo5DYBu/kIo9B80NXjI0SS
yWUhDYsGVhhXiLi3apGpXUOUAxp8pXGfzN8geyGmwCXU6bV8xno+lfj8ylM0wTJjgxjMQh/7LrXP
R2dZLLxU3LoHrLupFdicZczeRf5pLQj0GJMJq/wYtpe66g+3h1SR7cxWlAVp+qKifFqEi+0q+FPP
LW23z/SYDYXREjgsiNKZ4gkrwc9/AGdKtwxmZn7O4fzt/5AuBEFtWnJhi2ifgRdaLF88MTV+XhyT
dvcCThMFckZVCqpjnETuddbJHcZbHLVlLHJYTvRmo/0BwsONJkxEfRRVfGQSCZqNvQiENvQ2rCXm
KqEzLKdLigaTpE4eYsUlsFzRJznU6VNXDc8p9yuc+p75phc9m7E03kT5FDdCncYo4PR1jfbN5mEH
vb+9RpYSLMLLiF8+KktY765fzZieX9CeuxdPw+O/4/U6qKB2QW3yTcABVpq04hYJN8ODTkscJctI
LH4QY6nnGkSm8Bwg3GsZAzqmGzczXRhQcKQc55fjf3OceOt5qzNanCVN+IKgmjoRkwA4mKiTxZIA
Ebv8tAPo9YwOq4ArNDYWkLQsfNKlaVcs8eDdcKSFkBWEMFOEpOWFPrPXDT/MqPz2rI/mYSfQ6h3u
VSCvU2fUfU3uL6eWwLYMiaWflo+dxEuxKRLvpTWu20S1GR4UVwsAQpX4kkJvVtFXJ2f/0nd0HO8E
tuUajAhqGtmbweU1nm2goiYFmhA13IhDjzsgrYRjluUOzpHwVX9SyPrPNduaMyHcaWZ8xyrPv8lG
EejKf37HRZm0rJJH9smSsA9yRe1Q6DP6yedkoeAQyy5FwUuZwH1+fTqbEDQNUVD2DxfFrNw01Tuu
st6hSM8n4DJaA7jbd2uPXR/kwx8p8UdBOzU0ywNqbkIdwJu1b8PvfDR4sfk/WIj1hjRT8KzLPwe+
4R1Xv2juiq772/mk8dxxQOIEhK7eT+GYn6l0eoF4ZEl9BMrO9440+1x/9u5DW9TmS4bDzRBfeaH7
tbm8dTbj/7mxdHzfBY/rnibpsEyt89PlTC7UKpZA19PU1UByMVzTPbuRF4A8xAJ15WA1oX4p3TVj
VtiewSpMaUfPbaURs5YP26gJT/0A53H8nsCxxuXRb4LUqdwN3qbQw6xLSAGwjMGSnuHDDc40tSqX
Wn5M5XkrwasJxLpVxzi8xN7jcz+g/eyRC1Gv/TFXuqjdt/c22hEWhHGuGfrjGRLrhKBL+BCtSpQ0
gWChRKwHdUfiVou2JFJ657RJR2/PNubM7VIeG2paIIp9JyKO01OWHHqvMe328WKaVsMvlY4Vtj14
C7HaRlyMzz6kH3Io0c3VvXhNygGqAqIFltCe6T+hHtWG8GahY49tlluzEOJ9578aLnuqFQhd0xMx
KMF1wqxIr0XQAO312RLrPR82BPY9Tc808c4iuyWgH0WWZ6STnds1YeNRH02RoNdnC3sAWtPJApym
wfbb+p/HHTq2yXXhE49KAqlY9xEMsXGHwJAC0MVo1vvd5eX+XgRpuesAs1AgX/Whd4w3pFBt8wSQ
CSXP5zFzDO9JPl8hRWEp5/xeGjyzTAQ8CcPVEOnJ/FlaBfFLn0APwOU+/ZpxqR/DSDGBkjIvdZ9F
UzUAN22FBoFiuwKSdxrwteBek6EL727F5txI0+Oc676fsfJ3QhbEfWkJwdO5Z0fPafsTwrgTheS4
X+IdHd9GFb3Xkbk6iVIGj5OUifmmYcSCeZ7r43GXdmf1S4z94VLoeOBcSAsdID663K08ZcSdbKxH
haazWD7pbJCpUojY7ljO/GHEb0RryN4ipoX3HsA8m+V5j++ywg6hfzgppEevP7TZg/gcw8+ZqzV/
+8dUd4w4fSU6/C+nzbPR385N0063Iujoh4NBPmUqO6nBpzCGaLvgaZYK3gijRrq+Q8fV5OsxgQzI
NvkBt5l3SsbBkN5S+E7XzdeOTAOK8e3PYvdAyQ85/FMs4AxZ7Wfsr+xz7zmpjiRkDRTYrGPT0agv
lCFKHg3XzPlpak2+kWJdsSxSVWMPjq7RrAi6400MevCETjEvpyvHpLcTZo2PJONMzyBHL9Dh3ysz
qs/7UVEhvVQRSPINIVGcAl87RPcDd2EArc03S4IYCfYYzI2gOTatf5L9qAk2OjojdiW69jX+FCaw
RRpAuDzHaOebA891l/eDA59ZN9pUNM/zcms4e8wKQJyGfRToGSJa9tkrEAuG2fNU2XC16g+Jr0B8
iuxy8XiW4cyGL66iQBFdaidvL3PkBrAYRNXQEjywlNV5KhOOxcnApvz/9XZmYfZz8UqmqhWZcGED
No10RT0vz55nk6DLhkiygX93YEpVeIcJGCm6Y/LMCmMgFDsQ+UKOR75gYp4Oc0iIAHFDIqmRGh5d
Kq6PViOQN+gB1rCEFgekVgICLTD2mdn+3b48bgjjZcwjpxnSZlJwW1Gajz61eDI6AlRVzfI5ggus
5YkiCg2h92wZAwreBJRuxm1vekpnBjzynkE5W3e+hBb9l+Ei9qjftDTWuRu+bj1eoS60DUkeFoEp
oYP5Yxhx0UcViBOT6Ow5vFmIg3oSCBHJYao/rMkxdJhjc7rkcwmd62LKRMuDRx7pJWkq02ZR4S66
Q34hp0g+RiTWZu7F7LSC5rHpbhRGXO2VWTwbHkb0M5wDRdMVudQ81Eur7Sy379jmiWxVuJbAy7S+
058HAv2119xV5ym5hpUfBuwlKkO1bd+BtIrZdO7fh0yhFGmrTRq2t1J9i5/7cHxuczMOQNoMFSVQ
3oYlK9XHvYYWDEml+zhzj5Fdu8QZmgtVAqmbAQuraBWJ4X1bZo9ELBTRQcMrlaLRc6+fVry5QBZl
+PH/j06FQP0GWuK7EMp/lP4mvdYMXTTIc/+TblQGRemEzjcSzbk+BO6+dYv+oCrPsA6yDHNUNlOZ
p5/D6RqF4gnq4FK5UzMdHNL23/ALTyeltLWBFU8Mx8KhQ5F5Ky79SCw2Yg+WJ3SrQeDRhO7ATcBl
b2to3X3lb/ICLanjCYRi1SiIwVJ3CzRG5CeXtGm+KfBsmne9IsidvrwAdzX2aoy/abibmbQtJoJN
//8xbMK0i5Jzo9ZuTdhtNiIEsj4Q3wKVBDFTBsv09N0L+UClL3w1EXZpw81bt7fJwX/+7J+RsVsm
r/InsbtwrVji/BRL7xw2H4apaXhrnIfIa3ZP64Y5l2dPJCj9zfvC0ilYLnMf8LcCVwXqKJqatfbe
5efhbrCgoq7OAZwKnMdhsdPfAATZXWrwnwkMyi8cm9lK3nRlDnl5Y/PimSsJdWwI0Q3KR5jBKo5a
hra+pg/J9wHW6wHiCTkw/GVALMqkjdhtJlduweQJQGUL83BI1e7fNIRhOxyMQVj8zTwxmv33Gedg
69gyJoul8XTSRPO+sFeIcxzB2O3sO9eVrNtyzsSGCQe01Xv4obUwxEer3F5iw/7ahKdUXSy+f0gt
2pdMDmkXm7vJs8jF5WOFBsE6TdGO79axz5nsuVcxjUSsQv7oPMAXUufLWYPOmSp2Ckq6kHEWS706
AzotgfWfPwFmRbT8UA6ido4736Ot99nyBQtoMut6oUxX94soDpcoBpfWgn4Ie4+iOUmy0Ej73p0f
eWYrwczDAqRLX7/w0Fk7u4yBUzbM2WlkUvD/05MN9aKikRz4W67fXbX9AtN0Zc/G3SJ3sGlw1QTu
LwHZimeOJvSFKTiJRzU6zL9WwZBHqUruw5CGlutjTzuasTcSOU2DYm6LG7Qbd05jeRAAZ1V5yNp5
I9KJl1+vrpBdLoKZgIskqM78XrKe5eiOpIZnUarn2qvwCZKPLRkxxq3sDT8S2pydIuVwncyf/6/C
lCfB5bJdxOX5Q+a5jAWAknopqAcec8AesNwRRT69P2howhY2B61OhtCLiBPtLId2bGdJ9pnPVt42
39XqA92aqDL8+3uXj3PhZt2qXakFdD8umqzu2M+IDHJtToFxI4RdO93+Gv1l3wraN+3OtREfSG1Y
1rpYpoaPa1+t2xMR0bRSrm3WTTigQrnBM5MX8l8VAiDBMRNkacy7vRi65h9oVAdJ8UP4LS0Rnw8t
R48bul2nvP4zZWpJzWQxt1Uad3oRdIshPstMLMthqXoap6caQWFy6nIR/sJzCr4UbVYU6MYwJ6JZ
6fdaoTU/d36aXjdI9O52eHYr1yGEVq2rrcXy+FnE0tEFAZI8aLolCvHO/G/PNX2DeLm7MksjDDsn
F5ItvR680EQOKeSQcitoP5RDhUwG4uhCKSrPdoGvP8aNbgUik5GAcxY7jpN7uShw0IFl3UqL5Z6d
NsNLzC79FTdE0W025MlJG5SRosusbgfq8HmLSl+gP94Iea2wZKtmRoSQQt2td9aP71khNF8Wa117
By37HuaT/1fmGLjlzBfcveGDjKl6Hlo5qcYTqiSKbpRk1EpHw+KR2M/yzoQn59GGOh44tfbg8Sk+
7O6eFUqDOx31SKURyKj9pj0e2MMNSytQh33y8fi4/PNhwLSazmQrQkuIyIAZcrdzzL4XUYKOuSD+
RUFu2BNn1xDgnQFre4jYFeUvdZfvs1dXiFYgJdy6uGvZPVwrXythRHdF3spD24LZWJ4Jp3kzs6m3
NDYvOnp3bSAYADhULo3IdT+YexiuseqHUyxLBNuw6JQeW6ky3Kuy1MFYG1kDNrxDcyQl+2+vymeO
12Xptz0o4UKRix1w5AnxLrPP4p8beO6O2HKNUXcEXusaHsrSoCGYV6ibS+qNEZ7Q3GJpLWyGmJ3b
JxPgEUuQPKIkkA+Q+B6nWuVb1AkXw26nD4chbZZyVQbr4ZGYCsGGkuMTWOZGPSpC5VleBmaE5XX7
7Td0sADIXSrYFXr6wQA3crfDIKZ28hr6JbR3j9GvITp4Ld9ym97cNrrIv7kPC3D9PsJqorhXpIr1
ltp9ATWxue/vMsZvyr6YyDkh40uHVOn1ZDTi4MzavzvAs5rFiK6bISYODv+lVIHYRLU9d+766U4W
YgD2ThPT9mkISPGjuL683Wp4Mf6oWPV7nytBHglWU2m8ZaXhez9JShBm+45tRLSSOBWOObQtYih7
jAA+++Mssc9cj8Fygt45cCCMnJcillZXlwsN+1Vwry+ZotFIBchtU4hHxVNpItosyBqpHc4ocNNK
cfykgJ0hfMbG561CKJhDCMt4sQKa67LYk2lXKhud0OHU/FWcQkrRBlp7K21ptn8+nUIuARaXssig
y20Ov9fTRGwIz7PSJtmBA01Vtx9YiiiWh1lT2XbR2HqwSa8vRjgwunHVIpFVkFnwrzslTAZLk8bL
gJAbI3kfCeePgASnp9iIV6s11mzYlIyMw/Zsq5Y5/gJNTiXDUq2bNd8EWH/mGwblCkBcepeBR0DD
utYNB+Jmt2esRGZYOJRA0szA6b4uMi0jxSmP3eUDnSiewHEbMapf/MXZkwwgn4HfA2czlfMyNOT/
6+g3g/EGUfMDk8FygGdAkFR9ah7jSVDo5hQDwIOIdRTCc1R4ujRA3sqWqUxsaM71t/UzeSVQ0COB
lVSurEgNMPslb5pY3UZ6RWQqft5phEpvtk6MNGymVOaydlNYb8jYeBOlZiifUhVGEz3MIFI2xHbF
K4QvwMe7A/ml5hR88cwYkDRznHco37Y/r8y2dJKyCHLkgBV3ZF9jozwop07dbaHArxH+T9LS/aXV
KGSbCat3AUlu43tAyp0I2xYnbkPLSBCRo6Jcxq4brpPTZUwyowws9/IqFxyHZ2IQ0NM7tUhgyjKv
LuWAegjvj8otSy1NYYXSmnJLeUKfnvqrmEcp4x6NsEZjQBIG7TrOuGnZUKHTfzrgCNRKKBy51acp
SkubkxZVxtoFb3JNCUObqB2mkVssYjypl5n3rXAadMZXTU95KWPqUVFYXuaRgtA7P6+iJ44oPAQw
wPjCGZ25YznvLT5FZ7Q+7SM+0Nd75B6QdTMgDif8ZyvVX1uAPvXhyD/A70Pd4FfeqkBFtYq2d9Mb
3HR43JZGZxrH5wrShfd4vgdvoYBMyux9Bu8agxRJtJ+HWl1/BfzKoiPC6enAmpU4gpZYTILsIXYu
IAdlP9iULorY2K0jvL8RYSXPhX+UEI978ERaVhx0c+HS0e8TT/KVpZC25gzoTxlY7Fn0ZJIn2yqB
+cHec0m9Bbxqxj7ry4+c3FjBj3ctXxKLgsd00V2OWdytXnzlBod1medPZv/ZGzLoQccSDqCtuwH7
875z/npLPNGF0c1f+pqPfYPwadsCfTUvcyHIAu+pbI+41AV94adMyudiMuJihJn1W1hHDXmxytu7
SGnD6dDJVN/tcJrVj+CwsnRaRDcHEuv8/764mzL+V11tUfqOxlUMTRU2kc+iMOiJeKQ2eSUx1xs4
7N3mqem9B6PrCXLdWEUUJSHooopMupdzoWfeEk4YTJwAbd4TJiqwdWZ7RzbDx48nH00rqNx03pMg
P/GHqBjkALDbTS+IvyU6YnikV+Skg3Fl+e1N5fAu/mtJiE5ydOCJM7CKZz5WLC0bM8MU1fUQdD50
UCxNxj2F3BaHkaRdmBogjPhjWfXCriO0R2u9bSklaemkognedNoyNsFAbSVju9c+uBYB5zaSauVp
vRocHIdxN0O87ZhlEeYsJJwOvHydZmZqsLDIZ6TicEx0k62rpTNJrv4IiIyVaMvnqjrEjbC/HzG+
4iIiPAQpNrHQy+0++6dzAW31Itdm3DI32G7fEtieNwPJch/h8i+eXUaXgZtqVWu2fIww4o4Q6wZt
QVb22XFpLmQ7Jctpjb8p95bzBwG2QzjSQ3WCSR0OC5q/9BfiSd4oc6zCIYeDd+eaRDSx3hp0qyPd
iDscBEog34suwkYX3EG76fjLvltTsmnvsH4bkNofTZHucfURdYJcZI60WodnkUlcXYOLPwn8wY/g
H+GVjL9rsD08OIWbKiZUR8fIGV+EIPyGH9pWL7H1BgDScr0U9iprr1ONVKeEv6c+Z1fRlqGZnAft
uyz47PYuttjunmOMjiJPVfM0gGZz8RTAv6g3rQpBA5kPD4NMN4+EdLiaNn1bInBsgjDcy6TXMM8N
iK05/Nq99NtgPp1lpi90HmMR+vvTxyGsfDTlh5wruTCoSO6t+56TZ5N2FQ4+Ul9MPRje1Q/dGjEO
YGlCikxQNFGms6kpOpl4i7CtcYTPcxvw67hzbc564fpMRLBX5CzBje0zY87WpZsfRa2JzQNAfBbF
jNbi2GUgh+gUXGJSxVFM6zLqzo/ZAXzZtQ5FJJFDvJMhGBmmzxkCufPBQb1CWVu1BXNLDccvJS8l
ltoM0v2nFe588pQyT+5nQN2mJeBVFxdG+DSfuQdG9TNxO8SYv6QuKkB7xL6FGGfddXM3/SkLL1qw
E4GwWIPgOsWilhJJvEM0aUF9nlYVoilqGf0LAPkXCYvPmwlCvG9XJHBJnvyZTArjiGBcsrD3S3s0
RiCXWrrhHLMo7xcnPPuMF7imUhhor2tnU6qn0SrKECo1NcV2ZepnAqMPVQadxKyCHCwra2VhhD4b
8Pn11OVtKaPD95tNTfAIABwMQr+LNGfQ9RAM0siw/50mo7NH5ZVenz0rVBXIxEaaWAjs5EcanhV9
efnO/tR65ipDdj0YCtaXh3QncKJYPniSjFU+atK4ydnDGTqnPzQHnuR34unqrLqkX1X0nfP6p6Tc
wMZUUPwNHHzAnGj4SSZRbvBdCSBzJB7mQYD6FeY+axeXV/HCkcw/NDTbpV+gqXvmTJO51OS/deZM
oFPw0LkEjWOv39EDusucHQphFm7jx2mhTSIZUf82fyNQ3JLrz7jeAmyl48P2Syo3GbIktF7o228e
azoSgaehN1xhyAa4jDnIbqoXuz0ygoCpYyYsCyfau7XYSUx+vUoqJjHfu/Aj4BmJ/3ye5EOwzV27
549oUTuYaNgqmNbBzZLl0HxdwXzhqNuInuYCGlG1NE0G77NejSCoXx1wmlMFhj0jG8DCeyjPZ/CE
70dXKZyq/5Xx16NaMLSTPUeoLL1rtEEmRdxgbDacXMvS2CrZUTlNyi5c3ND//8+8tYSkEh++O+dC
msh8Gj9cO+LwYwG+KMKCD60p5e7mA6UwAL+g5kKg9chXaosxUER0wOjB28q2LWPvvp3dC8Gs7Cfu
/zKbO3/k4MFkixs294iYYvVD0Aq0kHyaCOc1vi+au9quR1kIT63R4JHew8EJI7BjZRmdvL0/tbvx
h8lmRGbkPYcGY5nowSac+IW2iR8TzrNYPjeMCQvOWtgDFDCgmlONyfSXaLB6jmu6qUKsy16bF/4I
m7rqabzNvTElRcf/Vu6IHmN3tcLRn/vpGBcArqA9ZJJ2pn8Z8JDWXiavYdFUOzZeebzi0kbRIsTV
2UPhLTX+NjK8ehHrDDHbJW7epvunyQ+BtqBhNHGSrLh5ke4XKHu/wERHKM44/4r9pjxK26ItIkDK
2nhi27OxEpXROSfCghQ9WbXtPaw2ZStBfj5pQAOlRFGjzGeyNWKjzruYTES9dXP4Iqo7qMACjR3+
3wxsMct7wQ4HMAhbDEFn2MOPXxUaMw5wCNhk7y6XZHutgaV5jHsEks8alFs+zIGFntrf0RgpHZJe
PqtfhojTF9t3WFw8sjYk3/Ur9ye4eBkspwFEGoriXuSeGktAMBQSRyPfxCrC8s0CrhOKNnktPfq9
dWltNqQ3Hhoe+l2y8soqAfyO0nmJpI2tdd0+PQcMKeY2wnmiDm0ODnUO7Wq3uzBRpa4Naao6wd37
GWqjFmaIMnHelc5VaDlv+pHV51hLqPSoPANa1J/OxYK2YwvMUrevUQMNHIDlh0xE25eHZc3CFhj+
8t1Xwiokyf7VL9AKj4GBfLx357cfnBgCL009GBve1Y6sResxm5EJ7ijx86ZziSs9wMCCEeXyNaOw
I2Vj8HCGISbwoCXp+KSQ4zUpwqEtA6lmJfhTFtq+ME2r9voL+4Mq2nYadiRc79BIKmEILC75LLNZ
wtVOlqDQzaay5nYNBCdOfmckqGoc+43eV5m0uzdCtpZIfmNDL/H9RtmIxb4DMXIfODZiBbbKhKUR
CfhTJuzFOA6kOSNK0c3vEK82KL3MoWs8vj6aI+eNqlBBpV7eX++ibkPqjlW/7RyyTl9jtwsr/6Ag
VfmnO16LA2kiPDxoLU+os1CJnu4z+H7wltLKnMGiC8z2DgXBOY94jqjqarM5AiBZWLGelcZznWq1
sgpWdZciAfEuT9h5uvIOpraNSDkcpAl0QFXAeBI3enRxk7qJ/otJFUvWwVjuZuicK6O4LtvGVM2U
V4pEM3LuvTKpZ5iNY+7enY80V6o7xrqAQQIQhmU0wJN4lBITGW4cPvAPHXkBROrDqBMs5cAfJfOb
g+nhuRKmVnSUPGSwLMcn3XIDe86p5Hp7bXxbx0UKi8URBeEDaZ5OWEgxpf5zqz2SXg5JLjtsIrRr
qNjAZZXi+LE51QmyTJEWgkdJte/LzYQvBqy1bgtT+OavKD62gyKjcBqh4gv6AFZR7Yxfi9helaQi
TGoXx7gcYayB2xH78uq/Y8v9mFo25AgMsO+8qyxtj4JCVCd8uuBtWO/k9NNh1dxETUPe74/2AdV1
O886MWAMHEwSd/W3puGl2E4tPPzSBbMFpYyCDl3ymnW8S2t1eRnm+A3qbv1IaU1tIQUQbtvx1goQ
vKGCDAeq8bc3m/GhWRAoDEORQ9egEjKSER+rbRBm0JRhGIvubekudx3DIvmdkr13DahUFP5MU+el
vAEJcKU5LvhaR02cpJ97qMfQ0HP1GWKaibfTiQ+BjfG38ke9+AjfyVi/sZcXbzV3Ow3SQ+gi4bEs
JppcJRXp6GIUXVKE+2vLHDH5yYxHoXJybSsVpzsjgSwMgBJC0hoOURwR5ROGriigTDggyqzUhCXU
JVabCBs9e3rli7kZ4nYt8W1kEgohXPqXfF6N+gfMTjZyqkHKoBcmQxGHtqYejz/q4p/jnICuclFL
eLYvNfkqlUb9/Dqfg7MrP5wuc/Dd1X9kkA9t9Cu667s4LbWcsU+MoFY94jb+N9uaW6k6bF5C0JVx
9gIuHt4XLhfcRexhydfonZzdjpmYXGC+CJPnpLt6LIefMcVzsbBRQTy8qxzCV7IgtQBaFEVUV/AM
8AhUGResAyN8iTSlfd/6b8kxOQUE+RFyZ5gtkXSNlZ8ndIVXbOZtkFM/SiZMWhAB8qyWSSrVvNx4
LtPkk8Bk8x0iRF4V8w8Mu/zCc3Crk8s3qTayK91eKS2xGjbFV5/m8GFl70XbwlxY8jiQ7PlDZ6Zg
7ddnhs3OtbTqKfC86y5XcPSMnXvWpBO88ibk9Wybl3g2Z2AzOM+YPmhNMda6df97m8rVDXQPuAOO
L1LgfDlYSe9nMaV+ezv4OPLDu5ZuoGFb621RKI7889L381V8+aNa3sxIp1Mga7aG4dog+IZs20Xt
2HqpvgIS8JAJPYJOLno+k/P1NZLi9lt9M6qT6U1iiVHe7L2HSrL5jY+p5jpRrmU79pB9Mf9k5qHy
T3mkFImAIynaRg8eeu6i588WIoHGCGzhZMZIBlchdnDkMsgJC+Q+jz+H/Z7LYhUPusy36ybsMmIz
CE49UyTs8Z8dEx5g59Kg+IjP3+fV2rD4oFnpSyarVqdoUZmhaNfA+oEfhoL8J3ld9eDZJNUyEMjx
Y09fTVNYhHFsMLkpW5Ahr8dtPEjYbbGcefabCyeEXI+Dbi1+uZU3F9XG2AACflZ5jnIxDplTWwgq
qp7RBLE2ONjOrsUdBOordDgUxcORYlEjgeQ8pc6sW4R99m/imV52TBh88bmp+rzioz0wcmwWkO78
+FeiVLXCbw/te0v8AyoXaqPOO+FCV6G7zEgLAEWt5P0/7QHfX4exFRUxN3YfKhHcJnsw/n4W1oHp
8xhcK27sYqhNrZbGkMRNxy/XDHSgp8bJDZcEosNRqpmTH1/zbA89j1kmykV2hlwm8Td1AIT1pSMo
ZW2YPgbij3hbq5mnMRY6q4BD8DCpC8LdTfkjKHuYCgWHWNG/VTV+tUKcq03H7JTISYbZRHwrR33m
TNmp9bEmXpbQY6D1gewzcYWLzYhBS+a/nnQIiUwwIaGPuFa/CBgZQk15vPQky4i0vXt+MeWH+5aQ
rJHHAmAPIARDWaRzELgG30qLhw0QuwefU8YpI8UzpiDZnahNuhaqjFDydcKg8voIGLw/X9coEw2h
JHDzPmgVZoR1ebgBZoef7mdz0mQPu0ctSxNxcUh5YTxAbZv+6Mwel/aym0RnB3FIuMACgiDrPl2l
g5aOGBTjohXDqXN5E4ssTjLVJEhltC29DJzqvSHrhTS2Q0zqWquoo5dzKXWwSV6Nrk4uU6MACwQ9
ImFWsogCu9MupRttDtCVLdikGMAU04tH4XqKsWzmBJT+jRi7vq3Rrq6NH9pYHRdhqBaZFdqNgeEC
P3DuIsfNQSlxFt2dQ8eMICNmhJMD7wEaynTxe0SQulvBlfuN+004RdmCJrEYgNFo2zW6HhmzpgWS
hTywWWIqvMQR3maAZvFtdKhx7/CpU1TKsNChnTrpb0KxQ7+E8wapaDhKSJLoXB9TuPbKr4jlV9YA
ZijHKnUSl3Hk/Aoj0zC93HtUfXQ9hll6VCC97hswbCF8/xtCQIeQ25CrczQavU5Puuu2dhzlOlIn
i8xmhHnTGhbHJGTo8sZ6Vrkbpli2uGm9vX8y9FGlDrlrP+/TIcpS5k+u4Rr+BWD7soiupDuPWuCL
rwb0cxDiFTB+RYWv+ONnLoDlI2YbZkcYbfF6QDbyy0uusRDAfpQ967jo1hz9JP9PA0EX2G0W26fT
ib7ueghQTkiNbaLLG6nkeXU0hs078smM0Dch3CLy8a5ujLAxcts5F0fvbYxc8zkOsm1VlT8K5Bh1
CWCTDtTNI1me9uIrtNaRtZG7L6vJMTe9Lo7k48jHsFsj+6JL6mGhwhnEeyMXYN6tKSJHP6mxJHM3
mNgReRrCL5U3R/4ntK89/k2oD0Jo1owqCIcNUlgzgyaziGmiHJQza7dKP1HvPc7+5oyOYx8J7bww
Kej+esiWYlruQcmjUBKaIfTYUPt/+tTpuqiOuBieot54+P+VvZB2jyM7fkXn3L5bzPKQzv7IVdR5
4qcv2Uxiv/wTz0r1RVEzb+e5d7lIggV/B8Ki2Vj1nCbq1sx3vihhqPqUT1A5UgFa9JV4jfXkCE/8
cU0+1aPjJUffLeMdS+i9UpjjeJmX7wZWNQntjOMaMz9T5fzsGjU0Fn1dtsNB0IF4TxQu2pRCxvLe
oniLFkonpAd3Tjworqy8J4bj+ijReLINxhSNEZIAhxAY4c+Eb0aq+9D/h7F/eKBhYZV0wRryMqkm
TjuMtSZbU6XYCZqTeHDk1Ok5+EhonaBnjiTd7Lzac/cEZxjxiarLY9hjg5IPggjr8z5F67BnhID8
TTfZNCCL6boiXfQK/CO49QcckbmimwizfKkWKv0D6GKzHHkhy6qukUDyscFmhqDk7EdJnHPELEgR
1itAhpQjOzcCYMjvnXQl1Jyan0ROnbBfIMUvr0NtXVXtPEyNLP1fS5TRnsEUTCSyHimI4nUPecIi
fvl6ZOcfKwR6o4M7lBRs8CBWO+qdbfOgiDDiXPbpQN4oilP9wxV4wNXfFey011If2LgNQ4QAeZt7
b6UfEOsyFZtL+iXh4mZb8pQQCiOuvkozP8TFqBd7GwWKdkA44Mfapt0iR6vHc462QcmL/LETNWD3
rOlZNKgGo7dgBf63cqSZLADQ7pa20wQ7BGr9YsL4z5igoE7kWPSU0o9NKRjelv3haZfxcoQMehxN
HO21uMxFDQy8YfQbazPyT/vqZHfI5xp7S0OJeJPrbglvHdWjcLmk8WYxUWbR1r+U82sS16Da9pKN
siht2Y6XJYub1ibxiW5a+VlneJqSHQPx5/2iCI8l6TV17ltsIoXKUIzrMk6OP271EQ74/OYlaZhQ
m1barXPCMR2h9V1xpYUDpTbiFVae8bgdftExgr5d8/EkMEAjIr0mQAsBqkOyjrx05B9qPIxs2cYh
yxYMzm8ij2nH1iyRqmwEgIHPNFee0muu1eW31nxq9T+io3GoS1NDDAggacNoItcdAdDAB11A2RgH
MIhbIOWJfk5rAO5DKmqANg7ObDIe7ArEWa19dgShgStJdOHV7fBEmhsv5WqV97GamHZ1+r8IcWQE
VbD22E2jMllcjKj9hh1t0Wdzb4cj32XdrwmYXMV2Sz+BUkPKxYKP6fUqZcaOw29Dttf2jOLGedus
P26PtOa8VzHkKY5kbD/1DXervnf+54lpSlDGJQbziE2wkugNYZJ0bFqfmWMdRRJNPfzkxmcosQsW
KVBoCVxXggZx1EezsKQ4tSXq/W8gWimHrr/WX/imTZ9j5YIHuHvA4JHUAw1oBakRRppoGE7M3fn+
ZVPYIC8poZvWFT3Bbb7COrD4zZBInlguHugmZAi1Ebhp18jzj2TZCR3wZ5TsSM3zx8aUR8BvP9EG
Cq2YkgGW9ja27R4+1eyqD1ewmSW3KlUyUMuaYLOxgFNOZHuDhkWziky4ZXvyqC0ChRVZfl4cOrOU
K3+kfopc/rJbYr6RVkFC3zceqdobEiF3B86G9XJrNn6uFE1BFna0I5+j4gfN5Jy0jsUif/G8AMDs
UcgXSBE3NaqPhJIJwl6UkD2syyYzxCzZpLYT2zmlXgcCxqq79oTvQvQs8uGZ6VGSkgcNpJsTqMVF
MGzhh/8ukqFToS70t8JSZr5mk5SqAErjqOBx7sCCqcE6ABD/GDDDO+52oNBx5IedEVqRDR5vth6k
CLTEz9qwbVgAqalNMnxjPtCfPMXq6RjCaY3W7zo8g0GeLXEB2UbB6Suu/1IMY9vw4dkPcQx+hmDK
dMuP6HgzRGGTDMEG8tXeLOnmYDFd/Rh99S6TBf0o0hciupogviBLvmPJIuQet3sPJRBWi/6w7vXN
lpmC8NH4yoQAp3le2Dd+BgUMYIZFcUJcsr9dF39BKvd7K95uAuruiDUpWbnV2EXYmnBMg9oje6GH
dxgykXrV6xyLvJRwFbQ8fjiiKgfJ963YjESellnNHPAAClK88naRbyB3a0BVreDc+WuM/jh9eqk5
ZduuFMIRzFPfc4BaEJyWo0/mf0YfcqiIgrdGwlI7kBlbCc906avRcm5KPRBD8roblePSkZJOX8sK
wfnFUYhig4L/4Ud2pZgeN++QnAuDVYeTTDsDkVFR9jK+sNRhsOxH8dd6ixq2HnaYZEyVJClf6Bt2
vHxUB6UU6TlEpq/P63NAPBd+hpQTIDbhCHEZd58/VIWTZ5OgPJ4vSe7njM5hJ5IHh+w1SSgrIVIt
syCaWimGPxzfWVjq/lgx9hqovUbGu8nWKWQjS1lAppqFAE/V6O62hyQRpjst2ufTRgTt0RWO3O0m
Qwt45sI0WRMLFMUEAUL48FQL6UuL4fSLrsfZVjqteWHOc8iACqEWNBM2vdz8o2tR71HTyRW3KN8O
SIXgC6tsiBX1wsFCPAfuwa+7vSh5Ihrw6+fVRGMPtDSDsVqKTwj1XIW5JtLj9dy8eWmVJucYBUdg
Ux+KD/ff9CqDTl/uSVwltFHlrRSZQdj1pjb9EEUUzv9hlefXjRJZ55Nd61VAfUc5n+Y9iRbh4kr0
lz0XjPCJopuHyfxC82ECnAdbqDkIvhn6cR6c+Njk79iHr3GVUmSPPRHcBni8RRQgJMydzfZFLKm+
FhU2ris/oaW65x0QOwfAkZSQZSCQqlPRuSc7yPppkVe2Z00xLReHZVvsYrPy2Z8iX9FqhkeXIDwJ
Fupm5R2d79EPEYl194mcqv6oFGqQMzJ5RAj78UBbHdSQF14deS1srd5VLivknMfwVTm3EpGvFcQL
aQzULel9L3lsW81bxsIbomzxQRQn6zPTm8c/nLcqq4a00Cq/A5r9XKIcly54IbBHlUmELieBTunw
jTMV/aOEd5gxr+/6OvedQHtFmByZpHV9/mUeg8LHClKZ0uB0fbbu4qCkb6984n58kxADyAt2CpE3
pun2n7v0kCYGueOfje1xWs4ldNt2pTo7jL2tI11aTteUnZLaW1+6uAE3rSV6hjie/3ktOvq5PkAb
dtlJQsvPunB3b+sOWywHdylk8y7ZNYg89/Bnso6i7yo0OSvdkMg1WjPAWMOyHGHIWxYIohzevKJW
AYcZX8Rb/A1kEIXCyR1roquLVvS+rEis6S3IM0l/dg51uzUBCpHW8JhC2W6Ym4BGkHcPkFGh9FXE
0OrZUQtUW6vFoALvalRPnEBlkebtSqpUVD4V1Q785wYaITzon3bOmSkZmpgzQBY5TlEtItpGfbtq
nzLWWKjhORmmD6miEumjQPTdUFn8rYFFFODOyb1qtAdcX/75lD/qoGbNbrIHdxRCy3yYXJpM/r9k
E8SDIUAFECBBvTYJeFYkP1PWAsELVCu5HBqs22aKyxk+RXauky2VrWG4vde+Z0ek7luLSZ0uFmlG
ip3vhrHar4ZtbsVxV1AjkDiP1dQ4AE0neOTiHuVBBTnck2yqRHRZK0LoRbs9w5Ys4kOXhaPqk00T
yLqgxhJlW5/KqrhA9J4NErrWaRYGHgefeLRQjwQ6Yahw0QDRZU0+ymXiIAokHwm3pPKc3C74vvAJ
ttVEklp7UI1th5xRw71oOsqK+0bLNMfS8dz1TYXUR1L40bynPklGVa4uOee5YfjTNZ3ZMoss9TAC
iebG89fuIUygbLNLGi3qP03MNLtuYvCuKB3qjpXx1zPMBDfrfzSZ0jQDZGYccSftAHQ1L5dhINpA
hC5Gpq/5eQZEpXA1kn/Y5Oy8NnQ7IcNULN2i/7Oab9FpCj3Ij6CUCcYg5ukA7Y1KmJh60sdTJSEv
mEsdrZ9HmZQzBiBImWG6eVcEUafvhEHl3LUTNxgMU4MMX6ZySwE6EZRRqv33jvKACeZlvqjV8dsM
ZpznueAv2dm0mTrlgLnwS4RaNJx5nSkwIfuOiCBKzMZ798P7OxNZ7/c+mY0FAEqH8CLnftUGzvAw
ViQrF9DfRb8jV8wmumXpQw0pXpcL43BY6M+olXdlleopk+kRZCbnJo/NcVAFIsC14huBY2Y/GnnG
hYXno10P4ikPuWtYqoShd8k+H4u9pomrGkcdAgIU8rIXk7JbWTFpRgNyz8biyz684jp2NlX8+uDN
ow+iZglveEFt87FYmdKkSQdvI1iBsE4DZh92NSPqrg/NbMpizwi33s40Enu/bRT87XKm5mZHywL/
JHaQmvd8Iu1NeYw4EXef3OIGpzL34spbzO+lqjwTSJ+ImNDT2Yw1Y+R6LUHYmjmDrV1jqWXpuiKc
WrSNscfyBCSzuVFBc7bb0UUg6e06W/PSzD4Im09iZ7ffeBwp4AN5R8H8POvxHB9/TlmSnsTct2xR
nPz2Iz/J68BRrbmWkt7/TfwgA0GdxylE92gkQIWyt52GJicnUnVXorQGb53PyZVhp6Ilx5hv82sm
hUYpY2EifJ4VmQJiwQNcafokB+L/B/n+N2RUwb7Ss9xFtXXAfcwPBe/QU6HAU4xB2Q2Y+i56tR8m
EhNtBouJmBeYjqLfTH+BvgOLfg/BsoBVB+LnH9CiUuDopx6d8kZ0l+q8XU8hFHO/Cz1GygnknHEE
09SCwDbrbpVb4pNNUNar25T/7142pVcz+ySmmAEv1c8QR6d7UGz0slYFr8myAjC1RaYWiutjqlBP
nA1Uq1sujnLBUDcpN/wYkplY7gG0wi7gloA7LoeFjlBHLc/k2Y2+t+K2udLP1ow+awBzWK3YwVKc
CyPbbbAuU+DDAyHx2igGIPdkgDnVrO/Ph49FCeUoceovimHbRrmbiwR7Z04hA4auv8H0zWAeDPTu
gCKdNH8PJra2HqTp1GSMq7uFq5sv38La6LAvIRPlPUX3UlDQ1svIltl0z70+iw8wC47tp3uIXwHA
B1SeqP/F94U4MgWIrgqdVK7RxduxcLopt1FlVwjdb2WASvuW2CvxbX2F6HFZA9TPK3+A+2FfS1ze
xMt6k5WUY0r8EFYmGrNwXjg4E/s0fdQPoFkPx6gTpVXTsuE5S7Qrypl1vPvnTuok6+Do6QLBSDYF
/zRm+WfYLUi+5rNdvqsIC/5ivJuYdEe90KBfUC4XqvEjLXpNXnzn6aLwHvS+W9iNxvwb9zKDWFr/
zJWSEeU0mAgmitzJa49kAeQ7yw0XOu/CEfKZv4a/gPO5OTyG8BtHFotiwaWuUNTmR/aWccZXp1PL
fX/5mKiJVvGfNwlOcXbti4e3K6I1P990waMCQqO8VTGDKTv6G/63/Pc4P+Dysn9uobzr5HmEoA86
g14zuCUczhyn5XJE2UUf2J+/Db8okwY7MYL3+Uu3goPutL+IA4D4wEWrXIRZm9TBmDnhq2aE/8/m
F8FjtwzbhphMkwJ1bw6U+43Ui1NSL7kYkeUFEOhgH6XGi3vGaJTwRNBkhxJk00dK5X1PbfK/yPDY
iuJhnU6mOoZ4SUf3RU5sOm4TvN7xgY6+yHsBNQ6DEy5+FASDRp6H90nj/i9/XS0Sy5d93tAI0DVh
rDGa1jFFyl7n1jyv44YW4gS2wDa/0NZoZEOcO1sZk3sqiI281yRpFsitbuPXo1VaM/xmmqmPQ0eZ
pFAg4bCT87dID5aoJoWw7gwDy43fmE9bcMRY5oEDrbO4a9hxGkKC2/Apl7ObkJbUbQz1x+GnbaT4
5xBO6Xk6DNAnxLggujAqb3sGUeJYJH7i502yzxoahN5qh/lZyXsw9OkjRFiB+kB4V6+YJrcrQmTh
f2fblL93YDmfjI/c0nDhMiS60exlSUpx0SPjE8veAzoWKvt35YH9YT0P3T7TYZAlCpOGzW0tbfaT
0vAoqkSKOMIch75o4otO74Z7sF5Y2tP88MkTqVNybhc63UbBvwgm8/d93O7jQiuZ5VsfYphEKApB
W7I8Sg/XgkQ+ggLM0IWa5OHB2fV+AiyGG3SVR0JgUU2fozMghcW13AZWIHojCtQrMwTHoBrRaLn6
zGFQMpKbYSz+B+E84GldTqTqC7ZOXnzg8/0f17fAOpFvaCoo6OZLPQo4AnjMggMqntN/ymsDjbKH
oI1KttUXGxTFVBWGlkvLxLOX7uj7cxf2Apmh3cZmUpEYPUOO8bArIvTeil6Y+lkAOSnfjrwN9IkC
wHUmYtyMbZ2YJp+j6TmIWsFyj/iZRZCAQmHTS+I4Q9Yg3wpFlJFj0ET5sXlaHVRz0c0S9GyA7Nl7
BKLvB4bKXbCSIl+bpNIFyHV8SiVh/HmVGghrEHDs/dnMknbQlMx6B8WicBHAMDt7hLDi200kO376
vi1D1CwvZnoqjbhteEh7UPFwXCBDs10AGGLVjSdiPTthyvTKX8EtgSNP92bjYM5FAP156bFwqRg7
qK3O9al16CbIe8HW/8GduXfc8MvTyV58RvH1PZ9ITaHaP37hz+9Q5bSx/ifPQ7z2rdr/mNMqpdBJ
yCiOnBKeyNsdi+n/DKT279n5hWv7El+Lp9+LluSYounroZcb03czlb3vkwSofbCWSvEA4z50FVbQ
M05J5WR7QzEetHG2yZPKm1F76/1kpZO4dhLDbT48XHZtnv2gHybpWZPQNXeQAGmKnO8d8vivcIl4
plzRh0nFnXsNGlCjBM4pmbW3IE3Z15teTIvE2SAv1eUsXbXjrm2+p3q7JSyttoVmSdSD1gu+tbjw
BsH0IcShlEzv+SG8NuLBWTC3p19wYnkx8Y/0+eJs1UzTG15Nbk8xrsCc9HSALQVzASAG3a2A2rGF
ez+/kC334mHKMy86POfcLeNiQifJK/r1n2sYmlSMlkg77a91iPMLpNsZzZA5lxHT0pA5H6hMxXxZ
QigkqGXIwyGmPYb6cvyrl60KCsKNcWFkq/WbpDE2LwRMyfWKACpCfFmEWoItStokD94T94QtQM58
wMqiTla3sD78qwdQ1CO/AmjG12rO0YHrwyjd75d77hcXkq+iMvmTaSKxuPzcedvRCXY319TPK4/s
Wwxm2QEP0/0v6Pzl+VaSZpmin03aX55Oqpav3YwCpTwTFzrpNH9F6u9yOKdVxolXaZRJ5R8u9JGA
R2AmtTr8QjiL1yzGXQ+umRg7FhdawFDHkVw2cdcU7Y+WtQdGOTwlL5t12XXbayCCX7HmPwH3aQIc
N7bmauG0bNtW3WYzB+9RYAo5dkqzfYOHdrGNneEOCfFmGqnLF0T6TQPEXjpcKogbI9GrKF0GHmRm
FmePYpIyy23UzvYLetyGtOuB1TeRZor0h0/LgkEJ15DM6ABGEmSUgcvuPSPs4cBC7WSuiFOxsX1F
mNFTAivKepO4eGsrE7u6s/fSW0G/pP1lcYEH+reF8UYpp+6IVXS0ytrPdjh+viRh8EVzq6hwGzu1
bWsql9jjnzzDoHhh7dFxSM4Tvt+5hFOCD1qy86ojJ6dpqmBoQ3Ns9hQPGGktrIDs1v/FR5XqZCuE
IehS6yW7ZWJohrQgIM6SkzbPfgJiLlH+P5OkUP5kcCGzNqPoC9mYJc1lyC3iukDeKCoTdD8RSeLq
GqZ6nd2BX747MCiuDWwl4hloXUc9BRhTelf5EmVUSi0+z88bwOZNe65I28msDTwIUPmKKMSqIEBS
mu6J6ncHw+Uw2nSfuZXuNsqIFXRuIWz9iCoxEd2+vZkJ6sz1kxOs9zMuas2WcitVmYpEtL1sGPZw
10e43nr39xKU55+zoGRUVNw3E2bnDDwrVRAIa2mVQt69pqBampWRoSKJ5me9shZ0Se9dcb149Ae3
uzUfMC/neHwEaq3duGyCo5QtjKBSxfFsUj69LyEzNVo6SnXbKwrW+UhBbVtyN9oYG8GBmjO/OQ7o
YQSAG0ywfrM/Mi0tQJcicjhhn96H+nEMYLLjmig7qOG6EiUQReJaSadH928KTYyez8LzmPY+B3UR
b8vOXzcX+xK7QmepSuEG+Vbw/moJgQXK0DNZvtTw705tZOHNUvTAdESc8lVB115TQjzGUagqAFsW
AaUfMvO5EEbYJ7pu7ue3vjoQ06Ynj6iNdGfcnF78pC2Ic59koCuXnMTuEiE2B6p6gEcgR/GvdAXX
Xdn1Vxe1DhBdblBhQK9csK6TlEZUlHRbJxGAXemy5ggtnY32twgswITk595VLbEFxD3PVA4M2N0a
m2dMKZaZ0ZtCckcEcwJ5d1GwKMb7kH8rMIUTlFZE45jO1khvDqyxz7AEcyzI+VJm9+oNWSGZD3K5
PkA5BebcKOair1YiG/jZ6JYwcggSDNiD1uzqRTvKa1IEIqmma39D/s12R5dpPdS9CG7+HjJxDAPH
14Kk2mVioF0KAwk9CDkKsL7MoOc+dO62e/pwHYGwKobh0XDnXzmSR6Cvmlc3YzOTR2oXVGNQ+MCM
sRPqVOP5TO49TKwn5A94JZv8d11atoLyoEgu3mjaHswwhH+s7OErJlw7WKT6wp5z1KFJFRsJbWv+
zG91pn8OTv1iG/y7LfyktDX2ctowFUtB1Utul9jZ2pK0xP8dBTJaP854wtMKb08vOHwM3RwbGimf
KNloryrDWoMqHZoIuKyEUr3f9Is7NFA7FkE6cGYApdSmRM7PsTqMqpeZNfoRutOqbVCCSvojsbnh
/7Yt8PT92wJVCEkJAWX7bdAnbtTYsqLUGMI9qfTQTxtVQr6x6NGmP0du+BQEgBz4r0RkQw7F4E18
cmu6vYl5Lbl6rk044gtHoT0yfY8q77EmGMI89X9NCKQ8cJ7ILF48IVZlU3+FEpjK2/PUENBQIsso
8JkbUhoyIGDLQ9/gcaI9Bwf52wp7d0i9EMM8QRkHNvy6yCxOmmvwV5uOBM8gKk0MgGNjdLq7/TYl
L0tOrEYcdtp62h1+xf0l+Ojd8Rt3lY3lEIUr0apdcHsdKlU9NXAh8qbCuKgOyk1RqMa4w73ktT0L
9/7OoE3RYkPzzpdr9ygMEAgWmuaDEgF1wlauEv9QvHz+PveNXM2M+lliePFA2Mt836v8Fj1S2+Os
1VAC2SdTA31hycUrkjjFCVQ/CJfwgczw9JXaTqx9kXFW2HnqhUavNk2FPPZwFwoaiOeG4Zo56VQ7
AWU1b4q8xOmgcedehKSjJb4GZ/IZ+h+teT3WcwdDJ+lDhwW86qBYwgkReR9nGsb1S6YFJ2MK8g7g
5gcSMymdwJKr4mQ6TiyqvUMOlDvD6wP5pmpD4YnSxJwD9Vgr93HOGvuSIxJYyreEv5gZxfu//6My
9DaYkHwRCvHUCmmMlmzeHzLlUzX9zeIGBpi3HASswLdbQUFaFBTAeiXLfnt3bs5zQXX+f/UO14rV
m39q/TWsgyH1JAJpLRjOhJa5lxIv7v5W7lKRU7725XN+5JGQdU6v7zcHisf5wIhqu63NiCc19w5v
oAtfCRlaJpL+l0zrcOs6HaD3avJvSHdEjzXsQaHxxE1d1r8CXNUsoT9w60/o3gQmYQjivrc8Oeui
1HlPocJVT+QX4hzzZM8o3w26jcVuO6ETvT9NgGFX8kSKYbyeMPkgezatSuyFiF64CD9bqloQhf7I
/iHNIqztXG/wXjN8jW8zM0LRLF9pw4Co3iXG3c+V2d6361Z9w0yQTyk1pjqXh6EqDGh3hHRdhdsx
MZVi/TZsgohrufvW+IjVJdIb8T/wxmZWjQ0nt25rGJ9bBwyvxIJWEjWP1MQV0G/NkDu8euW/ZLrA
55o8y1wYzT1b9bL1byLfcLk6bRUICBf4HVQPc+6DTxPtduudpFCfSxNSl7iUyuUj10ICIScKWhv3
MyOr78UVl5X/jdH+qUbyfP1ks1kQ2DBjiTHsKP694byLE0k7miOSQFuYSiiTeTYkzkaMfJO5ZCXI
l9nz1uZiQ0bkZgBwf8IslloZZRc27Hmx7BJP0pYdfM0Z8MCSdg/J7RY7AIiNKzbhdmrh0BhfoUIm
6aXIxAlQELdpqsWYYqZdcCUd8UxOS25IUF+ngKLbhAu42i/KjEmgMTj1GCnMgB3dxEI62YQzeTjs
b3hWtkCAPZAgFy8yFnGsrPoz+ZZd4tmVh49tM+GReS3mTYDmcK0gv4CQTKcGF7ZvwduICfZ5vd4G
Pw+Ys452R9Y2d1+eC+B367A7smavTTJrEsJoEFewMRtA3Spi9oKdLMkZEBTmz86NGksTu+IILh0J
CC1/jmCy3Bz4cMIHzbnzSSB+p6Y/sDwNnyAYaeyuNPiJ55MfmJl0kIcFtJnv0luYv513e1c7qr2T
NaiH609e/YkfGAVxpICEIJqGjmDcrngg3DuMBY0p+NgjUMbzcl3IxqLBxmthRd+uh8WPx1qpkCfu
6+BJo8/hIZYF1/qmFBoKiQpzirJM2Iuv9V5tuBHqZOsbtsBSRKBJS7QIlG7f2ZTsAb4IhCTSVM/Y
NooujZ9c35LW60mTqnT0t7yrEV+bDK4a9UlmZWP1M/o8MyYeJnum9Zky7/juVhnAzVB92mCGkCZe
4oOVMVNlgl5Bk1LSyKIrmvmK7AylB4VF53YCiDu6tpbHdAQQsWEqhLXeL/RhjG0E2+0tvQwyZwA/
75J98K+tTDuy/zO64w6FjqGk6GgoVFztwwJMJPR4eLqRKe26DP6IGCvF9dZwpyNA4jo5qnZiddrG
mFf+AngxPnbIAAUeNdIC7gNSwmczNJ0hMqH3KuDJ3ebzA+1MyLjWax4JLEIEsPAR0yAab8UxFnbm
S/5f+j5sUzjTcdCYMn5rS3/rrxn6huusivWC7NpJZ+GA/d1ehMwdlz/PUAj7loEzDHcvR0wBbF+k
f94udCTq2Y8VCffJR/79c1wFQbLbDCtyjrSSMnjS7EMvOOACBo0CI95JDK5dZvnAOLB41ZfY4SCJ
0AtGpFQHLna51Kd9/zFlBBZjAQkNVhgqrMq18KeWucEc18GKIQNE+w73n45ZnBDeOywemfJLIpSY
uvgUVle4HnNHgGyqicJrbfa908qkoZzlSOnI/8v5xHkmOtYbGyAKZaloABSiuet3+n7kNfEbyFNq
/T3nCAIHKMvGfwIbUaG6FtLoiSBWohOJj+BvGMrMGK4KxbQ1wyFXxFk1dqa6oln6ooof15kZv8eA
tDetvW6yZAFdocGXWTDa8IAe1uhfyScGINEb9SO3m59TFVrCvG/Vh6KchHbTB7cRpa29JJ0pkssU
GSGoq5r9RYNiBe+v9FGDDmVmRIAlY1S7/9QnaVozLHd3sPkLFoIJegNwrYvUYkrjIUuE4bzMoELE
OZ3AE5sTgI801y68CjRWBMIVmCt6zoVnlzFXeYY8XOrf2KPcr4aZOwQRtfO7DJqo2Umm2lsOk/Dv
hW/ER09UGMXbBGa/yMPumlz28PMvzzX7cvN1P57xx1d9EFfcJtV2leLMGVJwpM3YrGO1ir6DoMCp
iZXDy2HkPbSiM9k75QYRgATQ1SH2tA+xpwoHooi0JoOOUq39LUUeZWyOHx/5k3KIv5Ca3XXf29Nb
/0bcKiZNvsi6gjgn+Ua/DplmvENTYKiiuX7g7ASKnyglfDDmsjovzKpjL/UjmfLKzFwkZ3kGOcsm
DwlrSB4TmiJLNPm/gjluBI4Hk8vXoRL/aPC7a7pmHQCrUtVyM6nMLtJdyjYcuz+A8HYH9bZiDiSN
UyHehsAD3Q8sWuvw/HhglzbteYjqr2R6MnJRDYp37fJTcP6WxH6nA5JH7vueeinzrYjeNMT0Y/Zt
7dy8YQwJhHXh46PeKt89c+IodjdrMTZLsPoWYHXQsxq7tnyv95WP3WyPvN2x3RTqz5I+HKYiMIZi
9dAZbY31tqoSCuVrRpyG+hvQN3FI9a64RNOId9XEs7SQ1533uFnJ+CtMboyctwPipXf6j5Rpk6B+
J5xDq61TBKdL2Pt82nclWhr7WxyK1hwErsL9SVE65+pD9IonvCuCBOFK08j+RPF0dEt07OZKuxgp
C25QvktgRMu9XK9pUocqhuRLZgZhqbHuWzRebzTc21og2yd1WweGOqcXK5hTpOJ+56ZLWT14kbLY
bcQP2MjvlixFCpzL49HOF3xVcfDkuDPvOjUtft1evuIlpPi8zvv8MfMTOMXKD8qQGPpneynmBuvJ
SsI0BF/EYxj1Mt/r4CgCci+UfskFxbD5QdpaTMywfW716t43reTAEiF0v0MU8Rb7l3qZ76ComZ2U
Cq4SWObfd1aVnv1gtJlD4zccQstxOUEQPehecO1L4Z3diuGIEm9l6rdjSeFGVkCKlfXojbhbF7cj
0NEOpzWC5UyLF2IDvfRFnx9dEOx/91IUsFU37K5+dsJvgsYdpQNinipOuh3Q9WVPtvxoEu4fOWV2
m3LQLSlfhcbeg9ODMjpLrtYH7Bw6PgyjqqCvCQtIvOoUUi2+3njHvGkay80eznu/bvJoR5hDAvQr
MxiclEPao3eEv3dMI4D4/Z3JbebJ0qXrlp+eY/nN2qJPp++oUii2nTKPZ2LsuKIJWPxT7N8kHqSp
UJRwGuKfe7yRM8j3iT1BSd7/UPKEjgZkvfkrNRbyNFwAylMNmXrY4mZxdxyrKfLA0W1k6WqLPS+1
G2DvgwK73JygAfQfwrGdCI3JeLc5p9rDtuh6qOZ6+XcSf+SpRBb4xZvKLMRLiUncXKCfFyrU+gC7
tRdyRVFIUW51TUNvNHXpBVJ6FSD7eSslq8GzY+wJPgmWdAP/LLmmJXOA27x3ppeRhP+KqwEBcb82
VJ0fzgHTXVZQ09cOBkc1qXO/OW7b5d9YND8CMoyQJX0s+kCjcAB16xvAUpI6SWXzeH0ixh7oLG2i
4bqzhLz8+4FODeCNTSyJzJXQAdgYTGNtax/biBc38kHdXRhVukVfYtZbr3mQde/2Tki/HWP38Ftm
mMW5grs65QqfHJOE5gLzdi5PzpZ+6qe+SD9GwYtdFOqwHDDDI6TTYKqYh+4RDyHf+QBcHyIxeJLz
tf6GsiNqYsIbWwHMvPCNLMIfIh9Es8fZHgcZDCxNNhL1t285n/EaPMuGoqMfSHYlXErllakxTxp2
AFkFQrfcQKBBSbmCzLR2k2fAcU2bYb0FaY/T8QlOL2I4Jw9SYpNdyzZpbeP9lT03IgOrBkGCQFy7
39FAH9BRC3LzNeCyZwZx86VQO9QyRc2FaW7Y5uGTD3XRLZ9RXAhcSL3Z4cq6hE2HxL1JyejVKJd9
ym/3hOCvR1KCezFmf7D0dlvHC5FRVFjvwjrKRz0Prxu7NdWio7tNRpxkRZ9GQn+3vxC9ckaOTP4b
QzhcrB1sVytna8M+X+zbl3+W9qhGu3N1kF+4Paljvnfxfu+TstfRmxWYnfd8wGCZuEcdA4tYGXzB
ahq1hbkhchgrY1GdoS5IqI3cGa4XjHFO6yvF4lhMyNPh+sbYoh1o8UoLvhKSyVRmrRkHaqoS7hSV
pTEFd7LMEMNzw9Ju6U6G+HSJfQqMj685+j7VLDMjN9xfZwGk+cCL1MM94QqG/9KAHOqNS4PfVgra
jrYW5jRz+c/2ViL2lfGzgXDXC6FKaBSlfc1Sqrg2wdRIo9YRwzgpnaTRSrHqfKftijkNl0sRBijm
HWENq1OP47O577Med2HuiiC678S64p9oCVSy20xzY1iLQQSyLaeasJZA8WHlfUtvaVszodhrpjqN
PZjsPVUsTm7blEdOsIg7bMmpoBcNnaNveDN9KJpaAQyN0FJwVmlPzkWjEBahRPSGltnW0WLXtbNy
ARLhn0zGFliUVPV4rHV5QzPHl164YI8GBVO4rdbW6MQviYpApT5qzaIr99tmT5skQbszDM/VK9TM
QnPJbGkirDPipzyGGmhHF5tubrnJBcKd8odDkjhlw4RIf/l8ZXymYMEVcduX7jypy+nQihDwHVwF
MNEDChRvTjswj+dS8QwXczSrdtMvRIAL0SbiC74C3QHN5xE/QPxMWKg5/SrjmZ04GAkSNsLapkEo
TpQysuzdp8DNQRW7haJTc5GHDhbgVCTNsZqLwD9YjA9h6udZ6cUjhCjQ3/RntDDxebt9tpIqTBhA
JqRqHG/xZlVO5amw+BVcajtU8twgMv92iFZTTiHHBEinKbPGMIo6SV4z7J7K8hduxYwCsjNIKAPZ
zwTdDTfKWGs5HOxtDA7COrAqbrqlpeE77sRNvHImmzapWdXwR8Gt/LDmRzP9yYgy4npl75XMD42H
634yexcSjXJNoaho62nUY9I5xanpLKsD9WdAFxkNKL4HdViQWdL+T/yfXLaxRIJpiqpLDXDiruDk
fRGbmt51+3AAKz//sNsmfe+7C4lfabZnMtBDs+zK1TxT8YToVbiNZ9FJj8PPFza+LSgZRiC2/cbZ
17O2rMSOoeIZDgoXbyRFX82RD9oM1Viz1pUhDzN473JFYV4/6OlAHTQVw43WZflJFuHKa3EP49L1
CaDpqd0RL5PRYNtPQfPtlzhDrSkS3z7oE+e6OKKbkCfd0F2eqUzMhLIZn/UuF+VTeRmx7YHXXIjh
Izj4h0V4sIorQ4AOGwkuEPvJ94CYJCFW0HSxDFxRgU4SnYhcWWzQ/131pR7N1pnUoOMV8RVKDnLN
4ib6XXrEzpscXK94Umnf6qjJTkipReopRo1YB6BDvhL2vt39Sru3RwfxKea7A98VT66hK6ZuzMaK
7uR2REo71DofehFSMm+t9jtTcVUc7DX6auVNMIqsOC2V1FkstQYyZv7sf+aldMaruLafiOmhg8R8
UdDFbwJZzhFrSvuhFoXwTgsQQXVFQkZZuLCNBazAQ9ZeOmi5AcedlgMReG4Vnk2htPCXqT8qHjWV
MuCmAju+OArm1jkJA49g7O40kY8qkWsNDxxrG0oAIx28nRbptFCPJXTUo3xgFPKxMnfp+l9Jy1sa
IJCMitdiaRuTB2kRBQ+dZ5arzzyy5ChQ6QDo1MSzKlvVaeqOifFvqhQ3eT5tBHzRJloljzqzBFxl
mtN/ZQvG7wEFlu1lydPArsiWcmIaJ8ga3Xow1kF84kGPY+hovQ+hAhw2AltDs52Z6S94p19l9zFi
08KHTDhK+cSdO9Lobfb+GrXqPk6cEpr2W2/4xV/HYbJ64jwv8h9SNMjgwr1qnKIqQSSL1vuO/0PI
lOROlKoz12gQDJDl695SzNMSStDPVV6koaIpUNu9hW9vKD6HVxo1v1Izr83/ZSPI2dU2IzkHpvT3
pa9PTUQQn8LB2CRwC+evO9HD02z83eLVGKgOZvd3k7ceiRYLT/Z7qZhnMzsUgGIFY5tTfA44Y7Mb
1fBKXL/LEfbEGiBc5tT9RzwhFilySDd9TS5cQeR1ycJV3S8gmVmVWe1eIzCC8/dSEm8/U9mle3qm
9Hq3qYU/49P0wA75c+9PojEZN3vOupOoHQH3S1c2xW6AUfuCqfGifkh0npjP9arZqqFZZTjKDqlr
CzPLMnqbnjw8v5Vxx8jMHy49nAijHVdzIW0qNt7OS/LuwTOyOrZbt/ZhFd+90jIVYeo9KNrSy+Tw
rqqpIapXlLU/PdsAnBPEalOlYh97JFzWGsiHu53xrICSJ3znLs+1bP0A+MTM9ZJ9aUuNygOt7n8z
KhSkD3lmlQfQlHGz1/2xBbPzK925qc870ISszNLFGibdCAIp1hDbxY+tFRoQeuLpACpagYkIJKcz
5WfKOXrNeNiSgs2ETL9RcgRcz7mJ3hckeo7KBK6CwZgPZmqSNujI1rMNktx0QWWIW97+cD+L8TiB
ombcYBcy04Zj5NyhcVdMl/MUhfn+peoLXAeWf2dNZlckc58f3bKxCbAkGuSS7w/VnaC5iJmlN5zG
xABjk4GQ3/CisipbETqhsDdvQwlM50PAsP7T8+UnsIkHBOhrcyxkxdx4LOlgwrzsk0PX4pSaGKKf
RTP0vujktXMa5rdD9VKRQjYd7To6vcKSFjrUFvhCuYBCTctnIo+Ned8viB84SdtuJjvcup9xoUSN
cFDgh1fQW/c/Tn5FlqzVWcb+uMGtD6INuxcA1TfMuynsfG8idczj4yVcfRXb4Z+OSrWXPtdmp2Oc
m2tlO8GUxqJN7utKCJGj6dx1iTAvkEs9wW1jVHrN8sDp+2q+yGHPDhUmTr9KjSd5JbY3soyHjsV+
bU+kuCYKRcBDJxNkExxpyIFSR7Y13jU4En1luAjtznw/dWBVVfnXzJhmBzDp8ELocbEMG3tJWS2c
jgw3wNwItBZkRovbZieQ/Sfvw4/UykRHfMq1AqIutLP7DhrC1raKYI9EPI/Hv6MyZ2+Iv6/fw6Uk
QOrpm/F2v+KhrKy28Dt8QpfCO0JBPGbfEj2aruuu2l1yagTJdtGE5isBesHv87/7z6y0NRSNFlcy
SG+CddcdKnDtB2yk5vTx1j8Y+P6WeHzeNvc/4Q/bcnbPSeGkIfb2xnMTJowqDgGs7hrOkSarWlUB
lZwGNkhEYXPeaVjz7ijkLliJchhhclZ/GdTYEnCN9pOLvv/HkYgV9y3sihxdit4580o2qpVl+C15
O4LH1PWj4yEGLUVXiAJVLR9YRKPRI49f896Fq5UVqUa9pDP1++kYAggagzX1VyyToqdOGHX4kmQv
W/XTYrM6uBSbFnhIoyO2WlBey0zS9412rhg3oYJH8TzGtQmx/C98+QHoZkoY/leDsi/IGssNUQjg
GSnyahxfP/rtkXwFq8SYRZJdEP7fX6+x1G4LOIOCJJhsImySQ8E3j9UJw45+w98Ka8cBtHR3Tm2h
xs/r3v0tRR2CaOUxlgcJVRjmSV0yN2PRIdZzbawuySrpWGLkSMDwyzGIr7tr5vl1vhcFcUKLBkwU
WcGuY9i7X7dVbVB6eM7hjNz2MmxOD98hyKVFZC3VLcGDh0MUn9FfxUlXeZFqWSKPd+75/4MWnHE4
MWDxMbeIP0UqEgNDRWiwwZWEX4qDI2tDrv0Apk4p3HEXNAoiyx6LWSNeFlPEJLBte8knM2MpRTCZ
btuwlOKuCuwiFapkCFxARbXdTF3TPJrUTZ/uCtdWcyCrvMOQEstyb2b+5d8s8l2zdDPXlBjUImdH
14+Pk+X5qMVPtJS/xfDs2tJv7W2zeJ8QlzHQAHUuuwr1WcOQHjoI998MYLaJkgckIP+Lz/3Za72z
pM+eckte2N0EBZqT16yVCGf31h+a4P6USaaFtZ+irxMq2DmHBpoGiwOUWTe5JNpk6MfTfcManYEc
i2AQAisfmgzuB3V7N87SWdHq/4LSxdh4R9dGwr8cMVB1QZHzArNBh5nyQealHboQ+xCqK0yFGVM0
hr9224HnGMj0SycL7oedd5Zi0Vf4Pz3py/oMJRzsjlLLwLUkhyjX264AczS9srSIxMI9UIWX0IOI
ITysQCfO6CbC0CP6luwwucuC5ehntun+eDhLs6kJKaMOZ1KuxZaRb+cjiYy67sxYYaqil3xF9iK9
LJ7j06QNzE9WrSn4eOe6nwu1Gt4plWrtNVXrwQuzo7htBqEx+bVuhZDJAkXBZ+zM1xmzAHAdtIqe
lKpXaoMwl4hlpsctCVgSq+IMgPUouzUPJ8aMzc513t3CE3SU1gwuhye9SExOX6tray/ppE7IlPoi
1hnSI/GESyJ6qsHOP5/TVmJPkRtOo/czLVa8yr+GbCDsEKpNVVCaFvplp9mQgWstZIrJ/ylDRrDv
YN9410AdaiU7pAJq3STOaFgiyaUXgjkFd08Bzdy0OCvc8utojFr4i0gM0GzW2ZJmcX8zQMull/9G
CVnWLcxdPevyClXJx78y/XHkzqUe6+PcRzC/j4PSUkhsGKmmBUf28nDawK1AnZAnTaprdF+aixF5
Xlou8c26KsWCJ9M4gRT1QjK1H5Wv97TvzmWxov/k4CZyl1EY+mvDB6hAtMRyqRsXNd4A0v8FTcGl
DTSEEoiq1lQkuPb4/PUNSgIb4GSLyGl7qajtDfb7Fm6oYf3U3/PmRdbeRo+wZkNbpQwey1kUpIHe
QKPDqNi/OmsxPDxpYaSo/GoLVpnewlijC4Zqh56NMi7cpvEzKDIu6VOuksKhBltJ/vQLyXF9hzkM
6G2h5N0Z614BlTyZe3J9esBbMjOsgndbmHhfKTDIhIapWxGP8SIWdZKik12a4XAYMEm0vv9EC7Ja
QYa2c0BBYL4MEVuJv64VLStbIl8u7A6v4ZDm7r9fteEUQlsSCa45Ar6smJAv3IzXbVv8C7g0zGmP
i5k7TWu3hVXyIuMoGWRugvpZRN6x6uKVqu+whhvjeMudn6Jp4PhKGZZ+eq7Vk+k1qHsuMeLrZSZF
oI8ABAYi/613F9DvR+17o+7D4LJu8pt4YNVyhVWENf4v4zOdXGRtnZzTiG1SEe5jBSnEc1S6btrX
HeEYCrUXKQ7OgMqz/4ZQUBj5F5e+5tPwZbLL14XOb8iH1ZYnzpgWHM3gfwiPBmVAi4mzlKCqFzEL
z0Zv5oUq6sI7oKwA063LDuIlctepY52JBoQRGzEFbaUWTk6sKVhJGx7C6qpca4vFmtjBasPdsYTj
HzDWnHKOxqX2MZpvZutHNebHFVrKDGknaGiXRjecal261BVoUhRD59YYdTz8E/NXmdoy7h4p3KWU
xeiWBzk1wC6oaP+YwnuvdUcOig7lYzL0GJCrO1gcUwxn+gR5xDtavSJw8aI1tHALtqiLFy8tlww1
SUgLhjnZwoig2FKW7vtyUrLD2RzyudND4J4ZEPZ1kzxzqyzW8RqvmvKmRao1KxE9Fk6yfUrD0Igl
ffKD6C9O9lkABKIssLuRQ/diHHlTr1zIU7KIMGAQsPFZvwBkfeWVQpbdVePJsUwOwZh9wpExDbhD
zMSdeYkhI+Y3c6vE4K93uCunHALWLwVvYMNBLavZUndt6ZykrgVu8dUc9gXtmxOTJY7TGtsWmfxR
D/QnOoqMKHOnLDuIHHdrSChXzZQlzgssL9CGZaSIbhK/H9ZuKwcfgvY262mweVdKXw7hzVAERl1c
CIVp5FjnIRJKNIz/UyeRAhFqdiqJLXo9Zf9G4V1G1p5MRZOLw1wMsVctYl19kDudaCQ2YZsyLGvN
1kyu5ntZsuJ7/vcirzByytfvKqx/h0hvJ9LWeYF9/+ht6CuTtRWR4K2BosUJs/ZP6VOejmKwtkVX
gAimt47Md+CcMW31lM/69Ql+4u3cj8vlzXkIfO+cjGBx2g4qrlzHiaGAkQzGPnNDrkWtN+ygUh7g
4P/X+YmNJ3kUz2uYEMTBwmZh6PiFA53hyAPvImoLEd1pQbAjyJO1o/NGGHrV4mkH10HMo+9GKnQo
vHsHqY1hQoyRssa0G2DmzhLdA0meS6Z66K47brm46XWErK2J4MTkVWNH5PrsBZIWSPajXdLhYBtr
huEFg0UrIbjYgIKEcKiILIqmNc43cwLpMZdobppUa2I9E41vaOL3o249qb1AEvFl430eP49CT4r5
8qWsrkpB+2JsO81nLMxswuXn4HyDKstBMa/2JT6Qn/kqEinVew3T8zZHXdRNyrmgr1IakoKdCnVy
Twrcg3vXd0vfMHFVBbMnuANe2Zd2VObxv7BJCfRIpT9FY9ODJBRorNmFCuHs0E0B4DPSusY64xGN
VkGa4cM0KYMv0HHofk+D99kJQF6PXjJ8IaG5bLlZTPND3NeeycVhDLvtVhbdlh6FR57fbweC3POo
orrGlYdu3TujcLR+TXuNAYyZqLHnCSNLXfC/K45Naia8b6tDYhXLCtew10BlFUutPKbGPqvDPaLz
CXqtnUmSgVG0kxgToABEq5YkVGlyHAKchiz53QahMjv8qJuYbRyWIvieN7BDYCpPjJPDrJ8o7S7W
4HpmMpO7EFZMKtDghpXaExk7NQLb/fyQkmlGVrH5IUWHiNd5x+PaatpYJI4QM5noxbFl9oD4MuFF
gn9U39Jw5G7qc92F6BNFm5qNEEFjaz+r7ZrPdiSfvmONm51cFj769rNveT4ZhxoPTUNK01wIlcJh
Z13jk8k9axXjALhi2UZ0wtIgcUbQsB4XlFYW1Sv61jSz1BdiQbHzhjcj5NzfzE9GMj7jfU6/5eLW
481n7dVbnl9B4UW71H9wbgplPZe0g7qkC8BXW1EnIOKhHdy4DDb9vEz88Ls4Y7X8PCAVgoKPN/oY
7EsSN5Bw6+O2vtGxvK6AiiqXA3lbMU7vdzG/spgcvxm3wrn+m8pfXsEWHZmz4VeEqldg6ewC6m1d
m0fPs0Me9laiy8xIyF14kVIbIZUG+Gt/bwGH3WG8STt+Dr/gX4I/0PIjL6xb5ghsy2DWprrRMpLj
BYgD5PPjGFO0L2F3gI+/Xe0wURpLeAEQuIHPWMCEcRD93jp+tlvDF+++kcgGUJhcVMXNaEEMZTc6
5KS5Y080H4eYFiqWs/C5mgV3QNzxMQVc59IfixNpTg7HKiexlsk2LROoO4dwqwtPPbwrCgEZjW9k
GULg1j4MducEngYGybP8eaVVFZh0cVC78/bvYWuob4Cu4sKoc+KieccHi1w9Dy4pYuyJrSJjJAFD
V3sOGA2Hy1THTNF62JzF6rdtCFanUUI21kRaelpuiKzyy3q6FwY5vlBjUCLn7r7V8AvVjCNgJYD6
vQPn9YZ4VcNyhs4+qpxGk95wY64sBlQpJYdHt7PU74O6mR8RDLv9KP/u2bOYUDyLpYZtEYMLYqjd
36mpaOC9yYWYrMCvSfudceAIb4OeYRB9YB1s/4AhTbl+WoOMlxtipFZOWwmo3osYu0OEALuipX6p
RoLt7KrK5w7oH5tnHclw0sPNM+SjTt9gAdsqgiwFjB9IOIxoraEOcx3CwdTrSWTKxYyarR3EnrsE
8++kLygIOCs8lYrcvb9Bb7n2Gj/D3QPpAPFIMUSvDtdTOYDqyiBTV1lnnUKDCZ5+OhCAeljFJ+NU
sKNjUZfSxBbyzIavFPzfnPDFry2VqZwuLNcNaYPBH7i5lUcDYxWLZJjsdVbqT7ZZJj0pn05CyzQ2
tnSrnEiqvaQCRk7JC6bjVS9n5aDErz802e1ASlHvA5Ijh1fF+0+9w6qrS4Nzb7/AgKAk5QadJkZO
mJ6byUFwuIR2kgN3/LA7H0iKMWBoddW0vVh/59qZMwX8/b3JYeQgYV4WxRgSnZ6FsWOz0aceSWgt
PXx1EGZo5LdYIZBvssHD4+7KtH9X45pUzUiR+FIFedfdC+Ga35WpaYb87E5T+cyMhwwW20lrfsW+
sUGd1zRx8B5XXaeNwTCJri9g1qmDvUHwx/o0Hn1P+Byiplloqbh3FbiJCrG/l87fAK4QJ7Ay4L7t
nAvcxMeL/bhiKcBfsQbiOq8wu1mq5/8lvGr7yfRq/HVkydbMeACbCZp7MU6U+/gO/xFlNNCgSm55
rKV3u1O7NkR9oY/yscjezYTg8f/l5dDsA2rA04WiqdrzxeaPzbRj8XGJR0Z6cpuDqN28a34JIaxy
DdWm4rfgyoiGyTRCLGxg45jAXiFZe/Pkd6vNRbuBz7qFlKySMuCX4eC/o7oGC+5hsN1ZHPzZ6cb8
X+4iG+mMRlRo/8M0BL4hAmzoMFVLKk+NoZNE1b35hqM5duaWFlnEBtYCoA/X5YH5+x+7gDR6nRLi
/MWaXczksCCZCaFNNnXlyFg0o2qNn0bu/D9lYX0HwpOOdshLXxHyj7JwhZGHNR1wRd19pXhC8Dj2
CbLgKyzsWRQ4HzlPoqER8hy8VQsjdGWMY7R40fN/HVwrYP9BONRFCqLsXRncZmcXtTAvwevxX6U+
aWI9cUsHjxeobpIizpSS5p2CJfKkb3gZim2/3WiS251fppP21+fcrU8fJ3O7MQA9cHpHAwN1CvsM
GA+2HwxhsgNtRDiAQO6B0nyl1A0sV3aN2CHqpWk2a+T28UQKjhpee4LLNZaOaoxHZT4XJMrMcXjZ
4wknHAev+xYZjQkF90xZpfxjOqnrjjHYiJrJp3MVeFhilR2ojuTXO1oBUwjcvPJg0/ajlRRHGJDy
DImsLX06uCnyOyAZW0hPpJbObUtf6gb6FcdhvzrAGmMj8nNVzvZjwZqYu4x/rjEoX2znqXHHVMRM
pWgQdIV6P2GOSo0QTresYFt7otF8nQcZZzSL4ius7FmqeIk7ffKcYJGA7CH4n9cFQqB0Y6Y7qEbn
Xtvqnybzg2HbHRpgS6Ig0cdH6GGEvK7EAw6WE0zTsjv7WyNOuyI8Gf2viYzJX8CO/bPK5m1aa6Zk
m03FmO9PU84pheiYtYPb1bixaY1og6wOLSpFVImz2xpHD7OIgcIApKqS8IeXJS+ETx2k32s1O0Ie
rIRauudTFD13gS1YemVc15SpMSfspJ7yOydAB6fqBc3XjLpqSMaQ48AS/uQ8jWXWJ53RC+Ql9Mpn
iJxvkztRe6qRrQEl2yOoGtOXsPuVORNogBzMk/EgydProCU55PbgBx4y7YN/OEHKtFTkhw3fHQlO
BQ8Plhi25VrDkJXMUOl0jh4ig/rys0DKKmJeCUsCb2mPQGKByGadobBfFP5o0vZ2umBfEc1ca/Sd
p8dxtXtKVPM7fCWE+Vbx2sQRaHglOz6ovIg09AKme2aVzYh1TXfFArweiJbJEl/ubzt6S4rrgJVZ
4n24pBY3U1PbxK/+DX9AUmCPhBAYdLb8xb63Sgnnj5SRmSiiNjfAMvSZ5wa1zj0uUa2y/O5lzLPn
rbXS2IglP86c1MPuafSkU9Z/x0KophAcsJvVDz/ZyyRGAFtW1NS0oBu/jgl/aSx5aCYaT5y1YrQD
Iy0s2Fo7dtVpl6wsFw++ta2kTW2OSC2lbPbWIA6Z0ob3OAiFIX17B72dK5mu0/E7a5W6uG3kDKng
M+foZtA0hc68uAovD6qLt0e1O5tsfgMREnu7CWTrRMpBCB4M0XLXTiDIDEm/oBUHIoGIgSGd4JAA
AfJuhVRUpJPS5gJS9xbLxaslOF+OLcj/1dcuymRQMn1yTAkebPOEGcZxAWBoG7J++UqJp95m6iw+
Rey+0wxyNTJXFk7tAIirfj6s7+lIV0YaVA4Ld+XX3qvas85X1AMvm4KjcgxjnM09PxDafW1T2ImJ
XaNWyWr4t06VKde1Oyne2rvDzdhkAWII/Fn6gwpbIkxJ+Fx3UKCXR+I2PhxYDx4JCdLXFROrkZAZ
upZJVjvhB3LYs/lFr7TDApsZn8dWr9HwDxpGd3KwePjLBPH7GIvC+RCbpLLfwtpMkOA9qnQ+j0/e
uM/9wZUPHkFT3zW546QOtPko40/H+JIQj2VYdS8exO47eZwr/jqiYJsIWwbT+CI/4P0nWW1S9ISe
Y1xP37RNQzGOchr42rYDdC2ZJG7rieHR7hQ6zZKFNfma1ikByIi5r7l8qeuqSjPyibHC0DJ3671G
6sJZuVq49gt4hXCbj2K7OKFouOk0D2y8FU51QVpavso/ZtCbL0dEihdiVITFGL+u9bQ+sOrrDRzU
Mbcy/Z6ASe1DtSnVlDCc71H6Hn+MKLwpbw5nfIXhUBcQN0dHE1fu8WzNQJxCW6I/kA5IOC1MTtmM
bnFrDAMHxg1lAPEo5Xh5KCWgoYqmnsEOVBFxuv5dm6cuMMkkjCAqeYo2nI96cMWjm7VTGeK73d29
02+S7qCQR6F+BIZLOFw4xFQuoYXQGg1dEKCxsLS1HOt4hWEGf0UGFp9I7jflj4nnpJlCICdrJkUX
VqcG4Jt9NvfLY74WfMQjSwnAIrGHEzTFUeEjXUaJC04A7XSEKzFzj5hfL1hjtQw0pDSsZM60zTGL
F8hAmH7bkFOSFob1K+AtJjs3GOGuM+Rd8gl4fiFMS/VKHl28fPl1kq6JeV9/My+69Edht/+B9iP2
H4xmZnTGCST8tr3XlyZeaqF+OxJ9bQi6w43ESNUR1GxAQbXzuzBuZ7KIxgumtNeEejOeBaC7/dXA
d1Q14Q+9NLLWM6IaMB347UOnh1ZKZdOdGn8RA4QtLXXocYl6SY72eR84zD42yDA29eKVKB51EhVm
p9FBCZucEFOR1obrdzk9ZW6U3/v+jZTx5ZAf1uugZyAPEFY81CiDKede0+1C7rfiw3aenXVEwcNg
ODSuiiMGdB2KVo7cj5rL6rAVtwNwfh9wSXO7XhG0v728LbamF0HT8LulYJsAzr2kbhIzJeeaqmVV
VLm7v4U+l220waHtzs9EnW7udAP7IVQYZLnF7iKcoDGuXz2o35cqDMDBdR9w+jkJaHIBNZzdNNAX
13B5XlxT2VOKX4hmLOp8UIUEW2/Omf4xyZAVxuAVpYS3Z9GngspEICu9LvuEwy87dYt+xj3HdLnt
EOxHdbkZgid0J4/3F5R5MOt+jzqyCo5PbYZpRdsTFUhvcrluVPGUmN6TN3QDRzT1kvvEzEjZLUuY
rQtenhhzL30I1y+OHW19PTT2gin8Nsr85zQQwkgWSo2YUQ2ITpm2l/BHtZYWnSsPCVgH9U5g0kri
c+upgYvHN3Mnn+RZiBqp0Nj17el5E1HvCBx0ULwRbyRXkzZIi1PRyFfK1cvh5FAW9QScKSiLN92O
Jg0YVKsXzJo44HBHoUdFpz1nDs3buESEpNWPr5PxVKIbr91MgSAuDVCNpQyr84kN04D5UtXSDB3H
l08pSOi4JbHak+tJTJO5/z4pH6Thb+lK8YRDYvaencCnUT6zkitGgT6UhfJ7nApbUIrmhBII0ZQs
VpRFQGo0U2naFM70Jwm8AUx90LlpwU5SRLl7epzh7r6FtWHlnwrDC2+Fa+F2P8koIwwKnZPS7NIG
Sv/uKBZ+4v/TeQRVsHJ+6iXSQYAukNCshlRFdRTPC5j7wqhCx3gsnE0jfAOmSks7X+9/jiD3kfta
nC/YtP87ZDY7Qt5Co1B6F+mYA+FGZmerYG3jbO/TpXcTu5Dfn61GraUYSgf8XsQ/SkhFVt8FGwz1
dXVzenvfY5bt0FukeYWFyoeBA8dhPOMB48O8ZhSvhJqyWswrTAgH2MbWKD6EjLi5D8lWacTZYtEJ
sFsPToKD/3Cpc5ik2B5jrE1FpVtromNEUJhSjQj4cucxaCFyoM+DMCsqEzFGRQl0CPIL3sU2uaJb
9+y6D9bsxFeC0evrsQxsYzcvaJeYbCDsLGMEDKwlxnXqGYhDxcFLybArpxz2ku6Md4uva0vhhT0s
tRKegagvDLYgpOn1DfcyQVTKgLnuKAVcIOYwBDGfxTjO1o5ZZiA1Rz75gcYloRiBdsfCpeE0GsFz
PjZxg4dipQu2H1NBP13XZ0bSQkBKsWZXu+Ls+QFCttIIB9yiAi+l2ErTL10SHH2cLgWbVthYb7pq
H9lGeYm9y+suxwPw1xCDU79Rjt3/qgEA+KTBBS7qbhQzSR4sg7Terc++giKolZY9oUN2Okm1c9vi
WiPHvu8p60gKfr9JVLMGfmRGz/4BZbVtpXgZsSi1QRoQYDU4FCXzGaYS6BOFHF265Dyx9/MfykmU
faXHVG/SVKaoTxD+Co0z3WVYqri8d1ZjN+IqbgpUE+5iS8jdWuDjvvwYp3awK+6eHdrbMRJSwwGy
2P3bkUvJ1o1c6BfFJ21yF580cYkqNijzwzrIs0G1KaI/jp8nPKy7zM7gQgvhKya+PPV4uhoUvph/
/OLQeAWrv166JlkgeTj9/VAnvL/zZ5L9rKXBoK0T71gxkWl4lXrWpB0h3qGnfspDfeex6NzVyr2V
912k7kUzwmHbR72iyhYgozaM7T4RxORoBdJkA1I/+JbWKZUcAj/EizI3WEuUrk9ssxgrXs6OX/IB
uWOlkTicV6DZ89mhgE3K60iwBl0Mv/4129wHWLDdOOlvXyHijJcVKZCWmQLX/u/pbt/tE23x8RSu
TA9C9QEpTSuFr24XQVY+z/BztV37h+aAgoGBvBdp6HVFmIB+oqT9hHrSWJKng0bIvQ0cU6FpJ2eH
MVBmNyHNN03lMq+VvHPJA/Bq2eDqFB35rVxg9FTkrQjaV71bmhJtd+/ALA2KwzldY9U2lZ2S6ny5
zVKs/uEEkjQHy3Lfe1Dvac4pkjGct1QrxJZjcnR7C/fnnCAGAJNM7L/6q+RzPYONXZAE837xsYq+
0bogTrwFU7EN+Jx53KLB2edbqcXnqeOxU/9lmnObQsH4qlFUjNY7K+AfRBNdvZctZ9/iKDYIfRyZ
Z8ATp7KkU5U6ZP0CQIRrZAEPSPkty9BGp41zfqRkMROvJ0qUUO0+7eRAZrD+n4VscJ/lIHen5wY2
jYYO0tYtS/dOMVZ9gLivh5wyWk7orWrjC2jZKrzN1ydeF9xxmHz08XK1+6ygrEittKk5FJA1S4o0
UOFUR0MHhl8aa2BPapEromHr7egEbRbwYTr3WvSJ9A3nq1JVCadgKMVKVnsGhYOM1lqEfPBc8dC3
gahjwlIMLr8vYwibTzktqAYY7PysjBlwKk4w50ql5BTjLUBLg9ChfTsZbWGIv+/O5ZZQtyKc6S+n
vYMpV3sJI4uacUgWCIbf+ZgMZ5z5hKc3LRdkMOoFaCFxfHJE6kkc8sVLTW7OBmSDSuYQBNFUH+X1
XJSGb5yKEGRpL3TEaOH3hFsNcHpTY1vbifHRrQ+p64caEAmi4TFHO5Z10hDlgdv3YpnfFUd3XpQh
2BMDgYi76QuMM5pl6O31WgiR8CLBW9d4z6E80IMs0YwTLhTK+7E8HyfGz513jgvKjkX5ABNdVmOu
cYn4V34T8YVueezXKa8PB728iTsIBvMzCVkHZ0lU6t6x0ZSl7Yxp/BSUqbeXi27kb0dJl03/AORj
y9Q+UkYslFt+CR5HCBCVCyuJr8QC9IXkg22ZLK8BqSwTBUhZXvWnrwvXW/YfB8hwCwka0jzKEJWD
+KJVM7TaNikFXdOfxSeCKITpXdrmZUcdMUBRXjpQZiqlmd7PpivfnCdEcrEW8id+aoklsJkCuUGt
l2vof84uXHyVljX33HscGw36L+JQYgTrOGAeS0iGcu8Ley3OXqZwL5hKS0tJphfHaTCp7pDGq18r
iqagQPX5Qtu3KwR7GimyE4SHDIpNj0Qbu7Gf63JNKtm/z8R0RLGT8PHay+7BPS9pcZT0s35IzQQR
LH6jtn9pgDzVSb5WC+rJBsAW0m3j6I0lQ1xuT1xep7M+TPFKyo/AdQEMZp63kmH1jcVL5cdxVaSk
k/Mzuo6GwrEwRGkZjgrALeYRuVZwlA+yLKwnKyQ0J0tyqbYksKzaW0GiQlrwo/PD2BH8qKsTri3t
gvK3SSUjxMmCv0wQj/u88/kC4IS4HNS+iprz8o+nUIutr1q42jnQcUeIGbteRHlFl7ubBrvUngvQ
0qvLIjhVgQa4khy/Xf4wrJET4xRSOXeIFiJ+AhVNPtVzr57JbRNSyNWFGzb9WKdV3WaX3UF1PQ3G
N3BP7FoLqVaNNVPLNfdotpWt2l/UOuC8UjtWaI3z7BfhObYxf/ApxwWyP3dwvPN1ut0sNWj1KefE
sAxbGz/i1qBGBckApMYcywFj7F73q76g4WR1RA4g8hs0Ym+BWDByuxqv+I/eSkW5YnSt/iL3JbZq
jd0NgRRT3UC63WVFv8AEtskeDzj9RbV5rzZ272dmPTFWGdZhoWueTkhgPWAN06YLZq5phvnhsD3h
m93gfI8MMnDkgffBDyVoLZz7APy/Wbp4NRvKStV1Kek8ugIm2ODmB1GQDdeRmNEmp4jKVy3YlawA
zbCGo0n/AJrgR1CoKNOoJpvetkHuIb2aBNvgoHEjGJJyd3Z2k5lghhLinMC5m3iEFZsrlBKhhea7
F463Nw4omECu0d9QDfUEDeXOey38dtvx7gfvVrMbATtUk7PXDPHRWjle2KbZIOANJi/m5k+7j87H
+4y/c+om27NEkL6UqjwKRkcT7JQR0INX9gVLcKQUnrXirkTX7VnlpVUJjLFfFbvM9eMqMj/wUpYV
gO7gzEH0tYtNMvTPD1/Xfw9wqr96275WLGDNm99laXaXobZPQWC5NwOFmGBPre3U8VXAm2NWpG2a
ea4ww444QXIrDFkuNRM+ru3BiAYKsMIJnH2OYjqGVB+5XP0lY0yZjVOKIcGwxo7djyLcpcrn6ldq
gejQ11+0QhdXpIFC3fB+MdlxOe3Pyx4KRekupsK19TLbJ2HG0AZl8GVfqjIpxAfed4x58qKqnnER
03tWQuKpslP7DjyJWkp9XcII+byADycBjKrch8OY6FtgG4O23OgUs6s2zb17aCHz1ZwHvdZ/IIjR
2EWzHi1u2VqhcWcjcCB7eo6ob/tcVQhmaTrREteh+l363BL1lHjJTad0Lh5+GfHI5LD2greoYV9l
eU3dgkS/Kd08Itr36d6bFhWfpOklrBjWPOQ0IkH+C45lb3gBHtIlV4tM/BmMQV91bpY4SiMn1F2i
E7iiKIEwZbd+T2fMqEJnsU2+oKZp8TTr5hqWiENsZW1VJkJRbmXL12ezh8IIcS2ZMfi+DR22YXSL
ZjreC1yPBR9abisXwei/LvjDWvLSAqMxQdxIyVE6gqo6zU30ZNWtwd/lHZ8IfgvjG2OFd5aC3koH
cZGPya25w3Ihy65HTQHssGTPfGqD5TIIuyi5y7kAOMxsgKRcw94nXt4tboVRMb83OiiQRDTR0Gnu
AgUsVgUwybx7evvuL55Ycj1e6KP/w20JRgItPmafpoSsiI0unTJUX7Hw9ftbm7XMV3IDLH4PSL3w
jC2TNwOs09xJhjiyb4s0HsTOcM4H6SfTfHxRKLahQjxVNLMbbz4AUS/d4Rl4o6cHO52TgP4eP+3P
xv6eXgZ18aiz4YDXSoPN7Fyv+z9GK/sOq1O+8XF+LSyyABcL83tJz/KM09xVCX2Tf9D4lcfgL40a
TNuOI3Lk/BzQOvuQ9yt/OwMD9w2mC8QukfTL7Ejpm/NEPh6yKrdKlfXN9BYCcemcd00YDIr7byFl
3TzXHz5y1uKe/tS3i+97I0Rf12weITigzZ8Pm5XEJEn9wFT11FMQ4oX4SA2xw7XjIrhp3VcjgEiJ
KOx4zXWaoNTadmFBbNNlqgShhOgzlU4hTxoWITflSmrOEpTR9B2ew/h9oxKVo5r/ycSs5FK12Lr6
8r7TBCtGAkDPmsqh/yptQ8OrIitzSupz/1+d+Pjbw3q7H9KEHNHFW3rz8ydnUunmHnKZiNXuSUaI
C+UL+Yv2yPdKXjuipPC9GkCtWwwEmo0+vjRw7wRP+f/1g1HYQaSUpkbw6WPbR413fPajTb+tjxMS
xjeI62whUQfKV/HedoYpq/1D5ntNEjQDxFO5ZtchU1VYeCR4sw83TvEW7Al4QQdGR0GR14d6gitM
bexaiHAGiqgY/sfz/V+teOo67VcSmn8hGDPP1wojOGTzeUoz6nNs0iEPZzQJq2gQNEaHhY7tFpMg
cybEN4ZhPvKovdxf/4w+GdC9iNZcWSDzQbXtdXjtFoe0kXdlRSI9fN6cBxXgfTh3xaBsN82mf0JS
gfEh0lfoFO7RAWX7CFSeCjBLfrmdRIXKDXKKIPSVGvXSE34t5QOXpG+PJX6YLgoQjPF5R/iG6JTs
934Oy4m0yA0AFx7i442XDS8DVs6prTD6HEKPKuVD82VyAZGOX8zLVeyJ3sd8H3Yzl/ib+K5KSvA6
17hQI3kyL8qxE/yBT397W+MUKKJYaIJfadkLpLAgvLdz6vsr+Hrim/6lxfRrb8aEtz2OIxZFTb3F
t8zlcURRt3fzgmNQUmYp4pKLU6Cbr7UDEmuVd2PX4UdjGM3ow5MCaaM0cEHJEYHexF3Q+gfGB65K
ZmrfcETtJPN1TG+GGu6ko8FDZ5NqkCWxvCDPv9O1chnaYaBF8wQPuo0YCgZbHrSVRqfFJKNmg0pa
gMV+TEA9TztFSNFlGxhj1zDdU3lkIoHnZ6U5+Cq0A2FbP+0vquwhthP6SRsgy8qrrJ6gQDAnYOOt
W9RjHcyxvVkSzSMsZEt6q+1WDElAtwR9dWZ9eozWI/M03L/cUwHzOIbK3XZ3mAzDNQ2ldHRiRuFy
dB/RANavvSA7WlqfU7e103HgMHAXhQUzA5wqS6henOVb5/pbbX6U5vGCrx0IOJe1KH/VYtHzOPSg
ZQ4YEMFDS5c4Glzc7iRwz9nuAvOiaXw6jcp2gTJgoL/qkYI6h4Dg5VE8Dx58jjSn9G2rIN1b/JAg
KPEoEjzH2Y8Ga6mzd5OS/nddD3blAgxqt2o629/YsI4GyKEJDg4RAoM/sSGO0pdCYMMAgATuQz6R
3oJ/aOvavY9HOfAcIVUlFB9U51rlj0+rHNvJYlYcsexZRuTzZsUvm0XKjQ6mIqtqZLX3CnWEoNZR
q6jws5k4ZMEVZXxZO2yLtkMhDfqKT9wWEzFtnOQcISEUDqVK2TImrv5OlXqoFMqJJvIJ0eMp5BcD
cSouQesUFy6+Vlklzy2G8LB9hJNQ16uJCaN5e7bTcxU/YIuUBxRM24WTKPaY6xtKwGTZc/OWFn63
wxDCek+yojNRXJ6BVhe0k6Lb3wRXUyvNPbI1dko5H5XBRM19odLfssDrV0P0ek0YL1v4SJYTwnkk
z4+AOIJHpeOTnl/MAWSDMLl61r+sevLwJzWHljENcR/Gb5rwZeR2H5jAE59g8RD4UoO3lH8L7rJX
ew/twkMgEA+Vh/FLMGiiMUxIqgzydICbVbT1P2ZsPIZuGXuGk8Mt9CoTIucoKYUeovQcnkpxIMu+
cisZaJUJDO8BdLKy+MqAvJriOf0fpyHxdvBo/+JlacEB0auLaJqm7f/wr1xTRk0FzBgCqa8z0qvD
gTVLdc0tasZJTnE5IvZH+H/vV7B6WTOKpFYGg4DvqSX7CS/DIb2NalWpbZRio4PE/NXLQ0GsXiop
QxtY5YhqPYXH9PHalaYtQ2FN0goJ7OeC7oAS14w5P5hAOkmKoeJ9rszHhb+sLrRY6R9OP3yiDI+T
T13jG4CMX//EphCCDUWCdFwmGjALNvqmH56vW0R0WEKGkK17EYm8Js/F4Nes5DnhtFBvtaqNvFFb
vaI5KxrbuwWQLzoVdMMoRV4/n/qHj+YonaEwtOTTeBZnsDewXMyW6fweOcjCynhwRMtK7XyxBtYF
NDyltzUe+BOThmcgQtOfki/Yvcv1qNSTmBIReGgMMsoOh4qn5ZwOOdNBhXBwM2a7eYxEv27dCH5i
1dFTWGg7+PPa7r//RLbx/299IUb7GDifoAxbkbfYzTP6OqRmpkrEO8tXaZZvuvq0jHyh2R0ssijg
m5f9sD7HOK5pbwTJi8w44GlviKEaf6nZxcLhSwPpMe1ShT1RzPzM5L1OIZrF10JoDHtyCYu0HE4L
L6aME1RUYTBSMTX6to0TV/unKJLTwev15c6oUdILQGdRQR3veI7wdBffjIrqaJcqjrf8UWfVMyR3
YyPbhYT56IHS/Zv+1VTaCfYULtdoPGo4P0hzKjnyfOASNnCk1keFaFrtEo8tpbnZ6HS+FSdbpxWA
WYiR6gueT9IFMnEzQXO9NDvCjoDDziVokqJZoP741LaqNBkjMjvR7zbkG1gzRrU2PCyPbXoAAd3M
h+qDRWkt8qWY2StU/Z4YZzvdjGt5qm55uHbbokJvpEcb+7OJlRNTfYzHVAlpS1GyPQlv5b2JeQfE
bKaOo5VHylm8Qsxb3CT+AsOCoQDQ+CVX4O/3Wj6xAlfLqwD+lyYc3ei9SWSPLMvzxaraVberNoMU
kdL0uUjGWgvCs4iF7jDLNynpaCrsm8EFPjkqGac1K6AYbfULdhJvvgkA9Zz1juSMMSxlqXzvhEPi
4oeybrmAYolYHd8T4cHpi85oYCfbGvP9rqU3AvEEt7T0doQLNQWp5GbURXk16fZvCDL9a0/vwNtE
yabbxapujZO3vqbxg0wIBdmLKirzCLOXMY2ZaJC9yUAKdgHRiw6ui+a3sofefCWy37qqrXTlPNEd
TOtVFFgh9x4/Nfb966QkH8CJgd19uLKG9xM2cY3lsU+fua4Qqcjh+iK7t9LYDvEhUW9EY7XaV7ha
CLnD73T1Ova/tXOCTAxZIrJ7ZYseqcioIxJoXKyC3wKOyDekwCoNfL4pXA4J1VVWu7nahRhH4ESq
sEIcbhi6hY6evYDOjSyQyIJv2yAczclHDWD4jXnEFWNYWz3eqIC3sI0s6IoVyAh8NTjkKi7e6bs7
44iGBAUX+jrhnKwWwj2LCXimeX6Ynxul2+EnyDl0LYJ4GWjyZ+vJnfTgn3ukQrZqaFUNWKU17roG
59FW98CzXT1z/8W+BZPQe5QU8QqyV2BK+3g6BykJ10STiyXBaB/UTUl6xWpv/+WXk2vgYpRzoSYT
pFEWBWChCR1uv26X/yVl2P3HBiBz44CK3pu8WCoTo4qmL6IVM6Ob3NufMzOjLJ8ES6RR5d1HTsbi
ESCB8xV8xaKLJyGDfYwwnLI6AvYRJvihWc0GeFQR1WZBlbm44jyBUOcFgxfgIlky/bStf/r8DlzS
B/S1YfX/iBqweB21J7/E5/p9o0N4jQ3O3i16NVJ7cQ3yT4mphNSiKF/icPIVOzJbwxaoI5b+bJki
couqyO5mPowuoBJ/VFpKBRXZqBxouheCDjlzIGf/P6MTuSs05rVKEFHy6P1w9toEKsxwVBbllVc2
XIo2GYskeXtVweDfjY/V/Z3hDb/iCvzH0SrBHLQmmoa/3vsuxvDqcs6FpcZpQopROV5mhz5YB2u2
URVDQ8lN6Z7JxvybJJxe6dDBHfzVMfxw03ELUwbALf2TdFz+DjryJQeBq/GlTjGcDuE5nP24BzpM
+tk8ZDW5iBzDZbsAI8OYMtR9q5Zil+am97aDQ0rgYeRG3Yav88oHGZUmkCGdaIaRPj7kgvVT0D4M
NQnlNUHP2uzRGPOhQroTGYopp5w+c2qiNSPfq05IM+pUJuA7nY4hZ9siyofR/McFUcNt2mM5vjiX
b/f6TmEqDOY3ZA2E2ByFnnyQ977fqquko7fUSNw4yo0S6ruDTKqHcDEP/P3F061rvnJKZ88Dlv8J
UqdLzJcAK1kRArA6gJtGK8dEVOKtj20eryLja0Xe5plWZ2Oh4WctWKoZ81ssPrwQNpjf7E/JxqwF
qIxQiRdBp7sOwdm1T4nv7xdgy81skHaAdKWKepwl4XaWhusefVN8RYV4UPf16gg0xitSM20NHHIE
kuSKVoPs1VBTz0Ap68mZI1aYltEfbruLTHeHczGpn5rPIITYdwJq1lePoHhNm/Zz+s75IESeH754
56Kj+5AWa+nL6/obOP648xDUiLIDpZh4K8WAD022BSyq249fos1JxHC/amQqwgecN8SoWP0o55ZB
7q3/lbX/0RQEZjYJP5dZPWA8kBwL+X7ABAD9cJgPXo0DhD5B6QgIieykfKE3y91Xbj7auzeQmbdH
0hZpEYpqkRfZHhiLSdgRtPAtiX9TmO2ID4KpoVrBlRO/DUS9lWKEwBDlojXrMIoRDty+XTNILEfP
b1zYd7YxNgc9YDqOaQQV4xKiVF74C2YAcxMGOA39ePPfuIlt/EQLfiNnlF9bmXKM+qfy5EJQDLbO
nmd1rHv4w/HReOepeiKoT5lC2tEh6WtJfMXDOngwk+qDCvEeOfAihcJyiN++4GMVPuNYo3Qs0eus
wN0c82uSj4Fwp+dV2aUBlUKBGr9iiztjnMK3Ww+C3JUL/8UmINXnYHTIH4F7QmWsm14o5WZDNY9L
UdjEcKyNXROSV+CEo4c3HJqdPzf0s+ErOLUa4lpFGwGAj++bm6BPC1P8+0/V9JoXNXP4NtPcKB50
DyIvpgevbXBHRqkBrwEnBcyMqxSDPLWvFRz2e/2VjLUakbXByViZy0pvRebBpNl992fIXUkIpRg5
/KzF4Wmqdn0RUoo1kg3VOsrAfPHbkc4zSw3vu2lTOuMSPc2IlXQo6SeQDMfv93RBR2a7vIrO200D
8E6de6S2WRVI3YeQyaUNOKBpEaeOwT5UkT7gxHLtkB5rItN8Sbb8CUsywZnen19uB/zojbiZvrQ2
4RpkwcU69yvEls3/5iOukqkopRCD6KrhjNKJx9mjap7vV7vC8d9Ki6H584ZPTLZtwnu03mnhC68t
F4zXKVX4FqVauw9qqNDzPXP25R+vFwsKdSVrruDedvfFUN72kdi1+oVPGegr83S3Gtk/Y+siPtq8
KKKi1rQLe9L+XJu5uDr6gor0D+QJmenY5rNA1/fAOCOCUtmiX5JrVXUGGgAw8iPv0U5Hdh6uB5N/
lmdHDeLzdM2fgems7F1LBWq28PbtKCA4Fiy9oFrugp641bijSGf/VaaUeoPdn0ltdcljMpjMple2
YW3vdt/kNIklfzb6vEfGq5tu56eKpgxuNDoDKEyCgYO+uyhbJr/I/KettXqmu5MvXdk/IXzdY/ZS
UE295tXHisLhQmwn7HP8w3g7uVlSwlhXpOMpgxMLqTRRoHL/3AdzCKdlEBo/GmnaPnYP6OgmyUUz
5z/5TNoQb3q4DzFb1m61KcJ8mrcSUi5+h8U7BmwEZwwicd+OlxMYyBLmWfD2cZIeWgR4SzFjx0vL
GyR4j00Pyhh3+xwL8MBqHS9mJ2crgvAgdNbxld/lJAzcw7mkO9wvveUZsIhSh3JNFy/DTDQhzA2h
stySmq49HIb21wj/bi6duXbJ8QJHJSdwgkOM8bbAAC8R9DMMzbIF8i34DF0Sp3ZsAnsZQEd9PXA0
pgwTxj8ucJlLTAi3XwzGILv7Q5ItHO8BnHdflF3J+jD/7pR032KOBW2LtSLd0H8scOzllZiY1OTr
33Jz/62WWQYrslbYwywbuMiH9gfj2WhxryowJ+G4BES3Ux2Ac3mf06osLxQSZxjB4wwbP2sKWGXK
N6XYF4fl71xP97CjEt3nP0oFwn2jDZ8dSkyaKWnZZJaZrRKFfCzGJDd1D93onkQ95atdng5vKIYe
TE4GAj8VwKdHvPWFfEZKQmjq3pOFNiRPdlBfiDctL+vlhsEZIzACwr6WW0D1c1C6yVNACE/hGh2/
2A2KpPFJRRqsmgyVgJGtkFw9twmJU+reYPnMc9V7dvev/vO7rGvkowMhMMzqbuoFkUb3R10JtKoa
HhW1lFVNBKy0xEj3EBOQ+PHtksyJUL8cT0ucn1TXvQRtzhPD51yZ+dLic5iUSl9rxkSyAO2tN+Dp
oMZSXRMy90TAehZ10J86OSsOLKcecdoejBtMM0C6qNDeWR2BPfPTYn5Go7TKkLcMttvnEVhk3Pxt
RmwkF7ml6X9u1ReNn6wUW4PZIGI8cYy3Gh4uInhSurHnuVXAsWzJCyAgkYUe7IXEdfmbc9OnjTGJ
ysPntthH6Z2HX/KfcBc6Wm6g7Pnwn1SMov5f/fuarWQjeQXYdqgnY+4WPozJYnGQNgn8KT9lLxoX
KPt+TCIBdF0yMQIsEBrDx2FqzhRJAJOKPw4DeO3CxJxWbxrt0Kfqqv9z8ZDWPTBj/v5O3MA5SbIr
mHDJX0PfNAwNIovgdG3GJbp6+iCLMw2C5bvfcOKUcPuX8tmhFh07L04SP43JIKVPShrGtsY+a10R
uN20krMHp36LJagueW/s1ycD6ZIvFx27VtLclbbtsD0zjuclpQgKVMzZf/j6A04/hUI/IH0U1KVm
3CI+UfFlhfAKAKaAQKgd5mhQT0fblAO+PnDVVGpCAZ3XiXep8j24V97rNun6S8VtnIPqXRZhjQEz
uHa/QZs3HsznA2oOOsg2Q1tqJyl6BwV1Fz51Q2CImb7mxtgsLGdQObJz4l1gxYazaeySrrumYiOQ
8cOfuwRmjtyZuOpFJE9TlnnhpWQeGwEhsxqOtTWZGZ6s9CMrGdbt9+bOUkXkIpWzpg0sNMsVu9/h
QxZFgC4e7W2k8zLThYeamSM6Hmk+bYX5IPbq+syfeyFnGVUcI3ypCdy95Y2OPsD+BsFWEqKkQl/G
RTkP3gYpqljnokRIWXCA71teUnqj2luyqMkBNJdB4hIivghTrA6DDQLFzYnn2PYhInwk9SSuSZIZ
ghjxCvHyMYy2a/B1rOQquoD6uDiM7o0GeBylAv3YYPe86yFjnBoNwNH2X+8ki/WCBHoEC8ywoK7F
OTKs+XtgrPKIHZZA3a4hRAzrkdCbeHBO6mKD5vv+ZDvidjNHnEdz6ddYqyHCSsSjYU5fiweMoS2F
3SxUnqpdsSUQqh+nbjwaSteWymoaiLyPw3mE2WpZmvYfy/B3jb/ZV0hVRSQkbsGMRQBRNL54/HiG
bBEsmqDyG/l5LqveeY6QhK8tLHokZQkpDA0l/sjP+fRSgTinjlJJWwJM47xnwrhQDh4TndZbum4q
LvXuXw0VNM3Nv/E6Ml1UF7bOHuoG3bGO5Ii4kYRS8J6rs6IYTkuGqEtFaWBLVF1VlhUReE4pBZkw
6P46ZyS1Y1YyMzIWz9jKfXsjEezb6iH/cKLJVcFPd+BJyZu/j1Pi3zamMLef2WXp7u5zZv9cd0Nr
nW0vQAueOPZ5kwXxbukQslvT2F+Hc1YjG3hBbY5qiW/qmwZg2pStuHZbfTjK7naT4+lLC6oEipCH
qhe9JA/kuIPAsJFlrnE10DwZ2++A+vLJHs7f3rUo38eCgBRjjSSWeg+PtkYRnary4ff3yoyXca28
RkUkFuftQjF2jYZyEx5j0a6ic4IiSaqeFZOuM8yaR3U6PFTDeG33qvFKoKEOtMc+HAJ02YuGIg2q
eQVJaYr+AJ2Bfy3NCcUoynAxgTSokkMNLOryEMIZp8gm0nuXFAQK1XaV2rws5ybglHMXYNNDmK22
l+9Q5CndXae5NuTW/BTQTIFggqdMu0r7praSziZpazMC1476/+GDCJto4sIFUyIzL68CIpFnxDTI
zA2/gL8aotIMWBlzrcxXkGRSV5NHMgGjVq312apQghyh0iwBf27xOCkkR2pZAHfLDpu8BkPZrJSD
a9F4o3Ye64L800WAJllz86dLBYqvjGpND0uSEGcvXRuW5PQO9JU8EjTk+kZaSMbnWI1UAx8YjL2v
uQ1LSyNJktuOSfmdtDE8pV32A196IzJVgpns9UTinjpYh+GAJrQ59Dps8MMJvYL/YpJwsoki1bz/
HfrnhmntFdneH7bFxg/Qupw5sFo65nQoXfnlsYBraJe26WzYOOAOIR5mrYlqLNWcKSe22qtGVkvF
M2K/5yi0qw0UcMP0dT3q2zGfGXFq+YUNhvn1eDGaBxnbjdW4r4V90WxdAAWjMTzeTfihaTCSHjE3
JBWbwTmOjHLKPWZz12kC9Ls4K+sjB1FcVc5uWzK58BGd2Gaw9M5kJGQj/6sWmuNs1OKEej+dYfL9
LFgQ+PGTSiex46kja9pkeZDvvFRKhUlUm5ViW8pDWrP1Acv3dalbV8flsOGVKOJ3h7GpIjC0Ek6o
C514+BKoPaljn1AwZP6uSUQZmsEGBjeX34+/O8N3+R8dWqg5gbAbdN3CQdjEcrIwC3JCj4e3Q/FO
WOYPK7GyjrksVZDggfinbNo7dvb0RTsAqZ2aUZIhnNGVI5Fks3RVRmITcpsp98aMCpGsnFNeQel/
Kk/ql34AaIrMfUFTHos9PeYQO8uwBD34dR2ISdl0vH5oUv7zKgeiX/FhQzT7nos0AoZNtQRxvDsJ
o00kO6NWnGLHkayL/yegM/xXoKH4gi1PRIpnz6ZlPyKkK+yEAUKjSpPDHzvRPgZr0j8uPxG5wFpi
jg545+lappxcOkEVDdx4gJutgkkTXwXaQYGOkL0e1FSqfjqr+6mrtSGq3BXLLG/maj/wHlxfjZsn
VY7j6fhpLxecqTKjYcE7wzFLOH/jzs8JKWFeO5t0ssQP3dMcEYIi6q57dIWTh8ArmyqdfQMF6cIO
zzUZhI6SW/TEep5u8UDAcJk0u1MYa13lf82ydX+/LV1Z67FFu1hXpAmryCRfEz2Yk6zUsj8SJ6Xy
KEpQYgjfK32qs8XlMwDo+o4glOB6UWCauP4uckMFuNtWnOXWlb+mzxoxNkjwI2Q3k8DGkohOkaAQ
UBmlwqxQNxDhklXz/Ks5S1uW7kG9Op2S+kf4aE7NHXSeDSfct5vVBfXZ4zusOzq5awOMr1AmY3Cr
4XOZDhlVxj/J1lmSHO3YqUi13k0uRw4fh19dnmteM3BGwxprmkUjnyNpp+vk8JJV46Eg5VRkBCsL
eytcPyxyfZaZMRPopUNp6BBJrKR+VUnCkadvm4NWBpuARBegrXLRNIhSF7WcIoYLKOdE6j3hbaHb
ggPlLCNWbDF8P15pM3FdpPHqxBX1sOFr7uH0ilaEIycTGxP3U/99c0eEJMlgouxcohW5A2IU3B/O
3OI0x9/ujjwp1SWkbqNAs3fLhrgrCigbKh3c0cdz/jvCa0b60lem61kKWVfSABR/M38BIW4xzL69
kEShI2+RMnlEAzITJIBq8kN/ygI55EOS6k330xMw/L2vh/krra0QcxUcpV6TPFj1swjKc+JBWq7F
OIevBfvK054yaiO5KPh2TuZeFxoybR0XsiYrsL0tgmzK7kzpkqNX87DhzhqujZvIA580aB6HZr2Z
Dg38ytXfMi4ZnKv0yh3fCaJDdhESqzvoI/UzQYbv/xxS0Lqod1VCRgPjPjHRmLQldUkY36CJAVtF
FUaJcXZQpYS4Hmr4gNFQIEiKeAbnI8d0JHI2EnAPf81k9H0VfH5Q61Yp7Ylw5hR0mK7drQzXMo+N
MkZCb+vftNvq/DBVnasc8l3ctY8ywAbrYXWZXOn5kfvOydHCFgCyzVm1GYYcXDQEisXPsEFC8qVj
xKkQ9GnxfLBPNCO2ed5yjYXVibqHiyZXiNSN67FrMFpphbxZyqN4oAZaVFKuufDgHp237PLKgjwV
AboIU1tZn+7U2G/457Vmo7BredtUPMHSGEtAwdny06EN1BXGlsnhaW4BIs0nPb+8ZXK2AClTW5+j
eUSiKI2uhlqfaa498betagnxz57SIIiWAOj+dtwEAQKOMRGZtwYQrP8THNYLy9c4Jm6VbZgqSfO8
/OU3GpQq2Qke4sy5eAbC/PTn8dVHGThGx0psGBMKDzdZ8S1wzF/C0nZ66aAN00fjVsl4fZSJ6nCI
75IghweHVvJPzvUxDQaIFr+N7cHLLXO50CuiZY2Xxbn0mRqlx3bQbSLMUC2rmFqf1qfljoAtvr0B
51XPX/fFuJo9QzV4fiwyHHEbzKhJDUfAD37xr9fKsRoKJTrm7mCR3MsArqytlJ6XlJazDnZOIp6G
LgpBZBUufx2c7qbVF0K/KzwTfSFDdNKIxQhAk5blyexVf8xDMjlORKhH4bJjfh9jDj1hrfI21b0K
+ky/h1SzRx2GuEeVajK5GafxncXkSw6lRq5sB+WreWyrzL8CLJB+IjbFAeZXI9KpQxBUEkYRA+zk
zt+9cVwX6kepQqVGo8UpKvnZzfGNDcpkiNSfne7Hc3fHDbRH9X0smY9u+Mw7UkZ/HSwqU4wqzMu6
otvtFa1jPAlSBFVnFegPdXKn0qzLx50EPgJNwclGytkqJ2Exwq4v4uOIbdwmlNuvE8e4NDmZJ9vm
aNHzMAdX3DqFdFD+rPSGc7isTZZE+dof7zmH/cFd3in2U3Ig61Iytja9f/514Ss6Ie0rpFRRAd8R
TJv4AjRY6g8x2jSkbw5wzCgVWVKDU0Ko4HY0hYKAPV4sMi61b6PUkgzbEnEGcji/ZsWB+55WADp4
tgU7jo4jpVIIswzBixwNWCgbhu/otCC8WhdPGQR8jnQLwY+DnerDUZf6idolFjIssiz/8EAzsjd+
16AeT7oKDCOE7dCVaBORczJftBpy1iQVy8Mzz0fKJURHNOTkzKXcPxIQzVKxFnRV/qVzsApWDklZ
2LaMnusA42jqe81TH60p2l+0PyppVZlDhurldt7+geGpFc4pQPsRrBrajtd0hXDkOxDUtMGu9VA/
euCj4Ci0vcPAj+Z4+NXooqqt9R809MiQBNX8k7hJgqruwaddOc4quK1d24hbnCehXHxpLUVPGwvx
ZWEAdY6viBxoXThdLtSVbZex5cpnZYV2hC7Dk/PmCCUfGT0Y73GQF9ya5o0/VmwwRORubynGzNzS
enaiH1iNkyO1KDXDaF5+Oe9oQdJIjCJbtf4/Es9xuknn6UwrHICy3CsUNfua0W2PjcD9fASjig2F
QHLqb6meAixRm3u4FWvrOEQ1IHapNy6uhp7YuNOjxjbXfzBHXhKS/iLGTTMuPAqMYYJ7Y9eGzjcX
7CoNMlmyVJOilyR8rtvIo4TgpZ4gUrP8ym+Uss5T3l3wlcAD7MuEPebqtYbHsoKCpq3/sN3Odrrg
bQtg4MdBhjWPI18dIGxGTj3vvwyupaB3fMj7eOdKCFEntb/bVf6g04CmnUcLwZ2TDPnhNfW3RJAX
dP+9p4CTiytcGP1vf0vuQ2miIbKx0fapqVCipNtJmb4Jyy6ucEzgEH14bOmjCISk2DpcueMYQGsr
MwNmv7+Ct49GaxRnrnLxd1OOWYigv3vpdcdHcd/k1d5pa/4w9Kjb9JzBemfWyOFwFLCAeNr92BaB
VZuJD2aDYQpIA0laJ03fLn/iqyNsidzhdmp8tTfm4vFlTSOZtQ56RdRqilZjyfapWF3D7ib/gOVU
Z6I5c9hnC2YGTdzw0Zf6PTDSuxjDuvfzyHOaas5qx6Vm9soJC31nrD1PIdExzYRLmMkBn8+d5/Rg
FerIPbNsM/lA3/8jxDAOEkQbxdxmAdS8zb/c8fypw6NfyogQ1Vj6XLFyU+JaRNJCvPnfmI272mcC
QnHDgPTuG7IJwdu7HAils8A9GuYriaZ190lYbjsdxxX4dQfILlkSMH4RxsbQ52ImCSzFGU9dVqwO
7dUOh113Mzw9y6Z6nH4q0bd/q0/kVEPJGcHMujAaVpWQYUAhA24EFjDqxDh3M0nldpeaXBdon2aK
lr9liC/KE3sUznYHV3AbJTwzBqRs2tWlsfhfwZ/nxNhEA2sc6owzg4k/Cs85nESVdUsGGAWbo3Bm
5RJeAL2EOsoFZ4mtAFcxP/gx0YFaQRAREOkIua0bhSzzcW/w86y6Wvb3RQXukVaGiODDGEuPky7T
cT1GeeSmWcLMVtbY/oIyPUzauwzJY3oNbRpIOPkWdilXiqKYov+ZH7TZwcDrvej5gLO+PKO8DJJA
lARw4wlnZlzSH1QYHtX7HuJxu4/ueeWWQ+Nw94qi3e+UDSYae44BIC5BVG2MWcy8ekMyBWmlDn3t
9ksyp1CS5+wD9KNG3TANnadNcExtdHRfHj9KjcPPNFdkIb8na9Bd/BWc9LTnfBYKWC/gjT8Nek9j
R8t9p4nO8PC1GhylkZJJylE39zPTNks9H661i4sTJ7sHfV+wa18vA9qxenIYAyz7lGIrWA87Xtrg
OepITcEijC1JmmoudFa9nI8dLJCCAQB0Pwn0n7dmsy0NE17ulgAnpRZhLTxbDFOVynKndLgQsse8
kcaT94s1M3sbcxE+BcNR1nJqkAj2kHiYv+66/WKGk6fBQ4R332K4mLoEDoKBFJtYbIrQCcvMooPa
SQAm9p3j88hckz6oByLHytdUtzkR/NPthw/Csdn2qFjj8SaScdPhgFNyDeq5BDpvzXht7iSPumSE
l6Uom4TWI46iUSfRONicblI1rYwT758cqxRDygRyeD2fotuifKIXYwNxDZH+uNwlNR5hmlwTJ6Sy
0W2976e+zWYSUYlCB3pkY9IbQpcjNqOwi0rUMVQVzYqGAQ12BlfDTdEJGzKDHzE2xEFZjXb9+PMh
ej97lqfn1kfliFSk6NjaxO3oGUkeDakBUIslU4WFDBYM8oUt7a7JrP/CX73mUzDYCOv9ImrextfS
sJ8pwTEoxx2PSi0/PyH3cT9jgoBJi+xAygwhJ972ZpDEallq79hp7raNRkwShh3ZlGmzA7U8Ybyv
ZatSFytZYvt73ukIo7KbNdI+Oaw/MYbF5iGZfElqds96hmpGt9KywvLm+X6fuU0QDwJsBjTb+ShI
MtnUdyFc5qYJ13fk2zsAIINksirPglFJFjpkz782CytOF2q9sRmYF1mfAMR1U1MkSLPl/lx45V0n
FjGR6iN8z9+Htk4HnfXz2SSo/q1Pkc1HS0MQdFT/thdAMZCYNq2Dwog6nWV79mPpOGMbUhkcr7Qq
wc0YCqsHkAYmI8SnpU7LijWDulI8Z2QEdVVrd/ub55PpCIB8Crm/zU2pMd3SH0nLa8AhHCyUdXdQ
IYw1eXYpA4vG91j9yrAnsd624DVeDuUGCgyjp0C6qMCkx0U8SCPtlf/4qUgeeG1SjiFVDlSzLZZQ
MBsk8JuAIajl8vYCxhdFa9sYKGGNCucGYVfwbclbaI7oSDHyB4OPuHgk59VI9SQ+SOYkiDT9FIEp
NPP7Uw8vfdqgF8CgdUfQrgHa2wwn2To8mL707FzPXDJf56gAkeH1Sv4JI8F0IxvIQeBOu9nIclzV
mhLY9JIVaTPJSSKF/z4DWzOFYbpoO7xg1Tc9MzNWN9RpBTTpwy/bVEt24VskQ+jB8PzRULE5pS8z
umWSb9Qwvo2PHpPJzSX2fbcaV0D/8w85Eh0koprfKg97swHhiKN5tXi4I2Zcf960nm7ag1w3kHqL
GKDrhWMVeuqe/w2yLChY3iv0b6fZkS9ULPPPWedRQgfP36yYYKFzu8KIdvSW/Y1VrvCXAVnSRX1y
Z///3+b+KlxqnjMPLP894NAFXV93I9r1bcyjxg8wmQYKWcZnEfB5bvxPR0PJlOleRvldSYQlr3Ad
DPxpiDu3ATYVidtvfpnJVYBwFefvo3ygycHAK9ubIBvhM8CAG1ZeC12Xouaj6WCBFLeuNLCytcAg
vF8KQyXKZk8VamOwnUITja+NS5FIkWgg/VdzoPkr3kTO+lfrQma/waX+3jCOXSviXruKu+Wziagh
LqxS21/Ywoii8BJj08/PtVKxgFaIWgtWO7gh4q/MpjPkbiuGtFMLO7Gp7wshCinbR+R/7HfwAzNf
HK1XRcZNJ7LyZ/7ibG/xnh4x8zlphmPRuGl6YAklcsCSIcUdNrvob1zGeA+CVkEo9Zak2hrxeJsY
GeR2XbR+IdrG5aZHXI6B7ZC9FxVMn8JOyGilX9udNF0z3LDDM4GSZNf3FqmPCizNnAk6MzgHvyyn
z2n37P5qw944mKft+H0FY5hk/YHHas1OWI+63VDkFzupDHTR/JGhC6kd2hyPXGp/PMdVE6SbBm+6
1sp3Ia1FSDTci0coECYFURNp/1fcz6ie1Dcp/jb+lItmm9I0s8W4nwAQ0ASehjqRnQDa0evm2mE3
onZVwuGZSunyDnjh+jsEqj5Dv1yNFIXGRJ3veONC6NTGH+TUqxKPlcQs/aZ6a4m/+eQ6b/QNskDl
eYQV9Rrz6/5uAVc4bOGWswmqV4roZEpCe3TbWaGM/IfsGTAN0n30X2Y55m5wimamo6C7zcNFt229
5zs7mCYAWKMjJ7ubC/JzpATrjS/j38wHTdHocksFjKXpVUkw/9teVUT0W+uefro2O+qfiK85sxBH
LMYpZfNSJo/dR5E9iUxOA4QG8HGqlC8GlU7hv3f1eXEFscKjivBJLHsWJSA8e4QmsJOJBYMuNdZG
PLyKIOqlQEw715AIenXzcDQnhgW02adoMSngljWZA1QL5oCOPEWgdisMgWa7SEWkuV+2qYmfdnDs
mtNILersE5UsKvb7wx+B0xm/JXizKIB3k9hcLNXPd8Ci2pRs1R7jqfp3SHFLcJiXeE3pDJVn+4Nt
BmhgOfBnwufUlrJ2+JD43jJtJWDWF9qzOU1tTuo4em1wo7oXXINxrCMjGgy0wLJO1bxNin8jZWMr
BktjGZttPcXlwsxuVhivFQUrlOdReydIGbkImjpKpfrjdYZOvIyN2bFzekUmzRckRQc+fMNBmMfX
5+ecasez34xnLxbY9ZZdtLgPRyryrVcYIIVbxHXm/gxUKeufa6V0gSf/jaK0QuCu+yOtdX0Z18zb
lPzMwv3GYggb3E8rcAmOrEUm605TgmyZJluAZZ8gR2nHHWgJ+lj8dee9oSxvdiseRXQCIuQ2Ie7N
F9mZhfAGF/6B95pITM6JcteElcon1vkCdqQOk2zb0ak53H9G1MWqbYpnF3cneGrMDhhsfBaH+mwy
76pAHlSYCPrtaa4/iB+vfmW+8Yw9NEYfr6jLl6ToRzcZil0DeEIq/5cmFrvHPwfu1cPucTWGVH2K
HXogrTMGXXeyjOXK+SpdqPErB60RTyblA4JDLC927fQLIIniAT/gATPE+7bzrspCmlWqprhr08p4
4GnMzZ/1R7lljlC/1E3wkTqAx1VwEGKUeJDQe1uI/buRnRoCmyJ/DYNFfSqEs4+uQiR/0K3iOjOs
ODm/sk52tGoXPROCSjF4mCI76MNdnWTXk6B9L336tz2OFuY4rSdKDIV/lJu436/ZgEOrOkyAHFU9
M2g5RHohdz7ilFTUIsppig/r/hbDPQU0hn3rP+9tLbbEpsb93IfS8S7x7I26qMzB0VImFuCeetgS
E81cBwBzS9M7vgaXM5xnNwtByaOXc9j4cvZVg+n8jZUOqcbl+jFoACMoZ2j0SKXuOe1f2KlTVHWO
LKgO4V8khj/0oeK1HWfK8aZNoDwW/X1RS1PbSq9Zd8xVvdWBdFDPkd36vgXYD1CfyN+/ml2yg/Ez
u1z5W1HXL4oHf4NnDHFpYx+UIVWSoylJQ75IkF+3U0vuQyRWPbupw1G6YU/LjjFwG0nbSxVcGLkc
e8UVTEab2wC17SXv9kHewSoRO0LUYgOrThQDZt5iIfAOoal/OBTq8mYB2usk7vg26mL9Nd0doVhc
Ytp3hVgg85fQPZbX30pmtsVuStuQN1GXTdPey+yyAd4AJWoav37VexTAVDz/n55xiGuCj6h3eDMM
n5nQ6sLLa4SqSsWIQZ5NJzHakOAMEm3WETImLFAQFWW+TeEVFL1nVFIYc8ENW77PEyQF/UJcEKMn
X5vDja7k2D/XVLXPygsdEcKJXqu9f9RaA7ZM0m6V2G5/iFFjuEAQKc73w8uArd/mTzG3h30ehvc+
yzb7F1EsOzpCfx4kGVAq44kthAo6mxQmQfZmBezusQJ5eejyjmr7s3/XPMME0RaK8aB2fQWlB9XU
TXMkoeGPkP3K45L5sYAZQjmOho3YIxQ/xSH6UnWjfBVdlEpEU6O9UkKtg7JNc7P2PsRU2ZKJ7Yzq
DH6PdoiQZ3cZ81/qJ2KjZG2/5PmPNBTIhH0KwVG9qc3Ggb5wZr7K1JYkIHKUs7BfbeIZk29h+/Uc
BtiS/nuZYPud1TrZijJJQsn/HOx9dhPnDNdgOerpBanr5nflMEoFdcIABmbgm7b+oINZ6Ln7KYAi
peO14nIbzYNE9Nzz+Ik0AiP4m7HUupFJ6VWLvz5afW/gEMvhQW1G3iX1YiwyyAUGvtN1MxuMRvoW
6XGlac5at0j0jU7HpHg8cdEHPODg8nlNDWNX2ZJXSMyQ9YB7WYAQpXCmYxN5Wo2ttte3vmCX3qpX
yzH5PacUUask0bajr0AckTuVDxfk8FOgMjLynYv6kRBXPYJqwZUOdQ2uIonYYeUsdOti7GwZEl7a
t6I1gpPIDdygFMj5cc/qI8HVTLIuU1bWJKOQQ8C69v42bhi+sndD0XYaZiQNRuDjCN1C11e8hP2q
Wh+E16sTm9QePctNgb65c7qWn3agr8A89tyhtmLsKVyGfooKkudlp7Ul0JoiGdWXO991gPIqzRSk
+UCiSoLIH5OweKTmsZ5/9CC+RhVen2UItuA0BlYxw+by+TMGxPKDtHxa8hnoZBzSPm9QssYFx2/T
LEl1Dx6FIm2qnskELxC62bHMS90ZxNaiuuatXvd7NZJ+RobLpPq8IzVrkek+IUVzA9KGDwAlCPLa
kn9zetWXjXDZ1C9Q26sQWCUYVw5AVwCxLHl6aDZqNdNuQowfw3IxQU4yldDF3fO/gdvt/d79kctl
6cDT6yo/Y/mI1gICxom4sFbKc3aXEw9D59/FYQ9rRnXqp4F8Y3HXJBK9jC6IEKxfg74vWE7J89wV
cyoFFZkEDaRuJvAVCwpzLZ8BIRihFQpQZ+jOtvOguru3abvLPxAvbCVbZ9kzyyvZDEktDzL7jzfh
nNH4TEpHeUT78KawZYQr0/Kin/Y4bqVEXnVCDeEdsSYfcvVoAG6ZAGTgFYaQokTfe5FNBcZ0Vjsa
kJJO8d9r4yvc2vfrpWgiwg/c365LYoZ6cmUkCQMYIcV+AqsM7OXnEhWk4q5wtPnSZ/Bipi9QLd3v
RNNm3I3Dt5STDzlPGpdN3QQgRZeEuwGwJnlZcDPOl6eie0eKc8ZePV03zl5KzUxb07aELkMO2xJI
X/rbRdACWbIfI8Md5yoV7iUOYvNMxN0ZQcbDNINBKqwHJ5vz5ISKp8Zx1jUwdeH54xbRZb8ZAVqI
M+AqbuGHY9/q82+4UCU5YiGwlz4SMtLkwmwGwFNbzg1J2+IHikOyDFWFQAq4cS+teI/LCBgZ0+W4
sMtsVZ7WHhzLLimBCwaTwiF3iRpmtjLbZWohw6Ll5/f47rGg1nLqXaecjrZjdFNysP9oTzw9uR4J
eBBL77mrs+15d9pzp+juqJ6QZOnUcoljYtFiPhkODMi2HZlUUKynsZqg2VZuhTowg2IpMKx0fVer
pM3azRrVBlSUhS6kLMU3cT1C6sU9kHNVTCQvTM0737mLCYgsobI61l1IgPsRD7fw/h7IPS1BsO1O
J2DlxOa0ng8uSadCYjXj3CrY2l6k3zaaXk8K+dEfNT9g6UeiybSasKPkL7iNQ08Xrzi3hTdjZ895
x1bjxPykp7xRh8DUweEmlDYr3J/kQqGPAxM+dHKa3aYN1cba1encDDV3b1lTkS1hdY9WI+NI1FLG
33TvmBNH8ve72SJ2D4Ksp4nbbbifVyo0tSa0PRfvfP7T4HMwXyCzNe9HwNDhlwCcP+8Q09fmn9LD
Q4Yc+N6VLanKaudcnwRP8cWh1sWd/EI+7TbCKYxIlnjylbkCzoEHUxXth4mivkoADgzjnVZYg2TJ
I0Txx/hSezdFnf6HycvRpLmOwti/QBeJ8S2tGXZHtretoh1s+xPENXLx2gxBOGVnts2lLl5h4NWs
fj7kkm2jsh02BzrqkE7Be7YeLV0PqdToeM4A161Xc9B2jplgRkApSXh4etNw8QlmAr8u8aNrkL67
juFgpI7QqYg/RS+rF/2lE6J5jyKZk4SYfIrRUyUSFPqcqUhtAlejkWPVWBNlw3wVwhJLR59AR6Iw
Fedz7Q2ppA/+5L4p6uFuaD8TmHajDGD+vyPZIix0AH3ztufdyTnHzCC6Qo8jhP77kjlZOY0LvOpr
yZrKlnXBnYgckY8yCNNjUWf9Bh+nDzs6+68o9FK2P9DV2qwEJrt0uUZsqETUfjOLWqKjianoloGQ
qS7d5/hWqv5y/K5IDUFQ4jKQpge6YSv33MNb8UeAnm6ZP0RUuKmsqdy49uj1YhdOK3zJWZQoI/Ae
j6WO60MdZ9QfhHXzP9iqWjLIRoCPdlW+NCZesbE4t1b5uTra4h5E+8+TgIwhFTr64QQS6iW6Qlhz
HkPmA5Ueizrt/iJB8BuPddc8WOEdd6LrcZfv6Mc2FaRioli2ImrtnQa3EkBC9eFM6N0eVJuYB2Db
+/zt0EX7vJ0gjkWrWMXQY4LVp44gdzI9ruE30rmYJ/jVFsJg7SF5FWZMV5cuR7rBiw54DRGy/afq
sZKT5F3h8UkJcA/O3Z0bjv3wxdwqd6sFGb0Kd7OipPEABoaAKfRE3nk22ieErfRZRCgQgHVfeuAY
6w6hzjTn4FLifw35YutOsm555d8hBC2XzpxlyF3eFeTwi+Z8bPne4erKbBx4m1eJw55ERUPxyr15
jumrn4bD1eZeBpZSnBJYqktvlpDHBfd2p4YwV06fsFvWGDxtl0usRP5fi+zMyGEFZXiqqYQ+ut86
AV60jeXX5eRLbgQp2VtGCMmH4qLMeyQWYmTxChxHZ1RE/aPkEDJucl8zl+7fsClCf8gp7g7RrYOQ
auZuOigs8JAaUaCYBx/XYUBjbJxiDYusNCKAgElFkAQzGZXDlaDNDQj4dPM2aS24zwpAeqCe2pfz
zCMnmhWty4pPld5/2Bi937S4mjwgdbnFZTaqBF/husogm5g+noz+XA5b4C/eoZ+xokuYNdBbYvDr
MtL3ogMiLtbUxIhisgxAkx4zcNojclpYlRiExlcDyot2ieO8rYHxcGqnSskg+AVvCO2akzc61Vj2
/xBgh8KXbywOetCICZFDGChw49CWYWb1JA6YGnsOZgQI4Y4l3vf8jVXOpk5Hf6enRFlisrH1QcLM
OjPXxajYyrz/JClAZBc/mEtKWBBgo/VEv8UXSY7on/Lojjr5cUq8ZJHQqtlS5BRMSCtQIdGJDbMZ
Xegze9P1EgZvMW+DsxYX1KdYYZCVCu77oei4C+mfcKaXfP7eKnKLXDCgTN+gsQkGJ8T6tjvHe4gb
hZw5M3d1Ql4Sgy4p3oQLEvcA/XdWPI7HtXHJV99sEnqrcW8w2MLuTRKBjTKTKoKfLya+wvY6yeEW
gaw6BatA+Ji+88nDIJgx0KVc4OGF2Z84GH3839mpYF3y75s9aN7Qvu/ybXk2edD/p9/M4l4nqGpZ
duYEWEfLlAk5+v8Mwwok5RLoYdOp1oK+dytI0vbus1wQrYSiKK8QVH/pMIRRq8gxuO81DfIUxKWr
RUuvoooOxxZqVeE6ZRT8wuGTRj8kCx8BxA1AEFHD1qRsYjHab8N86EZCR4kIiuNoomTJ/nWZOY2y
aJA1RzBN/xGtsxyjiFAJzRSqwKHwbNVUyU86hLyzwEq6UcSVmiM5ti99DwGWfEYhNnL0Xh0SV0sv
tze9U89p7rJYFBJi/sZ4m7VucKqE83bJjXlYkNjSYlymk6UPJL3wa2BTifVzbE0v3WvEVRQCMfs5
crrrHzNTPmfzX6/LmCB4lZgR5CPC/hl/XXLM9+que08r196aHjkA/WQa9tyvzsai2KwJki0PYEwN
2SxoeaHqOaxBTi3Vgu6XCjX3O7mVFniMVsz0RpmPSS8Q5BZ9K7QtuzgsAm02zLMfami/3rr6LVxL
la7nIQOx2+o1YIcusAjaGIO35IWePZzKBTrVloRSaeLw3yK+efC/ikgmgCtxYPVREsR0pcNmskIx
T/qSRkiJLjoYpVc15L57DAFq/ijArT1mYpBdAmvtJl+tm75+h95JAdZK7J1UYBNj7/cUJsJoa1IO
/2zpypYTpYRQFBJBj7JtH01h8/DREbqVE3hdcX4N+kGlVLY6qN/UXMsUjG59mbfDV9I9ORZJ4jH1
a2KYyIHT4Cu+yl9sOCn91eM7yfRCTJyYdOFyga809m26DLwTRp5R7t+I2T5DsI3n3lUmaNRi9HK8
wV/mAkL0MLbM7GYviMricuSkoDeGymT7d3oArRTnjZs6C/lKoidhHs0o8o6SXUBRLqfh6mRSJwPk
VoGgce7JwHA6LWBDSv5AXBYvoV0ZPe+FiFrK1soH5v3BpdRVV1rjSR5xVzmxmJaMBM2TlvqUlKGR
v1W5D0ocWqKopbtdA+wX2XpOSoVKafGhoICvdZYPyREtxkTzRnSZwB5OLukhk4dHRGGJ6qhJlN0W
vytFZRxHQgVft6lFy96iSD2W//pEyE24at/YsB4TTv7NwotBRAb53KJdvqOTC40r3I+0hXWzTntM
QHYtX7TR1Z9uBczsa9SNHmCLCuZ/ZVogDPUZgoTOVOlL8sqlOASh5kZ986iCgcr0Sgz6aFajh4Xh
nZpDLtniKCyBiymnMRbn5ExWYZYz9/rz+erOnkLNdi8yszDLB1dJiy+XUePAasnvDQtXt5kAoK2U
tXSDDiKmL1iIITwxY6NQq8K9xxlY395gH9BJOa4xiyT7X5GLW/nneF8XsFQKQhytha0H6W/XF8xl
j01LET6AK30FPfD3hNEJcdvCcbLvBilD5H9N3nk4Udwf/N/Rh3oJggpavO0+5P2KR+/wSmChbOo3
Bo8xUOjdgX/fRlc7SpGh6b5g6P4mDnyOJMjA4i5k4MfTBEi1s6aWC0SR9+f4Y8VWy5QsSJELiOIm
jl8M9BGjxAuY5DljvnFqjZWBJQxc7rmMLmt73/tFzGAcXEfRBDZet/Sv7oDbdFrZZ5U2ly/d+jrY
WfLaAFwulL+lN115DsQZWYXntsBU4nFE6Rgvq8lYG2p+I8BCJHaAqJjAr6FTzo72nKq2QEtpPPto
4XLZ/BXbJhpxgB1mmki6FxUoZGjEJXDDmhIaNMPSjfzRLhSKWUFXXqZOVAp7D9HB7Mu5z1mZAQ8G
r5ThSmOUForEcldDlnUrV2+xPHTsRu2ClSDBkRx8aYkQN0a12hyjpLQ9FismFyZN7L2IMFHGXNFI
zt8etd+P0i00tkF+kemeIKbcla9v5n8T6GORqqWwkLzSgmnh4by0FQqcDFrJOMCFyPdHdrifgLnd
BKvTNpxdGnLyvQIhA7S09fpIw1RDgS0+tGnXKHVdmvbJW7W4x8afvM+o2rQrhhDnOBx8tTI/Oe9l
ZH+1NSEIhwvM1kJ2q353GS2wOnhmqaCWYBHmNKs281fkWZc2cOWiNAnZLJ7xCOOukhQDoUjHuKGF
kdbrU4mGbCdN5HHbTtSuJLle9VR5UEBk81OUqbfnjZCeo3MKm8ang0zKfHAvQU7aDHRIIIhmxXt9
/OBFDJaBMu9Qqv4SOQKMdijEiMRftHT+d3qwsnaBCB+T6h2XQqZyFIik3gxgSfG86V0zhcubTEGW
DVTKHO4u+XKerv99MLWffzkL72RZJCPcrEaR8msE2Y19voyj2omklq9m36DPjEU0mB7+a4fX5HAg
NSDPRA5jALcD2qi3Ajqgx22FN1U6F/KHMNsTmp6cZvAa3ZUVXpP3J9RftTBpw5ffYY1SUgoLO1HL
PPxdCcmxAUvRTHA/evrfZ204+Mh1vkUtxRmvWoaSZGPFvWtq+FZvV03qlVJdGOwBDOlz0C7n/wKb
d5hJc03DLMY9GnU1EgvLne+I4j2R9EOsZ5VXXlirU+6wBZREdw1I3QQPy52rZ5b+Fs/BYSaAgMyh
jkRFrEj6Pc8+Nk1P/NR+ERZXPrd1IRjpIgZGREIR/dhSBdcnV1SNAukOM9rDnKRgZMBEkBgbsBnd
q5RQPA78/vRp8Gzrx0F66bTb2RsUbyXkmtOHIaKZD9HRuIG+8sMsfavBpGthl/d9vts7/VggTecE
UoTXAQwQaRwQa04eQChycyUxQHjYW2ukBtgleG6COxHaTrRT4OFjTQRXFkO+ScVL4sKqObXWU3DA
LhXXnO8YoQs1hpQSFA1SW+uMuTzpfSrlCCLT+5fBjcO2PYbgOhGaL0rHu7LtAoJg8BuhqJyNax2Y
4LRa29DzkwkU5IkbiTau9uDCSnY89LWnFJym/I85F+9wkBCeVnQPktHIvfVZos0iaNrka8lNJGla
epGDAC85EGIx9hn9hBbHHndGGDsz6kZvCwQS0bTSMMXfLPNnCpHssZaZCGvcaOBJe3Rg/oUUyVXg
2IQyiWl/K8rk+COCcEiFo5JP4QQOo8+Ifg7owEXzkSeBvy5fwnIdNdtLM2z9pYSK/4G7qZm+7Cez
wShjaic3FZnbI4/wKuT3CsrVTH0sad+3fWenigrssOrGEOG74HxRlC85Vjm/3yR9drVlRBMLfHD1
0XykAsw+9S40Pov0hjpWnJ8X0gJTxTgy4Ey4zN69EkeeYZme+afxU54NvD0trRoTgoTnSxq3ifgp
zSHo2EPbhGkEloxRwYfFupIJFvfDiK8THSI5Mo3TB/2vPArSxA8ihsBxGUo19UEN5miLsnJRCQ2T
kIIDJ5OWjDOaRtQnqxScBFQYoeMYaqJUAhRMdVEanyrA2A+Mz0IWUxUdVPHK0zJuiMoMoidjJ/S0
w6RakM0QPaZ3EfVqb7ttak3FKcpr+5Yc+yWmqKbDFDpfs65I80L4rw4ybQXVRGv633H78lrpmswY
54Wy9ZYhvBW0q62FjUnM3z9ULkVLwn39pwEe7PgPtTMq/HOXL6SgMQok/WCw0w1tCujZ8jQXKti1
Vpi3A9WGXRhaJK4P+8l2n2lZR5nHUU9fVH7ChhengCbcRWJWbuOq1BWlaEzAWa6GP+0LmO3S8hDg
uhpg4Beqg45lt7B1bQDl78R9iYX0rn2KZC24lfEiQDfPxyqyKkuSOVpuc7/BT7UObReaZWOc3TQb
Pkh+/iZ8ZWd+/IpbAcliVx9FMDvKwPom1Uti9rvROjN2KNOvMA60kkgSPL+dV5Q4cvQ7DzSoqe7E
hHOEFjiJJdUGX4d44eZHji75nryUUUADPIu+7Q790e4RjUxu2lAEdwNyw1xLTWL3fvHu0DZTPqaw
S7GhbZmy+R/vSDP9r9R28mwmwwSeZDT1dOPDZ4CDfO65RKa0h2ZCP/mJOV60wHoXWLuDinT9w630
F6AlKGTiA21OKlfJNunx/xaWYtYMqtS+/wmDr4IdMHXuIxlbfR5eD+UOzuAm30E62GdePOSgoF2f
TwCWtt2gkNNPbrUNUZUqPrH31aJ8u8ixdpm+EXc7M21+15gmvdgn05KVVkfEvQtZ70YgXmywVtq7
9LQHRiFoU9BggLFVL3F6E+0YQtzr/584BuE3E8e9VhINRZo8jKuPaJsQpjrJZMneLbRr2wFNmRM6
d3nNNhddOGbfImiT7RakTqq/XJjkXj5McFB08dbHXTKHBcp08vI30yHl+smbGh445tvsHKxn5mn3
coBw2Z4uhoPl+YMDQefd2vWhSfXwl+ZcoDl0Rvkm0FLRjeE9jfu39ibs7nEEzRe9r7QI7d8IU29E
UKR9tXdc/ctePDclw9B6Dm7gyNM8Kv+Af0cNL1OWdAg6xbHtbrb5+0K3RewB1VNftI8Q5c+LikbW
Zx3luVJh0E9On5zxHkaoZzixQ5ixxqDF8XQPENkoi4VeKSTz37JE2b1yXIW3ODESvpsmjA0cVDET
uwjIeLvXV8OBriQ3D0r2cGZNIntdVT+1nR/NwUHxVHs2U9pvo8XpCNky59sy2+Td53In93bEJti6
FzedmisZ/yrV1/TeOiiwwRgG4q/WrfmBTxsw47iedBoUuKuuK0xmsC1xumDgB2oTkzIWcvxtf0tD
MU1aTUQ7jqDcI9C5fMpr50G7BlnX2NiDwOypB+T0CwMl8VMr7NCS6TCRD/wPSlPIrsAwVR2axuXk
oXjf/nLX+T4n75mK6lOGAkh3faw6gAL9zUuurX52c9NhvO78Z5KUAOoASqq0h9EKKw65FuNNfBpa
fxjGx0HLg5SXEQp9FeJRTPRF+hEH7NC/YgSfdt5bWyzFuPy2YHZLYjeAG+fznxL0i/xv8BafSORR
cWvHq7wRkiYq8uw/UpH1RNeV0ojMA17lO4ioAbGyt3Cp+sItFPpeco2xa4SKClEeHRwpgcpcBXvG
EEIinMhJzV/CCEpNcvCd8gJtVc4Y7EpVadqdZsvU18VyRa9PxU/QQDQVu+or1l2HhXm5mEusNmNL
zJMljRoby8/OrFVYmCmvIbqCa4XSUegmkFZj4phmOOx5lqZqqIoMlhWpAZdE0WYitpJFw8fqTZ6R
w2c9lVtiChNDVhG5n9nIaA+sENNSk8piZGha49yaa+mLzGzeHk0VUOiPDp9MD2xWpLpiKHCyuyfd
a3dZ9vOrqKx/MsaEubg/jdx1jc7j5bsud4za6XqxFKoVwy3btfMji5unObAJIhw9wdbLUJDS9BPr
5Jd6lzxVmzXq6+qrMS2gYSL4zaU7FCMLpQzVv4yTcNsvKWbOBgZqfA3uHhnj9HmGxoQtLAwBANdR
07ox3I9hx6FcfVJwzccdefs6U0II+tZ4wo44SNdDNs6BpIkGycQdwShbUj4ZI6u4GrHnwcJ4UlCI
qDMUY3Gvy9iS+HsEvdKQfw5tT9Vp1z5liTAUZY4id2l6IVhhPA7B1Mow0FWCdh3jw75bp3lLh7th
qMwTJf42YKjm1JNiDDAidC2g/uVVnFvVYuSuJtRMLrYlA1aTO6jHpgEgJtpwfoHSeQ1axM15XbFq
Eu20n0JznJTLERELqBt3iM9JlA4ZSrvusWJlukG/4V26rzuUMBpMCahGhq2d68MIh4xMMvx93plo
OIGukJizS/A5gNlMqlweyvfgqQow6A3abUL02NUA2v5vqGBDDQT6nE5IMHAuOojoVX7qfxbLpZv7
0WS9N5fSCIYADYvJVwEYU3Av6iIbyM/uyfTUUkLl4uVIyWITtncLYD76A3y2yRqZGeWVEqHDFoW3
ytoWFddsZ8EB9ep2yH7HU0/Am2JmIkIhKV9Lxyhvj90ASVkYelNzWEdULjLKn6Cg624/LVc/iRSi
YwIsdE9kwd+SkFt8ZaQsGknAwwzP8neciN02zB0C4pvYZ1D8AjwaU3Ks7zGPmvgLJ/754sdeFHdQ
nVHHg+JKGP6mvob2PbgWHd+ysYh8peTbnsLfYBGcSCTMaUITfXAmzr4gyVK5xjwxN6WP8DfR8/RP
13V3uWK379JOehJr+ybm/PkIqeql544sySiV+Y8vMiIJeuxHcKKwGyY1LMiJwYrt2OGVmmcNty2d
gKDlhfMNfDmPclfRREpj37QU7QYhf9w4uAfi5Te3sNfDWmBpfEDgwJtttL1ePXKjnGfFDTTDyjTc
GbaEguZKgm3aqmR8ysdaqGplJEhlRtd3LkN9Ds1fJgpFl6WAQlNwqCQEcSVfiTdsOlk/nfiYk9hF
8MvEG2MGmA20BlYhxNSVuIbaatKJUC4l/sUxN4ewNlclL0Y390kAZybZLzA3CiZ4t7Uosa7wgPlV
ll6bAXat3WY5XqD9uE9HLf1s1Qk/c11f4H+i0j1OpIBzT3ZjJbrpj43LCnIvuVi/UoImiO3qnUJu
f1LcWWDNxioP01mAAO8ZWGEG+Cq4G8BT2YUwhFpIMmAPPnN7hVfKETWPKcEn3D5ppuJ68LKjxLHa
GbInrqifXr0Q0cYVfVPCjX4aV1T3sRhynXggRxSjuoFHtTEqeTEUdeo0tWE5S1aM55bDXh9Hw3r/
VM27uz16LJJwWI6dJVfh+CMfwM5oA7LotdN/D5mR44aoME1qHTUxlOdldPDFKt0YyuJqfT7T+Pp4
PxqcNO4i0ABNM6EJv6bfCw7pJFz+weOTfvI//z2tIkzLwQ4uGOL8yEn+vzlY9e070xw5df0izfQD
yaL6f6f3aZZv9H+TInynQu52OY29ljfDENI4IBgeMUv/SqO8hGSHtvDjbnnJdou/kelN3KMIr3go
GzJl8uBvTrvUaF5XLNZuZHw8l5mZ31qMyQdSK0mFWqfC18hU4MkO2yZ7rqxbluaREUiDhLXd8ozR
czgwHjtDLMgEoau0Vh3MpwoLxB/WlAezKJF6c8UM3imfhc/d9Dm6XFbiYFD/XHFfCJyIEzwCKQCO
xsiJrqklwbmcDt7PZcEl1bUSKbsp/+G+1gn1nNOQEZpBYgCrH3xY6ZbnfzS8/MKkAwGVK4LF7npV
k6zCgn7aRP982JqGCaRQw1ZKb0KDVsmU51QZV13/oFZeCCG/mZ9Nv9i6K6RTxsS1XEQ7QPAN9Q6F
Nr1XDbQqZSTaCkNoviGzntD1yy5aKKNV01siJJmSR1zsyXCCdsBL445AGgdPYhRcpPqBmQA5GY3n
nmurJGUbtRe3seffI0XqrDoidhZL7f2Wd/3vWgZaovhAnbIvRoRd3pXDbFSc/Al6m43jAU2Qm0uv
bRwIWlFb+utvM7KKW561fqaOsJAmnJsdgxSk8JICvp6Hkh0Rq0TyUkEWsfCociYG+Vy9H8qNwfb0
vJ+GkufptW+rSoc+JRL52bcLZlziXHJxMO1goYkuK73b4ZFk6EU4kowx5gCpLPJQUU6iPU7R+9Kt
qoPcIDRPZVG6nZAfK3ib1DePwwQw4NHUyBlABZ+O2K6/4FbmAmhlFPCSPIXhg3bD4Hww2+1g4Iny
0eBl5Ghdj0YpLnRO3VvybrQIRnBUy3hZ+mroAlI56rKAMNKsOvBFMHz5CMYgTwsKSOP+6+Yn+1qc
SitLXmulPJ7FYCuwkH748tiGAav+wzvFz8GBr97nCF23n/5Ui6NsY12aK/I6YF07v56zjgPbU0g+
HGxFte1GfTLPyhGMl2Qw1mYuvBFlcHD+ertpyW7x0wz9Fjl/oQDihGSi+eP81JDo1ZWf5Lpt99T4
BBT7Ro1hn4bi/uNH89/lX9mBme534Q8Sylsu4loQkMjBBNN43pUJDHtC/iVyU3uqjmBJNuxgDH2J
BR9qvy8OfyU23w14n3EBAtbznQgAMMs7QxMAmw9RO69kYIhm4Om1jm5uxQkGR7OOyJh88G0e3fyc
n1IWwigtO4ABsyyHhgKzttsixX7OARKvoS+6aziV4mbu8lKcZmpM8T6KyG20ufRMCLf8FySd6wfb
PQNULsP6Npe1IHQYnQ2yBHSflyk0Q/iIwd7jp6yogdj+2wjeVxni3XssacMYY4nzlkwGdAhy61iu
SlP5yg1TuPz9598dF6xDln52le/puSbDTfDRaTT6Uv9IkQSB4o3+SwA8sjsNKhEHfc27zGTXTSQ1
TvIzOwASeGgdtFWvhWVwVfBDNpi/52wng2mPdakMP2QLdNtBBedOfnM4VJ/OltOIdPOt/ZPCizqJ
7hkYeDGYrwON4h1tlcSwDXWbBPn70pM+yk9D9mC4M4w3TRe77wxLJ7JIsNURi4N9V7Zn3NSc7L92
MNhOP/JwMPulzCRUT0pvSn6C/fu4anScCg+5SU21lSVMhZroWuXXZFmYh9TutpND8zd1vd60BU0/
a1ZljoPGu1mkzj/EXNHP3VHueFF7J48CrbEEncWuNy61M+ttLskEp05KjNu61HskZM10zzlbgArV
Mh26M5JyiQUVUD0IE6c5FsmsrqXynjE5kxVTPCC3WzunV0gupEA/ogAP2DMoar5+3NJEayFw8ke3
2jpCiBKCrl8aKq6yBoW06yUVaYZt9cDHPpOSWShlq70behptk+S5VZ5Ujj1BaK1sbzuD+MYg0ML9
regwdcSZgUjgYzNR2HYmltdQtbAAvIlzM7DvKrlu4WU/mMgvaMp//Dw324ZI94QyjSwB0mgEJD3G
YHvtK5MrSJ9ZXVg2NCk3oFG2wV20nmGKs9zd2ZrHsTy73Xemc+qkxNcLvkgPVKiQPqmPO4pn7U1u
Pk7s7q9uOOR/EviYPtXZg4+WEYIKAoCWG81P8od7MMcncHQDRBt4CfRUFsyAfeXIxeKn8FwEpgdx
xZJrBbbzzyQKZPrShkp7PjdU3XbSyBhb2zhEyTOkSpErt40hqdKi3fY6E3POkLmh6dPKdKX8dSO0
WZ85ZtEQBS4KNyYeRf+lXj1R7E/s7JvhHv7WcMGKHg6Eg5fWM/FtoxO3vMYlm6sksuhAShTfMpPf
ojlNq83Yz9+dOHc8fsbhENZ7q0BQwdvhXXreOzwQlcgHiijGNCZGn7tcNEYrVj27T1EAmX23YJXl
hQ/rG34HYxmmXwxHDs/7sNlwsYDB8xjn3kBDEAc9ZNDHN6wdtguKbz1sTCXKACHDz2jfEhSgIxLP
eeuPwKCwCMh4dRSIO8K9DxwDquO4sOpXghTU/j01DAP/rmhwPNoCcn88T0/toubkxiemEUUvo+16
edN/uvetG5rSfagTeO+tQbSQ6PpA3k/1vWnwbSgukvlWQ6L9y9yX1FRpV79H6SOfmMC+nQCDJcNO
9Wn+zClEqwtM2bHpoG9bR23RwF3zXkSvVkdIbqZkGKYijV3AuYPyVFshDxNcCSH9o6GBX5wFS+J0
0EL2OJvifVH+WiPGkPm5VRdpQd/xop/R/LRdmAZe8vXgHL8A7YrfJDj28JogXes6Jcf+OfonA5AM
oZGHG+VaiFDoTvLvpZX/SoSkoRsQyPa//WEl1RrG4+moaUEkWOEEqPYkKE78zt4aUHQJQypCnO2g
fvb0Gz46D8x9hDpcz9KkrxVsKbRwqQ2yBdLm1bayYZKGP8X+JxTieq0ZML0MyQg/5YIs40Zo0VBE
7MOljWFVgKU74P2ajh8/Mt7ccljAJagbxy/IkMJT7qqqkcZinwuqkM4CGOEGeId03Uv7YtyXQ0Yn
kpJ2fKdRfi32XXEiRsTOVVNhPxJ7WJbDP0klKCD0GVREajWmMngNWnVeEiLup73QBTeGokw/mCCg
HN/E4XIVuPu4mRYLm/yMUN+omhMK6Cik0QOvXF+226hjkZiCw/T1y8jSbfpOLYCpvYouMrvZfwT5
dKRk+t+2mB+85BFM9dSFumXKcv21YzkA5nKMUMZAFypBNCqqxh1pAN1f5nT/wf7vyUKuBzYv2vPu
Fzrrl0QLpPCWsKgmx8Q68//QUIsKpABkNe3COt74yQy78Usi3ZguCIQMtE6ZXA+tdlpnRJeRGV0W
MlLAIMvD0evyrvp8nkJ3hJF0d09gaGO3COYnQa76zQ7PsY9s9xtA4gOstKQil7fZxig3zMOLclTr
cZVPP+f9CKCoB0I4rG6mBkItBkfin9KIZtjGLCjnztbcpBk+QeBYEvnBZFvxsvkJxQAQRmWGaxuM
mjKZ0VudRyjwS+HMsLlvOjCzqVSQ3SWJgAjF3PdreAKuSc3o5C9TIqCrJBDjZeyYn3k+6Cd9iT/g
5yLgZ7cGvgW4ig71RyN/wJs7DF+dzcfCSz8fjO5+JGBo2GNbewSWmBFKwh5xQakONAahpFayjsjr
q+rVYgq75OJZ5nTtQnIUUV/O8NAZRUq5onYClkLFyuc4YubUb2fRsM+SuFUZGdtw4NPRCuhbkECk
TG6YKsWqNCrXBjLWylaGolUr1Uww3Ggsm2MChs1SJNrPEqMe2zpb4sll3PJpOhs//GerPe6Xu1UW
4QyzkM3u+JlrbjySxEBqcKGvVAxAAMTlr3fHlDjH68Z8wAjODxc66ArKXamOfvoOQBbhNViqXJKO
x+nOCLC3ulXon++nL68lUvw4dGmRtH2G/LIE6qECwfjzEaf4Fl1g9/kOojwpQk40ZdLcW1UIkboM
DK22BksuwFzSS4jyu3+ug8WTILqVj4PtVw118eQGT3z5TdM2Pbe3tZ7IWBZTQTn6LJ+IJKb4fqKb
8cDdj3cJh0hYtpaHYRQ5lIh2hfO5qQanTN+KjWWCUea2Ojg+3jiXt6I5RVbhPuQQx173RTLvCJd0
+aZkqFRngoi4nMaORnHQ3s3/p2HFiGkQfuAqAdTB7kc/SJECXrDx5qtkPdk5nFzOC98IU2JfY5p0
yaqqoRMmKQyK8FTMgAWIY2Lii7MDjSKCcjb6/460VBLBxFqM9libJ1XbsO7/1cdE87twtNlXoGu6
CTjlpD9mJG6hKa9jDcjBqKRfsvN0P1JCFxKo/mbHzFjqfaOlxdJWoGGZFOzbzzMMegdywSCICLY/
hCoVT18Ql/Ra1szSwjncg9giroDhwuif9zJVPxD2FKxypaTXg4/otkUBpVzmOGsxu9M8K254AJ+y
LQAz58wLAEd2KTDFJTXGjf1gPl6z68thheBnCjOP3XIbYp67jIksxcU36Nloj+lWqxz8M7ianGLS
b4dN4x0trNhflQFq4Hwu4Qn0ZUMwmH0D2/38NuPEZ/j6SiupXXBNiwLNWCSIE2sehXlvpQgKguLR
N6vFkudGK+l2FM98YcYyjduuemyDueIXT0ws+LADaVzhrhcWjl0mEAUpDj6lDQW2LSZyrZ5o2UKY
mGc1Z2CbRtQ1T4pN1ftOLeiqWnU7nywVyVbZLvT9eILo8ILMIEfd+5liuuSeJhLdLy4HPSoiK70+
wkHmrE0ak7K5XlwmK/nTs3OGhAEf2b7XpcvBnZry8BZCkWZ/pQ6FxaSq61y1OPvd5fFh293Xf2n8
Kgw4GC0hVM38fX3BSe9sjqBDBc9PboNN+GF6/TV/lduiM6Q8osmuxHQh1t9Y+Uf6XNiPZhuMp5gl
LLOu7mzrFEsVWhdO7nza1DIswYdY3fd4ixhHiZ7LbbcDeWvcpLARF1W82aFjXeGR4swen9DpHP1D
Bf4GAaPd+24PqAb/BOxXGKttQ4abx+ke38ECZ1wCVG3OA2Vb6v0ntAEheb7BGTWwGwIZA9SW/H6n
NoF9wI6KHACpHNDGbadGPj2eor2qzExHyZ92ot+ahEB8cunQSYrruYw+W7Py5CezA2oCD1pQSj1q
vTlhLoZ4ipfUcASwHsNsOPzlbEPmFxTKcCLqXhq+96RP8t3VtfEAe22EFd474s8ew8Xq61apv7Sb
vQ+Yg0nizkcIbCmVoXk99iovkFT2G+ZLdgkeEj3zBWcbdjfjq0X8xcrBWIs5XpfxvnwiX1k5W0gf
tQWQp1ejeqQwpI80Lju+bOmOEQgAi2ND4LmRtZrmrbCm9DSmfFx9fxokaI6r2z+yfgfb0SuJoUHX
DupXnclacjvrUhMcGVa0Izl8iNSY3lCzq7JcC+5wea68XD2nj8bk8+GAc5v9pTorQPRrpXUU6wCJ
1qVWSjIL76WyB49bEUV+UjkwEFG6UPWP33lQzydH+kpiI1hPwTd45V+DoI7MyepUlWCD0BlKWUqY
oASxTH/raPsTI7e2OF0M42M+2QxS5wgv69gYxRCpx/m6vN2IiCsNGOs25K3/0pcJtV/nyT7kCpFx
P1FMZ7qskSDoJLID5BmpKybVWvSQG1800KEOrIUq6aX2mN8pTRhl1Hz3B6C9xwyxOZtcpNm/wbMu
cHp7WhpUZ+IoFxPhHYAknNsQqPEX7zoeQOtb7iw0h0wgeMX6HfjGJ3tSedLI2Vx4YMwhpJO8WTfa
p7QN/63bhNL0a9+gw5fboexxyvAlndUVHtTGkZ60p7ZIlH+38exXjPdusQig3zMI135940UGCS5o
ZI9bV9D8eTVO7zPLJG4WXJzjaJtSe/BHUB+w6WMFdGYP07mWxuplOLXBG7Im5c8fqntN8ExktxbT
9OeFdDH3fg52OkY5V67Zt5UcbUcagSK2BIhV38a3c5BZT9lZcEeBQxgIuupOPAdVYPaTCcEmJYu7
XvQC/kVeP0JpFAHDbfYN4WRsG+IxuFN/dvS+C+xP/qSn7t//Jfl6z/c1ka9cnY6ac6g8sz+5V2tQ
+iUxroEwga2z9rOdPTeOaWCC1/GWdr7hhBsyGjoBGMN1sSVtzgUVnxWLk+a5k/rSyXRXfzvw1rDG
H2+fFuzTGv+Y/XZ30evYJ8dDj5l+4YcExHUYD2JZ1DIfTX66oRqL4Z6SFsaST/uqM2imSCvTLxAf
HPAa9v+NlaKILv2cyZaiza0dOLFtbo7fL0o+xYuWGL9ld6eqWCS+o7128ll763UHb7xzCgb8mtRG
k9qN9U0QG+91LA2TitPtSLrZD+CCKZkM+5voc4L1okDHXyI8ZBk7nuM61UhfMvV3J8UmcwAuSjfq
2XgZr/4CpYQAmMkF4eKpf4vLECykBtbn4gcVvTEWjQBWxaVUBxbQdzDl4zfWvYdAMzQUa7D+7QrB
1BJgm7WY1lZd8iblDeX9WMPhcVlhjoOfFiIBh4drJWGo+MKts5ZqOK8tbgVTKcPGM0QU0FYTx0lb
lH95MWz4Hfv0qX0E7SAe4gzwW/NOX5bHos9mtKxbytmkhQETnO85WKWCKmf26dDcdQv9of/JwyQa
g75KxWn7RUFHzHiidp8sfZRNZTGr5SzOHBq9WXiifT/RMa8oYs35hI7bSPt3aqhXq5qrLeawQzvt
RsXaVAWkAbPzL3QEe/jdO2a2Hy6RKmOkz+b2q1d/V27LMaU4BDX1Mu8JJqF7q4d5UDAur+Z0AcV/
t1gtCRUttOfNmi9/DVETmWQKr0GOkCLPVDzkVxlcCinW+Ko/90XrbXsFnERHLBBD4lL/Xtcn7WJR
WPtMD+KbqFv1tILVItNs0Zf0rzOWG8uzjXzSilgQXoeL4Sa7Co/YKNc0jLUh1Wxz9iv9UF2PXkmF
wWXhyZZ5c+FGQM+NSjP1jX2D/YMcek3VteXJEQrjhMSdG3FwJ2KOqCL2QeikoUFpDigp7KwRZAYQ
zC1Q7a7nFQil92H0tJEeMn2M6gm+Adxq5zGnQwvfIB40LIp5boZbtlcJYyK7/FDym7OMbOhXchP7
S8P/yDxy7YvAP7RDvk0Iy4AV3nQvu41LyCxNotFekDMt1B6VJae5T0zxYvcZX+9MN7w6+rz+b5dB
xNVwuNEB7VQiaObIVg90iV0ybYWIcDUi6QFfmxijnamyuLwht0zlq1azd4bT54Xxs0xMhg6O5zhK
SFLM+VnbcEjLYoFdGfNSWyhMc8hcsORNkZeoE+SSnFTG7d8IiNd/ROWXJvGXN4HbrMzcku13pgtD
q+kIavQVL7xVkXSkQPUkx4YvAjD4i1dFs8T4inn07YbpYnoth0MmpjCP9Hlx7VtcPDPm5iWceseA
ga8nRhzRNhDXvrwXciaRRo9gR9mvz+u7TQUWgRV7Fb1w2yqyewdRvby99uP8gGyeuPyi4mvOneMt
CcrR48B1a4AfdWICdEZBjjR4iLCzmz/1oO/wdRkU+hv0keAEyU6L+j8NQuoCVzZz7qIycTIveAYI
jlKpqRBjc8Gautn4VM1Mf3C9euh0xR41SeSCZU20Y33BmIiKqtXfFURu5pFghfuaHllAjp9AjNt2
dUN0OnjYq94SRWuIbVQrHTohCgyjH29GEAxwIWBlBT6BGl2Fosqr9cgF1dWrfCby020LJzvyy8oA
N7SiSHWV1/F1Gh7LargXc9fcjbRTPVSMgP3Yn2rGQcEOMvB9UORee0rPx2mhLqwxxfKEHP3bQtWQ
NulXyzRzWsZ+eQ51LpPYndB4oAFexw7MbTx18OwDvzmmXSeGFSRICMdH8Xugt3dRadBaDNIdUHCq
4Wi1EMfFO9Fzmvkr13VK0mKyBuMd0QGArNQVU9l2niEyW0rGFohSQ8M0Q6am9vRoOKu3TeX/8GrB
4/egxvhcm2jBROKd5X58GVXlVsW4yUZ8oIuDZeUcx2+TaqG6hWqquPtPapLoUJAPin69bYkdDFyV
o/vZyJKjH7W6ay7IVw4WWbya/mu2gGkb55T1i6BH1rMSoCJAemoXf4enAe6OgJkKpWlrTS38tmCv
NtYuxHy2VHrgiOjtuUMIdgc7wLkWAJ/zo7bmoHuA7yn8CFGw9YTh3fGPF/lS0/FLF9EbOax72ku0
PW/Ig8ckbsXYP4eM1vrTeGazwZZLpSHmFMuD2Jz3070L4gWU3mnOJUcQ9LjxWhwQVOyKGIy3TV8X
lz0mWaAX+Nnr6vdvvHIMOttVVkbF40yoxtnOWur8iJ6V6SjfcuIvAy+5oLGrG92l2xAT2/bn9KNk
AOwRE9hGXnVHWjaIhMUSN1+DOKaWi3EAkdsKZH3wbpdZxAo6SM12ZIYhkeqTOlDxXgwZHhjN5XAV
BSlDQV9q6Asr24UZYaa6JZlK74rPypo6c/Oh6SZhBBsEUAiYjd0OQPjvoGNqCi60wTeG4KZ8ZhDL
3woJ3GnAXCDfRzkWQzc9HwZ3Ksorf0jgktrqPqTdVzYR3h8M6ne9ub6OP2b1X6TGpN+6qh26Ro5T
dnZoK9RRTYgcALbrSF1doi9WVvutTXnLlZTyHSnpzFLzjsINhLG+dPm5WUK8C3tBM13PCl8Itxay
rjUinCcOJYsXoeqpxethe3o5AENW9iiBMLnxv/yovSYhX0qa00LThOLc/KhJUKdKSaW47BlffmsX
6yM4gCVCc5jMdeKbNuElhqFE54+CdfD8z4wdB5OoSMWgMx6dAXI+m93FCwxe2sMiua08QqZRZ0Nf
wtdlYdeot45zwJ0tgZOanNCTcNH9MkGs0IidqO6jsTcmaZ08hGKnfr/7qBiu5ANASaLg2CRMeOCY
nADx7/fHtTfn8T2tWMBovfUWpN/gztB2iPHSzcRnN2mDvHe/4LYwbq/r4A9m6wFxfRBGZww9yHrW
Sc2Jcco1Xx1PnyPZazQ1BRQCGagR6fV13Izb8E7eMvAqxZIW5DEgYHlys7jANfhtZ08OgdtYMWPv
NVFi/r14eHj5oxt/A4cEwZHQvTGnffOa17I0FP26ER/Q8G5halJrXq6tjNJ7irxzidZXkeMEZukq
9QDrCbIQt6m6e383O3EAHkNTQRLhTuH6HoScMBYHQY88sL93EkPuicRVuHjeNtbvP9Z5iMf9U/KT
1IFqKl+TNpoxqWYu6Lk0i7Uo5JmuEPp3vD7NTuAADI35PTrsd5Ln2/a8p9szuTTBtmEK7D6Z5yFO
gSvJUlDc3Z3tHPgbW5728yWh1cJ0jIbplQM6bAT/r17IahYVJXLKzMPxd62zws+y9vye+4PUXW4C
DUNXZDVx2ErXvf1cSqgFT8Tvs4njRDxyS+LXCsctiGAIfssnZOjpV3m5mGu0xKok4QRBh9Jp1JCJ
U1pxs1v/4WapkEEzwxp0Bncm0M6bO0j80U3i1Uqz3gdjs34Rr87DENH5+JxlMQFaV3l4FyodA2rM
xIzAZQ/iqMDSvw0yRzauHOtKaBvAwc3MqrU+jwGde1Epxmm17dyngm6yL+GQTQlxU2UV09WQk9Zt
lzNMjJbUFRMaX7U9kAqUZ/q93DmelJqfLaYa95O5cR7P8uYdIDbWtD25T+J3WE2LZxjoDGEw3vmq
1xf+RynVll5zdDcJ6533n8ZUparknhLks3VPg6ozd3vQMGUkikesgTDa2zZSRKCXfoz8CFwMBTq4
eH6xnGI9pu0QlNqHnY35Xv1auIvTZ6koOa8FDxVXRlrKUbIMOMEsKZJfG7Gy4v5LhmvvU4x+IjQB
Va0rsBh53mMEyPSPtlgnuzGaclDQA35zoG5oTPo9bnvWxmUTJAJwTanlCqCNaB9TCna3g1Yxms2F
dYmNI2/xNknFSPSviOJFzBeRoLdBAYdkHxl7HFUHT6R9qUcBw/h21ulUuDSurs4X9I7ygaFSaYea
pTPmVrbkWwQcbHq6PNwkUZA17LBiKtjL2bPKKf/os9gZVReTC/I/pucB6XZZeQ0FNaQXuLUr8i1w
+2nwsVsFIDUoo5fMQkOU/rNspKnFIYOXxl1Na21ZX9B2NPBl02J42lYYxYqiePXndZp9dVm3Yr9k
MWcSs+w3GrQ9KxN1aKKQfJe/IugxqbBghd1XuRYKh286rggk+BvB9Vmy5zOQsRvdflLo3nm9eW+o
dEBf/0vVGFv35NxAvuhuEn4BBZtkfKukPrvqZrk2TZlHF5WAOiCLT+4QtwnWjz3PZ1fU1Phxn8PF
u9p5LZ2lDLCLM3f9FztcF4Lo4viMu/y4kR8NPZoD1N+Tr0ktF7aTy3ZoMfVUEZLsR79b103UWzl6
bvo/RZOtVPbN1UP2yhpM1y/gYIU0BSnaCmosyQ0U8B4VGB2e/Dh/rqWaJ2kY0o7vEf51EVOlZtfj
wM2moGIIvzAyfufqUtNKba19749ElRzpALbyL+aCWW4DVtXLHsWa4Ro7wlhpbA37oSVPO0OIXehy
OAumXduCSWdjZcZ1daMT9JYdaylk4Tzo3eobd+WCVq08gbsxayaHXIE793VUDD/kgb3icICfIYok
8Lr1KhzctyFvUMC3D0+/MKJ5Hw8eNSV5QP9j51dx0rdiI5EDqIJqcmlW56CSutyYaH5U30QXRKhv
kezANXhxY01AlXBBmbfmN94Uc0l8uejBq2YrT0khBW9ZoGn6Em0RnoUW1Ex1ZIdlo3hQIb0/+Guu
sugJZRpOca79IEmm30GYb678FDWl1ecj+6OaSnectsinn8zI8luWpJq6JWRCHW6BYXJF1iBE6kdx
U+Ow/3L7NteWHZe+88SqP2zw5ngzcrEqefka4Vgoe1GPpaya97t0966dobw4+tzQWFpDBdUKM5Wz
if5r61I2+GEdIjF+6KDwBB+NzLZuTY2anzK66jk+0onsg/ahgfOrBvgK/i6UQr0ZAi9WTjOeWIbm
ovy6VgOIhAKgX5VvyKrJozxojwtTbs2Dz/gq+HqEzsDAWR2eYK1I2F7ZmD7OSFyzrMx9OZgDKs8S
uXMWE0/fmcGYUe9F0uLdeBOfnkUNVn/n3Qbb5S2+s56u+jIw4QQY+pq3lsbXqg9e/45spJuQAvQl
N0wdwFPpNNQwkWZqH3J4FfcATCPLW8udBVNzEmtcmeKP0dyBpVNf1IvVMwy1Wgh27WBTDvL1Bwd1
Lw5JXHZC7DWp9tsgoBW42iA+1RfK0kCDuybG2hJzsJiZ4Sa3SzROT8KD0vWtupL7ZvgExU1/0urh
KgNw1wV2DIrjwzDcmVd5BAEe2PNWmpMJ7PInX7nV2vAN6HhaimoWy2V4v/RMblfSVcJmUf5/HyHo
nnpsEuHMrunA6W2vhMfhFFg7M2F+veiBjhoxHdEi4StSR5J8aDolsYTOkvu4L83niBk96IW7fkYE
rl1QqglKI35iJW+MYB48zvFDsxWl/pMWjijYEowIiG+2YGL0cgGMfuYVdGLdD+9ZlIK/asxamF7H
tEK0Eagpp0KMXPgQ0zVt1aXESIaIb6/J0ASyeWxPilvJcwO06fB5cZBQaP8latfWC54BPLiWEb6G
LXNq+xZwIFmxOqL0jwVi0W//mSQ296LXyMpQmLuQfMUf1L0UzIHk0X8Fqf5X3YE3Nc7NxfrPP5XL
PpeERVl9uDf4LNe5OAHlChEus6D3cg5C1a0JhW7bj/hRwrHlozbPCi/S/i9yWhT89Q6f2He5rsM+
V2kOgsu9AyqB5TOSTNsLMVciSWkynq1A2YyNsI0zPsgJJNNUpPfiqjewnp9d47tEY2fzM3fdNquQ
xziY6+gNyUyZPvd3u8NbnRKfaqVcJmYGw/Z8g9EWahlFk3qGM4XDGLCEy7jhBRWIjTT7uMHrvNuA
aRtLysVhSklzyBvqNGDyr0ExbfZYL43vxhUX7PNXjKOie6h9FKWTDCRuH0BeYJFWw8ooTJZYMLVK
F8k6fyUqSkscC82tZk81Bo7A1nHAcKluwHboR/u/bAZbVllUK7syQZReSSF0p04CsFhzWZPrmWjI
c9nvPmpvpx/kZ/vrg3rjnDBImM2DwmK6cvrBH6FtCsQHhKamwNtrGpzftNE4pIRB8939fiyOA5pV
LpRx7hOj0MlAINP7D0nYujXSSpFgtF0rX1cbDAkFmufzlqi3yZ+E1MoMWSWagSLQF994aMWW4H9C
CiA5FEMePKBuKdQYAP0lKOxCbKLJreirUo0/IBCG8JHSUF4ChYvHbiKjsQQYIkSNaipgO5mFnABD
1W2+Fv+nUU3bHB7OeLr+uAmP/Nwnnj2c+ntekKYq3FkUVo6E7+7azWKOHPcPmUhV1gXUCiwWrP9b
FWmhqXuOD8BhNa/C5WFd8b5b4FiYRXKwduXVNZmm/2OcHDIgJSe86xy4F9I2huuEQ0NYZeH/XjD2
NATm4YJSm+JMj8cXZo096RZbgLqItzNeiTvbBPtMRqH7C7bkAjCIm+RJpEbx4CuUcc+2o0zuWlYM
M614C1MJen+Eww3XtjY9BPhdnC0/ibHzUwUrL5FJiZPG9/UCxbqoh4uEh3oB3c+FpuHVogtV1PCI
VODcoMM2N3+eGtaNsmOPTR8epRqGR6W7uhq7KxRWQE47Z9ZhtDfVgH1EoUFDSN2Cf23AC0gf+Ffj
xF1KBNf0QxlMmOVAOrnsMKNOw7WFl2GVNYCyftxLIXwGznoR9V6+7ZBaT097TdFYcaQPmZ+INDdb
ghZcWzQLCfQBY55dHcTPNe7MVUp761t561MT49rS+UvQ1I66KRC9OV6X1Grtpi+KCI5zIh9bUg5t
Nmf3vdxv3y+HW0KrBoVpARcBYgY54U8UyIRph60wcnjhyvPWQ7mhhFm0Wi8hn/prCX0GjMifsPDn
LDeVLngMEjYrWqAsEf+Jwb7t5gftxMxvqVJUaxJgRh/4zUhbx2JnvIkNbe6VaEZ6fJhnjBv36pgW
y/lTNa+a8G4kzVj3w2lwXCNfVwUGF6jDQc12PeZsNCsipB+xmQz1w9BDzFD6VB09wOOt1PtYWaj2
G9m/zE9pmPwks3U+V8U+aEc0RYBmHoFnlBfsiVUFOHfAhAsTFHWAoR6k1HEvWsRBhARJi7MvENYA
l1OpMe+Vt9mU+u6FmpIawzPtL/mrrlM0sZ/Htz0VHJ8RJxtiNggSeaG2PdQpWmbFwJ/YE9ofquaB
/VtJGUo83w64PJViI6Ul8ZkdX/dh8R8vCaKhEUuErGrQc5Wwny8kdnRd+2R/ZN01QrjEgzrGFYCK
ugccFQvXk68CbLot5GldyOCxAnUfTDmlBXqWbsLWUgrdWKKAx3kgurqGRA5qus8etSBuCk3EAaWS
lyrGkntqlFZxPhC53OTSvZErulsHmRtM9hjJ421IenQWhzPgdCxj3KZ86WrdKGSWTG9LRNdraNWA
qKWyaNX67xoMLTgxcDgko6iNGrtlGbvQkA18kznUogDql2r8dyA8XAEVxFv7APzxAprIOE9/INLy
9MgTkP05ds76q96Y9EZxo4iWRar0YkDfPLWg2pLTjOdTkue0YxJGFxHVGpNBK7vNnYQuq6G2d4Mj
XMjksx+QwN0CSCUefxqSUWlGiff33xVVnin+MMY3cI8UEIET4y0WWQgky5FXVuh9Q2DaJxYd1RVw
xNyxhrM2VvhFl56bTQ9TQh5uJ/mDKocAMcHv418QML8hU5+QnithV+nrNCxI4gPnM/jfg35OKx38
Hma0WWbI1qhqau8/L0VR420pp9bLDVtDNwZAKsdhrJ2tWcKbybNiui04DxofjqodY5YuhJvZKpGx
wdNi97+2Dfmstkc2B8F8P4KzvQkPDs0HdoHRyVOntASOH3zHxI2Couw8mRiz2C3AYUhsQ5laXIgs
pv89wletE8z1nn6i+fPq5hWAmzALtoYu9RI9eATSoj+yT+gXqBB9MSdUWe8JOEpoSOwPt23YcjyY
jcjlSGUa2k3lh7KFP8d2lK/KZx/CZ5LgpEF5GIA6jJwabRZylEE4ovezvp5Ug6iDip+nwCrL1b4f
g3s3HJ4iYTigeUBOKvrabbc8uzOYjkR9aOEmyxsE7gT3BXIStEad0ODYPxquerTXLr9Mj9sk99Tt
OlWvvlgz2RBVV4ULjhQkYQIQnTAMSr0nU9VIGCidwwVQV06ZWSOwjLOppr/y2dYFUmIgBdhIer0L
NcdEubSoRPPCtJQOK2TOo05BPpsr6KkFKhBTYXNCQ4I0ysEq+BAxH8do9x07e4Rp8d3DJLRwCrZO
AkjejZp/HXOlc89FLSSBd6GDMEkBDa0NSpxy1av6wHt3zCBB5t+VaRxE+i6rY3W+1i6c7QNvcbzL
M64iPyLFj3pnjJYr7NIDIdIE3c5TvLpYQERqMBWNlVS4wxJYi/jyj+drP1AURyDJ2U2olyHL9ix5
4nzooa7edDdzgUUWvrx9n0JTqDAn7fuGoz6YR9uvdtxDULTxlhZqfEvMLueJ7b4k4Zj2y1hl14iA
0ZebB0JIR5dcxwM8pXm2mejYOtCibApy8pZg2EK7klieiUWUpq88XCr1QjRuSvblte+T/KIsI6XQ
qH+OUJU/I7VwqnuuItOdsYEUistcbeWG62G7j3E3DiluMN8JT0vnV+LzabWr703s0nxLEn1DA2Bm
lAuWEYroA3oXBFL9CF1DkFpKY9fUyPW5WYOdnlChoRTz46EGKUjLWoF/kpP7IZsBb6TC1pjJS7IB
KQstJjcCYwb8VTuSRkgpcy7x0Lo73fryxXQ35TlrMaD/scG/T4O6ewkS/vdsdlKij0uYtpoJJo7A
2Nbx1dR/KOFuRdzv2PlWL09MWxtTNNlPskMwe46uzxXu8h6pS/8CW+sTegoWNzoOPtAR0+R2CUL3
FYRUty1Ad1S7Ade2i7t8HDVCApEQUXtPC59inPgRqUMaVKdibIvLawSapvntk3iPW3bzTFn0F34x
9QYIay7bWOVZ/G7OumXliOXS81l9X7boqhcyIEaJGDzfTKI2oL0w+8YALd6hdnNBrh/WexWCDxwW
DaR7ZKvltC1/f+DImHOlZSdCoREoFWTVMmLkXLXhXdFqymPEV9qxkOYyozAFmjY345OR7weGat5A
hKNA2ciuhWEK+hYO55FpzezQel/UJcWjrqOAm10ZEjg15Y3Ku+LArmlttwbZgCpDMQHtsGj7wIhl
6me/XLQnqZG/QWZN05DNgY7ebKJmZeMv8hsNd5brytRHnZ7DIfqx75iLRpNZQWzeKIHVTF26fIQI
sfupORiRnNKkgEgX67j/G+r13Y8Lwibt2v3ummHWViVMshRQ+BMsum8f/Atz29suHKgXissy/3HB
vFKmXohXttRZwdSx+nh84R7GTBsLcFXGqaDsIwUhsbbPjlU7AT4Smq3XVMwZpUpRGaCjlxOpDQSA
fTDSN7MkpqIDmKAT1IX91CJ19FXOZZOsAREzoPg482qsIg9UbajQ6u3GK9yD6AK6FhhN2f18LzAV
2nfXx7wIvXFD6eYehjetVqW34dYkpp4vnRegJJSCXavcKv/WpIjdjPtn/WadxOM3gqMgRDwHHKsn
iicKj3pEIH2S8qTx+Mk4tVmZRPGmIqUa6DGW5VU+N57M+e7n39t9VlulMmCYoJNQT+6DVUkC2Hwm
IuM1Cf6+6nrw7iCGn+gXk7z45A0IR9919U9gj4m2tDy+fM4BdWp6ukiu4Wugi+4OwKDN7UDn04aZ
5MOoMpxGSzyA/jXujlM0pNuz71Ud2OySrg9Zf2NcmasEqde28C5F+D2Ou40/PRORWYkAZWaAUdDP
G9QIDwX5m+luY8A4JdDFI3QhAp1bmjpc3Peiy4jvuSefoBp/aVcHpFTH51kFtTdTteT02fj51cf4
C9hcHBaDLJlwXHBRCDywdKtwnZIjMrfjkpX44SWl/Vf0EidC7Usv22C/c9FQJUDdai6l5mv0c9UI
Eh+BPoRFs2pCQbvobqrpc0Z9/ABccolj+JKvLumzeMT/Im8V/VdNJ92cESYgrsLapsASV/upBvpN
7A+SPmoasl2r/oO9YNdZjbXSaJioGYshF/U3e8foDOweOWayWSo42EcH+cEbml5EBx96nh40SlNw
NsnqffSDCQ+2xp2vq0OlRfb+GvXSuhEZwR/euS8n3vx3AqHlrb9hntLfih5hSFDc0S6JQeznBm5/
98yLNtxMV2JzSfsfcGilZlLcUn80iDTsrvH4x3HUulSOrbX+Sidx7ZhLQvVDfqjxdVSBFE904kLf
INcaNwYCcKLaoxgSDWODjgNYwjRjw8bq0j47J3rJTyuRcQYq27OTTFRj6S2QVlGA7QGl3+m/xTMt
qd4yDuOJhnJtlsjwHvsClz3TmYUd4jDOe3ux/tvT7DmpNdnm4P0NNSnPO/hIgI97eIzDhkPRx/NB
NFqRtYV0iOKqIVmypzl96F/iPpXrK71EQ8ukEPvYjh+xxB4r5GwtFiKTam6BJzEaa5yk0/wdByTE
9/aboCLl1B2AiZCvzB1xBAzCIBQfmgqCVw/lp6GblCoK3emqAsEVEDNhvPqsVt9ahF8Sg0yL9Ytj
6KmcP+pMPGSGeiHFps6HB57+sXF1ftnzu1VqqMdkbHk5OgeR2tcFM03gzBOs6Pus4qLkCWm99dkJ
1+KXAKw1ZVqjpMsOKUGQFX8y1Ozs2cZbbvBdVUuTzTfT3tsY4Ln1RYrtjjKSXZ0AUiNtFdgpLvzF
6iiQ/kvVxjRt+Eo4aUYna410zp6CYyFMP3qAbuITghL4+BApQlU3J5AsLn0M+pr64nmFfybUhu0C
HpP7vaYBXEtfQkIHzZYg99V1kRagcfofzkpy7VLFhX4gOSvRLcq99qUgPaAR3eNzshZS+0Y/iF4+
30YLG3JOXDGgoDPiIz4IJLbmzMVObugbh6jV2Ya0Z8NADJEEBCc5RAfKG2A3wcWyKI4KSxpidE6i
BwyIl6jMG80UVAok5wmqcpn6PK8rInTvguzpiiZFa50haIgcfyJitpqGo/nRG20dOC1Elv68jZnP
nQjZMIE08vmMxICX5nFfcJU32R+qWG7nKlq8A1CEFISLlVup3RVveBv7BZ2WEDFgR+FvKlhpAyue
JRDZ66aEPbAgvmu1/1K9js2CyIw+cstWisAGONeaHb0GHXKT07DFu0Uv/9GnfBlVAVVYyfLBnaMK
seByB07ln0St7xqSMkSt4OzfJJvJeuTen2SXkU7q9y5AOHb+1fHJmNuEsUtnrN/+bayzbbcARZLm
Mdq0ZNcd+37QFHwY81Xn1XINtrLoqrdwN+hGDVYOcWqGaQCg5vVfa4UgBLPTQDXvVNVFpEtVE9la
ElN8g/VxVzMHkDCFtgxmtmkui0cAZi8YmNzaHHiuRPmB2mbB9JmHlbbWn2todZ7yXnc+rmKnBTNf
lyyf10A7ABan42OFAsZVD5Z7Ue4qXNg54Ampqa0Ts+2QqkjMjRb14l5BD00kaO84GB17hMW/cdCc
sHuAgJpyYDICLOs/NoX6RbX+RStknFaZBZ2SBmt4Axvs2aZl80T2tj8+fJoty09tYpUs8WqabvYn
b/KclXTcaASt77MXOrq6K/E19DDdzjERNF04CIPYS8J6cQLdR0bNU1M2+G7ORtIejlUEaKSJVIk4
lWwHna8xR0kDp6WjMkb6G1vM+j4SpeqMuNchwcRSTWhSlNk5KiE/kRXHqNyaq7A9x/fKqwRaU99U
TEMWrP/F6cHaVyZMddInEyAl37HTK/pxMDCzRo7IeqiFwXHW5GYQN2tWWgIoYcDrErFUAFBB4wCP
8B6SACO2lBjfQQReRT4eVhjvcQTwmQ0DvOYoVuGR5XnEt3YdQSKUFet1WzgI3Kl5wEPsq3aMsSDH
iN4P6G2KetYevYbK22TPifyH4iucvTH7QyqUbP6MvqGU4Lc2ZSnFKFRBIPSi61AUCu8rVGXJPe0R
MBYlIrfoBidwr9GiD+s9Q/QyvnqKJMCva+efoTktRKIYPeGujNB9pVLOxlW2MIl6D1BPWaYqLf9f
/VMbvuZcmZz6R3HH3NIMvvBMqMFwWy9v2JYwm9SbS06455IQ/Z+N9+RzpSZhEkaZ9N47nV9R/zOe
0IMqPEPxH7gH6ApGb8na4iGroZTZrGxtIGWbhgwiMiQY9pr1s9FMq1C1VVYyVtw7xXat8CyRLzEs
lWx0uSZYm5+J00GRf9vp7zrkU4RDlqPTyiPTefOqeklBsCfVQOb4VfGagf9dqWLsFOFyZU56Rgbp
P2YjQbAdA6cDQajWcnqe5kQJ7a/5Oi9QbBVxIG5tS2FqaFj49+8Tg0ur3W4mdSxGsSjujMHxeSYf
Ljxc8y48X3HM/Tnt33SKMvKRbnEY+OwOaIkZzEcj8k9JyrxAwYgHNzJVNMd1K3m8saeT/mWDPs22
MIpxmxB2AgSO4moxIQHNq0BdIjHGJuj+J+HJJXMzKJuNeHBsS4MQbl8rXU+HRVwdu5vchAGHe4fF
jBVSsiHxIcPRIk58ig0gPXdwyRv3hTuwTwIF6hEbQDtlxPniZdf0JHGSxd8+BsxdSsfK74w6GZiC
e9Lx526om95Jd7jGUERjv5MQMZ2dNNYOC5ldfeqcADesrgr2rBhEBhf7ejhjeUoeLq1TSR+2nBZD
zw9Wgc3Nnm4R/oNWcTkelssp5rbQgFnhGXpwxpSuxXXB+yrb9+7O/23mr65QtQjBhP9sgowSH0yv
uTeKVOl16BULJje12qdq9emulrES66J6U3RmZ/jUQ9+C6xVm3kJiBLaUfL6pQWScvKNmz2m2vyQd
10fGBTi1/V3Ne4GDw4/nciR7owo+Fur1P+t13jUsrhhf4YLtNXFY62pQb4AcOb1nhTb3xUjAiyjY
WkRFM+mHjHeaq0XrnKfo3bbxEAe6g/gQ+CgR9uNaOo/1+ScrkJ9OLNqMT83IWehWC5noBOX8RBcA
ARePdYcMzwed9wPj4DaJvX8PTR+2/3fmQDo1LJoJGvbOO7WUJmdMCIwrN3NjOUb7YasgEMqvuAeQ
ACnaZ9/TIYYKMjdvYCrkL5H5mWO5FG9sMCr5lvLDUx9LBulSaPZDM0KySUnMZLvFztTS/Dj1oIcO
uMvfi1MwTqyjd2c3zaFliwu5/EmDRs3vWEDirW3J0/hoPjQCcYieWIaVKmV7mCYjhHMdnt+NALz0
kmV7sH7ojBr6Ft81H47fIOunw97BXxzoiIxrIz+Sw/TUkjeh1qks8TyXhxGWfP5sJuZMgbVZ44dw
K34aVZcK800lw0rp8rnYwaG+fwQ35EgsHUmOlrrxm81nXveGF3Bn4JzJJ8iS9FOwxACVhdjvsOtl
Wkng8bBhhWTVf3Hew8olAV4wqO5ObnFX27vdzOJ4fOOlEph44kjVrcHIDtTCydQ0dST1EdtI8RQd
OLief0ml0dQyZBbKcCKsS2kbRr5X5dU877pwR2Cf3QH5aXKOCCAVaZ2/8KAnT1+WR7MSfjikQM9z
vACs9xD368vo2M0Is7p0Vw2952YimgAtDJAeXRJzo474N4cLEvAl1yKi3qpE9U4p3ncirBr0j7Bw
NC/kFuEwW6UUUe9goHuvbVx1SsawY/rSerK9/ZffP9Asw1gsDE0UwZUoJZ7o+Xk9K+sywzqnEjxC
6B9kM3CjHgHLxXghuloVcHTl5Yne5MLKJ1YQqIANvef28hNkev0j8I9eIRAx/jF6fAxvIkh8r0X9
BIhHvEDbIO0ssxUTDFiMLlhOCKEH8jolQKxpfJTWD5Ko0kRH7ww6DSNrSKpbX20JlUSJ812khBW4
Ihu7GuUQIHHR2HfHh8yPKBShqeEHExPq+0biPCItLecWvQxA+4fpekhhfYLIVaiLAZLL2ihFk+l1
WDWH7VoEq9X/HWXjeH8RXaNt4t3PjmEj+hzGrkkSETifHHQIZfE8G8y4C2BS0H9lc0GowXDvgNHn
BpCXQYq8grMq3FdbI9xGfm3wXkYlwurQeT2TCEReWU9DQMi3yzMa3wouu2FkFHIx6r8n0A8FdZs+
DM/7ZqUwwZbMMTicKBwXR21GJLEUPxUANi3f1bsGg/2/davzTtLJJ1NDVPKY8F25ICdInqJx0nXr
wrY90Db5buRR1Ng5Ygk3n/tSU4IoaNI7A5XdWreKewxWqQIE1Jc4QD6TSCIMWswqaNmhfPo/NRwN
p89qYLVxq/ElRYPWXWym76kfVct9fUmc6crYw8KhQW9T49Mk3iQ61QA7hEYEvE8yLhEspH2Dop3F
sO/KXL6mGoVjRbAdk0r5cny6hqO3qNrwcaflOmiOYg4hVhoSFqyERXmTOlyjSXwCSIWcWzgN8HU9
1Iw5LzvSQWKsLzmP+kmSn112PiToSuFuQY1loyDJXJtiJCE0u2OY41YOo/F7QARkows5kPYlMgNe
35zXzOC/sYyCUPwhGjtkI+YKeCUcA+7FZvqfJ3xsTPv5uGXliUaWFixOZiECzIBKyqP+idVBkusC
aq7YVolvcEnjYBasZ03LQzKj17r5mWxPL+rafLori61L8buGPgUAy97O0bX0+g9/Z+8DSQxAJEmK
R50PM4o1UFjk6Jo1NexZq8H+9JulwuTDuIV0S7wiflgRSUXBapCEWc1T31fDznREQeyqEY9iqv19
Ab6zIRBjLE2splxpgxOpI+UunLy3df2t06NSK4oIxmfE3V8gKiWmUBLaOSE/il/t1Alz7RePByPU
9DbvND4MpwBDV8sG3gJlh5KyQIIBxWxFyAnn0J8wPFtFUnCIZKFWSyglme9W29YvoSoDO+EGRznq
rdtqFi7qMQVg5b32g0SAiLAfjKQcWith1abjOnnBq0FIm4JavAjwHxmasitscDKnj1JpDlQXublb
YDscrVj3jNE1qx0pwlXhMclnx1w0/1ry2jl8+ZF5APbDFtJ4VWRpLjOYdUl/ZDZImApl5pLGY1aI
nYInLpG3aW/4NL3SeqdercnfmvbqTBRolbrz/PytMnfovRHwVnVnrHn/L+B00wlgvIaO2l7Y28iz
VZVZLHueW6svdqw+poVlm+b9f+yUYEoMgfTuaG4JsIKe6DXJRtK27KbViNwv6j8bMJ3SvjnrlmGQ
VrbOxoGSk5sMg8AIti9TFut9sTsmwB1Axg1lkw3v+2fGDneAuxVZdpRAeEPj0WdCXF0PU6s0N8KM
4Dmi9SscQmtP5BmLqOyjme5xoQVl6vQD2FEGTM1GvGe0iyRnWDZ3R/fN8xRhGeYHDk9b8zKkn/W0
cS5C6Nv3Td3DAzTpfRecGVeTi9mH2H1B5Fu0EghkQS9hvW3dTxYlPX0ThQlzB4iJWYaT6Iy53tfJ
q4Yzo1qiyaTL+10lenlm92hatiiTIzDO4fV3xWfRINZYWBjrPSG6cg7juxtsfxL56EP2bc/socp8
3CLai4E6h12gxc62ryN5zsCHay/RIU0wW+A/HE2kIhmSIWuKh0dNmOZryQ6GrnTbQBYBNR2hemE6
kI3PZAqGeMDUIMj58P9lohGc4YeLBz6A4EkYErKNCKdv/Q7ciCaQOIsZ+VkU/JcOFx5+QNIvNeAL
YwehHyZpRvX/9rgSsibjnTwltCqEplesZkdczJAiMmplnoc4gx6/IauK0lv9s/R/U/Y84h/iuYCv
fpspc17ZqguElLOOvn+Pu9XuNwSpKnjTgS7gYLXFnVg6cH5Dwn/wlr2j5FeqH525J62LBpPOoL1V
tRlIJLLh2xa1CXVf2ByHQqUZt3HjrHaGThV9w/NGLaNwKyLqwDPafl3RKzfBThDLUJgm6djLIL26
DJD19MCDrgxyPNLNtUthvXzyl/v9MhBsGaoUw02a2Lpx1VC1b9swDXPuoDLZqGDfY2yz9b5bQqPw
v1BxsR9aSWHXr/HJhFuKGOCs5Ob2WAjZ7MEFcTgYUotwLMi0q4tpjBrX3m5tqijS9w1Drnvc/Gwd
WeZS5FVSykH993Qpqup7iCxOUT86bDH4Zs9Y7sq+0jCKV67xpDzagkb+Rnx1+5w2q0yQjH6roUqg
1bk3g/o+AmeRs9r8eLx5GztPahkav6H8ZSzfWOsurMg+w4dI9wKmbOJr+fPdeo1kK9SNKQqS7XbU
a7scupHiPaWb3T663Abmbiogo19k8/EzqBVi9/k8759ReZ4ASu96n9R0YDPXvKUyByJYbsbAme3/
+/tb3JLKs/kh7FniOcgxI6IdftgmI/jRYbu1cUHW4+z4Nve8QkXDkAmnDldt89izJLuNm4ksutV6
ES+4nQ8U5L2TqAVJIDlG4ClIXF58prFEy9+XFto/L3xdRS4tJARkzizgRntVFPWRHuGBnyjJuTV5
RD4+xZJSk3QTbYadKrhHW+dsTJreTADyoMORlg6Eh9zW9LrXEqFdchy7wHmunPvpm0jdSUadJTtG
ynO+uCC2vXH67pAkkEQjT620qSm2qJv9QD1k6HrK4rAAtujNK4ZzSBPiNydkUFbwBkadEO8FEzfW
4/Ft+sFXEoZ1a7RVsB/rL1+e42Xb6X89tplE/CoPfdF2YTY9lh8iFW9KjiTrBNdZC5m7yHs6DFmX
0TKau8eOE4GpkaNnAWYUJSWjSOtS9s+UbhFN3CKvdN4BRjHaF/a1Fcnv/ohwcuVxqOo9w9vk5zxK
O0KowhV4O//wGSGJTEcrtCis1N7G+ZWYyB8m3+NgG2gAH6BQF24T3Q8Lag7kxaRWxCnwh2yWnx15
45PCMVuv/95qzqiYSeN9PUz/GiY/NYxnjg4ntJKotDW69vxFr0bJzUmOsLV1P73ByYgTR8g286IS
MVeDvGwn0gzw1N59hmjg498c+7HstfuYgrWbU102ig/lLKztJ16ruBwrszgcA10kKg+kumOvPVWK
g+/e81MLWtTZsNIckeBn9/a7WXwwwQHV0ET9vBVd7UhktU7OmMTO7aQc/7wOMCJ9leQHYQYWR9Y3
+uJclSgzByPoI69FWfiD4cGkQrVouklkjVcYxtIGoRJ44RKl51fYVe1WQvwbHr8M0FB04SbFsa70
kU2hQbZUjZ7O7tCCy8nhkNrAf55YyJeKnr5o7jFAp7EGnqMeBi4ihS7ioiFQ7l10tqW45lwYYWoY
4qMma/ucjG/P+9w9GxE1Y+6naAGUHrsW5AVJtowiGnL5sRbZjGZ4rzjXiGmKFRUzfYUvZZKLM7xQ
2ONUVJGaLYB5RzklJo4Uf//b0tW9eC0AwEUW167n6Nnzt5AIGg5mNWzfMeDcCLGqOGv4TKEzpROf
0oV+OUNPE/2AXwA/jTT5yPowNn72QWHRYHrGVIrZqgGKlnUmmEj5ZnTFR5C+I1Qg3vpiXMvbPkY8
ed1dXbQZdz0mExfMJUPqp48RDgtSH4YuPYhJL2zkFk0O7lH49STK43cEPfFEWL16mXYn8nWV/WoV
VIotRCwof+4Fhk7ShV0kfHa0nv3ONq0jY4M2dERnUieido0E3gnWofoG/iqk4pI64VyD4qmjGrIb
FFxs9hhand+htewxlSoN60Lv5+IHy3tpMfEf6z28XwJAtVg9Y9qYepvnXydbPfO/+sQy57kjAdez
l8YAhMwestrZ9Is7t0WzSPugsQV1/7TW8+slPW5Xr9syr7IAGxOO0xxd0U61MbOagzDgPcL+OvKq
G4Y4RS6YF2N2cCvR5n3p5HgEiFwxQHnHggJSyGEdiIhkb8BLuJdzKBRVSSj5ki+o+Cv7eja5PfIr
G4NTyTjwpCd0JHzxPJqIxBxpyuYWoQCLjvIUwJufcflvGzbQ7VRxAW9E/srhedNH5QE58TO/ygEW
JAOgXgKQdWvIyoQyKN9CHfWUOKqkUNAB1Jz411ed0L1VaGL9aUxJSA3BMHPwWSu7V2MDRDTLVDMA
ihEUr+GAL3odZxBB7Esb1FL7YOgNIYizEgCz5pIF8vNfM/WJKYTdO8U6K3pdN4M/e6vT/CcGy0qV
yvR94LyDoeKL+06QiPBX+cCxllHUzdjLCkEtK5ILdPcE6VsPsl681BklROHhCMgBL6L5x7zejOTu
X0vm9Yar6p/XdaXfQ4o69fdCbDSJG2ZZfon0z6NIWqlnd83/m4b4TVnFyxebHtJ88DRQWEQ1z+BS
Da1fFezbUINCFB99N5hxcCWBZ8N7NACnKhjIyRhl7nN+LBe2DzQx6QUJzC4fzFg7mFuHlxrstNQT
jftlyN95O6y/rvMcDucAkXUpscNFPQ1dI3TWbpOH+3TatGUx3uFeinrKIjj3etY9LOEBItt20Ygx
yOL/Xfac6lCB7brQH4CeCeEJsdYWEVcCjI1eN2pUgvI981T8I8jd3k1jAQd71LU2dyCtzGxT7Mvb
1GI0jlGX0Wqodgq7f3YuyAF8i9tjkwuar6ibaeFkURjVvbPHsGRL7ru0q4FbK/KGtsBNi0lFH7iH
2bqnj/uba2s+nfyVuyygbuk9b2xlatNx9X8gtdL4+ZUM5eYEnUBDrr3Ee36MUK2OtVv9I9H560ru
ud5C9a0DTB0mCLGneUfjoOF+04eX8DS2hSxYvlY8Zrt4zmnLjuw+yM6lJF7hwrlZkd8EY1eyihtT
g4OCBLFJShsLmNKqOBKUqhoTFWABQkAHH+1shrGdbsyw/xcE+Sl+cIH4lsdIBm6kJWnib90vrRSC
BCKoE2FunoJo77LEghUwkjqiQdqleDHi3ZA+oXAv5EBBAB5PmgXgmiKYUc8lsIiwhEJXzrN4haqe
gDq5Muh0YiMVlCZNxnIf29yocSbDqyxgzFXS1T9NUuZwk9dknZuBqpSb2O3f7Ge7UJrJl8fZwIPi
VnZwTrtg1yAbS4Vvlc/dYZiPj0jWBjZoccIfAbu1fz5b3xZu1P+zcN5Ql0geoveDLsmlxPxYU8Kn
n+jejzwKEWxcPght33Ai9eiohfSe/7jlkwgkZ2d4i9auTNKWJi/B4RaIer3p+t2ke5Hsi/hw2qDL
yoxcMNwYzSAf15/RbGHE5USuBo9Ovh3WXnsO3QMjXywa5OtGtf/oPwDRLmX4u/VQHNccycz/adiE
vPELPogTergvi4OTSA/bwEjizLJsW4db7At70mGPd0sEtEULLTICuEZyGiFpXNZW2JbaOzVvuElh
UPQX2GZGVKQkjyf6qJJXrAfQtp5ItLMUVouM+qMvy6DHHanLWgKCw+EmOYbQKwzl9wMmsZnFf1yk
BQLPB10bYqY3/wpHkBe3EG5Upfo9bbox/Jgp1mjGa5aJ3ZHH6j4M0Om+6K9yqCnBSvt/E8FwsXY0
r9zTKmf0ShOR0iT9E7gdMIT6pF71ZeCSpFZPB0PbLW5HRzW4dsuxd++sXuuiqz352Z48cMbDAs/X
PqrE1dk3TahU8oLgf5bWY6ppaGcyYE6CO8U9xRxcLbrjEK8xk/KS/TGDYaivCuStLQqG7Dvl8+EJ
ctH8OtYw+5uKLc7lC95DkHH/2UuR1rMmVqjX5ZHfJ+BJOJ9ZAKJb75l8H/IosU2Y08K6lnbWEFMe
tCA7cHwNOI/uKobXkfRmLqiKmpjCHA/YrEmd7CW/2RwRG1gcdLQ27JHnMJM2lK6gIfuq2+pDvhoC
zLNL9zUtotLUCSPEvNgYyeHlSpG2kaVFc8tzSELDDj9FxmvPcOvMxhoYIHrJ/dGf7Fwn3AZUnUix
NP16LKeFm6mV8NcWHwSaj9qPA7a6owONu3LxeY3q8dVUe6s8xe9LUlf2FxoamDfF7MGHsVoqA1L1
v0xPErrD9h6OXeQl/IXiQtAl4r/o136OolXTxFwT24wV/i3EJq+A/SYhuomyqtJyIkgT5Rm0I6Za
a0x2f71SkR0X/9lYjLkDM6t4bCuFXrd66Ctql5Qwatfs1f/juDjmMUsqVCQYltViEnxwRQspgh0y
BVCehBhJny2+BuMS1YX8kSIDifzV2BWCleXEdSFxDUHAKSTkBGr0XxOyHzzMay5LpibsmJj3/k5P
Gj9UO5ALGYpCD7d0ulJ5NHgd3xKS0RuAdpuwMWiVqoKRge93Ai/iZ+T0sILB+J6CMPs/PBqpgtgV
k8wtAiiGRWdB7OUml2XIPq3rqWW51OFJbiyyB+oYleJ2aJktcZklFSjLJRI6MnCrWw1W+Xbsir6Q
ZoV5erHJbeSySXYK9f5JhQsnHeTUhZGIyStje+KVZxNkRjt9SQchk9n6WDXbj2kORcJqnjMruFql
hNBY8YgvjjVt+Vplzkw9MaNLUf/4TlT8vvi+8yYvA64k5Ko4oJdNCeM0jl9XQMm7VBxkoZbISfC+
HCTtsohFktrcYLhYPvchjff04yRTtmo5m3CIkAkck0B03/2QQ2EReFiwPx/9CW1m6WPU5M3OUiwA
XxSHICh+PnS0T7u1DXjNWojTraHdqGa1xy5zF1uYU1Lydvz5GzbNtllzHWHIMElyML1NfUoRNSUz
qToLOf/rK1hxbVAhRA8UJcgwIrPXDAo7kK2AixMMOJ8JLNieHKx+ALCH3Jwy8pQVEopN0X1FmeTB
SIHGLKWyIFs51L8lHFxWZzega4jLkaFSK9A0N4M95wA1MkJtKWfwPRv0x5XumaXrywWnSxJVDOJb
7oXEkG0AnKNKb+W26Zv/4P1sQ/eIVi8pbVnl3QfK6IIcGVWZbq7IhRNksP8bw6QEIafN+AKhAeAB
jLIpeX8aAIqWt2BYYQrlgFyVwPcbbnQF+bnBg58u8Lft4kNM7JAL4T04yxoWAvOFsUAZstvVUg1C
aIBXBQ2WzRcYxCEYf+gijUQ0qmXEkDGQpoQDjJECKAKR0h176jAbfzwo456Hn/cqMgdzkGaze16P
xSmQAnW+jJRgmEZvMdiD6snjF21XGWRTWkL+ma/zMV4D7qDU1YY/4h3zoU2J3ppkwWUgDAenoOVB
bBnBsnJwu+APjs1VgQGgbpfphOWwjfRRjDhwYkZbhikc1GnNXGBSMBTs9bk1P3bpod9hQeU1J+do
sHB7R1pDrPF/g8yag/tfa1w/Q3hDsXqoqBn6K8B37rF++McSsQ/9gRMWmvGcSM6tU9CVF9W7Oa/1
u5KdgGl4JsnufBpCBy1CpXITGY0g8+q3PtU3tyGGmoGvQBGvjyGbBnPiTvrWFkvARNHY3SRUMIjj
5/lWCKzbH+z4gSQP1XTFcNpakcjKOUiFhlEwSjcV+9FF0lOgtrgHm3h8+hcOi+CYRA0mGrjYyly6
t98KS99jUKQ6x8EU6Qhkq8GIG186RGbf974nmsOWWLBWLs7OCzIX8u+ABEdCtAfsMsyy6digX+H7
+YWrBTuP/C8EeEWKpVY/i7lQ+bcqXHbQlsR/dnR2rMDbXehFi/yk59rZvuFGoPC1lOsow9ucZj3v
e0YvhTnVXH85lGtWeYpByaIDDxS7FBZ1YigAMnyt9NA4/M34IpHlcujPEt9LRubwtOCrwdyY+7a3
R1x/PoUHrZoVJUEQNnF4779t0SppDiad9oZXOlkVCvHsWtGjDArvBuojPSTmAUKVbVN9JzLUQec8
7PbaIznQenLAECADd8ml6r74mAH3hcQul+Uj6a07sDVjhRAdjLqhDtffqCCDyIEJ/Q7f6DGQw/H1
L1J41vRKIn2unUiY9gCYVLY7fNK1bMLCl/SjfeTJIWr4lCOopfMF6qoh1Popr2G4Sw7r2koqL++4
0hlA2JlXgAxmZQzF5DVhaTgTn8r+z6UxjGL4SmBGMDXxyNdln30aj89F6KoeSLQwmPfD+l3R7wvN
TKKG+OpRrNkgjsJdQLn7u+JojpElZ8FkzwRklDIcIGZF4D91A8k6vajxYUcKQq5ZWBIFD2sNtuwW
+5eimt88LUHUIjfJAjBoGuDMcIg3tFQJZfcWi/gKkIsduHvIbNto6iWcvdZwtg9bFLQpt2zlvC+I
brph/IzKmCZAQbQUT8VKJ96MINu9o0QnVS0bGqsRBJ7I3VRFWmJ05pGY8asB/qay7M5b+S+0cS/f
XkzIl18GucqrefdDz8tJx2wiIv7pzPdW7B5isMQZTcuDJcb5A7u9nt1JQnGov8cloDt4IxU9llY+
d6RYUEfqqj4qOb9qqlHQ4AurHP2ZpgCRmF2FZU13dghaW669hJPM06QCD3z28C6aEV3cFU6ei1TS
FoP0IvHKirslvr52xTJbXZ1XKYt4hkwQG5Jx5AaSWDqXwn5v3deVNy2v+bneYqmF7mKRWpvThM2B
gxjMHiSX/9TPyFOo6apV9vGYbFDE+cDFvWLFqRZZsA2Y4JcY62b1l063Yv2DjC9NTiNt2VPErMAu
SpFQAO+OVQs9Xg1JEhGh2IhhyhYp8uCsrNJHIvBWDExuGbUe4DLJ9B6YBhUk2bNZXaHroKwS6mWL
lvXrGDNkFf6Dc+s4TG8i9rrIcZSTWM0SqBs5iBAQ1gkfRI8NTOktJAo0kr+lha5b/+Xajs1Z9QRg
+OO4X2qWbd8DyGKafhxX/tO4AIn7a106wQvm8VKQpf5xNTCqOS95suC5kNFOwprWSrS42uluAE4P
v0dt3ZtExzKQNbwvx+0ScXvp40deIvYnTuI0yg4/8N0RZT1QY+nyV7anqxvY/KwX8qev2nVhxejq
9/rsAQIg/ZSrcZ7i38pMFxAQVOonKUZxmTBbOw2q868K7pHRcaqYNffEiEnd58e6xEleHsPj+eMO
0ES9D2nxHv0KvtWHCTWro+M2DunFhR0nEJe0Y9fmhmdkmIcKPPjsIYpu6XxOXJaKyufjm6ULQSLR
FmUfglau2SXK7QhmySHOKDLnSzy5vi2ON70dWNb8VNoRn6VNfnXBVVGh3fc8GguVGxp/5gcM9f/I
QleiR5j6JVUmqqZWilvsDgfWHGPyFwQOvjy8pvZV2WQO6T6RySu2wN38GO5UsZQ3ECNEVUbABZRl
oFiil2kOm7Niy90tCZDEVhaRl86hcUfarmY84zTEmAucUtxJXeKyQlZjdcQp6RIJgN0I6c0vE0s4
7gpYPLSOm3uW0Ykf9uv3t6E0OvSfprWKLINOVxRUC4mDylxY2g35zTVDDXoI6wA3mqM+Pnaxu4ww
FjEfUImr5cVHzI+uDVCkF9kKxoRvJLvaP+kNBwr+yKg2G63I8KJ8ALQK4jmVoxgOMZv+WIj4D204
tS/ymTtTj0dyVDnd172amqaLZ55pgWlRYWMcarYU+4FG3HQ28FwVEZfxE+BOaPUnJ+6ZpAkGWHSn
/k37b2XoNgDZD1hcdn6o6q672ZpjDzsEPp6K0d3rRZFEN4Q3p1tdfuoju6iEGr/IaMM/03Nqh7I/
36iSVu9mXBzH27Lrx1fIZ82meL1I/Id986qAZD3uq6+ezZWEoziHYunPvQwj8+dSy5cNL5Ci1DR4
gGbNSweKmqi2Lo9+JlWuAoaCWYG8/4Ez/8dDc6THAgNiHs9PUHOnI8BVOofFKQMgoCwxp2nBy5gv
TWXcEex8rWXNfy7xyxPFFhTw3tUhbOMblMQiCqpmGvJhB5pHGH7XFW6cbRStQhk68jq4Kl8CEmx1
N+ALEi9mRoIJ8fcVDtsDrSS0hSEaf9HT5aIOFMXSkYsU59fq+HjA6HEzvAudRGedMdAp9OE0valR
Bume2QCQWnD9mOwfFWXnypF0KbGUcEmuNB/WVvLiab0570MkLt6bSsrRH5M89v4XSs1dE673FRqb
yppbzJXGXOuqU+yplmQmr11KCTgV+l9jSD+d0Eyu4ROnXtjjySWbE2P11Fhzu9qBCZgacfRglwEZ
Hq0T+a9wisEKl5BPBX3JJkBCMiOQBs/ZbBUpDDlKD5qHU4/6zZQv0vAlGcOH9uDWbYzCca184eDW
HZkgmGaKzPct3fF2w89OD5KZ2Z6eQU1Vn+ptLz5nGzZgXOo0CMn3078y5yJQaXTHDEMvkEj2B3yE
1o9utBWGRKvuaQ8WZN2ZxXJZRJPb0iclfzPMxyqW/TSA8aXGnrtVaimWPF5dN2FoYDgr8ZJ9Dp2f
hGQ42hlYOHiTBSRzhz8791baHvXlt6VzSIvCGPxEjADBhotBmtRjwqraeC6WLeIfy/LZjasI247+
FABnb4Qh0rtjuuTJfQ4HrSqnLE4Y2BVQXp3Oeskqstt+QTsXUSwE7UauY5GXx/IHwhfclisyj2qR
IT0C0H8WH8wFx/ZYz7YYoBYSCch+X9tmtXag/4CGy0Q48fDmuljTV9oaYFncSjCuQ8nZi70OkzKd
FcSHiSqg1yvadiMiZHZdwpgw4xEv/m2BLjL+59X344JNq/9LKGyjKICe1DkvsJmuB9UxfLl0tpAs
4iG3HLZaZlWrkOjc85FSKkp67BHxsdqmweJMC/QILa0TrNGhoWVAv5IgDzhUd5JqOECxpj0Qxyqg
Xn35XB9jC17hyeWWFQ776lYo5eJpKlS7+FrfuOHhYVOneDhmbs/42wx0MGTh0+UV9GtpBtsMyBcm
+82myVwDlZH77uRl/ZSOPyh1j/1LJRn7A8IZq3sQc0Rw+URqpopZTXVrpYSn8I/Ncc+6maM3xlqz
sg2hcwGfsOvfdLcUW5bSL7erdKZlJwZuCPSlGIsRX9P7X8ikRYzEGSbGcQklnWlXb7RpaewK8MYi
xBGpinq+TL1/yzrQuutim6vXUnMgsdx4tSPGRs2YggvSoYwc5TwGivTpPUnlB6w/yXuKSumdYRZo
BNpPA08IOA0tq/hNMlLo+Yy3fEu5ft5Niypo4vGvrdH7+sOXHqJb7j2yq10ZfKG2Dnm883/FtIH9
UC/Vko62T8mQmwXofnRNQkJNCpFPPKJfZmklBdp6c9g47yBsSWSCZwacrVPSc8P3B2P2gjuCDov2
op0w+3o4gSz3ES6bjLjpFwb7DSHVWgWhNuNNBs1hBKYfC1bCuWx17F+y09yn2yXSrTV+dBk+grp+
fRPqABPOmWjEtKls3/xFgm1uUOJXHbwK+fM9L8MtLvBcx9lG5DeHGwdeQ4JrCq4apIlGI+gl7SrS
OBVVsqhc1bPguPcKkxbbcPwa9wHYA3IvqyHEeYimy182ghK/+xtg27UW13zvChU77w5ikhwat0fA
HsiI+j43e9lSUrPxJi5bojquDZwe45Hn2YX++M/IE9o0YNtKh5HyWUgQvuPcRRIlWBV6Xyqp0zck
NRk+yQO/I8zoygEkHoFjYB+wdXrDXtBifKRmX5EzlSAXnab3a674Wj9aEHMr6+dAFK3ZGRTPofkE
ceSF7YAZrR+s8rC9PfrfHNGxjmDPQKr6esM/r4spM3OErY2Z5EFlyF2GHGsiK4jd0OKQ5CHAXdqj
YNT9MRJoxQ2z4Vce29bk+fL5zRtceGgonRFkj3h48IByxK6B12X8WFL3Oo6rUs2ltF5396NzTXh1
z8lRd5A/4wgeqyvvERMiHbswp0XYiTVazEgQK9YpC+srcxDVLxUipQoDy6ZG5I34zjeAhRqGALwK
54YljXtwuKJN5smcukTQ6lQvIV8cG+j34poo0NgotOPXbhoh+u09CJ6kyVh4YhKeQw2H7sF7Y6hs
JKie4W32gEnj/dbBiU7/K/IDbUq5veP/QegGRhYfKfooQWJXBEccYU0cNk2UZJKJofZfzjrI8xxo
RqKpEBZptvzGW+eP+cTQgND2os0jy/1fzHWAEK2N/bK3CIy/thjNGCF0ORSYy8jtCKcl8tQA6yJ4
MyCRIPC6KEFFqEsPSjf+lmD+6UztXmkGs7Nf64p2rajBWcN2fmmhms93GLuYiXVdp/2iuNhdxiMR
wBnjjqjCMthxPDmAiQpewr/Y66l0NbJxsWrEnPm5ng6xY92czn5FSFcNUI/1F+IwCA4enPHMxHC/
yFPojNRhgaVv4AwUsxcnDO2QPH6N0TZjuj3Kz5pG+bLRCp0Ad2mcKqgr/w9qghbd13+8m203ZnYK
8Wr5xXHbRi0Cma7g5ptnJZQMTKx4Fmz1tg6tWDjo9wbv17K6I4rhKybPZUtePjowlUpIGYQu0APp
30ynDXYobEKdHub8R0E/XhhZOhfm6+U3dPwYMmlJcjzNHfN25kNhHXqi6XofD4ubb6GR0NeORjbS
O/YqHpLQBKAI5mRErEGcEUFCzXhPxK58ZvNI0t+/uQMTMkF7fS0K5YBicEGCyieJE4Nl6pgBWuB4
FRxNbHU2VdnIJFpCofXZsKpqRIKpDjlQ0PvBEkQL0/xWqOLyxSQRQ8QZGHOQQZ7ZvLnbzuyO56vP
roAsSMGtqhY2y+6uNr8+kKYeZnlC/Eh1euBsLV5TpaYk+qO7+Mfh9DSVFMO19mZCjwWyZkB8hqUm
ISE2cxHM7XCzVxHitDrbEl4tXHDBEd0fXxdQ7oG+tPzCJC0dTHvGKifylyz4cpkofAlf7IzU6uXq
Jk6yg368ZfchaXBawR/hcAfSF12EFGnD7ePrKza0ZBJY/Eo6smgCFW32dyorti++sgeeWoTG+nHX
k7dVVLM1Unhl5hZJvxmkGVPS+R0yAAz2cYMDw6WqAHGUh2tKxnTl+HScm/IbpnkugPjwSYd97O3P
rR4OC0WZDHRTG8J8XCEJWbH4sCZHQ0pQbdgreNZGzxyq+hv/goYuEQquCNZ6zF0xVNZZAKiNFuZf
hA5TH5r7Afr1dra3YlmL0AORodpPWZTUHDI4UpLO+qgoom25WyEBjR5fNa9El/OlqStrVJxqSVD2
vC/W9dV5xropOLvajT1KWVqvuaugXPXWO188U6dQOgpiVzVrPcjMcIJVd7flsNK9Y7B2lVQHrdpV
y3zRPCx0Y+rpWJRKFG0LphrLZ85q1eJMi4PyHQum7ixMPUjz3+XxTkBCxMn+Ciw20QJePTHOmHzn
XnPfNYnrFPsV/x0ChcSh0jAW3ORna4iSbK10zK5Sc8dR6gZ5U3tLT5Vl9SP5xubhPRgT/C9d0r+D
qE5FXVb6J6Xakr62o5MD48gHem7m7G8hw+LU5UyCPCCBFnP5kfd0LVT8DvJxRPYthMfgMyYsJXCE
1tK0MljJJHDT+XbXpRh6HeCHStT4yZi7/h1TOJpbIOWoc1NvnHkOxO/LwYMNIeNDxDqLG0yfRXR9
bQClN2vs3q/tsXDKyRM4VFUWMqk8EjKY2ue5jZpCnasEa1WvrLEFpBWCM0jOE6Lyvwo+mTnhiwrL
sTwplJuqgv4o4g/BiwkZLW9GnxbFcYDMV3guuAxykDIRFzAiq5VOLC2XDb7AV665c/I6ZYdbWOLR
gpN889ekdrjoZ3R1gVT5E/Q4ck40QsPvv+K38BpIjZ6MgjJNuc7Zsc9nqRjFn8yfLzDyni3+bOtH
7/1kyjOS/d7xGVBzUxlDOOOuNXzhJefZXxSCvMTz4hJOKAxcKQE/kLpJZiXa11+6RhiYRXpYYJ55
L6iMxrrzHnpp/Uw6emeJ83m4IT2pKN/5b020I9NxdE/MT2ra3STTRwBK+rfxgDj+MzBS1Ww76u1j
9Lkwc55qLidnKT4p7de0WjBF0PQLgg9JEbB7PxZR5dy1ebEIl8/mTaA7b9IDDqp6vVke4kzU2i1B
OLaud9kyzgLD4JgFKiCYFIe71ffJRzH9nTdou4hYlcR60M34O45MXoUT5s+Q1xu+jgvW7pAqpUlI
s1HeaWMk4biZXI1oXmyhN4kQz1QudLkcfS9LgWXt5HEfs4o3uzzmQcfgaR+LrENXvfIQV4Dic+fD
82Aj5HPAO6hySsHyZpM98n/Byd9FbsXdMB/BHGeWxfnzopu7V7AIvIPm/aMpr0vLGS9eaoHdF01k
D0zLTNmwp0/M+cGeDub2BdQMDFM1tkugksf15nqfulIq2s9schE/JxfxOxr474EoIRMRT5okHpcb
kQJt0i4XtkoRn9O7U+P1zaHrrcQyOxDJc23Ms2uDFlataW1Gzs913lO91ct6OO9JkRkH6apYN1vv
6HA3PAHZMkL82ES7eF5EHS/+WvVZ1cO3ElHGQA9V0m3f8jY1/VU1DTQTzwsRVRNK9FDaZzBH6eAr
oy6Z+x4mJo2qC2S4L7J+Hd41nG3gnRD0fdtX+nbK/10Ap7iDN27auWriZwE84aMVWHNxunSovmJF
pgLf+Uo+oyxyiM4O3B13vLS+683B3ilTZfae+Vwx/fRZUlWR971Nz+y90w6yNwuyrrWEPQEhFJcD
y6/Mx7Hv2eoQAzbvefMW9Lj0DdNWX6C8Z990yRF2cT2e9aEL0TUSN3tXYyX7urbnWougH4hwOkDW
jkxo41uS7JU2N7vYyVu15ZFfIHyqXdknSFTFPk5ZX/OybmGwppkVXqeJ2dFnKKorU3MMrVWOyzg1
3byV2hQA9wugwWlfmI4hTAqW1V8+SzH4h0Iaeaocm5NFYgI1Ih2PPN08OINC+R3pytT4bmVOXDnw
d0A8ZxffOIeumadc/C8CQu6qxg5cc+E6e7vAx9RGGVLGbbbehe2FEGl7YZ8JziQsoVddD/blXfaY
HirpQ3gSFGzMgCxCI48GO/y6/x9DG5btNaEwGBdNlv3IfldQmFF4GNfYFWZ32z//o8hgql3K4iLU
baKqUNSzDX8eCp8OexcDN7CKihn2+RgSnIiYOXkkwRLDKCwSXDP0h6gYF0dqcg7PTyLt4GCCzIxj
q3ZEz4D8H6aOwElMrcMiV6hnF0EPa3CQ0XYNu0Usc6ISZjRaZn0PxkdCvdFmhv6Pfux9ATb/vkuZ
FDncUcykSgUFcWtZYl134qHrRVDrrwGpcAE2XfdsSO5LExAuMYF0YsJMcTJmNSz1gkXrQudxjpqw
+2OUtIGcS5IIajd8tyB8vrJjTK2FZship35z2kTho0KpTLMWIfj5gqArxl3KTGbq6NdPCGF8/cuu
ead/iYJy0WY6zldbBIsM/SvhmCt/TUab4ritSxY/KrcHutnIveLWgXLnuUZuySJ7YuP08DoeJAqf
6e/XSkm85TxYtPIgAexOZZ3uggQYwcsFtn/6k/Pxmng/rf+20OGExJpd1eyRHtCTBic70Nt3EKb0
F40xJY5tnotX6eMq8beylGSBdE/jkn3IsP0JmAvmI0qfEZsoQNhM7uyR6byvBpF/7mnGFPHGVGB+
6x9k7Wqf+J5pBHqRgCYO3k/Y6/wckIUg5H5A0BPmKE1s1rLzxEKoOKEjxHd84GgctFMEgATkzs97
0TcyU1MkraKPXp1kt/xUgyu4I1F2GiXCY37tVead6gxCMXdEaKA//soDDSy4FJ18ir5vrR4xdJbd
CFCp6HfU4kddOp0sVbx1YO22y/prllhQYQtkB6TsBvNvfeW+ucqQY+YY3u41M195MySSum7deeFG
ey0N9CVoNNGgAyHl3QCw0V30tjnyDVI1q8TFEhCYRxqSgeD2sl3u5CQON5JjGedX3vP2RflHMX2O
TLZqu0LJBaHb6vcgMWejUdlas1/PwBTiawgOoQyLVh4vX7ytCICWWVhKNp7Ch4IqH0ElF8RdBsw+
bA7jRWaLqSclb5/vohgvqh7s2nmiHhQIPHdie6Aocv30uzsxEPuJF2P0cKWo/ZgOqT7gb6IP876C
AUXH0FzZZ6CZlKizd/vnyUOYOvK7kmTLhnTcN/KJ3lrIj4JFUslsvKA/2/o7rPozQUq2QE3VRS8x
03d/uxNMaXtCHB0wPBC6td/dEFsvuk3cFSSyRUaejF7p/HwB/PELD4nRl2fsigTnaw2mB1JX1OG8
OzZJN63COjFgV+goGFe5n8UpZodJQZrSvgrtPZdD6R9B5h/405Oc3G0iAZRsZ70yKWnV1i3acmxW
UcCjnvZ4shqZoLXuobhEdylwSYTXC0QABByWR08uclKA0r0wNF2GlMTivu4LGx6OtD/nJjDyMGeA
HMraKRvBDJRG0j75CerwiuvKNciNi2EVS/ZWrrVZzw8HEn6ndU/uTI4zDcG34Wilp9ySgOB15nDe
eazSLO1WXQN3LzK0F485WnoHTVAJoLJUINoHZQJzEMkP7iNcDDueQzcUmZY14mB/vWyPiIoGyNEg
89C9nHtc6YncNNkdraLZE1jPEe0BaXv7P5QHPka1EGbvpqdCLdrn+H/qqc9M9nx5JukrRGToT4ug
MLINUo9vZLfooPDSNGr0XscTSOjpgEcXgLR/c0X4J95GToXjGFwQ7mszUouNJhUmSSrVhVKVQ7KZ
1J3t5aifLXk2pc9vHHt0Ygio13IiwCN6kYhwxslhuLb2769d13TpYbdT40x0cM61d1Tgq6jalA1z
GEohUP/59L7P3jyXztAQvNoo0S25bEa9V0A0hdlIIGV+BSI08ja3Abep96rVsX3Qk0MO983r+zPl
S8IXcQLEY03rtiMHu1Ctgh62ZCNYmFdYMYCglqTfjHcFcAnpwPweOltxNwU5JZ9DTv5LN9TzHuOE
djE92yw3Y1z5RHznC0LJQGpvk1D2n9jPq5Z3dksxK5YBu76hZZdvSaDQcIEw9H28PEw4042xlo2w
dcE1HXjSvDUdC1jnENctazQptPU5iq7Zz9ZwhYPchRfb+M9pp2y1DiSPVdH+17lzdaOFf7YuIZPp
LxoBW/ZEzSFhgzS/06k7nWISK6xgtn1DZ1KO5+eZ4rQPGJiCirfyPMP6+Ez8pVHfQXIQW9+0KikQ
gopU7SBqRMhIbPDfEoNYtU4clqjecNLNP03kkHXwLBblDtIo2yjdxaaQqhX2wh2BgxrWpBdowp7I
YtMUPinHrWkx6J+v3Cbr6pDlC9OR3HljVDjT+Xvgmvq/O2A3GL9VEKe+tGHn7H966Vejxxrel1TR
8gD64/EcbWhrrbF1U68I8lJ4pwTEDAE+OeJxg5HeSwVgcIrKTUSxEBDhBm81qaERk7RbN4NgCZ4L
RclmulTubtS2aphqevl3/4fVmIrMkQ+WypgQI+Uv2dWIyMU20PIa8O/JOhMJvUdpSNbkwgafze6J
+xr6lTZmJehyfm8hfIeL/lqYqjIJnUMJjMomLjnum45eWs3cG6PrURPyMBcEjUHYHAe4CN1TVRuA
0TzBbu/NsCMj53r0wHHJh+3XC1N7WcDOCMSEwZcUHfU31grmatj80TeiVaA7s3+VIboldfeKp/gH
WPrHZsRROslXnIh3jQBOYi2G2gui/Kdhir69QVOphi3ycxXkzBZNQ1BXf29pyRP7W8mPLA/cQtpd
VrRS4ivu3lOL0Sn2ZT3uZt0WQMT4gCvcCjUb5UrlppU8Q8IloHCUT12xbHyJEjC7XPK5pKimu0YD
NUQySg758wRMjZyuyI1buRdyMia7cI9iNo/oC8dfPZ5+rktHeVh/4D+fokv/YS05C76ZM8jdl3vu
7EcfuEECdlPHA0wJ1h2CKaKwcxHljY/AScJnRUHkUB19LRvEIMijzBjfGMKfzMDQggrjaNymiH6d
tvsNoKnQ5MAHasI2BPklYtcHmL8N495QDMl+Tx8oKcD4UiymJgbyf989v6vXp1lo+4Gbrjhm8SV7
mdQTf6Dr5jOwQ8e0PA1ruNMGmsKmhgIim1sRNbwoBd71wI4lt4UAA5uoWk+9OcA9umvzQfkZ8dBQ
u0aUgDvJX/hKQlgpdUpV2gBYkC1cjKV8aYQh409iuhGOS3daxMeFrXmOQNHcMyAAEZQxnNXwvSaI
Vk9Pg8EgQkB1Fah+607q2nE7w29GMzwz3MUYh6bYwfGZ1nO9XpoFw3YpQDNzkAnnJe1oJBRSPliA
OESOaRVYDQctYka2kIUdvt19On1qaVOD6JsRG2djxPjpyqBo5z6bJaYaoYIZnRKjOdN9HWrpL4qU
MtUStW9gV477qi2jx5ynchDEJ2A3ddLluBaQKB0bj56xmBZR1QoxbvaoidVHIc+dV1AWmV2awQ0H
bDu6XCfdNf+3EMhXIzVGCwb+P21hhl1cT1ucNZjtmCNLPKG7Q4WlEMB1CbPn+63xg1EAGf6Y75rY
h7hddu4pBlQJDdYwbWeNKilHNLHk1zmZk4BjzzrGuEh9HeONftgbJIJZsxZ4a7ezAq6jq3djb6Hu
XeC3pt6oaXBqZDyofplX7GYnF3fJGI3OeMh9o2BEwTivBGN6/qipGSniPkylPPvHFAt/gTESfMHZ
kRbBMKiZcD3GhRc9yNyJYwLnK0+VIFfp6jVekCl1eWG6DGP2fsLUyG/fMcxHFHXDMWp9dqtLsLRj
eTeGNjaRUGaCuVfN3NfO6VzDD+Dfh4xPutnPjIFMB//UgRAGZBUL+03lvc+Y2HEntziOB6cKFyT9
JX01YKIMiRH9Z7RMG6NBlzfBh/2x3B0NILZwztzZHX4LLDIp3AlqLsSHbBfUqKqRI1tOYCyzGDB/
oZuReZP6uPVyt2svS1cj78pTlUot+AYETWdLqQPIxwPKG8ANPpXWfc57lNqkW1zxq7nN5pDWI+Vd
U6HDjSNh6dtd4Is9hS0iVz47jPNd6kQgeWcM+IYeG9fypUZtTZrWU3jrY7XnAOe/JBWp74UIARk0
+fdEdw6WHrm1EEsvDOj/YtznCJKz+qI3yfhhwMM8jJpSIvelwp/hnV3oL+P0vzaxIuiWFrrjTJED
TBLT/A9Spywek+7g/1QhnCmzJn0i+BOCDh60kbeN2ZTSYl/Ik2VaQu4cG+8lOAfmtHjz2Q95A42G
WL73QVELZlTEqi5nKWb6qckR8kOLfX4giGxTA1wWBKVIj72VcmO7jeGt+AGUpbmoc8hTxxRfeLSc
k1t04jq/GYdWghmwDURDf8nre+6XXMPfGzGUlmj03cCtppExJnKjL0g5Rrm5HAuk0WnDPQMM4Dzi
jpkPrPtMlrgO28aFTEt/AH7S6LS1wW9aSzUqpSZxb485dSGMYrdnebtbfqWhIosH7JTuuY0aUtJi
nDTD6uo3RNiJtj9twPTtsDF0VSX8yBnNgH2tiofbAsv+ptOQ8D5eobkPnnD4tTCTe/Q7c7nieRJh
GGV0SeZLBVvjeVi0BzDY+KySj/I34eqUdNhHKTVtfxrUDSgSBi/aYMtJ3DvqXSTOJfowPHH7J1Tv
7UAc7xk0vZdvShqBtV65akCcUbziEeBQbXI0F29j8dzWcA1yg5PP1uIn1Hdzeva66BtEFUKo/YIo
H6tYXgw3U0Qhk5Jhevp9qghgk3CEeQDcDLQBnUjDVIv38ToHtjCJwKR1O8FVZCKfma1A8Vk0y7yk
snVgEsgRInULlyh5DDQh2OaleoD1WDM9tsvSeWJSshm7x3MUmUb14C/ynilvBw0H1F7X2uUukE/P
MUR3TMoUe7ywaCJpaY3FlQHlRkzuh+k/f2I8CTxsgcR2mMeJkIowXhdzvSGORMFNg7RVNcui07DO
fM35teY5XDUGQ4s5Ul/vrz+8N7yV2QTT1Zckc8rX1dw/mZL8gSEGbvAaM2Cm4XQNs4BUON+c4+Bi
Abpa9P4SQCzsJl/f5eeJXxMuZZtwwYHdBEfBWrkT7R6/tuiYf/yRrACd47NfmUfDMrGf3lZellsw
5Q5UvJS8IYXKUev21ek91gr1O9Pzcl7nHZA5auHbgStn/27Z6CBq8NEi6t4hdPbJkG7p7WykSl3V
EUWKzXY3+aBiVA25k6/sSqbPJ4me6sqIqoySnksi9nkyS3G2frJCteGA8TvIVflgGmfPm4FzM5z2
wrlhseJ63LmT+cNJ7TAyLxEU7nD7mYg2MrYDHQRluIMkk0pG0b/imG4ufEcIInV+NDoAhlVNuLMs
9vaPD3gycqd2CVdAaauTU68Oa9DTZzHzvD/KVfEQ1dIvvWYCrHvS1Gwts3OYfOiaaV9FSbIj0ml0
LqVvFYrPF+pachcGl9sLn2gDh1PbrHX/zY6e1kZJ75eFePRL5rIskZubm/ydENdzmfipDajNKohr
8joH/5HjhiEM+Em9OV+prESOX8ChcSt2lCt9I2v38DQ8DAE9GEHldVnTfX6tu2LqP68XS2y2bFek
kWamprFWMXBvtoHVRAalFmBjHnadtEgLQ1bjnpgLuNihGC7Yyjn9lmxWoWaJySYzfIcMDqyOkk4z
w3Di+VhCRyO7wMfRQi9Y5fvulBPj7Mq3Tkrdr9xskqthUx8EuEdV+TuyOmLCYxhY4zrzjXSmiz8i
ED9fyLeQya1FyyRRJO98zskUUW5Mzx3ewYggmwGillarOaX4lEbQIU9epKNWRWz5dKgkhDfbnuzP
KGpyRc8ZrJ0QOjwO7hXbgIUmOJNxNrJsm+mPmqDejFJsTA23gOtQ5XUjbBAmoRLzWvpsXIfyR0Q3
Vgjsq0zzhXc1g951KU/SukyOyILH9+C37HWZwhHWiAUDQ71UrEYtXMS/wob/shnJTVaKhubDNr0I
9EJ4jJ8KNM9PJ6z8n7M3J0LjN1xs04rn96np6bVjcXZrs3fVhi6pOvrCfUL2lIguI0TCDCA1rPwk
mujAcyby5r6peqUeazVHKb16D0wz5eCjp3HE46AnsnSglWYdDTIcdXYzRltteAsbdV48Zs639S8r
zw2RRubzlLWkZMg+Ag3mA6oiXjj8+LaIgfM2dC1gIFhmO5ThqVoe8xlDRLmRNDitDArqAO5+SOhm
6j69CUO40QQvKUnRmbG/p34hIbqGZuarCNPX8GLninzGi4h9+D1iu+cunoWwvtSO/cK4mDJ6del6
U98JHEAza6g/mbNtVMTUKDzEhxBt78RjKjqVfPriTf+9zJPT5Fs1ntiFpNriACXEsx/zyqBRO32i
72kfp8PB2g1JNI1aNem1LGIpRPQp27+P5VzaDFYgD6P/YSmmQBCRk8nBl3cKLiTO3ZkC4pwFIgKH
V5NuIkOka0eiRU5qWmm/2DpeZQ+Oe/kvJA3lGIRQ5K9YlaVCsdKtPTc0+leLpB9IehGsP3d6/q3H
d+bKhhnZxIpz1S+J9xjaVZjaFlE40eh1Ozs2MP3ItA3UkqY1E5LuzgRRVymCWKEnr+T8TYxbU7CN
CZMzMtBWLH9LD4BDWSUliZXvLUCPLBATO0Gy4IXZvbHbpE7o/LF15VoGUajVU1owPS5Klt+mK+vW
BCqADSPv7IwWjw0OdhRQdr/ICmM8KNHQWIhuZU0eAgHRZCsf/P2N1FoFIC3/TnAY5y9UgAbibVxp
Wqh11bNXLwnGOl9k7R7ow28tt+euEtMoW0aqzZ901WlXC5F1k5J+ZSUWOG/bi2JzzN+y8q7g3fhQ
RNJaLpVGQlRlecJYags6sW9w8FLBb0uDZWrlHCqdldswCw0QjQOoosfJs2rfRWnjxfVpSijAhcnq
ilVBdPeHmoI8qGZkrTi6MvHHCf2WERWM1RFchXgyA6QjtF96gj8Elue6pwCLrEqmewwelZOjSoa0
++jG07l0E2joAt8c27NIJgTDcnGMbNR9gyM2rdtlLXDIu5uqf4o1bUOAFnD4pY7h8gzc1LxAzs9h
+aRNmlJwTpzK+sqLmW26yAaJBBJHZdhNfEx0UpkUZcTpbcv8sNAvOphXxA84msfIhQsvhILbnDYA
HJD2sYgh2kj0Cy9T6VXr6mcBITbqXqqBgjgeTcjbMUC+fDRcFQtTrCgGOaAZskomUfnwD6WgELuQ
lpxRdDi3KLAgM4KAbG7D+Yl9503QApJP4CiA08+LpguoVdAC6SeEO5mwin68ZngMGk+SgwqQG66B
xSp5cxQqfSvH3PeIWlMO+pb8p15J4SNxhXwcNmDIgqBFVV/dE7o/dTFBlmT1iKRUPfLSE+G9DThA
HCB6qKbzhuGnrUjW6Uzw6CFhSDBdxpqb2OK198SJnmp+Eyu0D3yqg8Twhzik2FAJNTu2K+mXZcMA
hocbHrUW9iAGEqO5n7kJWZw72A7/d+4Eh22h2puuGCoo+aOsRHVx2Ihbac69CEc5sHWnwboEWhcb
GUDsvyGPkVASXWS99U2VjLRHA61RZQyDDL07rUNRJA8ui9KmRMFNeGnxcY4vXDDppVQy5DsNfHl2
ZoqxKcmo6mTiuuLJRqx6AEXS0YqMtkWsR1n9WuL9g87zW9Q14XjrNRANUGEnrB75bEtPRKAEWXn3
6xWtuLBsARhpyCPXeJpdF5+nV6q4RCPfKygcbjys0mST7i/TDx2JkmdKFEU9HdKqFIEu7T+y+fuh
zowbrWSmwJ5rjcCNYxAEx9SBon3seal+exiWTHhJRvdCt21ng72jtSRFOArM8u8R+NakpQjP2TGy
AYW2nKCU1zivkH706RX/v0OEICsxi1qlju1PTBbxJkTdrOY7qpqFEjv+PidXcMBDoSKicqdnOuCv
4G8pwi8HRBUaWscHjDfT4IUfdhG0/D+HKH09AxdTmyB3/Nd7kWVhGi8YDivi6L6xEGFdynzyBjFp
gFhteu+6rgQpDQovQ3X8NKfhjZI15+KnGuiLR90Z1bfzTGDCrfirOW0KeO9Ch0gKueCNQS8eV111
03CSG60dTGR/trVJlNvkUgGHhqBWtaSuzjKEWNVFFQCFfu74lED8eGtBtbmAPG4lwqhg3qpXIM5o
NaMUDmh0eK9v5xlGoogAc6BWuPqDFn+qws1eZtqcBkO6sLuE24/Y1m4IpJWu9C2BGMiBwjaQwIw9
ig6pFAZRnoXLKidGXrRJoI523d4EevaY7+JyZ0OLesq3U0xWwuajihm8zvbORr9OMb5j2aUd5Hku
a6Z3/p3JAPoE9h2TY8pYWo2eLBVGIMCa5pHU3mvX7a/9ZIYGCOX4wHOhMpmGPWixb3EUuocHPKqy
ejvOAo4Li2fWO+5iPJUjF6thZGaNSCI9qR58Brp9GlP0fZHBomzxoPeP4621wJQD/Wos6FPfByqt
57VjC5FvrslajeIJWiWfEQUmZ6Z7pfj8Qj2+vg+slEbycmmT3PDVH7JmbQYhmpf7t4RsfyOLX4Ph
p0dOgx9Sm5B+OrrmLwrRcW60gow35Tk7kEIe2NSNv9tJfuEtIm+yYldLUG6vWmmmMFxZQg/WgaJ/
2UYH9B9cKRQUbZ2XvWfxcf2YOT6RjiAkAn2TAXvvs6BTUlGevQjl9Nu5qT3c7hRwkzDSO5m2h1QC
x+eWDchkLUmbl8mmGqOipHRaVKOWLX4aEAkmSF6KyB9LMAGG9fPtdJ82TtKJInA4YRO2ZJBubceN
M737Suvj5bVyM7oM5Pfw/dzwoX7sZqtZzPDSRY/NEmQt+0kBAZH/SkMyXTixSYnTnVkxnQflUVc+
0u9zor/l8cXQ+cUp3x1AtiHGhIALPRnxj31tSU6glPA/WbAEN8RpyO0+rRhjtQVx/hdMofYeh2ai
BY8TxcDppDGCLDyk+09fKpmRJX/X5HFQbuFzekJfzwZO7C8NzHh1CRo8ou5R+5T/h1pRd+qiRemF
zfnlR1KbrS+DWOSjFA0O8HODRZgIsflF7tPEG/1dQx3ETLZ6ausKt/VIS/ZMDdvWO97B1ZlPoDyL
k1wS+iFH9kvV3WNHz4TOw8PzH9SDhChLPeotL7UIH+BBUBAbbfiDd1fgnYeW0/rQnb9jHPcXU4+F
TTm6D7OKnMZUNqG2mtOUlE0JrCMvIMaDP58kFBFYegZVJ4UFfanbRQISqOUsybgKOsp6XvRYzZ1L
+RrAInx1XewxkJTKDBU9EBJlUT5y9Sh3okjhOCJ11HZDA8aAeCvSCM2ZPUA+xYwo56azUJQI8gAm
b6bdazAKGUTNXThwk0SE/IHOkPZqyacb7hnV/GWSYm2hEQTDMZquZJbxXh9j+THd3EbXGGwROTgH
NxBLeeoOZo1RRBGB/PLwUOnJ3Mne4dy3/fqaKUxiqvT73nVJ3NhBTBEKenWRksjqWAmfCR3w0iiL
/xw6Se2nY1VXFUAHjQpW0CEOw72PqAoUD/5KAk1glvB4WDjE3H+g76KKFtrqFuKJce8LixYtUujg
0uWjEbUANtGLCmlUTx52ao4NfPDxdIgGsiZKjKxJUHCziReNvG7SEZhgVPen2/W9xVvaUr4FdAzf
GPRX20C/JmqXI/fZBBLvkntimvCwKs7XeMbpNX4H+07h4dFX8fmQEw77W/ZEmIjqdKCrBtzoW8gP
7z5PXq3teaSwxkkaZtdm7hHb+X98KxJ1iJMI9eREozlBbT6t+hnYrhoWrmQdx75roDKVNlqBJ+HE
jJBf8B0TxwdOxFswaFsb7OPPblcRjDHRLU78rXWhOFgDXPsoM98hHxdnhdDx/AfiCnDH2cJazSeE
G0xvOvKlCM09hU4Q4calbC+I12JUaULu/Z8jiB+r0Levam4/GMknP84WbJOZ12i/mAmaWDSKJ+hB
X+3/PDcOxyt4mvQVR15gL5HiP/GFRoJ57JtK1NKPY+P+5kKfszCt+4LbZeK9UDPnPxCyE/3AIPlb
/1F2vZnRD4dmTO1PaGPZX4dmu+dr5H+3+WaJ67akPWAD5Xp/A4pi5QkQ5XBuqQch99ai/seUIokX
/OLkbfxtb+0sd0xJCGREwGenN8QwAYvXceMEnGEy0KEceKHm6gFXGY4jc8CL6qYAakSTjqbbj/PO
ng5Lrv9Wroi3pmnCqdHaJ6iHa/GF3w1wnMAcqADYW6LtCxOrOCaOWU+d2ZTQvOO6PUtNviOYfBL1
+atB1uHAZCKDgHcdK4JgNKqgsnVjJEF2UfuyJdDfqhL43OWmblG3HQStBEiDm3NQjgzEMJ1bzR62
av0CRXDrsxFuRLr76V9ocym7nCRHiTVkaxaUp+LAUkH581q/FfluzfsotPgRuuiWWbyWx4+IZSY2
X9IBM/9EjobYneifS/Tudvfc8DeVJdyd56lFzforB7Tb9tyVENjtJXEGPMuzTZ5j7jO97kP1j7v3
KrKB3ewZtAoj232j98QW1NTdHskrFLISRIvP6LjwWzxl5qfK2fKAQOywPRGo2RCAjwq8eYjY4Cbs
Vshed6qGCD16Wru8ZQxhRr/zrfSlbfT/bxw8gKEAEZv2Z77UFs5e6rQzX7u243gj1vMTN7q9VR37
lr58endhA0cym7eZG9EqkTGW2K9n8orPhNIJvA+e6XhaSuhs5dzorAZSk1ulED9tVBxTlkKKmv2g
t1QnebGk4eePtQmcfEX9MKSiAZyBiBopiOvqxRzbqCDH1mnfcZTwEX9lXtE+l4c3myde52sY5nGT
9TSSVNTMLeS/aFaMTixsXS4+Qra3zwIc9fZYGV0uaHtN5MaE9/k6aUppkOU9+PtZpt2N7Nq2qd3Y
Lqxl1vaF3TjsANYgEOrouIyUJhcPY0w9sKrzyRLKGlACZvfOD6gt1rxWMP49LUGrOZNsML0hNZK3
4uXvX94ieSQBMsg3u7Q/OOUUOAqh2tu4uX1BloYQaFEe0JVZAzAw52fX+tp12rD+3a1ZkYX21LuH
ykZ3NtpnpNqEDLtJbuN1u1nPgZarkmxhJv310fXq3rBmZx7miIU0/EJ8S+B1lNklB1W6VtYgHXh9
OM4ELb4+0RLHWx0DSxkKxEkQOcAxLe+8VjhAYaf2OO4Hsg66xqBFzp5h2t5/cPyCvFVf3q7zAEu+
ZtH4WfGqFg1m4gueEOou6uk/dZE4kqzF2b9UZVY3QtBTlJBNzUmP7vVg0itdRfRqdxUhTVAVpqEJ
iJ2dg8f2+EzuNGcjpM+zt2BQX9agnJct/nD5kz6Tc1xPXvWGgF9MmCp7KWgEFyn+6/JPMkZVDlKf
C/GZfSPEFY/7iIF5ufxaD5mzU0mdCJmcrUB/UNbQiENZScgbftjaXm9kpibqYrmccY8lfQedfsAm
VJWtHmRh4+OehhusGc1WHqqJSWVGuHm91Dn4nQLWdj7QTKVR+L554vWzgZ7V+GWjWiZr1UUGw5Yn
mIfJw23wIPnZz+iKLHG/9n1WVtPVH4vaIPugEVyA70cHJa4Utv3Sx/JgenfwO05jQqu/kpzVk8i1
PKyJshwcJxuM4UaLAUgwQh7AbLIWgB+xK+Hv1tBqg48g7bHvvd1mikbKIeZGCwqXHEH0ImYrBG+w
kRpWWwc7jfnlZtJ6F0QhiErWYtsCSIzTkXH+HAGMYMxgde2AKSZO1d/jZTPsXuJjVGI0K4GqxeIE
xFTvEHGewpzFhequa1btH/UHQWZKFhjcPGQa8/wxhsL6+Jk2x8oVIqiwr3Iw7PrxGTteeOzldXDQ
HLlcjm0wPSvcFZvthqLRKbagTs0gIFE88U3pMbNtSrxvqpR7BKCNYK3rJLkH7nMBX4f9sg1AOsHZ
dnYZc33h/j4dozuQZfWAX7hjOsbIERyV0kWPgEZg3pYCBitcJes1uepB2JPO1mYcNbRFDiyke6vc
5WuOjkOrF9fW46+3ytzbS8HruMbFRwYPkiBVFRiOjp1zdqvTtsPIHUqTb2j3DYjxK/UY2XUc/1ys
i3x6ZfMJhXiJLytIoFUrOCYnuesi3b5iQBse1FTfSdPPUWqYNJMqFnwJGrVdN0QmpcgdQ2sQALKR
82HxL3QhurLoeMQTNfyqi3R26oC6IaOHEdbrPaOVk2H+iXvrG2J3lMiyUZpDskooEb4EeowQ+R8+
+W4w4Dzhx0Ypk8nqXWMjrHjha77kIOiJI12C2O8xhoCj/QD5te1Et1s+2gb/mkNt6obBLN2Qv1W1
6gZFgS/Cs9tp7rZ6ICV/ofGBndcog4J33kHWPcppQO0QNZBVUG7h4LSBGOxGa4LzvrYwOIcj0wmm
7RjVppaRHe1LdYRUR7ou1kEkHkLzhXroHuIa0Y7qyUeilWWdAYzF4x5fe2T2zO+RX2wjO1qJfrTy
H7OtnI9QK0E6QTOUrUUr9SeYw5wZvfeVhLn82SW1dDDdXSzgxe45BhRfG2i/cJrEqnusYkCMucCD
nVWUPyTKNJgOBy9FEmiwtbULH1RPqI32l6HUhb2FjD6tH9Y3UreEdbOCr7LGFIqdgshySU+wtUhq
rZnUjzQtu5GNiLlmoRSv2b0ABjn2IAELqagc1NIu4eX+1dzFgYHXFtXburWseHZn0lSfiRWwJilS
0mkjx2nCK6om/cc89xsDuZKK/YMViwK7EhavpsOMhvz/DxzHJ9a6jcRJtRPzy/ekC4Wot7XX26T1
cgD+QRhXC75kmK1LrV6eZaZwR/ik9TSugJfApkubnA7HW7BiCWtDdK0Iylga1zPs1b022QNTpp1a
ZlGkH1lcFaZIVVkIZPZkairjWkl8MadNNRRpbTjGiMDHAisT3ZUTpYH2p2EkvtNibvH8nYwVTLsp
WL2meIHvEKCoFwrY1PdmL4cjNKFgdhZQxJKyhTG9IrqKGdbkSWkXChIStzorcwohzDJlzB8e51BY
QxKiT6HSB0MH8bSzak7fm32585Xt1aliG+bGlgeW50ShEb48hWuWZOO9UJVnVOmPt8taQKI+pz3Q
p3UbQSi/Pk0vfyKew6EBfSMfoywIGQSM217URAh1TB7mZtrIs9awYM4PExn5MCdrX1v5zrsCOUJD
HjvyM4ovfEAMQcJ/YY2wWE/NEMH9Mah8p1fwiJjrChXygi5ju294FK1dMv0Ed7RA4MLM9y0gX3dk
whO45Xru2mnjoEwV8KyCQU6RMH6vsigQVWikz0rQalh9LLa3s+zcSZdJ3kNc4POZHpftVb2Tihl9
z2+GIgECg5sS8IZ0o3HOZ4U3va9eG0cI6JB9uEwc3hq/70OZJX8S5kFZ3SGe/gCaTQKqk+XuAhP7
JUIWEt+SySr50UAjzvB79M8v2M81NM8yUjfTcT5e6JV5TZ9+PueGeiWyZO/b+TnH1L/FxWLcROOQ
gRWZzdjOdjWp4PSW7Q2ZHrI8iOM11tr5gWfeYXEsAUloADRWT1hjrakK23koEQMQhYrxkP+qzsxj
eBn3UIzBLSpzC9EO2+VTJ13XPd+R6w6uydGoYu4EZ/IfXcW5L9vG37HOpABG1huJEnzkx8PvGxfW
9PqJ+SakhqxNxjElgBm2LsDIvCDUqYNLwSWJn48kBdHfUPcMp3LqtaU3eyZ7qhWc3664C/m/bkTZ
xFGC9l1so9AGT9avvB8YHEqX7O/YOSWE6GWsQY0WB/lVZIU9Ngj6uWTmGQ+R71HPGXnM6lyScJ5w
HKvydK3DXtMRjC6qc5dbfjPbSoMDvfbZBL6whH8yIaPqD7n+vh3vsXXFz/gw0Z8BmdKzX/soGDsT
gte2sb0TFHSB+TtRkQb4CsFi/0pqaZkDZy5FvJVw56FjTBifU0ki2jY2Nphkwlt1AINl9PNSJxAt
OnCTIxzEaM6cEx+nN8P/e8ZFTUeegOiCt1YsxA8cUxKR+BKMoIFxMM93phv8P3uoxyEBNwVlrEYv
wO8bbceT50RSUkmADX3KbByWhv9V3p5asM//1wAsy0utVkX/+9nzAM0UK9KGfqd4SuEcZA50EJY5
7pFarh8ZSsnSnAx5YSLnxgqW6EQFh+djJ7N3Td3lhP1Mq5sXCC6CYcYBVw2nUQXE2i9No4YnXYZF
gXSTq2uVjUvD1NXBNhSvsFb13nNhXprIpu/IV7pPuwumPp8jvh2G8ETLuxNzYEXOp/zQwN4/nAvx
oUQgULZXrDd6bg79pqp6lRS++G6/uyFY4boRdFsNQahK8Jq0YtN/k0tWor/UY/ZXICNBhbKlIZF5
dlfT12aPcuMTQ1NxDboo6BPVd/L2LLKU60bbRpgoHaXSc2ZwgzMTmiXtyBNB/C92JabCwh9JwUMh
zYzJZpdi2YK76jkKeGnw8Sfb4++PzNipDtt4z+KDQTNS/S9Q9IWnYhou8sK3MM42BL5IP8Oby1or
JIC/bso8xU2mBhdf28noK/TPk7nL97QWlg5DP5euUfwEKRchcxSBUqzv1TsPOFFs4lL9v7oBM2yi
W08rW60gdH2uosl4J6yJSaSaf5pXUsq+862QWg066QewEeqoVl7v9M8RM1wKVzLNfKkgQz9VZjru
NMAiKOc2LWewY50oppkf99U75/U+wzMAZPRh7+SJdryYsA+SF3sZqzh4amSPO7VTENgdUct9o9II
b249ECpNlA39gn4yID6C915BeMbUgmh0TI1ZWrW1xOJS87FCshtan8kKYY8ZkJJRF+haARHYfpE0
D0wppBrtT6qdxe6OI0slHkTG8yw77dpfhd+zkfGBcNNx/EZ0Z3Xqs/AxMLStCTmQglZiTfqj11yy
wjgbJ76W6HHalYQScpg/Wf9egBfpyR4ezB1vZp4IuL7pbsoFfovtw99naPcJGkIdsaZTWI0r4QYT
dHKN21zar7xleIDH6SEJbVkcjRYoJl3YN0THOv/H6E5Xd4XRn0wwwAQSFdPuZmmIkfep0XrIeH1F
uWMOtf3KadAYlBeqNOT9RsFmcx+6DKpfV4hZrYEmKlsQTG1sEnNcIVUJ8UtpekiTJGyk1i+EnFy+
x/8MmLsIXSgCjhRHwIbJkErpEqPtBts2jx469Gsh0Tl6FAiSfV1wtkKCX//WLoi9COQ2nNIak4AA
KE/K+KVUdc42STdBrYXukotO5C4g+EIoj44EgD4ESV7y1fLTMTz1FzAntykXDN+xLtdpFq5gZcnE
WX6BkQ0Eqg9UdKxh2Q1ybO3QRCe5IOs+XYxFjVMlrFaMxtGI6Lgz+Xg+iZ1h2SwFmYoEQyt1TKvS
wp69ZZkmpaUcTKegDnNMSOY2YqdgUJXBmcaUfw1LDnxFN9z4qlN05mM2tP+vRAFgSUSvw+q9/q4l
Taz0OVm5+wLnYjuOKADlqxndEQhrZdnOJFMAmVnfBq4/AjFUqNbD6xE9S2F66DD6oF8SB12cAyUh
/cq9Zlelj+7io+Kr1h87oPGF1T89b4yckGTHWfTi2gYWnEdXXUemsrDqcKFOyoT6JzZxvE/q1X8M
xQAosx6iC2rtB+IPKuJyFWsuC1885rqPHMeii73hLTdSzw34l8x1iR/brgJVJxOI8uYkGUGrJTQ5
qNbYXsoku4xSEB0Ep4DHrjVsEeAWTiMyoc+uNKcHFX6iwww9Q84m25uRbcY1kyAVTucxjjz8ZNxg
JzE4t6Qf+sI7MVkwObTIO3IZVmMICe/xiJO5BaWNtJrxeZ5k2h77dgUzxad1qEWrh6XTKv+Sa5aV
5yoGaoIt7ZqnqlM+Hm2OKXWBMr2Q8b2KD0FkcLpeMviMr7+gYGau5becwR09V1QK8CA5sptSiqCt
X4fJkLBbS3uK3Qqi1Emw9PIgWbJXtSXLypS6G4W6eCqLhkhtrr9ErbyfKs3Ra9WPPWx5Jo08V7sv
bW/jCC8JRVdcdfwI3VowMMGirpdYJWI8/gII0vxfNcz6sFRbdvA7wDkwRIA7uwmlKjfcTFW1XUvr
WWhpe9DUhvnLrTBPdGry5lYQjknxE0THQRQYuSj8Vh673WtMhGdptQbJZRvRw0H5oOCn5g3x/TO4
oMKCVMtb+fgMpip/c0ekHFzhvnac1R2ltf9K5p8NusrEp0iI5/shh/FA+xJdTZmt5pqcnnb1ZMJJ
cIasWJzwgDI3wlVQ3mJVkWVPJeJQunsVDmvyUNd+kXDV7YJZOu64vnzN1ZJNg/nPi3Q5Gy17+8zx
+6mXTcvxMVEt7Lqd56LT9DMgKqqUpgtMeFJ8iwq44w0Zd8JL2/wUotxkMNTuJhkUEiUc3kLKXEQU
VgN4tpB9u1sr35XBHVEsDewfMpOf9UGIcBrTRf+2FfsvU3r3Xl7xa0lhW/zABs8KycCNzRm7pvC9
aaUibCsWFSsXnrMBpibMddMK72zf91kg7bV9RgiZYi720/tF1JiLTz0BlkDZsxWr3EH2Mn1Codw5
LE6nE7WAsNhK03R2ZEvVCVD4nvXTtWqiqGcbWaB4dxXKUxn2T7I4SJ95ThCsG4mE1wMYxNH/zWKA
nKCZs5d6XqinPchhW5cDAFSlayrWjLl+geVsbVESYHuMj19qLNYo9YNeRnTW5Jy2z8G7VhKHQ3w/
UvAmDM+KxkTNh8m5SxNTQlmiiWnzzHHyLZhWmoBdUFfBAZKrqjMCkMnnjoh66xIfKogxUgSlMeKg
S/mMhXluuwIiv+hxJaad7sHXz0wX4Pft+kLCyL+h2VPp3XaclvvwWLydpqSvLso3bjY6ilbx7Rg/
PMyR7liNdTXLyRJxrWkXvM+BhjEyNDhtCCzWURQV4n8ZLZfb28legZqPjQ3Zjk4UAvWodyQ6CHdB
TIJ6a2mlJkJTSTsUESKKBtmBpZzndbOKJxvULFc4aM+B+wRvYrdxLVBr6YoiEEqAeiwgZR5Mthg6
NxddViYl1caOVuHHges2rieSnymE7f+orxlew6Rs62weH3YcgJMRNHe6MWgXrEgBxTAfEAiOdr25
UifybnJWMg1UfA0sTevlAwIoq+xQzbeDl/TH21QmH+3bM/P+9e6Pkw3mckfB9F7piYjORdlQYDnL
Yk33pJCRbfwjIJYHaosSaIWNEoKJN6fY3tsH6keao1rdXObCKrbZOmKXNPc3qT5SATSGSbgyfwzf
QycBVg7qMhYzh5o5wTX5oPxGneMqk7hZgHohXG5KSIf5CdJQCPBmkw3hBp31s7ThaJ7rMT8PP2D3
S6Z7ya8aQzwPWCuqjko4+DAmqc1asLcSwChwSt6OmJgMrkk3Gz1qjMRDFld/ZjlcCtsBdfoJ62t8
T0CkKr8jVl2c19AIFE0fpjcgfEYghYxpQrzY0+Z/suEJzVLf4hbuaGRdePkCg/50qRiF5h0Oih3x
SY0ohQDWLLn17Aa2bpISZh8vNCMyK1B+nvTufkOaO9k2pYR15/yPbL9wV1ORtK+O/0CzraeN0RCg
1ZcQOzAz482PJIWkqTIBWEoQK+HIOZUhbWwGkAOt3b2YcRxuG0p+cghK9WJNjW2eujD+MW5quXmb
QBBwTV9MyQRNtU+kxeGx7Fi1Mo5FYC6sWIs4ppiCGbY3hhwAfgui008dCqnwKE8Sko6f/wXIPJVP
ljGTAX/MjoO6p3Ip17JmydRHVOBNGge3FFfbzEo3Di2Ylm21pV2ySvAQM55KmkubXXCEixcrBcya
OgMHMdl/971mR3QB+DEPK5B/yrXALrjeWfPs2WDH4MLYVdqHZxaaejFpnPfwH5M4tSlvCBx4Lhox
oXsXu/ylwlZXEbrnHIRbEq8GPE2+s7yfYbusJnKYinTyQ4fvL7+JHe1LDnuQjo6eXJ77s1CU6ST8
i2aH9mHjFVhIGwKZ+IAr4E3+6qEoLIR6HTo9qGim0Jbbngqeup/rmR1C9k1UKcT60jws8I3FGxq4
lloBUXj/ghisieEl6O3WRQNYRMUjizNvruVKRkJZkq5NxhFLFVDYuL4Fhh2D4ayuFPWG7TLA7m9b
J0XNh14DH56i/tVfl10pdZRZksjAOWvlqe/3d2P4pNkF1IsBrHaXovIi2NeVQAMMoRpB2T+GGPDm
iJIx+b2Epa1mVoobxByTVClMOpDnamidVwShEfhih2H90yU4yH75HjG4b2F/epJyIKsHhoBv+uLp
vxj50oBLbGQykRzuBDGQqkQzX/yPubv8JVoo2Ay+jmtSaxAXjJoSBSTkBIrViTwd6f/L8dsrDK/L
Q7BJ3ab2K9XDCy9Hbalrkp1MctIxbnFTFvZLcSTfOFy2Lgk0htPd9VQkpDPV2wXF5tNJdP8qrzEO
yZachiS0SXSnyKlujuzMQvPrLLm9xDB00qwqJkXynE42Ij0wvrP6W22HRpsyUJl9kKAQ7UsmBq9j
reTWiAUvVBLU+EsVDyXbMnuDRCcPbcLbAR2iFT6H7BRYC1e/YAHjGelTwEYtLgr+QvRvgTkYZgYz
ZWcb3QT05Q292Hxo/GmsD3xiDKeEhjPOpnI128bOJsXT377muUbQ1IKsX/8+iQzLEuOBgGQvY96a
+smfjxSrKC7SFZySZBSko+DXQjBiVUFSIPSsoxZUJzEDsYnIjZ3TenUQv9k5V7NeKLfF5tep3Voo
beJT79Cv37GVZMeSjfdKRi/7WkdZti+AvY5yt+BUdsRNmblguAxksXjOmrCv1mH7ydZ2OlabMA41
Dcc8V6V/WhCuJZ2i5QJO4lFhBsbW0X10W+QzRTRej+3mYc5vP09O4XgVNZlMbn8J8Gv8bvittw+/
Dk21qyYr66RtoRJBjUdPUSMqoQKHOvz9ZozkGNSKgNxh3UQKcDWp3ek6innDsEM3rwrGb4OpMNPa
idcJaO45TMhHKVePqWyNqG6QIgXjIWyR1Wxylla0qGGugGDcdiWTxoM0zjLZDjeniHXsN2tAIu19
G/uPbU+qeYK+EcwGO0yOj1L6dNjk63BROY8jd/95kWOqvRsK+Gj7SFgcq4LkxaVES3h63JAhGfUP
s5tou96bj5ZraDXVlKYbX39myXSi75c5cBJ0TLxyJqJZ9l7Gq8asLq/Xnh0/9E3WN0rjV29nzQNC
s5E+ki8+EyAbUfclFsdUwqwRJHX9jPEdyXcwZFF3gRjNwGHQ709WEiFkttF8M67ljWcT78UgqYNH
+uq7i93txUcy3GLsWzYGwMMDnVVkcOWQNG4I5qtN4GhUPpMWkN92WW3rMkSJIapKVm/l61V+385G
d7kicLgW8UkuDCXEGNGK/dOCXoP3Nj/Us+rBd9aKMaqZ+Q3C13wjy0mQIquTXfk3GR4aM1UbqMUh
WV4IYqelhuHkxbQBccpEp5vsMmTdgcwYXtg9rZaIQdtQjsINq5VOeIkqHOJXaZtmdImQ3nMpqHI/
B7a2fUMhSHQb0hg+2ayv0AfZFc4z3Hh0HHhobzrXF2g293tHvmoNm+pplzkSYiHAdUhWUKnqDR9i
ZpU3osltDI+H9YMes5CIf9a8mejNg04FVNJANM4uCNAdQett5O9252BLnlIKjP1UjkY42QS9NOJY
cKOdC6Cz+cDx9epJvNZR3402mQSiiMn+mBlr/JoI0jfl3SQ0e9Zjou7aOzKI77wffAwAdZjVMb2A
LOD3SlTGrb3VXSGdrUbLdB6upI8lNBrtvLwyH0VI+gbDLuDI9oT6zlnpYZ04Q7pJPfuQOy/89MIj
i/fkXqyEKK9/Ls2k4GQCkUISgzubXDvbLvTe5bGOPEt4qS+3g2NuagxGtTAyKvWxNTO3EUw/uwOV
uVYrlVdvs69ww6zk68LE9gnlQTe1c3EdOtAvzsPtkq9GWT5P/ahgBNqT+TO8XlyPtkgdBhan1tj5
Rl25VLx4/tQtk9UpDzPhm+HnCJTngrSl1+/h1LGIQhJUduV+8gCWEiKPAGYkOjpdOthMt5Kag088
lsIl3GeUyz4QqsAGnQzFQJ75p+4bVysVspD9dAYWisuLoB1D7lDPGn5Yzao3PjIV2YMsBn5qcpua
qm5OqOCSNdkt/mj/OyWCIK4tizkW+jrbGczLHnfRfLV3L4WXOqGPz4phSj8UlJo5Uqq5wTx5duzV
AerU/ccTjmjucHDddiaXNpK+rmJph0q+PwdFuogS2Yti+4lXh5DRIz3Y3z8LbuDKhd4koT5hzHMC
jHPtrJCQ5tNozy3envO0a9uQE+LhyKX6ce9wPjThLBFjO5noPlIXXXSXtIJDQrq1P0uX35ljsWPc
gaOKldyD3mS783ywj4VQ1OkS9CJKJf8R4M3BQU1JIjONWT12yZJk5Wg9fh67V6NMbEf17uyD/mhH
hUI+ZZ3ORrggExe6VRiexy/FMkAQXXGYuVT6ORNgR30JJw/s0kbA+TpK+wA++sLUrx3Km+jgMKnf
WoM5Vrreht3QegoSFnqs0bCSG3zx8jVGsYna8sNqeKaTL7e8T/PGTWj5w0uYaiBApI5LDMABa1Af
YbsNZjylr6220Rk1++eskiUfxP/LvjX+sZcjW1bj+VvecrQfwZyE3xrumIjkGNMokraHQ2jYgGWo
VwRqlyDCJYCZbUA4w0EF7v69XcrOvYBuosh0w1gJxgxj0qT7N+1vaP0FaICJyGBUyKQioKamFW9R
KTbj/cXy4ZBxhRPCqli+dGCQ4dYdQEKH/v8WiK70HUCCwvXzTtoQYzLJ6FW2QHLdKKB9zVxX1d8W
pGsOjzx24y1qs+Nqa/nwdgxHJ3lo0l+NWbmXaNMjrZtrpcwou+oulL8yAyaAist2UVPoW+tzkZCU
ep6m2WOaMuEwwuoZO07uUFJj97TKk7TPCAZoQwj79e+BIHIl8nHVyPdAfq8CPF/4eh7sPRVEacn+
H/IJgtFN3wXKmN5bSldtkZ55yvscdOVan8cBhbJZvQfLEeN0cMqkjP4lJF3AsHweWR1GsIQUt3+m
hdyneSuQW37480XxxtVRZpdnnOvPCBFwHof1rXhbeMdfpdLX2ocuwxok1yMiO09Xal5/lO5cL045
10iVEncmBdm9aFBHJtk9Oc9ZK8ZY1FqBuScZ/Nw4l98vdEWuubVYymBlbdlpPAYoLn709ztZBw4n
a0ZRCP6iT2f766bggwZh/kadZAEaUVbtEWDd0AY5efXEsp+eUcdsc6SKnzq2WDHCzjEyxshyXc4t
SOzxFKrt/RB/K5aGDU/shhs86hX4lPyAhjHnzBLLcRdc13tDMCQ8RKhu+4EyAFQ8t5vsfkD5jRP1
WtCwleeNF7sQgXwzCOBUcazcZtJRC4d5TmkI8+yWCkHPqoQXSgfGoe9i8wX8m2H2L/cjwA82Vzeq
i1/mNSTRBYYOnIUHriYO+1hCsvDSGMzM1Qa73CY1gX8gbt75vwadMOg63lKemmE9wkaqlzy1/cP8
9AAv9x/ZBW1C6nkND/QMzqMWsxilpllkmbE3e11PCJP2zEsOf8hqVSfUUSsYwzH+g31qjgo0lN6Q
s7feEeniicwP1RJqlFSEJNE3IgFHyBgeN/mamKuBb6E+jFd55t4mHTVpdVVR07pCYTldcIwz8xvR
/RWlZQWBA4AskxHCuWiBRn9Qd31F87dvBDnT5lcwo8W6wXfQ8/Rr5wVUKSqhi5Cgio4qeEXfjC1U
B3plJriKM4TUqfxmjHNnsXPmU2gR9owIQBWH1G1Aq1N0wVAMe+52DBNa+LCiN/z261LARASFXESW
GkIT9YCnvMLR124xGKCRlc1f1oKoto/1GqIkulRsoTYIAyAkB88Lvgf2eEjQhBJF77sLU+yiyLa1
6ru9KnyzbTuJpRj4Al72AdcyxgNjRufAx1Uq8vmLc/Kp3zUxC3c5wx//YdBgJ/myCAyVgfbu9Y6J
pmyIftqKF8JBGhfuFv4QjJd+4/7t56H4qIQu6r7jYv05VfVxwe3rY6dfjijx08eY1zSbKuYCoCx2
ze03qAnuBP8aH2V4PW4zivv1yH0mkPSXHbT68cSamED/KAGfCebwS8Andwh1zqgzpam4ex7+IEDO
ZrqJKxDwWzChGRybvLE/INq38FNrsqVR9KrQWw+9WTnFZqbnwNS1QIeRb6A9dtwIqBBEg+svgGh5
EfiZaCXuurhF6okHi75LcXjU1wtM1iv4lupRbkrZfIHcjgqfpNUrCb69y2ZBM5s7MOpvWRSAAgxz
f3v6k7fXYBK/KqeDnHwxsLz3L1+MiOxkj345L5ff8adRa+zlLpLa7INd0C/PkXoD9CrgBITSDFmf
pXYXEZaOMpic65VHqCffYOPN4Y5ifQs7nWJawmt4fK1nwlfjYxq0mkSA6z1mz9rGCqxnO8kL3/mQ
pmxXO1U/8tvqlh9tiU+yVXq00jIY28wjourxJ5nz2Ectv66FBmuH8+j+tr5VNQ0+QyZBPQx/LpgZ
S8NXDkPHX4vJTtrWu7+2br7i7iGb6FUTbWeZ3y0LIGQxM0bFJfqdFibccIf8vON2vuzLiZgcp4x6
UYWCRmT287dbwcr/SOcbClT+YosMAdEBYldB1hsfXj3MD43+55IxJ2wqwO1Pd1Mcho9FPOqHH7D8
xP44fC7NNRHA/0jJUfuaIms3D3BRR/L6bZ3/sAADPRku1btPyHU5zdN6sh3k3I9HkNhB+Ol1uXwo
L4uaL6pSafEzJlzx5tLkA9cvrtPUzGf+4cvKAGyJO6wrfK9+nh6iC907Mk1/0zVlyBJs0PScblL1
P5oM1eoWxjhzpHRFtXZR6vzEWDo3VBYpbzmRB1fJ5p6QIbvdEq6Zk+90vU/R16oIDUuMRUMJt1ia
1tyMg5kZ7h1w6v58yMv09mnQbvgmXPwHy64KHk0lN6gIi7IKGyLRs3W5abCqpjRo2yMuS8MtQIhy
LhZieaNLtmtjpY2h89pL93OB46qeElI2MWEJVHl/T7L+cKUo6FbzlwXQJ6QZDXC4MEZcG4VAs11N
ioR244XkUlbVhYma2qTbNkjXtNa2dlI4ddb18df5/MF2xVOfyksd9ArmYSEVIS0LtfJMr1/+x4ax
5wArRkXKYrsLPdsiA9PQ6AeokfoXsezfcOYUKdb9xL84FNPKmCnWXbyhTjldRaquraxIOsL3sgae
ec9HXA9xuXzqOb9VIn3dPNXh46ueMS4khI7H/x+53WxBsUzrc4nzcFKrtCDZEgQVasTMk1LJqQVe
cAt7zKoVZ2hJSnZAiBFyCDfKpwIw5/s6FWcc7Ls673vuJZ3MPZBDQUJVHSiYEZLtreigq4WCJg0U
HRw7mEuBOJ5+eLxy5TleznAp28bK2NWFcPjtopNcwQLdg0ONbbERsoH2e6TajSKWozflPGbEH8jh
AeI780x+gQcFNa+SOcR1huOur/fW4zxuhla4MA0KIK1tEMD8bzDeino09OcNRsTSbVckNgtFzjJ7
MUlRxzWvibJBhnU2nANpVfHgyPKTk5wK+81jS5E90Xgw5rH/AZjG4ekzCYqFAlieRrv16hFhmBvL
URxNmiiHo+HrV+c367/Ixzqk02gjX3gRvluVZBDH/dvpjUgKx49v8MiD+xDYMSr7g0ECfseoC+hx
hl1PNXjrJ5JGPt7RO5BWZ4ciNkQ6QB5C552ZFRmlgjMmmhV6kKKIjWV2ons/IglDr6/5+9E4eF9m
9DLY7P4C1kt/7VUoGukKIn0ChCu+AMX6Z/5v6hNAiXYcop/565C2l71FpkMQt2DPP4FdkWogedGa
89P6cCRN7Pv550Z+14Ae5oGf1+Xla/RH4Ali3JndNwdCLnSEnQYhXVG5fwBUvqedHrj9gfDMf+Gk
meh9csDDfLrDloNwcjhgKnR4jUAHHJMQsdGSXA/kPaJ1wQs8adfDmOzGfxKJeVuc/JJ+/Ow3FRWc
HtgNzQxS1mG6zYfEuRcl4/jdIDquT5lJhsoousieV1/ewlBKe4IrA/xBS+SFueBRiVs+RRj4Ei8l
zHxuw/av7alxPDNAboGzUMEU8LwkZQzSUY5zzovWaRRJ3G5IbztuZ284AIBmZ7bZU3mjx1YzmitV
vjItCST8gqZmThnP//+oDGy6Y6cnjKf0HUM6qf30m2YKD9oWBNmRdf6wyXyzecrqaY2bejtRh8+t
JVy0Mi4yIRPk0nJVuxpSSNeGDwAsvRr0LVxqXyJwVHlyC7bb+MAMp2A7TDwdAlIuody8Dyt60xhO
t87Vik4fg2JypFF1TUO/bTrrroGrJfNOAS6h03/8Zc9fCEUYCjzVorQMjdX1gUm4aZlj61kql6FZ
yPyLG8iZMuroyANDqQ/CZThiHXI3NQZ7AYmxF7Xxd5zKvzfh7AkTR8FfrCvPAyflOUNxGfe6Y3rU
jHoqeqy3NsjhTRoyPacRcblrkpfLwmi5e7dLdtsPu6xnhzFt4jLc+fPYL02zHB3rV3xnO1I8kLhp
japtLLmyh8ghFeIX/8wfc1ND5yd+cEtVY3gZ3GyKffscskz3VmhjpxcvmhU6w8RSqdcLebQoqQLP
MacsvZTYpJoOt8WM2OUgcaKs8Vb5lzDItuqDk26MK2xYwMElbzJxyY2eMlKnjy1NASzsT6ew+yDC
h7FZ04kyU3QZpPYuuvZI6vTWoeo3VP+f2p1+8SbLCNtUzgg2J9hAKp+mnJB3xTwuRU7+NrBzMk/u
ojJU8ggCdcsdc9okWBhd3hFwyO95Pqwne2pXxXm0AVQ/0TEKipTVY07bJ1CBNSMJnXZUZdcR6Dnk
dDYCnICzGmbtlR5mU23fUrGxIffGhydxZrD0dR7QY2ghmVnKUxY0O020HhokEMjQ9J4w55F7rf0J
uW4ofW1/25So+9u4vks7o8IK+49pu548YWYIj7jfHcH1PuVoFBSopGpSLYQs5XAt6LLpzSEfXQVM
29wqmzr35fn0AzMKtROgfaRYBEWBn2F/2Bda+R4Y0JZeQeEN9hEYS5ilenieIPcE408k2roMY4F9
CSK5qDq71rHvPL5xWDODrETu4+s8xGht+sxmVUT+lgYQRLPrjmPjys6IqtvSFtVWCewy2Mdrg7/b
pJDZTxsfXvnBv4apUBDQncvB3vjjgKtltSihLiw8dUbP5hEPDtkR6KB919RNcxTB+sGfUpZV3IUH
wmVzgW+e8VeT3gXnOaBW3oVx+1eZKzlPfGOQldxz+uVlYcqiqaXnvmAgit27GLN+/7Rjb5agJjmZ
WtLI6xl057f8G7Sw4YvWlz9/lPKwSQK5RvRxprObgMpvOjnRlyYqHzmK0y6q/erRILwRi9fH45KM
tzW3CCAaGL0tGR+wScB2Y+87I1JeMvxnf/sl281teIZ96CJ5UIjO/JhGvbQBonhoPgNjzu3RTP+h
rnpvm0Xhi5jN4Tg1wtbisCHioEspEw2rxMB4d7UoA58SX/VnjGP6jbr2YNKrTuvCNW2SHbHKkqPs
t2sKhRXgIVP7+zoHk1IF4/pwGZUSZ1EiNFYBlvuyQ35cFL5EwqKwnZcb32LCB5VMBBGV+q2e8d27
eWuIt1c1HJt/0ficEAuwGG6jPqiuA2i4c2PvJV4c+k96sZLTZTriDEeMtxLHnouFoPXA7pPM1KSl
OO2+A9/fSy+Gf06DTRhIDuqi0w1+hG8rX5nw8tQ+eQg1Da45CFYeLSnwMbpFlyMaJAYG0EqhdNVF
wfNoXlfgvrVVm0qp+6r+vnB6ddsmNYi7tyg7aGR/xy67svmKbI2PGsPM9Bzn8yf5p5HE8WDrISFw
bFl1JqOdDlKYQeAth506H39SReWLzhKRY1zkyHFGDX2DmUowov+ZXoVX25uPuDlAeA1YtZFxDEXQ
Rd/obHuIIMmkL150yrzceAwlRTK5DGa0WIpfeVN1qsGy75XgHnxoFKahjagxTzPzCjxpAJcLCgoP
k6X+BS9yRlDQXLOUsFZWJuReirrda50DH7McC/zlGtpCYz11KDGtz4DCFM+V+dFdeV4wivk/wZWO
KMCE+WWSonc43N9NjdlJJp7DuB1l7z73lYDbqq30sWQ6wsu45tWH8RmgEr4YLyi+btiAIWCTYr2u
pgrsVf2Exx2xpY0FZKa8k3ADv4zqSXFs8AorVO8wJ6CdN/xLEICUDvV2+IJyBPbQ1uQ/d/SvMzRm
VjpESTQ/CetDy1mEyvgMQCXh1WplZsnVHP4pREnpx84T2nx8o/1UkDvukJsnz+LbxzOk4Vu2tjy4
3jcR2QGr+1yli3++1SsaEXsKnn4iVkVPpvY2skYqJu6BxiryXYKBQwxTnwc+jmNZ+PPPwUMfUWH4
M4JEs4iRiqEH3/GZxO+GUy8VR1Eguyg7UMFmtMelAe31M6o8XZNEts9l4VPYYC+WIUOv+43U32Mb
HKhxdlvZHEyZ00IxBQPdE2xNEUNWV0XUP2uXx/9w+bxqfMS3llNuTS5FI1q6OtGStoiCHF4WTDnh
PdtMsefeH2YH8MhgsZ7mtrlYPUiSXPB0iSHEG+oqlPLqNrPOi27POyYBR4LaEYtvfCtlwP0cpyrz
d85fRpwjnc9/fgoVhjOW2+rkBbtOsft593u105D1JVjHlfjvllv7qzwNuEADIHkN2VLEwQAG2Wsv
V7cn6OTWnwyMK4+VDqdGqUhSMU2s1zcIAKPdcClt83r4s94R4c8nW7VJnmc49QR6eMZQe6xXMYjU
z4SIcUB4yQv5xsSj/4sER0ash8dfwuTrtOkib59y8kFqgz/18UQ7+Dd0JHFkW1PPoo5CwF2DpbSb
zwZJJsrYqiCgP6loQJacPNNNLjKDZoFZnaVDrpnJpxMI8QBb/lanrFYtpkYD6MLNfX6hO29/TEXT
krZ6kEIoZl12S8MXAvL8+eWc7nqBPRfq3aU7MvSmM5WO3ib2yrtNjPeUgEgsD5w0LcAJ+oSk2HEg
LfWUHG9r/0jbHA8Zn54MMrXOkTPe7KO9dIvP6CTTr/v399+Bo5zt46XF5BWj8p7dd65r1App0njt
JgPc9N7zAW8ghZeWViVNPZfF266KmLdMetu/pvqL6tezUcXmbMx3qj82vlVCusL11/30i9/Rx0Zo
LJr4pQwbMo4spTVce8ssbvF6AGc4WGJRl1BztSnHpoefV6t3jMemEA8Bs93zy6HemoZeE3E6yVJa
2F0JcSqlAzp9UsL55Zy8jqPSoy1NiPwchPIh/+3+xAYOySHY0vAhBrJ6GZmgxUC3rNRnPo7esszi
5/I/m7xnDpPASlr83KWKInMR16/G2ZSBKLNBWx+2UkuZQvcWS82NGF50AXxPG4xdLEbjxdzDku4K
KLEG7cOzZaJbgLWUHwefIf4nNLnAT09OIwTyGw2tnC/jZIslm1utsumDgoVo2LabCNHW3evaddIZ
C6tT6MAEO/QJ4iaM187xXlBIwwOEmXH3OtqicJXsxSPJ49gt1TZaA6PRCpfUKJI/ZDEkL1cnXZ6T
n6zEYMmstxxvkxdpUB0taC5I91cnCswLTggzI/VqYw8yWhmyOgGOfdButpWPijbo+b3hohhKXmFe
F1S9ccMtx3KZxSLusouMtgypcJhzm7bj2umohhrI1iueMDU4uWWf4nXfJupgQwSw1e7vFB8EBMOS
CVQGIXBxPOnVJSVVH6HLrFHIVY0D1XnejmuRjT7v7gOAxHINsd3IhdOO0RrT8Oqh9StkBn051D1U
5Gm2yc3+AtKPMUrIbQMxrsw0aheEDEV5g2gM/NfmyByzMLJrkEX23C7o27WZZwUsmhqGJfQjmt0h
x/3ngGNelXNF0ukDVa0km5iOQfCgfkH9YfFgr6zktPEnf3Gxb8oXcikxtxkt+mRN9fZBlzKhrJon
8KlQHvpDZ8jZKLojIlzif8AozdDNtLsNBMY2Bio9GsOvgdEmLVBO4N1FMloaiaB3dSIvjs0m/F6H
5AAzAMhEk3qAImMSqKDekRl3Yei1CKBWANnPXZmY5hl8fuJf7dXMlHts5nxaLYY96zfZjT2wHcT4
piqh/mGecpaDeus06CRFbfU0LfqD1vXasjw2e60n04dMdnkvOfuFpu62fZp1OrAIdE68a0jQoY1x
F0rXkpaW+C4QsHitTdIG7zgVfSQ5c0s4c7LLxdH4C+JWahV8SKxgDgMQPnQAr8kjbpQDnrMCzhRt
ywfSMIUjoBhDt4XjbCAwowCdILbzgxeKzmd2t2BUdea2gnodrsqk4Oix/g92ujJXC3XPaSOWlFX/
AVgy0gTKgyNIpxkFIUUWUEFvrI6Zj4k6cu8JSJjnZK2KdbylOumK5JPQgORylID5ChcPBrdIQG9U
aC3lY0+LWQlWPF8jEolS/WyW5ert23SOWrPRR2CbnnojSatdXazIMw5P6BV3pqBPH/j+YuNR09/M
/QvYomGDqtfumLJu1bm+7xEd6Kv9Ib3Zp8H195ed3AySIuTube0bd+RyfGmYUoJvV91JtTGvfJEH
f580Lom/9t4SqWiKrW6+JPIfPjfc5iwQj1F3YuS7wKcnEKidGXErePWVS47vn8aUlnk9r/EY54As
OErgazQKlilTx5PQCx4nOTJJQv3wKYv9mAVT2O752dEGR6ta4RGGnbyBItL0aXBsNm1JitaG0gH7
ujaOAbo7sct5YBLKGxZkmqWjjBqKnhjWrO/K4fhXqqP367dnuLjIm9+WBcSQoxPf2DtzDU24Emn9
yV6hiGs8fXnMz8WhztizY4OyezZwO2pKh1bN4Spjda5uoEVyuyxoSycoXU1VE+F07/rbJpXtOdMY
n7CUjAu5NOsTOtb3989X7Ls5z1c65bGWkhtburCNHfXAsXbm0CBrMGpTfX3WBDkNZw8q9se/wznG
C++TrxQs8rSWO8XpmUD1R689TdTiQ8BPqSt3xR+qexXNgkA4xsnBTq0B1I9jYdtdsc78f/zGmWnt
qyX02Pz16rQ+NeeefeoW8joOY8022YMwI/ZM9Laff8cjQ/EXLgaRG+oQXYNIp7YpeEJnkTM0B4Jw
3Nqo4htTMJnsWGH5iuZpwdgg2DxbIsuR+iq6a2vXMR1NoRdGvjOYh1vIil5bHY2fpaNDJofRZYlq
SfZTKsC+kVFjSlVNKn5wgkCBXfdAkHiAEVDtX5I0dCCzCghBpOKpWbJfzkXpMRpXFqoJIfdKNAQ7
Qtl2M/u4KFxvX0ci1FjBYryP5y6BJ7gd55jkXVIWB0K+RhQwM0ie700cqKVqfDTqLrlRG4BXrLJg
xz1J7at+N7GpPmowBE970mzTVRnd0hD9BF1tJQj59Q/VXquLW+do5VU/j7yYYSaJwx2dDfejyr/X
vy545Y7Bu+PlTcBHbDRATfptbNX9EwCKlvHEVU5+7/FR9MlZ77YVwcSY5Wfei0+w1ZpkttTwO6k5
V1ZSn7nqYPcolOWj1VdAmsw50U1g6e+yECpfOadvPoXdORxkGc2f5ilFZwB0dyWNaHm4MrOTfxHz
gLRGYPaDuJXwFQsEwUErgHLtfb/3acqvAQbP6uvtKfWlRehYP0/m52bwKGS9Tfoua/vDnojAgqMO
hC8r29FxjES5jCQg6ACTacuZN0AyOTIkdgU4pJo3qIPUtqiG28w5ryiIFninaop3mAENPEF5MvGa
r3ICr8iJWjb/rDBY5qUDhbUPopJ0gEvWpxId284/BZLJh0grChGrJal4XR9F5KXmIvCZQYF47auG
gUIeUORTewf5w9KDlt6CmYE+ncZNwgCYdgm+mqpsd/crH1bg73T88Ch24XcZ7WXcmwniBg7DGzgT
bez0EzLvlgl+PT61pOb+QD6LnmTdCzNLsubomhxPx3Nu/aZ22Ai61lT6SeAM9/VbSDnttmCQGxg1
mlyX7a4NfPXGvyPmYoMd4c9z8BIXhQSgnmCBit82SLMwj6nv56Sk217LpwsJpQHPVv4SzoVeFGmh
wJGtHgbA48cuz1D8GlDIGPcMMYHUuY1NY8/zdl4tN9+Q9kcDEgPJ5+0s9++KjrkXf+umBQDHe2G/
9zvQh3KTHy4vQKwJPijJ3Of8XKVOav2aqj6tl/Y/Z5p30PaYr+Vp9UphvItpMqzQpHo4v58KGiB7
lN86bsCAI4Ggctc3YWqaGJXNA8NedW0sdhGNFsCgGwchCOXBZXbqlsitbmYO6asWBLIwKbC42ADp
vyHTJtWn859lktv6t3qnmeybU/fFv3vNaCObTlZEgu1sYefCy6WzKchqimgk82FOIEotoiEGBtYd
Y6QGnaYKUQq2LgTdLrC3TNb0AkHaw5uYSscPcNp5FdlO4/Yi2Y8Q8JXB9+2RA4W0x3jxIsH7fiUb
UhhRvapMoOywsrD986fY2M9O7BpBw0FaN9bS2H5D6PIpxSq9COHK1RpSo+cGDhpS7W/6kcOkFiaX
XGdL4xBtHZPPKFjOZ30qtwsiI0PY+HR4dpMR1wxxhIym9sw6m5nZpiRnK9l0QX4qBGXxFxzZngjC
ulaoQaPTNMTyBYX7PrP0ezT2VOFZK1nDM6Eund6mmbkrjp4Ixrg/waAGCf9WqCdhWdYWwv/HyMir
se0qwpvTG0eyNRUpSOaqfiTuT0SQzvpou9MklFu+sBKUR5iV8mxHjNZIJpq5+iltFgO7dKnPwXgU
5rsln5fOCtGtM68QxFV463TfQGSYL9u+7lb50JHVtr+CMXnD/vBQeYw2cvDtD+aBaB4BG8b+kzJZ
IZof6sk1Lf4XbCEzyYK3DINtEIrI50TesdZwjvbxEVsqKuwmKtVMVb1HjQAQdjL7EIeuQmxcUJ/n
z4beHGcN7yt/haRCrdlz0EUdEwu4i3lhcAUpMPH4iQygstWRq1UQUQ3P5ElB3NEtcMyRyqZ0G2Qh
3wo9xaISMeaMGspAxR5Gqr1HGxjyMnxd+i/Nvp83cJ8qH/FaeKmzGX+H0v0+2NP3aBJqUK0pbqoN
Ef4m87LoJ0gsNfx0luK2QdABH6NfdIxvH/jxanAI6fgLgxy6gQSRLrB4QfQrkPi0xbiIsRHWRGOn
ykdDn9S6X4MoTA8TGaEM1V6cG02uKi0a0RF26nINTJN1RbA8Cl/Ci8YquV9EHCdLLNz3L8JNFn0y
s+UHt0St7yLJtpQQ8I4mspVTTM4bEJSzs845+tpcXqwuKeOzts/IBiBUXNi0JnjjpLgQwI823LY7
nVmsnxh86G7PV6JIkutla2837xp/C6ZqfJPHYl4BCJ3OFmgoeVd6NjwVfbrT6Sr0iNNLALZqHkhv
pB1Avo01TMsQqqf89C2qL0GTos2ekna8amVNOkvC+araFQq1SFDQc2jsOZKc15Mp2CxKP4FAA7hQ
q1Ls3u0FLMIsnfSkIt4lXBoKPxYeNw/tdXiydq667Cj+uGzY2+Ueo6LxY7JtHAnThuT8Mm4NVX38
+G/poGeOETEalP+bFNSwfBEKO8k2M7hJpSb8bTdXul+Zd2tdzAyFulHK3dfny8UIipk5Hkxz4j8d
OdEOXQrx9DqpqZrX6XMQdTB+rQYvcLdUAEVJiGItj9Wq9q4oqE11MjMdOGMm58yIyG1M3XoulV73
xJgNGORA9Vnz6i6vbdfUpreF0WhTrlDSIkvE+WcVGRQG+gpfVZR0gp34T0XlTSUUiAGFsx7DyWG6
Jgmj7e+hU+Aftp30rA2k7XDozDCGdLzfYOGembh+U225xz4sU68efW/+849z0oI7hmY/CWMcnKlB
9Al8vO5o3QxD9YSycuY8Yj8ZxalaF6e8s/DBMrWQ2upoB5u3kpkcEihdJVtFPIJ091USllQKMMdt
fzmFSZNJ4nmyVyc3M8EV1GDZKCUc1mxwznZPiAfcN4uQjEv+0w0Ae9DcTZD3lMXObqr4V1kl7l/q
bmo3Jsw565RNTGFdYZNnvRE0SQ4/gASQyr9IExjm40Xmx24iNwSX61Zp82JW1Lg/FOiFmZ4aJexL
2ayb4ppxE9ItagoDkOH9OXczJnyGkMx09cEBRPbjZB+FKz/rG/7HjCXoi2RGafmFRlAlbnOPqylI
R9k/cgX4lnhbaCtM2JHs+lg6YTK/j+biDWNXwIMlPcvE6Kq8Yf/gXDHqr4pJvqvN0zrlghtnWY7m
zgNsBhj1SnVBd4qFzdXUT4kcT7Zh9nBeypBNSsdFiQ1E0+5Lc0vhZhNtaotc3uigSUxvZZvzyvhI
yP9ZDrO0h+8VJvYXGIarOBuB+8uv6Zl5uDa2TzPgx7fnPdN08l6IZLHBHH7rDISmIQukynm52sib
IkWOmjJW/pEZt1/wTI+Z7k8z8k/wJQqyQSFuiLJh4+P2xHZXmDJMUVbt3FFcKV4uOJZZAosyXj5U
RPIz2YYhDkVMZxypR/gIOhmWORtL/giZMJDgiWeEsXND8Cc6KJ4lpwngMDDdFHsdgEV0Y7O7pgFk
tQ8Xsjq6BcPc8htRCe6bZuuoZdOmC/w16iKNrq8TfzKvOIpAtfR/KcEqmu1DnUKxe+/YKFgkHBCw
gUknws2+vNqYbkmV2WqPAJ9MS5Kll/aHyZX9QqJ+e7JvVvSOSUxXBCDB4t932AmsnKR3CDI/YoN8
6bdUjuK29I09mmxSE2GAEZxCiynI48Pt684RfOISQdNjJgfvcMkWa61W0q8eeyeGmUOJQGG3blMb
Oh9t0g5gLtUGYQ8ncypDJ8Dd1Y//+sMrkLvn2om7TDY07T5rkPQoQSBSf5eNKw9FLR934R3WiqjK
d9bQIl6GqyucdosbBcZLTq9nk0VgoeJGB6hT2K4lU1fGLR2+S3UX5pmVSwts/j69v506lHr+krG/
sJhiXa0T7TPShmVsZsSq1B4yBrYydPq/eJZIkKYpNPyd9pJFhEiFKy1qwJkKv4ujIgN+l9yE/RkD
hDyOClLPck11+2b7lQ0oo1PCoK9CjY8u+4wKdi3SESmhP5dZNrOcb6UPVaujZsljQxq64MGvMrDq
mnhNTt+r5I0J+8eCyvG3fM2jB6s6GfWDbV0g6rdAdr6HsXq9hDWPM/mlhnVZrCP6RLM3oS0qArNA
J8/jrvM6LrOs+Xp4jOdHF//oMV/8RUIQbkr4Fxyl09b8K2ECkmC92tfQ8gSEi6o+GCfQgyBhhgMH
qSTTDOB+ghKbu4nmZuzMzdbB14BJZ40FZGscDceKq1s+Yxf4ldYVGt5gJjR8Q8rRiB5xQTqaBVZX
7gwg/gDd/Snyjjsn095d+fYegp7sVHwlWwixEHROJFqid3MyeLQCiOYqLHFlpOAgGQhGamDUzJrP
dpaWjUrgmI4FAkaxCFVficCbQgunHramG6tqAOFtFgSgDSLmTGNT7vbff4PDshQJgcWIN9dUYAM2
oBxpAT75uci3a1645nyX8O6cZIQJSKuijydtgSh8Xl9Gewaao+jxo4+Z9t5Yeln6D/2lg1XjxUD8
JBH6IxaFU5AGmlwrjmz/a4N9UHyk99Ne3FQrZZnvA+/jOY2APLdZy26VNT/A5hGMCgfPUYGsk97h
q0BcgKzkKeFSn0+O87S7cyLqzX4+tM4QWhKh/aduDA9qDGNWeFKPCKD2hTTemesdPRSe0HRqegF0
h0s8Ged9ROqo1AtI3fuObZuvO40hXg4dV1wUTfofBJbIRVjT70enhmqk6S1FCY5fdSQIQS2tGm2y
XL4/s/Zg2yhGsg530pJRipIawGUoxIsSbu9BMlvyk8Y18/WoVi/17omzfvhY9nDkUZp0C4D50Cis
GdnlP0h1TN2JULzcfUalQm0L+ukc3h/NnLmLgz0ysq70cpLtc/63plRpyKaNVmEAu2PwydXAZt6d
oKHTURm1vHshFv6pVs7jtEUr/xkOoc1Lk8GEUCMbnkQ77hPefdx+7CyvSOIZVGQQPGfpicZP6mcj
yXFXAdr6+m03VPopC6d+lG1HqwoALH5ao0FWD7PmwIJQU0tIuboquqIIY8C2fF7ZkmtDxLoUm8+Y
lho4o6Bqz6nmPc5azLrczvOLVl8mET1OGf3hgKEKuqrTB4NGZOC9o/4Vqm4+HJYzyIA7x5P+xGWc
2KSc7PuiL8vv/AH+jVU3cGRcq0Gg60IRedN0wHQ6BpGkzxJPHwRrx9h4nXJ5RVrvvStAYWj6e3sN
gwnCwMbHlphnyVde58qaPUZwGMluPrFDZbLWPp96n9tPC230ynJUw+syf9N3foUeMPBxb4hzensG
YyZmo5bryA5KWVK/Ncxp6+obIcyH1SrPysKA11oLFv9emW8B2JkiFz6NnnGTIc9+jw+VwOWzkYA/
ALi/Y+Llop64G3vrn7gtFmxS5FpnCuAZ5DDULa8zpCkdBDDMhhneE/eODiv7Y0MZ8KjrPWfffId7
brNyer1FPQCOmd1cGVUmqNypvAurXj0v8PcyEQ5y2wi9uD/xpaYjkc6SxDOiGtjrRFbfazOgIW5P
8hspxMVuHFaf7Sx1/c1ttD3gXTQuSA/OO6Q5XfBW1GJt80I0aDvOCfaRsEKJ3yUfhidyddkbfd1F
VLjq0XbDvs5bwYzvNu3163CPetH04I5oQFfRUq6J1YebRSFOHP5OhT/V/LFDYjvC5+En/xyqlVex
cax/HcGlRxA/+no/+vZnqFfH+nD0G24YFKvHlJNI8bzRnGmvfoxFZxAm1MgsKBSK+i0+y4cauVNK
Kbt+4mC/HkLxl4a2q8ZoGLMMUy5dLYZWjF+Tzt0ugTj5qKM2QmkIhsvpCVx2+XDAgsIrYw1prhiR
QmJEhqN3KiU548ScQIe1eaQEg4b80/7Nj+9RJ+JlVZXgSYnqHMU/ts3NKcy0f8psChRb6qTM/JvA
PZxrBVh7cljTtiK1SMYLpvkdFK1A+AcFDbTpX7SkeCOGqnq2uvxcvL/uCeacgk+PAHS6EEkWfOz/
V1wO44EkLnh/ayg3bBlYfA3fiwoFcaB3EUxMUzzT4xlLEcFicQpkXA550ErXkSykETP3NrwZGJq7
dHMDVeJCXs0IZfbBPqgl7lThtppCRQ7Lrmyb5lXBeVP4vpORUKLatGkpgkDpaWMwE+L/ZCehChYK
E+Eup6RdDvdHRUSFRYBhPZR19EixfG2M/hfba9b+KticuA0mCHpw7S8AfUY13gO0YqAb14ihOiP5
M7ph0WMYh3GSgerz6OJHuV2PrgPSQIpBW6o6aLkxhktzZFrZoQd3pBsWKefbPG1LU2V5OS9Fl8aj
XFiwmbkSpUQU2qjF37Xcad9NKKlSc7AmB6WTDsuyx40whTG8BiIO6Yzd8LFNURNZ8EAp3azeztgz
TtIR7Il0AgPVjmOeqq3YuJQGdKaUqrpE0AXw6aBPHgCEP1TcQ2dXd8vYCOo0ZdGcFnIvOPZ7x/gh
BCF7ffAoKHM+pxxlqFY98FZMEH6uOyc92U35TDqpPtlnS2oH2TMvaTTVKeHG1TdRpyd2mbt3+eTv
mTTNMXEPNAdYt0FYR7awwYaxB9+SviYUSMouEdXznr65OlHGGheqdLgqtHCyrnWGv4h7HO3SXoFi
JZlK6fpj3H2YypxZcNUBiCFsQr0r9xLatyhnaow0MZ3T0Dq/lX6UJtzrSXdzVOLDJowoMcg1VxjQ
ZYfdo2cOKtKL0gLKBsozDKTF95DpRqLwWbLx393CCMNvyOvKS/h2CGmciIVZ9Zgt3q5NXYnEzPGe
9HOKvYi4OVmpalAj7NT5G/vz3j1FnCPM+isn4BAl+F4dCoIni8uOecL7GlrvQ36eJl/qjeVdZf/Y
SSdDJ0Ih4ygWulhZ5O9f7GcPRociZPbvfl0WwjhSruPJW8ho2ACMMkVyDM5+2Y8T/XrGbClS4Idx
kKqZZHtSw+xoJqvJgP8whdknStAOnnX1JnApRbMaDs31TNgC+qGUIQjIl1RE020YY+4DxnU6c1NM
FSRg6oxk5HlglhyE+mGn6vChAA3WJxwDUOb/n9sNnQbp3x9DxJwMsIZJujXKtcCvdl/1mMmj10K7
8YvqZt/v98g5ZHaIjoBP4wIu9iOvbiQL+3lhfmR1xrngHzk26sH0gGrpqKxC1/FqQw3Bzs5YBfzs
qxDyd1EebKFykV4mOwg/7hijX+G30SqCdMP5860O3jaUC+HopIN4uNF9d5K1ByTklkhbf51/3iRF
AYcNjpdtXd6S7m9wvwj4Yxgu2HAbKMP6UR1CVygmwzp6OFqTdW4KwY4inLL55J4cwcTdLozXXLdK
hdrpOkeDHyCCgNS6rpWmp0px2ijuy2hL8QV9d4Rhg00KrZA4gkTwKfpHwLjXx/8LuPp/uZDFtO2C
RF3F9XmuWed7sLVQDFpaRufO43NUcCphrirgDwsQATGXfIzdYuqv09rLn14T1j/5Ao9F03hNFI0S
W0D72OrB5tCbrcQ7KKbhrSmAC7PzFapfNGY8ssARt9XBs5A7+MtZEnzAePPnjYFia1vh0RR3ePEp
WegfYd7YiWwHPunH+ZJUTDLoR5CxkmVAw9Wdn7gpRlDmHJWODRcmAQSpav29nCgfWESLT2wQJ80p
JabhC+Z96L/bjCTJca6vJpH963Vwf6VhcXFSyx0T/JVxdpd/uD5w1nXqHMXJgMvbHn9qaUYe0DCf
nSWEpW2OrjvnJxQ4//V6qGj1lnzIO8u3xbbbtFz+5dcbK5fBElc0I0Yofi8Q73pY1NT13rS/9Cw9
FV3uPQuz+iHmor+OgZXAj20og8d3le/br5Jwenk3GTYHHxDwY2YykUy5bjH0rHj19GTWvFcR7r34
wVZJTE4L+nKrojJptIT3E6R0ADDhPChB7wZqEeYcLU39QQ0uY5yZaZw4q7q7yCHnGpNJF1oUewh6
u7MC3s8AIsuc9LP9e5Bux20BDlRgH/piOTmOHFsidVgCpiAebS2z8WvO9Gsfg11zvnx5MKM2Ntsn
FKQN8iK16/lEp+kKGfbYcjV/YC+NPzhMgWPyRXG8aq9rY+Ae441OE3x72Pv7HFHKbRA++fKEngA0
XT5tgxSLRSICLLGwsQaC7Ka3mClC+OBc5Y0jwapj9FpcipUIlRVBMkDFLieHsY0Km1mkEe9vplmO
0/SVdcoSJ8BLpbN1yKKSnrRO8U8PCOSeRq4JxmYxKioBNf5jcA6EkR0pEf+x7QuJMEXPfBEeA2mq
LQItdKjJ9ut65MtL2koovznXzP1kKPvuoGYVpmLxEsfwtBH7IHc1JVbWa1kAjAmB/JMmBLG+Cod4
hpEtBrX/xAcgplxHXHoaC4Og8c/UID9RlJGiJdauI28tQHF3k7Zyd3E/+lSn8TbsLdVTzbMPsXvE
lcIUQgmw5yBAlgFTCNyfnjiFh0Kr5/VNVmFJHcdGjvxbjB4r/ta7ryEryY/Fgy5WRzoLCj9TREW+
oAZQGY/2+yYpeF554pdMohN0W0Q8qLg+sFDQtxmF+N9mvCtrlouxKrlFEa5ocxNtry9CKgYlooPU
rA+gYC8b+LZT8phtvRXB4JMhzqe7mwPt6oAlleyQ6qsN7JY3QLLn5z8F0HFWx6RtXSTEf28r4hhB
bbjSbQkDldpj1VrvLl72M9SwmN/3ZIFSaBn3qlhpAPx5x2yAVjClYFSsxyn7d47bK4r43IUwTv71
/hiKyw8VXErSMQZaoGnRwoSlyesvDhGEr3TIxzjkHWLZxmZsyC+Q0UDehNP4tHXTA0Ez+D+bJUXs
W8qmEyrza4s1QhYkYLGtgdTP2RLnANI6Vx3D2Mrzjzdc7C727LKt5aO0V5ipL9cgWHQvrqUI8nNy
5Sje3tJFhZkFs1ZM9nmXGJWJAiiUZRTdhTWvAIJfXIBJB0X3wbKX9otpi3/fRA4UmQf0aORokIuJ
pIrygB8GAFevcanSk6v+4AT474r0vBAVbYTWFY45dnKiuntWqaTKyVrJCe7MULvva4ggbWiZt70z
VhQpHpv5Wf65ut4nh3jajCUugxrbGwHJYf5FscQqH5nCEyT2WRTuWUGtW8Qh3sxUHqnIg8bTizLu
GFE9eQoUBeHI1wYNdI3wc+2EgwOa2vQmPyLjFIabGakAToz8UOzBU8Bk2+DYRZ4yT3OsJUto3gbr
qcXi+Op37rvydPe7lm0fCnqWENPltWxhMclEMyQw8CWy4HGvkCfXgJxfHo/Warb5YrvfDnrf1aJt
yOdcY4hhArdY7FGr5zEAHruP5pIR5BZQR2wN96i3NkZClfrKnwfQu06c+RGC3GnXvVlYEjoRVstA
iIriIb0nKiGyWyTvwtWox/0AYp4Br4RrGrMovlOQecS6YJsi/WI4T4T8D9uNaNucRzRl36q/C3IW
jqQLNqx68SnxtZMqzt9mMcEN/f4C5DTizjQkPWHdy+I0827i/mnWQFQngXBQE6HcvKUxFWwj5pFf
2QSrKp9y6QMrUp/FezA1rAVmbBW9lzlGnZfdElG0NP1YYWlRUHZ4K+MWX75i2R09DiidA6LuQsCF
+lW/zPBBgDQlk5lRHVI+QCeCrNaJJpScM+vlt3DKaJY2Zi9qGoeIb2ytlmvPD/JHv4m+OH3Sun97
hnQnVcjwi36uI18jzRoYve8ImwnvzL8qnncyOVclUdTwcoD9Rl31A8YtN/uosNxGM7wYzQq7nMQs
GkcdjVXhvOTUb+ST+pgrSsrZwgX4I7yqPicRK5hUyQAM7mk50KD6ZO0o6IH/yXDIQ0kvVSM/zd2x
fwAYDgckq0wYysrQ7NNFe7ii3MxU+Olfy0XESB5I+sN9rfkl+rtZhJ94CKt4aVz/4J8FDgviQRpY
Vmt+2QTB8H8KVhKHWYjxT99ZJ3J1Gv5j+2+SzR37CzH+jgmS4n+25ZOf3c6LhBs09+bZ5+fYYsIl
9yJyCyHxMMgDfmmkXjSSoW/nfQ+Qu72udcllmJDyOJzXKrSFhyZsr+apSK1yV/2/pYzJZYaFprlk
zbcHoWQ6Ukn0I15Wmeb3lO3mk512VJ0Au4WXBRfapcoPgXwbjVgKqwcO7qH5/u6LlWHJY/CPEuZ7
Sc4YswfIDTngQ+LMcD8O2OBxEbjW2D4+CHqfRPNaXhPgbN9RbFwCS4yuUjhElW76rptPLo2XiQdF
jpkgX16rNlXd083KG2KGJAUrVc2oAg/kmfo0Rn7aTNUoeYJDcZXXSqpEHeU6p4MJc67pbkb5DFK2
FjGx1/2JnS2mnG5BtjpJcxolPH6BDklY5D67OOjHb5Bw/GA32w5uY8vxavJ+Jb463bURBusJtNJm
e4lD7g7qBOX/hp94FkQlj1Ok7vbh6+XDK6MlI7OkfTatK90GJlQEuzvgFExMAPt89jTWypIFEgYu
+SqxzvC0egADzRv4ebmJIDlbCAmYNe8eW1xPEOuX8+CC2AOGQ+Lo/jUFdph1LDdPEz5Y/byRnTgM
ztH6tqHExHZWCLe6PBfJgo17R2ewMHI7Bw7G1Qo4lxypyix62ZDCpfgBJU6LNJ2Vs9xos0D1KWBN
RRTOATdkQYDz7oD49olBrioDMB+XTbcSOUDlGQzEy/K02yHULRfXwNRTiDE4E+l8kGR3dIUwUdxy
woPiUt8bzGly0GByk9ZS6/5BamkQPJEaYmcdiwCjqR9r9u31bySBRUef/NsAu8d/zbcCpr2/yMfM
YR0VTjVlJL8/pDSJiw2AZRNJMJSZx3vOCzTpyJmDwcTWyhXvL+xHYiHWDBFU7NMCIeAxQ6+TCkXK
q8m0mQ16aJEr58LybbBYrsNRS4vwAaJS03BJwU+JWt46ujbbQIa2+sW0OrqKCLl1DuILahBsXpV6
e2he2K2qscuBMhNeOL0LY6Ksm7JPuA7ElNjJxwGZboyie0aRIA0ueJ7PLdaLphxYytXl+2w0ZBmc
w4TKs6kXSO49syDTd3TBwid5l9PZ+tGOX4MVFFJNgmXaejkMiqJIxQKjIXZaCfaHlznMkGdxLVlS
aFCWtiSCIDd8Jk9vgx93fD7TBZbsUZ+h/Lxg0mmZjWExyCy8JD1uPyr/3FMWF9FaO0qQnHceRbmU
J+c4AfxXaVdh/mLcqtsrqrxcFzZ/eOxNaYkLzPhvuHBwA5WcNVqX+lL/9IyM+ubczUnCO7HwyBkV
DxdDpXaJIvzD4vfdO5xYdvwL5Iv/GYPM6tdcW6SCe6w2tzdMGuJbVNx7PUw0nfasCjxdHbTgXpab
T8OkiEl7ZHS//db+PfZ0RTuVrA/GZM2nNRQklOUhNnQWxa8Ch0EmfdYzN3SsMa73M/yfZfsK4xXa
Jger41KDS2qUlHnwpWAEefeC7NYI7shtRF2CbUUiX0AGLT6Ia39+0I1ZDhcDwOp6M0ufDhZj8ajY
RzBGmnZdaXt7+i7VdwSRN80T3HGovqSNrHvJA2SqjWHwB314Kznq+woU9zOxTQMdpQlekJ8CyyNA
Mc841rdU/ptf53z6yNrOMvcWmy3dxKtTPRLnr9WlznB2mMbx7YSH+/c2p1oNQCIJUwP0m5kO63B0
S5lCk2FHsXxaCHqn7LEuEiNAfOwx/OlJT+z1/wdGHW/373iJvLEnWKZAiQM4Oie9AHlqhvhjTprp
4DwaCxfHPvoCJ6Hf556P3oWyyLqeZJlDJ/AvLMImf+duiCGpOnWGtKUevIWdSyONKnAQa7AfREOW
cMF7sU7cWY/U09bxWqc5TwXw5XACZcbHEDkoPgCpMYOexLyb+ybmu8F3lx9scMCzLtc0eQNwGUix
tyDvqknNmSQKXs/QVI2OqKI9cHZj9rvDR9ronV49SuFu8/28FouD94vr75Uwpl5S+VSjuvAgtJPP
0TOpJBCTibcxf6FrCwtVJe2dlsOnS4aLQWFjFweIWLJgCBhyCs+iD3B0i4cF8qkMeWQmsPFYPpaR
4OLAzAztXeSmKZpwuI5RKXx9fQIQjQYBhRp8Zbq/kibBduRsyPN8SUUXgXh+TeFRij69cipTFsx2
qmGqt1/o6wmsFybUCvzo6IVKT6G1mKO2cXiLcq8fZbJPXWOYEo+85/88V49IPtH2wl91rRyODOfv
zSybYQTlmtUhQDtV3DCnYkSK8+EpNkYnpoN+nSYLf2GlrqreZmVyTVEDlB/SmW05Ih/jdC+5E4Na
XHn3ZclNnjWDt/E+BcCSxY+GoeHxbUDxgf4CxHBizD6JQwFDRnCYceqF7Q+tkwEWAdGERYYWRF6d
dWCNG9w6cCPozgwW7ITaanF7Xp53PgdMs5g73zYQ5jm5pdeW2Cy3d/HOPrpO1XLJsFg6CVlKFQTM
2QOypgdnhjFr7FIaxytbeglH8VYpcf+94ynIvrVS+6g7HnQpacI+6sMUHBV5ypn6ql7Gye+fuW0u
wDSmO9fKPgfKQZRJE/ZfOassrHvUD3BWGyGmls2bNqHO9chWnlLas4IwHwIi3nWvSFEP+DqyApJi
zla236Zizt3YqObasrtFx9bmJHHkToinSL2ThlgkHQtiuVn0gLDdZ31sCleb3PLXKd65KgjhWS7I
WZ8k6nVagzGa15WD/dNOJ7+EcM7KOP+EdO92ANld3YOM23Wn/3qIuXsVZ1fr0wEd6YodH6PyPIcR
+xURqNIZ3N8yjSKmr6huY5teSG2ty3BwoOKpZjo8xmshXRe3bHVW/9qnDDN4lw+gWi0nVsAl5kKA
HRLK18KXYGve4CQEaYiMsDUUjmai5Vsw1+j9JkBuN7zu9tCdRzFH1RAlhtfBk1TRcXSl8IAMVPw4
KHhN2/6zvzvnlcifdKf105XazqzEEzgAVelch8y1uD2rgC9n8H5wKgihGcM7gKXKhvqzQFbb31pA
LSQyepJ6jjDjtlVnjz2pxV0m7V3PFRLdVXtRutSbM0A7voEd/YN8jQJwLQmLre3eFIH4NxBfxMb1
rU3lOcjwwnFA8WLNAnPeWeFpVcY283kXDeIQLz1JiN4WpatHJ6DXgyMbuZm9A7O9gRxG/0pLTcOe
2jIreFIaYOjd0kBf8rOZeJIus1f8GWLfM32TBvKOt66pR0DOAJXr5OugmeCG83I5p6qCalpoDaLn
ykJhYTts+czeVs0uRjAT97mbzxlL6fEIWX5CKwNiM/g8DSSzW7tEUgFWoM43BFJ+3Cz8YbrQeNzp
NvDKO5DGAtmy3h25nrI180V4QtEvhiAeg3L6kU/d0HBdMy2MNulJXgs55oXqQn1mhh5bvCwETA6L
qs/NgezL/9P3qxdL25+rWTAee3VdMutluS08Q6un7DzlTNKNB8V0btYtflfAzFgW6/gDu4XNrpPp
83E5/B4wYA/4810umv9VqDKAYdSuekVpdD5F5zVmRbg9mGeTfCQ1aw2EWIUt7nq0Mf/f5B5fugPX
fMwqO8aLSJIOvOoiGEMFliedPzdeBOHJ/VVxcCJ0Av47wbwE1qk8H1TYMAxoUa0NbNYiZLNhY9KM
P6LbVviXZiDiLTTqttf/DVRUQQ+sQ3xmOGCy1iUcAzf82NzQ3CyqETBej2B5GbxkyUBrgrZsoXwd
eK27PtaVO0ICMQ+4MFutJ8VBe35JH0xEpjAb1IDQoWUenyvad9qD77qa3yf2b+rH2MluuITJGgHH
XAfotchSMx9yBFOQ8uOwtWNU3QA/70nqSUmpSN/pxOPnHHiMSh/GHHc1NS8lN8htBgKEYo+UMRbU
xRPzR87q7vG+ytQSQiilcGrkfDA8MfM3RYofxSZKwU9jSvgZWr0QHE80pz9Ed3sNbHlXLiYc8h77
2CDnq7n9E1bjYJbyGlxSOLHAxUQNExxJJ8q/6v8qbLZ3dyckP8dnd36GF1c9ApZeoJfgO67xE9Tr
ydPCHG15ex8JPFAIp6uEP7b+YDrdNLBKyNsyoSXgnmLl5Bh5/STeZm/IZVOiB+bReTZkXOPEP8m3
5/piOHHJpc0GfIsa60LItP8a9dNOcPICTOliQMORdnhDWxGiXjMTPaQ/Ui8vq0SKm+EfmsQdecdg
zQ75guxng6uOQiOsib8rOgznZfWAigbWwgCfYncdNHH45ut9ocNsl49DGubOyeKwezy1wPh0nTCr
WCvo1yJIcMGWsz/SIBKmZRmuVt90KeWVexywtNF3LJAnZhMQ3xRfHpHmQ7o5BHuSZY3bDlY+0W2+
WxN/LnVaY/UEg31IIUO09/9vyoG7YRD0Y0bRRTE/56Ky36u6pjZQmfyqArcsmtn+jvb1oRBPfFOA
GFz/asTkHYG7RYWLxb258x2iH+6lsL9RHjgCFOX20ehQSiMBARt8ZHjqU59X+hNIyGerQcYeCDbo
iPNIqtvRMEJUZJr4nv/88/9Z7rkgU6mzRRFm7+mc1guHmzoRvC+PpY6yLLRQkEGb9SOMo2jstaXn
kMQbSvwzDXfun5YomXNSN4/hD5/C+Jx0+dhTixyEGrjn5aIeYDepjADix3XILkA/RMjiA+gPkfMz
KkUTePGPeOYsKZHFqYpOFGohKh3hsVJoGSaeJlz4Ol7v5Itfw/raZJeCuUtPPZ8NXV2Vmae0yO0E
URx2ZuHqcAQy4G+03wyqEWWQQVX0KZtLEy1OmKO70/8/bT5AEi7Ac0lxZxjqAbyrOpW1c62hCCdF
Cy6qpTXtVxi9CmAC2mnI4R/beEMcJo62IN5OmzASx//0JP8EFxcQQ3eGSLxqINKwT1ejsysUkiQX
5nUNSMHk6sn1vBPL/IMC8aoBRQSKNBMw4gqb/cdPnECJof9R8izQh1DIriXv9e4A7I29R7+StWLE
MHM2wv/Ef2e3Qt+lAwCO9OIcH7mPza6J3QFNPuUZ2yyQPLPKUT5FqVpGAD2x7uims9csjXYnjQ5C
eVNfFVwh9RkILNF6uAj2+tC6sv09pqWmOvpkDHtZtJpG0aUiIiOaXx2pFgVzUV/ZKM8kp1eG0N3r
boM5Zr1uEGv/Owwq8wVjy6BxJCbocJBlNukRF89zgeAIaKepXrV6Y7aEp2D+ECKIFDXy3gTSI9Hh
6NSoYMBOV+9HhHOQN6DrEQu33gq/QYnRhi7q5OLoS3tzxXnfHOcwh9YSihtRnG9vO09RjgC8Letp
+bk8Def2rZ8qRVlSZYiUI4hqppRTmXbReN9Oyjo0hqBrSL9rerQLzoLfigG6Ccoq5KkN5xLNsO9o
zdSWFm5mtW8F25H/YFRolhU0PJvVqXSw7v8hCROopBVhOuDIDdhj3LpRRo5Gd2V/nShikgvyEfUZ
wVi8/zHsFVsjEtoDB1BK4q7/r7oTRP8Qoij4m71jP2zVjYeppcH8IMPHTtVDDzHyyH0c0dCQgrpa
9BvD/zlNgjzx2/qaCs3WAcU6EsY0LdXBkWmZkx7BWjqSbxXz8FRH61Q5hsA1tmUmdjWcvAE4B/Sb
U8dOcj4PSixuegz3lzbREmS8k+K2jJgBvAKPJ3m4nRwhE/Wy9tRH5ExNd7Ct2sxrOzlT5RFruG6Q
aI3RmnRuTYArlnmEbEuF3kHLP3YYmoM/SD5GEJy9niCk0mfrHv/duiESCJ2PaMkVgOPRm6wKR+uD
U5uwmDYfqGi2B3ZqF+J7AeSqpixuQSeWqgTqk2uzPndYGAG6gB+MOVcXZmlNN/hwGLpAf+bFSTRM
jdCqpmfuGtPm+Qneq4PD40o7NFLc3PoTR97xP6Bmmfr+/Z2JzeearYcZ/k2UUoLg7O/c9297Aupq
80T/NrlnQB005MOVoqp4yHsKuaKb34W72V+UQQDh+qKj3EwLU2/hZ24dM9nQFZcloItry95CNIOm
GjXHdpeN1DqNzLfT08qoshkCiGht+G7RidLJvW4fGExmxrKzFIq4DJc/rvHx29zbrrMN/rGfWIPo
4NlAirDnChwoTiCx6b6Eb6r82tUunHSq6BAbIL6YwWg6xO6uQx7EovoSEW/VHzrAkHOhFVKdWORc
uVEJX1RzaQwNbGfmCLH3IAzTXhxnNYVt3BT3pGkXIJt2S/RFJPlKCqSxVsDxV+G/wPhsAxWos924
FN6RGHiKYSSi6C7OHPvdCH+8syDiZKCQ9B/k916cmxLMPp8tHycC9BeJG0m4n0hh9/71uvRTIlcY
jsR9Xvp3Xig3puxCgQt+24FiAuPWoXSxUlzxGJwkGHm6al65IQ5Z+uDsqETrAtdjvgc1PtArNwn2
9pWQR/Np+l9otshTKhBxXA8wn0DMIETmE92TRY1PAhpz+wdq1WOvorLFdh2iAq+xzzgfd4FdjsvG
/p8EVSXEFsVmPkXU7TPnpzCVAOQhN8qR9GvlMVe6ySqt5oOW/e5obx3I7wTfZt21D9vBZIlCbliT
7bWDiGLiR4TtyN0Gpca8xvW5HvEBqlC3SMp/0dTZr8ZxAIg/3xLvW3EFAZBI0GS8IH/+x5FUevHt
xyjITWrv4/nUWMfHq5SReuF9UgtJxgg6KiAhWsqfYzYPRaHr0JLlVHvODTUkH49Hkbcd+zgH+XYj
wrBBryuQ3iWbbCzp/qlcfqO4SBgJFD5dzvL8QMoqEEu4mHwWR4dy4N1jpY3v8varwT3cowxCXMr1
Oc4Et1NS80MiijrppJ0ETAuL0hiSKUVpeGZLn+QhAvRvGhQWhdG3UUPEnBfb45bDf08qZYThnNk5
y6kaDuVREKxAvzvWr+qYTIku/u+XjcQuPJSS6dZTYZ8U42zrco9SevNYNbYk+TzVN9CIg2Et1veA
TmO8AygXmcQ3Ale+49fIYf4g0iW/qD0MtB3yCQG78LkQb3nFW5Nx6GE3fGa1GjC8qT19i8oGbKeF
IozGPR6D3e3kQsTDoKVTMOXWQn5w+g/y+U/Ii2NqR26SwXHNrvbO13rJQ7xbnbuEmMZh50VzZ83p
Ku3RVFkIp0A5rY3XdiMdhraqz8JJpjLEFIeilrNncgPoUIjtSOSQN6IioZ+RUx+OO5Xkez4l4I2o
QW1L6kMHjMLyhpH/NonbECeYi6nCiNVVYIInbM2kVbAtoP9KZv/aMD0HcQQHtqFdvKtVKcq6JYYc
NixyzhGTrcXxd5wD01EfUZwPSAwchCXvUAjz5gIDk3dVMq5lmAqKhXbW2v+Shk7HPURUoryToFAf
J6FJAIAT/RVVLoIeB9KbYEH90kTVeyVyQ1QB4QIX+lt9h5AGbEwh5czB5kX/dIQ5i41cSSphJZts
9rsbPM2vnVwuJ4h4aIamnW1L6R/lkuo5E4qY6gFk6wPuJGACgkS5u3DN82EUV3R9rB2SBp2u2FjJ
0L8XFxTgcAxLY6XreyCOEX9NjsP8olLc/cXpHTewKHfxYW6yAQQZ1+HU1ZVim4rMWZVjEOO2K6HT
UFVxD8l4bfUkrurTQOlBakF7vwGTh+9DD7hUVAWgowswe4Lwn29ufP8STgbhWo0oxxAmGFXtt6Vn
h4xsVhMixx0DqA4pmGE0ghPJkLLkHUCAYlqxPK3ZmaESSC/zdWWQCjWIcnofVnEJJvHPV0waNy8g
zeExb+GE7pr8aLC46bKw4LghjUfSgWkNhi1hShdB2u27nFEUEVCejdabKcGoV9aeYkF/PtbDEpF6
L2RrDTmBj+3N+xCWtnT9klDRhwaYZWmOAs0q1JGGOzAJz28XYyM+arRluxiMRSrXPQT95EKk6VbD
QTZbN7HPvXIRQegP6IvIRkkLz399yjKLbP1+npToqXUcGn8WGtcm/aIOa0JL/YPcKmWZDIVL0s9x
ctaZzyFgAJDO7SZr5kLQU/bVTaGR+KMsZ9SBRHLEeahMe0eSTpmxLbzh6bcC6/hIdm3QFSd1ELp7
EmBaBjuS7GDg/3+h0RF7q+wN0Iz6gV4jEy44tKp2YbDOk4Wj5bFcqVOPk41i5wI0BtMFNRLCLs5c
0PrGkWzHn8UOBNjg+oWqVZPbdxTSGPP0O0cFck3q9q76pMM5CcgnsWfJk1ch/ZL6dKJm0XRtdijI
XqvBS0b70qavhCAng+b9/fUGN+aaUZGMwqJpkRq2lxEMFibxLWoYVWF9tSPXtSkJPe0Kh3LVpwGx
PJr9V/ShplGpWzVAbL6TynPTxCMxZ9TxVjAaZtd7fg20nX8klGx7dhMZ7JAMWOzLcLcIHxJdF+Bk
5QrMbn/dSrNaU+KP9A2rccrirYBHyJRFT0QEJKpBNjQD6cyi9YakiqyhKAYBQkPBvqMivKV2LEr4
q2Rn2fUBdGfDxHgc72hQJGVHrHOa69COWmCuDDcRc0bXBtNtjXwtC1IkWSGx4sFArAM0MM0g+FIq
KrzOIhpFEaNqcWkajGL22L1I8nsWdnwQGY7AYu6UtGiMCN/sm9bomt5UVj8+4z5xl9i8aNdOwhv0
nTFI7Wvqdrj/IrCc4Xp7wqpxUXGFeMtk9QjtRvB29dG5l3agLRl/PKVwuzgGlCBsfDgxIE0litkc
0XRvR0fb5rkMIq7I/Gj+miGiUGDW3sU3gLh7vh4bxPT7tEeyRapHprkW46w0kdwUmgGJz89GL1NG
mwLrLnsg4daP+b/SjOd43gn/YZy47aXH1fkE/LC2ATpagtWkklr2yMfE06f0TwK7GFJqcKOsHkIw
ND7b8BhfTC3JPN+t8fSYbGwrIG7aBPVpSVeclBdgCxL/d/zuVToK9pH783TPb5fBd1S5boLwfRmr
RcylNRF6v2YcHVkqpR8PLydTdNQAxxlixjRCEhAIXFB/h9XJKXDgBo/ROWmWgGNOFfQ1d7PXY76u
AdfMImkT7cmCJXtt+oieMBr41N34zCvARq+nErgnYG1nc2Mk+RJlomkx+3CFa1A7QEdiq8u6oMMl
9t6rgz33Qo7DmJ6nVvYw9c6sqkeLQ6KsqRcY3S3Tl/3vc8HlxggMF0fOFhnXEvinZSr3P824+nDT
JJAIco9c28BrDXbR3GfsABRQf/1tOHc5ICqXefUuLahHNHGf/35CFImEdiAxc+6yB29IikkBcmEY
wkg7G/TdXAp4FlXu9xXej+xFMLbELuXAGZGSInhIijh1IW1I9/0mi6gQwSQdb2H00adtehlIZmre
wPPm1LmddwFuUt67Swy5xtMmOGGHfHzXYXntBIl75qIhM1kyqR0IKT83Fx8Axn4r4zdrvoapJk64
SvIWju8tJ7gi6kAFHW7zjq18H3Om5SE3bCr0w2KN/WUBins+pV5PcbonwNU//VSJaEVq1hemxIk2
Uswb88W1YhMNnuEcbL7GSL5pq5yf+3wstNXuKOUAwW5VvgJozFgDn92eb/wV3sKtTlKrQprpJeE7
DectdWWIHRNpytlVdGRe2FND+gwFIYwCuv35j5ZzMdKnnHxPTtKNKzbVPnFszbiAMDslvQoXJGxo
eAHdlpHR55dmXqw/YNx7vUBMGL+nW6fsskrS8wR5za3OH5gSazNCcfE5nb1nH6i1VtIakjXW2BV6
FE+qojfuGv99p67ttAu3gZl/Ldp4LO7EWPbbPd/p3BjQGa/7Nsx2B8JcPQVz5ytRstG43KzFvBWB
Bad/nOCTxbFeDDU9oVlYy1IyVLLq/0DiOFzUbzPeiwo2e814wnSD/aa6aFePIuvq/3Fk4sx/x2zq
R9jC9XcdEX8E+wnN8F9jZHYMLZ9bBl4BCyhn/22LWaOUE6f5GP3bcu3KaFK6f2h08TgGPIel7AVU
57JH6BmuIuYN4Yc+dNFOUxfXwKRJ3Vnxzvr0pj24QngmURCTHeS7ZuiScvKDnP2WwMUo8uD9AKO9
BpKizuYa9qqt3J2rFStMvseIYU2UAKNHjrKcs5vb2NTlgMi2kGUw0wNHxfmo+3IiZnic5mIKetXl
JjmPsvHJySN+/2m2MQz150x1NTAU5SD6XWeXHMB45fD2joh38iZQFM6aD7ojWSGNj3D5gW6o2YWb
6Z+kovdH0ETukAVw9SmuTF+tMyQ+9XUvWSmDcL0OaBSdJhPBjpe0UaFRuvSehJhXja7rmRJY3T84
K6RoYf3Ip6t9G7GadarDrrMnn6kO97+431Zm4ZAcQXicEdAvcaylUCzLyALk850qzUeDPtpW419w
tbaNB6+6E6mduUuyroW3LOjTFCDG2FM1Yi+es+wn9BLyZW2Z5SBCAKvmrL88pzXBGVj7y4KML5PX
XiYWEfP0dynYiINtSeI9ncx2bp28RqSObiaKqr0YarIHtzVeFo7ZePe4W+pFvNKhvS4V2i3GF3qi
0D5dwTIX8necGrPEhMWIXHbkH5jKaUIiSAnw34277h5rPScvH2UkgBRhDgHw789zVJG0OPMR3o+H
Zo0cRMkCxCF5770gkOb7wrq3z5uypcMxYqfl352g4fcZ1+7Bp1sIendzwgmyvoo49cw1AjM5GfTs
3tJXzbwFNWf9bTvxD2SvrcFerBhrGXGa96Yic0gkyvjnvOIDAsWvug7lZ+PIcD3/gb3HPBxp+Otn
z2vNu9kn+4iv24ion14d4mBH7KpyuFuPIhz2K725Gwn1gSaVYdmE7hq1MMHjbfsPf5eceg+5R4Sx
c6Q5bVuyIP/CyjvzQLaJKVmTKY5F51xSe0wQ5hG0FtvRU2JxY4CydxKNoDlEnYgjqNZ52Irt2nlX
hLe0gP3zjl0HaKAcy2F3Dpyc/dtRCAnABQMfCLrsOCNddJHV3YM96QmnlCXqEh5eNNqRR3SnMBOc
xOaoOG8cOmL6rDzH+p3izqccmhxXomelkwVwizYLAu5qIrPQw26AJuY4FRZ/9HVCG45JTDq6aWTG
bZ2cNdbR1TX2mTS4IAghR2mLgpl7PY3lxs3iP/GKFtubjq/Z4z/zS9+4hJm5AxmPyMt1gSxegFkk
02jHvj8tcYv2bNJfsYzwdbMev+K/xj8zg8x0hQitYGKov2sXNHSfYnHpd7Pm5rKulbqfolmfFrLr
AzaO5C3w/glgFNQSwbNGjomjI65ZF51GVf5XcZJXsMeJLusviEiISOAEJojg4hVkvfep6QDoQEV+
JJ8+5/tu+S9LQR6+u2mB2dBB9qkhp0HdO85SWiBeVeqnNZT3TyWQayrxQYjGsogU/pGe+/aPEtac
XyxApazOAKPoxJXns3Nj2y6EHOCYfxcfI1gDZSUhqW5bUR/ZbvaLZzvM+C89n3bg8tj5GR+bpVSI
h6pXRA9nSuitoqmBN+Foc8S9dPs3d41aoZhdmE0PVq39/lN9bD0RgA01WrWoUqSlnt08PiRoJRLa
+BoAuwIo1KhQxriZBhPBdKExUgEpQrxy+JwCLoCjeaViU0jnubwcC2rl8aWkz1YT4fQIng3w6FNR
WdA/ivCx6nCIQnSoGEFaEklBIal6IjD9EbgEAw0sMVzmx1g9m7JOfG2EvVr3jB661OoY9oEAygY3
3Sc0cTUouKJxdXCKkhi7H/zoqyn2iGOv63E26d4+/TWdOLz9V+Sujw8ydzJytEqrIbiKHahHvoEQ
n07CKpd7QYEtYcHriOc9Ngn68bdSYzm55H3zjRD1v1pmpnmYQ/21/nPKBbAEA/UCnAswYgo/OBcu
lzurEAW/jR5Z1p0agTuQMN00AM1MndgxN3cPqCBBHf9jWMN5YhJBCl7YG7guLv9K+yB+7gy0MHTA
Wo1q/dASyWkPLhmcmMdjnJU+Z2cLjeLpHQPsOjbHn3ebFDxiFLDQkbN/BXf3c6nUGI+vnnfZrdjF
3+gYgrQd6j3tN/Tf5GTNiz/4wnvTty9XIkxmMcedxglEe9Obb45iZLL7c0EzTIfqTWR1tDw+dyoi
6lVUYAXPhJwFO3QJj/ObrfeLNhgQeFmzDZzAFvpd8VKxJYScKRreRLIX3aDCbMqD4ZPIu9Xqg2WR
grVfC66YxGLE3xJw5ihaJHk8JfPBQ5dE/Lpg5dc5Vkb8kUz8sFenBQjDBsAzSpgQlIG812Pvmomq
xlH3xV86tsHO28uPFkCf96w0pG1DYri41BDUJgDjHSkTgpeflhH0FGX40ktwkJqr+D8Yaqwy1KgL
ko4rFXeOP71cPk7ex3QXaHMiuMMykdmjSxZMmip5FOM9Ulmngwc/gR8Z680veyHKGOx77fyb9g5n
CxJCE6NZhcy9Bd4J4vqbtZmoK0IbS3s0Ah1WcciHdtWEtrwosDbSC/RkVXKX2UihKUcNS18xerPL
1mshnjtVjZJ0jPS2ib6oXd7phaY1LFcopBOFoZCWX+5D51TttsowXLHY8fx5eaJy+3ChmNYdCkuM
S8qbjPFR5+BzGeaSRRyQc8bkThQ76VLDbjfrtrZSVj83qwebXrwILi9pPHhvOskevydZUDhJkiEo
BfuerbEaDxiuq/Vvht2Jh8rLM+R9fwfOmetTEbxOz/IY681tJVX5LNI4J3PmJ2H83IdfzmBfgWFK
/83HWudK//HYOeN47c0Ay3EYYL0J7wML/cSnywHNibvl2t3C0YLVf8knGvk2q/hVqkCCZ2yIBDrR
sytPRPrVnm71J26kh+wcgsm0BEV6G/Q+Hzkh5oBxjONoiY4qD7T9hG5UP9IwkAbasjNjXHttst6l
+kTI38uuFau2/wPsnGN6WBYQ38ppS0mwcvaAl+yCkPlTsC/LNXNwYHR7N/FdH4KSd2PbAS57C5Gq
O4pT/5piP/rRQyH7LztxVFffj6PGI4IL4oH+Ag338T9iXaVMqmzKbTHy5bzC0/QnmuMo2NasOa9B
2zSMhoh8ITLZo6UOPTJdjvIrYwYmxpRTgDwiJtLNYVoYtQ/elu8DNZl/+J5ieCfGURf7nPXsmPSD
Z2UzpNxmKo1JG38Qv2ypTle+rFnqxlPt0d7HCjNuxsVDcrgwuWKBjPFPMx+sbmbX5+McvRhXpdaV
e3meskGpWG8PiIP/RxP8KllbFKHtl9Dwb29ptLyhIS9PkXKQ9lheehyyHpmQ2SUve5UTo+SB/5QO
A1rbpF2IJbb69VU0hMJR71ap/LoF3NgUfkrkzj8dn7fwLCmt7MCLknMkQ/hn2YiTDt3wYcuLpLth
K+nTzb5L+C46ti8yISKh2CawiDbrJ/Z437WSI4c7z8rCCuinIy9Jq0yo199rwwQNcj17g0JMHLVr
HgJ/RlczLbUjIUSfC9svbB3IWjhY9HyoFNTIeRf84XJox0/b2WkfeHi+rb4uf2SgMts9P5UTdFzk
AMpE5/HUDqDFCnfohFKKC9X15exNls3XCiNRJ4F2tCE5nIPg9e46e+bqRKof5te09q8nIWJeyClM
I4jHW36zd4pBlXELVk/jakHGRruTMp3X1MBziKnNqchADDO0tCvkE71+o8Rv6zeSXtePAYXY8wL6
/z/NC3kmqNeRtF9ecA1wqZN7fWbjYfT3Mx8K11twDMc0bgWscOVYTLat/xnCnFwY3vJD5b/D3Huc
0MKHQJDQUxXiEPs38bNnBYco+4f/ZLw+pDVrSZy8z4/1mbhuxzxwAJECjYg5xAx0RrOeWJMY5lZX
HI/dc+w0mW9aXJWaP9fTTu5o/1nqsCf8aS5A09H8vTOtbMGFdZZ6Yohiv8LeAKcRYH3f1onmf1DY
7OhUHQPbP6QFkd5R62yw1kH2eXE4LZ0MgixybA17fnGbJflmzSZWVAnOgUOz5Hs6fgV4gxx/t4iA
w3iCt7cBcOLDD1Q8sioMcafI6870I/QMZKVkbwsEQH1wl+YG9v34axg7Wn1LThoBo4LCI8zPvwxx
l8sD8wDbUDdFGdUxZatzFQYtG1cFgVmGJl+hfzBvaSj6CkMHS68VlhvejJCYcAwyFmDctWeMp1Wu
rnYG7K/8KKOFvkMHQBNVpwkzlNmx+TjLpPWYlxGBDuQSU6LHoaHRgbc65Qbl9BT4Kk73IfYn4o80
xO9+AYL035Zhil0jJc7mvyExn89kOjgLcigG8AJJNVt1lUDC0CHnHwgyefK1ToyImZWKE0Ts07Ir
ufrpKxfaSMwjaPU5kCF1u5GAkLKeZ0V3blTeHhESDRVGf19+5ymfPAsglYm0o5LvYl07YYiv/+30
+FzSEyU2Jk6AhLfzytmaV6wWbAI5ywL2iOnpMJ7EDIkejUWRI41ZNNX1rD7H860SVhwpBW6srGbM
fSNQxs6JRkMH9nmCpYuxbGMkiorfCM+etEXDIrIBiGGYmf3YHp2W2W56ZVVtRmju1aDt/3L3NQYg
O6xBeO/V4hpi8TB3FepFcpzy9sOBh+d5i9UoouurR/JyU1xNvMWybMxDShugrD/chYTI3F8Ejucn
9iNo6G/sY2nJi+nHYYLjvPH2nEkGLdA3ozdCdE8vx/bU7V1+C5CygC5ClgS9tgXGc8gxcnJYNISl
fUBjWupnc4mnK34oIP5IQa7rPFLLaKnzTV74V0Fi8CqJpT4S0Mx4gxZmIHRai9OcttniH5VmJert
xo/PCVbQCBeLrY4y6yIng3U4eAZYZmyO5KZLsaWlWu9hk6rAAagNPVq6yVxE691z2kAdGbnqiT5g
YSXe1mRoNVfQ4iNIFGgdazpixuVaRFHTiegyahslwPPEEHIR+hy0ulgCLONTg4EDsw4A0j3rjkRQ
RYGDms8ow+dDZ1q9EQa500cKsyDboJBOnhy6+drT0I2OTwzMhKHPfXN48YXZLkcGnxf87G2eGOZW
bi9qO69GTPu33sxrkQ5iGMxxLma0m7KZ4p1UGBVLPttnehAcEvtLTve/V8zuKqbVt6hOGvGQzfXH
LAZws+l/GbF+UxEBgX2rAaxAnlbdTiwb2MS9+fTrPWKHQblI4VQBDGRmOI4/yrNQcavSdjQt0y6D
u6htqz4BDcFCpRslnHUt34/QR4BnPpAfgdD5mcmaR968KFdx7YRcvU7VPh8e7Yc9ajZITwWp/huE
GE35S8vNnL0vjpNTSdNiQjsRGeWGdsbheF9QeEpW89yafxEL3h+ahoLgkKktdWU5PPGzrTFet1U/
ZjhCpq64t1Oq/I6NgnZt9NTFVZ80DuFfLFI/MMyOElDFCeijjCPJW9rjU0R+u20COoOXu1Cp4MBA
WRBDYy30ugfNgfiLpGt1jQOM4YhjFssNQCGzcZNSJo65NkUeToQKVfCPMFrP5+LcooEJLCpEdMV8
4Lg1jyFtFbeuhNlTs5PL/DhQ02UIuCt4UNfQCZNAMT0nKMkJv2bxS2CsO9uXatKNZ5PmiFMob44+
5r8QeBxFaKiytDoJbn0OSbbbNeiL90cw4KYCYufxTL+UTveJfcX7mJrUIV5zlMaTqjrC4N3TTuVU
9/oX2+5NxD0aD55WNw0a4mm1uazsuu2IgPzlMk8YpQ7GjRb4ECFiGJ9kOGM0O4Sj6bkl2pLSI6k0
dONfVQh+jdqrDSoDLwmFDUV7sG7b8a8p5fpe58hdGaOQX2GE1jQX5quNUhBrqPchiIwL3RPL4k9T
pKdaTjt2Wg6D4X9rk1xZ3xqVAGrlYvCZTM051nOTRism4nI5QIawF0h1nveFcnv+aoTSZTWpSaej
9x30kct30hFgEWAKAG/7pb9yMT9bexG2e4qDc7AXL9Rv1VI97Zwfv7ZdQBwvdb4YUscY9v/zR4dK
gWY2Ww6KEefRs41kGmcGIpx+PGv0BazKVERMor7NOB0Vw0fQh+RN1TVPl65tHUA1UFtAxfkdn6Ug
/nzJWyfDc8TMPBQGskQVfxGMZ5Qstn4Xz+38jDSi2ex88Pvkf1mb0056H+MV0/3KsZBqVOS/De+y
fQ1tvQ6TzRTwRGMOWSjNPC2bsWQ8498B9Lv2HhCve89X3CxI59ZQdi1iAEBjqgZAu4F0oQQ6phwN
pyTuuqhSv54TvNLVxRt9Zzmc/JaEkL+UkzmQ69N+hlsulcSCM7xi85CenMWazyRoC+vVwXyMAjWn
YhR6eayp/XZSYxfc2bBNLK009oqfslxrktzu4HAgvvWvkbwHBsTTSMiNvdafimL/3Y3B0ClKRlil
locVUQWfs0e5XzM4s5Fvimqgk3dBs2UiDNkzkXUmaSToYiqHg+mBn1PrezhKJXwLeZQ/HnTzv0rk
EnmLRbMs0q/OuvAJhJsHLR8RlSUpJcP/7OFAf3KgGawoCfRW085jRMKAU+JmP8dmsmhvBUjwg2X6
hoYpsDME6hSmviAteZXOKB69yivDQOC3/+SXvwYby86YvA7WpS3gho/mR1hcjnaMtiN/Ft3ssXda
52e32rKnjhTAL4ngTOtMVcRtwuO63QvGe3NHCgRMvDFPjSN0NKWU/m3/zvKrB/wlJ+Fnn3K5pLd6
21THe3uhWigCTu/i0Yxvi4kCPtl18cyuDol6UPsR4vH32z9Z5l4fV/UbgNUnQfvP6Yu9LJZYCQKf
2NntlPhgJV/pbWPInj0tugDZjlsRHtfF70RLEj2ucQWsrzRdYWvhkQE/6uCMxCNt/rbXRJBtYjmR
f/I7PdwsdtuP6E0R78Dxa0YjVFmhNYsHoY710QkvtNxlEjgC0PeHD4p4w9dN3ljb2INR7KoHatkj
fejS5PnLTnbNN9WSNnhRoumb0WenS+bHqkeMEx+UBDnl5ra6eBF3WYQXpDncAG4FegEfBNnCnkwd
ppjQlkB2Z5xB6SQlCp+8nyTNGTAWBjLfSYCeMXn6y9FbXvUNbovVzw3T6MlS5YFCUR+DVxtFZrKT
mRT48RwxekRFoNU5sI05WIZP8Zwi1LerJFFzXIXdFkMDtlTQZLJ7kgXi9+t5fFBUzR8o0S1HU1Ne
aQR1Gu6Kt81MKAvBqHOxWEAxfm3KIyLZ+s1MknekjS7LYwh8gxA19JUYSlk3Lm8vdhyXHUbZQxK5
SfvZJ3NdDs1ZxVBc1X9NxUYt5TF8ltHsLHqVHIJyPm0a//EBIdkApkwhD/8UrZa9CZ67jtjH83/W
MDv+06bhyk3TPnV9qrCUUBxKRQGBNFFEA/Dnsl1ad2jtyCqCAKyOKupqGCGqnQ/6nbUhFF8Xq7yF
EscqSFaxPpBWBCXOSvSL7TktAw+lTsEEHvX2stjlQonNN1DKJZRKyz7MMQ1N3nOvTn2X8U/3MPdv
yF0CuC9OfYJN797D9PoCY82gEq4HguD5NQwgy+7ZOIjbdH4qrH7J58lZ1r5428paRgdkQ5TrTC4f
SWvlhMVoehBtxcGo2eLvJ1gP4IW+8g3U/beEJHJkV+h+Whs3D0XnQN9lS06KQm4OK6UPzrO4+MV5
PAw3gdGMZjA2j7JTtx15/iWNDu6fPVN3looelFp1OkKnuyQh9hvTJQiZ8f3991a9MMtAEurvoRTp
qD+AQMLe7SsE1UEGfKJ+p6C9K1NqHo0nqnhYighSFjbHJdZHgK6F830DrfsZ6f09pV2Vcg2St2ys
hf+YsfOb1yuydCMGV1LEywg+yeJbS5LixAOCn4SrakJgCH1/XHEkJTojw/4AOCeZ3XIvsOWYDd8X
tIbkPDFt+fHXbNcjoVK1VwgRx0PVznNYrokt4FjrNpxfeVtnjNRlQlaXdCgcWE6imztx4Y++TNZV
/OGGmDLvo1cCQoTEgwZepjyFkaqcnHHT1adIua8r4JTRaCrh37ezgi1tRhbEqnaO7usGUXyaILZr
WKx5gDlx7cQPmIcMe5H/koV9t5S/O5JvQux3J4UoKu47T1SmcIyWZBK2ci8Phlr5tdEa0DwfuZBa
ik2CN9pCC/3UZp5Tk8QvBH4nuMiNUd02XNg0nuoXrCN/rPmNPuF64ANK+doRpAjLBf+dAkV9z5tu
4vMhUUQ2U88YSL1Yal2Bifh0kA6IdRptCjAh6BS/Fvod6W8+9NNJfr6+H6pqcG0t3K3Xw2kxyPR9
RUkFbVuUFVHhv/o+pfEXXoecgcvjx40mBqnSWpVqrMqMCs6LdSt4t7iXJDhqxFYxeay7GpqkyTCK
C+4W3PXlTMkJvlR9d70WBaQNEbuzBMSxClyNcE/YtCOESAZDBqeGcRbzqkuiuPDj5yu+wWc10Isp
ZVnovENQRwnYC/dAJlfrNm9RXhbr2f4XwRmwLwy6jIVmaHX/rwMwa13GG89q8fDdG4xxl6HtWnN3
45rx0ZqYkQ6qrPX089r5BNEb4XXehOCzNZKHeAE8mITXwPs8GUmFF5WqadRoGxXufs93oqkTyfgB
wRxwHSr3ett6U27DHKiTqLIn4VbTJvM+GOb0zXHGt/nZxi0gkLPy9kxCGXuDIwrG4ChPArkRyw/4
hG+k3kQF3pbJkCtDvHZL28wXb4I1L64gGeN4JZeC3+LLB57CnxcNUnTd1nRCmfoJOEpSIxmH50OA
u2DrneD1i1OnrVWecofc74Q9RMxqL75wO7Fld8q5Ay1eOTZRdgThOvPHQDwWNAmwyNwQS1aZZvbk
mU0605zO9QUauSTIxPQvJl8/m/1I8WllpH6tgBntVQOpNprwS4v+nrG/1uXBe48/ahhe9JXKofP7
I5I0Lo54We+3ZG3OtSOJbRvQmmUDmQ8sgHvDl5upYGCBRZ77Lcj425ezrFEn+0KQKrttnDeduuv3
d9Uyy9FVgMKn6YL8FVTn+lx0VUSn9yWklcSpC2Saai8ak00OOZnR+vV5CCCgegaEeT/4ldESxz3n
dOWGSxP34Xz2gDT1UYdzb+m1VU7NpjzUmesmFuybuVmpZYlbEPpPRpEIqTW1QpYFinZ350G+0W+N
BZJezpNXcZ8ib2QvBM9nBwx1D1Z3GYQ4OzV1tPIF/oPii7NXA0ysM1I3HYeWqajTdAAE/6/eUQT7
MIcDcBKzhPwTP/AAGwNGgeFy+8zcklKI6VwbXvMe6mwB/7agW5gGwakmq0uww/3nXA9m/mwH33Le
pMeV+C6pKhLKXcnNfnwWViskrPIwm1kUdQe2T3YPG64e1UbPotr9oUko4S4JI+Tu1dcXkvYFKTSV
BBlUd/pDdoeoLOjgZkdoyzLnuQnZ8Q7Irf8DI8gCSo7XSBP3AX6o/MdMqSQVeZZ9zCHjaGkm6qav
MhYoeH5SwX7wmlatnFe45s4fsegAwNjsaOJofRumuNnJl8q/F4/BtdawMie4z/W3DA8tgOLJS6A6
+nUZqRdNgqf575FdD4w7ZqJWQ+b43RvIZG6hngJUcouNyKpS/4VDMC6bc5oaCttDLL+Mc+Sa6HOi
w90/Lw5xyBRSulsAzUJ/6q5z0m5R9jm4WVj1AiZscCFK2TMBFU3sM3I5bJNIbtgtxRV7EfIdtkta
UGFH95MlBQmdKqihoCP7XM6KgTSOuQTUl2v+6nW4AhTCkPixlUWH5Gj1eFosMnJc94U553JFhCrr
v6EVJUw5PxSpUM1Jc+8PdIDXjsRNKHJrVqDROPVmwnbeuGTG83HaQIBfa3YIv1rP/bVTbzjWnVM+
Qc3foAuk1/Ejz6QQ3HeAAg8duWgeXfaxGQUrZH/alXCBy6RQRV3Tw28bF3YS6ixV9hfbQEPMtCO/
S2GQ5vfiO49uHTYBg3gKAcyS4NB534coCvSsGO0/ZFKJ96iehE9TV8bROhW4fmTUJzYL10soYfco
GHtATJcFXMVYpL468SdKFrw1UN7yldFUdM2Cmh5K/+FXrwT5Na17FWe0U6dZHcEgIo6O7CGizn4N
hdzHykRzPf9HSUxIwAlZTfYqI8UhrDVmGx9UN9UbylEk5KKZL0EVCPffYjtMvlpAYbZ7TBsyHOVb
pLy5Mqq8iA509fQFtm6t7s9jHXS/HxYFqm4YfcJDi//cUlGm+37c38xQXP8mRFU0tivLRWAcD5UL
VfZVntDnolKO57JwjQ8xTf/7X7Z9N4MvfZiy85rmBRrldZnhXgBUWqH39R52tjqwS+RQ3gklcM6P
uA0G39DGVZavjKfo0iNOziMDbGp75Tt6U2oX8I/Rmy+Ao7vfz76XwXYSeQBTYmVGvTxh4vLVc2gW
02ns2X18OB9Kzo0/a/TQZ/z1MZdgBU5idDp39JKPZ/+qjf95rN4zueS1xh50XcuLDmY4dn55quej
XIZ6AUoJGC+m+M+FAiwXxMCvusnSLufU8xAZ9vwadxZtUwo+3AgEGdTtUpTa9TVt6B0O/QoE7f0V
fB9i/8OOaBiuTbx3Ffl/yC0p2qr0Rtg2VpLYKw6M7Ah+bdE60TVO+17jLSX8KPQmXg/K3U3vy7rN
XXP7mf5Ub0Y0zIi990JOFadOVac1umqKs6ArEQGKzYbtAS8i4mZpqS3HRTFpfuNpFX/5zjID/0GX
w887FZ0SXvsdFaY3Yp2ctnhrPcttRILVyV955p/hyhh8fZDS+G5ZFPR/Hpkb3VM1DrcVzQtJbnxn
XGuHHVicmBCPb8ukumjRxl7Zk/GKV4PFCpTDsIXlvdUo3lLjljaN2dUOy+P8r8LspYiFSgLgfhyq
5icUr35lNBps6m2aEp+FuGJaXHCutAGq6xNhB/BSPvwKURbf8pyhn1AbWaLZRiRxDTG/ej9Y032a
SEgBelJeVOV7pNVn0gqJO0vEFKvIa7PVELNb5AO6HrPrh1j82+8fvUtRYLU/3KNfcca9QnN4BP+X
z7i1aA6f0ShMgccDZo6px0SR4OnuuHc/YmxwLurDLKzhs0wbl8q650QsgC26nHKt+itig3m/KHaM
zBVct/W1TreX/LL6TjW93aW1sMo5I9h1sO96csSH5VoqLX7A8+UDDxi4xVIwbp6jlCcT6wSitwty
1RInxGHKzNqtmPjByv2/x+1eAGOI2DTp9KNV2Io+wAjXHxVaUAX0aL85tTCDMHAdR37rgkKsfWiY
aFoTEP22Lx7NuhWZrE4ZF/Du+Mz6tmmYwR9EUfbJ9VbDWG1gsOnjl4DDlHADQ6v6i0Y/40UHwGa2
57kT8Magal/wYyVuofkys4skHbK+/XJrlw+JYOP7f97KmbZ8PwHJFibV9geDdxeEiLXFZi9DWGVG
cvOrky2PCTNRfVjd2Yfx+8GmHlRtw3vfdMPH6fV9cQ4QNuXKYqshetfBxPXTM7fS0CBpAGSBdej0
GCdr5Y0E48tvI7iXSS7ozwV3WvWdSgsN61X0iGrEssG8tnYwxkl8ECmuSxW7bwueL03LMZkCSeLe
aYbhyuUZZDep2XVQnT+GgNoAg1U3oVqq9F9TsO9ieU/E2N6YN5fYb+xtKNZRhmr8xMmF/pkccqS6
CMXF4zF5FoeAJYt/7uQcAzwqBsFKZTCT7+BYx7BtMmychIWmFHPGIx2lEJib+oWgsq4zTaEg/8Gj
0xB7cu2LThHBA61v1ZzlqKiFqLD+PVVRpmvLIes3OGdfrDTxOmQb7zKKB0zMGnAIenk4GX0G1JOH
FG2J/hpCfLAwFT+T6YKzdyhL/DXGSW0BJSVDYp0N1Du/VhgDsSWXItuL0KmvZxKF17z8DywF/43T
rf7Dccn28BTL8erBLzNvkU0uucIVg85n0h0HeCK/Q8+z8TOMNJWHCePFjd1N0Li4R5/o9JTM90zo
KgrcRKLp5nAntwLhJzfHCfwGhtTXnsbADid64Ax3O316drAh8RcdTx4SQcz+mXm4IMU9xYKCBins
hAO+lGgx1sp57poJn6ThAIqt8h+zQ25ca9YM8iZ3IG2RX8IVp508xWP+lZx8uTalk1dZVs0ok16J
c/g6q4gD5pWjYwLZx7RTBFSuqos7krientVbNcrOT7JfgauJiP17VetXgi3emqVF1vrDTnu1TAUS
ysU+NG7rgRXiSugJQKQuHoDt4OLIsgUporfE/foPR4K+s8syOIpw6ntOxCBZm5kyht3nUb6m9oia
OzIJOL9qEUK1WjpEbjLIWVfOS9fwkUHgKuCXWOreMKwuT6o5lFHcm5qXn04bJ2o3ovcF2StjHNXg
Rn+5nJuTDPdt0mPMzwkKT2ep6q2JwUvXd2IcDTgRgqU20ScMcHTJl/oEB1wfFG6DX3fG/vct5Wj+
Cn6LNLCVFkeZ1k64KMSfWpV4MfwsDpgCACXFAtBIlesDaIAeLIqHCngoceICpstveakqQSJJGvOa
vM3qsEyF1wPzlwmX6tJniYiTnMsQ79cZdKt0BTKHQj9z/zJIeODJalND0oLbc/J+tc99lokHpapX
Nw45e/E7JF1CXTJgpmzOlCDVBbn32LW3REgTSJJ8ECsS/Vkz/QPsl44zUUUB+JpYuV1zydU+1Mj3
+ntRd+by+mMD7I8biJOz83AVkpD2bXTtKoRaHgSRvhTXHn68Yulw8yxmBpEk59JnvJ2yBDjPTgA4
eHbTiPUhiZ7oHAPO/b96fRUvoylGW/K6saeKVg1CC/T9oI2n7G5CUVqwC4JDyg2J6ahJpaSebHiA
W4QrBiDENvX+TGaVzBbeMadTgViVqYXQDl/DBC1YzQ81Ymk2cp6Tf7od73LMEvCffsmYErqfTmdy
R8OCS6I7cjuYjg3eSzEkVqouy9OWH16RswJocmhy5/8JBJ7dIaYHqF9gTTIj2XXoCLwBsKQW1UfK
FlOeY22Y/aw0vbSDreHstKlDrBDTHELzujCJY0OMOvRhY6mMMB2dLIPnlJjVhhnC3huaVnkYA20d
8D2GuwhJpOzg49eOA2vWtpwdwMCD/XmnhpLgjbJq64ILdb63tbffRbfOiqNpT5PnOpgaC4xQT4bR
uTxKQWipsbixtkDG9c+DHNkwMZTVx8oyA9eMXDceOpHSEOv+5jHE2Z5fl27orMXrvelVK6dmZvB8
ZPHLhwW8TuigAkOO9q5Lm5/MkEFN9sEzTv+f6/y5yLBSnOHe/WhB86fSSr0GFMqbD4rlYwaPaqC7
u7fkSWstFdgr326NvgPLVdRm5TBVmmarPx/XYSC6YzQjqv14U4xA4Z7dfxIg1IaTQ3iiDYKMuY8S
81jlwz+V2iThzbgP9YQGqrH8rmMsbUQbQZfLGV2p39lnkb8PEYHeizO75186FYRTcynuPRG+MEeI
gfzrTiB/p0nfLw7SPjez+Wzc+KOKNUXVO9Jzoh1ahMQRV0JYgaXuIRCMElU9sgGUlT/8qPFdGqSF
XMzizFigzzzOlA8aXKS+xEQD7yTWP3cXxaz+KiuU8FgyGu0wAw4ZeHlL0kksiiBCI2AKgh4v6cN1
aLui34ixjbwMWLJupeMDP/H/uCBpPcuNnpmN6LvF27N6rI8lLd3Oraq+3sYfQH2MaIvQWmo0QMUm
3edbm1nxaQImiztZqnxkasdYGl42MP6Bvyu6+A85WmK8RlDHEBV7s7iTdNgYJoeTol3NMpmY24hQ
44ld93LN33KQ7yBNgNY/SX1ocF70hYVKkzSTBiZo6a0k5KJUuG4LGaJxsSkdp7t3+7DnzG9UDWq+
oWwiJB7M321FonVsGjn/bAP/uJLX4uZD0S7F4uKcfyl6YbY2xQgkJnUBTiSvscZUYmyOnZo7V+wm
txZb4iErrcfak0V6XUa8kypncSbkZ+pZpUBwIKSGM7484z0WP8lVp09xzrXAa0QXYxN3X+Gb32i+
7//7keruaPOs9V6i9FTakOHejMajCis4jtfC/bbBnkRlM5VMNi4yoNo6uldKwSPlgW7tgmzu9Db7
0LWs515KLzX31ICjcSlukX4zbiKw7XdiAQbWkgfKKlgGKYED0jxfVV6F10/ZExzuIwQGqQYp/2K4
x7JQDyFwUQtt4ojwRbyd5Nc7ghGS7FipDnytU2D0rScAG0tcaynunmkuhvMbyyJygdW9pYNwE4gC
FinU3j1FfvFUvjDOzSwBQKC/ibhuGqBpj0J5w62Mnu++NxZcecni5xZORtPMppBRl7kT8wit88SY
Oo5yV0E0C0PMM9Wv46r/omVZIaftaJ74lEdtPWULiln0ZdM1DMTCC41ivKVfiBeiLBllrjMvCnq1
jl+BUo/4rssHZlG7P2o8ip2fmFhZ8w6tcouQVIt/DpXjPibm2A/bL7b0W/56fVnyrcx+ibemHd5v
dWBcYNa8+psKhc+JZLz379ZgTUaS3+t4gGRdzA3NPCs1Q0M2GH/+4nag+8FwwdyqeFqDBvO/2Emf
nqwnTUf5Go4n3s4EO0JG3qxyT2UBaBM4kouzx9oVA/yhErdswHwrB08hajAJ9SgmBGV2+M9PvEmt
p+z7e4KbB6cddWeoBnz9uyyef5Ozbn98CYH/DQb1nT5jRq3nNZtbyjgWKsKEXfjjwj7As2EPA6Zk
b8FKYlUSAzhtYqoeoJTEBWyTQ+Y5mUZedQDMy72tao+mvt4q7DQltdAdpkJ8SN3TEbuM/lrbeQXR
NhzuLw0OsELjJOCWcpFAHA1V1FPXctFHxFwCV0zecrNXrl4IUgHuM8yNodx+ZjIRS27z9Du1R+OC
Bbzfg7dJj3Nde9MjY6DW6tS+4wnoaBjjxMcqFuiwvWFBbZiBUJACWIMYYDqVAnDhqFmyTzrkvRk+
QrwiMQf/4jEOYdh5uxmA3hnKIhCVhVg+mVF5+bKttHYOLmf9PmNDA4EK92TxkRKt5nZ+2abRaWI+
QA62ikDReqEsVLazWDC1UKVqgXb6yOEz4g5rdYNMaLKpdjacG4Q3DtcSfDTLLlcAAA+tc/2tuxEs
WyWc88HlDNrznR+ustD4rJCVT7mSWuzqHQmxRdunTgciJZCQDZ+tiv6Ym7Iw9Jh3BitaIjAGAM7Y
yT7NFupyfJg6ovkNO6SLykn4weFneI/cjdzFETJy6mmaGrAsr8Cdy5Hjt+VYPfm7bOog4GX0bdI2
8gLx8tHNUxJLGLBk29Ilw8VjQseqhIayO/9KUfP1DMweRvT8c6TqZ+EI9iEoSHIk1sJk1GyDyV29
6nsk6GQ7PX+cA/fXRF8IJgwWzgxiSt4WfLyj141vMU/i4RvZa0x5SNj9TDkQBsKUrtsmO+XOk1WI
SnTCwLT5MXMjMq/nAbZQ1oPIPMhr/0M9M9wX0wbn+vALs+ZsI6wyfAohO4WGVaL1cEQWGpZaHe4o
v0w2nsyWAp89oQEZzG1Ob5wtWVE8qda0i6UFOfFgfGu2NkvQSgdJ6anpMxNYYzr6Smo60RrQm0O7
ULg+z36M51wVIgxdUOvWjeD75Z+UDRBbOPPVmDOTLn/ccMgO2vl801mGT7ZLwX/FSTUGivTtemx2
SGd/7UB9z154yjgHIBWPn39YeUokav/5MfrwFcaQLss/SxUS99XZ8Z20qTquSEZ3AjRy/DraEJr6
Nr+evGsZT3qReGWoXycS+rsEh5aywl/cBCxDcRZKLUesABHuZPjOKr9Rr49wTkohmqJTdFZf64lA
cXqB4+pFmseCHBQqRQPKKsJDs0uyWleL2AoytGemDMSypSQk7O1eecM9xBUbW/ZjZtZmaBpBwYAd
DAwRBnfUD+Oqq3XY8kMaSpiHf8BmvS80DDkhUOwnNnSCRMbtxmwC38CW3fogWLQ1lZ2t+idmeIGo
4TIOnPjr8EPV8izyzee42TywOpYKtP9jgeZE5v1UR/KVkLUoWdLTORfUlxO1/HftfdkesQyj+ovb
cj+TQhEv3Q8X8dnVua0BUOhHZSsjj9mV0jBSmY5MEjNrXtDaJMbxv3AYw5gcL6bwyQJrn4Rky735
Xmjqb8j66hDX1qVDjPRaIzG1cVzIfFrjmTAtE9r/kAX84wvJqayp9Z4c6yS1U8VOVUv+H5owi1WI
3MyLfR+MebOA8hx3eZEWULVwmkGcUaeqdVOCtO0D+v+4We8X2QVaml/HCGPvig/oIDHxDj4fO8iN
iQTM06THGTrr5JzsjQW0Hf/OAAidhxAc+vVXEEcnfIv2X4efMCsoGeQG2hPGlpPC37E0yRq6r7+O
jEZyWXz//PYoPw35vmP9GoHGkJfRcCYyJTYmfa42o8PdwB9IfSI2vzkcH7GR/FgPo823FjkcfNRI
levmS/Vd553fZZVsyGD8lFFklJFnFe9UO1j4bE/cf/T/rFycBHIZoLlNu172ecHd74fZSOm3AYrq
clk9E8dprVkpk4QNsFgGAqNswMyZA76WwengNmz1aUMJbyfp5BOJs5TRJwTyU/IeCfTnuC4YiR/E
DeyhcDkRw5aGjfNnTc/cIdgAzbKvMU6RydyD1/+WaG0DMXpzCp5rkROtzFMHRPl+t0MSqvtyBpH9
BragyTr9WKupBEiNiujwayC44lBADyJrmq2sa9iPQGtkJ0hZWB1Oqi236GzW7tY+oQ60PYQyn0+f
G5jjayruSSPqBIf8mcjtHHQaqnTE4unpj6En4D6ysFthDHWAVsuTyfE2FOSraE3VA1fnqlyCixYK
k9OI/GhrY3IRCHfISysPt7n0j7DvD34T8yjt1Kxc3tO2vHXnSEtfFyuqtRE1Wsbsp/LfdCMvP9hV
3J2diSPyW6QpYE5AbZtLgKc4a12yUtOfV41AyNArXacb7fJMeThHAMYojjfMElvn/zzD/8TYsAkx
aPptTVjDSKQeYo9wtLR6KLRAgi29B8y3bCC1UVcBVGO4p9yG4b2j/J9AZfLGI21w9RuVU/UbTfDu
p7ixQWY14h2HOxVqqvZQ9TwhbNQfk6gyflmDcchCmMlgSlrMZU3wTOl/rmo8YvLQSfsXHIpURkh0
O5mFWn8x+G3Fb/9sNgFV0278eVa7ImcCc+FzdsTzcxRH1A3JGwtxitUbJU04IFeMo9y2A20xTo9o
mkIQguIdOsEGuRd8P1Ih7iAVj7+x5YtY6d7LLm10FpbAq66cG+0/qkZmS+bU5SzPpiyfkYiKZFSk
BlSl7OyJhX7cTmtEaOgjtuJQE/bNB9yk8OIH1TNHr2VLhmJMbre4UAovTjpPNO/FT5GnhXZ5Ag84
Fh0otJZz5V5C81lwAQLM07smllfsTfWkZ00+ib6bo7NYcpon/XnR39K8k4lLoFja+veXzg3tfuL8
KPhrn6m0Cmp3BAqjUb2kd9OrUcbL4TEgjMP3xm6ySf3000NF0gQCwDrb53NVkh2E84n3xsVclNdB
9RDxUkWrwGuZMLN8QyZA0kwS5xE9ABiVN9tm3Q6a/j2Wrj8OOIAlvtoSADJXVbuM/EPdBEViz+H/
ihfC+q/oaSjj9bzKZN2aLcWZj3PbwArNYPduNAW3WKHcxs1/UaADAyP5rfdd/DP4EzHrP517ZsHB
ajkKw3r3ASBAD5EkbD5D93k1I/23IPhccuyHdfc2EbYJlcXM4zw06qUM+xQauXh1WwRvYSGRoUx8
+Q0Qqtx81XJBMfNWaNQKoJ28fR7kvyvrWlGpJ+slU230lsKesVyqJbpyDYEzDDAqzqJEDSzkWDA3
yFUbUZmfaRwX1PVkzvsPlmVyl04uojIhPtkpsYXhswHWeT11F4PZ0JGAZ7f4MIP4giF9s2b7HRfJ
e0NRUhbsDMcvMI61NTBEma6akYkBBiJ49emsJvDoFaPKi3OS/lJsgJjWn/c+tZtsdbY9nTx6D97o
WTetG4kpI6Tmgr785renO+Y8vk5cymVLz1RgqfseAbh4vAHmXMF+MCZwYkGEs9EBSxc6KzTouHuG
yTdqWTTWGz68PMFHmTXKluNl1vh9anThirHyGGT3e8eqOibeC8bGliUF+je8Uy0Qd2l3zQuOka6n
g4zujTfI5nQ80Vag16OygbLrUm/W6i5dshnUm6nC5mZRoh/cPxHyYe/dtNfP3sa9YPYBUDKs0386
UIzen4ndT1RpVH5bzPzSr18IrqkrzdnAzP6Yluj4qDFlA3CwdENiBRQelrvWQx0/w8GEdo7ijN8w
qp4EA86Bucpddrsu9DEdieNULWtY8CN4hr/gtxNpqYlcSAb4tIk+r0C99qqU+cMUzjCVQg/OE1b2
zOEonb/LvyT7CzJYJyQIX1mfBz9G7cOmNP2V0KYU2lslMHuTqYbvBiZP+T1e5MUy4iUrLc1rEIvq
ztuSD3rLheaiB7C0+oESROOJDX9r/TceHN6wuWe5G4Oid+uHroSh4HJfcd+hrz/bXyYlqa2Ake41
eClIN+oeO2BfI6EPBqTbuy+U43p9oTzSKX8KrXPSpdNryw0Wy1E4DlGi65sUGCQMA+RrncLoL4PK
XxkRagvyplqAb5N/P6aBgNMPzPHz3fBxjqRd/6VQwmHa+GROPis1zT1hZSVU4mm+bmsG4+0vsomx
VfhYNpQ+ootgZfV7feXO9Ise+NkGj8kq2itAH6zuVmqTjadyMS64+8jxPaz3spg/F46j/kVjNWWq
X3ReqIeBxWRTRSdF7By6KkeKrhSsrQgq8+BXzWVrGE+SLsb2Fj68k+l2LkkA/8tqE21LOOXe9OKS
CzFZT5f+5hWQvjbozPg+crzubDuCC7VrexK92Eqn7Wa2zfReiMOByAzh1ZpanI/jUX5QDdEdKu7u
vaNOTtWGvWWvuxG2cLIbN2y562F0WeajRH6xEbo4JK/SEx4/IidqiSN0AWFYb72NZuZ2Od3i+5ms
ZXLZbopzyMYKRgjXIApV3PwVnuQZsxPHNJ0Mwsrhfv0Kl0pvd2yqK5DT94UmQribvRgPh6nuLVIr
VgnJ2aVe9vf2oiZBDSExWTn9qtW5xfxEEa3Q/6gjkn8K85drUZs+OH63NzSBdBYmjFaf2oeYx6fV
UCKB17KF23AxXO075nV30ETtG1g7VsbUJw94setexJ6Y9oS/k2FxdjB2HpCaPqBuqr4EpATinXb9
t2Y/cEInJM1PYmFwW1b5AA1GOYcvmKEaKv/IUZFpYiQaevQMcUgQndsvlEoDlzRN0jfsvA3Ra7Ia
OVLRZ2zVPBATsvekmliajTfoXOzoP7N3xpnK6Fqq1dYFQiW7t7Gpl19d9ltf9RHzuvKCpTlAskrY
x8QmPuA5GpDvUwRQuLvqcMCqLKsmL0rgwvn83WLimbm86QwvSEx9D99r+CD8RyS6rKwEg6AMKLf2
FYQgmRqZT1ZEPZAINTiPGJ8C9FAqBqgCiPONg4QG+nDu6lE95t/Ci5V2LFDQp/+n0KLZRSzs4Taa
fQfPPqxRmjmu9xmOGxIOlcHb8rb57SkLMBKTlCsy/+2yC/lrc8yDe9EPsXEsVDAI+xm2iz0LbLQO
8GOWTa5CVgSq6HxrvOTusc8PMpT4lv9hFL7NYnh7LkS6vL0onwDN1exBBOQQDzp2tBVxVknUtt5J
JfVrIIC1/13q8ccGS/3LtL0f0CyAIzmudW5/uTY+xP5jSpKElMjLGpCUbakpLpM3BLhNEgkx03Iw
F0YMIcM1ht1Pq2e1iJSdXlxMB53IYn08cPZ24VDUuNFUf3pkU6XEb5XEnou4U34nJv33KQ86C5Hn
WiXl7lMnWkMzHV0iL6jsemCBpK1gFfTD65GP0+QEaaS+sWolhC/3Vs3OtOoYMtv32JNVw28Rw2mC
pQjvA9LD7J8TSMDrG3Mz02jtb3RoxpBO+wPPtpJF+88y9iyWsH6qro9vOjN48lkd3kzoZC3/p9nx
zLErJ4NZqpWvjojWuHT/NOS4fTRIGtxA0JwyhRgKmpWSGpAIbytuo3Vvocvfslv/iZMOeUEX9fH6
yqixXD0sFJkYfO2z4qt7GsRHoGcUKP6u6bS0PzdATWVnCUbR2pqUGW6jRSj8lO3v4/6fWP07NACT
CRuaO5y6po4m5Fd949vj2J52LL76pv775Q/Xyy7IQP08Tx2AmSTIJu/9tu/wanA+Bu7zBrc9LXaX
mHaaCfq0pWKv+C8G21PB1HPcVRf3apSN2HtE5vbfI5hZlg1mW40rO86R4SeNBs4F6xvhhuWuXHhh
xbo94fdnOsbYpgGO0a8tyon88lYlV8RzOkxK/lc9uzMMQVZCJ1MOt2CJTmeZil9SFdINwW4E84wm
ULuTTxJkHkW72zyElFFpwcT3NtL6DfeYgsz/LBaPtO2joczIEfxpLlKBnzxp0kKzLcbOtHObt5B8
coGEvPW7WzSleC/LSAwjLqeOrEIeyuGxrN+QqLW+OuUA816EYAId0D5jlt1PoaRGkiScyV6nX34z
lZf06qOR0vQDWh2zKuMebfQLWHGWi62KwMB2D+ESmrMOm37oDR6FvxD6waFQhenXrwwRzggFn0up
8CHOfskumVQ103/Yf5SJPPX0spKB4IXfS0xI9XVkfJUCDnkmaVvM66T3yvtl6qRT09Gs1EJZU1rK
luEGHrPWHPXsuGNp1S7ILCC3q+2Z2twf59ergKdRSDuu6FIsyOh3bFQmIAdZBfeYX/+Wthpo4JUZ
1lPQ2MY2jRly6C9BpStGK2WJQagg9XSBKiH3f1TZVEcSWnXIQrc9y8GC2DH7ly2nq4LXqC5GvIgX
tWsUtvk1BszyeHOm/E3TQOxTkr92yGB5v8blGjRjaNVqYVIInkvj1bahdIUHipOVGIrAVX0mgeEw
JzfC5YSKk8bECVfFxIHTb06cAM2EEmYpik82kmSpE4gYrWbQxMeAus5AQF7nMtV5+jW1J9Zw0Trh
IOtZY6+8kdeLbTd3x9LR67bDDSo7DPN9mXbkyYbidP1gmxkJRs5L9z7EnqQyPc0evPTEf8wnygxp
EmfUe+xopuvGqK6xmmcm996g3Lo6eF+/NlpRF36ejdTJA3OxIOXXatsTVjrfo4RdAsJO3iYCDjJv
jzPRI49Thzo9ZzLjCNK+/Bj0xmcEFEUOTDetjykhMCfAaHui/cUNENZT4/B6PWAzB4I9I7AgJc3M
M9qb4u+bocb9v45qib9jSUGILDabuJsHuuNjf346cUOXPmf6d1y7BFVHpPz3a7ixe+Mi7/fHpyCg
w32aNHi5Bnf4UpviFCgFYWF4RFZj2iIV3JdTLMKTh6lvbAS99swE1u2WPQeKVQvZPXCwDybDHe0i
E11Udu2YPpQa221h5IW9jid5R+7w6vW+vsLM84CvFIEreQFOCTZebPrLL3aPRTTfHNB3v7zO0b4A
WdhOUBjOns6FSXMssBpxvZE+aoWTC3OPhdX84FtLRMSJWrcSx+6Mfq4h8ed5x6VrGdVa+9qtNFWo
QVMq8XDk0rqFrHDXZkOx2o6MWWDRuMnJBnNvc21PS7cR4p+D6sBJNZ6d+cgfu56Sa8sVDvAoZK6O
i8tzSwkD3scITjv2OYKyhOnEToTs/uEM7rn/cq99bD7jqRxk0SvFJaqryMpq6DDIH+ZHPx0OFpWJ
p4wfVeyfBte1RRUY4vtEFgDh5tjGkUhuCMN3k0JMTBn+bb3QZiP3ZVxBN2cFuXGFaS2nI8tqQyXe
Ss+Y9srnkzs7WAio3qvSHzOjHLMIBsOnBbdx0c4TNdEnDD1HAAFjtrqPNfeMe/lijHliPib0hP9k
wDkJOZaUgs3P/Gn4MHaaC/6vqLFJ3+0RumA0Tyx/xJu4q/j584+qUmCwccBnZEFUah8NvJmXxTaW
MSNXj9Ik8rSGpQxCkD+8ojOJak7xbatzjxZAISGW1Wv5F/sr4QZ91jrag+SGSdr0eks+CBI6twFC
C5B5aoEfHFJ2AuRSORQG21OpQwPLmhxtE+CY2FKcdvmPgmKCbQAcG/oEBHuPvVEu5mni3iV+bvqe
h2sWDt193cNmxdVIMNKrWpghafddNnPkxjvqqkLIAj7pOefG3ddivkFRFUQezKV3NjIZlIO6h5LJ
MjBTo2LvJSwWjmhJXo9pCtuKgDjAJTLjW+tekGt1vjXAVLOnfq9jLZlfokAIT7Vxc2LPMaKWbGPv
zCzczrT7JBf/YHhkzfEUe/Ry2oI+XbX7Ts5Urva73+wzS4bgmj5i9OyvpQoPAwof74bVC3jVEVqZ
Yuq/trqLnLd+LZi5i4/n7jAJRkohtm7AS+teu+i6tf/+Jfevx0eaezp7ZXPscQjEd6uT7xgZJJrn
A7VNjKVsKZ71hUId5R5W8LUX6F1kMUOAMADryxDOJ2mpfQZfEdx8OWvMNd5EEvvoL0/oo84A6g5C
fViK4SoY3Wh1QnZDW3ntQPesxn3pEOJ2677nW75dawPS+5ekdXmWaiBuhtmQbJnjAzjPFNw7BEkj
mhBxgXRdqaaPlcOFEBe9vtp/wqRNsLOnuppAkA5rcm6XNIfBgzn2yP9A77AGKvdzGFJ6levAkKW/
5cly1a0e+HHfrnVYs8Io85oKTyIFJqmTR/NMESpffBTiYIgaUyBU58uzg2cH+D4H+Xx8elav/j5x
vMC/3T3b28y0ERGfL4fLIjhpxSXTfUjmEDBl/LKSVWQq0nkzmpoCC6UzydrzRVZszES5H2K4ugqH
68aK6w+d6BPNhjm7sLFUjQORemP+hzWE+4+Z4A7/27G4/JgLTrSJSVWBgljfKilK+mGa7VBFHaKs
HHQyDxPHXBrRjQKDJZg7eM1E5LqrNBpEDFlXF2s30l6uQQBQhIv2A0hLdnneW+V77Q2rAdL/CFep
XzbCR/OTW2fMPlVx2Jnjl7I0T15Gc9nXK6/p2kBCLbrjPYJXn9UzV9zCQ0cpgb1/BHSthWcrdHpl
716T6HJLiRNwutgkoX9IOAe95Qj9Tsl/kxIDCZPMS1SnNXp/IosCNSfeu0gv95e41STL+x9HdJh1
RvszX++mUiu5zNYZ/r7DyqfXpmgQJELebkY0IXlShb+6pENb1SFHWrfOJqHJddroy0nXBtdiMT+S
7WKvHIwFOey9Ed40d6yKMYzkVcLj8qiij1UGm+QovCQ1HlyQXF3a31eSwXnd1oCWcw5VaBMWySjr
mrIJtfiNRF6vfb/dUsdmeuydyal3n92JsT85nFnLqTrTA6uoXrWf+Oh/mR2cYyMKmSf+bcmhgJHn
p0YTuHFA77xaKUPeBAHN8XFwDVCE22yhGcCzlsdNOGrzeMe8OJU7gbR8HpHiz8RQIxz9LagztbZK
JsxTvkuiF+H89BUbApKBxYNxstVi6s86tmtMZZmnhub+FF/gFoXS+hytbe5a43W3LF1r8ci+Spuv
9qKOpA7/fzbx3WaTwx3qetrLWjbDBk4fbATIox7Ud4wU7n3crI1UuNSj/sxaA4UwblNcGSbwkeJh
A2x0qDoVvLah+tCWOQ9lv7QQbuTrvj92RnbGHSIxdq09p1x3104fcU6IVZM8lALyN6kSOxHn4R05
oLR15GGTKXHjZVJkQ34lnKGX0S+BayfzPdWM4lvwmPh5VkYVCvSIt4urCgwESLZFNeeolDEpacr9
9RjsTpdKbi+3xDX7bgsYQ8lUSjJR+j/crqnMwQ5Ho1XchlsAYETUr5t0KSzy4AnwtG7R9msvxNmI
S2IAj7TzKMXa5Gvo4Kh4Bf2dGUahUsDcHvFi2RJ591l36wtLXFshzOZxHXLrPS0gitivReyOrtnO
oeoz5XyQIDU5xXjdIjyL15uA7rbogYsE/JEqy/ajjS0s2SCjPQiWO188zGTvSRQHg003fHQABGSs
8TFwpYZFI36J7wI0yOkpI+9zRgcTW+pGYsspQiNHoMq7jkhWxKNmonZnznc79eqJF9Comd/0tKGU
YX9rmFj6TbdqEgCcNGrzd9I+AKD4IMEmI3aJt+A0wFLsDYLIsq10idH6xDCHmyDF5l7twdbzwNGS
z3I15RUGrPn7TglvGuavBPLTSY1WrMolzoUF8i10oH0ELiYUTvtCaZ0Qrd3eNE+bvdl64ifCeaTP
OQPU4Aq1JZ4nzxFsJR/A7SjexhKzUrZhLPLwI8duC1Q733qJOHawg0MAmXWE7/wKhL5NtC/c+trY
eWzOFWawPR6+jOsuhL0c0NKXj2mAXlgKJ8d6PGXjHiP8l7GSz3pXXUqP7BOCVUFL9gtv1gR+Kmun
G5EGBKUeeT+F728ycWitHDBZQsf96s3/Py7J5aEgKnCD2qgvwvVLxZJednqwL4HXKNmcJVVJkXTe
vfbsTAE7V+VeMbV7KAFZYFdwb9juE4oxtwiyLcfny9iFlg5av0YYp/LM37aWCy7LZDtGKoYbVSPD
Z+d8+d8u7kVtoJVlnahwiNyIYzrcAJ77UIZ27xdNG4jPehufugUty3OrE5SLu8igTXgPNc4CFByp
R6cdGH6gXRJcrKHiRxVR30/37Dc1852WnErwt3S1uB9n00sU4OoWZ9DSDgOF/exbswjgCyccIVR/
8QgOprUYDp7xhX4HVV8vKpeR9tV+zswQCSesTyZdGUeHnry4f+/kjRxPLd31KsrKgNOKwiy5vCLf
h1qSnbhx7J3d/WqB0mlcaqWErQve4yLWeNzP99Nu+6HVVCWSpXcH4whCLnM7nPbhJmxdvrSDtH9o
XKZXF1Ijump8O8zfK5xVnmLfeTqI/lRIkClRPgVB9HQZJoG/VfBdu6HJvSXGsLkfsR1M+nC+xOko
ApKXKtqbDV0FUwcDJrd0wnCU0zamR7w8jMJt1gfeT6fVxdg6vg+MZoXxViVFVQBkFZEMyCqt1Adx
0pfinxryr1nGJOar9PUAcZUrscsAihvFutM6gjtqKcBYJcgAb9+MBYQmYQt7UBsW5EFo6csxa4Cu
eohN97gcsNhu/gM9aDP1eS3RZ9U1IoWg4vCPtlEmBspXX/y5Io00+xxzdCY4BpISGzh0y4bJ8TFs
nklgIm/vi57p4AMRbehDHn8qyaG2PK4LbYpdvVLeYrs/Az+SFDgpoLll+TCPUZ9J0WMrTyupaNik
2Yl3JryAMVFjGjcpoJ1X/NH4RHwVSui+Z5OUzKG2KGwKig7dVicprE3kX5Ycimpmv6asLyVtxt15
KRg9C4tXdvTSNVEnetSjgrl2DILFuS6kd6FIchhj4bkYi/OsAh3lcFAul/9cMSLqxVJlY0ChxfIp
hHJXCui7WacBrEhbfqmHUd1PO00FRARswy2CBQP8PgvcyebTqXiW4b7Vj1SNauPd7Ot2LuKtCvN2
DqqqQliLGVz0cCNjElmo9DIa74ztE5INc7dgLz+2OknY8WKE7iQjvMP9vUoVzXa+re2Emyqdm/GN
ASEzBRFh2SvNwYrC1EXKFaOCfGoboEUbIWMNhgikfkzeA1LqpSJaHUpsnQgBx33IfJ4wRn6wb6LO
q/B+5l78jyMuI+nz9iE2/dIwO6Xu1zYBCvsLNf6S8zl2Gse2GG31+fQcKKr5WPzU7Kr7neSl+TUM
DLmrRIOz0yHNEt1YIk8G8FIlMNN4tyHupQ3wDQK8rpbaftU+PLRJqlQoY12Ophi3ay/mTdULCAog
zYh/p3xopnayrLql2j2cEfkh3lnpNb3VkeBMUPowzoWWz7LlnlrdELCoDI23P9mdZwpdP7b07vD8
GfmXAiRHWDtTiTBt2aLffoQ7A8cwxru7AyY7xDfsai6TBOsnV16kbb8wTt+ENUqRanqKHyKDatbN
GPU09/+w+UwPdorWWa2Vh4YPZNjOLfWRMunm/4Vz1DOs0KEyHopDTlLGJcG5okyAUY1pH9aMsGyI
lBJmUpQTDH5kO94AcE0+EpBBsWu+q/3byfm6lmxlmTbStVhGgtDAHJx6YC3+EPHHSZgXHSzW0thU
7CVdz+6M4XblwlztT7L4P264hoCWPPBSBVDI660Fns3nv6IMnjBzwdVh81K/kBGtZXVQSxFyzRCi
n9A58BhGFFJ3OtXrwYI9NOMz8ApUkhcx1Q26YaofjLFWOp8OpoUFGvGHCkSMgujDgtseomB1f3qq
+Ray/95j1umaADKGkmcugddJUZ+OLdDOgrOgFq0xJ5/8Uk5L2n3nS6QDREEp8jeE6IVD490UE79l
BQhVKOB8x52nlh1KVPY7bTrhGx/6Z1QItBlQ73JaUthr+7Uoe/TpL5nA1FnD6YyKP8v4pMJb8Hn/
3o0Z5Uo2ZfKQsV7b8QYWt8D0iglt6T+Lqzc/IRFgHwSOHa7DZmrpmNn57g1X2U9dOniIoZRtLcj+
jQKxZ5F3nMHYa9wmnf36uT8lOd/ARiKESv7hJOsWcBxi5fOipG3Me6XCwEmtvMprpBqASNDUvmIZ
WeVwW2mz7JhN4NlmA5Yz5F4/sIZK4wvacGWan/+57t3r9ewjObBrrUgRzoC46pkJjEc4tRFhJ1HP
QS3F0W0M2wp4mGcR19YMfTCczqiIc1YTql5QZZThWfSX6rCOU9QBSeWpIkw0z5NISxE2sTyBrcxM
QDPG6Cr52rUYQG3vkq4tP+RG3pF3oL/7uklXdyFSolO3cRFen+He4Q0gqGb3OBiPkPd7WA2okSkH
9WQHeeSBb4h3hdmtst06Y4khAy/1Ka6i+l9qaxIvU5vQ9KoD50djfT08dBpDSMSoBkq43uJrYEfp
tmShunL+Otxwq3BTCCZ6ahyt4fmtx0ZMI1ESRV95AC+zMGuldlfvVdqIgC4R+61T7PqxlVtSI6ym
OVTpKaF09/TVd7QXJ5vACuW7b2+lHAaKAzGlM29tlW69gEMUN+a6sA6KqqEmbpZhac9OjXnvUA+p
KD3FCnF53p2hY59DRGDUNyo0NnE4M6f6QhQRhcVKpIjvc8IH2tyylFkMaBVvA1E1wYNUYiXFyads
yYRiLuMBRCYY2Z8UYiPXTdxvkMry3NPRVvCadkd0Ts1o6S5o3DGRsO/PgnX4vQ83Ypc/NscymIJb
Cz34SJ3dA6Zwhvs1ECS/i/gyWTRhIbht0wRJIiDGO4PVoj+2N4oE18GQKM94cpkMZyuXrWe44m26
oL+l50pzUfgaEWgZRSieASEMgYaKbNGlAv38HTGjm+0UIA07kzxf6RBCjHmXR132VjbBbvs1Fdlx
pypKPEfTrIFjsSVSmatlptWMUjKU66iqwM7evaW1FntI2bC5ajD3K501tRM+t1ZFnHGv4wNoUjks
opokdykMOXnN3Qmj0HgF1fuJu2F2Gm2tDlXwSXmsRBC4HDyN844+ecNWOognVJ6Zhtxi2WJ/O4Jz
FYhB1sBsm9BNPF2E9qDtjVNO5DjvJwEp/HAaZqJNcdEXUIiv2+oQCm7wXxb8nH4Z8qnH0FSLg3dL
QBGFcsDX0uIkxKGtrAqXzMQLxSlaxj4xfRVQQsBUSOoYa0/dTWBwGR5ZKxXscAPhQEke+5OwPi+0
63Uui7RtD/3h2dko2RdI6iMSRG4Kt0Cs2B8B9dPyq90Ivb5RmxT5S/65vZnD3q836j+9xNFGcWH8
L8ffopcnySOniS/a+q0gT7o4unEfiI2GDF1GJ9b9mBwl7zpX0fsoBhaWQINKrJdr+B7Ib8ntXrZd
u3ZhRANgsN+m7pNEkOb7PcgjjquP1ThPY02B8caCQolTuRKrVS8djlS/WXCFnN3DiD/ilDv6kr6q
eASlQyoYFKX6jbzc3gQCAU6dWdR4BsXmN/uD7MzIKLPoHkH+6wrG3ADzqtu7q4jjQh1ezt6gRrTO
6Sg+LAH/TD3jAarI0MRC10PDDkWWpQz4zFCBAXdLonv2GPi8H8BBtRL9DysHIAnvbYrx997oNT9F
6G9tYXP+w0TZNW9gEmz0G0Fn9wOgeZdqEhC3DOHeDgX6S6LVzVw6YN+WIP6pAybQBIDnz1EHbBpg
+mGT7f/Xwc7J03lSlL2rT+zb/6MImjosrxmyfWa2atrT+NPWChknqqhYQzo5G6s2x+xBxhjREscg
pnW3TUiIQw1X3d1z6fIqCc0uQtolQ0tysLMVtfNgJYEGfT1/ZygAUbhh2oJOJHuYzp4OuTWNmJar
Ui3az/odhhasdS/YztddimtOQSkEzCOmzEqHHwFs/w5Af45T1Ug2B5EbwDTyVCoPub3l6n86O/U2
ULtc/XPsUUgHTfacfjKGw9d1AkO99nK2M52+j+cl1f3F/VGISUoByVlWFxr8vzUzbHINY7mdMJwO
gF6DpfGWs+S6KC30aPm2wUU/r7hYLIkDMFACVsJj4H/XokT/HPkqD9m0+cyYVVxXi4CdMMw2+/em
O+b99tW3EGoj5A8JZoqgekYUTCdlDxnKUpHB5ZL8xP9KnCd3l2rbeZtNxhHhUWDY5JLDgglTZzHl
J6pWVDQmgf8qG9KAH5jbGfHLo480r6Gh63CFDDbhZqY2AEGJ9PRMFTYHdnlMWkIOGqI2bxtEJu2R
x+lKbsHFmMJxUZoYRI1A04BjL3DIqlWuUkJR3dt8cwybet7YFn0gY1cv5eb6BzfxEaoVj4ItHgb/
K8QDJVksdM+RhHHDHGyz10tXYFTjpYP5JnrkIFTqRcB6o1/AG6tQqFbjP9Du1ZSoQ7xdQe4/Osn1
m5uOk625X9Fu/GU5VRLHn2pGQia8ZkoQL49qyO7WPVS48vhv+PNuC2fdhr+l5/mbCCTvHs6wLucA
Gx8ShuzTChDdWdplNVoGqaxmOL7lVDXZwFRzZoXrtlZcDjc6A+M4hieEfuRIM9fXGloZ5MRb+pqg
yaSw8TW6JQl7uGUgSxhUP4Qy+NSCC8xQdx2in10OuaFJ9y63VbWTcYh+CMuGaRQgjiBojHQDaQqu
LECLz59kLJPGh2vM7ZahuCIlBzvDXyjhR7nZgrM3bo0DeiMa4JwtR87KsLRQvUaIpTrklOzBT8cK
fmIpBjmTJJJxIh4SyLGWXabNbkxLegtZCmYOA7qX7pX5dxvqzMtsMLqEMcyia4CvsxoI8UEwByzk
n+wDtlRpm3SEdAEXaa/ZnqhF4zSWtmKnH0lDn/OGjNpp8okErYq0hlqqlDjOACk3/au1x2jpK0hA
DNGK41ZIPp4IXWzLdsfNzOZJBHdJyB5vgAPlw3CGw753Bp7ewu4mj8xBTsmxm7se3MTfDqUw0Pxj
TX0+NlbFU1yokXi2/WbxRMpv6Ed4fhMEB7J1VbO0t2yBMHYsEWTev3w9/knuygz9gC3+QjuGcP30
OYqrBtOxchTcWLre9e3VrZPFWyKEdanxTMdzOJhJ2shxs3tFadNw9+6itBuO+LrhDicFocVHzMJ5
DvU/YQh6Rc4BGlMYLKZ7Iw4vgdGG/1fcak2XqzlUp2eTGbxKt31Cp0YREEvWsmBPuMNecnsGt4uE
CzQ0K1LxyvRpCb78bNJcbF47DqzQXd/r/ae5BFwIC0yOupvuCodscKgyaisOcGJy98aIs4pmwngq
hAb+Vgh3Sh13VQvrINBMRjpoNt028el8e9w3STIwGh2+Fg7Hwwf3I6007wBrhqzLf2XH435+1hAA
UM8jeF/A3KfWVLCLNieNb/+sYOd97FIO0SrHMA7VSBD+fgPQ8HuA3zaWXcrNw8u5BHfdlybQAuA7
RNBWGE6yT3QQoMlcUUyj00/yqO91uMxwHFWZ0uclq2vjMIvCafhUJmup/FiAW3WRj6VRpU5sM7XZ
MeZ9UTHEMraUF+81UPl9WlvZoe/uo4p9442DqEN1/snsQ7KRZVWFzwS91gtH6THpIiZ9aNZRQGpW
UQhlB0KucdzWpJJXfPVnwd3mf4e+DxvnJfxim0Xit9X/KVIGl+CYj1ygT9yGH/+bVcey5QWxtShY
sb9GWyFiqCvOm60ubQ2cRQwzbRCq6JjQOIe73xLSyiha3j6u8gxJVVRWctdODyfatmwNj+ipfxqU
XDnG0WJd9cpiaFQRE/StLiII3BpCB92fXhIRKNZ+EnGCuqWJN0sUMD2kGAVnpeLMLxcBjptrRnFE
d3NXir24lwlSvcTAj+OBIgRvRPDObrShj1NBkbyV2HLWALnDtSeE2Co32UlMVolgFqVhVKnz2abA
n7Np/1JL0QMMdkWTODcPpb7G85iuekR5Wrkn1Rr1v6uxGDJyTSyZZrP8HRYqGkDK+MP6I+l5psH1
vgcRJ3I9bTUmd4YTKWQYTrSHBrGV0l0Lu/33w8wQAczOzh8wPswc5x6mexcS1gNDRpdYfLXHn3hr
qEDShJTRJmhuJYGcWO81RVkv2t6Y8k1J1iwDPBIJo2IqcN2vmXpy9geiywXW6wCn8a3IwBqEBqo7
o+SgHkjBefQ3v0jU56WO81pioa7i1IH8PTmx6Wg7UMeUyREH6LmQ7hRO4z0wMXs9tXP5Ywsv0mFR
hj8a9EpMKmmCGKQ/sPy/Q9OTCAMuPcSD3+bWYUCRf/pgXJzgn6diln59OObZmEMZR8EWOfOEQ2o4
KUysO6ALrUbL+Llljo7a8G1Gp1ZHeGrrj9e/MeIg159wAnint24cituey7ybX7WCu0HyqyTv3FE6
aRakvNvLSmr6tKJY+4KNokZEL8bkEhOA+Qihr3ZLUB3IfSx5rDQJgd050L4HCAPJMjM+nMaXV5vY
ADq22sKji0z44Z4mvAlriqiFU665Anr75Td2sgyKvnDhAaVCZBHnBbQtk65qL33vddfruoJVk+Ba
Mvjo9moT8e8Wgw2BFrU8Xyr9VtrNueeCTvge4EQaeUyH59sCjr43RuJUzunXlOuF7M1/CjZ+JmN9
h/IZEAO8OT06eL7kyRzLSBNDVP90q3bbKlM5cZuTuxG2w4cKlLk4H4Lj04SpYvjaoK74fhzvpGXI
2JwMRpiwKdXeIR08qm4l8ghUYjEXuGJDKSxfdrHX1H/KjJODeR4KC3ELyiI1l0gbKkwWpH7YGR1o
t4iioXye8DuD9sJv1D6Orxq8zRM4C65+4pj0OjF7SfCo/ufSyykYYkohfL0Z7IXsx9Zonq5+wX4R
Xk4evLUd9uNfIim1wxI8OCqIwANTWulfn/0whiULinu++FqU6bZctJkWzO7YMBm1mvn/jW127BJt
5HFx6hkviUw49BaobqnCtNg/PNqiopY1f7jXjqXLBu/qX9tmryXzBS7Jx9ms6aJU1Mn0RiCfiON2
hR3l9R99bYwJlYlPcailSmTr23BZVkeQRiHxniF2wJsoPu5H69BNbDGMA49XJa+kVTexZwgi8ubU
CYgTORgTPbeGglI8l49k1bwdilPyg3b2f7ZavUvO1mfjqYxD3bG9enr0akEP0YFFbtDVDBOn9IvI
3USD5dKmglXH8bT/JtU7Dy3EpJGa4b1u/i2v6/+e9uyKBLt+ZGCMvzGxsH14nCzS4j4dSJb0C69J
IUVZrjKYJ4X8Dw0YptVJq5PFn7ygSnksOZ8lMmlWnbbfEzqhcB+AtKDAWtyqbHkDfeEbH5n3oaH1
UYfkSRL7yViLoZFi8HOUt+zTb6U1i95/2VdTGsbmWqPlVU3O3lgQLK3lmevqEvbYHNtkQFTmCC4z
o6iN23ehRiN8plWA5FHw8YdK31t9ybDq67DWpdQAMkxx+DBvEWeFyxMIOemxeDSetRM83uQsHKNx
akNsdo4Vbr7eG92142qrJyX9xX8HfHy0bgzr5ZECs/BSIzEr/iLn96ZGeepw38TmISt9usqHqIYs
wamy1uxGXZx+Em7MU6WwDXqkcGGao/tooi7gDStMgcGnOBejJ4FwIUoaoiRUcRMEBpVKtcd+CEJl
1B8YRrDHHq8pPuOgW0wH9GZZGN771Et+lciGvVxHjNbG7+SuPSBFJo5NUrlWbYUOCsMxfwhL2oK6
rV17gEwD8Huj6oyYuiFOeVmP0AYBdrvLXOGbcDd/Uyhyg398+DJS7GZ4t1C6juauvfM8clds0Ux6
8O9bmkToEKPqWAHkHUl4CgQUrjqXNEwWEtmjFHNOZDYinJ68z7z508steYd1IvDE7wC91euMuWBf
xDN8UeJwwfCxhFyG0H5xRMfmmImg3EE9Zq1S0sDLVB4gNZjUjG4WjxHiPZER7a7AHdvqprZ1j4jN
lk9K+1jW/t3Ewr0mtwKuWJlr08Ex/TKo1qpUpLXXFAPcvoC2rUdeWN6zMArIC8jVVS4SrQeEsatb
h9equkrN/nKahVRB/i5+bUZAMfn8DmOumyW4hxUaP3UlFEJgfI1W2GzE8gXTFGb/yuKJp/UgDEmJ
Cjsmwt3KufWX+G+HLOls2P/a5sg68nRuSFjhxPXaLVBZSHb6nn1Mh0+UAoczx5tPEoMSKhXays3/
q6K4kjt1i8hzEUgSrgx1ejjhakk8ALMao2lw0BoB1neXaBWl+AgCVVciW3bB2748O+iR6tz2I5X9
uhULB313btpyLhP+RV1hL5WKlOn7mZwtyQhU5u5h0T0+Wk2Df+kxsOokhfM/dBdpsPgoWIJZpKTg
PGPi9ztSPoNi2qbX9S8RgMXf+E/cCgnL+4hJFclESviJicATo0zma7brBs2GksFidI0AG85AXCNr
+RW3Uw5A6W0cR+ugrPmGcpZh4mEZi1dih5MeyRTXwLgyJA2vth7gGKSM2v2VU0tGFeNzx2RlB5vq
xhDlGk4pxtSrgkb1NSeg2N2zdpasEr5GaK0b9UkcWCG4mjWU0q0E9fA6dudujqMTw1hQzbQ0LsQh
cYpZwDpxE+PFuwf3TX8QoVIC2/9rdKhuDZa4IV4kEMmMFth5Lv3TnWYCfP449iidy4ONcy0Z39zS
8znlb/x8K7Lu7ISWDPdjJxsSzjou3rIYXt52cZOm95v9kBmMOzqzozQPnR8p60+SW/+sfCEaj4X0
SXYljuQGVsMQ8JbQv26EeXfjhnK1pUven+XgnLfrCoVWa82VWjZyrYRjIqSqBh15FbDjsdA52gAg
PaW4r8nxAFg65nZKWx2eANryHuyoG1HPOJ39K0R3GpRMqihxRCDOmj/TxiVnaCz08I8tLbwtslkB
GH7G17F1kZV3deGmKjWSU1FT7dYFveqpyyKOUswd31IV7DsLI1cJp2IqYtVj75Gn+Tznw/vonHSj
oFmnlJBAa2ZlyeMrGBxYuoC699ZRJY+nn8rk8RkflP2j3AVB1eJWIsM5gVKtoAtYvt6qITyL+3bl
tzk8YQ1L0Ajrzhxbcp9F2SjrQa+y3oUzOQ8sXskU1w0Nfxvr1/ueW0FvmAPqUvWuCuJWdXo/tvIt
I+noH6c/L+2uSOAVSOLWQukxM8seqUjzz5oamNdwgnrs9l5/mAIvGJOD6YseELbrI/uoFnNfz7Za
G8lzu/sjskj/a6YbEjBIy7yWYxGTL+zSraEzJ8CLBh8XudI+YhCzlpKi8X3Fbf3E13ckS84+jJoj
4F3zOpNTWj28WOrqPlTeFoRXCw/HgwU9ec70EiL1qxpzn/nGOFtRd2LNCUqQvs5BE01saLb+JC9A
xjG883RRJa0zSg9TTR+4U65xFfFWnz8as05U6wScnO/8bYPi3rFMqLEYsuEo6IPCQ7icv2NFztJi
wAwRqmU3iaDfejqs4bA845AaVRtMUqXc22WgkOtBdVjJu5U6px1eBkG+T3bEYr5LrpUJ7mqyX7nw
bTKM2nIrScXHa3/yP6AZRe5vWtsDT7edMsmWNxKQhduPEUJ9XK7sM/5NR59X2RR2BnyriWRNzV9l
4Fbo0PFIy+mlGGqx6I1MVcXl5l+U9T+DKypIZx2IMxyMxUQnDn7ilm6PBCpard8zNAUBkC0+usP7
DP3QgUsMmzGQKTjOF0uTV6o3ilfPLd/dPn1bBezhVsmnW1lQxLThvNHIjWluByP9N3pmtrf2lGnS
K6kCFWt58v+8M+81/TDX2bwb5YKupXvtmv3KjKkD+JC0Q8QKUFNLxB/87W50W7Ho4oE6XvGVS7rp
0SG1/iQKsEyjmDCztdgO5Uy01QlvZbpypmBKNodaq+he+fuLal8gKc1OiRzAuEU+yDBCstK8rcYG
oU+VO8L5GVhqaVhpjIibAKftmv2AL4B7oTFR/SXR0MqG1qe0HhFhEMnVWRqSQBj9dU8AaHd/zFxZ
thhS7nh7h/x9jt+wGbBIzFZw5/AQ6zhcq0gviF1wHHz4auH2y+xsmfK2lXRKrRVJZJzCtvzQKq8A
0kLSq+9QY2VuD7hYc7xApXOM1I20GkzU4Sej53WvEpojvyKlgNfyrhOyaIg+q5wmDIeD8iLyvcke
sTFH5lk2q0Src5fsL/7xYkBThA+Y/Q4wWfQqrZQCMS6f1q4OMU7eb+ic3+yyK0Ow8dafjo5cOxQI
fQwHQYU4jfw0AWCLMsjzu041AytsKw4w7c3owabb2LT3YK8bbhAyoKGhAfK060wMBypMPS/NvmO6
Rj8BlK7gAJM4m5ZUJY6GSCdBI1/kqunjC6y9YIuEd9Tk6Y7dH5bBUvB6PQpt1lcLoWh6Ps2/NPEN
jC7tXHMZ2ebzy6czxtOvVkovMc3rlOGbnDQBpqf67lqvF9kXexT0zXkCIMY8tRU5hDlAtSLIU5si
eCx187wp8EAPXyENq2DMhWKn4HwGWRdC0FoBkeTTVB+F84AprPPaqcjTKnlVi9iTfXxvXCN3126j
f9f2G7aAgQeffplLcSn6ovoewnoumQxigJ1zpPEhFObS0/Tgso2oURw1Eth7Ipqv9x6y+3QbvueZ
PaQhcWYxyaI6Nz/TeSbxmt/Uh+stTyifVNntNPcWoHJQl+yFHxh63OAv8mwgm9TD4H0F5ByzKQ+z
U8+38ZKJ58U7OknWRD1i2PJXRVVVmJAZKlJNRJFVVsY3/ls9cQWi/HfyL20zfMM/+iU4d30Z9jmw
sHC7+gngFBr6OqCbfQFBb/GUoEPoug7VXk+SsVvM6uy2pd/RJ3zLHFvG8hyOBZOg+rqgibghmGbU
uXcyhqKphdHM4CL1AHssl47fjoc9piYyZQckt9zn4+bzetRE7bT5VU8QKrTm5NeATMjKHRzUPEQT
fZIy5k5n6+vI/HOAoi3ZT8/mHyO9tNi7Cv83BQ9eGoWGbgLkDcNKFzUMRCYRwUONW8zdqL2ERVjB
NyQV32p1J4sUEBAu9dUBMYfUBzsQUeLwsMlCWxNHXfLQX39RoGTp6OAqYSPB/w9ajN5e3aASLZGR
MCm/4bcP+pX5wKya+2h4DOXfF2dm1H6gDOLDnNXjXxeASPHJd6FmGtoGW6wot+DMK77C120+qp4U
Zmr+LM2wZQc84H7sDxN6ZHLAwbQZp/Yy73Fb14mRIvoC0EuLK2XkUH6rPOfigdcOJjVml/GlxJoA
0ynqb2vZ13libkmhWpmRi9vlm2HM7vjKMI2/57a+PEM6BpLwAeaapNGHY4qdFp/MyXI9iaGZjEnY
TFoSmAvgp5KHizXI/qQLzzUJbNPC18vvSi44t7plaUyGbakV6HOshATv7G2TVtdX0YsILk0K2sYl
3ZhEZBwkaghDV7noA0dAN18/zf+CZjhsVCn3t1QaWujnnWAh2E3xgyJqAg5F9dLYWLKn0bYF08KP
PUlTOjcGieGbFqn+zMYZT7DXqKhqAEiTkBpW+OpQ6pD6jQNqgKDdpiNNtcagL//b9WdwrSb83rIo
SB3qPQu4J1S8Lq7kcZWLgD04Q2wIUIEL/mlE/ws7fVtL2YuTgbZZR04/cWRlfKpXU9wMCzCo+Qrj
ln4TDdbSVWt2DbwWHjlAoawxJCuQ+Er3J60InsREFbeTy2lkTXd+r73yfR4zUA8nKe230TsgSfVQ
ndNTwsBkAUfn5atyjwLJzjUXonnBQ7roH0aExJ/v6KfeAYN5D8AplsY9IO4J76CdfUCPoyrt8XaC
9HMPU2NdlJTIB7YewmWEi6Q+3qS0kphLj0QnxsJwEJH6A1iLLyCUzIT8rVPSqOCU0W8AqxOU1uLn
NxH6hHcvbg1o5ITBru87y+jApxth9BXeZkxDWIsGiNt6o2cBZZ2HyGoGV0dZn21UQgcOY3t81LCe
mboFxziHN5sIDrK4/fd5Fa1XH6sxr7AF005Yj/XWrpSTQUvjy9WCn+qKmfj06Oro6ijIFM3lFYh+
m4PPcaTF0mvtLkh0TO7ib2NJMwZXQMj7k57+n561/vH8U3+N7WwY5FIDGnNHpwHHOY0gyeQ7zUXo
0eqKlzBaCJ0UllS3TOBrrtkeS+DLXIoNCRBxHp+pu7yQJ5TttxC29dZNtMtymOxuY8hzt4qsumQ4
oY5EKXs+GTZ5vN7/aPyVof34UY5ocesaHXFfx7F/RxnDu/6nf7PkJftTcXCj2f7b2dnqOkXhvBne
K0mkD2oYPV5Ir8FtIAlObUKlVAF8sQ1zMYHSE/0jbLVkeQA2nWaOaqZUrE8SAVEWb+bXiX09oMRV
JER0b/ou4PjrJuAGpzm1iPXeVfkFNSYEMYLNh9h6dqnPFntoDdwCeiCfoXJjjCCXtQRRIb70UZm8
Ir7M5yLqIE/Idrs8uuLm8I77uhdyezSNRdc89or2bVdCFHK6jv+f/9aTA6i+bNeITCGRElUehW6K
igJ/9ylQady5aUgIQ3HIIVH2w4HDKS4iR8arLRpeYY/V6BG+xVau/kQStlXgtgKbOQ2ABeNBhIfB
IgcnGEAN03XWqfON1+pQiz664WNiUB9N3lvNbuoUT2eCEbwlGTPlFRTmkunYl8FwrFBMW+WB5qvw
CVheK1nYcK2KZEK6xZM/vrxiCHvpT9auskZYEA+SFtKiuSxrpZaXpxCCM/4k2pI1931nsGwum2XF
W/woqyb/V2aKPrHdboVdKL1VCaOkERQ7oJHJD6T/Z+YldPEuZyNzdYcsT10jnksKxFUup3LYGT31
cVGnaEhJ1prCF+FTOz5BTidYljeYNygM8quutoORLfqmwMN3F5L1W8qyr3pB6vFRKaYjSfyh1sdW
jcfktaOuyCsMRMkxl3SIS4C3IQzT9TpB+ebSLoVihDZof+dnBab0umE6pZvMNQAfWuwRN6yVvAHc
AF5vfur4HvcAAvzh0blah0vYE95vHw+qSYeJK9LYFREt3qmUj2naXjtQlS1ajmM99tyBWkTq+PR6
8tFkvau3OeovlbsQzGIUEPRMjS3QRd+DOQqQVTA7AfOPr22XOgWyofuIGOIivj8AZ/yHUyB+b5xc
QszmhJ6BiwwXA1jNMBBv/+vA3SWoqmicRuuJav7j2ptji9rzSbDipve1Cogwd3ELh/J0pEqwLzPD
tvqMIt2/PxM96+ReEX2JvjVX3teTi3NUaqzYAJLtbkhdTIDL8a2u0jdUacLRk/+5F+y5zguqm1VA
ctLDOWckLYqP1QE3IxzDVHVm4nHdE41OpuEcRC4A1CjMllofwFHEv/ezgoOBbGE9hftX3QhHIEf+
qU8lVOy/h3/4xQQ5rq5VUv50Tc40BnUNYIzwbLv/7AytE88QuWGSad/JWvn96rqmyLz/4h1JReym
ohZzd5K1bnxLHTEQY4bUN1Uy+bioorly+zu0/o87lgbeVxJMr0arEYOUB+IO1cpYySpJ7UUcLyfO
AcFG5aO2Rt2U2FXYYl0C8bcQmvGy0Cplpzj0MDkuSyGJYK1yT8xL70V0oB5V9LVHdt9oslEyEYxK
XhdNUzRA7p9zvu/KHDHu/ZRXuqrfblj1cwISN66aenDlBWEFMDoYPxYxgEke0bgCRgmRvrJzQzSD
XtqVOicP80xl6C+L3EaeBVEkwevgsJ7MbG/daBNT2nI0LN6VZbKPNd1iEh676KDpuPPZScX8fNlk
NUvRg9tjmqOzFOcf2xgk3vVYxUnfm+wt0u3qqypcBQ2Opbaha6tTkNvNJxCDEk7nhuKj1dNTE5+v
D47cF2IkwTEiftmAsNR5e16erygriQQMmTNsSdqCaSS7wVG/zbNjP+MUBfeRAKnezZ2bDFicD0z3
iGgnnmbDFS897HUQWJ1MdqdF6bQYmxKzrWe3hjsYzb3hbuVugs2YfZGhys9s+oREEsaZ73fpZN0l
YSHapL8Si+ERbPAz0de7q+gryCQz014i+br4HRkgwa/aedIgGKtlccyxDbE+3sQN1FdjXZyodAG6
AyWCabHcr54bQqSPfB0BByQ5uYoGwzeRymrEb9j2ze4fr+kIGuY2xYy/Ppcz3WCBfxJlMSHyL8PG
oJWAsguALjJEaync+hz863o+PXLHr23ribMfdzrAQG3nW2CwhE6PXkX+MjTGvmL4pwWE2j3ZfQSg
9t/vHzGGA26+4TcnZiI/fq97Qd9QdB6OIy0Q1CTvfJ147aCGrel71F+OxQ+wd+oaPU0/TX15m5Bv
Al3C91uVesxUxiRFtCDubCdZ6FQXUAQGLvNPZ6FL65gFCQ1ubLWTKNzQIT8tY/LE3qwp6h7Uc2Te
0RUnyj8gZrfSxQawbcVnAx6DDGC7ZF6eOJbo7VYNQDd47agItPaA2K0U9e9WQ6KZ3uisBerx6Nie
ie9kRK3sfWt/WxpbG73SAX4PaotTdScK/WWfrZH5pcP08GZr4W5z3RQrvaMYFNYuIZB4fuVAhX2c
hgHvlTfWsKJmrMLrWx0NwsKCxRyxZr1ocCepMtoHO3j1t5JWXmaAd518tNHG0mmriaWsH0IqGjmr
QhYKUvb9QKU5JdNrFrq/nxy4IxNkOMZ22xaEK0FVYhQI+h/pKgDZQdcKxBJvPqRxMOc43e1ygQqU
cIw2Ny2y1ywJHnl/OplfJ5ip2YfBz7h/25ThO1zg6I7M5K1yTT4kpTQNt3PAG/S392UJL10eW/z8
ZeIs4l8MvhdrR3iEwDpmpXjulV3yeYHKQBQgUO2YeWRNjBCPlxQeEzmxzkwu6xCk1K1Letv2zJr8
DbbDCKGyG6JxOLZhug4RZNFh2etZH9uQRKzRiLqR4y9z0FO0Z35+3BBKUyziArFv5QVpL7sOVjy+
NsPoAHxogMZXhsOdxhe91Dl0XHxFGt5cEF+wO8YpEZJjAsaL74YEg+EH/1uWDhYBPnwXm4aW0+Pi
Ks3zoG07ohHLE9GpF6/vWCmhrr6DenFvqFXdecJe1bAm8NziX/SLPqG4U9dSIbMs9tLAx0PhgPEZ
IpstOO8s8Pi8l7OOYaT3Qr8/Yn/amzHTZRQbE1giwDuC6nWINWuS2UuI+IPU0rl2T0yLWuX6Eb6E
8SzJu0u2Ji8GTBfdPvcKWCi2QCNbiOYsETGEeCdGoDGZ2tfBCsb5SzR83ncw45ww5lC6B+mxo+ge
0vwKPGSfBJfRWgkY3ibDta+z1VBmaF5qRc+6dUXQxSMr5WZ6krbw9UjAdwhm6IP/ua4vC/vx8a1u
CpdXhHJ5Fgod8+NQsd5dpgBmzXqVhIv798hZPvXyaJ6uqfVSWJprSp7WzzsVhMIo1EE6btneW7Qy
ysathLsuj5x1/xrA3nIMjID/z1/G2mwrBSV6pp5hBdK9sRRztGJEYoXWvatu4Hx0YvWJfM1aUR/g
nITabf5KW2T753xjzEgMpZW4VV9fjqdMDGCok+JsWKfcpgE7VIzHb/3omY7dsjFk1CoCEtG9Q+h5
APhU5ZDa+8//MtHYe04/nCXMwscegDAEvxccmJ898YseNSIACXvH9MSe+npDfcjbjO3UGCsOIGsi
OR4nQCNUkxOXSxjFaEO/iWO4jGQRzptJotmtrgSRDhK8s9CpVomPfldGBLOX9cttcKwR6E8M8YLc
DhDkuQbkcpOsK6KWe/49c8b+5HUS5q4roUWyDIW24sfQKrX7mvRkn6ITrW81bYqKK8Gv4UQ3OtD+
p+Y7S09ejWppGIvRfpsgOV8GefAU3rBYyF3sAIFYbpWz7NHyAbxtXdv4NOSh7Io/gf2x8o3Dx2Rc
9IJkyimpXzkZfIkh++Pmx3Uk5nLMzXkxVSz2OwAS+AuwlNEL75t+rzbqjt2CHD0K/ZN0phVtrj1r
USvwTeOYeBBzKwqviEIKADXV58BhaniLPyGbXHC+GGHx8Dno5s3uYLQlTMfS5SLZBOpBw4XBfr+M
i4isL6rZacHhUCvcIkuCajq/7z30Kj6wUj4UYHbAFNbR4F4mcVsnhEOrCw1nhDkjW9y7nK84ZBUw
uDCkBSp9nFhNBBOXZpUN5PYXnzTBdS+RvQyGM+5LUzO4iap4pjpbaHkk+78tV7hP4BJgbmieCEWW
OxbBn5aXcwT8AeCw+KxpGv9R6MSy5wlRsa96569S+P1QkfRzzqQw/M/loQQAwN+ccGf7VSwX5yJR
oJ+UC1y41t0TDw9kmiwJzWNXCW6EUMUsgZJCkRRPt86ONmpByiLICxbMPnw8egdQNJxw61sc0u+l
k01s1i+53L2HteVez9tbzmGqUQ6NxLVlw8/Zy5SXKRAwY8Cfi1bebjMVQvPzoyZdaVi/CKGgzKT7
aJwtFC7FhoqEtvuiEVRj8WHD+nbxy1jCEuyurGDJoLJq5/nVeW6CoGaerXhZMwEDxLBICTSkfNky
ghE7IzHcEV62L/hFFVCMjNsjU9BasYVoECgTrsBi/bHTzr0Jo+yiDFxpX2UmKuh7Mryuccr4mSvB
3XU/EiuXwe3cR+jz2LFgDol7EIWnJp9GAkW5SbTp8bw1wwAV6MkD32MCBdhm8M9T4rc0sbviim62
gBZSyukpLOtza25H1koF3n+iNW32y+eW6NCpeQukm1CZ6MjsDHfP2LD7l0UV2SrGp+PzpBQyKOjS
Yu+QO8BKjy8FXwDxP1qH1j6WqSTnvwwLIq37LT34dT+v0zEQQ2TSsc++J2gTSL4Yj1M6yKoPa2HW
Lf2uByGLZm7eks8Qxic6011Ey9N7STMg+PWM1FyVCYjGSCIVR6nW7VUUMUGRLM/WhUenk2fhSOe/
7KUok/fuhUX63Aa6Yo8FCdh+gXItShN50t/ulnPo4Fz/9XdKuBHHpuxfI5c9Dp+qEgkXXzH2BSSn
Nvc7Z4QcO3uifjJU3/KEQRAdtm9BEnJVCCOqbaGggyFPZI4LqjzBywVVDiqtarQQttYQFhMZY8YZ
F9innCkK1wCmQE+MDDrek5b7we/fHHXZxB4sQqL+g0KV4vYk+rJwQKGjBz/pttZk0EQirVFITCEd
kXK7AUl/Oy2emIBk9JlS3IlwTrBWD9J+Gj9Igg5GuAMueDaqpKfNx7f7COXP2m4k+1qVGJB3Op8u
0D9+t2tRPQDmZSE0Eopjg4w2Lmisdve69J2iKgJBiiJyFYpgNpVeZf6qp/Kn8kAenLQpo/FHnEHZ
Z7nvJkTdfBKuFanX4alF8W3OjgfY8x5T5K0DzTh5ceIrMRXJcMIMgH1h2hltHyzj4d5kYsFHkFWl
XIcG6ABJJ3VVsAop5X13MK5AiTMAhPdEQAGHbysYWJxothMxLbsFi1UMDjBgbc5pk0VHcHrQkMjF
/YTozddZxlk42m6jQfbjDWpmHhNhUSijqJZCn5gbl8FH94LDUoO7Qw7pHL0wV11hURVKIBA01F1M
95ETkaMNqMctrXhsGrtjaiywVyZrDOs67FJjxC1FrgKVbRI4X60JrMPCPs3lo0uTSMVUjh08leqn
6CQSVzbiDE5KhfiFr/j3dd1TfpNmgmenjHDVmo83F9C5Jz27fm/aCeU/IkjwBuysvcsCU5F0JjUz
0t1pJZKjGYD7a9fnl1zAytewNSrjD/JPfQQxeDrW5or9yAkdkoY2FHnDJi1UlxXY8SRIAIoH9J3I
6mJ9BtXSHoMzbGvacdACgkBawnv6jxHbT2/19taRIbDRkiZZFo6PWZEOseYiSSwG3M3qVd5NtJth
MkrZNFyWhXPXTuH/yGwjg/MUHUtNMMVWa8JsbRsa5IxG64DN/e1k8J+31ExUQR7XCP+9xpfRZ804
JuD0meahc/M6qo2kTpr68pYlT7Y+OsQqR6ZFYyCSQew4QD4MZLtyclG6wsWv7iR+wWBitN7JNZMF
C2rBeYC9FJALLS7KtHi2ShhGczGwT7HWYmt36fWYsy4y4i4evNNwtPzYi5F/oJNHqH74HA1L+ky0
E0kgYJLXuqKSU7rRg4aDBDii6sKBnwk9OkiYVeQJfaL82gfQ6cWISaEiIkyN+38xz3qPV9heFQcX
7zhXHJIHnI39awbXEwp9nimIq0vVio9pYLA+hdkZ8Usa/uL8tzotyzLxkkT5SkXaebB3mBlBh052
XIWvxLU0kajJCvNZjEn7eoNp7k+QPpY1nzZTZxbDZd1Tzjp0EY+pxQXLV/lgiXHPoDk08hbABRiX
yS6gqqcgTl+0nltgEIanqkhC6nIZO1cVo86KFheQMqTOz19yqnSGNwrrxdeZdhVuu0sXyxnlt646
AxhVgMYwFVooz4rBo2KILccMp7UkSyn5LCungdnneadNBWu9euIGHeMqeD5un+Q/2HKuWjiFyqlE
CP74q9i0QmmgaYO64x4JBQ4Ww6MQvY2kc9HnBATNbVcaKwoGCPgm2IeMRiWN+QkL5emZkAhofeup
A9iMTlCTYFrazNY5a3PMr0JDgckMnM4lYyi/657pwT2EUROd3P8tZVuzxgnppsoKeommrGfZ6vc2
fBDkGITdPvliOExH47edv5xyl1Pqh8gUsJEUO623/LwJQ5PK5WqTNmzL2X+rP6yKdNCpq7Er/hZa
AwADdX3adwnw74DAU+wO7jP61wmFtEZVR61hnQ9+mpmE3dwKKDb0kaiH+8Nw1HBzB6RppMMtP3nD
5oN28r3AqRaAR7EdWENH3dLmw3uX1uxsJ9mF33M3505c+JUoV+ZKXjGJllrGBLS2alj5FlMQDl7c
gglwyQl4XaBE41nbLKpfbm+hWBMQeNs+7mMzj0M2tJ5vBWhfy6Zm9cl8qA14eE8kO/TSKsOsTQh5
an/CTzX1NaxxYnE4O77icODrZvk8qR00ijUBQZ+FznYOQBj/Y09PHiz7n+MBGPUX4RVmsS05R+0J
UXI1NYSwe+JUepukRw6r50JW8UgyCFLAaszEU8xKksCou9rkeHCwWy5hhtDoLLuDF3YZyACDlcje
nONjmTxcIuP8/tGqg76Tr4NRZL9Z9zWi/TmEnfdgz13NuVSYwYK8w6ODzhZCoeMcfCCqkSmgDEbt
rlsZm6+oyw+2aPCu8OFms21ffeo7VB+i91E7H2TcKigf/QyrwXUr8nOuk3p2rssj7CNMNzTcPXnl
8pmyHOVBvMHzXtY4B34GAjbnEGdQORejx96hfP00nDJVRPn3T8Wr7w1xt6ckfShE/PLSDpsj8dcD
U6jPEV2TDxiTdL7q0QI9yVeqfb14H8S9oHwtzMHalEz/TK+HqC5IMsuOzEYlAb5KMt6xjDmQlwU8
4NkGc6mul7HjKHNww/wYEvaqiiwgvcnUsSQJTpgGbN3hhmw2XNgFfjnq/kV8thY2jilwEExFGumi
dyaKsXd+Bo3hXcOdafp0xqrWzJJBu5IBXu+VrO9V8NTvkTJCpHPbYwyZusyjX4qxwKhYInwjpTfE
G0P2gFA2tJ1AXjYNl5A/ra9wZrJt8u6cmLmHEm+z2+OR4z++2SM65aVYexFXv26cR5BYv8nQpBcm
JUTRiWGpjHRRRhO9IW0V2mEe/2zj2YNx2sNe2lq/V0roMJPMC/A41faXjNxUNOGpY8iD74dgwyff
I4eAQVrxFN4wnXF1HsQvA3IFgK1Su0vB/b/mKE1Svy/n2L2hwUJsHfxZTmSMVKYQfzDED1nUabfl
ilr5EgW/SFWfjTNaBHmadRXlFdZQpM+qcRpa0vvFDgDzxt09A0qXY4+Fx+794Ts/YIjJ6DWPdQI6
89fuzVRjMBB2WazmIASPyX4uctwzqvMaUUAMe+R3ggVXIduHPrmgNBf2h7S2UWFlu6aDU5/+HlvN
0xdkVKQ0dNo3QE/FGbK/DLjuyLqUD8lmq86ZRkUe0DvzsDNUMHDuNTcg8CtsbIDIgxoOp5+puF08
VsExU9pJpZJyR+3T7tOP8rEBh/CjRqg7Ox/WA1QgdoQZ2oLN/TEuXfrJkv+0JJV/WygmyvldZ2Kl
V2cwi2CLEPJV5DV158fUHkXhf6+Gh6sYU0JQOOQdbbaavOhzNU3us6q6WG/jPyyx6oZ5HuTQaHWi
VoUusG3y+Lvxl/6q0HgGswuXnR1C4xJIMFRFE7PzIKeReV1nZunoaLlmmHDqyfQyjpqc0JNKXsuU
kJUx89A30fwbT3rdEaWZBoIhz05fwAYnsJqcOMxlAN31hZkSqq7ezAPGdELOUYHBl+67hmSDcUc2
LD6vvZMmFlMSmL6vd4BpDATemOKjTlwZ/QeAE9YMsbF0iD3b0A7A01+gqYhWpxnzjH3Fnaor6CsQ
sF8lXbnToC50NO8TN6+ev1p38P1AMirl6AJHyukXH3tLmHNOyNCv5rsJggIIk/4JobRjSfr61wfO
7ae5Fn6rhBvnrL7UHhX8OySE+Y1geBVgfGEqjykCEUeqB1PjIrCx4+HxoAwVMnJKXwWydwb6lHxv
lDbHGzDqiCfP1z8TlSfjgCQ5xQFboQudPvFFRb/TF1lEyUDL+Y1hg1CzVZcO6nYGmagL3Hhnc9I/
nQ5Rd9mHMj++GhpvFw1AJ8AcbN5rgvvik91r62T/KK97QH/nm4qYS4qTdtRTJy8IAPAVRULbO0b+
2MYR/4/BfLOUeFSmgUhhuFZYrtUGtqroSFvZp4EWnunu72dufg8srgsBkrMmGbnh1akwZxLKbF0e
8ZyC/gHtBGtrjlzD7MRZuraaZjd2kLsiJUJjV/XuHSMuzdTey2a2KCL9tcE7oNIwUUZ5pyebEGLr
9QCjgJ/Mv/xbfYsmJeeSmspvTSYiAmbRMQuM0uFX1mhlakD7YkQ+KcZT7+6P98I6kltEaw+K7wCD
MRPg3AuznecbttJwg6v3gZ/Ax72QY2RJO+4wJN+tDLsWG1YfJDaTk5Phzb9MgmDWQXGbuHJgHBir
UR2WTWsSyKfv20Ckv4eSdXYcisRDzLOAGv0WPm51ecrIa9fPC0Ugh/kx1U9ANSj/L4/hj5v1qDgx
78/xi64hjtb127TJ3IwO4k2Ke7lULC/ipRcAlWa5NCR2jmnFJmDCCAnVFuDapfqgCGq8Q1wmtdsn
g6mn2PIKL0JQ2jsUhNnfuL6StdmT50zFQbIhgfeDAKT/5d2oWJj0VO+/eAYyg2DHbTixtrnpxkF9
AjGXwoXNYo1dhWEhs/I9fyVrTekmyMu7vvwTfAKMzocHAKcHjivrj7wSx0Aaav6P+91Zfuog/zYK
qSBuVvINzhdvG2PUAGfZrqx8TLHb2IONcIgn7yIZM0FX1vQh6bLnGChL2+FviS5wtk/Ejsbjy/YR
/DKcsnrcZyeLOYLMymHF6azm4/CLbPcFy45fPkzQqjKixOltbZfBKrIsMckgjBiT9q/s2DUY+nLY
JzlxkBqgeYVv0TuDdpDu3yz5kXdMMPWuxV44AibM/RQrN+bP01j3G56HSSIlxzam3tUYMTrq5QeR
shADfo+o18/IG+UCB7aQMzNzNcwIqezFh5XuvqCPHojxRoWSx7aDayU6tHo+PFShgsWJSdeAsGuv
ypCqI8Z+orzzcHv5t2G96OFmomrEnFwGoUvoGvFowxc+BsY38tE2xCg3zqCzpH0SHFuTPbJyMzoQ
hEySwKbZIjJdafFL3cmiwnfFqEqJ1Antt2pNA/f3d9FjMj3lLiagx0gZ/vfxELrT0YAa9YdZGwx9
ahHvMdwNqmZATkfMVzwomfXyJNPfujC11Gmha2JDNFzxgsyx+zQgAUxFiA49jQkEtmltJFzdKx9q
5DJtZjk6Of6qQ8yzmaKZqLsbQ3kFOgMJOHx5VgGDQqoWQ85VCLONGZ9Ihxu12ccMlHzeIyuDe6Ya
Xcr/+s+qkEVaRIffw+W3yiLc+etccR3HyQG9harIomXfnF5b2BAIyLGUGNRogPnwB5vCvI4WJl0W
DAz+vOJx3IaQ607sG6JGCPVBzO/vT6jAIiFWwXpnJCxRyjX1Gh1VuH1W9Y4wxz6voC9S/NH/xQPp
rcGCxwvRkpvlYnTxADdYfsSun2r6nTmwrQ9fcnLE36Xnykf1ei45NTUSzpymJzWScZRIkKiF0WhU
RuxK/3evV/n94lqdViXcP/Obc2mGYcQn9o6n5BNU3Gt14EE2XabAoL57KBErlLriXGAvC+BpHiDb
TUl02RcGEcalPeNq7fAMzyANNdH0iNOlqy2FEZ7J+foio+72WEl5iDwFNP/W46a3T5BEAbrm7/DD
QiHlOdrDv15CnVw2iyq1Z+17/1EE+BFXMJBz9GoaAuXHevpyxhLrGzRLerknzgIs7hccpjXIrJ55
96kPl9+udwqWa6FZfFRV7bPKEbUmZg30GfNfmxYP8fQszXxDw+SaLWLXCMBojIGtt3rRWIF2ZVqs
OQe8j7P7Gr7jrUFEiTpVj8fw1WQzQQSpbpAWNrI9hq4dCjvIaUOhjDt5lyT62Y55ba3+H7U/NusL
fEiOivAt85YLFzTytXVWPsCwUpSrxaW+UH04uCuW4lD8xGDmat3zWi9Am7JuKNq9QAz/hjijJe0w
zDuESKOEBEXKL9qQ/9lvLFfYnE1t6O8QqAyEQpuIcm84p/5epBVVnqTrsong8Oj1/3XJ0X5PeCSF
+abx/UO8Xk5HUJyVIbmzzqT5JFdG/LC+AJZX0NOAUXmHTr9IBuUtZXIyIa74khQPSnhALjAz4smy
2Imcz2hXOGWsiL+63Jnvf9vvgSDNxi5W8j6lGH7hnTkKMd0lpmhH0mNqWGNocjLZ0furTcBUCDIx
GctkgG4YZvgqBG5JCUXZbNVh8ZtQSVdr41MpjYmCLuBzITl/lC87Tbpkwl/cEfozuyz1pibdDzro
CnnJ6bIKZJ3bhB3DqxPqvsBBDRV/jJhAFgivLgLVCtGXxw4+zPmpphLF4mvQa8hbODtSi8tmw71E
oMZCW6QGVG1Q/+82XDS/yVnJ3yvYWZJ2z9FYunx9BGn05ihsvsCOsDfHbQMe65IruISWN7GIXJc/
px0TSUmJZE4cZ4PtEuVd4cLKiyzuiBc6IDspjFat2QKPje2guWOYGYGAu5PqJ34ozEaC6w6pX2+f
LLiGgyEE2BEIqGqhWqf0PDqkNEYLr4iO4RwgMDoxauLjJL3cFkeVbDcyq3cq+pMqiHsCJIqDFGCi
06MDjvOh3XvFdzPiGIs7aG/MznqTiDcRZRJogw+qBuWAuqBawi3/gLaSHsNr3WA4zjBQY33QP4ed
WAlnmheqEOgAnDnzl0XNu1ClZoNkyn17AMKokIzz94VBmjWRbTDVjZcELoFl5Cxj1BvLAupnKreM
syaWzkwCPt3zdS4/mGA9v+niIKlgSHdqV+2xDtFaAYjhFyjK/9oEEfhaw2DtwM+qQAJwo2m5WLnc
WOCCiTnZlt0Z5xBEe/IPY0PzR4eQB/08NnxNkPwXoTD/2YxYwE4VMxeDY8BkDxa3MMv+1Tk0YwAX
yKqDOyl/6zLV2/If/2QCfHmJReadiUkdO49kDh19IpWQkGO+iYc+EgNo2vZxxPOvs93M0N/qozAY
5N/4d+ebGdhxggLIxSDp2Egsh3F8J1i7Hts8u6v26RnK27+p+6BS8divfVtqt2yyHNAjUZAZLTd1
IrFSzSo5cQbpvKS2Fmk/UAts89K7GRLxRRP+4LOJ7+hwh2nyz/+xs1jkg+tNiSextoUfr75TorTg
IS9rfapZqxzXBVg8wVsEXJPGSqeXsgcMirXsVeWL07qb7IG0xfzj9x/LHd87lP1GBaxNasQTkUtr
WjtiTU2Bm34t4xjr/g0SkV0uzdywOj4F8DhScDUa/g8JEA8WDK2sxiq/Xj/7w+jVamNFW6CGNbmO
mYKWtHuTpF329z9ATwbWzHnKsJxOaZhhCX5tWXdHrAUGJbN/trKPA7mPOc02dsXPUxb5A3IORRvG
JHfAH+t0CGjOi0NXdITUYDzZqGIFbiS470K9xcuDPut9Kna60gh/2bM/UPLJv3bjjWSW/u8jYXPJ
9ZMZdwQ55VfRxLgjfspsznbEt9tz8sOZd5KKM42/d//w5PuLWgQkac2W9IrrDAJG7w+omtHC1fEw
biOLarLTwWYjz0i9fqr/kKHGhTRU5rmhXiO9gbq+3fwd7/qf7odAKBho5V0jBpWUXq2zdMF3m++j
A0kwX0bnzo8jsAo9jq29lJsCvVsEiXTaXASAdwzshnkxjiziPmA9bP/FggUW5x66KqgHZjUis3uw
G2BzKKBf++GDAGHW2z7AQCT4pi6u1DS4bMwm972wUzPlS3tIC6pOPjwTwUDVw7KOXopTYvklQjOq
8kpn9Dyx68NLGCAVI9+uDZAALwu2nP1vL4CglT3dE7X+8JY5DWeR+M7y9tW9G+8tzjTwXFyq4KhI
7R4JETECIfBkUcZHxGr7ERP3kU6KWi64RR53vHLwkEqi34LdFU8dW/0AiaEEaq5iSUa4WOL1LpP0
l2dBrygb70GkVhvsA+CfqiWi+OI0LTuTP++MS1n4e8nJzD6wkAXrPFfbNk2B6v4jW5ZXuq9ksdpC
1LkzQ0GQ6soLtQE8Ao/4UgeNL5H+KMGgf6whh3SUR2q57kF4hyiG2SQf8ft9Y0OXIbmtYkNe9rsZ
J5XuZPjFRhWj3KVgfHYc4T6d4KVK1JvNVvcxd7aTFbV0JsT2EmPwHJEUKkX+Ztpf1GZ0GJa/b3/M
yuE673ELerFNiGOTV6iMxUHswJHkMzgc+fs/AMXcb+1zlrnOTEQgFSX1cGU/X5Sd2vxxaO+DUH60
QAtp8BRCu3iGmUNBHOCziYVs0YM7Pm3dA3fQ64+tiP86WTtbZiijsZI1pgoJGofqJGxbS0yvNmdT
iBmqFHajtAlKHyyQaZ3AXGjBnFTLGkOZe0/aNn4ugYW25fybUQcpPZQB+47Jl7+6leQVoUkltBis
1vG6GqgLrEcT01gailb7xZXK+tI7uO/HfpJbWETL0AEbWugVIYM1qaI4Qm7mcVO5hrHGXOTTqoqL
foj1qs9SPM8xxz6aClhy++/ZgE48UI4bxejZJlUelC/JRHH/TZ1eZg73ZOOHj+DrKAGfXgn1/fz4
mJ8hSHFRfBipFcGCmqdQFBcybAV9dWuhRVZUaRkCDKz8ui5qKlzYNTGlhmBgi7AvHiFfpBVNEupu
mXO1xZOM+9/5CCbqwgjmLkbA6ipNsc2ZS0t3N/VMpj3aMTqTJaAtAPVnwdWX8JUJqv7DkELA9wke
bc/gHXqEkRD7pRypAq4tkHkbZDGQTOOUtkx1HumKczEYpohpsXkfTA/ZmxDtjis0UfRMPnNuMfjF
X/izdNJ51aTQuld6xaRIKdCNg7/lURs4X3Fd0eKuBwkezfVO2C84z8G63YxhezZ+bPZe5hd4AV5w
2HR40wsLGQq19bL51Lm6IBtgHV8cmv+kl2dQfy4xZPpHhiEl17aEHLpWzj9xP6WBUPUay3DvemEV
5XU79qUpK7ENec4bwqy1NvVrRVRE13T459iPWW2Swi+eYmZmTdc+ZGTrvSN0x3sgdwp3dYPx9PCA
e4BKQth7wQ/Cb7Zgd7uaMiVqZHOIsVQxVvFKyZX3tQjMHjEQgpdTiQPBWdhXgAxcSSYwfvzn61QI
kW1JFxeCdGq7ABOcZwZ5zw+XYWF7kX+D6N6juUNVxh1TXRO16rxs2qotgabsN8Pra47Dp6YAkNxN
aKmg+u2cmjdrOokJ1tXWXdKb6lXRZ5f8ThdaqkDCz3xSRfIi1nGtRbLu0qZIIBb9VMYSkwFvS8Dz
5pJBuwxoy84OUsOz3i6ef2jR4u2Lluy99COKfDoq1NziMwza7fyyX71qQLKaei8RAEBt+gMNHo6c
35qgbGcB0mv7qN8xnvpks2U9uvXbxuvsdn7sY6HJRKCgLUI/Qm87aFKOp3uds6CthcaxhJ1WgyYj
FsG5QEO0fCK6UmzvgkuFzLcRyD4qs2NxdDb8mFMS8fAM9zs9OKEaHKjVTL39zJok2dBZxEJxp77n
Cn8PA+JuMLhtcOZjiXIL83YanL7bM27mQPtwJWkIzN2pUjhZeW6aJhxVm7pV0j0B42xjM8Mpdh5q
Ts7qXCN+JcLR9I2YCFiyZj4xEr1PA6+6IbjbZ5ggEZRUpXGGEmeafTyIUEdddqF681HleGjCKCXT
lZOD3H3cLQOV6AP1FNpwG4rk4C52+xJmL6HuQFQuQD3Qgu4vu16gKOPmnB02FhzvfzYNktSo5Vuy
6vnBQEDA98D2e7pnUIjlljrtAoDuSDUmNdQHrxQm4rRN5/C1+mqgbK7E60fP5Fna/VLSDsZHurAq
QWBQW05q+MkP2fBjsT3VFK5WAQVg5ZtfPkufnl33v82QV+EMDQhJoSCrNYNDmZgKHUU1H33putJG
43d3bGfM8Bk+Xy4G4LEiQfd/uJtc0TNofGkYCIE2gxv7t66QXk/pZxk+vmeGH3GdGheRHG/nEy0D
wiP2uW9GkKGRbJxaMrvJ/QgrfrBOMUOHuXFj7neHK5iJmn7Y+rq/Nq1VD2dc1dGToKXiQx6NFndL
s/Uw8P0OrataW2ye/zLaOM/sX17cMU1teADZA6oTGEE6t3ymW3kVVMFhM6lmquN/XkfmGis17iYC
DZd7dZpy54M6jmZG/MIfNG1cT1kXn6Y900M0Bv2D/gSRLjMVNNp1ufRy0/yn5FHsihm9yr/5diVo
4sVoHNM29irZeqmgDE6TB8O3OrHFpHxV1mMpiqb6xY6kM7YEML/dNIh34CGO/u0t52hQNnc5ZKox
gPJMJPomP33c4svUTqnvStJEYgOHJ7GLrW1IAksIR1VoDQXSk81yWgaHFxGucQrtCpT84zlFBHyt
iYEk5zlA0BuGfOBKTCInwr2IPky1tI+hkgWGPL4ihZX7oxwngLp5uj64sVzj4RF/JFIFijjBGR00
eVcKJaQ3Yp0qawXrE7H+dKsSZcoGQm9K61sxcF2BOHZnZ5jyuz9NoJ39B5jGy+Dq9i88jwD7NrUw
JRIaq+li+7utWF3tSLq79+BLRHKANrg40ioJMGNqSJHLEgndDC2GIe7YSGCoWJaBCDmsvjddtHPK
tTmvsbrqdeYxFJWe7m889X4ZOzO8TiT9l0zbmauz6ct40ReGOXU7d/uvgvV3uYZ8k8KSZRmiHUe/
3gDWvE4iusBJptz8zxgpBlp6PObuZMmrqq0WAfwoFqCNNveYzlJAFnox7ZnHYlCfP6tXPgHxhHlL
UA3tk8bNjUU3ZCtZfgkjAXidbLOKFqH/IDtIqUE6myeW7gty6vf04y3IKW9pDarxpTrXAUzO9GcT
FR7ln8L0yWVjOCwQqVDM5i1dVlIrVyqSVArlCC6+OKYqvOsyMCD+xckItdcSKzKf6UXeJ1H0e7ZC
ZKdBPWw20chlqcSAYBb0uu56ZKg/FA5ThUNsnKAfuLW51zXYmbOM/X5avKJDDX2vfdClwrOJX6zU
3LSYo8loANR8u9exVxO927xujdfQ3UixDwE1v7wd//dUdRakJSzfuh8l1mtn94oA8gzblUNQi7wv
1lV69s7dXu28G0fs6tg9y2o+7nX84rcy2ifnXg0XiT3gVtOcY9eorF37N5/PW9kPnfGygoUPBEo/
WquRA3/uX4ozXOXxhpZP+HCCwev3jAZBmiJtpwWpnZYkciZ3kjm5s3F5/ySttLKIbPIO82BR5jJh
x6C27E6rGt72oDJLtmzMNyXr2F1lab5h+NhYTzieo2zYBYM6tAlub/vSwFJ8n3+lXEFKtP/wPs6V
moMNlhyMOfWqkn/Jljt6cx3q85DsWALluPOhP09ZlouOIe2LvHKD53qEc4di8IW1YGv+TD+oq5/B
CiYQSN8sWA6saPLF3WzgpXqBYNdIgYVjhRmuCGSUl/dwFf1RE0Hhei9Kvjnz+pwt1nTk+pQbu+iG
VYmCFUwMdC8IHwllC/+lQtI6JEJXYDYKKPmLcjOByJ2k2Mwg9NhKg4L/2R9hLQaI0bvHYKNSbtPc
LlWCPMBPnFfwrryVFsJKk/6sQylHrNEX2e1V7DFAmxha2RrtEsru2hXXz0DP+iuggW3LzeuL6xIK
mQq3SlUwOLjtiHf9By0G3XbgRruAGBRf0RXGbFo272aQ4/Ry+NLn46kxs6fWcwhLu4JLHikQV81y
e/HddaBkC5DSeyLJCllchZrPPiYlT59L9ZlU3hrFVV43Qej3qRbncJhMUdsMFzKipxIIMIXAGyUa
12ItSp+3Rfe0HPsjqM/PzORGrY6F+/OxCI81FaXCUhKz6oskZFmhsBRDRjG8TGvEP4kIfexP7yZj
9A+3GQJV4ci1QPkJULCl6QtFUi9ESQaJf82xrbaHf8pHZh3xGoSWtUvoy6aJVfUlOVBcwXKbNaZx
J+raBd2+Hht6pclxBC+Z/GAVlwfUZ6QJrqjNuJgqdaovUij5vknCLAjaE1SEk+gYR5qS7qy4vTe5
Nsf1eQxsZp32cph8LrrIxqu5PeJB0O8KryDwToPCJeockrikTpFu4qtx3rASlP4zjOeFXLB8rs5/
N5C2Q6YJqF0OFwIyDeNrg225RfyQfakWJpPE31YkEeR9nXumwMq9BRSeV2obt98F55vuS3TzptZO
e+sZWkBYDUGJdBjCTlw5WB2HZttMbJd6Yd37SnakpF0V9gCLOLiC6kGulsDPntrGSXdscAx+A94A
LbgZTCjtDCntnzBwZu92mypv7UGQG35BVf04xQrWufJ/xJrvNQSkJa7cqqII0u5ePrnuUjQIg8bd
LEA+U/sop1lc/cejRaEzdVivwAhWELmSO18I5WlJf9npT6ICdeYt1+GJexgo0stANhTaisLNy60/
BJByfOmnBpA2qhNmtJ5CqNoI1rEVSgbR9KezDgROBzs4o/41sAAQUyvKKRUrujLr2h+H7QPRWkqj
FA+jRPBQmFdazX0ZpmGKSI/u3dqwpNYRfBC2MdqjaoIZDm9ZeAHTgIqtTZdU3ini2poO0j/MYw4x
L8Lss3OHcuqta4vBmeK0I1Jr9c+FidFFZp8cUa9EcojtibLZHQxhCJROvDocLnQqVu8LSYVOLLhL
8loYtuXzsM8k9YBdSH803WTB/EI+4HXu1rShscJy+jk27oFAFi+1h3eKSk7Bm2Ddh1mGJ47xvUFl
WTVZfrDl6XOQR4cpFEpYjyKs19PkQuTSj9P+O5yG4oqvx9NSJ6ZCG+BzcaBv8QV9dJ3wKfEE7yf9
Tk82LYK3tEyWtH5Rq5f82molw7tK3AXPQN9/dwXFqVRsjq+Rz1i/u7LjQTiwwlMMBqTFm8NWToCA
qExEdBLVbGr7Jp589blqUY1JB7LP7Z5wXuUQZZzDh+7ObkcBkd4l0KMcU6oxyPf2TQtkxxQxlUWN
Mf1REpzldsKs/F1/50BwIIYvNkQlxCO8aB6opZsvxbCcdekh9FqYRrItUwf4w16LUs0j6QUwRaSY
atAKNnBHww4u5Sc/inJS6jGYTMBAticjZUiZD8RKHv6WGFi+yL0z6HltSeudtwGD6G1kFyErB4/g
NTb9Iqa3r1lpcYVZgFwUq2lmWjEebAe0TPwHxJglG8CYxq72fQ3K9vrXL70NKMKLtveoZxiOlZPz
aAwLCCxGSTnGgVTIh+FymuBKZKKqMXSAu3/hqUEvKPhKY5yXWP7IoC+AtCWlxge9uTKKFaACcXOa
bKHXYYXTJwLgmh5OuqxEYOfh4GCbh+Lhe2jSk1c7CpSSI3mRoMSpp62R4KK52J7Bpu1hlFIp6lRr
nQh9k5r7CkKqepyagOfPeA3HPu5z2yvRVz3rB5K3xQkVfOxVKAO6N7ndJaUVOKKybXPudXKoB63j
j6InzX+XBbRMSXlSCu8oUEvdfljSQGDlNC5UPayrB5YVFdw3pBFJBjsNDTSXca0ymCUbOeLe5ww2
Y+X3vCAR2xCae8KSdnKkYYcwY7V0wnAKr2ykQ65QLjGZwSsIhzA1sXgrPyeJ3xr5rLL4vkwCDHy8
REwm27MJobrFTpNX5Y/t9CYAtl2KKqxTlosjrRV5LLncyHcxXBItmGMvUSsd/pYisrc1mi4F/wVY
yBap7BZe4Aag/ysSxdn3n40Wn8ay19odrlzKQZ2mvmou9Ui/hj0PUktCOmzb0KRGiOu2yCO4O8Y9
ydU8kd8jRIWGwst4N88VTWLV0N/j+5x+jQzsei8mpVd/dxYbj13b8xE4uy7Dtqwac2g5Iz3OwbvA
jDPRrm+IncjVUdX0bTt72lE4pzPpL2/Gk7XKYXFwz4p4qfgo3Ee/eEkVWPBfkfsOkQyKTiOUtqS7
YSHzn/5y1CazDa7l4fzw8rRdu1vb5FQFaMMC2Zt3mUu2hvxTM/3rZjS98sqy+g0lkZlALaoYOemu
JE73Cwh2ajlWQjPdnyTzfQDhfwVnfhKAA6MzjogpQCsN/dj0OYZtg41euWBqsET2Amem8tlOCwg8
HvPK+zJj8v/Ly/Am3kXP+ztecUvooTC/aSDZrqcBVHrc6XzclC3kgyk2wFtcUz3283HTnj8dYAEt
lNZMr38VWlYApfMjlJDQdzD+i7kz3XlSBnGsRGARl0LXvFcvpzwBfePyJCg1JzQU4ESWAlE8uAe8
zJlIeYrCe3H2yQ4J5LZNFnfn0HgsfmArFbKJiTTZJGURK7K6r7JV4D+xT6Cd5gEfFVltgtLuC794
DEgsHdOVEtsQADA113mUGkHqkzwJvNuuBLgCTpBK6qk1eHUPHGR4wjjotBiOMWa1BxMQ6XSZOxAk
snApezngHLnKx/C8/tjL0rJu6m2Mme/0/oebWgLftG7D59APFaJtIDZ8Y3fdd3LZMjruzCfUM3/i
tp29FwotbomEiU6TqIsq1idmH+DqCWc7cyXpdUHy4j7ysMxJFq+AleXCoRT9VXS5LwmL04G19+UX
ECodCeYZpScUEW4AkWmc7+33TwY8kfO12vCocez3vuNeY4uFeXc1TQ3pnqlqNwYOJ5qz6lE+PVEB
C4zEcr1SmoIMcQEsiHLMMO5CqXk67wVhh/xUzonfY250yFHQfvkrZ3q93WBZoahc8g8/p/pRTFT6
WC/kk7Rt/yHYYKCx20HH7swzoeTF4lWBealVUP8t5E9xRuIM+/Q+LsneeQwjJIcxAnRDrbX+AeCy
yIDR11CbZKtdMTGfYTXd+JNLs4GzSr/HndpvZOdyPqbbyYOWCe1xUCDMa5nmSCXNsfzFdTDL56yQ
9WmEJ0/JYrbJRPWNh9DBbe+dgTnJILhAiLkhptov5q5FmWrTud2xinAQrWfys8ThWhhjhzurxnAD
o1LXWUeJ3NYAgJXJvhu/iVM1G/102aMNMkQWLg0Q8XXd3MdRaTVNHgBB85/BphbtGCBBpC+0ifk0
muAngMzIfk+/cWWfcnSULEFAYlll6s/4q+pJGla1/mBP/3mR9xNxooA9vPxsQhkZJnLKmxohrF+l
aMGFZFd3JEmGcMxwsFD79Cy6onVk5l7Szwu0AFLq+BFenA/SXVl99SFrDdhDSiuNeKVDWboaextX
oSpNZtJ31WjdGu0Wvv59q/RsPvFauuptJ9Vq9zf33C9LFLvp7tuBJWocyoFa8uBnLm9nx0oFPxeK
Vy1x7aEG7JXGBNhtNglBWsZfx91gkidjnYxyUHViCwr07m+ea8U8FKGDNLzdCEcMFO1WfdABOiFi
cfPbYXvsQ9HqpMzF2X6KQg15MAMU/t3qM+Mu/hGKvlmupVtkIcIKAAny+pTdCUJpW54QXL0iC4P1
zTirL+bqaxN8Adm1ySpUKoM9SyMI6kP1+iESLkH+mbNncBUeEoRO8HftR4ZafEKJkSRh3lA+xMSQ
uI3647mmroNkiA5Y/uEixfX6iRbYGCnb8gTQIOml42IMJa2uoTqUr2wvTCZQa9NWRAUTefof/nui
9nDcCEZw9GvQL0HmoSxR7GsG3AOjWdCTTynhQ+s8SffuFegk1+9GOPIcqxSYGschElzFbSJvixOx
60iVTyz+ci8+rzjoO96Tq51v4szvFPY6/r0jM9bKJWcsyGGOaHp5f1jsJvewZPVFPnJ3HHDUJKq3
03fu3A4Pw4uQkOa1P1pLmk46Ez1NYWXOJDdb0Vl2Rv83dZBNMAbbVX4tnxBBWyAKKI9wOEjwE8C0
nO/ZLHwLdozCDBXKlulckwAEJ9UWXB4lbJrkriv9gWy4jSmxPrAaFi99Po2L/dtQbh0EISQXPaGQ
/pdvxdKzvQmFM1pUVTDARCE6NRu0ziRDb18ka9Qg41S0XfykTGq45z4tB1+74KR/zPEI+LZXOY3W
tRDBarZnR62ZVjuOQQVw3Le5oW4szKMWY12kFNkdUd696iy/+7YTn3SXZKn0ERwHSgYgct1pb9RZ
71L4zGgMHx5e9zx424bLUww3MhGsftJWV0pcMUYO6CVvd6TiBUYd6TI8dFC935s1wg0wzZRkCZ5u
D5I2vB9X7qXuSsch8hZM4fBP4IKwidA7kkk8S5Y+PvV2bUJkHEZuXvuPuzMEa9alp1U7XcCPVAmH
bAZb0DTAPB9Mb5JFJSDcaTQewcDGrPYzvOcJ18pP++/ZahjoUd/oM8TUWgoCmA/NXkQhTebPCT9W
VkABv4pMWKMORGXoajVuCWzPHi8G0SfWdy/Z3sYC0p3Dp0bQD9IWudU+ujwwe41ovLVDOs4FeB3C
FSJbYSqS7LFXhYIXdw7oSAlBXYu/vjCNC2qVBOuW+P5+Qn4sJ5pqdNuP1RV6wkEd9gN4sxGcnKzu
0O6JSZ2jG2bYt02Pf+Xn7O6CbJY/KHwLDU91oARgV1hWQVuSsOQMXDYRmyAtvwYUzwuRSr0QXz9B
lZWPJDZGIHBsZpzaf/ZY6fOiDy7QlNzG+kLCl9JhEywnwtu/f62g8/m0A7zueexmBiDrBDsiJGsH
8cZ6fbtiKvc+3iRfvFZHFvvXJyNa4Jt1Kt8D+8Wdd6TbYcA54ZfoHsTZfmxV6tokV1rz/P5pwZv9
ni3I+iRZZBk2Mqp/dmvjwmRsgjgxtAEbsH5kCydfDMhCy+pz+SAREz3uUf1vFOklR9z/iwVcGE12
QNM9i179qujLg6IjLn2cWC3rybuV9jE2ALM1W10tG8UDgKIBjNgrav0+vb1GSgLCIa2GE9HLQYuS
tTyhbJ1awj481J9PK3ueSpksXByEwxO8UcczXPTFt2Af5L7Ai5e+ChzB/NZLiw2j+fZ/VlF2TLBT
h3wtdbVm3sIthkPR0YLlnxyANqroCk+fwfjEzgEGafYmaA0lWycU5AgZzwLbiHlmoKN90C9Z0nQG
oJZES4dq1mva+DOILwgIqMA5HGmrSFSeTFPDovhIuOWSWPZDW7BBYh41+VtosJAE+oqdBksM94cu
PKUZCh/kHamqScd3Pfa22E5G9kSCdjnn4BPliKiDqnjUfoAaabzKYnu3qmsu2xpj/frgFC4uIuZM
/MHiAao9SioumV0EmNA5RJP4VsV8wGEyWuZ9qD4ch1sWx2Kt40P4lZ0Y4uMD62PCpwO3Rm2eFJOP
hthtrMqlOiQHbqiZP/gpcEHKZgGEnrkPbJysgr/gDL7BdYdWxSlE5S8WGGArykT3TSKE4n/cXPRF
veULKDfSaa1gZyElNAy+m21jsDaFBcUugBl6GnFrgLtgXcPehjYPphoa+VRwPmRvJ9rDebPJKj6V
vXtL1HR85PTobogCl8IotUcJgEdf5CF7JqSMoAmltmud/qpzjDwDcOilQbcEzJvEnRALqYDkOrZy
7bEIJRodlwamAe6cEtoG6muorFJf1Qi5S9jroa5ICSRHXIDcG4v1zpgqtNP60L6F4ROpBehAp53K
gOa6U4o/cK59qRyG5xPrrxomtmJqf8T2qupCIC/5VYpHpoemgPYK2W41+/unFoHajNUfBWzl0dIW
DC8kWihHQTPngCy7nHEsS6B1IDj1/y53aUHQxJR4fvC3e824f0pwGCFpJ0XSdK7vICb5fhjn0R1B
d2QFIo+frahVR++9mYGc0QenmH73M5aUBTsnFtIrwM8M0JomqBowK1lTOVzAmG8yJ84W4znzZWJt
9Q13QA+I4NIxclN1733t20XREScGHJKYmDVg7Yi1wrRMQwkQxEOjehbycXc+hAI7HdYjLcpfjR7v
6fxiCL3AKxdrc39ESm6kYt/YuRLSVGASUU3kXEN47wLXM7co+FhaIGxtml00M90uX0wN5LvbqhK1
Q0aWFBa2tFa5VGr0dosbEl+Uhp75MnQIXfnHnO5IrimLEkLq5QN4FKmqxclUs51D0VYOkTjoQZqZ
j4lUveaxm489Ok4nHMxfsosmBkyp9s3bKssw1fiURpoTswrr/3wMk228N9n4amTKb+nKb+5V5HFH
nk1agkuD3pFsLEYzQtWMrBAXBjIaDvHYiHrOvWWkiNRwa3iNG6SgMXrSTXX6n3twTrhkM04V14jN
txqXAxI3ucMnsRjGux/xy2kmsGa2dd/6RU87SA9DFdbuz+h1wgjgutGIuctVn9tkZSpBujsCG2of
j998K2b9KAbrEl6T2QBVl5yJy2jhFHk0rwOEgqeMxhcGrmXiPt/ofkg1mfldzdoOcqaubZbWnNl7
G9T+s06AZqu/XgO91zOsxHutYqPTV5uXXENwDal20UqPM/m3fSmg08AhFLQuNFTAVFFhVfKMy+cD
HrivnhgoKO5bkdaKdGRvkToJ4R7PMBVMxv7FJY4IABaBISU7hhPVZ9IR2l8ORBRUDndSJ6OH4OTY
T6om1Vn0oG3/Gajr4KaoIVZq5mH1ByNU7lrRiwSkVWwE1/9e11YwivRyBClTsViAZbEP2UgnC5rl
7pAoz+95mNn8ZtK00mQS+TWx9yV00J1hmEI0qLjzMWf69NJu0wxRP0ddJSLmlPuh+1HECedxlRk0
khiG2JW+xCVmjKPyBlt6a5U0X4nU2jZTtspHaaYpem3JhV5/N79gQYlTqAUo8gsvJrFfuGaMWBKD
Pk7qrP7wNd6V9+5/R2wqj+uqvouJr5oic8NUHcAbB5i9gQQTGwhkDdnR8O6kYNmLMehcduLPiVzR
wWBNYEp+AoQqX7ZHzLPWD5gqDBgq/6N36FgTCZ2Ed/bjuq0ABDe9/vn3UAPChdh+5Ha47KsG/jDR
6zWxwa1rV6YiYvP9HZ5eHO2JxB1LSZcvAfBCGSkXqW8Icu5H02Nky3bXxS0kHXyKeRCKVEGtC+Aj
ExXtu32aglHR0bzAJlx9taEXEV3+MYOrvK1qTNQ9cnDvRWDaWzlx3r5mfZl1sKK7V/dvBwSX1dBz
g/h2QIPcO8RnRY3fub/2QIF/azuZ3YavwJ6vYWN7h30aLtVwBViaOCxoaGPijxk0vyeGu6re1Knf
Bv2hWEEDAry5zZO4x0RbRNGlrMk3f0FlkRyIW3mP8aFrVtawTGwO15mREAtVzkcLnuTTQhRhonwq
S/sKFHIhnx63/hNAhCkKtjDnTAHTqmO9n5tpAhn8VOiAVoRDilvm5Hk139AllDzdmUYNbVrw60J8
N+3ousoEt6y30kz/C6SXxFUw/inwkegn9KRcYr/MO6el8ktpIVsvOZIR+6djwLG9G8VkQP+G7FNT
XgSneuWRcjT4E3Xi9vViD4jz767BwFBYdCF1syNzdr2DhmqG6o7XX/c0FKm+yL/IIJvoctm0eqZd
trLLqAGuL1rjaH31DhHjbwWYX0yVOrLsXNnwjo0OaAgWUdnnJlh45FV2GyXl5qPWSWYm8b/N7Mu+
Vb4eFubJRomCOP6Q8odkfFKotLkwp5gw/rRZ8IhA/Mz5CJ6Sj2pIl7TGenRmwXgVS2D4rfy6Q25m
6XUG4DgGeaHv/mgqf2eV4b4OiuW/Vscgzn7NWSpCLI99vAATmzOHyg9iouX1EANfiXGrsRsMmE2h
8t0U7MLe+XutubS1+I4J0eqO7yEJpE7OGxb1l8e0gCv0EpOjJR4Uhi8hML6X7Voa+DkwURi6/B8W
TJtD+n7mQnSFTC+qpyUeF2SRaBAbiVSPcwBT2h6ff9Jf1dGrbuUwOBtAU1LG0fXiWhsdFBGQXKIc
QFA22IY+KsDTe9IAdw40omwaqk7tQh1T8eR/mnIzCsNFCj2Tb/vOsweAwT8bcX9xUvFDSv9RE2y3
WAy4f9DhK8EE343PMeicBHAsqz8bt9vMknL4nl3RpOZoqNVbFKi6WDS9k3CHi0XNyOPathauRSEg
e+eNANTRvfUVQ74SewEZznaaqe9xfVTDbXo1SHT5x5dqU3qhzdeQEVlzZyZTbvWz1H0bL02Q8xsP
5B1KFfXBl/foeHQu5zvTZjxVKRkamYvXB90F5HybGhbuW+nEhRiYv8ojfudWK13g8BDbK0xzuhwC
Wna4rLgSkNL8WTZWV/WDtOwOgYJpbjZRprIvfXV8cQ54bw45G9wF/leIy2YU+kyyQCpU7RJ4o7eD
pe+1uwt+tfjgb2iKKKVQXXSl3F8RyE1K3zhEICHCQTxLgOnz+DYtEZ71FnRnEsr74XWBN/tq4imr
1YwJlOtO1XeaW5fI93pEjKQj9tuYAEWPhHhseQCATTHEcqIfXyoVEjwIOX0eGjdYEfi7hI1NpTzg
NApZEqERD04MkItVQmJOPxXWXse3IO7G9fFBZL2mgtbVCw3ufgdBG71/sHjeiduupnXqqRBp5pNV
zoF5WjOs4qxZMDBepIZfRrr412rCD8yFNcJFOkyTuxsb0UWg03BMd8KVh9N+zjhW9AlUtfnERmfT
QQCdefrEfB/hIFWkN81cHv3gPOGjjLm7JKbY0qbSQ6hQ8ew8xMVz4VVSsW3Nb44ZUQ7M8jKjg/Js
Y6tUdAgVuuCFTpHWWM+YI+3x1zwJ5WJVVG39A/IhpfzL7qTtaNtvHRdZsiVdZydW+BUJwJ7Nsw3G
0h1A+TGyk9s7ZXzClLdg3B7HW4H31fivufF3sJaM7W0AOfMj5358wxwsBlThZDEAXFG5+D4e97F5
GZutm9p4Z4lxCqce58WXtdjUKYHeEMS3F2j0g2XPtqceUaqH8pz6TMtOUbX90hgtBkSP0o7Y9yp7
aPYO6bPqxaMqArvWbXidRP0gX85ooxa29cJf7ixqSSUfWc17zwp28BM5Oex5w2C+mag406qQroNw
TpRyNl5ypb2OFk95jJHaagfKbDX9KmHKdv83yPh3qivuHZI0p5IEb54GXouWulNhS4L0OPK2yiWZ
9Uvh/Hw+8Cs0KeWNcZc+AlOn7j5r0HQkrjWck1/9S4WLETCCBDdbrLvzzuOqzGQVTE8xxzq+BDYD
uyEtV6AFoV4xcn4hMe5wC50xajL2bo9/3x6h9dgbi3B2F5sBpZ2ink59CEqH4RaYA7DMIGYEiSGz
oe+6fFFHVvN3jLbgM41bZSECvBCa4zaIbv+Su/wZ0ExSsxNVY/t6l3W1mOtrDGqfdICWaHZEn124
3TnUjZ76OoxZuoQ0dIJ2ALr2tzhMnV69XCSe7lQQwn+n/BiD1G1nU0cheQnyK6vKZQkPnXtFq/Ip
AgBpORgpgs6Mn8ExFE0fE1wjJ3wQovRZGLTMMqrZr9Xe6lL7PtpiCazGD1utAgH5zUdydMANo4MJ
u4hlbfeYvrnbvdtCPnCL6IuUsDcI/8py/BP2aGht5YNe5py4D/UcpJFe2V2vFS6oXpBrgF4VFZN9
76JT1EylADt6ApnhjI9BVYXdkztiXBLXfP63ldB4xK+BQiOlitEmd+exnLDNz5vaA+Qt4wFWNHz1
lZQzFBN8a8pRrw6QlQCzytGkVFHoc78nrb75AA5QF66iBtRAkSpasAyUw1hi+zkgFkqDi++uWQi/
r/Du8DwVay9GYlHv18UlLZjBRgAJ9TaoB7tJtFiEIl9CvbE37XHpF8IbEoPRlmxrFU3K6EBOfz1q
5VT2x2CPMcqMJzClvDarOJHF+fwAqALyVrSZiBFHZDXjTIJPOZoDPcGJo86jNZ2VOPARrN+rWy5N
TIg94VlPV9xqmcvJRm4buon6wriH5fsxgyFK3u799mwvJi2vDpOOIQ4GdUp6auPUI7shqnJ5bBSe
JcOTCSBRwpsqYblF3dOqXogZYt02icPqK+UVL1Z/SLAqnzD+rXpjY95LEHgajhnJu9XEQ+KFVzfL
vrQ4C8w5aAtmhtq3PqlXwDEUvlLVcBUdfmJgnmkUiLqkB3DbYkAw40ci7GzXyVPgwg2LxnVjqD53
02hno9WumRrKXAG9opEH9BCcd/BGzzvYEUKkbCwoJiHf8lvwPFi5brV0vrbN+e9V9hlVtNeiBj3R
naZxDh7C7AV5xqKDpuiGJfUgveTV8jYDy5c2mGQ1QWaE+nUiGpEQ1lWG+1HyS/KnzEyQLc/9Jch4
ws0+kvkX9I+OoX+JvtqXXRpopNlJkYubHJa323rvuZKb8rJRkz7cuYGtQfvq99Js5q/RU80/W3zH
nK2zpLcIZV/C1Vr47tCRUfOo4blX1aHos8/6Lk4zeygZ+oer6c7poDkPSwGCzGmzrcaLxw6wF466
gVGTuuwgsjiven46mtDEThXSpFdmnqblflZQbWWENaTjMDIZJfS0TkWhd/bdEtt0k2mFDInSbXfq
eMnSjqcKX5m9mLh4ultgSdge2TYyasvhe+kIvcH/CHEMjoZ50SGS4sSlVYNFBwiKsCcuhNI/4kHX
KqWfTqmdK/WL/+fWcduJLdaoPRiqSEfbxZgdUfGMe8WgEXUaTdlY/ul+0A0Df9I2Gwz3ydMq376e
v/6eXUo0b4XXh8gO5Pjj/sE9QL++h9q7B0TCGbHrGMKGJcXiFUf8uUcBnItrfTO+KEKD2MF/K96m
lvZGZ9m9An4mlDzkDK8LFCS3TLtA6PZPH00vGxkB86H3DsdvkLOosBqxqmtUFS7kFvmS6WbF56MY
ZpRUvoiTA50DUiFNMmOWLhpiqpqTjkv5LKY6BL2L6Ge+DHNN8IS9DPFkxZjgO58QYIeYRRJ/z8n+
BCfPjE7NJkuVyGnGErX/GvflZ+Q4bC6AdMzU0EQXnqdg14ZjZva4eKICni2WPxR8lfx01p4aa7cU
8EhFbDKyI3AYSbml/mVLoMSJJy53n0KVWrIXGziWL/IyMOpnfqcGBL9BD715fNP/aG9Zga0YxNtZ
DjFOhGe45bgk3I5iY+4+meXNKd4Vz5EiktDx7EzLsxNJ6Xm8T+/fPPj3cYDvfJNmOLd3Vv0sMlsp
I64P7XAflFV2DAx/IrIPJTAq8XMnpvIF9BU0VJqD1J9mwlbSK4LCFJVgr4bBW7WdmKs+87ksGY1Y
TdnjiPVs11D8IhBFwfwlRUmN5KMifK6cGT+bfC2hYYl2TZQdUGNUNm6wJ+entiUb1jmoyEacq4nh
i6eUXU2AUMkbw1wdMrGwiO0C5CU8hacRO0NjGHzv5x+eY4AE/qxUkajGLOzWGnR6VopKpJYSIsum
vY+ahhZyLzUNnMTHRrf5efdQPqLJcNimwooSn3CAe7KqapPzqWICz9/bsIka6APL/BAoq6UNbQ1x
ZnibmZ+b74DC7+UyMKJulf0N2Ogd5B53iwf1HnYB2qBjZuEzZkGPvtLknF8Dd7BsiMoae+AP1rZe
BKEUnbt5E+PJZp+1UR/qASLTUmm2layCrVxqenv2TanjYmgPS1LrPBSIZ8fyDB3mmA1knC6h/9uJ
YdEPIjGb6FQI5JtoQ5i2Oy9DNl0v16aQLAwTm6PN9oL0UPJlhs7KWJdKXyVSvKaPd8RINPF6aYHx
gxKoA1RSOYTRCvI3M2irborDMPKQYrDJACPcB+eHk9UUVepqYhWH69/yYa7hCnKiEsagIh0eB2dR
N6xWjrpPRGMKMbeBUK/T5g+/P8ingqM1HeXSkUYAQQCT9vutS0Uh4a0O/IvENP+iNiYd1t63uznn
eg9/lun6O2nxrCb7Qe5F+RPhTq43F6AWndMfvFRNYI+zCToLgaXfIpATLxYMjsUcexKUQyv1h+aQ
rjw18a1csch0hi/q9/VAZ4knOD6K95zyAVCjO3lYLB1CEn27vc9ScQM9az3IxPctAF07eiD3xJLB
IGpDdM2R0u6FHPmo4j3HzpHwwY143IhME5WyCzDoeWQ1iBBSVeXRixtLsq8effa2hFUyF/lHU10/
34htiOnnLMdi39cMVdQWZsF50/K6qLJUclzVkEXeU1a5940UsrK0BxmgsIGIFh+axYQUOe0O5mRo
lIG2p4Xn0gvddLZbHZcFqj8l3UXaG6dgAcQNrh3/5d8QeEjfY2nGv5XPsT6WJVpiP6Ij6FTYxnTb
9xZooyQj5TFTCi4sxgOtgPK7h1NopPpXMWvofxCTMHTAlRYEh70jxnPs4x7FedQoHp/7qm3Hh1P+
470np6FCYxZQrD8gNg450ipbUPW/f2zp7Ue0dMtrmdVOomLX/vZvvbOfs08xJHdEPfctrYLqaImv
7si1tUn2UdoxkuQu445cEFDFMD9ZRChhAFGYz01Y8MNAtGB5Xu+oFdCjqFDva2bqjAhdv8okz3jG
mt33McFmOajkxVQS1m/A4gStcYqH14W7VYHDnGxuk9WETjYMLlvMgM/2DpKjmbja4PbPerHE5qZ1
4EwQNyJG9+aK+4/md2zkCJiYDnG2M+VybkBeMCFU7m8WTMNOFXC7FVQb1PATC48XNWTjunbSM4ho
HZYamWYa0AFm5yXV8igRm88jo6eWUog3Nkw6xt/M+mT2Pi1b567dbWnu4c0yhX79JMBJfU+DTRR9
a0tz+SoluAtSPQlYdQ+1dSb+q+tS6bnVGG/lXoGusVQKp1PydnJNVAoFTHLCuZQbvlOCip26xeI5
jja+iAlD7umgsbL5P3c7f1LAKA74JM4YDHGFc4BffdSyUmeGQoDVRdecORvZd7xxsY3vYbjjXN0W
qOYhYVSjQ6W1+LQrMtv1inySUIxQuK+lHkQnf/dh345Yzc6/A2qmZK+xIAoXyQUCCvagsBDBhtnH
+fPH+bH1VGIH3zQtQAPGLuK+UiGPgk5dIx3bnQ+wLC2c8EO5bLTg7aZGhMJJZoMtFj+ket5qKRwE
5ceaoU2xEB1RMPB8qHeQcaDmHcpeOwif+lmO633eHT4wPvLL/fzFqh0hK17h9osvwo0G9LK8K9o+
nQqNaavmhk3/acbaeo97dJSxsIK2/aR29BRXqUBtliX0/Iq6XjlclmVL6EfPL2xw1EstVVYVFXOx
6vrw7ysnEoWNxuCNcGAh7U0oialYVwX2ghgJzKpJKI6uJTVhpuiLDX8fmGL72m8Q0uQsWLaRsdBJ
OQV+cvlKKyct/BrI7UGs31Vy7PdX86OPaYAUw0VFkjqgS7on2dPdv0+9gUuthvljIISYqgSYg5oi
3lolCI5UZa9gPYicwt1LMF51o8lmvkiKSgZDa4BSy02b/r8YRCWNs82xUH5u7o8kkMiFTustydBH
6IhGuGF3eFfh1kA5ppbTkpamEqu4D18Vh+3U7bfel59I8iWmlv8IHkVfpVh2UPrAJ0GznB6pAnue
pXqKLeikNTVHDfyrwd0IalAxHrHryjgvNMQcmxcUBC4/yV4Vrm5nOMxTEoKwfeGA4EiUD2n330Sp
WxyrXfcFERUunPw23K9aiM/rAbsksM1/IojXkhzy9FXaybMNv8tY56S2oajrXKrN1cQpK5o+IARi
O9zxPrmwrexzZ7XCgjMuK4P6xASVP+r6eJnGN2e+16BmZWs3/uHWSErmDJyppJJoc8YkmgecOIKT
JQ01ADdkx8sp9XjQ1G3SYSnYuioauY35zcclp5Bf0NRPjW7T1gWofBEujchb7vvu5va4OpO4AEVX
dzZKRI1TsNNSa/m+KDTVVOpQ6ExzbA1tp6wPcY5FCBG3ABVcXh2xA4OWQxT0OGtsUvwrb4Ye1bMQ
cXCoMuJXs9fcCd3Qdk/VOsKd/0pby2o0gAEi9ap81fiaGEwq3Or7eqeQU9bXcBSulk4EVTKX8l3q
jS9gKLCEKIHZ7Dr1LeNfVepAbNa2pKzintY3cTqAIxdmdSrcgOx7gUfYwBXYH7shjtqTHirJPsfW
Y/t1cVGJ4C6atsNV3HJneftRn3uZ9cpL+UlVHZUlse7USIs6gaQ0YBJbghbi00ylwkkEX9NhCR+J
KD7QoUOIk54A4AtKglMx/0O+n57MGxkpC1xyOtqtlPK+Ekf4OrLyDJuSISjI2V1Nr2TojreVAeQt
egNtczRW9sa7UDrt7ET29tvy+qTxu5k/JXx8k9PcOtU+4+Y0IHA5zi6xpbxJv1c13PWckCxIe1Rr
lAT3JBrlq+iSafS16SYZYayhRLf+DVMeesqnBcEX5SQs3+i60Y7wl4hAyLhuEWNMgQVF2DiwcMOC
Ixulz6P7XFCn/4yD/0wI98ugzgIWtROg85oGxCbK1nCUlnjuA0dZmsB3C8pyBzISDw5EiOF73Qan
QlMjY33mUdkoBl/J6FrO7+zeWj9Xsx1Gb3eCsDSTPRDbAqY5zTq6Rid1+BBJGgZm/Ij2AupxUKAi
CbG3zo4I4pFfeBP9VjT8hrfDZ75t4eJMkBSzXMlcDqLc9rSan+Ldg6Eq2z9d00RLGxYrDbOrNzwo
NdhUlYpaAxdNjRq6dMpcK06DTvWSPGKHRjtvS2BZlw2xkwWNz+Ja1akFV6Xra1ecMohGcZXYHLsf
DB4RxRjS/V8ImeLJBDYLGLIjkVqPMrNmv2WrbBfqmK1bX/wL8cwEo9Fra0ug1kMQI4izdSCRA8MP
+dmUABvGWPBolF3Lyap2G7L+M5NX6dQO/E4QfQ/M9UB+4lCY1kCakRo152W2jaBbz573254hsA05
SYo8GURO6gRBWoi8AyUfGBXoVIK0TKuwIJ+lQlmyIGP8tQke/rwA3L2tveG8e5Uv3pTmweylyW03
/+x7bOzYLT5kHHNlbPtY3XlNdytYhWb/fZRdUTuw0BZVsR7LaIn84MEZP883VR3i8nUqxIWqokX/
PpyrOluQWK7+uEc3fkIqSk/KYqz+JFY9oaUq8sjUlmLVv1jZEvtQFDwgOlV9zMrfQwIgnnAfSaCd
Duh1e7372+Qx3+uz4LGekygQODqoksTqL72Wmiu7ndx8aPnUDeQKNJyjn5/OqOExM1ChTkvbz5Rx
NuBWuJnig/MJJhgexWH7VyDKSLtz3bbIpKZMN9WA5sAILgy7WwdI9U5LnzHXD7yuLaUEapyksMw+
3eMoEeFwYv3RQRSHCf8SgSo5vKWnN8qixEw4rmTDKM/8MI5Dti/ZrFpSQCoy2J53QBB2c1dbe0JL
cpEI+H8voEQx4PTwrkjbjpVbsQdd4KSjuASwHmymIcjJomSLL/jLLlDtCj/lS+22ukoDMh3WClSZ
6mkOC7wrU3nYwpozm1trJhehFZ0QMrHwDIWVDhZnjff51eX4KTyc2FuzQ5DJZWMKN7GZAfx3NM6D
jofL/tm7rqKr13bSpeSwYsyyYxvjJwmroRTR+BK40VQFFdbZgLGNv4qL/7hIJNxQx0mVDgi0YAwE
IGUJlwxrrF1qn88x8uk3dv1uYxt59m2bL1AfK0PKhqVEIS8UdkFosj/+51mCC6svjd0G9AdYEfKO
kl5wLeISjZ9e3aYljKGnu96bo0aEerSTcZy1IS58T3Xpe/75xfilqqlChSTw72+b5H/4WkYVb8RN
4Ev0RJAN+v/yhLyOq5jtrPOL4kYNrIp1aFMkhfiv67+5puInDgSf//LVPqjabN1ee2fRUfTSBqPe
xwo/IO1Kig7TmqqwbUA7U1Cg/OKaLZ1k6TgvtCzrnKvTdo8vL9yoWQuniVFK+yzfZwMtYICHCcP2
3NTtawc/Qw45+8tBpX2m07ULAVX4R2OXmEF4SCNFuvzAkL4iIFOeiaZ4FG8v2MWxy3ola8w4+sb4
zOT/3fFISM79anaXawadITi9kL8lsbm3e4IWKl3iX4SepCvQBL+uXTgtWS/K1ymYY1vFYX8Q5hrI
ehkBnXNRs8lJPidc0gkAIxXROf2ZH0YOBrOo1Wn6SQ9+U9XQPiO6q40j/IU7V6N/H0jLAf/8sVvb
YXhzn1gK26D/el51uiz0g9zl4rAWlk6Hc4nNt7hmuKO88fo+C2mJB7jnxFQ8gc9aMQOXYfXoWwMr
vmLZhUHs8Bp14SGhhK+gt5/VZVCvsywmOIPny6zMguCE55EfjrDpDX/jILYz/T8R9CwIJR/BnGhd
fme5+Ta1n1x6Q1PACf+XMNn47SuDcSqiJPJVwjVMoBhHe/iq5BRMK8bFWOIkp7Mt4bB9RotY2ZyZ
FRXmpqNq5QkLeVsOxoFic/cbAfVEQMWpklyVVe2hY+BpaTTYDwL7zuzBq6GCO7BPm1lXqDQ9U44S
2cFucNLnNFWv7Ag0+AfDuQIbnZ4gi5yLvLLxTPWxX50IGy86zNDlYPgSIp+yP5D+s0qBXfpUKl40
WrWOv0nIiEk2OGZWwZn8Qym/yakRQABxqz0uw3eNPc4h80+Coxy/W4RYEOKbzr14OgrKMC6Vj/Nq
bEn1EQBRNBEVHJKfFWi2pnPZZMHuhYvOuvzAVkvVHu7PFW4FNT+z3MiIvqz6ttPMOYtn7yJjkyc/
OBzv7BPpTZ8V+W3h7VTCNxueW7/ox4BpGg+PVO/SvwUD2EIoVy11xaNQoOriBpHKE3ZvmrgHcvLm
kA5v6OCdYJYSsWizxy6/kqxOSO1lwxkeD77hzV+0eso12EbMglOGHx/ixJyLtfAHLvSu0CsBS6/a
Ks01nWhqTMZf/QJSSh91K/ZTbbpG5iDtBNIa475CUeQGH6BaFh0CmqOK21Mc/cH9eYsc+gAIZefw
OLFWXY7k31nACWrkI/z/5XN1ONe2KSD6GoLUql8CoBoh1+x3hmuoPIBgncJDhNLZ5iHnIPh7fiHG
NmqHX0eKS9KpxJR3DayD/blu1oZtK4VD9znXAB2zUcC+4uCISgScjphtKK8Kp8+Su3hZEh2tW+tG
/BaN0UrBMP4s+Xaj0FwG08ooSMW6RGn20I20lvijTb8UreRDP3/FzUHuc/iHOCS0htSgnZLs2x2/
5Gh/3BnfNkP1OYD0MibZyoGJyigaNCxeI4d8Knkvwptr5+Uib41otLcu0T03stlhZ9B/HXetPgFF
PcWnOmjN5ExIy2utsnNcqDHoVWP/ZDWSuyPQyfvwk+9VTAd9JJ7nKKUDP49K1yE9WPViOHCKOA8R
ugdWP7CSSawK1fSVc3DxKYJMg8yRbNtreOVjfgRrXSIegD9RK0MMxyvcviqfDEs3I5ZG8pbv2qm5
ghzQH8UsCKyc38vjre8fF4KGhpYi9I+8r2eaAkZxVFhftsJRHkySIW7Hj/uHQZnPqyY3kATu0XE/
rdXd6fEBmCOujSgVcobU+9eu04t8xGiy1qJsdcHas5TaRqclfazo631R5LQx+bJ77QIEYpCUPg3N
H8y4GsjkyXc1MlG58GJ/ADVZxpr6KoSkTbj5OqnCcpb+kSTiFiu4HySwmuYEuJUCde8MS8SIkeih
bHmnsRuyOrq+oanogoMdlO6N1UW9Gf1PNvQGWomluCddp553oP4m4a3YQwqL6LB7Xc69s1bOikme
O1TBWAjf32/dfVGnROxAcMMvx3ETjewLb7YIOEmZIs7RLzUm2pGq9iE3Mvg84SuHEmyX+ozMR4Zg
FtdPlrcix2Js6xYiFb0Ar2paQka81x6wa/ynWibXNWef/ryaziRP4zpajFS2ed8lqFbJVGlz4uZ6
zk7yOMbHoFeKPR52XWyRXTI5jORfg8Xn9pU8XzNAH58VEaAOEWl2s//R9CHvktMiYjz+ZqWDeFW6
Vb3iOJhrqG3sJcQ4302M1vi7/A/G6yw6RfGbJk/Sh1eEjTzmedamaAYo9PxtLh+UVBHrhNIS8B8O
Nl6t4psGPOdvDneRJkTY20FZWwlKIto2q0vL778g2hDIrggN2MR3aUAkjBCNY3UNYmUfhLUDZhLx
zBpoAk9QA7Q72QO64ZhRVxzFBZlYkrzVqOoSrouSFgIfEi6H+r6mYd+WAdXPjCQlEOqVU/vqnJlK
inorn1jd9FrDd4IB0xgE3urYDKIEg6atiK2gZWdB0rkx2plN12P8qhrJGc13zjnFqkXZbQZg1KZl
qyUickYzmYePtIZwIKDY/zzqxVckhDwwmo/bHwS2hSPEc21gr1yM1zry4o+4cmhCRuq6D72PvF0E
ToMAL8x7xQ69+XZYQdFkKYcXTlh0DYCH0eYBb6drzbkdncI3ThSR0Y1zxJtJbGivsE2xO5PC6Q7/
o40QXxFYgijbQA5hCWl8egL9+nMVS21RncgNqj5UM+glpxqc2zqOoQ4/ClkxueKiZDihO0p+D9IG
NItHwB2TNVvjRUWIx8eX7pqDNv4KWIANc/CVClW2N6wnaY5lKcl3jdNYUKNlVL4Y7vosorMRX/lU
xQj5GUSkW5tdfQRzHbX1OujDw4nXo3Zg1AP3TTbVpIvK+oUQAMtn4DffZh/oI+w0d425J/HW4LDR
juDkm1e7ldMCpwH0nWZKKdYbmclu3x6aDWX/56Hq2BocY11x8io2fkatyYCWaM5Sw4peRrODDaHM
4/zFM3WRoBT+V5a3vfDLeJXCv+5kGwHaAxTQxF4OfCMqonApw6NWwJHZjXUBEH313I3buD9rAbHV
akxFLZuZ5RIjSZLGj6q1nCcV4lpLAZZdp2VNoTwK71H/ATmzTbL2Dadm6RJ7BTaPijenVNWHQ1FV
xiY0W536JNmzVix9eEVPEzldQdv7aP5BB6Hd87fcAMrl/pszzdCYEcZonBglIQhe1quoLEr218BU
KEHA0ukz/XVRRA8WRkQ8t5ZskiyiBrdQancisNzLeLa49ZuSwgU9SwTPYvKcl4b5HmT/J+My+3NR
/1gty8QPxl8/LU3D5waraCTu9kU0qmwt0Ac7LwLM27G7+GH33zZX/mbRw+e3zEqfeULQ4oIjNw2Z
m/O65Ddpa2NL4HSUbDYiUbWoKcxdBJZWl61B1pH5/IUVGP05TZcfTUocAheiszeLzpnv+GkXzMb9
NTq80dfwdYQpPMNc4weHDOMXsoxpdVzHDXkIdDdFbOqgNBDj1MNFXFZhiguKU2j+jJpiksyZJuQ0
cp6rU+sPTOGczF9wRWLfTf/Lcm64PVeANKLm1BmLD/zQxmGWO5XRdI9HTUwCravlQSK+oNsesjsi
RHm21IT0aLpT95JpVnnodz9xnFfpzUQhsdi5+pIbfGGrlvDzOjBpEkiSSNs8/RgqFB6pAXnIAhWS
TxFRMWRlw7e1vvUW8qeXP+mxHdkrA2lh+KAlFedE0rJ2t7UaJjnsLahf3hvkkjBzjOM0aGQduZYe
j7Kh/2jeWkUVKsA+88q5F86tpc7VAd7zh7i+771Hwq3p6lU6ONqy2bhaPTopHsSHVNAcgOUyI1k8
jFpvIyNlDFdndC2txC5kuTRsjLlpEk+Is2J9rur/1WYbGLZNI9G78sxaoQfPwCgEoWPxg4efKDBS
7G/s1yFt2WUwkykuL1Cop8nP2BonCT+BKcFqgTF86q9YppmRLtKfAOVon0LuMJwEQqFdqdF6COVx
9Q0azWtG5q2yFcFq4A/HY/PFrYmuW9lJTvbQqbvXbL668zyiOT2yCqY+HWgKrZhFe66BOr0F5fer
Co2ohR7XMm5t209UEZ85tA7SrTYNwie775lRkJrEjyAU+6Kzmb59Ck7goDjg8/yV0GakjZUAsLYp
SCvBCtKn/buvGZDkF9gaxrLRa93OA2k5+3QDWColK/V2rFMFcJyVCMIAu+yt60qNFI7Os6TK//Ql
g9R9TwFw51XdAJIwmhIMC+A8Eaj1R4LDKH4ZoJrGdIq7SisA/V0jatybEnRyhMaBJdcrJe/J6wef
crrJ6Gu5aj0Kkm9JA30oyqyy1gflcuQrTzqxF7s7eAgNyYmfHRT3kSD37klg+rJbVLX0+ENV9RJF
hn1AiVtv/SmQ4mhJpO7G/4mIsdRdcx/ONp7co5YYpHx2yxiETU9E8b8dbsL4YJcJ0lNnZGMDZnaL
NTqvpznygbdqO/k9nCFQeE+d3lbxYLRxLwGzJP7MWOCHvsd9Crtg9ys0q+gGlWKgs1pO2dsWbFmJ
JVBtG6N5prfTncA5wRWu1daGCx9qLkKgKZQ0RDLFWo2inE5OuwsYUUCTa/3UJa057PXlk3TBPO0b
lb42vZt7Gf+GcAAnRf00prUDQPChdW6OgJQw6O/W8NqDFjkaX/6XGqjyqJjTxKafxRCjTN4QFsWs
7NRTSS38GpSdToMOQrZuJookU7Nkfp7fNq7we72MMaIuiNxPbtJfLuueqxP2Zg8yxB3LeobJPO1/
+dxdIinl6JffaPKumEowTflWl9Op155i7ysJE8WWreLOevTwS5oTrA3ep6fLca9Iot/5Z3eqrvZt
HJGTiBhaKNl1r8TJ8BoY8fuEexycIWhoQymqxPzG5w6mVRW44iLdaNh1hsgDMwbVu8Osd9rwqV+y
8ytrxt2NbQ8Ms/Y2eXyev5X059SGPoTNfHwGCTEI2mx1XvtUV0bgXYIMo7/T0pdKBVeFfrCnCjFF
GQvA55OSOgXPTWzwHd49iG3zD1vuvojDEL6HQqmkFUBetcOWUuwVHwxmBFRkKQ8MYGcuzC1RUK2m
uZO+GtxuXappPWFhyqNz7cEQuemVFe+Vj0Vc1kU9x7qSonx51AnpeHK+uIxFpbkgkLqxizTSiDmU
+aFvUVrIKYZ4V6PTBBnRSAHFJc8mcNCtFphrUgKyxgAOItKX8sFBNTHZbTxz3dnVjH+cS26SUWHe
h6rF78Jm8cLC9RGAUJ71JzharYs7b/niZ4izse7CxVho0KRVQYGmkiVgOVa78ScXUyEHaiiCMsyK
zITL4NdTvUONonODexCs2/7zojQBgdMAQudToOPveGv8UkpIzpELWKvMYxFCkTnlo2gD0R8T3H8W
hYVu2xMKYyIRKbI7gAMzLVLB59axo0TS2WqWgNqbLteVqsSWmBv9ez8lqyw0RnYBoiRolYyX8qu4
vWqXDwE2GYcdpwERKYDLrbGcgc+VxRj7j+Odpe212xBr5nRFHBo8Od4nd182J5ZphPQAvgAfmrPj
xZZAzcYaRjWFTJVyNuJ1xlV79fmCWLkvMFNXAnJYoB9VB6BVxOC68Bjm1vKu3erUGQpp3sq/r1xP
HxDVrEim7xdHq19qx4iBHvsS2NmxVjFpKa3ezKhIeqhlkDigswEyJK6QudiIJ47ltV4afULHCOnA
hFq/tkjHTz+mL11wtCWaFs1mS4ClSGJ9aYSkTlgRo7rzZXCDyYZKQMNhB59euxTlcK9nHHGZjfNO
qQoj9HoVfPc2havqjL8c7b5y9Hhv28gNAEhvy/OrD61oen53rR8WBKRcu3ASMUD1LxjmHKrCEYvj
7NJU0SU4j0xCXhvfymvvSv52xqhmLfmfUwVJpiBWmMBgaLB9PwfClZsnwZNIFbodiDY0EZAHCU7z
+tR798Ktt1rnu/FYHV3TMeBPveCwTTxUkSFB1R41GM5aK898ZSbosAfRi6sP+JvT0lXUeyfrLx3C
15qmAok4eIvvvKc+19alz5S3kS3jCLTNrfqEOF8VCyUVALJSMWoxjBn2X+Yj+5rE1RMUFIWWsI2a
Zvig6P2UD6PlpC4gGSKukgUCJSQUpg4ObIaUSCH8LU0L1W+rdZUV8QItNhZwhuWOg/5PdJPAgP1N
y9PrfEWE8Ytrpu1EgDdffFuQox3lhNC1eqyvka/dCF2+ef7y37rk8rwNiwW7KJFbzU/ILmhtSjbs
EwuUOTU9S1VX9G/N2CfcxGXtgFxXmDgu/jCcTTge4brJn4uDnqicHn2SyCvJWxjZWcGGjC35a/dh
Z7vf0+Qn5T7DkybGbwbe6TaD9slckjAJm/Vbtw64SeXI5+/QF4FCnOp5JOJwBLupTxbZk42dbih/
OpRKCS4OC73/J8rkBN+cSLQtVAwTXJTa/QvyxLTYgFWSMyyKXurwhkr4KEgKwJFCnOnCexC/x3zv
V6R31XmHJ1LtYe9rKFmv1mOxxOymgvY21GQOi1uJQacgLUXMFNiUTR/ut8vKoVUHVe1kro4rxr0x
tFiVn6OegxtY4NmnfYP/2VAb/sjwxlkppJqMQCsIqxOouhI7AUfP6crl6i+mjDSWDE9x1va24xwE
At+ewe4oxyED/s9jX1u9l3JG0/67zS7rRA5w9fF6A1LCN7w3LUW2tmfAhr/WXOl4FeluHxDhpdAe
UGwtJeXgVyrOwCT1+qc/WdMh3BlfSSKggrFjTMUOAlLcZawIgyK51Hj/B1UEjQddKiBxWf3KjPaL
+Qsg8BlwFpC5wvcw4K3WmM5U/6wFsKIauoCJAcZT1Zyf9jT9RoCUX+P4cmcBHRx0EnHwy1euOURP
Yfg3QMKzzfuqF6IXYUr/gi7PJpA/rtzEbHdeXdFV1prTyt6USK24n9ce50zFb65Mcq8qm+vFU/oj
k5T521BBKg4jLFnmIWRUmFYg/pxxzQ+5+/avpj3vXdXydjBbRRoSJ9/BqIfBDbz0SLgGcCs50pfo
EJhCAoaEdbRmkIxp1JhRGwu/b/gvFczyU3JgCDG8sZnKKRvxL3lVjmPi1REd2mJo/ba/l/1k5i0X
/Q/f9SHW2IUfXCBd023w5JtAaGGEQxbxwfREf75OxBKJe8DMTyZXPNk7Kh1NEoTcA+gwzV2tAuwl
xubafgyHk0RrLtMwWNdLUZHtQtT8N4DhtpowzxcwfZDIL2wOrsD9r+6+rK0FFkytbkOTsFgf3a2H
Mz8qjD2+cq0S4uIXMEXQ+1xL5m2YS0jX8sjc+G110SaufXeJbKKZYn+1BomU7Hz8Wq09Ok+t651U
ONlJfxDY5jeSj7QnzKfjk1mpbNtTRxk89TVkCnf+hubKNpHG2otwgNZZePYiLC0d0eATyOj+WMz7
Tg9tala/wV4P5ZbxXHpZVQkaf6d+f3CCa8zJTztd+gC7sU+O31a7eeXGow5oK6UZQTwDZSZI6gXG
kMldg7vv6Epu3tGCpbf4CLjEwBL9+jRNJ1QQ636DNN4uui6e4KAiP53ZskC7KhrR1FXm0+WxHlP+
xn9aSxdH4YSm9LlFOhMPDrt0Bavl1S2hRPUSeoYWokUwxnmUmAfUpGepLeIT01W+ZHxhL3yc2jQW
iN2O1DvbFS/N/+PCnqvImPHU/F0Hbqc5UCBdzAyRxkAQSqKkzmhMRRAySKLFJ40dmC2hbAqSgQuQ
rIYMLFoOh/dSWXvSCGcsi8/bCv1LEKFttkjGJg697xwouKmeXeZtVOcB/aGTOhg/0KsvVunHUOBf
cAyZabKmRvgtJiimAxRLf83rqXjs29nt2YYu08xa6lMna5A7y1lJli+0M1qUhKPXrI+m2d+UXkDp
ixvU6Rw4E+WT+H3ugjQEW/wh3JJumcRO3epr9Z1z12mXjEndHeLfPRrWELy4vD1L5c/oqasmhnzE
vl548ozO+CfCSVAqgnQLjaB/VfubJvFjiClk00XDJb/SRIxmgjRtZ/dSKXDjb1iQAPN2cVsnK/wG
3wKI4h2L2VNZ0PKCygKKGPKjjn90IUAF2FqdmQ77d9bzkKbN1TqYM29aQ1tj+rdQopzEJQjOY/rF
G8qNaj1dSkxfjV4vEnFTW/cZDccPS9rc6738ijUeGoIUHsuNSlHkcBOp/nygS1P5WXjoIDevOT+i
vBcRm9FPAtUBVXRPI/Zd3QV+jw0/5cw7xmzyGESAsyCTCtiALnP2UYYyoVd9DVd/bur9UnZJmxi7
6n29T7lYbcasEokv09FHddNmNQ8LZW20eGgCoj2sAOoThyq7qAWBDFBdCmqoerUvtzbaEKFoqFkv
vGja+0zMNS8l9vltyL9W4eiWdYvGg0cNJtLttTGquK7/ettWDHfwdX3hSnTZLLImnI9tYwdW4NNu
3FVMrpkUhhBf3y9X5mAAh+yKcAtHThvMuFiYJZM1RoSF0wMSjX79+8+oPEJ1FnbM00UVJliPWY9X
neZ8R94c9TFV53oxqepnXuQ2t2UdSBUMQnEc2qsnCGorhs42j0OYbr8n3C02vj/4ERJ/2/3OTYA/
DHG+4MPV6BJD+p3EX0V67U72unR+hgInFSHkyF4la7ezGQaXLkLSRYYHEBuQZcU/ClrjPeyK5Acu
2Gl+iY3qgPFs46qVtlmBdeB8U19fhPseBzBoZYv3FPDLSlcqBQMr9f/jiIObqwEERvtLL7GY1koH
YVvHVaRJil1zdW9mnRGiXhb/iwFnOk13z6gZgLIuW5a/UPmZndpFzCCSjYziy2/4mgTFyGtK15sn
GL0ODZOnTCwcZe6i6BPt8Cls7/8sXE0QSFy38vCIJ6c56yWJKTflBrvsSklbIx3qoCk0C74J4E3w
lwJtGk75929S2cL6jdIRCIA0DGM0226Igxi1xUaKYHKRMIGbACc0qBVCATiYHKpdPG5nYGjTotEa
TysMq8hFGDkEQMzpKeQ3jNyevM2NbHkGlxSLAyJgo/BeW7kXKQ/qS/YH+kLNNWGFx+DqEF9aSp6L
cs8zVMYWfcVibi/rOTXmwL6Kok+oneJLUaahcXzNklZ3b0NqpARRuPb/i/Z0Tk78S+wwda7SEKmz
IbkS1iYNvX0WgeK3Ka7Eu9zHlNXjxvHBpzSkQF6e5LFINW00q3rGopBMHG8cB5R7o6lGTN76vRDH
etQ8Z4z8HquRkkV1xg6aHX+XxRY7vppEoWUGBFdlm/6clO9rDP6wpTUk9AHBBnJY4Lq2mOT5/ZEy
mwcjLa6IdxK/sc+yRLe2WLftARDDsPT4oFEtOMJrKIQUR0xULtT/kWr1neUXVMZnEcUd52uvGmTB
brqVgt62M42mdrImflw7p9ue4ONvNQzGPRSwVB6ZyVDc9alUUV65C+K2fFsjj0P4/esHt9oYGfjC
1t9K/Vi4Y6AQkn8MtlERPNHR9bri8byRW/Ob2bN/zIM8x6SsPbYErFkS7eLZyAPMrc37K3iNaHNH
VI5Hv+NDeIN1GntnCpcDiBZn5AFQMZY8FCkO/QnsA8GNX82hMiQlv9MjfAd3yIVYheOIKTbYa3U2
mUKKhid3UEoLYcASHP2uZ12xPSC1PskSE51lKo0e0D5d9BVVICghq+TgEkHUXi7so8Fkx2jxk7Cs
7MncnVX7vvvJgS7iNinbYNaLyrV0RadTzMd7Jll5IcwMyUWnH2fHzkE0VPT8sqRyWOK2euYwSy1V
a8iiA4jUpc5GEgdyhLPyzk0XnO/+KmenwxJenpS/iWfjMuD75njHH9y/OKF97cE7OV4qWHY07l/f
VdlySwKAkF/XLA71NqpjN/8GK0aRHFI96E8lDeVxoCRpSFZV0lJB1f2ZDwJQChhoJAwPcUhpqlDj
JWgifYeDq/o3xXhAwbwQTQeB4JEnF2+Q3iliK64sk1bm/QJ4DB26F0Slw8brPhG3sF7DH0BbgaY1
yCh4vJmEoL9lHKrab/rPc2Tnyi8n+NvPYcGbRBs2OmKSf75ATWDB/KJ52yplqCGg6Z6hLsfJhPOE
0Sm4W806dm2wJheT4W3r0aVLZEsAqW+uTsC3W76aP7mPS5KhR5WdVM1wld1K5O89zs3Zsh5DP2XT
lKtpljHIRXZVlf7WmEKMSub40yc92/5q6hMRDT7+biid6/7+l/4f1rlqto6/gOg4f2nVA/4vKz3t
EcO5cCBeYrdzMdVvbHpehTfzVP5schp3p2LEY6WzZvbr5LH/LyJgqNT8HVgrkfAcK/Vn6omk2xHp
np+topnZ7yXmOTZn+Jc1Zm6mvG1FCwImlKWE9PA0ZjI3potvZZWLWQSW0LzpCrWDMFohzDN42GUK
HAVLLhmWqepMMj6u4l6WaT/jpXxXQov7/aSSFWKO/2jLWDn/PdbnY6JHxbjQtXOL/tMo59jBj4Z1
WPep5Vtm97e3X+bucflHpRiCr+CPsDOKi+fkowm4lXrBK1GzHpV73EXpFcO9GttHaL2CCCtpS+Ur
oFsiT1MEdGH7jkJKLZ67cTygRIS8B2ItwfDLlzRjv6EwQBxxH29lgprc2WIYwKANKND++mNRyu7u
Zay59WbFaJcZSOwLL4Us2G5lMCfavS0LQ2wt5XTGCKmkb8GdyYOkSRRv3mXpTTcB8hxr38+4Dc3u
t3JhNn6MxBtOqJAFkCgk5nu36CmZJI439TdX0u9BDnISjBLseb5iH8CpxQytf4QDnBtNq3g+JyU+
I7MwpCNlpvHVStrFoZWZNr7KhB/2jfzlKFyZPr/LdmrmQcc807svSQ71vPRxg7sjS7+A9ESp1cX3
plPDh3VsfRp0q9qoO/ECpX7LNZA8WQCU/pXcGVpWBKvAlMi4T6eilquILDKuDkje0v+TuAU/XYlA
WSaRtguxRmJ5v63iVKdkiN9DjBaZkTcygPwKd0033AjFezb4Ojn4TeUrGUahRiILqRT8dfHPRz9Q
GHDqRsrMj1g+q8ffIrN8HstBo4fCYwA2VrycfjovrqKdbUE+G10nureBkJCIfLqRwSnB+dMcKMPL
S9/+aBnZbBwgbIrSlHXYTmmQhwdmbXsuz/TiSzxeoRyoGFrgwOpL91qwmwROoYHHB+px740fKk02
i+r3bjobuz+pjoK8UMQNm4km+lnKeB1dF6F/cgMbT71hoifKme6KEFVz5jD6iL4FCfp5DfquVzde
NcmkiNuyaFivXg2n8YB+YtGjWOb28waeKwmtQgz0sBcZvaKQjrSJg39Z0cmfHc7M3X14YrFiFash
vgUKfr6jPkZmqlzxxDA+Wsar7VjCh7NcpePu13MKGH4woStR0GcdpzMgW4i+92kcghV1KimFQTn5
tegrXLnAg0VGkgo4KrJuvoVIDssVc6K8edyVJ0bsZAv+JFBy+iYYsvHDWuHXIJuDsFptGd/tTRc5
x5IFMzureYU5wu/tZjcDnYIrFChAMisdagMZFgu/96c0bKDeg204Ognhuowr4IGUoG5JsTsFg5bc
IUT9J4TNZ1yQwBFSKKlS8uN4Ym1zDD4XrqB5kPpeFDr7dsvAI6kJ1sDH7Qg/cRw6BtgckmfBdp4W
+H9YLI+wwFT9pHJGAkDRwp8JSiMjyMJimXd1ny+xS40hrDW6c8epL9kPPjeXQivrGpulhpF61qAL
hvWbIcv2otOtifspMbpub0ryUKZPovqRZVtt4YLxrIVu2Q8QPnVSFGqw5sKAA5ikB42Ww8Skr1D+
ctcKkJI3CeYpTSiycXk78yxkUJT8lkgK0tfW8dNEvwzEGVniZbVtSxTdbw5TUfZd2ux2jHwZ9gLc
ZqObt6vNqvTYsuv9ns74CaFoJU3T1KCWrJ0+ffM5xTLSHlfr8FdJW/jhfspUh6bDiRtxWPi0Xgpr
OkIahEdC72EsqbAZSUL8tXrLsqO3yMVz+8rhmVeeZV9BeVitzXiyOfst8Pc9IYAiUdrZ0JQnlXHI
MglJ9yfvt/cI4PYkEFivRgxllMBx5+VpF87kR6vNs1D0J7A5UIBKpAkJ4tXtxlN7pIMVF2JGWk4k
M8cs0StYfx9tKpR29TZaFrFIHQ6LqYNrZHi+6Cz2rmt4xea4KTBklY69DD9QYQS5VZ7ldVK8PghC
uWNz7oj3BKPMbR8nHZNGvcKTTC6c5QfCDU/zUCCNFdj6t5uQzitk3kOJme3sSZ8kbLtrZZGkYg+C
EvujHrIGhouKYG3aKC5sJ07hkKcWksJDdclzCgy/0Ol6jyMW7OY5lBolYDE2ic59Mbg2HVQkWNmG
bV2lskSE/ujzH9jMrzgJ/S+X6q3q7bzYDWj+X+KBDiiMTuUFyE/aUMp77Jnu6EAk5FwDiPWDXhmr
J7lH5yz6DUKtWlL1rW8ye/4pk4VOobxHZv03M1b5/bLCh5DUE9NA3RClchyNX9yhWjsEheOjCk9l
yu5M/7/Xl/LiifNOLM8/EtwPOdN1cJnF0kh6Hf2C+XllrB1lSxtP885Yw/gOUulVniqiqArwAap3
BeqD7+CjpDpozWAmgtxyoq+9LRVsm9SKtH6Izw8MJdy0EeXv5RSapGdt4tgi6myXUc/3gl/KTY8H
6qnk0Pm8atGTP6IHTyM+mR14+pJw2Rb1tBHrELDytvfE9hKkFdSu508vS2eI1g2OBPTXgfrloM1I
DxG83QUI5MmmI8LG7+sE3uYNabJixr7m+X+t5YMkkQXMUT7X/9SyVcjlQYcOH+swK6y4tPSXQgWc
u0F6oXP6McIFagY+aX99RjmFwOHWMMzl3rV16ejbCO6XbHXzg8zHu8nA1VMSl/DwVCtsNeZu703i
F9d6miCmWNk5Y45klCVyVJTIypXiGukaW7n1hDjB20YVJHpu+TBghTQOH/IDklYCi5pLUEQ0c7ee
wJvyGWm9ioYzJUsCch8PH2s7pAmDcWXuchAI95WBpTvcu2h596J1fGVmTIWEvwHWbekfDpvS7URS
0ytPhQOJnN4ZFtswR9U7vHjbQQoV4rf/WCGz7Yu9/MYRa/dB+MrXL15T2JIzW7OF7NwtukkArm4W
n1AOsIbceOiLmbcVOThdnGrVrbsru2NDluFXkCpWSKi5EaZPqz9vOU2CZNI+/gtpIDF1FL7XfPB1
mYkisIoWkLIwId2Y+b04uPwelsS/afIVYoWOv/XW1+Zuawa15EL1ma8PTOcpsyxJPTRuCGSXHRab
maTfPsyDcLw6jw06lXM0RfM5zwWDLzoMd3nJ+96tGA9ffhPZV8yVDdKQnr27TcnEzBwN2zipoqRh
GEHDfG9lSpmfdM4TLYU/rrDAzxuSt/90gg4eQuSjWVb3ilclA1euQWS08C2qUBLqsBywfUPPyvvv
9AblGs21UGf/fjc7Jyo38+SFE9DrWVDnkwl1LNnuwEDW47ZJzTsMte/F1v+hjwzkGfUFd8MJEzG9
pLf3fGCKgv+undc+kzFELmnViG7989DCnzo6uy+qWV56xI4y4HKTS6gJXaCtBAmfBk326nYVVDYc
QGIAaHrOARxldybPCmEX3eoJuMfq3CSw9hGcxz916n6VpsXXlhTOwIXtMRzC0zX5L4qii1PPKEgO
jw6yvSo2n/LI4yEPwnmpGTYGOreWKWkCU1ruRikDMjzRkj4E78mmgwZnOHz4uPFdLiPZal+BYxNl
d35zZAU9+OJ+zi4Qdfn5juoJlwf/BGMkwWrnL7tNYTU2dKLWPgUHqZvbNxrjfCG/EC4qr24xQgJ9
8C6KPlcc6z9E0vk/AOxhtG/jB+Y9033HrQ9mnG1pxkRDLxCZI1/i35QNwvl81tb3La6tCG5O8nPa
ZGGWupVsV0CaJ014hee2JzBTuY59WtfvVUXRJf72Dz/zCeCORKgk72G7Nd1AK2Tg5U1agdxYkky1
WbFDqfDO8TkV7/d/qWF1QrOubcZ79E+XnI4wKaUgn99QLEYC8AhdlL0LSVfeNskpFLlBruE4ypr2
YPA+E5HuEMJs/rveCf0Ujv7+GG67UKP4NqajxGzKTGcus+a19atWa6S/OSNdQ3Gdyob57I5RjF+k
vpswUbKoWYrXZDqLqBquC36OUVElA558+U088zKun5XDKRaBHebYBDLj0eMk59Llr92FlISK2p0S
SmiNX8xeGzEGBFUvlPusEtoCPwrZ0XvqhYU9haakK4AFjt9vFREYz11W3pUM2r8+dMUkHd0GAmdn
REclJwcAsoX+USdd3aNoKRuE1ab3SWgNEwMXGjtvrunlJ3AhZ8fRkKZMwdj5WgHInUDlEhOTFwYa
LAOFyK3MrBF2WYbM6JWhM7K6lnncqGElY01R1DFHs8c/TsavkG90xOyRl2GI0+xd4Bz17z+mYeKb
x5b2qjAFqgZpm7Nql6/memRl8zyuASDa86BTUKvpIKjQ1/s1Ug1LqwV12rT0pTDrNiSy9xmmaZXo
c573ZpHV5DvjH8dHB/VwxyznJI6WN30AlVfKfDMQEh++WrG21W8hoS1kYwl8USfFisKhmlrVBmWj
MXQyT4A2KsamwywjPQNC5yu0y0Q5B38I/Ps7+tse++KdZHQZ+pxvrredY/tQeHrdEVZbFITXGkB+
ZQFYPVsX/F1WKzhgeYM0+rzsSU2FZitFs/01ux+PerqivC+XDj7+1207dc+8Zup8kxGfC7vVtOLH
+82dckBP5Ym1RcERnvCULuRLw3RLCizNH1VhGpkxmDVm7o0Zz8abTc6Xo7qG6LVv3rLhwH61FSDe
CzUqsDRhj8b/P065uZuzHRB9LSJzZ3KlOzUuaF9c76A8S1zKReoQV6YNlus0BRgr1hb0P1aBAtfY
llTBYhUCnUakA8vFWC/JxO7xHkMxD76LYr8LCOOZustqZyFNh1OOgODDWCIf4a9JME3IdGbU4MrL
33RBMfol2Po3wCLWR4CvGLX86DP+kJlXJuB46v4VXcZ2nIOVD7OUj+kH10wWA918w6A5lJ7x7NTK
IAXH+qSRdw9knIeLqQwtKASsy3aWYElh17ws40vgsqAnAyMRGVrRq05oNSBowy6tmIEYGTEN3mK/
FKFAESabb5Ddl09DxJg/lP6+hbA3qvxS3cD7qMYw68+ai7gfOW0BHqc4u1CQgewNDomtDT1aSxxP
uMqly7D/aU6GkaAfcNaXZbciTGmW3ZaQrEX6Nqn92rKOMXcFMe2pzh3mgOxlhmikpK3qc+2kIO6f
y6CmnJH3xeb6KYovY3Z0FA5FK/P5BGylrA/DzSWELSGBJZwXrp5V0vpL7EM1NTj+2coJ8MkzWHlg
SAnMTPgPrQO0qzCUNs22azRlgTFcQTLe7JBs89YghXZRlNgU6oe8nmySG5AhGnXt43zPAP8IjEeC
VMGLHfoO4nF5/noUqE2o0Lp7cwKJhuB2IAyRulv6frK+h1JZ8IlmFAateTONYGuOmSXnROgGNsoX
yG4s9HlXogpO9GfAlgieQe3JwQlX1AmoSxN7PobmOh+CkZPtSdJJJ3PDoPhhVfesC2PpjOm3ytWj
sdaRv1qcR1Yse89Qx1OaoCQbDhwGULTd9wCUSgcH1q735UemVynMaSzF7UCesWNDTESuO1Ix5gEj
AUBvorA9oSbjwXaqg1qoQuvndj3jpZPLhbUmBhtYkLzg+/gQALyIBc3BJmb3391k/PYbg/vGVTz6
C4U49ihtPxfWhf3yaOBe5pSuP0m/gELeJLOEd6boQ6BjM0irtQa+VDzqd3D1Ze+RBRgTLkaCfAUg
Cf1kZRH2VUrENUdBXOFBsLpMdJjd5eLgIb8Ev2Xkymbtl7HvaSMzGb/OYDewdAhWuIki4T/dZVcV
fM8EAaLj7A0Bpd6G2gwJEk0fbT1mcUNZMlKDBAE6QWqBI7Emh7vRYKMsRjWr7r2PwliyByKi0g1e
WC/U/TrYxZuiJKSCkP5CfBGPodJmVC2kdWw7MlO7CKRKGyMKuVWW6etNhFvLTZz79HJPwh3n08OR
9cT4wJ5ALj3Y5boNZckLFT7ngOTFpyEWtHlq4zQ8WoOV2HozqP6A2Q982oDylBZxc7OWbbUt0wqw
+owZ3yX5P0Zh5ARpgpaQMXTtsyPNKG4Bg/isb79536GDCRwkqCnZpPQdU3iDongC3oS/cyqpXhgY
AW8cpYZCahcawsjKrjGRoi8HlE0HGnJ3I9LjNJbeNPoaxwEBorb3rLSGVTitvU+yGljo/ZjGuutz
UoLqy85vBDt8qBDgQiCmOIsy0OHl9dWarzmwfehCpnJrbh2oUdAWnFEhjc4oKNJV4xW7u6jXo4Ug
UB7uBCU84p+TUHHDqr3AL2OL/CAekz9H4JBUJ5zXtI1mpRLjkmKxCOUKiOTQXxmE/nCfBBFXAj5a
+SGzdkGtDRvRU3M5moxvrPKSKKP/xenq7V7YiUi3auYPuPkIUDX/OyLIWu9przI/2ibKw7GZmo5p
I+d84ObtN+Tniqqrr/0HW0rcIRO1tq++zmpUc8ehj1cmFHdUO5ZL2noXUzUkEBq+9GKUI17ZhNT4
PQCTXO3diJzoc/aPqSXg2jPjuu5p+/OmpNJn/7lKskwXyVK5A8rK2UN26cwco/NY8k6+SnzbEdxZ
1ra3ofgoOry82RyvY/kVsiUM5NFXYlfDUcQo3FpPmoCE7K3r5OlGPopZ2hN4jBVhzNp/KxWn7PpU
fIizHVJbZ2amFw7Q8DYv42UtCnUD6b24N3XY3P9dKkoMN9dcvwUjRXHTz+pY1nLwoZSNPCUnd4T/
zUIXWeEew4YdIlG/A127pffgc1zSBWw+UnPT/fMjpEzCJ4YQWuJEzKx/KjP4I1BQ14N+mVd3y2Cc
EqQ9EU2uOVioFTrHR/8SnoPeP449wQgWFxH9SUjoknxhbMLeK0r5A64MPrW5b9cDgOcm2dFGOEsa
BozU5IFb84sA03kI3K0YuWxLePqKffLhzcnvEvgZ3cS2BJll16e24Rz5r030qtfjTM2rFM11HHNs
5LWVqySZlmUDKKW1xIzXFSsIOBZRUMkiJL0LiyA/f2L7FXERxLCxrPZOp67UeuIjYGNUy2Am98j1
DarF5fyDxzU8sF7YVsCo+ZS21670jPcUpBaFXSngEI1EUK0X1X9l8ZGFkCArML9PC2BEkeEuFFsJ
d6VJsiStyNNjL439CFQ22aR+Y/dOa3qufIcl+o2oIeMxtmiEiYcpE3fkQUt8Ja6fUwYCGvIxaaSV
rF+0yu6Q8iMorVItHyVmUNFmTYQaEFSrIMMQbUrAxRYh9LP4GBYKVRqvknV3BMn2tkGmA+A7xsT0
/VVdyvP2QFSsuoKh/2AkXIIvzMtdNbvJmsFaC2egd9EEEOO21dLVPbq2dwNsAvVq1G0m4uUKld+J
edORfP+EKZRC23y342ihPkE7ThcRZ1Y4CxN7Nx7lEiAeMEHGYyDkPRE8B27XaoVvpxKjQ4idzQdo
v7ycS4DeV57/luHb6E5E52BEgcoNr9ufJ2M+9woZ49hL6LrK/ToKqv9xl7S3pfkSKk3rURU5G4PB
WxnMKyOj5UwqNCoBHyN1Z9AAZOCIjhWNHgMaNBmgzdZxpa7gaF4VpEKRgGc+IjwejOhkN4vbk0RZ
Kqhs6F29d2SBK60V/mv7E7B22HvuYKTKn5ZnsBpyRWqCC7/VgeSJs60wgI1gkdZvhTXVTsaRInKk
DUthxdEgRTl78trc/paB0T03K+O/tApOd5mNFuSp29LgCwHalXIgtA2PfFkyRllp+miduoYzNq/e
lQnJGqa4Xun38UtBdGUvc+sIA3T8lUubCfg2REGHFntXDt6tIjwhHjEv1PbxXYlxknMbTiovY9GK
MwNYaVaQlO9kLHUrNkMWPOO3fVvDOKfq9xv5Qb2lI9NkpjYQQat/c681WEhyfVsndEUFPX9bHO71
1R7lZE59CaRs6wj9uDuvZwL5hUjz/dULP2wYHrIj/F4moZu694qMmUQWOHrM7z5vomm33MlIvZP4
3KZkaV5OLsMVgga5VyLeSkOnIi+aRRPaVbWeQphft0NEpMFeodSjJ914AIYAEDRMt2Vk4f3Inw41
sNe+45vbGDcH6suRMw055uS3V9KvRzRHjbB4FpLcrQdJlJjtXqdcmihgb5uW89Nc7vd/QgdJmlMc
U63O2AU2bW/2/nkIj0lkOWCJ0I5G6wB+GoMhWFZEqp4bVTdsVGW1W1iJYdvn/hCS830EGpYW4x0f
hrdjlbEBhuF9aVJ6Nv6s8eAFK/D6cJI9syrtvhtPIEvHXspf87IUCetl7J987R5U3aGnrOnbEygE
XWei0fAAh6y3E0yp0A6hMPzB89dgq8CviDJExqnbK2ZKa6x6UxDpPvHwwScvO3Ph/9dFtGqAv7G2
r4lZsrPkv/FWGWU+pIpBeVY95fq0naGYqBfEuRc9nqtfq8KPJtEMHfAwh6Rh8vxGZSr13+eDyL2F
tod1XTr0sc3KuDn1TfyYqvTjSZSJX+gtVBgN69p/BYRmN3vFxiH0AUMKsu7ANRJey2iTU5OGR9MY
ZsVNG9KG7bNI5Cb08YTVu9rEjUtozVcQdnzawLxyyBSOUnB1LqOONNbBMir2zziT91U8nHtnKkoA
6ORr9EESylUeh2UBhiCH7e7pUSC1V/tR4wjXXIgZN5lvMWkJKc5jirMGv/QIN5aycO9dzHn3CoSA
YsQVjdsNMbD+V8H2S78pQNDlcfQrwjDBARaIxF3a0msuQlr32Km5H575OYVFmpo2KGNbNM9a0xoN
BOPXSPn6ItzwWnMjW+sJbODON3bAJYBJr77u74qkOG7cLaUFwEsepf7U23kFvDmU+axzKMDOjWs/
suBIqHVdj+PjzUPisgHwG5xA6KXO8YhvGMnMvXCJBHFO7Boz8128hCZ5273u22NTFo44I0rMWtzo
DiLZ4zSKxo7FLSI5k9EfVD1aCDn9p1dr7lY+ekyndq3qzJIAa4hhFrXzkIBuWE4bcbnLnj5FpxIB
9mHEuH0dQBAurwv6MPbnkSgZKTHs1x5qc/RV3wPkKRSO1SwKKRLle9ugH5nynvqZSxeo6fCV/sev
XCNa0UDSzdzjQvADDEU0G17d4zZZEPXhhBOREmNzZHDFzAr+6k5p1LHiUTkC9D5hK/eytVxQdxip
hqV7xekNRtE3EFaEj09Ahx+eDOgEmNc1O7eMQl6GF8CmJmB5ChC8hQOm6ANhdMx+xPPtcffa3QEK
4tmqt1zyppa0rbn87ZEN9cnCmujXLeLsHDrG73uz7pshDgZkqzCPWI6MGfZdoG9QVJJA4Tar5hb2
WhA+eJUDEDPi84lX8dSTAkdQh+obLOj9sUBU4A5uv9i852hsMpLdWQZ2oELCnlWJV35ZcfJkaVjS
TEKYnXY+GhwUxeWbfG200SrNnG4t/wcGGfhO2RCZi04IkGD0wfxq9fF8QnybCJMfLuMobHp4CL2N
tSdJV2AH8KX5VunfFp4ddwWkd8AdAPF8cPLMSoWIns0y32p5bbqmfrWhrz6CdQI+xkn9I+USvHll
EwMwjpGRtOCnc17rTepQMpNZuXutDy/TsiekDxeOqoTMpsIbJNODDTZLk2XqESYiJC/LO9+1LAX0
yij7V4c3HkN2xS4czE3vnxHbnGeousFzKxeFXDfWbk3OZsOEmCYWIAnHY29hRsv0rxkMpnyhHZiN
fFdlsERjdBptvPzfl1fvOUC4hXGSfPLGwSyhP32hTS14d8SbXiHiz7/DJ0+5463jYTtD7R2aE/2V
vhQAu8MlCL/q4bQ1wlb0wBBw4tIPiDsSmiAC97vhW3TiGCLD2prRuiL55DwRdIS+/MXueu5RUjCC
2DLdDFBlrLxjORWd/J42bri71Fv2IFSgwGBS8ZPIFytorEZ3mwqxQPbFKIuCbKq9uydUnrQDHoW7
+/5gXxn86HB8MqFi/KX6L/Kz0/XrVyyvzk5cXr02sG1+lcMVEFLDT9vFGMqqDjwhz3uUHeSJj9U4
kDiGsFkpTMtcndYjL14Eaziah2kPSC5lWKb7ENNzuZgLGSVV0vO4B4+CujWTuNJxk9pCDlOTMGHY
epkRHu8R+0EQew0CnKYvXiuq2FxaQmKzTrLN9fRpkNm4G3X1utwlSw2Sel9OqoNMP1jzm9XCO4LN
COeVIURNR3diqOlZvS9zxfOYPF1lJLIKH+pPDWTsC6CnHQDL7a/EwgQdyph0EPbul40Av3w7IlXa
Zqlp5pmgjAV5NJ05G6Tfds0E5NUqLUuLnvSgQawxN6gHw+mtjHO6joO6MShtjs7QmyrrDMX8B/wI
92dUIVnxWv/ny3rTCx+ckQR7ce9/Naoz3qeXdTuBdFwwcNZkTNOib1rtVsXW4g7e/Qf6UZOb9JQ+
o5j0n8Ow1GjfSAeVodADic76reORTHc4XY7ILC2qEmu4Iud/bUb7KZrp4tc2FS03gv0SNE1u+giK
CUTdQzwE1tqKJYqMqQyGJd4gj5AtIaVldvenQfpywtMAk3qMs7Fj7cJYLt0Ej7oPI8jxgMwsUcQ6
fpKMMflRWOvMZGRArLFV7Avuu/+fLGKDa4g9r6ZdOl2lsS2tWlaOKkSigAN9WZEJZzOMbn4Cm/mQ
0h+uMzmxwmJ4yn8F5tI2b7on3tI5YdAIfdLb+9Jho2P28Iy0Ucf5dCnTL+wTtV7PjgBF3w8eshZn
GUpVhMR1QpAvVXVjXS9vj+u6ALePm7qtvnkFtcClj5E3dZr/+MLtqSEJKqzEzthlib7hhVQw3z8H
ulBlfzSOwlc99XAqN67jP+4kRhhEDxRIMAgLm5+Or1h7TRwXfNH8pZYGdgdXSl9JLNVPyzy7oPlC
qAgEq3nOvB5j6pc8klzoOL/J3C2YTqr85fBySfHV4e8wwaWO2rp+3nxe72syVM+20iC5XIu4KJna
wfYVGlS6KpMufrMBlNYX9QKSgQ0blNc7XsDtJADgQf0MsST9b8xGKv5h/ahV/FNAUpufatJiiWMw
C3gjvOXKssI58d229DXylGa1Ugz0j0wHaz3uxmAU1M0qpi2AnM0srf4wTXkwM9DVBLBlYtQVkzH/
LpSp/LKMQxTWZjmStJ16ETeKoTaXcC9A/veQbhiBZzzYx1Mw1cUMsGlf0tj6+xaSc5KVLrWATIG3
dDsUjCoO+KBIQ+NEaSju7K7ow0MfvRVD2N2h9rFbA1Uu+QL0a2rCLWf8jizF8yInen5PHB33G52W
5ipYKoWN+n4gqQPhiOv/21QvOXbxEHiBpZtNsyAcionzEoHo/Kd423ywgBKJX7jNkhZznL24FIW0
0uRKnpKliD99ExSdvSvqiiPsIWdDGMSZP/Sh+nNmfx6Uu/GDc7CcKf9+twmLN2Zyr0jM9+TAuvNt
5Tt+Fz28iAlBv7I4Dg43lw05CFeiSKdu6wUKQCTzxb6Mcua7hg48SuAktKmcirOZvnTNkU7Y3HEc
E1TikwAb5AVsX23l6BnHLMsZpM8xpaHeieDfp3u+P2ZAd2q6FtyFTqKa+1u22X24PAydqiXKRdFc
uIr9X1PodohjlPeEWmaLgy3N6y3el21DrpZY2iCOsTEX16f54I/JKASx9QMZSjogo4KJRnj3Yq0o
k3qhileDRwZgZJHVCln+mxBcragoETGLy6MSvWzDB8lhFG6oCejFDNAPWPh4V7jrd7RhZWGlxCmr
YVlqbrv5TrtwIM4+8IMlXh4MscHa+3Cfxg5JYjasuy/JGZANoaeQwwnSVLPY2JZleF8aPhutKkWm
U6DSd9M36qbW0w3O7qsdrYiey+0BGqODS9ndfiCop3MQHWNQfdieS8gSvr+BTjNg1M0uvr76ZdOl
DS8jgZnJTWdwdL2ZWONrXefGXoNm7r/g8oGEOK88UCO3UnTA+YYloMyLUkxmQNRkDCvanwbwCc9n
9fTbApOA7zTaDVwS+2TTxrEduBVi6jDHWnuN79Yfta83Nu+Aab7UPPVYHDT7jSzH2hbTKCmyVab3
JLdjoE8OfL1fQCEbGwut2476A4urMk6y/EhwU4outmHalh/88U+N5t2hmViSrG4HvSQw7MhFdt1S
gcGaVsxiJzpmx23SmM65iSKKznSASxa03VIaXMRc2DxBKtXipuBZa5g1KZwpXRNtP9m24o3Xl+Wr
JW56h5VaDU66xLbIUlAp/f8B9iTIEvw1oEgW+3HMjM1EJ/pfc/Qf/AVIXHTj9B03p5ItAbcs5ZvV
6ZGVl/iJU/auc7RNjfLf7fycuhMYaf3dU2SzSns6nuWZGuaibNItrjFtpAcJ/1IN3Hz4Xq4dFGbB
/Idk7YQ7rHTdcZM9WJ6NLXYJhl0iXU0NbD1C9mIaWlZ4s8UPcCny/hrF+tRvD0RDOVFCI3WPnOG3
/chfsKZC87dXD0VhzIj9ZiCkHqIxZjwxcjgEN/R0vbbTEoWg8s2qYROP3bza/iYIwbd95idgfdbc
G6AY10C9BEi/yVC3jDmFOc0kAZvapMOO2Wh2DxIicnAVqg4owAgLKxOz2D1iqH4vipUTB0OwgwIU
ldHeUKDQEMgT7YbYgGHgX7QJFiAC200eRd6FTUafGrIX4TXUqgldLf2Xx39pxxgfN72huApkJAin
QoXehdmdRnlguCNvEL2RKqwskxYBCD9wBuXuXCCeuinbEeOEm1e3cgRi0Vwwd4NEkinR9lQTY0Cw
itlgO9WUV91o7kNkjfXujQdQfZZcv3ltX2+iSEvtlZa/ynj7vUXOTDMJ2nyLETrEhlG1LIwyrBq3
xbn2nTDTNaL4AR1zEoqh3HT/cJslQhyuLO6EjjaHYiNABBK2v023E4mKt8msS4Mm5GgDgwyJKonX
ddeMojCzRNU/dOy6U9LJZhHfLaIaJbibeHOxJIUKPC3w/WhgaMK3XHMqRGsPbxEvWfCTBufBI9ZV
8y/HViR1TfKCfBPpQheEyGYPqof2Ojh1K/6f5Ams0GzWxOtQv12LPc/ECaoohWcsq3f73EolpbLa
zlZ+yE/IowMNpazvnpLtAMkbjk7hzcmg12yjVxtEe6c1sw4IkjBloG6h5b3WcTJVFdXTpPb/aa/d
yge5Hs36YmSUCPUJd5euyG+G0uYEPcbP9GLmhQmznHWOpEvqyF6qGYlpo1FrXM5DNEPztKPDnXYu
I7GB4oenuOWdKcj90qjLg6otPROOiml9NeXG77LDaXQRgKyjENMZD2gqai+Lc9qSVAiiD5jrxjvg
MKFOcZ80ZYgFNuRF+0We5Ec24WvJ19YJELM0o8sriMoAIZ8QJmHn1r1Z/NVmLnuub/n8q84vfX/M
wk79Z0O79jBNX6MOrQ5nvXLXjTsv5dwWFe/rFcjXHaLZ8zk0U0UKC9O2t5ZPflfdb3fnMuWwIsvc
Ew+BfPJcNpSCMO7PEA+pMfShZSXkXt1ZDZuxXSI50txdsGG6oib3lXvFDaHROX7uy2D4t5ido/7E
7+fJXKOxLKGMmufxkw9vqiyXXyFoFXZLpS4v/A7k/Qdni3DZxf4Ep7CKCarZQjRbfiuFgLPV+XPf
K7o2nJN3Yhhqyjti+MSCnRcvngl4hO9HLcRzB/g437cwe5vV0V3/7li6dtsYMHinUZm1Uomh3XQB
BO/WLSMiziTru2hDwnPuGOo3ydtMcjeY348GaCbjzwBP9kCnWPYk1Qf8aVTNbJnk5EkNnvSCxRmT
rEvj/56N2X2apTKt9glisTAGE0yfrTZVNKd8G9FuGuahvL4EmpeY2IBdqF4CgLgTtJjiwpP6KNk5
XLbk366dUuipcyOHoAJ31k6z8ejseSLJ0S5aZb/rGF0kK2gRecLT58KUDIlVoPapUyZUraXCqpA2
II3STpRgOPNcv4+I+oTO+a5C0Qkcc+F3LIeK50GfyRdK+6xwoAcJkYdvZAxPdWwxDFqPTwQeAbpF
8NlQTMAppjt/N/t1KHfQdanRf60hJ9FcIeKbQWf6qRU0lPt91qKhvYn8xnF2slqqtlnBoDrebUcE
Jh0XW2p4CmSGC//PujSN1IDmPYdBWZXifd2JVjD+RNPwFZ6vmsqlcD8rb0t/RuiRgP4vhsqLONTE
XpCZG4k+VWwBK2UKD9LxVtsiSpqWAu6ws/dkwrYK6dPIxqFwlYeqAanhG+EgTZuV9SJ1qGabn0iw
JVKOeilkbjX/2qczRMjx8hlGWZjyu5VWHkCxY/XHClv821mKJMPdsCc+iQ+syjp6kj2OUpJTlNsV
76Z+l2LUxqziOBhTuHt48cPV8Zs5L/9yiT5gAhflak94URB8jVcpl0ovA0Bzk1v2AdYt7yXgjDR6
2T5dPWe3jMTipO9tM6a+V/lp9qIDkY/nDo9GG8Cg9xJKv7AuNELszCklpcy//zwvcsBwcAiUH/GN
c0386pMO0RRUbJiNo+PSUQoG3I8AW8JsKzvuqrUXGg6SXpxz9bfwxIVd73AIBtrutX442WiWR7zr
LourDNSshnt3sY8yR4pPEJMJLYzWq3CZoGW5+BelqfdeNm4MLmAq6RZEF4VQwd+5UnQlpTEfzY+W
55wYepr0reuZTsqYBZ2jEujfUt5DRoLNi3cTj+PgYjAYMeZjxQTZ5I2mZHC+H6TB+iEn1xBqk3mm
n4/kEvekZdqIKUDfFj+3X79gSPpg8D0lX2MMCrJ+1pVUevn6xtvl5i3uEqseDPjMncGg4N7NkeNA
qFrFGlo/LuIaoD+y7PWC/pOPfmHxDLB8epTvPjAnrF3WTXNJ7VC+8fkkufODGDndYC1XKPCW2vqw
rNiiIZ1t3jRuXmpyX1Vqf2CmJm1PnVkewJbPLbUtNCGOobFGdAOJGPDhTvNUwjtpu62GttVizZmK
sFwbSkxPPchxX+Ilx/+DB3gzJU5gUzzEK8TCX82P9BaE5s7dKl1S4dewK5UBAvM5rYuwlkfsI5MS
u+/Zt90AlzvXZS9gdoiYtorDBvAr8p4mFjPltLfhHuGKxKJpqB/abJxhKszj7IDp4j5AZH+L13ac
2EeuimVGLPCNB8NeVluwJQJ4ambvulmnoFKmL6CDfGUduWMMuVIg4wLihzSbOJRK91crIL/L0qk7
utTJYi8n/egQ6dMBtcfSpTSGjG+B5Pa22aIRc1fc7eNxa8kUJpsLxJnnO4MPhDG57vOS/4/xOKFe
hMmywQXcQ+E5hU6zO3JESrivMj4CQRC1vanwXCLw106V1yDrqXwp1ZWJLOLCr1Xqtiiaj78edLPk
VBUJ4Tj7xeTTQQ/qWv4YMCvHBOBZhM9M6XeMYcgWHcR2KlttPgZ/ysPtt3seG/0iauSKBFmxQvjX
AqlYQ0TzYE5C72PZ9aWFwQeTmuFiIUlvuInYKCUzb3lJCg5EBHjB56x3XVlxOOp0NBxbiSmQGcbW
fV+wvyzLlQEDdWl/ylXIQe8PeEHUhqrnVcB2fvxFuujt9NXVAW6PmwcF8pZ6hDrKh/ZKedoI1wjd
XHRdBemOd284PAHmM0FZhy6XEpi25rneymCFlrReZQX0JwZ4X4fYj0FLndSXCnOSBiMIRR0kvfiW
UR39mEhDR4ztcHYMLVLYLqmxvyZGz9nTlfmViX3dXss9vuIRC5GsarwBUfk4Jf327jUL1MTa1UNY
Z55z48wh68lAPV41+d6+Gu0qgDxVkKbuRTVahBySyI+GC+mfRuCAf7aWZchI4VYShfOlJCiBp/pM
qG1/t9kmQ3HPC8+RCD4smBFV/V430twCe8hFZ3ZEDQVyYi2iG+IU/7VPiwDajPT/yIcS3W7ZWsA2
VxrCQZoLBUkxhmONg43584wcRngKtwNWSd7b1IeKy9iCce/D5eMkbsVPr8rlwT6bIgvaKLHEIf9q
kRKIdln0zCrWqRiVjk94GimolSjFVBV2QGgQAyvB37Kh1p88Af6Sr0fhAaLTy9B2vV87jEdW34uZ
1vcZDoDBP5aK2sDqp2XKkM6Up58DcbNhmPA3NG9BTc4UXF61mk/AWyZrZHtf0tEvEgZbthy63mbO
g8BHvZ8Il2TsGq3XQl9NbboiDqj7xuNxzTe8s4BWRaV/lT3FQT/dcaRQOup4DFYDgCrSYn+T+i7c
hi88ogxgu0xm2a/0cCalGlkfHvTz8t54i3Z02hlkjvFEf00MVTwZ8eq+7rCH6cKj7Q9+5rf1SgTS
AkLQfJk1Yjyr49AQ+2NOjGaSrPux4MzB/q+1rgE8Edzu89aW4QkPxypVRRqHQM1OaiCDriFv1mu/
dbDiwa9V8rI29Qt98x0sorcoruVfRTujPf85W3O/cuFLsh7eQH6MIjX8MTD1houJwJzNz9+XNNQG
Qpnh7t/y8BjJXwWDxmKPD78I7XKiodbyokZ5touvQmEHbIPmR0F/OeSqVz3ZoJbwPmmVqJSDZrzF
H2Cx/DmadjKfXf/+9hwFKkGoeq/3enm62XqibYYqx3oFZ/ze2S5NqoOp08QF2eH/I0gCNzsCE1/v
mdVnJQIoyKhJ4toDibsab9gVcrYQvUWh9MCoYAUCpJvn3+vcn2/tGm/ryneiqwcEpl/ux7e43xib
0eZhwITR+c2Y0tVwBk9LyiRq+cWefdLZdIWzuv/xL5mM3/OgJz2YI1dCODKlJeITZIAR2tiZmOMB
a4zY0XdLG8bgbz9oqVgEiOQMCRJOg46rqTxvm9dFrm0z8Ws5Twa69pUpdye0ENczxeoABjwt5hpB
xDic6hBz3HRXnt7xFAwB3phjVwDIApi04qprdtBsHCeDmazOUXhPAG0n71DHytuQVNgNnwrrs4UD
+illrxu1X9d5w26ekIFdJAlS9iQC77DfANkRz5EK/bK4bml+UjIKGtQUZ/emD9/fFvBk+7CB34Yq
dTKW+yysbV410dn9S8pjWyXLgUw4eiiEHIjDNjGJWUODqQx8XXewe76PmoOoHpE+T5VUKzNrF+VI
nE6DEwiO9QqfJmHTmbFE1zWZBXtDyOpNzmduNCyfmMtwXriWwQbVQ/NKQG9desiQ2LmWhWP6TxsT
p8IYuNykfRrTRaqonJtJ7y3Ck0f0SMZHJ3OMvcjR5eKITVCOLcsNoCLSRrwsXaKGMw7wRPtq0QBf
R50uW4SVwUA4JDwXjFH4NGaQEziOy8m27TsSqwwKheI9zxebf1JL0cLY9Y2pCxMAbYMXgkPGw80I
0gpQbukRu2PGACEppFWrQkgMi+2K91eYJu8OVIHJHZPNsVOR8grT3i0TnaVFJFExPCo7rlOTNLCn
fe1v+0tZDtey0YjNgCR5qCqRedWetkigj5vKiXhmZUBG+vRgzq7C2o63d9cyy7i6C4no1b7lsEOu
kqvm4i2VdKIr9Wwfy3VKB7Zh0btUcsOGc5LcHOx+LuvJTJdSW12RQGwF7QFHIUn2KZDDLzQ+Czzq
BtKdGgBjHWjO6T1f5CEiGzeNHq6KbVuxoOkTiNdcw28b8+6W1oTt6TafTsz/yHq2uuO/tYHvsyGL
c/MVzbw3sS2S0Q6MzKlwR3p1mSxlhveP4QlmDZoqvlrPHMeXj8KoLWbOWhK97C1SWMjyYb1ynLkD
7E1PxtHOy0UURqE7epDEayR+AV4WFaO3qr2aHKA8YdH0VbN4kD7iNWvrPlVewXGR0cBt+eJtblYf
vOY0Opv9Zokx9oEycIh0J74l9BTec6Vt9LraNDndn6MVM6vbnEIrc1zfXKeIgPbPrkbwC4wWw/Me
LALZbuo7T+y5wqLhgDso9RIRZCwK6I3zEISvpaLFmzXg8dBAQv8wakwDXh55i/Dc43nGkU5HlKQw
z2/TAVaH7XxrlPWLWZncfVrLh5cp9Rsa5SHpoui1Hzwtge1YqyOul6Jl0HsHEum26HpF8qGb5qgW
QB/yFWnjA45xuhP2H1Ga2ibz/msPhvHVry6sgIEQCXY1Dg+D3WbDGoIIM5drDZZD+y93TeM+x5rS
0gtJsL44eBImtiPMltwUb5vfDPepL6/Iv+VOrBMB0WXmOriZS81dshqg2auru8fQS2VV1fZao3Zx
EdkrzMu4wP0zefk8cb+SeZ+fLaERXSFFawBsVfievH5JBgVS3q4w95COfNqASEJr7B+wCRblyEgB
xSRLTejx5gUREaXnPQfSz47GuXkZ9Nn102zcjx5J7FvlrMwcTWcdPkK9Ra0QSHYvK9VvySLHln7g
XpX5mp6jzEidoeMk6j7fP/UKa9Ji+fSKvId/J2RvpTGJ+iHwnVT5jbQFkR/dTjiBItnMm0Ln3+nv
8HyG9RZXtjpknLYvdz0PoTU4PRvNK9euw01/qst3aXck07Xclkj7Gn71Tt6AEtZwI08sJghVS9mi
gcF+hQzhaw0EgIWtsrsk6PZtsC9hddzVefjbw+Nsjw4qE1goQtpk+iCe4aAvT5x1DZODBViqQLnb
a9tSeWzbai9bfQRHRlbF5d2qcleObvPXjs7p3/uAFX92A5AkRq+kezTZxCWPIMhcYYLCntC15P2L
GXXSJ2KCoF0nVkH0zPJLiGUtipbHTgDCFSeT1OuuINusSFF6twDAHTQ0tPJUPN/d5usHS5uaUrhU
WSui+L6vsbxefb2zHdJm9j0c5xZc2d6D14nhVRVqd3FYSSN0nyQdAvf6UQIqZLeA1o3tM5VDB9HR
jmRcXcVk1zkShUh3cGN/epOYvPy4MYkTAMr/9TBMKdrx0r6NBt3f9Q+7KhIe+o88GfiKNgZkmgLp
pZquKjZoekrJIGAh7oX2WX/5u3pyuU1IzDsYCRaklzALL3xEiWlhMH9yPExOuOFH3g3qQgBqYpb3
JFexyG0GO2cque501Tfz0h00nqGLkJ8Lz7kQYrPFDUIHkeDgujNkLuqnL/sfZ0yumVhZumXWbJUA
CZrzHx5VLNWQHoIYyoZ14WkCrz5NVgzXyC7LebB9w7Meo38eEi0wqEt0C5vLEHtbBk3ep2N5kGKe
tDj+vzTuF9iRCZwURU3evdj71KAAWoN8+QSSwKBGRTSPLshxgFaWZgYEDB89QnfZ1K55QQ5QxqqU
3WLtMSZUmOPWNnaa5B7qXOw15lZMzaaEMHDNec6SUZ+OZHJtyP6PVpFM9z10sSk721HWvO4yveI3
dPt76ULamuGvIpdAO07CW02hf1jqjjrEGRIYSBPdPyuBXTcNj4ORxrVgNqXwaQyVScXTMAK7MMt/
nXc8hluPZ5Bajv3P1kJKO0Sd9jlnk2R2ZsGSAoJJ1182lF2tI1AFt3XqKL8dJYm8VnK7KE72+oU8
Ub0qLvwNAZrwd61LPBmawfvthj3zPF4xy9DDvlmIyCnNBgrxVgd5cbYUV8FQHJuQdgXwUDACXfit
iDy/RfZoPg/6Hwebahms6dy1I/5bjEO2pwkgYoCHFSZBtoGATu9wdlbK+V9KV1jJMGpzKskZ15ZD
h8NTSkZXS/DnrHZTjZF2/9xtGpDuvtbcWR5uIF+wMfMwX/LqExv9qjY9++TFqyfhPkkcrAe6zQJa
Z00AJ+u23HY3kHTvfNeOTVUsxS84TfxEHH5F4zDF4R188fcTZIaHSbAm08UbuHy4LvMrlc+zYCRS
7Nt8QNBakubQw949SeMfzA7TPgvO7qswJsQwf6bG63gOsECaJtTPRZiunIJRHKhcbQX768agtyUs
hfHOgQ83i4t8rZVsgR1SHpY6z0Mux2QnF1U1Q9o6LtotUKVVBGAUUvcK3cKr3zSOc1BWgWFoaCvd
NtE7EVKP/q0wxMXMnK8EPyiTRxzD5IkrM2/2WaNxMk8dxkGDOCEQzKuddBT/skzD9gc+fchfD6WU
pT6t/y3PuzPELUGhyZBRdyp3F0oVuzHW0lSvwlwHRso8rjukcaZ5jPDjJtQCcfE2IC5j6w2r+Zj6
6w+gSG2hcj+8D8epRkdrx1DB9jQL/7yzi0tWOWezIfgwto3EeNIrZScwLfPiq4yU6sQ+Ref89MZW
Of1T7HGE4/GCT0/j0uM0+1JkUNo/jnn4hb4lt7PEpaJn3kC9DxQ9ZsOrCiQNXxKo6jtqevGfSgOr
bAysV6xEmrbMbUCBqLB9ZThINRQu9BLWLpiqv1THupd6xUi++Jp/W5oq2e7eu89TmGjTpQwpxN9L
f+pceEWDz52XH4fNTsIAyfTwiQdwh2iK5OcUL+L1DSWDDep/1Nwi36OuZYQEjqK5ihcKDbpPUCBm
yGuHWH2Eem9TTOlBQnJMoVHka40s3fV1mIAzoM5hbyo6eyKeQrTmxG91W9zFvX7P/MRKVNM7bDjE
SW+lxLrsQUyuAJHMZ7O9NM5Lws+PmAnF2McGihl62vslKl0E1aVG34auHHksbsjkLVXFpZFLrr2L
by1xg3pFNJEFGWaT4U+xqpJdzuYw/O1SMRatzV9544EwTPvIKw2mgJkbA/I6CrgA/uXYlbsu/+6n
8QGZ9mPYI7JZhPfLO7I9FRjN8GCWLd+m+nFHh+lEuPY0Rc987NlV54+HYTpSh0YNH786qH8CnyTk
YcBzFBK1CuzGCtVEISwAv4DWRFF2MI8Fx53hZ1Nl5u7PSzMZvFUHS6UpxHHt7077xb+sIKy2sZVV
ffnwQT+iZknuAMJnKnUEHA/kYm5hticXZZ2b3QILP1f0f7Uvdb2a97PTjm8vS1RNWRXpStW14uVR
Huzi9R68RQBFazK2+99FqCoSiS2MxLaeMI+dHTgW2LH0v5LhLQQAPzVwEKZEH/EDF75srC9XbFug
PbSMQwbIAXDsORCBzjy8DFbpOS6n92/3yGzUA5WBXxDVJ/f0IE+fkqct5d0wk29ODwxGYIF39THD
Wzk1ss5pp9PdrTQ6C1mOLapKPsb2DYIU4eB1QSUT8vmAK9ZpJFEz6w6fsG4uqskqK8X6O2EyYcBx
GJan1Q8IpbPcPxSsyLgs67dK4rEaDU9/Ut3CjUL7hIvNMPKv+nQEnMtYpmnrhkkumYY53JvphOx7
eYyORwc05YkYh01WsJvY2WGwaf6Xo15ZNhShf2OKv5VFE2dhs/orS0bF7+e9r24ScMSScRLYqwXj
s9RKHI0e8UnlKz7XqJQxe1Q7jrZLDAR1otCxDOiHCnZXTRhQy9RwYqXeNTfhMaas0DX2mqxgE0xy
CAHdEgQQgPHklq6AngnqY60EavsfUNryxMlWOSw2hbnuc/D7C905Uzsl3omTp+H/C5XQE1C6XR3s
MlZ+e3KTFPkf6Hhb2PEtzN6NUwA+7mTWNOOQwGp9tdJMnVRc0K2eRQHrbGaOXbuY+DcrObNaP8D3
EKZXv8CR48AzJ49TbLhlRuQLIp9e6ujLs7bTxp8YicFBqRNnyTdaizF+EOEVWUNxj+xfP6Lzssys
tcHJ1+BT6kQvuBzM+ZDMtbaj5mx50gxtRIQ1sUl0wHsUTFx96d85wfEI+J2I+k+WH3iARkXe6MKP
sU1ouxj5l2ktv9WR9im8ciNEtxHsrGuS+O38SR3c6qij1hoAoQXWLxqwvqw3q4WYqUOB/DiNNXsD
bjq/Ox925yZo8iR8ndrCncdG/kadnCelTXbiSf4TiqPwwPaOSwxWaRTcjatSxWasu6UpSP+USWwr
yDFNeZHP51da5w/hTRIXz5hTBQryjM2khQJ3Lfrq/1vsWmFh0i+n1eNiXbmMU7Jk/IqIwBBxzlrk
OcPNbUh1xg1hSkJfMoMfU2iaSahpRNbsEMLwOuovEh5n+wBCK9Mcar+EoBKydswwC5EJ8oT/vAxi
ymFqWea3v3i3Ci0n85/300prgCUiN94CM3WqCMSHHgg8Ni8Y9lDjhMbat3Tp0tJWY4gLjqmWRR+y
/m7k8MQNrQf+R7R711Bq2Q5RPuIO6vhbyI6RfQ/GYJ/N+XcwMGjyDO1RdsuGyPE1KZ+6aBUE1u4S
OM41485pwZHdHMHIDUswMXXjuKdrRYbIh2q01oLA+q+apWhqkpvNlwSWwRb3OIFaraZOvvPhsPSL
wMOrc0Sl15BBIFD/UZUfXE0wM7iRFaCigwDv9lR2BklA10kv35hawHssmtxftjAkv6sSsDfL9H9B
WmgWjXaJif7miZS5MiZRJMd6uEdbt1zMqIZhe7/47ShQcWPMEDhUz4V1yL3XRDTk61suL6ntHju0
GrOSy26Mr9FId0ZTvmV367kKk3TbX8x0Y8cEHlYm9L4Z4zJEHFxlnn3PY1oL+RCnhOPnFkWbT7/3
KOABQunE0hYh6enKuyB/0Iu3ek18ujFPCH7MJaZ1VQb2vAuwh0752ikf8IrYoMgYDUUhH9+nIDHo
zdEFmIWwuUG8bUPgTARZUlXtO0fXiNNUHX41eS7YqWUlBBcP9gsYNRn43Jj/cyYDOKCeZ8CJ/hrf
NZjPip5FVVoGNvX7zfQAgLRjZeDDeq++WacoGMatE7fg/bsfr/wjqyAekJmz7d1X6gF9kIpACEWD
FgjG3qHRSzMuz4wzT/L6EWpi2IFqkpyYQ9KvQbHn8aJ0M6o+jWt8+Vtq3wamho/pzTh+NpBEPCQR
l8e25Nn3ciASVVi6ys9p9YkvlSotCwnN93TjQ/HZbNGGgoXBhYklg48v0/clAweawgG+VCn9PH9D
rZ8JyfVrF3I1Trj5QGqX3c2w3HSeIEVtzM8OuSmhI4fKbusplSAJTuf6DrUOGowLWDdW8hPSqDTg
GP6zdpdM5BSDHWpMd1Ts9xUfQcYBuVFGkYNqg9X4qJxN/6eBetaaYQyaYQz1peDrXjshUiwCi0iF
DST0QPV/44ic3ONvc5RgHIC1Y6RjH7nDRpuHz7LDzdHcq548yCKLBZ5HWZjjUQPLutjlT0XLETpf
Y4KhRWn4o1QTVcHKSsj1UpDxLZQ/bY3PK1WST9J6nVowZeEEpJC4e+i5Hy6j7BNDg+R2W7Kulgl7
v4EUMq2brV3ox8TNTruQ5AXLKWx+3ReJIqvnXSOhpBLhI1R9SKKERkKP/HLp97wYfE0tIttieA8x
IXZUZAsiaK3wSrqIoDwKRi2yYL4z38UgOMhP3PIaJ0h6j+4aODfWDcqGCEjCrkXJIYafG9NFygiP
L4EGgf7J2cRPs64/m550RLuOkC4R0ULwx+8jfPs2ZfyapkzFYn8KXFLY90wE9aDk5U8pdZ9OVYyD
cKsSp13x8p+TyHZmlzfp668kBbNJBld6fW1/pK/dhmj1iMdb5eJ5wY7FVvqhBtGilES0bnSonVLn
VIgHkItqASllNpSt8GzPqlAPWxu01KhOjVyHKSXKnXS6LCVJuAI7zS/f7B128hEaBLGIz/ba42CN
QvqyomO179b86n05VxL/4vPljIwG5Klg4Jyb7Ci32aglER5r1A73uD+wfhi2spBNN/3ruf+qhbiD
T/II7fgJJKpVIOB6fZ1+l3GceLTucQzbbQGKm9644CWwFtoqrEh6oGKjJ12GBbTBTTU+GF143S1e
NwSvT6nwZobg7+YHzyRxeyx/XclF/klUQwszIa/9DtlWFekpQR7iWzXFYdNvD3C/k6Vvhk2JBOZT
xZIBSL0q6iT1vYA1LFUFdZ3AXbVlNs0QKTaglJJfXPpQrCzGrdkdnLSoIEy0C6/odHY6atsFiBNZ
pqPZvuCvXwrmf3SXrTu5osOD9+pRlWcT+Rta4C+Ilu2zhMpQI6tCF+TPR1a7SvV1XsCwu34tOel4
HkYqXMmtX9pcDovc22SZZ9Wm20x3zH71crq5FmjrkxopDg+6m/z1Vfx1lfZjATsBacexvwgXU+Zo
HndQrNEmmSPZC5EAVMJVo14z8v6l4qcF8yOdWWE5IVW++MQpCJLtz8FMnpiovTmnZv/RVyP3zHZR
VXASJbbaG9YuPzJS7a2sOZRHNEKIR4Rh7IDR1bf2fx77O5O1GEhe+J3qWRwr6R56lshs+2P2UdlV
iE3x3S7IfRYXgjfX5Ka0p43zGbH5VpIgN2gDr1ckCgwnOJAqoUA6MJNQNzSReA2e3sKQG9op8vHC
+lDj/YYnY4V6O55ifKG7J1TTU3bDFa0bRYbfTHZL0NY0aCmvntdTVbdpWZ5N4NUdpqkCRVyG0yqb
cScJPHSW0J36JF3heaSXeGjsALB6P9DRVidLOYeTsg7Ze8KMENERBCDEP2J9oTe+iWu+HkLj5gh7
SC2LedDn+gjPMtsoNES6KzMqZxmFHEV9tpnvXD1Dsw6wJXE4fjK52my29Z3f+Wo4AIjx2+sEHagb
KapFk+ugpouUKdr3+ssgcJfjSan0pA7vGNRgPRF512qxWGY+HOjot+oguiogTqlOA8zAAQQ+GeOu
ltRRsaLhwv5i8NQj0w/XfYDCeuo8jQFJ7dFSofafboYX7F+zX/FHWQbS/rTgLCWmCHiPVupfWE55
/2f09xEnzpID6+gWXMxsl9D1pRiE7MiEsN7Qi0xEVT4YW559lE0yRUfDsOs7QPO8ZD/KQ0qB44Sm
oV7un1pkuiTogOK0hsoWD1e9q8RUF+4BQ4+YwFen4DJdcAaoCeEAcUfVdZPYYd1Uw+Xjppw+Wldc
jkmgrrgVcvE3ph4AGF5ATor9O8C0T8/TiQLobKQknUIClV1U4/V/ZMvby2nVG9c5cKiQdg8bmwoc
Z5oELy5WmyiO+sMYnFjdyZlMahtODDS0QWe0Ns08aFt7luN2Cu3cExJhlzv25gL0yX4Thfi9I5c9
txrjezdiSYQU7miThpWcRnCKmHh4KAdbzVwn37zUpop6KeSXg9g7PsC6wH5zM8ZYT/fx83lM2JcP
44mDCjgbHOmONJSPUv5XSYHBoclDhEz4EHU6f4+ZfftiAIttM7RsprGC+LlrdkYZkohnvlJwpHEg
Ycu8Ba0g1/PN26dB091Qt9pre8iZXRLJ/eaNLznJmjJEMCY+A462b4WPDYSU6RCq5LqH+XXdMDhK
k+HZpEKedti+VlA7GVBDjgkGarEdJgw0gsH8tRSjP6q3yzo4USaQ2dEjLLf1Cagb+WqZKsATUCBT
sBNxdxNDS4u9TKKG62LIPfyXFEySz852M6w9oFSG949/j5Hcs5jhg4DjQ2QVb7hnheHDzBmENxVZ
gR6NO+sG2opdLDjpX03qAKDq9DeZWzXDf1gGuhSB52sj0jBQMl4R0AMADu2NI99VfTRhShlHNUkI
S00mOHi/4Paa8nJAUtj46Pluqs6oC5Q12hJMSmPj1kN6+v5tgEHD+E60Ew1jPSTiBB1E2b8l5+0d
gd4rrY8zjMTVSH0gF6YBKVluTG5Vl1zaHHTZphIODb5SvmZwp8fPxcuC7/07gWiK6o/1x1E85ZRA
QAultAguDbsaaml2+9wa/GGnYWhQReEoU8axaa5RxLEoEBNgt/LcW61YqNuiHFGWHr1/lGKuyjs1
0ruq8vYVzSbfcL4JkMLRlPDfN2157yY+TatAItMOsKsoeJMycqPqIZJC1SznZpwIE9fNg0wGPgYU
fiiUDLBlwV18V8nZH60RjULgh31NQIME1+wRGGKLa+3kb5MZvMtE4T1Nh+M2eR7xPySWw4WxDkFD
7hGN2Z1KOfSPLj3q1td7f2K2K1aBm5FH4RnGdI/HZlbzIfcyT1Tl5qfUmk2dNwOm/7knNVuuy00l
fEg6XWALSPw5fes7ykkTwdWi4M+TpFAenLL3Pi483SB3i+ZRQe2HGACA4TiWoVpr1IVAw6Iw3NHe
5A4Edep8JLoOjxhSUfOrKFlodzS33g0YphvkawB6DXaEV1iYhpzqYMqlSheHRkARcWqvJwEnkD7z
ufo8UAhQXkyioKwq53sYMdyqK35aodZnICpueUIl9u674MfmnbO7qIwQJi9KwxUQN0Akw3ycXNqu
gB5kmQqvVf7dvHxjDMZoa28s54gNTuVmiwfOJ5TrAMquT4Ta4NbYnsW9GRvwOO3Uclx+vWOlvDHO
O0UlMYTO2SMVlpD4XORSlv3+bc+PN42gphTMShd2ILCCZe+ap0h0McijkoyajEqXldlXT43+0iXA
C85qGhdx7MAsOYDpLWFqRWHQ+h/vfViE89iNFlSaZioSgDLvMWcS7Cqq6Nbfk/5aJ+5v6vBGUlhc
gi39u2IfzwM7/J2OGc1TneDQZrOhflir5Isx5svHywXpKwfZ9A7ofCdXIgvMjnuiSuYC/eyby8qV
sOXF2AUBEuS2n/C6ZjkfIp0YQIFKwUtV+JlTGIcjq9X2NcH3i0dDWCb8FITy3++dTQn8/Rff9wbM
+HhKajpA4cDdmhzpk4BCHRe1UYJPgUHL7y3MAKVClG+5vwaykZEFwhI52a7TOTYu+Fwp96X5/zrX
0QRcwGaM8Zjc+lJJXNHzgSwHiHC8bJVG0AY9exR0zLM2RPCWAE1Vuv0jM/0AiCECXcrQxL5paddp
sK/RixPiUsjrBq/5yizeKIKzXeh+A6ZyNbMr3oCuMXjsJtvmt0dtLmjhfKPS2IEYvwpctIC8k6Yp
T/dnjpbGCgCJioH2MDpv3dY+KkvdEJ7s2DkBRLetpHU6Yy0ZIqGQIX1AV+IoCY+w1PLFCAa77UTd
VJXHzgY8DQpVWoq4TwOWZ9DznLEqN0Th8DxHW+6UUBc4N9bRFi9gesGNMl/C+YgbZsEd3YKTULbo
elFwJF7zq1vV1aYo35bBEuUiETqdUvHq/N4jlBns/WkU0HBg6KudhWnHEsIMRTibfT7nKC03pBZZ
/1QNSx8D53KjKnNvS4kd/U+YGJ2D+k34LSHKdU/JaOpclZOKfmiEEILSIlA6CQH3mCX1ZFj4Y6co
WsGmJTff/rZL+B5fOXx6G+fdptNy6Nn4cljL7ld4LWQwl2BUGIXxDriQB/aRtmOfXz8G3Dst3BRa
3TTbY4Jr7+k9U0AjmuBf98xb2F/kApJTglh7SV/SnbZzaJVuUoaxxEb+tTqQfYop2Jm1IDWN9HhD
PFvOm7iec3ypMvEuROZeT/u0WbxLtzkQA+lmlENiCO9M7lTKmQyyiheHKYZ4+wwmyEMdVIAnbKWL
GgWuG/GVXxVBRC3SqveZVllkb7aXZX5KKaHCFcIRxT6p6eyDfAnbkVYTo5y0k/xkoPFHtHA04Amx
rETqzeCrziLUMRCAzazSffXvi1mYnM/r/wBRewzrPXE4bM/7kQT9EHUDdAbCzEligAASpAS0RspC
REyn8Z8LnGvex2xOPPcjhVZ7TEF581ZsaEnQmbUqF5gLQTn4l9D/EfHSsx8F4Y01n/IffLAi88j0
Hj7Y37MXpQQo5YTwq5EISfBCwq7LaVyL4RBY2PCNTJMcNT092na2t4DS3VkLFbnC9ASw3MIoUshB
xSxbrSusoQJg/FSgf2n90wPaaJVuPEifx9YinEkCtbkg7/BHvEd2srKREZxO3l7fqZ5Hc2V83njc
4qe3bDHSl04RbgJeLfTEGJCRD8rysASgX+/SOzdzlHM8a6eImNMfKlBOoj9Jgr6elFVgGAuT/+oi
r9J97riov0iRCu9MH1V51eifYdAs1X1J50iequmGpFlHdatMcTHE14HJ1NeiZJ2LrOYo2gGUi0oV
X5hBt/X+dAwiSIGEEwEQVLQaTlE7EemOVArkbkvj+loAlBdJwaTNViqQremJfbjRuI/NwJ+2RsIX
kij6oHmrumO5GQnBWgoyt8q/aCMSAbqzTv9+cjuBjGPRZyPTiaiRoq2ogkkdxGkifkKocb8YGBnJ
+53OVcY+TQPuxoxDFZ3/ziJIAp6ZFwajBrSzQ61P1O7T+KUwJQ4eahJWIGj9UTLmmebTbkmO1mPc
ztSBzmGccPoAGHjhxSraevo3mpm7fAtzmNp4D5T3oBbDBe7WYjH8LtJwQF3SULKmkaGYknLWg8gp
azlc9DLOb3hNDBkbBk9trXW8RGRhlCLe/b0S7MPMyknZcQbywHftfn7kHPafWN+1s6SniJcDPnpG
1Mlcci322Z/6avJW+N95xjOhuHzTpuG15pouXukS8wbDJqKn08R+UoUr/+n64aryu3Uj/IM0abI1
TGtzk1WqI2fHMITzMLwAsROruT9iWEps3Ib+0qhnOcTFNlIkPRfDk/FJEVGt5ITw7l7UklR2bEIw
6ao9IxRbQ61pbxe4/O2EnqEvOcwuDitclRnZLK/cAxyOMLxspTtEWbSYhfPYQBgVpfeOhbjT98Bo
N+HY+J3piuCt2Am2eZhibKX+nJyT0Y0Da2ol0jUWj96lJVL4IyUJbYLKpCxJ1sZz29bmSPxuS6LU
LSSjTM4Iie2MDOxhNwTDOVe4R5orPUJBZnrqwWzAY1pnWOGa0XLFnyr0LnxeIs1MY9Y3C8QtM75p
JjxZhFS+pzDy8G/oD6IKnoVyqvoO5510gDlic4a//l5+l3IxjMbdy+i4wmcpjnPP+6q61Ma4XX1K
XGND+xriUjLlLGdWXTUntRi8ZhUe2T/mCgRfLSmKP8aCcimYP+eGLW+WWW5ZI0MqUF+eVew+2Dw/
YZYteSSYT/ZhTtTYXJcta/TVCC9ui6TwqksoGsnmutzlHEN9pa4+UmcnVajmCXHwaXlXJ9exg1/6
n0MGikP/8XWdJsDzqSI4sdJsGieemg+YeL/vFxfE7hk7nr5wEQTIS89dAS69ISTPvTRsnMSgObyN
kXubFXlDIAYsIKFLHRU/IArJKcQjJ24nwMwOt1PZQJC9CsjK1TnTlg0Lzs+FcKSHr4RGH0gbjXVN
Je3F23I4Puf2abCagMt7dQjQyAyOkmXhJSzsSr/A4MLO3d6RfiMzmpAqf6J5fRGcWM9bV246uH1V
8lptPeGx0FXajmhtXvOyn5t4OH7wwqqNfWr510fDfh9gGarPFoYLscm75tNGZgcq3FaaCPPHo1Cw
vF2xRSnv/cy0FmVyd10deeow05G8QoOOHoBykmw3ufJOslhEqQXiNchpy8YTlCayQ3aORPNW2uck
q+mSyXneyK+3czD2XLLaNIcRUVKZXiPmr+9vrEDxNtfvCJ9y4iR9Eb01QyVdHq72is/o9VswlYVa
L7fjggD02Ca4g5DdJhgUrVFQv5l3N1VvZVQ28QInazzZgwwT4t7S+cA7djCUnjBA4EVH+YxXTTJZ
Xxz5rCsbDDngtH+ykDq8raNPXe4PXxMNaqMP93wPzVSZh/XhZ09nU5Aw5bYIg2Wi+tr/a0ghiX6m
RnInG+1dhk+d0x7V5kcvbHI9hWbclUaTw+o6EASnnAmJOvchVJcfXFqBrWWXMI6rcI+Za3oAPCt7
yGNY0VPaj3zGqh9wWiWDva3vAtIKDbXT+oHxGaeYpfuRUSzkCcfy1+Ca/8ZIAqkCSIRduN998fdh
BCzpuIkLtnshbdEK3zbSNVlQfWHcCcwQPjz+wRA5oiMDlJhhkTo9nVckCke3L7T+Irzo4Nlx16vU
jC6qNbOQz57biDbSuFKcnOQdHZrvJKiVxsLyKPOmC4ubPxO8C7ycWegTWCm0Wbx+VqC5R9HVnPLv
Mkvl2CBfVcs7HBOYJXWIYLrzNzcQ3jHbBFapYttd+VUkFL84MsM8Go8m7gSd8M0qdadiZYr922Dr
Ub9/yD/2JAgBBeASbXZbKOpJJG2JX/hp010lyAGRk6BZXkROH3gT2ap4VdoXXj9p3gm9SQKLSNfH
c+GKqQ7hCxxTREYV23qbSSK64g8WLYvd4ofGyCM7fgC2zR9KqAusSNs3IPNPMiGhOVmNYUAfZXLR
d/eMAj9AqOW053Yk8R5M8t+SuDWGF7pFhfSELnadmr7GfZefr/NXIZGzR8h8UT2ea59dbyXQXkCB
zzKC5YXDR8yUJgGJjn7jUWOW+dbjEyNwAczDSBWImw/0wmDJ/ZsFNiZX3kgKlddTn4gDq2h2tmMY
1GGoHCv4T3RfLZ6aISCK3vbR5bfMamHB+If4sOFQSII5PZE0jiBl5+1hqxU1rdxH7FgVMBHTUWor
7SnDqaaxGmVDCc3+HNr51qLMVD/J1ybFGLksJonnpNur9poHQDr+YZbfu4S/GXN/XViu5dt/W17T
0hkyYMggNqq2B8Ex99YXD78aPow6bqAOP4rT4tDPolp4yqJhduGbSFCX+SHYRaKejna+o8a8KXqu
7/r94c1KEU/EwOatZFjC3dJofatZBQ2ACLZMuHWi2lBJ96ZmqOgHlZQi5CoYrRO1WqMXG/9AoShp
mFGB1UxQ8QjRvHABoHnjWU1R8anacj4y2Gq0gzk8W0D5PxephabopKn7r63RwrIJHDLbIBR06gGx
nd2nHOLrPabFOFfiI+/jZfzyMzLXvmxMRXCvogU7KLBVQjVfpCx0/7OBy2Hi2uKvHTEvnZMDCxyv
yIyRLp7+tH/9YUOIBpYrIEqswwJUp2zBr2hu+w59Y7s+US/2oV66wYIzlNgLv+rXD3fKdKVjnYAY
xgwb9P0xEf9J5eol4WawcBoNbpQo14hn4jiBCzEDxVGSlfw47oLnIjmh3m8Pv0EHy1ryHN8OAVBu
oBTKgJQZdTfvLZDrRxt7svSm/MbnU1U3iexphV6PW2UooxJZ556inyZh6Fo1z5zFob1ZfhA+QOMp
EvAh7N8ogEisU+ZlfzRMVpqbuIZzv2QYH1G+RKdFJTUPih2Jzv6dO1BoXYxxTT/SL++6VQw58SG1
Pg9r9gujitGoQ8FY6emEEQv1jdHuVBQiWa9AJ5sOZ5M+9TDNuDL98udpMzI46CpjjZ7H4T6FauDW
j1nAokBb40Ry4na8QTozCQwl7/Oy/SiAcIoHhcVTKYh1c55x9XXUUbcLCZpkCdAwpFXGI3M513Fu
UGZDm3OFlzSKoWx4ymyDiSqez4vjzwslcSBmErgGKuWSrZiwi3eCTB5dX3wYJkHuXc4pefNjIckC
Z9uD1IxfWJGJojOP2/N5xIkYG9o0av8wSlzJoCiMnmsduIWEeUJlnRrS5rY6uk+ZorFAp2aW2FXe
/w4y62TJss8HtxjEBFSdKHBUqqf8Xv/uN0Gsr6Q2r7odP5RiONOiLpdtoc9fCJBJLCtEGZXjVrHd
yBFi4ftPTFG2K/Rwgbu5qLr5GvIQV7q3oco08fKqCPoEkP9ktNs83kLhedO3PQ4gnfMzk4SvpOES
PyOb0R14QnqPabiM+Uys+LEKmiT+6VqLzwClzuhSN+kcQU1Ru5CM83bU3FfZh4JciABZjEARWuAg
uqGB0HYe6A+smse+4H+Q8OreYxEyXqCegI5u8VuLYTJVmheAr6zP5z+OwZB+YnzqDAT7Qe4gedTd
TJN+xRyuwD6apIKAjYh4d1RClBMsBhGKtPa+Pl3PeqbfXQz77CpAmRu4ns9p5cuuWUkbrle7jcOV
/Is+CXIIEM2+EeJYfxFswI+olm0AVtDwvworRhA6MJ8k2ual0Y1tciTpbzt/vnoYVnCQjSMXaf/x
B2LkjJWEgcyaJPMa2byKJZrSG86Gzr2yQkY99Vlo57uuMOtglGKMJRGNVDi6LJuVkUOE5buGnj4l
yLPD3HOxm7CBffMDAJym9N5yhYPtw9fCya5iKfrfdw2oLaAQiVWHvsDMDjm/KzUSzfICYASYKDec
Yt99ML6KEyP8faKi62EGvOghFZiZN8YFE1epGbA2bp2b7QMdDmxZ3/R0Qm/2kVGJTnngTFTHQRaG
qGDFiZYf6YLzNNSCT6MjEuC0uUdS6I2sGJ87HhmthIIRDTQfqK+Aw8mzKeKbRthzA+/EuradyMQG
h1+az7VsNtnAIg9eAEirrP+MgT/Txav+RtE0RbJtLOY9V+rpKNOev5WWduytIcYXTMOA+JH9K4eD
1fa3O4d2owK7RL97qNUwEiDvJkiBXBW/czuOHbtLq9FF+2pYb6GHuQoQg4k4sYsn6BmitPAw15MN
sVK59Tqywkg0R+zB/yjhJPfbbiFWowYzP9HAC+/G5sTd5NoeVy/5W6lBiZv/s/DsLadvJZCI9i6h
jRa7+r3VvpzacClQ71rMvMyqNce9v+6qKuolZkD5ClroPtmspuWeW6c7VfHXm5Afz3B54Y6TgeY0
HmnPuIwbsCbP/yhyink1U42YvwDhSgyb9kr9+uvG5OKz+azn3TBoSzICHI+CkYhZbS/eOQGT3gP5
eWwdqWEBFKyrS+l/jeB6cySiiwz8eOJPTAAIP/uZK4bBW6k4YVglmbY+VuVLBRM6bXwLIXXsjldl
eRlcM+Y13J+TUifv3CsabbFSvQr8gunIDkt1pMZavocvymeY2ZjBKTu7zbB++WbF24ilevidG4aV
OVmvy/52bxo4XHq4FyN11zF4Gy1j9GBZI7JxSVohJNlPFu0DIwp62yOuF7SqF28gE0D1/JiQynaI
BaCcMK+W/kDAUdo8euSE2RCxYz6gr5UZFBu+f/iBfl8Mmsfhn92Icg2X1SemKC08zHeO/WqMeX4c
AYMt0x9FNjnd39c1SfbpzxW5FPQ/uvyVqQHG+sXX0eJqEDRTRboiD/NOF47MrJQYvIGjq67fj75F
tof6aIWuuvVkJIPVcFX3ifUVr3Fvh86tE39t47tXP7HbXDnUh349g1gxEW+X2Vsy+miWoDPPKjuJ
e8P9/4v7ItrIs8PxN0D3YDfjcXhs3wdtZtgD6VsKXMQmTjG9TJKBvhrOHCFGlDz17k0ZYj/lL5hn
vnbSb2ZOl0ctQNpDYLr/YdQZNEAYbflObVIH1yQ5OAEhsC7bZ4VXP+gfQBMVBvY/PG7gT9xx0dwJ
Lm21WoiFvZ0bLo+1CZ4cifx2ufXyC+Mhi1T3CnlZCqaenD1U1zbJ//EMEcmQmL4PM8nF5EYzBH2U
8ag8SdFAshPTU5rDiVSurwp1xqgN7fvxvqpOxOfLEnm5RggBJORjkzMdUd6y4bD5a1YyvO/Gb/0+
uMR1CeTydp/QFXYCUl9Xfb2EAiS1vVz19OOMvF8SoDOxg6F38nMrSc2ZK3z5FxqtcrcZc1lUTdSj
nvE5z/30WxouxaphqzCIJ/yla8AwQB33X+OV3O6/Nue9jgeHd0mlOGtAQIKOwDSJIum6i2cE+DcA
WO6QqWQjFZVmzO/sOVTUkCZj2UEbqI4/cmF0s7TE6Nhw/+JIUm391Dx4xRmrMuS/uWNGl3hzJgEN
36AcqzHYhxc7EDv7bwALHEDx9mSyYsqnPxocg+eXDmwXZI8IGBRtyEtCFRPHeBiXonpp53RBHkzq
V209vQ21/5U6vNGcSFjaLiaA7xeJzuD00iQzdgaDlct10XPtLyGBbo5iUU6vWogiAMDjhdlxpKq3
X+naZ8eoVH+B1iHhxbEmryv7q0ZPoWNAR25uqxC2v1acR0+jICUG+BblcffMLbVf3CIJ6uN6ZsSE
F2M7UuNGsGPjG+StHn+wyOER0EvxG6SWFpVAUd+fIzdz4Etfuzoqkwh80Ckw4DeNop9kBdGLJ9ha
iSZvNzgWrOB5vJVxUn4XRYtZafMgqCFM9zZEa+bTJp8z3oPFGpG1yjhDto2MMoj4Hl3dHpYGS+hM
5bY/rPvdKVtSERX/lFPUenVKi3Dc5yH4kzhGUNyLML8aFQ46pITmmr0UKDYHqOMGVI3SB19ujzOA
7eXMb97q28BvFIUk54CUQEAnvmXUQQ210pn6nJZJz9oim69KQPd4GRSQ5m1XD2fgxASdWrxJ0Z5P
by0nMOnh5pkFCNbMM+vnzZlmL1rWw/Nl8ARZrp6QP06oiwWPI6Fs+dSLCHO2uh2MI4uZDIA+yEwC
0d/1a4MrTDZ+Zr15BBuHI9ATGtkA3mC5yFOB1yiIpXADNaFY0jo0hUkzaq68Mv/6xe0ffANHyqxT
GbPfc+LaPP9FVB9DUK/smhj1cfqvC+5E/HgCoTyLADD8yofjJ56fWktrxwUDiPIG8r0R0ojQfTld
lJHB15aqbQCe6W71LliP94LD2NSPUftB661Sqr4Lmd/pgAHpFs+6zJL2+VhP1FdXrgTOtZxziC9E
QtDKBmRNORjTHS8xYHwXBmFSDmGVq+1NWETv1FRaUKbWdVuiwNWF2Dhxd7l5h2pECtHZdxrHwICb
1LQUcR9M9xaN186jby3HjQM/IGI4AJazfXUI6syEcjgt+5RVBfFlkz6FLXawBcYQe8cABzC4nDOJ
WogEGZEjeQCd2+lo9ob6YE4KCIECR4+Kd+JZfxrTsoS1SBDqxDEg0H28S15udozy6kx9bcg07cIJ
xmb3cHfVeZ5pRKCoBB6zi2ptoddxtuuqTQijI6yKMUE2zz8gHAwD5RJnb0rdRCzHWcHTMGUiYk0m
p/aW62/Vp70PSJ1jdBiKX17zfC36wPylNC440FKqMxgPhkZFn05NaM5TfMpOjeyGUaTNX21KPzn7
TuX+qpMPXYmkJpt+JWoTQaU7pwY7sAY1pa0wZjIN6gvpNMPTOO2C075cu69vyQIKYV5/QHEm4RCX
Lno9GsCDE9vxEFHzeeo8Tnv4wSZqlPPHHKHBIpH6ae10DKFtF9dHWYJMqCYgrW0hGwIqzqRt9ySJ
200SbIy5bJw8YM+nntOAjd9oVqrTa7QYolZve8SDkqpNmMWpByCGK9i8TUF1ykJXA3yLF4d6qduU
jdNxRKqoYkKA5UZVMNIywXQxY/7ALfGTr9yhaf0bS7FbyofjwnBUtpx3k9utdNew8Zz6BRLoT2Mv
utyKIF7ZMYYNHv44/trs35LTee15xyNWVXj+/H1zudLj0wewNy9tOxedH3y7dLWpCzKOW5bo+v/d
V9AiyUkQQXV3/ajerk8ERiD6s+zbzH0XPSphFrRz3DC1PcSC6LJmXEKWBLiI2bgabhPzCKoaT+/T
6KDzmzS8D/xpJFPSY26DYcnMdI47oxuIVRwyU2XMlcTyiqUuXHBZhKf4eG9d/OSP7j6PrBXOQAXa
4DBUoIw6MxuYYywXNGX0Zq9RV5zGh5TOOh5+GqvO1hLIbiki5aEBE4Pr7/ittjZ5RA4NrSkyDKR7
bQouO2q976X2Zkph1923uTVXwzwj6qUPidnxZHPUCtoL5YOCO6DBX+8gyfH+TKfXFSEPHmEB4rRj
2d3Ekw5w+6j1yRGzhoi6zYexSuaWABk/u1g3IlxtBZBhMhvae6aa6YoiY3VsqGAyedDvCqtTI5Na
rCUI63hOFtvQfdX5o3nXVMKuZuLdltJDIoBczSI4c1aSed8GmaWOZBpIJzrxe598YYTA7x8YY8XS
KHIxHVRpMYktu0EkKcy/bDx4jHKwIFYHXi+5pcnHcrr/e4D1dmMHObxF5/gy7wyKkfvisjS9vcdv
KV5CmHDnfk39H24B3/2EYoH6zdWLtqI7EGpiDG7N9b2/oSMEhglsy7mTQuXkQnEjaYjLWFpL3j19
r3JhmdioekEG8wx0HGJxJXwA7nwDLHDZMZFGY/2UOYMjvg1C4hNKV9iJr1zVXSosSmWrRkb4SbYe
LG2qKY6ynAnlYfaflVFbX6+TolcZTl0y40n7s2f2YSrX4rv/apOo4uc+tpMKIzSpoT5oo9xMiBlo
1mOZZvYlB8DUavZPHH5IROzA158fDFc3sMj/f0PMwTSb7kgrGBSpNq1hZRtjIasUnB8ohoO9Y3ma
DdaYVyxrL0RgBQlXeBV/wejKikBNtQvpO+79uiR6qOk77Fk4El3L2CRfnPzxG0r5tDM7OXycr4t2
2Eu2HD1zCcc+aFf6JFdpu8HD+q708SO2Nv1EjN7pafOE2V9mjmVjLUel4ZvXk+L/CJrNp6RhMR+W
Hck/16ENL059KEoSIdvice2iJiGf885lnAJU4O0qqlJ4AM88wjCFwZ5eKLMsRf/0mdkYmCzJnZwc
xqFGbgtqf3CdklE9T4O9wOqUxQ1GHdDTiQoeID0037pWWNjAFbr2QPW2noAMsimcEpmP6+esN81a
13i6QAWS2OYbz2Ui/TWDmwkPZIADSglHY3ymlB1uASDl+ccbhbQ/s0gYjIOh07RhvjcdgY++LSSC
TNlfXfoJs4G9bADLZwtRiPMzeSsJX4DVJg2Yjf4wTGA4W18X9uYcDmyh8yKabpxEeAtJ871A9OBY
cpqM7p7LtytYh/Ho7yN8KxdnOyKM6SetbcFbXbK44WBOOmxLcQZsRRl7PV+xq41j5Gk2/9dl33bg
zfe8xVBDmZtLBIOOgunHPgbVJ8oMDm+yQQ+gwQBspPzHKBAESXEoO4qYWQYFAYspKJfhudBy7Abf
SWqy8xoGLqMwdHdlxPvB3Fdd69R3asf6PfRuDKFUsD7aOhWQs0L06m/oJV1BzIbVkDlr/KCDspea
1ADba1Hb4SBmlIgOTxwBFDrpj/00T3Vcp/9GmFz3CaXrYjG66VjfCnZTTfKnbL+l0mAIHa2MXkWl
HevfrGoRXT5sUqXFTnyyL114DBE9GHuHf1JYoTTkip88ChIJunvlGvGtp4mP8Z7v50i6O81wkJ6H
OOGS1+Xzn1aCX52ADPbzAHlrJR34yNpYs5ArFzg649wz9ZZi3so5NfDGLclvCcwhIf7cCCyUkYX+
md1bcJezbrqU4PeKStOQ4RqY3Ck4c3kH4y582Qrc37tNe9Awpk3vpuGc8QI93A633rULkHhH/EfQ
7VT6/aM0BvmLFZOQgTisA4ujUuXvactMjYsPRtZ/IMt404S59ddNC+G6fXaRHeSvy8zx5GUUQek1
IzeRAmPfpeoKnzX6zkGbxocW24zouJfY18XozuBmecFOI/jPX2wp18RzVNa2kjqsmWA5h6FVy5dg
w1cUQjgvFAJSHsl0uMI0WanHxqyDhQaKf41zQSSE2rKChUxeKylKaKNO6f/377oZd2bUNd/PydlE
sGx+yPQwwcwjB4w14jnEwQc6ZyRi6FDx7ydF1YMPnWgynnUr8dJ4xnxrdgvXWdsBTWvCHCO9ERF6
yDyKOrzteR1aXflaFH0cYqqNntxILA5ho62dMlRydsLSyDDCnwCefF87wFv1YGZ4/9JgvvsdbmEz
e+JZajnPxRD53HTxWkO1HYUpXeXbX44IkyQ0c4+TU/lXI+SF96RdTX+pxozoOYqIf4Aj5gVwCD47
/vr93Os1SkXEZnQPEIP47O2Zt2nDUnG438ESVGncndmGlERCzbLFgZNmw7JGnVLcywKe1s3HYilo
MZjYvFIWFb3dbAJXiVSbkHuFkXpCkTPyGh4SfbJBVLqswCPngp+ULPItOE5s2fR6YvFXQuynBmuS
laeAlNeGwh3h2y76gPbwR0htu+fBPQvJ61Q+NVLivjYe3Y+aagadUVYER4beQrm9Dted8l1hpl/k
0vYU+5XJQRRMr2ecJ9egdf5XDdLf8ptDWiggpkA/+KraoA4DqjADDxUzrk2GK308bbW+l0Z/mz75
ktJ3crdKzwHHjm0mFrl+7+tXrWmH7DqbZE9NdRCS1mVA+kTpq+2zUp8CNAMFjelWsY5Ln61ojQzq
WlyuaJSukSfqzt/em7KIf3pL+HfniongTAsXocn4p7ABXmmqBF44vbL2gqUEv1E2vpISSI/urMPQ
Iq24Rfb0ISV2W6bhKX/+ETZWFHoWZ0I31bdMrURW/u+0ITOMyVrq64n60Af3io5gryD705FtykyZ
DqWp9uCQ16h4hZyYGvPbfUenR6pDijQsInPZC9wrGsOb2dQ4P9eAv4RXuuhJcZOsI3F96dplefl4
cAf7nY8iFhQtTuE3ZByLbIrAtmvkbvDF4IUtnuGpCQ4EAST1zIqfkwWsgJvv2BejUZfwGjUcvKY1
3yX5Ziqe5wWqPi+Lj1kj6vGfd8taKlo1GM2gd41xUD6dz+bzlvodc83CZv1LASNs41m8VM/tyJzz
kOME8JsYfRxSjcUpAceE+a+CBtOCjhaiSe2fdbY7I2cb9gjZrl87ggUhGLW/29xqb8ParBtJmnuy
L1d02TPXdALLNcENt2Qbc3MoUNL7KYposMjz74hdqaAOzH06fYkC/hIIbEQ2YAx4VhH/PYSZ6/En
GD7pb1+h9m5n15ss/98pUgfaFX6v0T4pvG0lHbiPLXas9eaAKzGgMAuR8Xt+XoawHvQriuf18qRN
EZWKkCB7D4oNClwq7z7qlCTNMABAqdfU88377b6jLUmCLiJzWhSU91fnx3MVfKazjGWXaIYojfLR
zKg0hrcAUJ8odzrH4IAuogKEA0O65DlNpDRlvYzN+YExHMum+IzN3yTtgwdEiCGSxsXKyLGK22Vd
lzilDBKgu9uGSu9YiAVw4H3rLMPbZzJEmB6BIcrJy4yy0/xKiURBJc90oxHEyykgrjfhHlnKLPPl
I/bhybnyp+VL13bOT5Sd0v6gZeF0Sq8hdQjvbQWJqsHZqEQgYryBu+uQHA4wni04sHbpKakgryuv
1i4hfaieS33mY7W0KzlP4GsJehLX0C14ggb4NZkN6HiShXNpo2qXu7iR1Oe9+nEJ3FpGunk9yfCE
YVml1FMy8qbd6DuXcOH6g3oWp/AQtAJd3LaI5g1J4+KUhREpeutZJpCz6YXTWTa4JqfS4HcRySx9
tQ8PSWfllNlBRirUdManQlq2aRsAXABzWRSLnbOsNCoSkR/ds9kPosYqr9vPJIZHtRyv7kGm9ZHq
gGDCgDqDbwbJb03Mb4nsSEcTFib0ocyV7rwML6GpYMhxGeuJIxQuq3GiL3LiuF2Mnqqu1jgQ4fug
OK61cuKo4YS/xw4EQViLg/CtOToObvtICY8xko5VxwhW/2xQztqrMM4kRrmlHOjfsN+CK8ffcMh+
ctgmstDi60STIK2YyGYChYQOf82AgtRutEqVRRaImQGJAJJGzp37rt/XgSXkOsxTQWSK/A7t2heN
nLGvweTlPrf8Xh5vOVpd5ofiMcYLpctR7XL45SsCVYaBk160q/nKU1aP9OxYDbjnSTfYr+rdnU9R
SDrQql2sJDC5dDAiIIo4/84DPaRaHjJOf60l0W4dOt4zgEpO53q56tlj4tQ7eqxXnoo/7Fe3gBnf
EyCtYEwdjew/nwaj1HWo6SmcjR2cGz2+9EK1s/jgkxeES2+HRzgSULh7+iy7Zf2odb1A8CQM5nes
GZ1DEezvprLITyvN1jo2ROF1/cu2+GeoJxvCD+rGRs5N3Zi8OAZaCckmzrpHHn3GYYre66Fj6W5Y
+Txec+cDw1SAP2aZeq9Hax8WICvKl99pA457KBC5dEJMjtYawPffjPDoHHxUSak6cnR42lkano87
AMxQ1N5WghN1xQwRaBjV8QvBC2hFVEV0S/P2YXfbIvIdCTY16bS7GxHyzrv6JlsnvGqpECdI1RnK
bxh2BfKuldEPqRi6z0l/0dcz8v6AxRkrHAwCPcqkKtD/TRs1czofZu4cwQNGXferdRpTbrivk7wx
YYTXptk4OgKuYy7C3HxAnXgirIlh13r790azgQrP2dtomy/3fCB/sEjnRanrWhIlRljxgYwrD6ia
G2uPgIlbk2Q6Zl7IYoUlIhporKv1pJvcRiuXVARUY/JfVP8OEfxEczGZufwEki5BBvfyb5l/eVSW
It7c695Tbm1Dl259DXM8Wnorng9y3w+dZHD1nJJhOZDcuAMImdhDbdfWxUjciNoJeswri9cd77IV
e6QnwO7wYuWknkTwKw0+2z4F1s6tCC+A3YetSs+9WksbrDYDujt9P/A1jy2/4GpUzkNVLC4PU/3b
YlBB++o3FzWWgJNtX//EgS0hDwph5cNxauJm9fnMeydHtokUlYDgzd3d75A1JlPxLpP0hQTP39ET
5SVIiwoPkX9RBLowXwgiv3tRZ1DeUJ3lavfdN0ieHMpsWFBso+CCpEIHg1Yqr2cxSb343tCyLu+0
HGswBYK5mpmlPP5gduVMom/CdF5P966SnUMcKFf5+4NhCRPRiBW7OCdgEcNEHTa4wAgBUTGGlivX
8t0TWJc11zrt4grIBAKwMZtzIDyw70e1cL+9w6vgDGj1D+dey2fQM/nG6e9Fj0wf3f6BiumMQRsH
56KyCKt+yVhCUFrxTCw2paHHJV9sVigugUIISSJfUR+gVd98uxmaOTY/Q2L2g21XAIKojy8CoEgT
5wlRQUxPIk4iY3lPx6Mm3DIqh6MAI1DTlo28vzgeJzTpop3mfVpjkQZQYSIdql3O3o/UY161g+te
GBvm70pZP6WblHw7MevYG3AMEEk2D3SDLTCPNGd2DYKYb64daX358QG6y17LUnwiSd7f1R01AzK0
jdFf3JUunohWtmx6rUqKrzOms0wUrKTCL4JWBb8dFDYGp2WPnPZWUyQnSk/YCqVEooUeT6wicqWv
GCGyaKohGbFn1VgQ4XWX/0xUGSkzkxhbj6GCDy/kwWZEWDj1K/InuaZh9+x4CkFKS9VZBnbDhLwr
iJDtnJ1rfh6KB1+I5rIO2gqIybBpJdkTOoSASGKWXO0upxXscTj83De8P2vOT7uPX11q7IHQg66d
KswOHaOfOKW5NboI4jA9I6EbscgZP5TApF8MGad5L3A5L7I8QfwAJS6pyWSoHm70/DAqjjinwDl3
CU9a+/JqqaGeAgRQkgA1NYmHpmz66IcESFcoBh/xs/aPwMfc39sx9DCM0e7spwtkEE6jSk+KIv0E
QhEyE4PxLlN0AKvGEAiNDTd8ca89a8nGpldDpAqhaYXzchmLMv7lH6yKcQLv7VatwGdpRVtUkOhm
y/ZYIDGzcMI50M86W2RPl7CektjNpxX/OlrO//KBez5AUaTVNheEI82xpSCi6BOyNDiMEAeE5/re
wsenA4UukIxeSHtIK6hiIZd3nKZYp0y58QNKNPw1lquQVYvgdH8afmjhVjXPJw0IE/ALDE9C77VG
q41X0LbbRXCsg9qIcbsQsyjCbGuA7yfC70YfbPbDe6RDO2Yo/EcCWfvvyGBDFMpRpIbY1AH2e08/
0L15JmHJS/7ZhQvcMTRPuaNqp/tEVn/wqt72UKUlfU/8XG1sIDKIsANbJiY62jz31ntnqfknsdWM
v43YSVNYaX6tgzYKyU9OyWxyVC1ZOEjLYV3WJ0uWNZoZMbT1b7OFoklnpU3TPbm6e9Uzd0DvOSXi
299Dg1cmRGY5B8mMXkj708SuCypZ6cmFp5PD2+JAA0JMsLZQXfXmFEc+/jsECpmSf0SXXUqygtI5
PeMLibAdkFWFnwWkAUvDA1TR+a7XiF6EOVtjXs1ml+Tj2JwD0SEMdNg1b3186i/TzsPMGuy7Qg3w
jq+0VIi6TckO7aBaG7Ol/Vnv/ks7t7vVH+67Hekvc1DBAoS9olMYWTVDz3pBJBlHqK+9z/j9Mo/M
0DJzGKZUijqXa9HKoFA+088zsB/gATc17MOo5xK6q3bb+2UJ/dFJEYajqsK2eyxyiaPhLkqY/XGv
ufCsGcAT0o2A+Rl1YiT7x6g7W4fSmCzDhMc2RUZ64YNjsUwtAXrn0n59+XNhaahjqL3osTGFOraq
nBwLbCSjch/LLTLnJ9v/AZIf8KTsRniekqTsDMmSGpJChcDHuW9Qwcdaknk0Bgzrf7BuplX7D/2V
LKF05j3fRkI6VDYHv6IWZs2OmcDckZjbqL+ylY1D/80dzBvyqX8sKC4sW/DuBQV+8qly90kO20/I
ptOoN8XNencrRgBmhKWz7reCeTiOEtewjD5mS44db0vuSGvKcjA2QUK30jMQLdavdG2RjQkEPBTa
MdEGYKTfrcAyh/uuw83Bqx/ZaWkdeoS+CeNvqrRnoaNfTjYkb3qbkHAQS0iBzOcDRi0hJt1Jw30E
5yEUZNsVfvSdw5WG1sHJjiOPbSSN0Ye8iVtVDc/ppA4uuli+wKH3q9vO3fzThTxH2sVaqFVNUXMl
7YAeUo1LUokGHvzjlfyJrjij+AtvWJief+KpcqERxWrrWKPDXzkLKHMZSxh4ZeDpL8taQZRNmKRq
XCt9NM/bo5rJEXoETC/ZHYTmBQl18DwLOsm+Jlxc1beV3wrCz0dcSjAkCVDR7Le2qBK9sR5cGUHf
27Ny+t5qDQfw27wTFG1seGCvt+ZdVujFRtOOUgvmQffrJ7g21BOFXNgOhK8WjecJjm5C0MLqyZxu
WyaKqyCex1oJksEyN48WUClZHPyctyUa1/0R0fWLtzFRFTd6/A6bvV13rwqNaNC8fq24miEO9oLq
jqdQtVvLBUJy5tto52ChRUQkU7Xa6x8uHGfkVMY7yLkXZ645cxg+3vwF+WssUgReuqJXbzJIXOfW
O7N+nm6mte2rpZGFFyAmxgy7jwAQmh86jEXRcNFW1/+EItpnxz5Eec8aNMM6S0d5AJ2oOAV6WbbT
vpYlyFE6cOZURzrgCaKjYgmio/NT20MTkBv03QINkTQsdpK0tbozoVw8z1mvY3IzHwGqRqXR9mFh
2npf7PQjP2VoZUccNeeIZwbMSJlLRkwTZ/CuAsxAejVzk0nZ6k8Qi6HaSb817EXgQHEyLPdYCoDb
vPsGgf+tLXjbNzt+Y0QwbLw0nYaCnVuweXSC8BZpi78bdIJ0mk621gigBjQksJZYSx1ImoHVjcpe
qig2zrD/HvMQIG5dueb1hZPiBxvVqvTb3cJ/s5y0pChRV00h/+2ZHkXP0iCnrJOygXfB/6htdDtH
1fmM2jH06LQB3pVqjF/yZT5PmvHEQeHc48LEpLb+XFifgCTw9kAJUdzw6vvR1bmS93bTwNk6Iasa
8RNhHOeq2yHGFXPuxvMrmr+TtE68QFuGltGmL7oje+VGBAI/+XFB1Tv0t1O/dXP9xKO/cVz+g+KY
dpwujIVJccd9lIA4mgy1rAPSPKEr1JX/5cBISk68RZMkEbeDCY18J2OMd4GRkEL2e7kumEoSSNpy
y+gHgtZUSdI9ACaRnahrqh0Sg/x0QYOFXCSLJjPV7nEtmYsB5zTaLjD+N+TdpjfSJEAVb164pvJi
etqbVli/JtvSWXTSMNcM7J5+hXkuS3t3XWxsoQuoEr5NtlP9XYsoOuCHjtksW7wVi+AUwX6RPmgp
dEUQnksYBTWByL0dVqj2xSGXYI15DgEJQvE/oGwOlpJxwAtyW+Lyy8mgRvaDhmPDRUrM8aOIlD9I
gXXknGzcC9CI10dZQ2r2GRkZ3PEOV9o8/qpHkQHi+6vxqhG93l4uMHv4qEA9vtT/WYPdXU4KufXR
WH5n3n3otFUl8mKLtXuhMkX8hF+299Gr01D4ubqgER+j7cG4dx40RODuL8EZJB/HfMld4xEmu7NC
a2GwDrqQ8aqe+goGLgcWMtu4ACSHFg2q0iEmOARUm3mCQ0UlTkrGNs3ZmuYpE2qcLe02xVAMlCsR
EnBVwjqkZZxPFX6MGuLO3OtFZIzxc+JaKQIeoKpNpNFIFZbucCYIE2n759vYwiUUY1P+0b4/br6j
PUsEgTduNIGbuiU8ixfrNhaPrJolAaZUeYKpkbnwtZoEhNBBGwS/Hkme/ich7FbCdH0FRzcea+jL
YplufaroomvT59YKpothYNWR9IAw3Ih5DMCZ/v7Hr3aKtBwhCDYqyxtGrrxUhAgey2FjJuoFTt8b
4pfYofzM8qQMKNcITJ2bu0mo/HXxxSHGnCAKX9hqMjx2Uj/FPFAjgxYJfdNrkD+Ff9b33Pg1HLI8
CP3g8VV/gQtD3Ub9iL7E9U+GgUYWSh1+6Ud//U2O9TbZDPn/rbCt3+Y3KjRylQj2NsArSBIKiN90
Mi6ktOr/N6MmAVL28kMZb9wpGuD+4ll29WOZ+gjTvwwSbPrPBBpYqkG7Y2mROpUT5JSFyTMHUsh5
0ogGJDV51+C72gnNPGuEIUCHwuurDVaGSrPFIgjXBSZniLJKR19RitZ5nn5upbcBNjyEB/RBydgQ
3yz5KmCrmq9eG6hcRQBsZ5N3ko7I5mLaSmlQ8t6ugVtrxZ7L0I6WJqvNjIQr1f7sHdNOOo7dmlxN
bxFLWITgaT+RrA+MDUeLZx/9MHpUbpI8EShW0l3Efyde/fI/dSylRmyqmAIPtEBkc/eygZLyfcNK
7ZJmQ1Y+6osxSPIhX//hMCeIgqNhCbw9xGgCN0eBdHbooeESoQ5NyCa3mOGBbVqerXKmH8RNqBsH
eSHxCObibSCHFi84TIS541WKl+lIzlSqCeBNHmQZB1yezEQVlWu7cF0/ccDNCTt00x+nsr8/V4cE
PDs467QzTUqQ/FA40qprKzXsHUr9iET1EBGbGpmDq0HZXaRoxyfmeB+WFUFzItFa2Je/l7f3eMRJ
rBJL8eyxRf/kOrs8YC7vbzyhfycRH166nPH+jAh9HdPo0d6FgZUuH9hb+4MxULyDITDSvRBp/ez/
hl/iPrcx6jSdC1DgE23hfv2oJ78eH6/qnaOIXHQt+n8pm/MofxxolpuRBOm8z4K4x7VI+Fd/YRdh
yJ/oLMHRrB5MN/cHZwYaJ/L6xbrquKQWVM0OIHFn/0lj3DLMVqVbziztZYs0EzAaAYNjrr4k0VlY
AXe1PT5ky8wnpq4B22an1S+1kJPVIJYRIwg/06+L65jjzu9yWh8g3ATyboJkckJOh1LSgkn2fKdz
NVIOAQ8GEKBxHVvJpgl8gK41ZijlbnxnhmFOUcIjzwKonoczu7A+gppE2zbBkeE3fWIqq/AUGXCy
tReHKVo2pKf1bdS+R1HCF1FqBkoEk62ms43mkyJQmc6fPUceqwrprWigmb6fVeWwNqIEBpwa8cDJ
gI6Dh9+awV1M/5A0k1w1bxBhKt7PExHDFbqTNtuWOU69dHowCVYHOnJcS5KQ7Jj/lEVr7eVFSdyy
S0H+ETd7uJisQNsetbyauFbbiqPtOyR7TIIbik/PTw3+EKPrxb5ULklGGJjhO9MHhmW+sgWB+eoU
etbe3k/5+988KqSpJIcQZJSu45TrCADFqpVzW1XIdSlA+rWKTnOzKsphjOq6U9q0qTCKdzvgU862
nkm5J+OV/hAroWHLQVzcDm9J03ySw/pIJte2m2O8/GekZIYpFDtEeVaBh151Q3xAH6xwZEgnXAoF
/a85A+UrT7DFzWuGcWDYphGD5XOOvOFuCpV+cCg2QW948jTFGwp8VmS7ipj6s1JqJ2CIfBb2ZJ7P
s3tDxLPwP1CRzXvOJY+C9EBd70pzmx+EaCHJsr0iEOUx29yZDGneQcMEwNeCKKpfdA3RMTJjvCta
odx0vRwR12+YP5f1ZTX9ZzUWN/kcBa+Wjs3kOX5ZSdxc5Dj/WbK2t1uQ9eT5L5u+uNkqv0+oAb47
xYYUgBKF7XDF3UcLhLmKdnntlbHr00SYiR7Enl4gty5xOVolFqqTqyfaeKNqpefLYVjKJoACBNAi
HbcF7ezR/xo7gO9LoYCxE50Ah/5qZj90W7rmBgnN/dCr3TGKDHLhZBC8Yl/gtSUzs+6zEasFtX6P
msKBAUBa1wnsXKELGsDmHyml8peeFrPbeyosmu1UcsK5wZM3IFQhD8fEf/rxYQnDKARcOHtvMpgr
Shb+Q8uFKR1ceMohoPc1qODP00WH09b45SvMue/bwGmdI6w+xJN6S50Cs2F3PZoCSlOjXNMCU33+
5yv4n5qYtwAzhDBcJb6DropGOLpXENiWPfNytBXM6RSk8AmreI3m6Hp3XZHwLPc9oQguOIm9KkYS
iU2899MITS5DdHcoM1g138EYdeBXGT55Vj7jmb5L0gK7yFkzKOGMklIJTKoCVyUU0hNdJZwXKmUU
cOY67+vbbKQLeG1XXjZ3sZRD7wxBoTuvXhfC7VW/5lNpNFSsaWgFeTejZy41DbDYClX5hb29x1i7
6zCFbOY1CsOhQcs7eENur5TOmFxAkjuBLIwz8rnEuZT5r1CRJiNu3ushv05p5oIam3065/3Vwts8
DNR0oDoINIh0d7cmJQZHJbK/2jpSbn9lp7P6WDdpV97BQVHaNG9Xbs2H+i8jGAzIBCuznzhKChq2
Tv4G1hX1RbQ4z4MxIeJeu6euGKWHBPdzYwDpKePRsk9EgEwn0LIj+j0o/tuXXLdHRbn9Yp+p6RII
ORaogD2Nm91/0JCgjfLggr6mq80m4MUpMov45kNKI3xyU2Dsks0mkBEazLpgnG05KM60TMQGuBkQ
lY13XRTjcYm5c9MEihPCwVo+eb4ODPeYHR64Yjnk/Mgwh5rZ4xeYaCVU/ftWrbivBsaf6jh2Ytmi
1aQMlt4zAXVZ7Ozrg9okJpedg01jv2iL4l8rmK3VAKZ3EbCxMMXBm0jV613jOLMQDMzwvwc97qzj
cGjSDFGhw4X8W7oF1KCSROuqJyExZRzQo33ZRTaKf6U/w8R/l1/zPaQROG1XWTUHAtKSmlJKZ7if
g2cN0bKnOMD7ovgzv5qYISGZR0GIFcLhFcz6oeyz9FUGU8YDQnezb0RKlTnXboKsdSSwvHv4f/HA
GeYVp/ZptxPbmSqia2d4fpUymumqgnP0fXwK3XhI64E+i7BqeCuDjuRzWlh4bBqbD5DRsrlGRw//
5tz8zYZQNk3dSHxHILvyx3lBYHSkFYbWv+knW3mhglBUlU05QTO59Ylq0eM2O+uE6xMkAWbZSOSE
ptVxsadnL9otqkT+Ccj5yzyQG/yNN6bFJRU1f3pBZ4K7fQT3gHQoZuHyEM4SHlzETvUAk2HWwgdo
qUs++e2tWnPKAMDx3Qa6D07mlJbnwIC7/yW2NVmw1pfIx+56RW1KirXyTERq0m1NJMSMqzIvc2oA
Z4HcSTlu8vWYKT2zgU8xdjdkiFB6z40aiAGuDDvTHssg2BQ5iLatoTXFpnY17zFqxd+kSKlsL8Te
AQ19jRJ5rTp/Z5JxIqxt/nqqnmFNzNDIDYvBLcRgmIltu+UNZp/V2DAb4hru4TEM9N5WtX5j8cvk
T5wzTy/53aV/2wTvZ5V15WSedfGqXLQd3c7wTV4fD/SBxfQfJS/BZ6VP0U/OxUrT7aEPlBo55Gz2
E9boYSrE1bFsityvIjE6/xGNxd5Bx1ub0d6smwbvQ43+15S0LnSungo6/Y8JPrQp9UcGCIldZZYf
pyQ4fNSzgLDi13OB7Zk02HXFKrkv83BH4UU2oHRqAZhynGiZ1BV+HK8a/85mS8q/farvaKBWscFn
ncw4Vou24hi4EBPOJkl1oIGCuUyaflq0TQ/hdvbrRprajtGAPNBAvYppukt1xSr9hfeHu0ayBdzl
dmOiPDxC1tysOfWHTxEoOrRXvOgrikEn1yl1n7HXNU5wEEJXH13cVNiu4ufjpm5VuISNNJmZBW8/
AKlCtCJMZeKJwaCUsI/4AVuzFrfdNnqrPaUzGxxUVZrsD1vPdAkz5yu4GkZMyUn3gsnbf9V1+907
JrOgCPcW3Jbx59//WP5893IWcsG9wNbjMFzboGTfPka1iaAq4jODAJqZ5bZVc7QqrhGPRBMmfQZs
DNq50Jk1fLGXKddUcUiEs6jYwc8Ab95x4/l/JqE8SIX3Jo0YwXNaae5mj1mgxQPkgMtIb+BV7rST
TUhiosPyO2vr6QgmXHp+QK4ya+nXShQbUbG9lEhqK3IbpGf85l3eGueyh3s/sLELVcKm1Khd4n6L
3+74rwNny5ciI8A9Ec+hWQgrOw7nFytGAkaiB/sOohObVWfFv3rjcT/wXSsDEhBXXvH6HYzqXhFt
KLVx4Ow1K1KIMxnrQEwcBaOLUiTtJataBRZKdf9x0pF/+qbTtRtEdQg5+aecp+/gCLbLFteSR62l
7kCZ8ZfiQR62791hV0gaZiYHbUHU3oHqouSNtq/RVk3Zr308J+QJ4J/nQswfaHgxw2FQ1Bth2Gym
WxoASVaAA+3BCvbNp0vagKtHucWLTNkzXeUFKyzj+b+faSNbU1iQ5OOGNYkMg+QGGqhgDsZTPf76
EX0sHpCjVQx/QH8t9kaznz6zRy+UFOz0wipgJwM0zxyWJ4Jc+/E0p0IO3vXtoLnNek1U21nXSCb4
2wzyD+WgBVFIk/Oad6/c2LrYq4AHRLeWfB8xZN+1iuF92zbe+t45TKVOh+9WpEw05eaCvmL6jtsc
7OyYk363xWSR+6wR/A02hGCy3CN4dYRE3L6L8uUx/SKm1/yZ3UOptAqUga3v64VcI9BHjgkm/wqj
aPWhWnIKcEHF4e08meAnfp2kjv6+XeBx2l394RQzRJEc3jwcnCe6pknLYb1u1oBBRp6newAUVtRa
25/NVa9QS4jGMN7TVaiqCCt375coWKWeDroZl4L88y5QTsFZMUAk3YoilZdYJ22N6hUzT0fHEWmG
tSgfzaBAn9CqnIySF3VnOwO8PF60E7dhCDZPX0nDU5Qa+LYIEO8H8A89LDQomMiKjO/Lj95P4lE7
Gl7/tjfskeZ0ymWywZtMWyIb5DBMxvuAuPEOymqo+TBteTdqMxtFjHtVimob+8JlXCjXU1jkpZhw
IbUuvMGiAOkGT8RvO2MDiXksyNWew6C723SNHzdZ/ktJToP2b5KCu9Fq3qh6K2/oMlRBJbqawapu
euA3SBFNmnSzd3cFIawLPG5x6BOYNHvkvlM1k3qPetXYY+nDltjo3XPSSsjrKhlJpQgBOsx154FL
EiHF5LAb2iIlwP/jdZPDiSEsV5/UR8L+7hPl4TxtvgZ5oQQq5pk1AJ0AAEvWo5HCZQOtwvDOfDzl
jXfoRAEhqNLBIeCFmnrRZ51BE1khWOvTiWb/C+LAeBlgT2iI3l0AalE3P1Alshlc5DDJt43iP2or
Bdw/JRc0BNZdlt9Vw+s+cqraBFsS1IipYcGHDXK0m00hfNDgUaTTzFiy7mF3psGkeKNBMPGljYIB
MSL19di1zIYiLDwciGlDWpHLgHWAi8EM9EkTCW+LR57UWlmkQGjhGloQckEzce4qZHhOpi9X78XG
LPSRPCFCLY2ATCz5SVwsHLZmHyaxDVK8NG3eJlO3gi165W4MJ6J7Z716Z3X7nRGgwQWM5YryvLJk
buQ+hSiIo74OzodcYokh418ku2J37pJZSXO7bUk8GVYKWjDT860j04PMemlgCKX1YFqCD1Kp1lNX
MZS2pFwb1SCutPL4R71m7s7CWu6whX/ycBKqXUi1zUC1wyvv2wItjel4+vnzCWl9F455Y/FuYuyH
K00o5bx1q+vY5PSixaiwwGsIugrE41FAwpyDNHwDMk7di/UZa+vdsC73BCgMNBQ9xGyvPBl9Nu5f
kgUQVMyxtHqFgrptgWjAoAoQYKcEZZOt7XmV8Hf71oXoqfpkILwisfX4iXQY2dQLTe5aQWyQWRJG
rkWkNH6PecRYemDpyRQxQWEWgHj1afj/sf+7oAP0wVHjd/enG4pHM70XFBj/pUQnR/7VaOQBkW4o
M6lg158DjKTjpL7fg2arlNB+xYQB6fAOPzJAsR1sOJSUU2lIMUvt7ck+pVA8uWbR+4OVMxmjEoQ5
QNQ/mCyfkAfsXxCx1cPAzflqun4IYNEFO/OgSGS5zFhE4aGFc7aXy9u1+OvAfNB7XlgJscHnl9mi
YFFw0J5Sg8xYBRlx0HFHztqy/jejK3s2fWlIsZLxeHaRfaFsuE7KeGpWW9O/xWUQX+wtsfA+he/5
YjIbbu8wx9Q5lOgNL0E83mn/n90SwkoyVsy9phmvfI6MXuWWnZdJ4ddJk9gH8b1LanpLtkvR7q0n
Bqzy96cJxet0qbknk/46IfG25QzjY3A6Owogb8c3QalT4pB8JRLnculcdOK2XGR3HnlBvfMaYvWc
ezBfpqwPKZ4bDHX+NFXdC9gkUdSgxP52WMaftTeyOV/VnJ0xCsNX5iF9viRjdAqHLtT2upYgBepa
6CH7/JG/BVcvV9LhbgeslUzGfURqQDKHZ3+7sK8zvtyQExEegKTTpiism13OGF41IpoH2MP4MYTg
S/HwoByfYlkm50As+X/SWfwKk2EWJG3D0nVYOkZ8WGCJV9ZS3De0uUZLSwQ8SXgvhzFIRCry1z3K
s1/dGrp7fTbvc5Y/LEm1ih87+1Y6iA2Lpy1HPJ5u4Ha7p+72ZJxzCSBJlKYmPMrl80W9a5X4ubx+
Qbip5qzoSRVRYf8GtwcDrV2qQ5FArXsLQSBY+1FG04Y4o6E82rkb7uuTPz/32T0Idn9urSJeSRVx
/ZioAtfMM6H8wEkTJs7RMNdepU+ePq9ZXB6nQCbIZp2YrrDVAfmLilJ9gmWckp5nDaOhoqRMwQwR
pqRIWDYGOS9Mr56Xe3yQpDAea5a39JDfPkwYcOE0AgnF+4L/sUg66ll912vu5X9MoAiYmiRdlLnq
gCnSfairht6s5acLm9SuneCZbEQSgSVfXmGaCZ03Ufs9GGDQ6WpnZvRyxOP0RV9LnLB/jhgzJ9qb
FxnqnC3gXRwp9ymnx4lf7JICbd0IXeLi5uab9rLGOKBMaZM6zK1afdNgKln9TbAC6UxLXxn718Cz
K5enbbxLbCqLw+pGvOUCM+Vsi9CWBL5+xSSiABWgDlvnewcEp5Dlul86mrv00YIyoU/dQdn9zFH0
7DAno+TB9AXhs7Ba05YsCaX0az7/VzJ5xGY1ROabdFMS7zsmlj7z/BOL3u+hGs4/lB5R6UyfKc3m
9bcU0zhqf6PsPAd+Jx0GT7FVCDZOooMNIr5wtOP8z3fb4ORuiOY6CAGZOoP856L2G6kfCL6YZzZL
hSoWE9T6d0+tGHM6tQ44ooJdSiEr+N43kNuLKWd8HbZBg6gM+njG78qrujG8UoHFMZlaVTJGAC54
XuU+79Xs7daiccUSIGj8iFHdckeYw3keztW97GcI+g0jnYB2SlbQ+jwUohY2fWY7IWj59QSBJ3Vu
ZjHyXxARIDfY/QDn74aU1ru/9zHYI04Ona7tR8rpS45MLAw4KRdn7iJx+anefRy78DQzEY+Gytev
h5SSVYdiYwqqWAq2s8ypRX/eNmTiR/u3FPDQBLN9Amb4Ja2QnQIgBC47mYRf1MwHBMl/64Ss012u
7LeAz+V70eSTqcI0TdDJ0MeRrrFEw3AMcnfH668SM56Lb0dTAJfME5ZvewI2EU8N2dFu/sj9OW1h
cqLZLWUQHki/85GRGO/cE4vSBlk+SkiuylpyRZze9V5MU3wFQ/PT2/6FZ26d8FdxBXEumcKaBGRj
hm1dj83DBKd/t/Zy/Zqc+ihILr3cXt5MZJdA+wmZz9efykzzK7i9cDc0YPl1lPJNU9n75b2n2a85
Y16lyc1UIkjkJ+6k4iCKYd7/AA3C5bz0pHgqgOXFmNb8OkNe3z47AeFALTtggzy4goBBLcohZyTw
g9f9RVjBjqJQNCDgCQlMPhIGOqeUSALS7HP6nr/02t93qph92qh1X+db4bLD3NFfO8eo5BCvEGS9
P134XX26DomORqjvI4BKjkx4/dXrB1r1xvYpi4cEy0duP95pzZnhd+HcPz8lZSDypeUoNZJT7rqb
C/5ImTB9YHy8zPvyEFiHzzmjoIzpCLE/0p71Cd2ZhhLzo/vUPyWnGEgVwd7wLhdAs7EebzHYsl/M
MT1y54dXN+m776H3nNIQLsnyWYx6flv3YRyeC/E9GHsJgBDBv0Dc3yVVHRZVrBXQZc36KukdlDdl
W8FSFcz9q+GssX1nuK952eQU/qYBmr/VroctACICa2ljnMDMBu8vEDLW4o+2B9GpuSQugDoevWuG
C6l0tI9a9dEs55gSr0fOqU2CrA77gJZfJ5Mz2Fv9VnzZeRjMGYBppa96lbsftRBtZ5R1gLA3QeRm
/9l+tBbwG60/sUrmmsao9SW1sZCFzvoFeGi2WQmqMW1Iwq7tyvaATx5KIBsURTvT8PLGIUjQXpg7
jpAHwHSXigha6lkq40SYVUNm7I4ki7rakS4IuKQSKbZZKiodDju1yVQsceICb7naczaLfJJVNBLF
fPiD8CqgHcDZTc94420isLj/XShOBVj5eZsLf3MFFxPs4605dIerp8FLBqV/UNx6Rwfo9oX3KGR6
jVXUHSbl40le6fOFVkx/UlK2tNJ0dAsmhcOFW4NpJ/2oxvh2oF90ozv16I44cp0X/C4LioZNGBPm
38Dz/3mrRQqS0b8JMFpPW1fnpE2LOKF4Bg6e64C/IkjsQyHej5EW8sMHcvC/WOoQz6IVfWpN4C2T
BvXYML8dTfQgxAmImDEF2kKlJ17uxnalXKKhsuAtd84islzaPEtq4coBkwGXjapTEGwuHnlk4N2U
TLmCmnd0O0nISQPvivE64rGWm79O6SdKyB0RwLTAIlE4yQp1EY6InqMJshsEEIO55G+UHL/YR/xp
LWopQJ6yWUlg0CVdG2nbLE9AkGmHwe3e1IiBAqcuROBB1KC0qjCTuAEJTxr446lZWDJZCWT1BYeO
Lcz9MuWheI38l4D0wYICi5TmCk4vIWKPXLmWr/yk0/LlcXysV5ItkVHXORr5MUPalqvrFhBPHXu2
LQ+OVxeSIsIekTa7RaMdireTafJzyaeXsU83lHO70WiPBZs0gt8eQ5kBtIrMg5nYtGPt6QzTZxYI
9Bdu14Q1QppQ2mB83QtWM2KDVj6Xqnkpv8DBMKZXbOignIPKyX+FMAIXKnexRY61255JJVJzcnnO
wB3DQs9NxCnFEEYz74DVjqxzSEIFR2Nj6MwNV5RHssh4hWWtI9JwumnNgvm1ead20u6FYwoygMGx
sRTnD90osT5CWJLlQj2rq5B4A2U6484PpWkiyEDdPRQuS761gcN0HmMJwJTf63TjEJ9TFwUUq0jM
VXV7uPy0kAD93zEUxKcTJyzTRq092I0m9rGvbZQdA95SrPehzvNMo83yWDfOtrPKd+bhlppQvjKY
EjqyUg9ukxh+WVt5VaLaJpwU0/OQzL+ZWeeUthzSnnl9kN10zF0FMdDYj/bohJp15ayC6sluuJJR
gWtFxH5t1DMdrn9BQo0jgp99B3y6WbTVauxl2LHy455v75cwugddjRt90aug408s8dtxuJj4s/66
Ey0by89+ruLGtduw5hM/ceZhQylBOXqkuaFitt2ql2PVKQ4/pw7NRes06ddy2IW3hYzIyV2Iu6H5
sikyloreVLltgTRQ+Z822Bak75qs3RR1EkJWbqoAS2CMg2wzCil0yTY+RdY/8FHhzF2Qhbato9PD
P3a/yH430+gDG/tGY5mes9lUlkCKFnPsxxTNk30C21/lj9jiRqNwtzqOfts/n58ZaTuAyGGCgd2j
LsyOxB0pu09T/CnGt4zA0x5YbDLvPXK6bTiba6aLIFRwYzDOnqWkaLXLEbkaKv+rdZ/3j3JoPXXP
kc7Ugg0xd865lWNtBdr5uAKfmvfbyKUSyclPFWEv3CHpCi51bR1/cuGUlv80kc8/nOXmeT39m5cd
i1juDVA4JPyaKlD10J8cFvhLLxLB18R4knwwEXn4B7ugnCKmH2uozqYZb8eexnulqD6XN9qnWK4x
r8RhrkMo1AZlE2q19pyKVXTzlAvonHC7awt0lNdRzzWi9Tk1M9TOpqQj8ZIBSt+wLgMV1qCADZNq
puXpt3g+rEdiYPWQmtX2DstDUSRrMUliDg/0JICF/Id7/TNOaMeUsJUlaCULQbWspVj4vLHic+Uo
RayLwpoArxYu6903joPLmg28VEXNEuP5cAlLHoX8lYOuiOucM+AmMPI2RQzbjvrHi12Diuti6wRX
/Xny3rJyJSvl7XODCWNhK595rC9LlT4Nr9jRnDGMoCGrDF5zcIz2toop/zlPOykk0mcZxoVekVIY
+5zrNnnB5sxXF/EW9zNj/zqH7mVhRRUUzNw673oZ9KofGslCtDcTT7ffb8IGjGVtpiH2jBs37RfO
HozAo9G8UKPuWhbS/m17qNIoCi4LqKns8Pex8dmwvkBxg90TlJaxZU8GP762YfdvWjd4VdGoJPkK
MdfdKZQRoedYlgtZ1Ql5GRlB91ApurFGAn1C0pjRlMt6SfXZE/BjhhwIMziamQtxknB1c8t3ogap
rL5f/9hh+zqN1PcgIWmbJ2+mM/RD60LhWUSMVl6krhIw8HPZhQO2ew8jezjMmuFi1ynJpdDWlhn3
FRSxdWrtI9IwyV+4ha44Da1FaoNPLHKc2/0zaJAxtpRXmFKOmMyi5ysDdvgfMnU10iIfXyN6PVIx
w0SBpGsTtoEd82fj6VfgJCnC+lR+W9VDaO2ij2o3lE3xiYhZ7X9lJ3nzpuGKOQ2zTjL6knHm/Dit
cJ0T6TibGx0jlwBFME18oQxaNBe0lSzhx3Y7w8HFjs01+MNaFMI7K9Aql61dj+qZzfb5et8I/L8v
xIN/xk2MPjTaQucYJ8XrwfON8mKXnO/PH7mN/zH/M7G+XBmj2SvFRx9CuiEuTeAkRZhyYcFRDXcN
lGjJ2WFsm2DI03dK1KKjtf6U9/JDnca6oi/PSSjZ7ITLkpF/N/MPFSrABLbrQRr4dpvy1LqL8Qbt
IJIC4ypuUAPuLB66MvU2caSa5Gg29Fml/oRh+Sbpwj+q1FLyh+w5I1XzX7peSJLraWNM00Wdt5XH
DnhMFjGt7ZCdyFbmo4QYCW6R0R27MavQgxTLxk1lH/uxrNXthKOesn1TBjb7cvNmyxyi8iq0XYqk
uiufkhz5GmqSFNz/xdPDj1d7NtZFV+1+DfKKtEy9llvXv6el0W2kT0hyHOSPiYuWipExjPfWKa0N
5Z5CoNIQWCq24j9/yEXMsNacZypxe3MGTWacmt/BfM/hWnrLFg7tNy+BAoWlDrhtXOEpZAsW8Uih
AM3+JIQJFfEW+zNjkO2yQ/SY5g4WdsN59h3rOE+VOfmumlrFG8ao9Gmoox1pXawnSko8nfFuVoNs
eujjW9LCG3kZiP6yKoecwSNMjQBKNNfwi2r/xdLjm6GT0xkchJiN5HaphvsdtU1DMJBKHjNlSdtK
GGBEEze2hCUmXkeEk3zE2z0t88OqjYwSykz6fDqtstobKTmqGMYu/VcT50UVTBylG0msVnKekj1U
BfX9wWy0I/ez2AcIrRRQWF7EGDa3wZHqBGjI5mQJM2uKgsB1lLXQHhWSUdOO73HrfBFsQsmgOAQv
celmJcDr75eHFftJdAIbzVw1PPcRihH+NEFvW46VvJ+PZ9Rb8rGJSS8kKN+G1D7PZVyNRDcBk1Yi
Px/QeQglrNd8cX/roHxTo/khu/TJT0LO/9HrqYmb61fVCHpOaGgqaQA8OXT0ZDA2BjXegc6FoMSI
0aY5I6pkpTjHSpgexVdcjllGsXPSTD2QF6lsFx3lGatnz3WQJHnUykrxSgEN2Hmh8EaDYj8LQHiR
DqrtxcOLulGTgoNSGA5GXk8IP2j1OUIRYn3IfXWj7P/fvJ1jZiZzT1PBQ0yNvtfjd7CPeik3noRJ
sB4TbEl5EO5XGe3EV1G3lm+OQaMHpWmnabT0VYz/Ks8PHHImD3hg3y9oktah1LgfZTdVCxi7jPJz
k0Y+TNgx7RJiA1silcfnvrFomxy6mZJ4C6bDHBNWBeTFwaDszEsL94x46P3NRMtKfEa9VrLoxHoI
Va1jhMNd40UZvXI9MmAiy87GURgZTcw09o0s99O8U44Nj8WECN/IXldvy2ZkWpFV1sns8/rHi/nD
KHFkAJ0Q+1XMW7+wOUP65DuvBFlLMri9nFOOdN4hDSu3JZZ1CAloPD5swVoy57WgP1W6aWr+Uxdz
FG4H9tCqRRry2oxjK1/dQrf0/Btmn2uCOsAuLAmXGBJei3BsqpSj4gPB6R6V0nMeGR+hKhdW+JZx
V2wtB3QYA+y05vVm/xQFrl4pLrb3ItVk/3BAmCSed5/EpBC6uWLaA3/BgRXfclz/bb9c17ra3G+N
WyZG22E6VVk3QfPlB+I3LJYW13KZdgJ9sGW2uPV60icR/Q95mKsq+IhKG3JM36ZM9FCdkQ8Gc2mz
k4+QpV7Foy2EQECaakZmNz5gcZY/Fm8M5faMNBZ92lAtahW79X40ZKbO4ZA3BBV9DE0uX2eJrniY
mc/a5MdplGtQUG1kSsPdJUTnd9JRKs+iUGk1nY8vfIo9ODH0jGMiDRksm4kuh8XEn6bc6xYfnBm4
7slw/Vn2m3WdOpLQWUfMXzdreDCp8f6Xs9FWVVUYRnrgVyR0SD4sCTAxg8sq5VEVLDGLMhZz+CQB
8QhryWvf39+roi6iF8LS8C1cXRVC0VgWfZUTl3gpn7Cp+vGyklzYVu74tX+9grgFn7vke8PlhRRr
o04NBsJRti/af1iI95uW3l6S1rtndUtlOxC9J2gB0qK1qeP1dGgaFkB6E4lZ4CTCGfePZo5Qq8KI
1UYsOeA/9/lYxbHFScuQmdysRHe2f9FF0lBKYi7JyTB4SRv2Xm7Cy24oIGSMSbJGFXIDdM1IodAQ
SA4I4dmOveQ25L/88QW0Jv0wZ1ni5iLLmiFljM5fq3h7wPWChEXqxlrvzvsw7Q1eLJJ/YWvW+9Hm
umbtJrv6pK3HZZ3g+bWEGfiIEL6tnNLJvwlpfHOQPojA6S5+CSEyx53BnV6v45fnljWPA19/NikG
7YVSFYUS0OE/CND5vWrnOwNejYYARM4kItK4yH7LoS3eQOGwx6CDDIsBbMkLY+/QVGUiBUXsxrk/
zvU+i48DExxPLie4kDzqzzQQNZV9Z8IPj2psqaewGlP9sWqSIiXNJj8pgJbza116DWstS0gg5+TY
F6u9Z+injkpX6LYLHrWCB7jKRuH6oDw4C3lcfwEIXDy3ySENrQG7TuhLg02jBPY0nAA4Qk+jBeYZ
h5/jcLpJRWUML3VLlkTnYMqkmXtDIbRQ9Ki19G412E2THsV8YZsq5jCNNlyY2QJ0aj88hFUbJkr6
Q1vhiqL9JPOWMEVwLAAfmeRjlI7tJ5HEQ1/u8v4CaR8PbDTcq7449zXqfGphL2mqLsKbHDsL60Vy
+wbNuTjugHzkhS2BQwloHqPQk86xnDL8LS80bPCK3CaOR8H5NIJpGi4fFd1kZpSpAc4UGVBz9xLO
4aQX3acl02cN4rL9y+764QXdCQLc/gKy6Pn3hkYHcmte/uZYV2eVDKUm7UgUavRn0jo06QfEEXIC
Obw+BL663GQgWt4HQla61/A4ubFiRBghgKkCrBEQjKai0rLObFNw+mZEQohEVAtOALxJc3O19IH/
FFYqJ5MG59Kdm2NQ9i09XaJJi6nHz5NkF6b/IdQ6cM+vxGGNaNV2cUhq/mmZRGUj1TfiKb2S4sWg
j10LjEn3Q+sR8zKBvB9d9JdtJbf4GAQToost/j3HNSIqHZ0fHRP30iMPG1kNpi+2c7M0hHyFNN7a
tNaMg7QpDzommoIaeCWZazDwwbqODurgWWUtLnhb9Da3G/PpK9bJs5GcVJ3+a5HjLM6DwJ9eJjLA
O7J52HhxS1f9saCBb9S6Wj5hIJ1ZicjgnvIzYAUJcO2UwdA/dSiyhhuaFQuVdanYGn1ULljTqlCZ
23DsdoseihewsfOLVXNXtA3GDz6wALe+ycX/v8Mu+L7t3Aj0OZA5OzHHCCa/pPMP5zw5/6SlvR9E
9GnVrAJyaUVphEzh/UvKbOuphw3kUWMiqcfnzTLV+Rlt1IUrPtStJ2NcCKyp1bpd8WJ+JpOaCB5Y
PCKh2VljZBXFbCxg6HpBoffRe+TbW+iAC89z6irxzx/MjsxuOqbT8+JBxYZY963G3WmY0wklaMMg
iwcDGvIrOWGOQKBzFk+ynAyGjScmtnktNAbfIg9EqVPcp03ZLlm9N5AgL7udqF8V9q47Vw5u2Nhv
UzsrSIsycdGRbf+6ExwVUXjHUXyEDdcQit51RwY8T1K2cAyzDISaSzOx9eyfvHRc5IWyId9qpLnS
zJlzFlKvtzZQ9dy2FtX+OSdVHjlhUoZti9BGA09fz5Sjr6DnlzdGY78NKVWki6D1lJBMUPEIPFQc
mneDpjxMPmUlVzqsbv5FPxlB8H1G5Ou/pMa5D9wklImIdOkAG2dGeUTjXzGxmdKgAxLaZR/xI1Ss
9F2jbMPy+DSK1YZwIb91hqnA/qTpV5Nn6YM/qaoGV8iwbMbEtH24zN23y8LPT/tjzkk7q49iteKD
qZ7Gh6S+Bpmgx6FkbkKbbZyq9hn66ikpU5CvORAIWMBYAudetR8ZB2YiCYdkBBA093AQAoO9vpe2
VBDPefS5U7CHskeS62pyjA2RaI0vLh583cDupE7Z7054bg2iKDsWpeTpSRTkf4QqjEW7MBQUEOZX
aMpTlPRGDsX7YJx5TkqIUVlig+gsjw+c7bTbVa5gm0NeawB30m47HFVk3NPI7ZrF3yIaZuVPXDC0
lld7c9EBCjWhO5mFk8UMFLtqkHFdKxNVY7hSAc7jQcmm7ME9vXtpeqHQ9fXXdq8LpUjEEnWETa5+
+hCSNZST9NXThKb6pdgdcgXdLdxhHTPyyqnB79RlA6vLiS3aI3B5GH3jD7+ae+aNO9MsP633sNtg
MSI9vLaA2mFCZJ8dln0P80dQ8wYzxdeyXNn67SdtXjjEW4NzttUiKxOWX3EmF2y/h4dg2DV137Ik
ayggxNZcOqPORdWzyUhPTl1W7dbWYsloIfD+og8WrN2Is+/8r5yolUWXfFDrmh8S0aycvNPCk9da
DRDmQ4z4CNDJnvOgBUNCen6yzpplubO+HUXobrcsxEFN8if/75M9dXXPPJ/Hmpm6VrkMjHWj75P3
Fhq7bKI2nC138dnMm4T5EMtDU9frkYT14MSxclpBeBOrnKAyoQHhpPfJ4++z7H+tawV6TAruU2pr
DqBdD2N/EsrczKDjUuY9JxPc9/j+lfwYEN4UFmkX3DFCXqA8d4p/Ia5C8PjnKZHxG2tC7oFjKPCd
qOn8abHjzFigUeqiGrnnwF0+xTktwmgmmM2geBjFziZDNeaul75ivZTiqFudT6rLDdYZlhaHJx+v
6i2gCP2q8qHsX9TOokvFfqYTmjHv3lmo0vYnMh7hcMzYoBceEs1rellhfAw/ixIaIVPgZo+kba4w
L2KHZAFyXHpqKmfximzF1yOA+O4zS+PY97WdF5vnt30CuXnwi/7lkN6U/zH7FZu1PpX/aFasTrQ4
ktypErmK/VRfIHkRc9rZw8OI7KY39d3qXHinRMUOkki+/D92TCPDFo3ArDoDULycos4C/Vc1twbG
yT8RFPHwvkJgv3L4gZ8DDNDKx3xIaBAY67S8Eg0Hg/423tJxpR4He5SJIn0QhLCRJFRFJxRpcCmv
HvIGtJbwXx5mk4eS5l5ufNKmmLk6WNB8euGXdrjCvXoYw+OWdb3xpsD4JPPYmAzo/sAncO3FKy16
lfop87JlGmtNqNXsSE39SZ5LmWaB1jr0edjdGhEq67b5InWwi+uTybkeNEFsEn/ixMBMXNjw9nQZ
CIGOrQcXepBpZ+JQ0+MzZnl2ZLxzn1zZm5YFq2Kq3KN3FKPgmfuapYJ4fMWiETjevS8XymrOMEMI
aA+zpVDdCAfbINdg1iSSt7RlgO1otRicP96Rt8/7dgOuXePJe384VIf5keRLg9OWkOW3IpYr19EX
cl7RMIq/2nXEWfmp6CK5NkgOJdQy/DLQe/6YQC48tQo9biwN/3essaV4/tAp0qa5ZCOFsPI1Yygt
2wHXI19biUlcD+h0uiog4hOo4vGcTj3sEV2kllM9SZzKvFwDdlq8w92SSmGIgbOMhrD4hvLivXUD
5RBWUPqho0nFc/WilcjonRCosp/eq2j3+BYsrkDf4t5Hm/t4MaE8ubuTs17GvY1oIaCVMzcsSCAO
u5bx+M10Ph9EfAkuHndLbIZxv43esopsRvxrAspm9HnPbU58cnmBR0GRQo/GvBbX+kMz8zUsuFi3
fCl+MCzwz+BwxFt/4UFYVFsTaCC9fGEIWFAAf5O/5N8sUlpohv3XyM9d6qj6SNvx3boabccTtDJG
/gJ2s9vJxaOWXX5pudmepVX8XhLRMXuwH0RpM2KZSpsoM8SUIXG8izXk1n3B54m10+0xsIOGFbtG
sRzMv2W/okMcavziheVu4zmKgxaAWuRLgyxDVsTM+eG7CwbLQygtYaIHL6gBm+n8ElqT0ENGKhQX
R7QFIhFwXqL4do++lVr4XWCMDPS3UvE2a/zp2z371jvC+KIMWcXb0RyuXWKweIbqFjasw6GQ5E4R
dBJC4yuD8BLLgseajNrZ5yOAv56zdCrDMlSGpRLBg7jP68+h6JO/JvrRzK1uMvdrt2PO8heArEvv
A4Hm6MRqbfpCuS2c6PSt53zsG4s78c9pnIY8sbIezJEIZs8JqYfmKnyeaPOZ3ZxAQLO9flHsFOEt
sjJSzIsEdalkcVSmZkuKceD+H7q/nObAfTWaGK5G6jbQmwICqfbiEPRfiJ18Sz9428sHENdW/UfK
ZlrWCJipWjJDuzEaqw0QEH48jFrCn4XcxZNLytDazJnNxHo6K9dXS1HeZRKbX3C+Yi375S6dIzMD
ftEwz40ZDv+9c9scdZWZzTAtk7XF4laHJbksyb84nIZZY7CBvtPHEtnpDl1Lk2g8c3s5gVbskxuC
TB3YH+W3Qj4uyNuW1sliPmHN/nIhBMb2XWSIjzkVHkoYULYliX0YIfmEm+FBSQmflp5CczDbjqGW
XJGnU54rh3OwdJ2+LcY8KNhFl+zNuWX9YhFwmfaf3889p4Ova8+YI+FA/np/C0V36bSYkDDuo89O
GkCmJyayaoZgsu+lICZlAeVVFt4SN+7NUX0v+ssei68YGq8xEhsJcQ7+mHkpTcPEtIKmIByVdNQX
kB22Er5inCyr20FVQwHVKtt0V/Sv65FSaO/6Dmc5JZ0dL5ZlG3TpiF25pVzYrp7JrMr91MtQ3Okb
Hgc3lMA5Nru4BgqZBqFT3GkHhA/qVj4nXKyxnLA3k13lMFQMjchuvXrQGxIx9ja0y/Te879fEF01
8F5FjsMp9KfYoET7OI13KLvmFpYP8qLGeS22C/kw/7whpL0oJoxrGhfb348I1tmFblMcTldut+86
Dz6AYJmwfolLOWmeeHrxEmMkBxOxA3SixlGgH8+UHjSU+38oSKc8EyIBvll+pDz2vJLR8nI2YjVG
5rw+oiLXE/E66WtIVIHcsw2Pbffd6QWQR+E+e+pWonoJS5sQuYuOu4AVHoq7LPb6lELHLOLog6nE
J29xfC33fiQKm+zVuWAv5a4zmukdFB23diG6xA9AKi3nMIW4Ssh2hV7ZFn2k9gIfseCG0P70anrD
XYZxobZ2OzQIGn+e+wOZNaN6AL6VR98bsKC6Cngymz4fS1Oz6LW8+iwNklufYOzVCv5IBEiaE3BM
gfSWSSRk80izT7JDZDHtTqxx13AMSXJb7oSGYGS0lsQXjdgFOS+mJtpWBdN9zmZHKq1Jg7Oy7NJT
GUhWykEWQCMp4Oo3XMRPX0BmeYqLpcsMW0OMe+MjTLz4LpBH2yG1dCTu/X+42a1r2bceuDc9M/Ep
TefjIFD3nAvmq6M/pEjr+ZXtnsvpqf3tc7i0VfSUKKScGKUbIrfBrITHZN7cZsj1hz1AAEvpVU/+
PqKJLhPdYFdoQDXylXGe7xYNei4xy5iwdZeMCz8n0WHi4Hqub29bcwmxvvB1i6JbEGmKQgnMxvHN
FKrEYlm7YvHYpF9+pqx8z8tuFVe5zkYfT6kLZLKYxxoDzD85ckjFMsDJi9rwAs7Nl55fVRjZhyiX
4K8MXmGZsdClgFBFTWV4xREgfebvEcPQdkv3LDt+1OkYmZqnVvZDL3VHCD5A43YDhPjgyl9ThPYQ
D8eNoCIk0N1n7TVud3fG21FADaQSdTXmFYVj6qmkkN6J5GjXTp3D732D83CEbi1AVdgZhRpSisk0
7Eri3hfk5hR3Yn8utq3Oe7bdoslY+zNxMvANku5WxghCMbL/uiew4AZwM/u/MI5ZQYcjx7+Ve02k
bXxqHH25pzcH+3G0UbwCnRldxt+xF7c6qZ3lkH5RFrc3Vv2PyJNUDxITMjjqZB3n7GvJGcJEL7Z1
hOZC7ZoYBrkDkpL4thvaMqH4VRPIPswArWCZR29awggvvMeW4m29PoTrngB0/XDl2jZCiYaHuTJd
r8DCNIlyCXsClNQWZv9RiPfKn+6s84jVQ63x3o3AfDEySAKnPlq+IdOKnTO92pmltQ9jjnHGA6QG
vjYxk/lhH29VA6GUiZnVds3P1PiLWO9m4UKrUDNa8quz2bGrlEbguHpXH10MXYMg8pY9W9m4ZblP
ei0pvgM/7hPPfH6cDahS3fQLOeWavKfM0cGT5dbFWf1qv0+BUrE2JjSBk0uqyBUizTPCg8z25WQF
r4oZ3fKrn8DX16NRAPegsPIKVUlY9+oXw7nFU3/FaI8jj6gmEOJwtqln+rX4Bl22q3hdLt1bpvO5
CCMxiwYFbhJVMIk0mn5WtFvFI5Z4ZYyJfAXf2cxfpdxsZfp6o0xRxS9wQkQuylk5vh9B8hsxkewX
GB45jkBHR6szw+GU7MMGa1D+aOn/HYLyAq8bPdO48DkhuO2t6EUK9wuvMV4k7BcYq5CEbaV2hTg0
bx7lgerd+wD17Xdg+22JzVlCFJ9IKVb/B2hlz+WlytywoWa1P2ZRBXGu7N3BalQ1JXqovdxzLR2u
aAWWt8D+zFeCyWO/zfTnSqnpEsk6vlHuAsseA1j03ax7kjt5xsA89uzd/qK3o9+K1K8IDLP5P+vF
SKcDa9ye3Q7QE8OGaz5k99JOXJxCMMJukOs0PEmx+onDGKHua/mSTp4f+faoVPjXNY3dv9nBMlfd
ZuH3jyZffImE0L/IEhBkH2c6PFjq/OD1ofkRy4P9SPJDJy8knfMLhpCMvlj5q/pv5I7/3jnmlv00
weXrVUbPg+z4UV3mPI55ya5lmR6HvfutdEWJe9hs0uX2XQgZpne4GGe+j7RXKS/oLVCW2T44pumU
qTOtUFu7KO7c+rQvDFaUtDpezSvkO8eoswYBBIUqpLA/IWiLj7f1HeR8Ms6fUnke/sELmwn+oG8Z
L2vLHR2RHboreadbLha6WGRI5fAc0EYH4f2mo92U7UoGRAHLqd1sY0lmYMmC/fR4F8DJZ6yj1ZLS
NIiRD5uQBX/EAGjJrEi34P1gXCTeHIo2c41TIehtdNTO+jObFE83dJdmoaZvsvgUiOqBwNLSn+bh
nHUUrW0e/RCB4u3fL55cp70Lt6s0SLbqKpLd8HZDFRqAUWI7uFB76FLKECRtf0muTPKNoa4qsy0Q
jE86vKnzy6tESx6s8zynnkVcnuOoaouh95weJOeF7qMpcEZiVgw6daQpbM4HBCxpYmI1NaHF4T4Y
6Umo9RM5CLHUDHKzXkJK2XP+jnAytO9y8an3sud0i3z3XVlK9JPteVOOflZnHw2VLt4B/oWtJlvF
S5LP9cO6wQDCPUWkrwPBtu5CQaP4LtnE6qOT3zFX9/+Rk80MPPKkMagGvbDbPnMoKXnJssPKXBbE
NMClhR2xyX921B2f1TEI2o+Wyw0hComih6XjeonnUltCYLWrhqMNXC4WBijNcUfYKhv2BlaR+OmD
UFFtOimsgC6KWV5TK9DrOEGvgL7w0bN1gtVOonbiW0lUDJvz+HUpMcyN4zyai/ENqpHnqbScuYJF
oU3zMCVVcaN9IAW06mmaCPz4pm3xKnQNZrik77xdK2HTWW582OUQhjTBFW1YcPPiV8dzseTgEEtA
D7gIKOjBjvplZDByRcShmwzdsSNudrAm3P1asCAtLIPJPCxoownR4YFXGfvc5nnvSJ5bCu/iSWsm
AEziWJTMBldcCt44+beIZ0y6t0+iL160+v+UfMGn6/tw555qkG2w106yZccqBKEwOBYAVTOGCJ/I
MQJXRP3jF51f9/OyI9wpJWErGhH/iQbSMvCUKE/IrAUmDK0KQPj+3jCjArlVMh/EI7mqwWJmGIwb
fIQfg3NnfF6T8RMlfjx44dHAyHxu8Pgz97sng4R/xERKudHYKq+ZX9ACwoCQqfHylK3Si6G3F0X/
4fNktRLpv+ck6mYsW1AcN6JAL7yJC+DUb8DpbgFzkK8EbCsCFHFfbto0XGPrWc0+7E7jRzqTHUxN
tlm9xo4uc785e5pYWu/7CLjl8sG4qc0Lfhnr45X4y6uAKFwZ6P1XtJCRUCcHsYXJVizhOx/g5ZSb
KfHcMsd+3vvn0d0dntLbRcFNaE08QlELVgCAiA8hhjW2aUML5eRpc3JOlHQy8eBWSRQOZMe/SYPY
XS/SQuCWsMkOK7OCUcFoWOggG+NXqLnIorVMo9UY5qwfF7xumiRGD23aVKKamIeW9WJqhM5qk1Q+
QlEaQ8hlf2FYhOzn8+Ox5Ds6RB9R9fmB8EUpOEa0lntP/VTMadR9RvfDhQinOfwJeEXo1jx16ROr
FYmDaVB2ze+R/kiaontGOhK96qs0dS86G0pILwuOuVXg/TZ520hXlvuduZueF86iJyJiOBVaBh7z
qMUKZUqIEs2X+rm0+vzFuOq55sWez1Alef5V774bdf//ktTu4S6c4dVA/f2Lzx9/BilEg9XKwcyY
zcCyBmlKgfBt8JYmCDwgCn5edvOqSVA930GO541KZNHrelv7PnrSibBmAv0J3aK34hNzx3DdsTiv
+x/31F1czDeRd98eLleU74JdGjjiJZ0C5rHnWQkMdjnGAIIR+m65XGIWIYTXlSNcGxYz1M/uHiFp
4Zxgmi37fWXJwZHEmS13khTGixLjWk3ksuycCpA2kR2wHRlrrvc9T/GQY/6SsEit0pm/y/b0SPMX
Iln1aIW6tZyTnYlxXCNwiL+NvZXDryVaoZj+TXS5Nbv12ciFkGILbRHXJ1LNpJK+BunTa6J6Cdr0
VR0hbMOV3Ambpa9p07dmkZaPZPoosVV7ixn0Y2FylFPX/bh1hLkVL55YqkeW08LSp1mHsQueGrz+
oqWieIyq5Seveey9TBtYajCabdyr3mCQLNJCFAWYdLkeoFv6Vq+d2VkSoaS8kbeim6v0+HToSrUa
w8wDpQk8DO/EBWN65Xd9tuAB8KrDZgfsGWVCEENSFZJdyAJQKJwi8IHRV7vj8RE1J6g0PIBvz0iV
tBWoIVLKPcqVK87WC3ULgYgIDKNqmkWL+aDbDktXV9UXuIUHtaObmO51w+r3irkAYXYow/nCEEh4
otiBgR2ZhRyc5Titf0AvVPsC8EGsvgI9u/iiAv1KhETKYHibFFh5zUPQVnW+Bu9cGNnXlcDGPxQ6
5YugXWuKi/sj7k6FD3urM5692a4L9feCG2NtBujDluOkggt9MDeQIDGigJu/YZ3smGYMn2UwZP87
Pcq0O7Bf1sxZN6iLnEam3cykB0a/tirIshBI6PclYD2h+trzcNKVjLoKmbN4inkD+0+pmwZwyDVF
pfe69nJ5zW4oaurJHljpJDUF8s9agnmDYNbRqo42C/pv9DXjgZMX8pJKdFcPdQ1rqqwu/mA+2onO
aOghGrsjmY4zk/cfWxgDGTVBkRMYTSoUCenvOsNiZcqXhpSfHW9nxwlf38r41NRsWkC2WqhIxf3E
hMtw79k3FmTD2znwDUT0j8VhhyAai0ORsSIw+Hbs5j04VGZqdf+PJkXcQNb/QDnGEDp3t2rXcCZ8
JEZJ2kaPkePwSJ0UYvxDQu609xtqwWCddo1yOgeD8q5YjOoKKrq1KKPAo7G80Tzp5mkVK1uK/Y02
q+9nMnXtf2HKxgWp6sWsWLmeEf/m4obOsnXHVyafhkSVSbQviO/yJA2aq+ji6qXOtYfH2T2+IVot
97yMLN97JMGaOp1qDdFg3dYeMkY+uwwZfnZnniFRKIHdiuTeD/3bL6MdoJ3WOIynsJPTOm1K0nDH
hJR2vFfBjj0YZsvD4DKtSOSw/7Q1QQ/1NTGkx20ZTCnvJxuABN/DHUtakyRNb8If/9w7oyNdGsR8
9MIX21n9tlr7HMGOMjsUvMaFFPmmq3ASTQipKjzylfL1Flz/DfD1yOBIWo4Yb0LMvKZFf0i/65VA
0SyBh8mTAcj8V1GzXwuNYhIN9dULocjPFrXA3FPIES3G77WDT5g9lvnEuMMMYOZ49+3en/RlBhxE
1Hsx0sjwmW56TYkgTTCsFwiYiD6Di0NgHcKvDpIbyaoJeygv84YLQ4NkfHvGUX0P7N0rOP7kFDdv
kAXImMTAvxyR9w1DUOIPfDez1Nt/BnQHVrb9ZIg47OAQ+4slnEez+w+NxM79nROLoFl1mw+UfUqQ
SYYkVn/1faYDqAtTdanvi3+f/XkAJhRsvSxT7UvVtxAssdEvj0fgcI3kIf+UT6K9/m6Kl5sD/dLZ
gPKcrt6xmu3r/Kgw0ooKasAeGPG9QLdYdxQZJ8+7jIqdypgQBkw4k3dD6e1NOiB9COlagbq6GSjj
mkmJE0ue1sz7U1SStQQq+1t6tIQ4MngEJu0UHvG9UIIbmgJjvoUxEfjWa//3WtjwUwohYD9bIk3s
RnBNykWU7BhQVkVW5DCAbddFFmoFa+dk5W3tUknCV+VTNeYQm2LTIXi/tjqYPT2TVLQZP4xU7/eG
4gkgsQQvsAlIwDlqQ4qwwZzP6lfgGWU2qaGZBx3WQ/emAu3B4EUGvSyJ+GIydzzMMtxtIvPK6lDt
wEEA9vDiKrjxwXlqCjGJZuDVCaMp5CLkRWH37q+QjCdGRJgNEk+cfdIxa2sQTho7DZBna1nmYnRz
d9eo6lmZly9+ixGbyXDOS0aU096bfsOTxYUcC/SD56+86X7S2K6qT/HWk9GhVY71RLJXsWLM6nix
KImdeu8O8ogDdMTWCwq9Kf9ZIAg5JuAmlidT254CADA5wFqsuSNqgCw5+Am8D86h7qZpIA2NXqv+
iywawZdd4BYIm6t/AgtWLBeqMzp1RRvOWO2Yeh4qaqOazypfqqxa9V0WJhfVP8c5YTYbm43/fSHd
fnEprJMjjEXdEW9Ao6CFAPfvjOu/8oTe5BJP2twgD6hEJXCIRa48krwpDCXpHlx1iWcqDl4V5rSe
4VZmNkR2Wf1OiDoYp4dA9wXOmsu3TC425ic0J+gpP50MpMvJZPCzCSIqmILNPRbV2N4rRD6uTRTO
7f9xJ/o3twPr+ut2Jy88cPkTU+3tRk96OdtiiONeahetVD3ISn1tvgY87h1BajyqTNk2cxDqsI05
/sRNfKG2EGx5K/ZZ/UXfaRcnzkjHxVbbX1i6frtq/2CoPHQgqVjWayIYBD4CGWI5l71s76Dnvo/z
WEjggLrPbG+Pe8yK3I83N9tJbIBH1ti1rwMVuCXMON+3xvM7s3QAUSbih09vzF4wxzHo/3sFeqr7
z1zSCw3TkutYPeiDh/kF39RjeoSG9P9K51AGpRwTs4kpPWfgEalGiA8bwGYnbIaJHikv6x4I18y3
xUxuW+8+kuYwpfqxwk6yAhipjmiUDkVa/0g6431FB4fNwN5TzDA6SiRfDnPo9LXKTqSgraAhMOy5
pVji5hrE00JXX3q2lKuA2JmXBxEJk5oBCuSiWN5PGnXzGIssaE5lwXoBADdMnNFoHeKL7bZUbGjJ
06FFd3TYycDejkCwPTKc3+fmTmIuQd2QCGhYQ+pvIWKqgcmlj9uBlbO709uHNmtqj03//u6OS3nY
Is4KfYRvPoToR7I7pTFxEreZS8/jK7StcuELt/axnP0UuCC/KtJ6nw/XPwscyi0Z+FiXZMwj87A0
xiYF5RKA8akfFzpjcXm5u9f3sm21HToOkbsrJkywQpkQv1LlufNUohc5zYhskK88zXIf8TpRH307
dvbi/kNcaWInwJpyMDdF9UC86ROIUvK+mwN3/+YjNaZ6ZAaBp/yDzK7vyT6xriFcMJMXhfVsMVeW
6cn8toYBRxMh0c/Kght5Wr1vTrWhLluZetuvCyiksfxRzbe16JGj35pyndJBWIXsWnD7892HCZ0M
QX2V24mHzgDvnSEZFyJ79j8b0LebIb3qhWVuk9smTU8Odu/ycPhuBOcqFktKkIOrqvw4BdaKvmOt
lKOUQAsxvnvPMOjHKfh3NE1sDVeVnd+rTokAq7RXHVXX7JdruH6unj+tjEBTRmoLvNdBMVE2tplH
1PIoGeBklFhBAkZrpgp2d7/zHALCeliGO0r7FvKec4jJ3uwDn+PtXt/UBMfL5EXw7cKCVMo1b+29
8gFCC7u/5zPp0POlg3CZoLW1Gz64LvrZ8RgztCQ0aUzcHpTwqWYg74KCKhT/XS9Dis/hCKuKTJOE
3Y8OI3QFwjA+MPJivFkRNgNdKyi5qEfLqmlL8hmyQojYkKbNZ9fBwPidouKDr7/3acAOAWGbAFgq
NBHPKSXPORZsu2pksYPw4dNnhmHVmpPFK2Qefih6nGYi9e++WgGrQPWCav4L0SqN6NdQx+BDrpI1
6UykKHZqu+HuDOKaUWMke4QejVLCT+rs469Le48cx7M5XFUP9DFxLziJWhJr43KAaWIEBqH+IYJd
qRd5JvJQHk6RxzIAXGN66qG8A1VrIUbfI57YjRotA7rbQIJvFDhqhvUP2kksSYABAgKDumYCTCWI
r1U8UVX+POhHHOPruftXGeJddXqySPnC6ItYzu4rMZqt6+0prdmrn9Q4/sXvfaRPCKXptTPM3oof
e5RQAcH9MAqJVQYtEUt7UPtPWNTpEzGt9n5O2yNU1gFI4T+m6L9c1idYTRTq2kHfXizyBZ/Y6xDQ
qazqgFm5t6Ha6wvW4U9b6YxlJW7IBFg9/W7MErR4NHhYw1OXk01wQdvEhUqkSsPsThovAbQ3ae4Z
UNr/NQBBOjRAJvsZzmBrR2dotF8vZAhhRbQIBz822uihViNy8qL2LgMGwTyOXJ9stFRKXOI5e/h8
LUgm0n2atthi7aHikSRSQnhCaJ2GfLxoV0x2z0hOcbwlJxhL/AIdb/nds/jxqtjSNpb+fqbXvj2Y
m8phAZEcJg6akWKJ5Dq3E1J6qBMg/As1Rw8KOG/12/JTkejhKdA8RIT3eyAvHkGa44y67zItipsw
NwSQNazOYQuF6K8zqQq58b7+ihsNbw7UAHYuQ5asCGmpvTBSKV7ATUC8xzuHB1Be4XVrz/DkhWqY
i3ecjPe6FwmnjX2jma5xUZFdgX2aIsDgfeGra5Cm8t4LMtr+FtOne65iZbI6LrqtHX1vymxPoNGF
h6/lo8Rsn/DxtBzs0ob/b1OzTqLhcOum5ZRndYpypTiVBNUum1bLoOO9hBUrOMm5zzmjRFUAt9rG
qzTODOh4n/LNnczlEXLT6zZj6FgcHuP0sjNAy+urBcER+ZMbbjBip8C6qlhDZERDA/YFy51fmwu1
v30eVvAb3O6Je8H4BkbXaKPKyzrqDunwUaF4IPE1XdWiWp+rJojSDX4qBWLFFOpcumqKq1J6TdeQ
uzqVywxEvaZbgUT54wdT7eWfjDyJ0CX7JJlzREmFmcxNDlgmXkvl8UPlXPb2vBZ33NvK1l717H4H
iPHtTz2AGii8+Kxx4DcQKF1wYoAU/TjsGUf+tOlhkFoKKC4fp4tKzWdgE0qnzjisPJ1g2FjTHXs6
iEt1GBQfKcrk1VOH0ZlNCPIIzk2EGXqmkzzQzIZwkFPI2c043k1/kNQTAjxAAjN9EyHIW5PYdob6
F8cX8+qDPv560VWQtdZJSo9fRY/s15Bvq1lka0RoahAdRKYJhxprTtFeJEQQTlJDp0N/FiAyfW2t
UfgxsUcN0WCw659xSj0virvAPi/LvfiVgXroXM6LAo9tmI5JZt4JSscDXHRsn07T49mu43z/iDHJ
GQGdewR0hlL6xPERJfQTt2yEJluPkyZePh+uCDsApOdd4BuhukfYiNEOUMK0qDPOazCxIdu8s0nF
aJbFAwfB8zWiBYG5k1NySoiMpepq5txyIldeZP/cUKcLaoEgkz71QTovSwfspoKaUry3JNbb6tz2
9LsyppUZDjoRNUnFEQ+KUhCq7NST42BxRlxz1BtzKUXYz5hQneTPdQIok1bh4c3SwRwE3qAica43
RU0I2lpwGtvMs41x/RuzDmOKB7/r/0OarIxy6GNTeT6mfxs3zop50T78ow+xOWd/NMT08y7AuZrQ
wqSkRC8ac03j6UksEe3ZTG22yVRusk0b/ykyxli4Reu6qs139EMXyL2Z22KYDMIR8wQVTKBkZ59q
2vct3GjPs9+Gm+WPFOUSM2Mzv7V8XcomqzW6nX6HwxYdOVdadcmO5/ssbFI3PgYYrI50sddx5SHv
CMva6z5IgVwnUpfDu903ovHRqiSy0pbh1UC7wJis9BybzqrNKQEo8VPogt0T6r78HUAcPwkaFasc
BAA5+gPATHqCwDha6apuq4q/5YRcFIy1EWgq0WkWq+7BY97bWx5lt4BWobL8kj4wWKA7+pRayeUn
o5Ex93RD7AeK4emoHH5UrhTT/r+bCkvGOAhXyL/CnM53IM9+OfXu9CjzywvNeXEP9PIDay5tqLpT
uFsNpLB8pxz2PNsyHI/RoaWFsjO3etEP2xh54CFSCxo04tb2XhRPqlO64iLxDGVob+1pwuyuyfnM
2MmLgCiP/bkLwDG56mtmq69F5mwcPbs8Q0mCWDkA8zjby022zS6iLhgFVQB3NhHJOV/1RnIwisVo
vOf7XLFHrdXwD0B4Mb1/ff73ey7XmT3ObY27e2+tIXr6sO5dkJwvKpEIV4xs9FluH5laQ+BB/cvC
hbTVLTJcS8DGTsauGzQU5OFxJpE4rtyhT2waVV0YIndJ1xbJEsV/wIS0/qJXAiXJ+JqEaYnL5EvV
XXf6uWBfQoAcUYVVbdeJcDt3/sWWPbI6iKnyWnqdXNgAjFLA8uFJzs+LdIuZWMa4alwCgdf4ZkB7
ucBy7mYiKPx16KHWqvMD+2nihXNkII+90EOerbkCYZyTna0IUB4GAYxt0IrsWnZTfceffjd0PMFM
y6iukQXc0e84Su29wbJFbyDdZOOmRrZqsLua8BXw1GrJry0wrziLzAf2LCp+6MG6Ccg22vTkMel5
RvHtpwTJLiuLutPMxkhqHwRjgdYjuETvFYq7mKZyrONVsxnB6W5QRBfIKlKIg0ER5NUWpxAwtRu9
Go62BNfhFIkgw1AObRUapEJIf6ZwbWJFhKXAHNjA1B28301YMEV+DV19LKHOpNZ94UAmrWy5Uev+
l/hHR9kq9b0xivzUJZj7d9GYOt6yTXpLxNpU4UjFcJ/1WwJ5HhAP8mmIZgQ5V5LSFfPFxTSeyGmk
D81PAfxMYCnxrC+ONqmiwwdjl9xq9y/0VgRoHAlB1h0+cBaofFR3rN3ol75iHPsQXZLHoTPUzT4V
3R3u+t/RxGXDfAzPqdB35qvmr0/RMamjGsYwzoh+0l/9hWL4pKjpW/RRupisLDpnVV4SuU0HvB0M
CcUL/JzdiqyieE1UJct+6U1T6wW1z+W58jOBfL4Hkunzm6hzfwhJKILtXEGmXLJm5nMTwlPAQcdn
lEv7ddzAofv2Z/Wbjhxw8INJ6pT7ctnPdX+MD+bzWp2JmOHvwmDgzQYV7i5UwmITToIueimS0HAC
TVpJYZ45KssmSEtc+geKuTD6ulZ/YP4RDaOYg1S2UlBmXCeQfpliHXGYIK8FUNTTNg1DucAwpSxf
6NvPcvdPFJZbnWf/QH/X+ymZycTFQibBf/p26pzx+EPZKgK1aXlzSSp6WQ7vrfq2GiX/C1KQrNtx
nXUtDw2k0Bdvr39Avr+B6qGy4PoOJ4QuMmNAIWpSKwDe7EibPRLSyI4+2amotRwh+MvFWinjridC
xopkJGTpmASx1U50HMM1DTARvRkfseDamFHIKeHZXIixPG54qF7c6zlRV1SCo6FQ5iC4bYRANpa9
/glswqsmCiteXHvEJV2DS+HcH0gsQn5jU8NjEZLti/x+djK0un5q+v4oljIXAfOD3szptamfzNma
h+08dnp1emwZtOoodt5E4VRj18niLEXaW45fayaTOuDRmFU3gnZq+W3BORikSieGwVKCpL3gCUgp
jTaIFoHFXQ8w0/zRDKwfg2mm5/GFl9GkK/yFYbihSsjXfbgOh9SvAheGCqdMkjGww3LLHA9vo6Ft
uwlroZqkUBbOPxCuU22oTeqh3fjENK4HqmRiFXrWZUIEY6x3xeihd4F9+VUkvDjaDbaWPxCwOUII
LjduID/l1qndom/Ky1R7B17tvnExpDZOXBfR0u9ph4+6OYIUZQXnXvDOqD37/D0nVuAl59NbrSvf
I5zFxxZfhwtcd3CIjHoJkYYx9FUjdHByq0OiD/jb13xa4iDewv/F5+vcDMs68X59hukeFuG6pYRZ
wpU+A83VpQsABb1t3xLDypMPCqrkbMCgxNy1yint8H19fqCrcfQdgDKs4zgI2jKJBnX3LmYbVscZ
PL+AKVqhfV5BAncbbX4+TxbDVQ9j5YyNDn/DO9gDipj7izH5eCdE7tLprnL+iy+CirqAxHC14RJ4
kJa0gx7tfRRj1hMx+tbyYS6FI2kEL8UEKHtXjn7MhrVTMvONLY/xpM9m52+OVjdII/ZU1KgCXovy
zvOV8Lq6nZsv4msbU2TIwNCJzUjKDurbmRNJK5fnPyEpJzK0VrpkYFwBYFl1JbAWYaxVngEIxT7c
LYMFyeuNHxHkFisJ6prkh1E4thFkoCjr4vD2GuvAFkWosMkFoiJRT0pPqbKAkJF4DQpFCQ3BxIAd
+H1R8z5PFrIUL8tPv7GUJ/Le7NaaH24VDTvUV6lb11RDD+k+uLlEYtN80/UM5UC9xG/0wmYLEmBw
q+YyrdcJdfeT/YlGDtZhUEUrjL+hZoh4bXsHOSAnN2rWoqFZhFvtqLBw+aXvDW1+jk8zad0Vjtz6
RoaI7FEko2a89WFXS+1hiiEKFon2xpBJnb6YRtWQt2nRusGTRl73Khbx5xwCD6NbIxZuRTcJ2FEs
iAzBj1TqFmvQ/p7DwNAvHt24X0Z0kow82ta9rB9VEdsx2dp7zZkXUTd5MxtBlSh3CkjE2op5XV+F
veEPpUB1HkZ5b/s58sWQ72xgmUbvK9vbx8L82bgMVrWRngwYrnN6Fa13zQz1oge+nPl6rTRXfPfo
LOX96fylW1aLCD+VyRcZHGbFYa5MRwVncUo9e71GsUTWfIp0zgQFdSnPKvENGLpnsYB/i8tievH+
+48SGzvhpAwWBVEaf8o4gagcOL5w5PLbXPeFuyHQ77is6MCaUk7/0nMkvcDz0kVqRjjz86sfU2hB
orN56dYFMZMLM7zuLvFSp6ukWJY3RWesRGgVxUkVVAgTFQgCFr5lVIcxsbTfc5YI3eZLb8CJVPtZ
oOCbuB8bleLkiZMnbP/ZfUSAhFX2eIIvQJuSQP12afF697ObWJX/ohIeKpW44Rr2DMWMMxyPKtT8
oCAdKIgZd6e6KSG6eva1SzQX0N2CxWR4UXyYSf4NBBPJhGwVKSVwZxELPVlOWRHa5cxuzNgqfx0K
SB9bpBlpmUMxecr67ocv787Bo1UMEmwxYT6oL7GQQCPbI73h7DIOeaKGa7jdg4XUcEzp2+yuiBFe
6Q7EEP332rVddwAoUG+7tP2CM2MBYQ6tDdSJTpzDMes8K0DDGBMnFmRrwKvktw2SwB0rxgtXxGhg
KoI1H3mG2/egHXADG/WWDW7D/6FPbiNGn1SiBJ/SoPOlW3mOLw2xHaE+A0wtvDqa07rXzNB3bGHk
30C8gkJNdA9S9NYs7CrnLmpBtjzyuAv4q1pVi3b7x5MOx1vw1CWsV0nWd9q5Rzt/rRgIIdnHRNZp
NqeKBITxL3Z++8qpD0IrIxyzw1ANuG7JkZuzP740okHKR9oN+Bz9/YS+AhDpCBdtD/vOTFGOL96q
u6Z7Md9wE5ii5bzVJdX8V7HzuvQ0BDSNDMdqenkFrpL9eedRXQaOnAj/lNvl7AQmjSZT/vJAPLAr
jhRNPxaQjJ0qI0t4wvQnrxOJ8upiYS80ZNtVpNIK1TNMTQy7GF9jDCkT/R9mP6Giuqz2CQC7zHk0
F4bBGicq9nBslPPxs+r8BvSKu0rzmO5FP8/GMly+JSuzhtTjnL4yykYbSlPlkk/2t0i71CRpZyQl
AklRGLNBykXlz2K2dnFbcNRI9C08Wa9YC34YalA4qEiPBL4haS4YT1zyeCm6fdto7m4cBdJvoOHk
wSRuWceUI7Bj13QZDb6yF9/TIdB7mEQm+ReJkjjFKUuzyocGyAAdj4eJnvi7P660TEY3a7U4AQG6
FMgRfM3gRHM9UYG76a5pEmRZT7koF4nIe08cneTwIWpVAWTCVR8bl5XzprkThI/7r6jr8MB76ONA
reMKVE6w5BmFltebEAlX3ChCVqeBn72trM41nSrqI8zgz97JbX0We5de/R7vE/gGXc907vruXuGp
iOmMhKBPqb59G3eI8qAZdltXdnwjvJyCGFDItaU6t3f0gHXpNiyEx23F+Jf5n3VIwYZOMgGn9DZ8
0j+xR4iHc4MSXhQW+nHgyiL7k0HxNcmDed6uTZ9fJ+TMKR8H+RAcEr22CTvF2nMM3Zo3rhguQjNg
MpIfElGSTGzYDsBYtwbP5NRpRGTVk12eLARCj8Ve5p2BhE8un6oJxD1F60OQtZEz8PqcgE1pBPqP
pGErxInQhmUHuCclpaqOFaS+zKvSE9zQGN4qaCQO3ZCFEik2wnMoZ4mLNDTcMpb7Z6NDsfi6+wCI
+MUvq4zcuET+KssOeGl3o95bu2JZEfsBLZ1Ft/WnGQm4hkCq5i0bUSOKDDxK/6EAsYG7zqeH7pYT
PuxHkZZc1VRLMf9R5LpaXcumozfRTu5HpkQR8YYbhe9uQvQZb/USHS86wrqiwGimh0OOm8gvqMOj
cXUkcbp0yZn1zu5hkhTjYg2FUTa0nVgxt10IuVXzfotN9HjeKdSL/mzvzK32J738TD/QdQ8oCc9H
goIVL1yrbeb0dnDdgBzXSPm4dDXi/+yh+d7KAToUi0bdpvB4CDbdeJMoHgVcCNV3A9dSYrv/tpN1
TsDQSTTrGl/dVCd0mhAcDoMcQCXL5t8YVYkvH9pnYaLHdOe8orp6ZVkix+DKdYSuMiB+saP3X67u
WTvqevTXQylvKdKIn6blRCA7cXIGMheWjcfwJ6ocPku9ylYdyBrr8AU9Fd27uNyIsKsaDvI0ICH1
fpsfztqhbDkhZHDjdiLqRO/A7J3EuWdzwXoUgAlAMi6StMc9DvFrKbvVFsW0ilFNAJOxwHhIhAKd
Ot/FjPHj5Mw8pYteG7n39F2aflzm8cpx2g1lIPzKt+armBCd9+Zd2sIG4PHnBkhixJuNTMD+xDRT
/TdFf93+eo28rqqz6v5FHe8KVpklBL1FzxNYpmOg2qe4pBRWPyaxkEyhVzpuhQaUrfNRj64MRnI7
+c1YuqrjqHvJuWPtcCK1yuZxgfVhhejUJZcm5Vd22KOitNm7mCw3YpZdEMqjlNsD6+PKSpylvnX0
tpPBBlGvZe9yQXCRP4qaNe1BGSu12eTEZtO4OagivKFXqj5hwP4+vBATUglnpPIXlsPlv8mJsO3J
dOcHoo1Ykq8MG0AVWmCz9y+uBqpNcgal1lXT2wMG6Az9ulr8kDexbKxkCpH7/tXZO2xRE+qL0b7O
A+6uR1PuEQwhZiu0jQkBjHjtodpBUCnRPpm7CHwpuwgQHdw/ap73jeSS62zmMSSbS2ZoVD2FPycr
BJ4QfpcyYJDYlahATvHz971nzVtxv6miuzl/j3V5sa5JoJNH46G+Zms1b0Z7RvpBZO7aw9wyraCg
YxVLwCQVjvXRspcIJ/EhgtF1VFyqLleXD+YKIkQ92BfTVJR81hL6WUrjegDfVDm0Nsz6OSF1aAoI
k+zlCOC+UeGAGq2l+VpKwgwm7xLqd655+Ww1qv9IhatSO7qKd2Nbvo8DsHKLq5m+TcSxrzJ437ZO
uasl+Cd7KQGB/UdjwtV5D8/XDquowIWDOIH9lgYbPFOriuyqX1xjFd8HW2ke8PNmjYjtBCwQAd4O
ssFO2fLmR3cc0Q8f/EAKo2pelIF+B4VResb/GQgUah743uv1U0oSMQxQk/4yHC83tRbBLo4XkjIE
rSLpPzlXZ2OpuMDp/vePzhHL5KbHYMaC2cj1NchL4ctYVlBlZPfJ85Aui8w8XqrNbNJ7lgfYh4Cp
T9ZnewoNft0mJOOOuFLNvCBd5eoUI3JMqPQFxgiIRpQ70atQBbNrHHYn3TkCdhTlhnUJlIrGY6Nb
r46CAdjzFAd8iq1R4IEDC9sRqzS07aHNgoW5Kl5IKAKSpopgp9wMHN4BMR0AuVwTbkq24NC78tva
iLTxt5PQHELqbRsDU5rclVTVVWGyb3mbxiMbmq4b1NFWHfmyT1TdJGDtCW/1xuBDP/i2i4A8fB3t
c/kgrMiDOiGM+51kYkDeUkJzPPeWR04124yw2aQSAhKcwt1ioqsS6cS+W8BNhB+JGYlKTwij4QOW
naxZYfHrYTcNIpxWEFoBtojmr0SmWV0EwtbmlvzRi1P7lZrZp0YD3EJuVHwp7TxfipztQI/ezxAG
vKXLtiKq1EPjdFVipdFazqJBl1RzDTSc3hl2jnsrNnq1ZeAfStoxdivcWTZdS0Z+2FjDo0BgtcPI
b8yYJHtgvGmHXuPGdY3RE2xFXxPbC/ow2x7yRYCGFFU5F+cRU9VwXMGK+nUhksnbjZsw/f1IoAkF
09RHb0j2MNncsfzKYxrpLoHWaZPoOlU96/J1fFFRk1PdkfhIyr1n9eNTWP8N3utkc6PsF2TFCjHo
1pwk3m1WnS8FJwCNylZydopmqbsINJucpI+G/EEzcHjRpLfqbj/g3eJKbCqJgCUv9mnLEErnVgTd
Rl410I7yyJINTctg6oXeyYdgtrsAbF3pq/RWCkD7+20WnFUzwqE4FQYEwHQj/eXwoMZY3+U1ioF/
dGtNyn/E5KrYndv99yMTc5rADnt+vYf9aOjYUCufITeLr6zsOdNyu8G43oLcECQ+OoOkC9lgAxDv
/f5PTds1bs/nGmrDpS8XLGIL8wEAdk1k4fCt1JuRZeBI2CjX0HwgkUIjZPxIb/vJAy/A4BQBh3UQ
We3UbXvL3d88OzbHqh/Jdxl6ewNV1rSna8F9+Zk84L8JmxfbNMUWRG/5vRJcb0ZyRFn6has4oOo7
5GnhxnRz9IvdRTik0DCIgNrrUIQe4FWfhPRsuORfhvSytI0/xP6nhF4hbAGCHaiqlGmC8+OT1Zef
DKcfHk1epoTWQRNF6CEwFwS3CVlNCoLtgyGXEJmcV7z9bTwjyZ1vMz7uOrniUqLZm3xET6IgCGtG
abvba0alh9gYjpXc35UzwjcKQPSc4hm4bU1kvfCZlDoQvrN7jz8bKbyVg2P3dD1H5NGrnoHkoEcq
4Gvydiq4eKiAGqw2WdaCGSdJYb79hWu6xb81aml/Di/c28DI7j1D1htbhqw9qo7/8L3CtSu8HErk
Ne2tcUwWdRPvAb4vpdVcyRuUPDNHEajAl3GYRxARXyupuQMnI6ckiSyJnCqR+HhjMh4AdM1QpZO4
JKgGLNxtY/eh0s05o0Kz7w0Kg6Td3xhXIi7I2KvTLGrGhcSFIcfWK1VGaU7oSParDB/+c/IgATWQ
MOIKZKB0EIGL/4sqlFaS99q1X/2ytvUpfcgMXgCCDVNMbsApfIQ9QVRvueIoVAUqbI78nqio40R0
DmOdgMdWhPsSJ6GE2/oLVdHlWpimjLFMjWABuTY5AePMkDj9KZhwPXFb74SJ31SFeOxiuZYjYWS6
vEsj0RxPNa3O3rF3ajjb73Yl6FVBhTNgdtYyG9gS78e0MNmxmbzabvUfVT6Xb9kxqSoi9HgmLY03
XyHAB9nyn0/NEF34xcKfdxvv0d/hEtDY0ovW+LwShL8CV550JhkESTrhEFutoWR3DXmv742AKAFG
htR1zWxwlRvCKW9bRbIwKzdfqX2yfl+FO34G+ASefliBZoD/sop/HECzaH0mn3oO85F6j03bv582
uKvT6gVMrsK5NIU0RxekIv58yMugQaTSR6zmWk49S8Y1g1mxMNYnwmZx3PDGcSf4U+ho3iOLb7T+
HHB89xY/bHtz5GGBoVqMXoAJN3R69DcN/BGlI4l3XkTVfl9YQbOmfUanfJiV52Yich2qC7Ky+Q0A
zkh2U5GaiVsaM3Im/N51uA0xKfpkEYLEfa8FXz7XWYWf3Rlt7T8slBIj0GcyWARVccTgVKYbFJxC
v1XZLQvKSV25xfL6HTLhM+bR7UquHmUe8EFbpQub/QZYXPzu6ovnJ7LcK5PzNZ3fHsoJXXaDpYS5
AlpDALIKa9Z9UXEmXpNlMJ8bmbb6D+PfcPXiYDrNnRdiPG08X/vxy88mSz8mTWU7Uy+aew4RauJ+
/k3CO04OxXsx4aUy3Ugt733O64f3S85usxQNNT7y1dF5SXj3YgWGHlKPUdNUHq5St8IoAieQhjyw
bLjhBcCG/9mmGdDWBEl66gAl+ywsJtTLoEGTd6L9gtN8dWhV58g4kNq0EPINpHzaW8gJ8/BLhSTP
tWAeIeQ+9Djx1oZfrtPrrMh+1gq5YRtgJFlk7GYyUekG5LW8ZuHFd63gzC/6+yV6bSqCUqzA4Tgn
XVn2d7tQ7Hn6/qei6lGNixdvlIMDLH5FMODMel541x5Hw6iaJQKEiU35J5uBTE8gHykM4i9/XLKd
aA150PFb7Ng7jBfECPAWhFYYmhC66D23/g4xkEeeFt5jGVpd1qqb3WLFoyEOazPKTMtbsNCKiKqm
BQ791SJnctgvatHvg1+P0ngLvSuZqZtkTYdyDsNotrbONYO807LHy5Pj/gOMJGGwAS5ImMplFduL
wQIEYtnZ9ENG6pjsLShpduueu+ymNHVz433FnOWYSHBgsyw5fyNrN3kMH5fw/6e1xUSLCC+NAZgJ
+KpP5xl/rdWdJj5jT819Q1ytuQryO09j5sTQErTgvpK9u1ntkQB7Zy18nXBI3fzVx8o6Pcbgfcvz
RBo3gUMaTPVpOkVsNrJufvT6GujEIifb1Sc3w8ME9BbficA1sLzosBnTRVh9c2nHivKoPwS5usGr
XmtpS7/nZ7mdHAMHhV+b+NsVFMCSBBt/zua5P9xq4fISpBymUNe36LhJn44xCwYofgbmKHA2XF8D
3IABceUHe5fO+65pB/DWD7tauFh+UEbkhJ1mM/+pXB5w0Rw6/sKd6lj41ZiUdfKr/e5LH1vfY9MV
DfGTp8jfO6906CJJynrCrfBf0O0bF9cC0yDkARnCGRUjU82cK2cj/iMFANrI/n5/MKQ/vxCF4n8i
IjW6higGtX2W3wY47RIFJfyu1uSnZS9yqIVlLQ8RaSA88+K6X/ZphOTjR6aD1SVX+7fBPDWe6tWr
NChE04yc/diViQrA1diE7qRhTNZ2L+7cvXa/I15DqzVpE00WFSRsKimNRcKPP4//XqUppxvDIoVX
v7xN/2VTUr1SgXYjg55/IiYVd6Bt4LFqXumXVqYYoyjSiNrvRAa3HxbTAb0w5EFfBOdut1Q7aPIr
/F5IMlQRcTjHWUqYJqlaJJJQZy/4TkzrPVjJAnDCPMsotFieDyCAtYnK4yPLELOAHyyNZo0fx2Q+
HVUI4F9+DPsrTW91lpDRPURT2sGUqh7fPUr/L9bqBDcfCgUJULzEbuJGzfnly0Bk/HWb9FM7iYeg
0FYd5YRqL+Vsc5klU42n2OAUVOiF/od6Ketv9UYwhSkqtOH6s2Ki5E6DOnq736Uh9HtFa2+8bJLx
maWr8+r63xLW2zXsfp/0gFhZCD7a40iBCYbd3A6/74o1LKOJdhwX5x2C8AYgWQBrWuiMTValSiqn
I0PYachlL5S2m90F8pR+YxkHLw/ZHabeX8glRj6vvS6lUoGEObg0gSIcV+7Kl2e17pXS4Rv+dg3U
3VfQIkjAl/itByKSEtqqE0M7NZWbjJbqCC4dShlmU1w76V82cS8oV5j+Yqrxrazjh7X1qVUDwxiP
W9teHZMXPbTxf4c690UI6fp1C4dT+JDeTvhhB61LyV4iPTcQG4h/KKkMrukBSi/08EzJvEGYfy23
01106BfwyOCNwNHVQ1bJ/WikD1eujf6TOC81zFTajEvRcmvo8BnktGx0fXsp52eKO7IEuf9nKpTY
jmHfdzKEsooxrOczBRDBvO/BwQ0iltdlBOKpNojpbrhulXpoY5S6Lp/u43pgOByO0B4x6FABAnRt
ySUFVXUReFSFjwoQ4iGE+s27tGermP/X7emaxzU21RWu3g7n2a/6+4BKdIWr8tszHMhKmvTJqfEM
5vEFcUEY6F8y+i0J5hHjoiwPF4elyin+7geL35Thv58ajxcI+TkzL6QqX0YNIU6KuVGyhQSGIk7g
Wc42kZ01slbaKFo5/mhTzSG4TUwQdEcSQFydmAyp7O20NBuF6pPM4myDYLkAzazqKykP+a/eU2Cg
dF/bC7VPz2oDkzwFClZ8NLc6G+mVr5F/yYvPiewE04JwAEYmAcBCHSvaJ7ej2qvcLybpeqrj0lNB
tjempCTuSWD40akS1DQRBRAotfK+fEp06bT/2MZ7S2CbvHSV4IzW5brklL3YghM4Eq7iLwFd/8Np
/V/8oZNrt6n0tgwXBhNXqCNqeW52CIn5E/FiiOsYrUvlXqlJzfOAQz4rzbCjhhdcXRwR2qydkuOZ
5c3fV0nnUWCx85NdjnHB1vk3L1tnlBzdZV69kTaAoSakbbqTSeS180AV9t8uYxiY7hKGCAi0DXsI
HsYte9ARv6fKbHSm1kNNxNJmmQ8bcJbFMk8w7+5lXYUaavfjO2eJH5HAM4v6bf7QbJz6aB5hVdp8
bLeCW95ZQ77jgzwz/QdjixPcp4Fz5z7yTTFPg6TQvsfZfbA37l0xTc9Vd9e+o6Xe/xbX5PYmt4aV
U+NSj24XLg2f3tLZX07xWYohR/L94+hMshjDjwl7+t0Buchzehju+YAeaPFbCWb6GUkY6CUjLPux
nuwFJCrlPLvTgu8gvWhQwPfsN6CVk32eRqoljzOX8GzWloxHMA39v8Jv4PoDCdBkogsOs0KLKdpX
vXzsYPcXnIrIu24b4mPYAylNFRArejI4Ux4/zrs6JxKEZsPTxaBbHs+EKUsXjuyq4MdOy3tcwdVA
QOomc3bK4AlgVCcE7LukSVYXrPI1BepwivAosz7nfobzP/38/sVIUV18SI4Pnf/LIiPGdL5ZzlOf
fyutbgE70N/33bq4TwlKBHt9AWU9ESmEhPBeG+yaro1UpgwIQK/qnBuNSCCM3TOV0OLT9R/Tq+uP
O9oUMfPu85M1laCb+1ALROqLOvi4ONA0v3HGWMBSv6jnUMIM7tn98L0pcD1hCcsRoWN/IVulOLZn
qGu3Q2cQprXwOBmRqQ9HKfBfokPc1E8lZR9uFrk3jVmffTRVP5vITlAh6YP4sRiMGb0YUjQ/iyFU
5iZxXnKMMq2tp0TmyxEh8eg0CHZZYdMFp9fKnvWZ/is3KdLxKebiYCT2L9Ppjrph+R1d/NXZ6lkx
0+MMUxPXf8I63NHqqCH+6401w+KLX4SKqp0u9TeZDBtb1i2i7voWsUoUgAo46/irPCnPOaGfQocV
xoMalGHRAu0Qc6GxUnHKDQGirP7DigGHUZCmy/o/2fsw+4nbmV8xD2Zxsf3BpmnrW31zu+G68lqp
zCeSNwS8fo/jZEeVZcebsrj0NQUTBC5JoJFzXKpRtRZywKofB/VKpdZ6m01eUBL+JI9kdnustYJx
mH1uDzD2bD1NYEY3svTkLmLtWY+oA8oSSqI2xxWsKhXZtoZnCinnvZHKeUuLeKw3Vipsl3FoxwRa
fijeMREjn0kcoemyzncbN1tUMusfAT4AIXm3IIkrNUxKWHSStWwXcYnKjceM2lhMI6Frp38mgdUo
MFNLH5qBnz7gT9JPqLLDRClQZWtFYG2UNy16ZpyKP0Y5xsmbqKXuskMoYiM6aQ9kOTAgIvZ97STa
70txodLofuI/pR/PMRZNkjiTJslOtHzorImpAmWMgdB0tErgzT0kDqJkB00OYe7+uO0RMgg3Wo9o
p0qZWWQzGjIsIqhD+3ZQRQGYPS5VNWdXiqOiDD+rzFJ/09V/FZ9sgOtnoqPYNYtGlWk7zjNbib+E
TRwRAUvAuZy+06TMIcZqTYLzEfFsmIY9V/gqWLTCUXftq5pso+6i5jMq3P8i7/pX6SllCJ5pDO8d
D6U0oNNZ0H0Ag7PvvJxmpPVBNP11Ekq9U0oHJcCd0uei954v9FcBU+Q0CafTXQSxaNS2onn3IjUz
qmeYrBHZI3SAXrjZOFVr4DbFk2XGsKzfGhHvVs7E1iSmQ/kw0r07cEHT5ufORfil/wAfp+RkXSeN
k6Yo6xmUW5PXaxcJmxnfD+pyUkNGfC9fSHDiAGuIoqzCzpQ1TaogTb3XHql42EKeXgFtS9lgbRoc
nUG9ilttjNbC3rDTc4LE6Mtdaf+UE99LfGBHxqJk8KeAjQPrgbzq+nSyG/uj7arA7rDvisqd1oEW
yA2u9u6Odsoyx0YBNdFE5fP0Km7gf1AeZkxbKN78VnF3aJYmvHrZjWEgcgyoTW5cRsDz0M0nW63j
6m0ofUB70x+jEUVqFC/dO/baVJqFeSxRCfCt4nYnSUaP4+Rq5FtTsPet69fPj0v/djd1zgEPQ/C+
i8pl8yVdOcL+QeittWJEdSqUcCcwnSgGzGQnTSonm1FmNrMip8KmzVG+z7PZlmzxbIfKGon3ZAQd
Ua+cv9y2DDZ2H29Ocnjh/TkZIy1nWQHgRvb2E8PnXkBg5IA1a3bQ4CfY4w7D16cQfzxlrqAKHMo5
ZOuIMVCx2fuJRvBZUD1kdlYNr5F9qTkkMl9uEED4NS23TASMY/9TiNFcC01Skh3JWY6w9IzBCzhU
kiSmfWtckjyHNMxOrnBcvVcQ7lNNn/fS7Zau68KgbVFggIuaXQyB5H9oaK7euGqZBv1C4KOwNhfk
pHgfT04fWYUzfxN9R2CIYcs/nn6kpSqhfT/QnCoAl8GH5qJ65wBOlnjnDukVNEcHTeTfdieSCOxp
39WPHzBBbZYTU3sJF5wv+Hnkx2TxkAvZLJXTU31VOpkd3X8iCeo0g5NbCfqFArSCZH3jKAt9JZKb
OYrXcDwGpMujzZRQnH5u9QKRWw0HXZAjjzzGsNIJ3Jis2IdTuLykPUXkihffgNy8fIWhWrnoyTh7
BSfvDJ1y64aa7MT64tMktBi8szSZ6RLi49eN55vQqu38bItA2FiI/XX66h9U7AGPKHMFw0DUYVL6
2yxhiqCST/QvOnBVG+ZdUnbSLzSKsqqftpRID7N5bqW1yHBLxIiGx0N5L3yO3bePtKeiAS/O5OQ2
3Eokoqw9lNVlwtfHxftGmtRDi8GUPXk5myZPHqxn3rjXS5ivTMai7y8aT0HoZzs0HKWjgr6qMvBQ
TxTdkaR7ipry2lMu7fn0X54jFAiBKl09ufUNuezV3DzDdHYq8OdwPxMKZh9xdJUIIcIycsxbgmzy
KA8RJdCsSwc3TyuKDUyD1CcbxgjeWJasUD3u8xkPmm5og6XzvLooVzVFajAcZKILjkdEoXJoGQsn
ZvR2Lo96oqbR45rfejpprTJTuWdT6iEp+tDN1b5/L+UmCf/Xwx3gqVdV+wSmJS1hSBBlVfbncANn
jmKfPqUE5+o+lTqFk3ZHjiSDb9KIlTph4V0Ly0ttFJbQzEcPhzM0eNtQVMJ2HJyJpfZMHtBGFMRS
oy/ZW9tebC0sP5G9657JWFnZRSYphm+gIY9LF3cQ5BFH5SQ7y9pJGAPd0HgK3rcZe11SN7QXPYXz
trxzi0ghKCBvHGVmYjSyliujHH+vkak/Ha2FLabUd18x210eio5b+UbdvqpRZvOgBn0388BORVzh
Qcjk4jNikAwb0+elNPT6OnvKJFzbejTVwvcFuKgwmUuOFddxNWG9lINMBbFzxvuULYw+Yj+nT50l
os7+hK3MGaTb+h58AT+dIwiaJz5rjIvi/CZFSlZjtePYsEv1H1kwapXfrzepH4s40t0+z/Dxb9H2
D+M6/qRCSjL7nG0VLWYOAmNaCocVbWqFCv0m6dc3AiZD4KXLMKT4bbGi6YpAO1vpimS2Bf+QDHiK
twFKpjjuzwA7RWvNWpXImjWaAYmA2jrS6TJ006hl4gRAdrvq4UTHlpOqi8wxgSkEiCNZM76tphZe
bOvmzZtka9StUmVwq+ohxvP7Er2s5OSYBxSMe/rQzP1rzI52QB5jiWIu3YWb+RsUkHktiqYOiODg
atS6uY+IPZw77B4OmlywJnFEIaj8JWJYEFHMtqfDKs3lfSw3Du5C6mCDYKPeCm4y/wGCA9TJe5dK
FzsXuy9/hQiP7czzdxlA9k4Qbqz6m5KIR5ZuLVzoVTDdQCuXO4KZf+V8VdVC2OIrSXq50EQGmjpQ
M7D8aVSy/JVtqzLgunsaI64jg/jZNidSCZ0MChtS4zbHXetXEJ78yEay6NacWIFHdVwdXuIrRz+3
gVJpCGSXDnD3q+bYtPeNnsyex3NtBNzQ/z0qgQHF8d+GkFp0oStiamwU+79J0rLjLvMRnaw95pqq
ma5YE0ie+mcFRtlxU+dcOQRqToptgUWa/xSgUnqGOaU0skRj8TpTNSHP0Dzk4ysqoHVD2OZvEbnG
cnm9m8Q+QvAm+XlnpO4XZuhOPOCmK2bzUKZNqSQ8aZfLuiCoI+RGz7MdzTTAwgx9/fDe/4MAevLR
Hpb/IwfH3apKjZkXs1u1TifU0A5iQYd5jnBRIlZMFpp+PXH8hQhyFcvpi8qQr4/hGVnqFPvZq2fh
NRrH+pks9/AQov/xOAbV0zQiER5nyn03AKz+/FW7K8GmX/+taDGvaDADXrplkUzNWyy3kLp575wR
OinNEocfA4OfLRzchxf7925cb0uCKK27b8SVRLN4Rt4VrrgXLKbxFGwGF5Bm6yxjUo4gbA6BIzIM
5qJDxlpnWQRH1UsO/ow63fjHposYsBCc+mQQ4M25tW/CS3JiNhf5zFV2obQQl22n8IgHvzDAptg3
pv+/qecvY8utKMMdzhQic0Z6ibsxmikY7hgE39kadVz0CFqQLGhy/QWnETbRmUxAk4+YoEfHmLkO
pIEgsVYOYMR9yqS6ASVvi3FZs39GN/XVEQXGCst32qb7tTvvquJcz9LJC74Q9KX55iMd8SvuHt/r
rdIhuDzYFCxpmueUHhKk2UaUJv8Pu4E8j69CZN2m4OQ+89Je7/Z8KbkPRqgXSck7Wwt/IIbtC4NO
l/OaEWCxieadhibTgwOO8gTQB1OZpUZtxAlmlDWPPRSxqlWydBu5sj/1vygxyKuPkUDJgKNynoXh
1caDIrTPou7Zk1O0N1rr/rrxe0J6pWnQkHqoI0qPfFYs3pkrYm9JP0MSh0TLjGXVyJAan4xEX0o8
ojGqlM8h29i0VS/Q6htYtoKSpGGF5uJrFCUgHqvJZYbZRjacEhyul3q3akd/kZ0hAr+/6H0C9k8W
WJW0jfeZVOOJFPgGl4B3BKBxrfsp/D5i3OTMvqHaFAFG0lQ4XVteWnnVNTTFc5pDdtbskfrCv7oy
YbGmkcz2uZfrm0ZZEEAafqN70d/sZHu+z48NhmaTmiDnvGV2ePEu049ruTc5/c3LVPYA1+em6saF
xJ3AvrXH7ExmGjI3GTTPCtWQKfFZLL/H5hnVCYQPwBG6oivZizaCaYWhH0G4O60UVxDl8epW5zP0
D3lLhvLkb6QcNJTHyfF2M+nQRcYXEz6lZCFTvxRSS67W3ebgRoZhMhnrM3yh+7sN0blTZ4SZ/I6F
wRH8xETYgqAiR7VaGCCFVoI/1JiSYHosL3wEZIaboBHK6b1tk+FnQFFsC9UdCP4fjGiebjTvnx9w
WvV5I2Osy6I9SnJCOg0ellkUWYxDrMeMqiSjyMSBCcEMffuu7NUfE58813isjrc1mGyxylc59IBW
IifSSp/rQrw0ml05bZtiSTRMMdQ1vdP0ciYf8sttA6V14jq0CzObQVoVYwm9N6tC5IkFpTg70Yzg
UwavVKlCO8EsshKCyOKxLbO7UctufYanEnDXotKCLxftUPcRIaRDMcg+fjDIT4P1iDu4AtUK9V1r
r67+8LWU2s6rSphWcpg88mmjkvWQm+7eqy609wHhUuVMbLX9YxLrXsrt0nxgevMgOci7b/SBHdIo
VuHr++F9lZBrTkhIF0YyKJTDBVcbC0EvFmSuG3Hn0jcRMM5fr2QcOArcf1hDu++TSZRhu71kq8Om
Lb+YKpkrcQ11swQNEUtz4LSWS+dNY5voL6JIf6MxXaUiYnIDcp5ByoRO3Ltn5LwPYRJiE+REQGqB
ukgE3oDfCMloZqIXYwYMHg0HKK/BgDLB0ULEVdGnJU13pnxoaMBgHC09CEOl/RdnLRYC9G5dUwd6
0Uc+9NUZHqaAZBWD4QPTwcxay17zn05ocV4KjTjAZPJalY7HXd88KulL7NCsQTEIWyMoVvMKw0vR
HUKbs+iX1QUNbUoKThn9r8LOYb93hdnBz88/drtU0q2XRP+ouHiqHwW4ibX7OEBdUU6njORdoWJZ
CMw8BD3ViqVV0ALqaIax+cb0B8t5VlFrMjyMQ0qgTT6uM+XjfnRe4o4WFjXKn9qS2325Bl14QGrX
KSJh31xvGbOxnudPsvUltr9lldpMX0irxMDwvjLBai3diwL4fBJRxk+xhyaqD8/dgnWw4eWz+jax
ygZgCGioqzmzPQtF5a+F+usa6CSUx4muq6HI478BxF6drdHdo9L9hOIgWmrwgty4yiFbFDEyRf1Q
2dxEnrHkRSDbFwgj5fqcuuijJBPaNEcDeaQDDUFnN5wM9gS3VC8BGA5QzTMjvg6sLlUFgfIqYKoW
B091gfnIjfeXy7CMARfFNcsxEqSGoPVpg/gjY/YPW+h/Im14WW4qdJNwZjywz4sGfPxua9JuHASz
M0EXMXFDh8CAui9F9qNUF3gWlLnCfpNIifvdTBYEB5Zx4FRUg4/oF2j2b3t89UA349RWyg3ZC6cP
ESE5K8jO6L4dfQ/ydFi9yBnHxlbxd7cK9LQTL1z2yLn25vJI3bDGFBx/yZJU6QpLyvFOp7raTUcv
OtdC7PXpy8FYnqEEYYodRaLtc12y+W2fg8gsaFQFrzl9c4xvKLKkCpYGnZnSfB2lm9aNWySwudQe
8Xx/owbT3uXSz1k7Hp0Aqo3+TEJkps0Dzqvh8WFZ3NlEYTCcXkkA+H4ZRIBNP21gp3BvHMoBPgxM
94LHJrjw3U7eON0NFwp2iR4dAvwMAdJp0CLhex7EgexZVsfWJMbHyBAaKnjF15AWj6QQveadjVe6
UhOzzJ447wQqdM08fzLcfcbtIDIY0Fl+QXX3zN7xrh9MX7I/9SQHR453hvzB7fWNeuFZdx2m1S1M
EL0cjyOL1soBjb16HDh3dwYlMcXV9aHx6tQvfkJ2ndohXYb0tGMRMhsLMxt/EJpdCgMMsyaM7NYr
VKg+1s3KoNVHi+QYJDRIyuRqyFgzA0YpRqxJEVswNsFSgnQaHHpAh2h5jxcGFOq3ceMIqcK9VULo
mDbMUqtHvWsFz7SxdV2hQbxJeb2BcC4ylLh+tVJaPkPiz+ymoj01VBF3+VQ5qk07rGgkH745saGb
HwFi7GKlH1FcNIaEHe9b0CF4pAO3EyVm2Ou6WbxGRsHmXHxOV41/MhYXwCPiHZPP0k2lFQiBTlS2
pzDZsblXCVskuDcdKOSjb8u/O9+k3iOTzopVbmgh2AkbhSI768JTxgReWJmSLOph19EGO2PbbxmL
mrhad4w927vjDwFHlYLVpmMYQVQjQ1i6EpXer5wkTaVbHSyLzH2pL2HK+NwA1y5Yfwd41La81bHs
KWoR1WOaVLUF1dH6S6L/DQHX980rtxY1T5/E1ROx/nbJXgbZDTcOcHcD+lRo/3XVo8PNI40cFQgF
k0EpeCjZDAFGwTSDVhcxiRorYNdcT/owui2t16t2YTrA35xWttEpl423Q8ly41O/A/peirJushVX
xgVvVk493KbZTxVoYbDzyOE/sMkjVHz0DfMO1G5KA4Oh3lsLEcDbK5QhdVjI4GOnEwQoUf3DS4wy
qiee8NfDi9aBKXQXEb+GGOXZs3o0cxpNzyIs1H850Jt9qnhwt8tLL4Geg/tKH4uC1ZSP5504SUgT
7SU2W1Hdhd4f4LDC4TVxxnpd+CRBNdoq4wft3XBsxNnMYWLU+Eg2TRlK8Z13X7HZfhOqCKKdqWv4
+9+lTC2UzE9wcuhAVTBw4pqnMTXlIVao5r6pbu2FyzdQe96ewICWyp4HY1yNOGRL64wQkDiQe000
BtEO9hFpDdvr/xneCIjcNZLtHfM1GWjbsCwiXnbSvb3v+4Ff9e+2xD6J3zvdzGQkSDg/OIl3dmt0
RFYDoUTU0paVOhySnuuuFe04TB2jQ451fza+gr5mzBrKqLwqzKuJqoBon3Ypo1st/j9RbIlKtlgO
S7YF9Mp04smeqaGAuVjjZ3LPzBIx7o1maKRt8fxaHX4B7BE1KeaHBqo/jc9wLBtcFcjdYefFWro7
ccg6saNg8HX5szZJw+UMaxdDK6fSkUdwF7OZoE/mfYkdaN//U7yLG4i1we0nc9rmLHr8GNRCsEyz
QAIEqapc99sxXEFfIWTt8Du3e64ZgRge7zNJdE2J7oKxEsVNYBuE6sqK0D71Y1dHZd/tCT8nWsEL
ooGUtN94LLm+UFdzAsvIzD4oxmHYWz+2tET+6LdeDhhxQgkJkFVhnkbO1k9Z/RY74MOoMSVaD2Af
SBcwvwVdqm50FRSrytDL1zJ6A7qVxaBy9VxI1+tEr56V9juFVUFeuemCES6Hrd3U3bePB94UFx95
7MIK897aizwRKHSIsOoGUjaoQofdhWrCoBWVWurxU+96Ad9s+OzWhDJOuB7owDYAYtORPaBipjW2
FoBf19/pgTw2bSmTPYjUlfw7VO6b8GgplvbCRbcxvL6DG8igCvPbKDC/n+NKEtNTeuEiz99w1HHV
3WY78uRdnWvzFvj4z9cndAj10kl/mgQTFURPK0bfhosUBsXv/MYKc9UHodYzfZqzcS9TUV7eaNNo
8dGvrUUuunbzXPLsS7OYMUny3/KyXkl5YXttCZAsAdIzRH/bSdXhkp3UdgXzmohcu6BhR4Mi9Txr
Pgz6x19fKibxI85gTJOFOSwrGygrfahb3E/BgEEzIYkvurw7BTuUaCPg84QFDIyYDQOAEOnN5OC5
B0/bQ9aySMPocf1xX/adqvZg5222CSHZ3kKH+ZFqFdO0vRWLTQzMkcafPagFdHj01i6Yrb7/KRMR
iyfHdCFj/uGDqvWbgIzomalCsxcpwYuSak8ArNzoRehWwGTal+mONBYJUXj+NzOfyrnyicUJ9UmH
gUMcqELDK/RShirr+I5NRWFz3AC7yDqGcebiqY3Cbj0krl98ZpexC+HItcQPdpDRFyuaULQs++VK
l+w+N5ZG/Jo43yK1pxbxSJGnH86mCAJ5zHMLObN13cbfvbHDKX4KNPZZ7uJQhPYjBmyQkpSnAE1G
O48Hy2zULLu+7MTS1kXLvfP95fQHrtosxX8CIKX28Gu7k4zWU9QnxeXH6ODs1JtkvYGESh1gQXOU
UEyQOWfyfZOgFLnaPHgv6xg83j1BIsF/T3SLpcglgmOHKAphyvsXIxq/9ICQDbtwjVmdyK3wVhWx
2Zun+MKG5srAk5EqPV0Su8Mk3ZI4N6Mt3oIrZVcWINuOzyL0+WeSyPhRZYLA91Go1/YsbAEv+KMX
J6D+mhjuMfh0GK7C/bQbGIQhSgn3scbqWZ+FgMm8CnQJsDsLPsEw2p6zacSiSrA/hrwG6aIouFka
FS1y9cwycFhCZHa7zKyXLmMmuXZMtLO/P64VxgOfxbrYqtLQhNqDbilRyLQAydSBNgGCIefwS9Bt
H6947W1Z+hJxULX4MDiwczZr5At/JpYToX3o+1fIoZ61qxBAwMXnhoaoCE+7DyGNxZW/3TJORSZI
z5EH5KO/qL9GW1x9gFZ7sXFy4g+bLOsdBtmN0cUqNwbP3fqQg4OBSWWzmoTsHFa4RwMOJMPlXDVG
OZfMX/wXNQl7Xxt92HQwfzmPm8QCYA4tqTbIvTGCNDAMLZFK+b0rPVkNnwR76Umh2xYSifemh0pu
9zQA6IVPZa5cUs9LWW5FDzkmIFpU6xhggnpEVFSnriFMkevj1wFTRrbWQvUWOCmSTI63DJjJgeFz
cy6agWXpNcO2gOLu9SQJEruQlZv82fIQ37f51Tbn2fPVSJWm9yPXO7G4YQbnzUTv/0mz2sg+6MG/
iPKt8wdausqAvizFjJXoBLidqItE8GUKZcxJfWQG1cj28rgs6q+gG5ik+6pZBHl+KfhWK/7vgPkz
8rkmyVklL7vg0qmtDyVWPjv4WmzW3yd47qTHEcsatfHsEmpP++6PzXeXwZVlsyOwR2ysLFgXwENa
uZVNHaAMkJiIzsYLl7wvqS6u3sBmKUr4sllPD6jQFO8lv9ghmVNqRHOHvy3rsQLSgiKT0xSYYlXH
JUOaWQ/H+wg62ypDkzN+ooUFM3VhFA3rCy2ppHI5WHRd3s4fqSUbaKxpIV0htYLYeLNVW1gd1+Wg
JPHrhEEpK4gtYGciMMvfEAuV81at4J+1RuxUJbLiT2uF064qjojN0cNSGTUG9h6fqX5IPSuF2Du/
G5s+yyUnmB2i5ZQsCEv1RQ0DIpaNr2toBjbB5XDybWtXLvUEI+JTFaDsx6Z/mdVBQa7jhgS6s3FC
tHjstjT/uvfONrNWMQ80OwtNiY+hbbUeq12VzskfNPr+4ACKilZhL3o+/RgkKAwA0yNbY/ari2rf
tlrsuvv02s+K2qlRokkN95/V5vYGh3lAMHcL/+jUaUsKV+a3StKSsC9erlFiGmCIcayHoOs1Yjor
lUcqV8XttwP2o/phEEUtre6wFua7ZGEpPcOMpSFXEgvSpphgu3Bjpx+huIx5xF3Rq66iqxuqaw8d
7oeGVcjUQ/V04GFnQYVHoX8+rFXStXrSLArhFnwyQZoxv7luR54SZos/dDcCZUxr50mi/JUlBtBJ
yM9te/B3+RpvSyAx00q90J97bPvun84061Zy+kUlOmMeADDq5X1cIYqEBkz4Mb6rnyAgXG92Wz4I
I29yNrOOCg3VPpjFNyKgpHtFkwp0vTYGp82B01vjpteJ0dRLJYPZs8nrEzoqs2v9PNztzgoXy8lF
Mi91bBrYlbFR6GtRGOoI675XQnk+ja9ZzuICtyZVHTFSYZy16h2VJKDVNo0/k5qebdlp4NwccKPn
9keWJNyHnm1UB6uq7xIAQ890nM+3u5HnIrLmCDFyeFqeJLRiunyZXUD0aeQanw/z2x9RyxQ8y8t9
gYWlarmf0KKg/48wRt4WB1Y2+IagWp571hEWPKAjZRO+vqO24rB46vPnA8WeQyYhgsxKBT9cdhsU
wRmUUsFiz3E0azkOEYOiLm9hzbOl8euU9gUU8hSbMgOSz9wATN3bMwcEha1AxzDprfQ7X9KxryEA
dwL2dnWX8lu8PaydODe3mcSre7XM7TL6cM7sKiW9EBXdD8UXznRwb7BCOjbin8V0nTZYt7/urSZv
2CM/XVdEYK3xK/c5hPZ64x10/inDqkFbCpotk2wIc37ZFXosNb57N4a6eu6anOYYz5QMALwAhi3p
VgYxC4k+HFUwVbyqKx3e9UXXu67gHnifUcB+uNlKoy2HI+bJ1Hv0jyr5hztjNQT7P3YXnTzmf4Sg
8d1k6Ex/eunJVYFMQAgdUzwj+I3gXIfSwOzjAEtnM0KIMK9Nz/DCM5rtNiiDlfhEwurxAlZszayx
FceCeRTxnfqjSESCvJzjAAkE6Ov1lqS1Ot7cCXGNP3y1nG7nTpOdqE3J0dWVW8wPXZQot8r2KUiG
w36Vl4cQ5RBSXvNmThbg+zo1vpUWBRzH3QrjMh9Sna5UIX16Was2G/n+ou9TLfKJ9tHeQSHNPSmZ
MSphIiZTtZnqud8kjgR/A2skYNU7PP6bCgqtu6CUZTY/fBEjI3DYeWlXRq06c/nZtC7oV2W7IZv8
YFX5sWkiiZyG+C36d23a1co6ayDcF6Pi7HfHSLvvbGV+Rb4+eNdGy9CnnjbAm+rF+sv7LPRPfjHB
CswQmReua2gk957I1c+KZJvegYHBWw2CFHgQJtb7lnS2acXqvjEmJPGbh1sCzLixcvdrh13tA3I0
ClkVa7WmWRFXvOsXTkCeMP5ZYj6PMo8iWGpwvUK1WgxRMG+EKa7Oj9jX2crSbXop/OkirZz9gaal
3kJYHqdXrytX+W4grBZLW+2tzJ5wolt5RcxA1e4+mWwfdmZsIfuehzSorFWqGG+Gffl1fTfOs0g+
pC/4+kq3hVz3j6e3lmUp7dqLfzEhC/tO3trRO2y5D1QUmj5PZ4t5GRiM2Zg5l1ILzBYk72RHfITD
/WALOviqBkYhNgKN75nqhOo5Gqhx4fdcq7wipeCdpx+Hc52vXksASfxaSVNKGMnqaz5wNW7q/ZAu
HhLrDzs5ig0AytVeJXYcrIioud/FzvHPoLg3cY3cjVcizuVrhpi5CvVOUGvlYdo0wnnPCA4/0jfy
ye7s80yKN3QhxLTwhIfgp/SvjsqnLBGs1Wy8tJr6apSCjOR9Lto7Yw6iBIfc3/ghBWDE5KrtWkvu
pj/iVSA3m7BambtUWlVPPLSDAbluN2onlepRZujTclYHZSpUKdJRi0Cf2tvkTW8gvKiIr8R3VQnx
qAEro/e+5gWVc2wS3+rDFIPvgU983lpmrGIEqPBmAfIt9cmjIyYcYuxpPBYRFjUUIJiATkrsiOhL
sFULMmy8JDVzGHLj56BVJL+Jebq2Vp63lN0uyP5yrRzrkSsjMTcAjayqI6BCmKs5pSPzxYICfS6a
fWufZ6gUrtz0+EhyoPYZBiy5Mj3by3bVnsuD8byAAvAIy0j2W6KOsQFIhiU4HXQG6SnsYfgpSGf0
fwlrJ/HFXGLOwtpefyRaCxqLv85Xkf+4jWGdDzFH65sj9JWI2PtANOvQoSEOpTiF2pPIqtAolxQa
I6FCU2bi/wSx9rslNDVZ54yaV2FnBFA3BLfarX+83yyiuu9/x2J43ZZ+bLt/oxUQLfWwbAxNThnA
yADUJNIReK5VHSSiJxC3Qaeu6YmepObipRYHxt6NkQT+ZaEsW4hcjt8Ky3Xnv14U1PkLfzytmOfb
W9c3GbqojB0/PEpZtkn6rNMXZ5pcuMCMXf2dSX1CykrsQZL0MerSUa2RkXuyOQqS/Q/RqXU6gQ5Z
W5yX0BbHGsmm4OcxBvRQH0stJk7nQSDWVxr9ty5kuIJx0Et2RqujxopGnhKq1aREY26UnLz4Mc6T
t7R8cXIxZv6gowROwFjtWMj6N3emYeYn8oGWX+60fpGCKRHkUGO08WjAZEljTIadSMfyw9RY5dGm
F83wdbImhPghHU43CKVGmJAZKZfUYSMs6FBq+1Y5/mK4puVcT3djCi5KZq1r5eXAHbVf8+SXVq5X
+uUmHxoEto/JRcsBm1YLeYLYewYfjCJqZiAfXT0FkTO831ylnilpp5NwU1uAk9ZQijFUKb7SuFFR
ptEHH0S3Kd5w2Oi1eIvDGDHRtcyN2VYNGIYPY+5zC4gIAUlmRmwDCEakStR0ZmekSF3nuWr+zZiJ
G6qt6SuwZggx3HCksPwipzyO8KSd0VHxZ/3qbYKp6F36Z3gSaej56HLCYqZIluP15r1XZqYVcTr6
QAoAdr/VfrnCA9M9RPEFHtLyxaxwkuKUyXqBbrRMUdew5cRAl5zeLJbt1D5oHPlzWNYNk//VQbUZ
GHVY0+PMEEDLu++Dzx/Ged9iDysaHdl16oUBVDLxjGqyA27dw6Ew0kEwLDixG1fa29NFz3j1XRHg
pN7VPfx9iBJ41DpvxgOQ559aPDzMYsDxqI1yOriC3ILfh7WrUQZSUaorUDjkqfMKFB781eOJhgGX
v/EP5eltiWG3kuQZeVZMs05IFrK2QDJL82R77ljbwIS62Lo+2MFpMjeilLDsaiz1XSYl4cvrKo06
H25dk9FyUJy2yrUwKYSS4shig2lkK/sj0lrugrD1bdIeBfMOnVLhFogshkU9FEmb8QmQlfV0IGYF
0zC4p5hePqd65jQoRxipCY001IeefZcqwMcRn+UU9RX3ea63ZJBnYF4qLfvsJNmwuxJdtS8IhQ73
hKag6Ap5yKas/UJOb7uAClkk73xhW+wwk3xpx5FC63s4u3OjtLWzHBtfopLV1OHwNC8N981RU8fF
QhHGitiGgeCVFpXGZTq6sQxnr9ROyLe2JzMWLfECUhQKdrVC+4hAhuvGHzay0wWDU09vivDKiIuq
TL41Nakez4IBCdJ3FqLvTW1krJfKMebRNYs6B4VehqSdnJ+r49pBTb//4MybMcoOUMpPlDauw+zW
hXrV2joco3HPUZifUs13xKpFXFO4gvHN4CVkedyNJsdcKDrJmDifQKt7VGCO6rzp+R/eu4GkIRop
XCgvj+w9p4qvmBghZW35LHr7w/gexlquVghl5vYTDH9Yh+lS5bNhasQv84L/LU0NZ9bnJC3rw74E
zcMPizpwjQWntF3uKkxeZnRv0K7LkwSSeHPXLBHBjR5WJGFb0SpSJtOazofuLC7wZJPghGCtUVEH
OiL+oMfNdwe6MY4PQXQT9b0DATh+7YVQh/NUxBe1fjvV8CGu0elt/kuKZccAxgnXfusnd7/QfBME
JTY6jyheD5xcQ5143ajc4YdDQADAAK5aROaDERPaZzr9HOMw2gCWwY+QktRj8HMtKZvH8IdHNZBG
fKyb+iG34C2x3SI5/z9M7mKcWx12p2Ijriha9oRJ8bdpnYRoYtgWIe9gh7KF8xpI85IcnT98LLjj
sKG4i7K+9qFYPEO3RzaPfEqDlUCcCB2QcXJfkw1j2A1nHOnLqhz0zx23b2PtE7UORQhgGww9PjLB
jfe+wgZ0iNnlcOlhorFFabJYzVSc0B52R2Ss7ffeuPvenE0F4EVuPIjYDDKZGHdUZjf9CTlPXlwy
IDAhbHYrhpN++MDgNTBPnhhLismbcs08qQfo4s/CAt///k5K/Lc4nRqwXnVEwhmZaJQKucfzQoL6
1zOpd32jmVV2HFFRcMNDA6zxd8FV+USKIoAPYxCy1i7PTtGwfR7iC/6pG+GG4sjf5tuEet2+j8DA
Zj+kFsjpxkueod++rkrty2AQGgUvv2+qetlH4Q51nOvGq4puEmHisc2nwQedSnkRsCJsFkTbnBJs
k3TSnYAoO0kUP9wKOiNMKHgqeHyHsim7RvkMFdd3yzMXeRhtUuhdqj8V4iwsdVLE/O9eVL+oSJCQ
iEGKQx5y8rcPLzpv3aCA2lku1PyqD3E92RbLNordji8K5YtEc7FN3MoRF8jx/VPIsdfOHP8SJlFA
P/JL33q1fSo+L2DNZ2vLZAAlXr7IuDykDHaNma69WlYSy7Uv8A5+r5vfhfgVjzBJFu1al8FVf1+f
rHrTot8Ij8IggOWXnyFZuRkODgWXBLFEY7/SBIJTZDnz7OL29L7s0+YHtWCoLnKk5F0lAgeZpKs7
4dzEuDhj5YTJXn5jy0qLNO7tdsJQd44z4ZMRjW0xeCPP1ubvBgVyuxbV1Le2GhmJhE1h0/KvAAR3
YjN+J+V8PqrBwSe11+SJyRRTj4R3DhHZ7uIrFizcA+4Wguea+5DGxx4tj/mTnRAhuhN4YEtsFkae
uA7f4d5dkOijuTUdhnR+y4K7vQnLUf6oILVwR8fRqCb3DyW/Cr09uTzG5A4aj8GRqqB+QDCiwKPw
erfHdEHy7+Ts5Kv5xLJG+AqVfuL5w4Phy/dMr1Tfs/EidnkqMP4HoDa2H0B7t18USH0Meszsi06C
Btl4roSUU6mjXCJFrUK34Amq69O+Sh/8vKR95JI8NLNuzQ44fz3loVKbG9BivghkpkVXxuBvSoYC
B6d+t5qlbLQnFZTceTfPZnI0MN4r9IqzivBucYUKE6Lq746n8Dq3NXZovawBYDTf+aLhX8XCjXM5
Wrcn5vhjVAlN5PDRxD+UUuNLG8bs3ZfswmXCle0YmqVtY1pKGklIPdhYzgBnPEWWIkmQRlCZxS3K
pfrh+GLcFOwiqSq5jL+G2cKWhLC7WOLFiXjYFgOxorDZ1/XMlDQNLe2v0ZlDCyaLnkaUzcJ1VNcL
WlhUQyUldFbj1nL915LIcvH14Wqh4m8xM7oNZ6BlVaNsmS4eUIhXYg1iVQjGKTrYsqK4gqv0BlmX
dmKxWHnijvvoNCt27KSxiorA/chFQRKIlONS6j9PIUygVHRojEaAbSlVeaxvO3lIHzIDKisr6Ylf
xQCt14BenayD80HZIc2WSxpMMLMczcaczxlEWusRZDIMUJXkaNnis8O+nYVKHHNLMBGmfNc/KRom
2LRA2lp5MfgVmyiyLN8lw+vFiGCpcellWoMeaXUFmtV8b+fohpGs0pJnjEi98FMEvMxLS+56hS12
vfp2bEyHx4Jx1LOtqFaxWkJAYPvb6pxEa0lWUyHEhZxcJJ3l+O0emkHDNB2+XBLgzkZI9KfYwoX/
U0agFsZd0qqNt0zSx//gMndBT7PXzX7bmXtxJ1JtjCpMztUfDa1+r3e6E1JA1s10GOflZxVXS2LW
2tQWQ/M/XjfbBpbUNZvbz3gsxjDbfmV0fUO0z21pn2d95/VYiEn0WWohkSVF8jbUGcJVuY2zeDfM
1yY3145viu5PyCqssuF8phy25VFiyd8Sk7kcxrv68445eWGi4EzZiGHve0S/32l07VoLWJA1JQY5
mgNMLK8QeSPMc1s8wOIyE+RBqmtRv3+I54WOwQxOK1n/vL0ucLUZ2pRRzicKArrZdukCmJzH7SNR
v1tBM0NEZSFsPOx8ETP4308FR6nmbSVfvaAkvpDsuNGObTrZ63gF8JKbgoukNlbYKbXAKLoRx6Ht
kdU1nfkpo/1rOgJAkI5IGeybvWYcdpOVwVJHkRVTV18lACliiUBhan99Ikrzq7en8aSmj7eUgTq6
so3DtKdUWHfGQDfsH2ps49dZBm9ioKGdcyX4I81Q+LniLtWbIWe0epPFmfRWSjQqPliPdy8N6XXO
fslR3kiA28NvvXA1HarsHE+FkQyTiIBgJpfbJHfJs5hgL8tOhqnYFSU2k6UphzyDON9RrImPY1mL
XcwzFFY19PMxODNpB9nhyXq6e/YLmUmu1BPoC4DUU4QQp7ykfAnv5uv3C/18ITQ5cBNdqkmQI9Ce
U1TZBxSMVNokUnFcL7IUxY1jGBK8uFexR25Hn/24HSEKHGqq6w8BJO/VVN1YDWz7T6HRcBh/DwxB
i4W/ywAU97+yEZWc0/Po3tvzbzBCUAQIumK5TyNLWjsLPu9nokfrKVSG7UktP+4Yv/Gp2xWNC9/U
FcLpoZfyvEm5xyUOPJX13hcf/G1GXiEpKx/3L6MeqPl8jd3Gz3MecM6hIYSJ3HmmAG5+JybmWEbs
D882o/mIb6vEHqgzXa8TROOTR7qB3B9auvmNZ3vZViwHD4ogrLH3/oQXvxptgF/AAsIwe3HY9Z+r
EJXRsDyPsYkpIo/iZCwcySUsbZ2VPYI+V9EsIHASPCmfkwKyE9vlnbz+wLu/sjd+SxcH4s7Gn9l2
1PQ5tiy5H2U/ZCzsO+95UctW0SkOE0TAUwKZEUCInYVroQvG4xb+Z1vHvNFEPr/478fbYtH4nGKV
j2oSEQIxnU/iukzl3TnPuH4YcF37oDj0X+JaA8eNGB5pis9Qap65Wus/78WoJzygf5i9lVUXu+ot
/agq1Qhw7y9w2QLlb1QnsPzLUtRTneM+6zMIduJl3Vu0ltv2x5K2i7S8+Kyi/SpVC6GXWHbLaN8D
yMCnbnHWQF2c6e8kKhw1lcX8clv/5n8ynngdF/730N8vYN6SrnTQfoEtUlgJ6aO0CYuKHk57Y635
QO6+liSs7SNTgXQ3oaY4rP7i4wkUHK2OxAc2VMK3+QBi1DbF5A4Jdlle0xMBllhLSjs8PLHujnXS
GLbrbpDuTCsjWncmjoWy13Yq5bhV6cUlYhC3zuMXe1S1zcLoYHVYhYVTdmZ9nKmAoXdzUFjz2kmI
hNzs52/VH/uNcug+kKZz3Rx8z0nF2vowSKFNRxi1oN/DLjWPo2ClQgFGdUANwcR7xeAgvBXBwCT+
3dsrnAdcJhmVahewu5sb4R1hpzBzxBSGXM4oubLKNIsAsuRNdKExcZaaePa9rzRI9IO9n7J6F+oe
a5HkvdTLk2Xn22k9WhI9jvsxlm6CZSktUNOXfUGj/BAEVxROCbmcM/rFdsUzqrr17sbeI/XdfKbT
s+GsW4QkRf7O0s566zfTtWrPQL1Pkp+HkQowLUlCUq/+rtQFn6c+Tf827anHZIsF2j0B1F7CPe07
uZpERhC2sydZgom7WeQyqoNRtujLlNsFy7B+5r/sMoK2UoedmijMcSx9SZ48izaQtcq4GIGkhTZc
ayxYyHpyjgjszuXAvprRDSXFpH84/vYfUiyvjOtKdepjz2Kfyp11byC6jYlpPb6lmyHmZBPbbqk2
JYNcHGUpE8ojMS0pP2TXhdPbhbqiaGRvRgTcPuRJ8hPvNFVPKBVQ2Xp+tsuZebeY5u+NChg2q6Xr
PexW1Bzj3vzwxrIsXXsTUQjTT+fFWpLSnmT/2YjhmG+unv+uuF9gt+6KzTOGslsikcgNexIfb2Aa
1FoPmxixjP4xIUZQTtAJhCmGu25airuyEhYZ9PY1MrbEY3poz8koZMwwb7t/LXADCYtO/MSnT42B
rlv9FJszsZoSYcKSDULqRF7VqNv6BOdE34CYBms4l2sctGN0szYfRYlsCzGEy6slOoFPKLw7FXkX
je8uXFQGgHM6hsFWtlpwPSIkY28XLt5cwKLmyHFAVFc60K8Wyu1dLogZQItv69UahqIZfpouft6U
SUF9YkSXgIJgiDmoXStqxMPVLr7StEQpid/e7cwbIyuc/Ce9qKqRnxYYZfAZJBaazGWobWKYjLRs
VCenMDC0RSoYT/cae/8G7uJL24+1+bwwqzLRZZsw5Yn7wQy//ZCcWdKGqXD/bAu0c5GtGAII94hZ
kJHeqlx/9oLj5iZ7DNvyjT2/bff2zv6xqh26HwIMdxLcsz9y2Z1kbj3nQj1ftBg4SZNaQf71kDe8
VqRyiK5kuH9Zq2foxBOtXrBbRMtXo4ER+0oismJDwFQhYeS8MOmkNsCWYy862EFBz6cLBQHP3gcW
aYLlcppUP2T6pEiP4Mwh+oUhUxs6uvW9Uvl2eD4vrMOp7WHSmJPaNlDj4qbVkMbXT2LA1pEUKElI
e0rFp/0TdLq/XD74uF4c3tzaQRaatMsze2C3K76rjLVPvk4gN6oCEaY/Uudik3vH8/5SgMypp+2u
d497hFlJ/aarMk13mb3ozTIjQvNhFL3wG8dXuKjs9yiZitFk1iSoHWGafcHAjFio1Z5a0tmKBbDr
BUsxPIpHqp/0N6ifuN0Ml1J+LymOzAnJFElQmdFbqolWKloyhykzDOo31LDeRJD4b9/8PzPUUK7q
xEX+h33ZwohoWqFVJBJkJo2YFtiAoh4w2yiHIKKxLUhYowCZ/ZOHK6+DugNomDDAToFJdf+BW2EO
1PndbLAyDWuKdrimpEAo4bApAbH8DoAbfrLvUCFkg/fgtp/wcRqCTncpGhdcMXWsvEE7yaV4S2NC
HcGAqIAFKge4v5GJY+xe+1g0lXiO60bQ0dezAh+cMVYvkwXgrxXwV12svAdeg+ji18GqGFbqqVZz
hauK04v/Gwp3ZtrXZltp0sKAdvvjDqbDDO+QtvQ+NDx6jQ281lDNTVbjTpkIfcjNpzcXCWoytWnD
6cjQXUFMaon+K3K3N/t/yWx9TSgpCzpYoO5nxedoSwvoOtoiZCrk71ptnIxP14fRDonmPk740vF4
z/lHYwP5E7clqONQbsjUCqkOFsnmZmrvgsutmPYbILuR8QzUOHVpw/Gj0KGqzoALFHf2NdQu1SgH
iYQbugwSLfOJVuYroaowUUzGTj+6G5PdH9tlTaD/3cBJ7Ff8TqIMp2CSTnICxtVgwnheSC4NG2Kt
ru2l7lfm0azreBFDaaHG+big6WgCHhzgjvwcvP/zCap2Q+Q0p//El/wu6XWWfjLBmldAfzOjSgH/
1S7DPaRuxME0jkIXkPYhMi5Xvfojs7OyQ1AJKRZIy6MXz1L8WcV25J+IQLi1hWpJ13ySuCgEDkaQ
hgPXVx8Z/sBbzOuqPpseMDhR8WrHlAJ16fkRCazfnQy7kM4golbqVn2WghxreMTQjj0/sqhBG7wc
Ed4p5Vd/1b7j5ggSuek/qpQEH6hvK4eX2rQ684tMDfy34oDXUv898er/BE+pcOiDjZuQCCOvz5MQ
GJpQuGYZEX2R9LnhPADJe7W9onOSZ+FaO/WSQUNEtRirHwWiHcfXVuziQwWFjihEeBqbDbClZwmL
TzMQqkvaIuTctpg5qEH4pXubG2Nzwws6qNTCYbOcmWjvvn9TyF+NyXswfD07DfuDr9k/Dma0zJFI
AkCiRnOBimSovhWvwnhOE7Xbh+McENkEytZ6O2I4QteerauiZ8bLQrjz2uoNLZcyp+vhjZeJSljJ
EF01xzXHLGNKyCZpa0EevzmG2OOOJT+9KgiRNNpuTrvaR4q17VIs43XYuzDYWqbNyWeezMVZQCfH
hM3BniDC5MfY1cZdzwfd23Rniv6XLtk6K42VqHLm4zhgRuwTujxnr36QSj1zLySYAwDuQCHaYCoC
vhYm4PYGD8MRauVUAcN7uXXNAd9hAilduP5AK2FBKesq0Gis+IpfGpYHrcj91fGt1tdK2QlU8Bk0
sffe1bBEhKV0aWj6K0yPRWEXvT/sgP0AZl0rVzaBIqzdAjE7rRTnM+5FUpC9EjnLZM6Khn62ErH8
jtYueZ1U0OmtS6gYbXQAxHB07M5v5gDNDUvkCtG0HKv4EfVS7oPm98WUmz7hhPaPjdRdvXPO6FBz
Naup1Thv73auyu0ERUo0vLxuDUm0Oh93sQnGceRJfYWqK27uNxdblnlpr2AvK/REo8K96mcZeLoI
K6X0H4U70idPssJAI0CqsueHauPK+0GF/RKPLMikDVtF2wLRnOTEMEo5CTWLNkkbWE99G/IqEXZY
HJ56mjONi6zHl8tEEMpn6fQ6iQOwFThDtYJZhQC7p0jsDBfFq49rO1CRdxKVlkuQk40XZPTJ74J4
GBBN7MnhIEi1kSMUYFRnX/lWMJufPrfDWiDIAsgdy8BIgBlUB9CzHFqlwlhMMC9e2YYZCUAk3LWD
7EYf1bsFVTgEjdIQEWgh/PHcfin5aVsM73/eiYSFjnnJ5pl7gKJ3Wnq8H7mJIKRVk7sGjzVsc4JO
xIGKc3s8XbimyMQyE8udjbgd9TstvZqNG+BvPNPVJuTBw7isbpheW9dncEfiuBwvihI2ZOPZzyA4
krwmYltdYiAF8yWXjtITK7wmViNPI/1hpVsDC29cpI0776Smpf2WmEIRXFtDZJwO46dlkwhVoRwy
a6HjM1Np90NQ0fAXB16m+VS0cfS4pBNhRE3zHddHJ6ukGMHBAUdgvVfrbtCxUr3QyLQxtSIB3F2j
9sQr1VH3BEWTzSQihlR36QrVAEZHUj+ow762nO3TxkpyuhVrUCOR/oAnf1Zqf/o/uw7f7eGRXHVr
PydnIqWpLlVT5VfNxqEmfdYawSghl5Ulr4UQpGevJF7hVhJYZ/ZprNAb+o4SXaN9aOkfJlXn6Iok
9kxjs8T7NRHWGbh2AHdCXSpclpt/ZofkniE6CisJhi05texYaztkgQPLN39dOh+mEpN527atQJFc
xKS8+WDLGi0eaUzgeNx1ysUpNomu+aoA8k9bzOTPvNCGqgXRnBFoUTM8hWqkNglAULSfzbioSSaL
QepM4XvU5NwNr5QbeTsqs7mjBfSkNYwxGckkkGK3R+Y3bCGVeOtdkyOr8ncnycm64BA09HRDP55i
Yurv5r5RAm1DxELNHN2Ecbn0XvS0aOmVqPYJHU91kMIh7VoaBs9JKljCUjIJVESsCI88YpKJQFfM
aHxJzhi03+W3na9P0LxXCYSczXvz/hamEPjXZ4OU0yn55/ORhPuYk9d2TnTMBXtIxdrrhQvitBdX
NcFUVEyzhRCBPfBKm9Zj4+NKvg7dFNAHGHHbMchmXEBkVyLUYHnqjCuq0gXLnb8IBdgVkD/wxLQd
UjOSKfs+w6lKE2uCVrLICg7hfksYB9aioLW/gLghAgrguRUVDRcCTfoXH/8Wi8rwE5Op5ILszwCN
1kNMSEXcM0x5Cdw8l4T8mmxiVHKQLecR8SVDcCzE4nkI05rHQokzH9zwBHg0bi3y0YHuFpgaPnmp
otr0YUFJqQLEHQ2eHWpjpPDw4P9pwmTJtlRznLfLXzjhxbb/6z6wSwRJozTlcZAMPx++lDToMooC
oBeHaWa0aQ7rZ6HDC8gPv6kgPSB3RBoWOKXMr9fnEY4d9OPeNfEfGTCtDc1jG6D0LZIO7OLoPuwo
pykB5jVpa/H+ZTWiWfGW4MNMMOYK++Sz7DMICCwqrVNchWj2YDRgTFv13yp7f3J5OcUPliNMe4WI
gDTdZKxwdGFNC9LP65mEuE+yGIDtVonztCZDe6G3WfkOtAC+neQYbCYXyqCsru5k1+Oe0C+CGce9
gesT4Usw1m0hGM6zCZbAkCYc6Ahb8X7/pEFx5C/VEZWVTsXR8nttBYITkxnBWJVKKkC2oYv4iCk0
WR+hXBeSRiWuxB2enaY2ODpFAG+6KxmAN+Tlv0wZcdhh3b1p8PHrLBlvjKhRPdoFJGQ7tS/voBXv
g2FbD1Er3dESZH8muer0nLjLPDvodlCODd7UnGG9d7chOchh9JJEBvEj81Hbm/aqnsC4gxyT/jpI
lO4sDrrNsgLOunqvJJw7v2QUFxqGUzIo9rU6v6adZkOz+DL1rJ1K4kZ4OeRP/Hxsl75Ay/gH43w4
KRpn2kP4YFPFnUxcTD0XNBhst3TtVt15aLdzsOJUBUFbPlHda/obJm/z2lhGNbRV8/iJjygx8HeC
HN8fZB0DUc8Kt8WDqG0R1rstMtRnEG2jF4xm9iDAGyXV7X585v84803KJfv3ErMrpW9bInRvmR/2
90apdZc/GoKcP07n3gjKKGHyETGTFzxcDFs60n/gL7xXSgfMrc+rUUJ7mJVb2Y56bYiOYwbRO7lQ
HHD+PGU1wUM3WIU7+lsxLe6ErfPDdhftQr+yMgLEZW4qla6e8mrbwCxi9wAxAMIp2kfJ4VSOzHMU
YgwccCkSmXLdyhSdUTj+wyssqzmyWo3nTzbYyYtI1t83daZI4KnjJAIOtm58xRjVpU8XOp6Zz0qs
AXQQ8uKQT5GcVpIOov7Xkyl6bc6d+oufgFRZTNGw4EgqI5fA4M8qxE16Xlf/20I/6rmDNonci4hn
bBoO9/29+LHrLm6xKklq+RzmWSU68lm8aPRSpRSBrK5V/x6N/3tXQGu3CGLBDyyro30myWrZSi2Y
Se+qOlRLHUgLUQ/UZyEuEnJ3J6WR5glagJ4XL2sLDfcvUZ3GdcJBszi83slEizY27ekzPzSGJ/NS
iZuFuH/grz0KqZbJAlvgDRKcPyJXwU8dDz63umZJs5KKt4txcHmNMuQ+NqX4V7ChFSQBb9mv0zUv
4WUZdXr/D1UgAHeIDvZ14GcgkFr9CkfUL1gvgPNlkrHgKj+ZaoIHHya7jniOgeHXW9W4tAR8AboW
c8CVJBlwVkUemJD+nr4wzKAQA+JKGRUamdmYTmcKuVnDyjSHK60NJwkaJ+bt5FlBKB3ZGBiTr2LT
HcrdsHLQoSJPSQ1r3+HYFUY0Gvqn3VB8Qo4LOhScqzaFYH5lkYG6a6fEEtN/NFSasTYeL6qaneTF
bpmbmFLPggjPJB9xXV9P4lpQg18SjbYrR2IMi6ly54ppmv/ypM85+HBzcqDkYQVpS2D8YYJASiEs
PHxgswOEGgGhgrZhRKE2AnmFdty/DbKRlQUs4r9SfNjk6oyvgYYCDkXIkeGTRVpnVGDU3JhtRq7k
NJ5yqaL9xYcYhmT6kiQi/6oSjBY2IUcfyP/gQRudQ5BAJH1SAnhcKKkfK4Wnzl6s50MvQySxcYs7
hnCt5yq0quXyPoCn4k4pCXTv70LOnDdR50j+HKay3DMXEXgTd/tJ/O0LSfFAxNRR5fRjtTYg0Y1Y
qoUD/IqxL8DwReeN0pmZjr0oxkMFN4h1SDCAi+ox0NXuH5dzyRg6kDrcVzdud154zUkgv8uEkpFn
d2wFiq7FDvOZhcGWSbL3Jo/tgiq5EXdQS7v0hdPyJDpZcFVAZkR8hqm7xNyWryDM51J5miE/2s21
lwcDoojrt6tbA+HP0TSq5fw7IXpma1EMCfNpsrUMXwy1zwhy4om4OJdUh6Uxsu1Ktne0rqVk2fOy
gwA0PnHTcfxPO6PJEXkE3mBBEK7b0VB9iced6OQjOcTChDbvPXVBpfQKd136twOufe9h+xwEQqN9
lfaMbxODFEFHMk4JICTXJp2dEPJI8KtSmYLFxGOe1N7soklOOGEssAfXVHG1UW2trI3YSY9X/S2M
bMvKjS1URPZDGL7XQyKWV6gz6ZLvUZNcvDBpenWdoEXqD+MoohhRTk/Fy4uUAgCjHcKeRWxMFKPA
84tJVFWJEvPbJYxikWpTVfMWYZu4Vx44Maol8kFBjD6CfC/xrJU0Rx+8Am13g/VyADMgpoNPoTh0
yj+318V2IO6JNTpI87wOrHpZNJ4OekrEFT6T1C3dydyz/9FZRZ4eni25W/TCrhatHyM3lXmITdbr
sH6e+pSDaHVSoTKaiTr39/2vMHrRVJ3WrIDKsYYlZhadBIhkUIs937geuP7oKiXei0vPAm5Gj5Tu
KwhZZGAt8kZm9Vn7RSrGjADTi7IwMvBfHV/Z/J8UqhAzosWz0Q7MDDXQl1UKNi1ert6dDaMqmy3y
ni+RcbHC1bKa/8+YGW9si7hoTfY7AykAA18XccNTjG3yoMxv/55ZWT5bvHl0itMv+vnrr+V0IEoJ
h/Y2LRuirfsj4tcGHgDNExy0OhsHO/Gll9EBZn4B3eV1mg0TwNLhhrg3iA0LRhS60q3VcEOZp7Zh
U9EaT7rIPOkzaxN0Z7EZdw24LJBjmUAi2yx0wQXsus5bTqys6ZyBc4ZOAiy8NdvPPSa+aBOJJinU
rZgLymzFRm3+b2x/Zr2tBnr283EcQcbaQGdOSoWxu1dh6EFHr4P/qi0B3PMXAgULpGXDKWXZFS5S
dvOBahepcFoGo6PowwSzCtyLvvTxGp1iXJ0DFjjTta6ga/6wGnDVCU5i4pMByUpTm9ZOXnYEhW+D
ngCuI67wanAif5cd8f04amx0I3hao7wRIYfCJ+mLIbDEaYTFxnt8K0c0QYh1ded0npfX5Cs+Q6h9
NbSOIbCi2c6ey8DgnNCcGCFm7SCYLrvtsHNICBtD7leH7vHrzlphwRjHNjht2zpXQYv+OOczPxd+
9Oxn7DzcarJwQ1JF02P2OC7jPo1UWR8loC3cidA9wnsFyboaG3SXccS3Im2A9k2iDNbkKlPncMvk
nLIBwITv+KzZoHXqgxSzQ9HrtAqKjKYcCdL4CA/2SPHPO9Gs5+RSVZo1+4eC/raryP+LzZLEgCw6
kZ5sjuacl80rghwoIDsWYahTTWwLJpEBapzfQr0AQ5ilcNuTxLoniHIjqWPMWYXc2n4X6NnLr9+2
8glxcbT+v9R6hN+JzcJcQJVyzZW0pKZKCS0wxFDdXUjjPPVMSrAzhptIaq44/3X+Y+BF63VhElE1
VuCOjmrsWArhnTcmDQaO89JDk3aW2NQmqzuemmjZYTgdHATPcLjp7uDYQdMPnDMVjwzLTgdxpRqQ
qii0AFwpcqE1tqMg5HTnArOPnZYJ/Pplx2LoPjsY0VJXMEePcrEt36gXUOiRAEdw+PuI5eToNWs7
q7LM443xMrFIKflbyWxDDUv7znMzzxaxsyw4sKwzVIxCbH0/ukdZL+ZahHe+WBamYvO5tHthtQj4
e9BC/tHvBR8p+iSOd05j7C093em77jSke82r8tANaq0JHbIw2QQFeMAk1EXtQ844p3kKt1dA47m1
9A1od73LCuw3AT4FkJkoJz3uNXEsGyqZXehbnRkacqjhmqPmIWKftrH0j0H2tWsC04ijg9xuZOI5
LXAKFdaKCwIfZnQpmAJQgNsw2xNpp15Jv6f155CndSpBuUjZSR9liSKDdGBKs/DMtxLoezWVMqH8
c0DABZpV3TMag2RB2/xMrQAyYvXFaroF9JUzaKpTpSt2eoL2qsZ08oiMPkNHWjz2yxtTWiM2o8eI
dj3GJ3fGmD1fUgp8ekFH+miP1If5t79P3neincS0lxYhALtMeAQtOj2AQesw04fe+ceETmLL5fkw
AmNvCsu9bChHptqQMst/CYLRLI7/r23jJcgvtTnnaDRG9VxLvr6kF+75O54+c/aMwTHGuoZjpdtD
F0Lsdy3xSwCQgsA157uxZD/YyZkv2+HlmLF+zr5hgCZ+ZkJ6HspKizglZH1CPIpi4OyU4v2KSWvi
1Oh6HSZuWfvphYhCSBtVyeAbscHxS5DAsBHZv95KTaUkOyc1+eYV4jL0rr6x8T8DRV7O6nBObnQK
KdaU4omRSuKUjmOl1xD5OWIsB3l8L1dJqwPxXWL8b+vviKmfHMNiTL1yf2IJk3K8uPCxVSWZ/kZ8
tKp+woFmX3Wd9mTS40lt9u0r+xxlrDRwOy8Rs9tCCYvfiOUhUdiH9P49gWxjW52NwQsIyEIr5WHX
zlSQhV2odGNutCjjdhjPKOxvjB9lyFUC/Nuk+L8PgStg9gop3u7t1MFERgPUUw3RmINUkysxpN2c
EovEDP96RReyxEPidSayUJNfybou3g1kv7JmEV9KHMzn+RQ5XetOmMhOziX3Tbe/DYcqXiOpCPkE
v0ok+tbjZ37UBo5cOuRbSexhR+yzSW8sMOs8kVXWW3Zi6it2KUO5xQzJR23qc0t98eDpB0Bpnx+K
Ini9A154cNs7Blu+lA2OLh3meKPE+I5fjOUhKxNHNHr9quL0iCQFEpPfEQNvY3NzqaVXMeqZwjli
USIBWUPu7LgZgyrN8Z2iBKSzyQPXLhvce+yYxJ1FMt7Hhx+PCpwBbuo1UpNtNCgr+4m9y3MnjpOD
r41PmFkO7ZapY51IPiZIHonnefv3dKDcfQPFif/VHP/O9K78pwSPsiHeWlzrg1gATduAkfBbbo/Q
0G1gBROKbdkrVmn+SOyWg645YeK8xTFI36DHUIL8y6/XJubQJpbk8oBVfIyw754OBJQF3YT1M2md
zsCRoUZ2AK7yJsiie7J3JE9Knc9XSUr/vRFPzZ7Q8u/lR9MEfXC12w3CcWfms8JhDyFvrqTnnlKP
5LU29pfvxYs7slCiEdgu+Pffj1/BtACmscRRGBQ5SGGVhn7DHocHJYSbt8c4xCXv6NaLSpBHfChX
b1VBx+O0MpeaPOhXjGa7k33NWxB3iPzIouVmMvNTODyWLdUD+cFAtLEIwU5sAARl9j3IIjqVvJYB
OE7oqiepsKIeRkvOYlLQ1QDRpREiE+9ORkyCAv1V3IJNqeYrzDphuHHwtyzQxga7YJ819yq2CKBG
EgC6gZLrsgzkpg/II+ip4XOw6Q7URVNFvRx3MYj0c1GrE635Gm9aGlh3aepZLm2WlfewXQoMF2Ky
griRC9X+OSFxmbotoW0nNjKORSCWZkQvGhAe4KemLY38r+g7Xzd1UuUUfDBO+XE7kCnxUXnRfEPl
50NG83gb+IGHmPDz7XYI/4N/KvRT6c9aHwA/MIxlti5pWK7SrCqlAzcVPPbEChTZ1JwcC8+544pQ
Rsb2Tixq29x4xwfgSLNFU8uxVp6+2fOi+60NJgMXIrEc3qdpLHZD0WjNSkBnCCE8+N+tywH0HPIB
6oAg+R2lP94zIAOh2exxkreD/tpM2jhyR5mDUkFi7saNEEzX+VnePJo3jjg7E2QYNsBlalJxU9k5
hrubQQ57uh1R0R1aCQaubOOmPKBY/TUs8kNUS4gIEHJ3uX0uGhrK0/49/14zJq35iJ94cCCL2Puw
QRXKNMQ4ffw+e5vtH4Smdka/8RKsnIxYdoDLtZanvXjpS//U1bCHDZoiYqI4di0vtlTvBWaQRNyW
FLml68yyzZ+7vV009Fj2zIrxnlmEHy6J4oVD/zGvsQmAjjq0yKI93rvNmrEd6LK9vzo6bIoSdrpD
PuuZi50VzCEGlZb8owAJtl2F+rGLieYoCVW4NzCHntydYBsBXaNaVsEkPbs493YlqcN1sTtBPOdK
qd7sFg1fbar5n9eX9cQPWrfFFSlsv3Z99cbZyvOm1iknrLxeams/9MRDQ3fMXQA33ttMFPOvU8hX
uI46xOQji3RFyI2qqqGe08HSP+zhKJKbMYcuDN8W5rVGvJ8hx9JrgzUHhf1XhE1LXxVrAQl/KMfE
Anc0zESpA+Inyz6Bv3KEeUMxaSsklh15c1y9rtz8znXY9YFbOqm2/vNHeU/Yp2HHSWrVE1lw4uA2
ArdrFs4F/N+hETpYTqBhWjf8HUoxkKH1810uv/SlYWK6IdrAy6ZQuvQqAi4cfnw4PqbSIsKDddZa
qgDDkhlPt9IYMkFMnJ8EwwLPtd6JJcPSRGsma/uBMXQXTst2vksc7AUl2a2Op/0l+H9U2qxg5vUr
8KDu8jus6d3PvqpUAWUObVionUXaqMmdDkYmMUIuD/Y3ZoSYnf+iG7m5eEpaSAOA225iJ/bWoaTQ
aEQaM421TRR/hUE9MFei+2yWHczdW9pAI+ItqjeZ3ck7Bt9dR+fjSQpk+chMNr78jrmCheQ/iupV
hjGPNMrFt/FOGF2Wfw+tGAc2iI8l0KNy7UeiCMJoGi7MLOjwnwfQ6QSW7z2ehjjHstn+OcvERpNN
SdbbCBN1aDb+fHgQc9M21O6EtW33JuRXrf96a93p+CJ1SjOg38uY5iTCHKiDnfM9CF4gKlALeIDL
DdoOoIeH1limYZoxqnGaU/2mQZRIkyx3wDwVJ4lMrv9yOiBDxOEupw3JGwCqat5j8QOfF0sZ8Yef
YSfdqZmrnt4sfznwwylIBlusZwsdWONuyONxTNSEMH7lQRg29yNSjmJmL02m0YORhdJsPlvl/eNb
KhaSmP4AWwnN9J1SkdxSpxRCZfV8KsYoZIiYSmxLfzANnn3Vtlr3J6c2xrLwJcKq9DkuisTxHtOS
UafqE0PXPr81W2xizEAbiMASDB/9angds+P5nyjTo/lPg32/SqnKYlzHuDHgGdC/w4vcu8pX/p6A
gScnIVy1pzM9FgFMm3CWxQlsuAV947d+EyiFCnBlDr2Fvh5KV65+EV4m3fGN0TJfEWcDnRrGFk+I
+ml3DPJTiZoKdC8SW7yteFLnAEx0g1uYFB8l8mOPvLaFImT3XYdaIGCJXsBBjlGlwHiq970mqEjN
OJuVYMXIHaqcVqEkNOjNC1yB665hDLDtkxJmHVI39RYE68PWYUT9Q/H0oI63ub+wJfMBHmCJEfyh
oN4nIvW/B+jX6N7gccxzVq5/v/Opg9tc5pi5BdgMCjQIEVnEX9ylXxzmL2YVxvBcox6cSyKDNxu3
KucTwWvIuXn9oiS6W/l76BbJfBXC3vZvvi8ZoziPwNPwTRZtcvG2W/qC0Py2AWvxMR3W7MmHPzVd
pTNSKMi6P/Hs16piwEMLfQmle0rpt8h9q8qm2jiIwi63pZjfuZZv0cEFt2VIHlfVeTAFSFQGn8zS
E+NA7AHb3BXtZBKKLeJ9HiSyEd4QXNt+XrUJHqbLGp0HEsnd46t2onP9hmcCzq9+MYa1CP08ATFK
Na8NXhSy3alux3xCXo2HiFqQhf/Pgqz8CvlDSsRfVF28rGrqBhCrP75b5k9GEnSHVi2CMAa8bkVH
oCyz+89Ws1uWway/nrgWS5aN2loExHZ4d6H5hl1mHCiB7Ynzaku4SujBh9mqckf9RLcfX+lt/NVK
P8CN8xh5oM32Fl8GbqhzzItm3w1IcQhQXdVaL1bYqtAIqHMH/m+1L+jRp8Qr4oGwitN0FAT7USqe
3vtRroCJRqEwz11b5zUcLlZnx8cWmdGtj/xmg0Q0erH8p1UIZPQo1S6Vzb95iK9YZ6q6UlHxSkrl
q795vybnrsRIpmyuDy/pQZjHVzNWlf6FfrX2Vh1zzDLY174rsvaLzVmBYIqR0TAMzmXQ2VwxQJyu
I+PggnX0cxe/CGssTdbjQxwFmyWREDocGvht/I36oEe+KHczgVzpax6YCGXT4xOUNuucBj/CV5dG
DcmZgQKDfF+pyziHu40jHaqLk9t708EPhSOH0SvvS07Sv8A2DTWXMVzZc0yqlJ5gIFm0cWSxiNkq
xDSv4irOqNtGVDc0+W3mv5QivnFS+cdu/oEBGfBmKVuDSF57yOYvlajNJvtoRaas+2zMVisEYE/O
9vUpwDYZ6oUG6SpzOgz/35olZz9ALjh6nSDJg4lsKZcpPskI9yeDTITVfxlwAf4l01ALGupsLRtK
DZ4+jAsfAs2WcX/lEhjBol5KOPMl0HocFvG0BaBhg80jZq5H0v7rTv4o7lXt34z15e8Kv3Kve4N5
9Hdg7k2TgnmrMd5YVk6twAaeDZRm0auPdHiaF0ZYzBs3Mmu0VkJxGpNcpsQyMkhS+duDf290KSTO
9NhiZ9T235/INqm/BGrTQPJ8D2LixOymbPUya8NObYrgujTBHdhH0gxXH66b6oWlJX6GUQIknbyv
vFPl1pdbXLRqdI7bJ8DmHlp54TUZTPN5qNjGSAjRkwuTyBTvTQxAIB3+npTW/kv+1XEvZlx/j/VK
NHb5Ra1ZG38d1PCoe3R1jBmB7FnLwGS8vb1Hoim9SWp0TSvRnHkrKod1smuCWLgmZjAB3w8lmkYI
R8gpaLkwRCYoKsifV4sCp7qV6J8+es1G0DR7T0VEM5+IwMKGnRA2XmxOvplVesetKCXwnV8tvkSQ
vtRma9mUisa/YNjZ2ZfrQY31KxcmYi38EWg4UBZOKu22iafy0vSjIMaBoJ/jVI/5csq0c3/aRzrF
GlNWzPtNrZQYFT1OWKSHyRLWhx+XqsOwmMI2+LhTmi1Sq7lpmZfW2KD4eblQxBf5Z8uQkFbYdStK
+aD8GX00RicCsnHLWgX21stkC0yGTcyWmu2907lBrJjY64V1hNCAw8oi5nQn1Z48EC/+TXbF2NVW
lGSlduAEE+66BiiXVf1kjALoVA0hcGCbKzBPh51TAkz5zFLZV0t1SnQi7DP1zqkPegNVOLu0if2R
t7BXkAYrCsMr8hax17NH3+CsqXEaVv76iv9mY/DVJvz94xPNpORc1QY+g8N7GMGa8wXHFd6OdcQz
r3sN23DaizXMQy4XECj9cq9OAPydhih293z1+efCBE/47usdpaRDev/OwjcuHMbrVfR7TqVGVPRN
MYwG9H0FU7CZB/OP+VhcwsoEUlWeUJRAyiQo/8IOLpEv3u1UhedkuHvkBPA3a6p+IJmhPi9JV0qH
HTQsdYfSrP9+WIW6a5/I0XrfS7dmIoVSQP2t6fjLfFJtunh52vm4SSCj/W9C1H9hkkmy2D1EIoGj
hvmr6T43jP8cReRg5MvdunoSwBuGfPOS1Nrmwj7aFY+5wIekTiXZnOzOIdmuUhSLY2hrEuX+mjP9
qz19iQdXD46NIkHogHfRzWtCCoMCjAWtEZ85Cl6riKMZEgAlofDHcSiwT9Wvmcb2BzCpJn5i2Ush
qvTBTQaBjx1VUra+DJuDVT9K2rOwPpdmmRELVq6IOntpzUPptj8CDcnxrnYnqQyDllBOZUuWNiLD
zqxT05G+sY0uLhK0AxsHagi1dOneIaJGqMbVu0xYjdFFDgyRshv3p6jIOkVPBayUMK434HskdhRD
qv2xXg8qdDMipTYByGagJ9yyFbzIvHE5vOPRlS0BkK+cgHqrKHnxdv2HRmAZ7bsP+hV5cwSEj2dl
+Le4L3EqOc7zPt+VjUeXLDF/PRh1IshbrpxUGoxK8Vb/uueTe4ppLnOMiym5WumFqgBxu6+mWwDY
uYkevq+wJAX0dm9ZDKBU27uo5My+ca/WRwyX+2kgvpJZa7/Zprp2glwDPSGUcYHnspzGYlhRSa/v
/5FOJTwA4tCo2ZyUHcXWQPvHhtefxvi3gsylll9sFitaqfjCkGMIJoLc/JS5i7TWjJHZ4qqYytFv
6W1vmPVnqGsHvf6+jFFwz368r2t7pnibj1FHU1aA4m+uOnZEu0iaoWNgEYUBjuXGH4GKHNJlj2YM
883avDr3y/q9eCJD158ou93xtDFOkJQjfjGneQOYd6YCZFFMMLviZpc1BNFueZGbMGYRl4MjNcCh
qsdGsIfP4FYY+OrFTXCkpUl16etALwMIMyhpjABuzfezzaNzsaq3FOECniWpGG/oK1pUd0d8nXlY
ECpvgkF12BbGzBORZezCoU31xHf5g/+VFNPcT3JmURItTPZeIIh1gIAC0N14GGypt7h6CakgmDT5
nF/OQr56QVeadjxlMsJhtmlf1DjPRPxGUwki4yMcaDoJZNZvG/s4W0I3bJYQOR2vH/yjY+ppRTch
d3QEEiArx2FtOJ/ekcRV/L+qcI7uY/3wyAo2BxbwKiy/IMxIIZj93jw+nvAXctWCuT0l+RXciKQn
GjKC525Mbe4mzjdpLOotTMqAwHQ9VNVmI+iZfVxwRv/zb7cRYF6wS+Zy3s92uWh8DauXfcYFYJ3P
7e29CW35cpC/WRbEt1t+0MYlvWuiMgUxGEYnTxivNRIncmwXyvIwZgluCTeJeU2TQcNnUayu1/Eh
kTzqRPSL/pcR7xx1XtHvrsKegpGAaQZ7mADcTfgzrHAQCFBP4sOkddoVYR0IAA36E8kWAm/PUkwM
0XlO5rImWZX/1HCsIA4iz9/S9dWTxTMs8drwxDpvPgJyUpLw3MsSh9a0nhydsR0uoUkeIAnf9wcP
9G5SxaQfyBzEyv1jBHe7Vp5jQ4b1fKna2Yei74woFKI8xvX4GCQTsZ/0Om7N9JxiQRkhzndPI6OV
xshi23ah7LAUcYJtlAfeOo/l0P8TNvXxKNCMApUxLt0peFL5V4lJdofeVB3lksBwqHRi8s7hNwqx
OzfIJG0SXZ0D1eKZyEIbXB+CP/Q3tOjkKFRUbnh6kwZ1ipNZSTuxpslHMQcMZl/zH1YqFZunDp5R
78D4g3PfROo1ezd+QoPIFcXZHonHU6HvfYjyXyCv6/BixIVmaLdbhlVpmtMJnLecRbFyxt9vN6F0
kwLxw9D+8OAc9Vsd9a0uz4zkJzjbpuL0VEjxeH4yrykX+HOaH4WBICXQDveNQ5Fp4x2uy8pG7Z+n
9CvG1HBtepet74rmepOdQh1dRFK2tg3DRJ4IiZdoZWi7fiKtRpiHPT83pl2J2NBvAPrYyi45SYYe
z2+mCDa6dSzuLVVF2RSAT3jpd22yMJd3Gr7bnAepWpmB5+HaQGKjM/1I/HJjWOMMmLQU4N2UCUG9
8xFijLNFysLBL3ZzfXMqUXl0V8tt0j1AxVw1uuj2OSvLSVzMILy1GdtB7lG8NNmsvsA7+p1DDE+j
QyZGK3TksDUmxradNzbtfNjWtvs+wft8dCXiWQIeaYmR7kPzwi/3J7Rg7Fiwnv1WjBneE8b/dhu8
oc/zDFn4CIDGvqDdLyGAnHprhrYrSurX9Y+O3lO0DSZ/eDC5pWAJNYMuUB7A96mEFzZLoQqbMMUj
oW965Huk/xUq5HOpfjuObVHmuypyG+/Ce+zejqeaZPdIyFhx6YQkvyRKPF9cZeJamfnC96K5xwTG
FcBK2kzsHlNP7fMnzOeISDbRbUgDf7SUI6HfsRqAX7xITs2MBriQP0Jb8/Wu1lhgPceWYtnzAQqL
l03UcWofn9NOIDqKm4SfnwS/XJ0uvOraET0Dl67B5GEigJfad5lUvdpEZTwpq2VbC6vijnI5CTmS
9rCY6krOx0DtV6T9f088I7gsqQuA+92a/We8GEoybLGRyeGL8mr3xNdJQbX6H2tR80VyCQDy/iOU
BAseoYVBEsYNSe8R/fbDbhusB9KjGa0FH/WLM/pU2rahimSM12S+ZkEcQq8ykfMaKJZGovh34AVO
mWVClmO2u0A6cumdXrO9IZHjnxkr29JUdCrMj7ektsRWDeOmWM+PqQHcd6u4Gmk1nVAEmaHWfffn
29Lv+DxZMPY8KQPhZH/daLioVa+XXfLioKUObTbcIAd77RlQJgEeEB/nAZzP0Wmibj+roMgLazkh
ZegRK3HRK0s3QkIex8Xt9gtvgS9DtrCi/EiZX8DlygviYNou0I613XjLGntDN1j6d6UDOkvBPRYU
Voo4hA6lisqbYlOuhzdEP/Tz+a2odHlyfiKpGwH8OeEIalnHg/voFInVxZeoul5E90YCGziXFnXy
W7Lv961vCSqR8whaUws5WmC1SWRU1HbdYOu4lBRGWaOBSd3vPnxBpyiNkr1teN9b7j5p4UTdabun
EOPppi4yhRLwE7VVECRv0pk/XPOwfCy7v8oNxkfalJq94jSoubv8kkUp71UtTmthCxTHlpN0VcJK
4QDYWvoSOkegPg13yrZRzP6fTC6ubQnOOD4LwgkS2Nxhg6L/d/vUbaeepYo1p4XZ6q8XQ265mgWW
bhVsZy0mc0ACL4+JaPeDZlNVBEXCZTn1BiMJSuz1K/Yd9I5XLdRc8nK+wJC6pp30kKaRvRBsFFem
1oNgMg9UZ4GqA2HRJSoTnLsLxJNrtGaXKZrU3v5hkcx4av7vi/dCTArHYsBBr7vz2fqPY9U5sf04
pVdh0AdxESv8PCQ6dghRoOuT+1AD/9mZGHDzk8Mi3Msysa4sFe+NLI9T7/tSAhCQPAuQF5yf4Rgx
Ci+VV4M5LZXBOitLrOzy6zwA6UbuJjGJSqfnfItm3JKFNipKLGwy1bvoZqPdnFZJuuSUj9bm9/oY
rS1zpCsYvMUKJDiSNR4sQIdbt8DEsv86EvGPq8kXgKrhJ9LYebwTwa5D7Yg0WVZdqP2gMSkjV7Zm
3cWz2w8jZUBjodYSgvaymsT0LvWAfd+jGT+th7gRb7TwhRCiilPlJ3mqtHWO+m2VejBqYYQ0K60b
UK4y/F8aFWFCXIAq6/5FZt66tnB18HR1Cf8QCYUvj0O2pwEFCpekb11mE+HaqFiGcs1nElZa24zp
b5stm9NpfAcKiOJXoN23HcNpFG5pKwx/O6brweTOh9Uvv1z8j3jJoBtn0T/txMsgPSkXIWvKKmkY
INL/vyILleRIGJwtc0R5EZQhqP0wSTwpv68ZDmVNnfCTE9O+9m87Ef19tu+8xeCppETobPQoOcLK
xBYx1lSpl4dNepv7Zb0pFkWx6YP0ayDmiv4nXvYhoK/rnWBqjvTtX1dYhZV30VBOeV1MlRCHjDfU
Jul29boowY0eGN2TgTRDlu2AId05SMmbN16/Sm3yTHNn2u8bSAdchcaA7p5hIVTrlO22IBZ5MFJF
mVs+zoAK/R9rgxq+/VLyqQGvw/chKsfKSfjx2m3y5RxZEUzPRniGnCxTXm+4xEJ2cuA3K2rmmOrQ
h3cL3EAdX2L7013AxBPNkDYR1H8NPZwSGbWpoWZ4ZDN83WmEBEgqBWqsDOACk1IN+Nu3/8fkEupU
3VX6mrTMVJujan8QSUQ6ziXMI2difbGz38g15BiuY4hzTm1bd25Thy4RldWjJ4GyDZa1TO4CTp7o
Qv2jfabJ3G3YyuehY3EFfd7e96kCu9D9ATBZqNaWsOV3RatPQBVwN4LEPCBiVpK1O/Bds2cDMsQl
O6vZMv3sHebLMGDla/VRqDang9draFAL+exlQ2M6oAogCysL/cbsRRNlDPwLstoCJBIu2gFXVPxN
Ha7ZCR3veS9cdiWs/7UwlId+05a7MIlx5yBjhUJOjpX3yaJMfqQPmOVvrswWH3trE6HWIZecLCoq
/ixLbTmB6M1AR58Gnz0eKBoJpaoE2yyR/ZsFMB4zFN47IzjY1PJOzpKibP3gk+tJCiou3akyHhZ7
/yvDG17bMxLbeIYR28AkaMGW1sP96vGxPhz268plGWj+PjwqTvrs+G19Horn6AatnZEtb8E7Yg1X
RPeOplJuO0d2988JoZseDYSzpBDIOL1ACdM5N6t24QiMTNEUdyn1xU4iyZzsTz4BT1SvEQbcWeHz
koWxSukMLKTRnHviC2t6akb05JDYc7dt8BLNmnCrr8YcyiFvxppCmO7jy8hRhCGBeKPoBYuM1w7q
7ENjO9E7lZsVUfOYGK7unRD7dQT2XuatIR4b2IKuYuPEn85aGxkNVskppqCGmEwH27cN5Z/mH59c
BE4xcYy8NqKhVkaGAej2W7LZu41J3IbT+bxzK95YUCmlB4UUyupp5sRySFOLZvzvy6CkzQuwcynt
/NgnQYZ61+PtnHP5cTHOzW8lz/p77LeJiR78FGAf7/2eOUTGEbaRjeCIaXQki14CkB8KLtFWNX8q
NJii8ujygM7TmJgB1oKPL/EYAKajGSn1S1I4KOUDBaey6AZfgb+TpSswlDm1j2fyPegWU2fcbVtI
0G3RvBh4xi7UX885fQl5Av9FLiiBsM7HRjcmB8HkGkJd9qHHQu3JdvCnz5d9gBC62HxwolkhqLsu
OFWPsiElEzqGNdRxUNMzLlTNxD48CVuE7llGhxSqEEj32e7OO3DXlWSgYg9m2JQZxERdDYSxsqkQ
KydqsIFO2cjOgnv2SJgpycDp0I8kEJ+iwHj7f4U733Ihv5YsP39a6V7ghn5bzE3oo7hSFuu9FsdV
vVOfSPS6LoSpNw80L/tKUWBzIVEm192rK1f7agpn6XgDL8dBMNgLmA+sPPD/w4Jo/DTTB1ZoDnq+
9Nfj86vxnl7KA4cxpRfe9MujbSkc9U49clwDTNpenHdTm+aqVpD9C1dzIPcJWo3EYb98iH3wSiwY
CMxQEN/w7jmfa2dTODVtJ5m8FHXc8aNyIBtt8TABZUblh6KpUUDbp0q4mkCjQlY4QeUScm1Gv+w7
SaNh2AAYc9a5GbnsnfNtKvaA7+7yaMLWs/rGiOAJpj02NzR1L3S4dDYREu7J1TjFwyAFEGs/oLxI
7KiZoLIsL5hvI4hlhzONuOTvcek0wHepLcJd1JXq0j0c3Sp3A06p0xNFl4ccjZbwAdZDQl9WKkHT
ua7ePXxxfMpZVBheKl99CojM7uT473T2/g++iBkCCJcqPWER4vCm47yB247XgH/RpqFWMDS+DoO2
1vq7iK8Pga1diW9jispwSHei6Fh+wI+TpcPtnLnUlwAmAfjjETn2SMA8ieC1zsxxa9xPxRcziIG5
70ErksFvE0KbnNIeC3gliapu8Z3NJk0ZgSD/PVbjN5RUxAgMrvSHq2EOvjk+pAfwkx+pX3a52Yi0
vyDRKr3gDH8prdspvZ1YkrMLBrfoOlcyLep8VZaE95hacqyX9j1IAERRLdKejBPpl/SyLF88+YCA
fZe6dpz9IYvqa7gv73v0xyu4bHWMZUFvCNwCk5uzsPVfa+RKcVnpKZmZAWJEpild+GCxFQws/4Ct
NJVdQeekutCGfjJkBJbaHlaa497RaMoJsKqbY5Ux75uORLIfQH4imqg+PDDJrjkcX2v1Usk0KxLY
1WdDvtozL77eG27G2eYMZE2+H0BSguGelZj0qzN/W6f5qveQV/NmoC9Yx1ERmRjCPlqMk8okrFAG
k8dMQP72BFg/0LVXIA8WCaIVdvOjScRIDiJxhURtO/MpOElpXt604TFR5tIyV9yLBC37L7R1ZsUf
eVqybe9VeqLg8zfeRHuF0mQSmo8f12ZaN9/TTcIk4Imz+rWlWJPkNMgeu84Ay5jW56wcMjHpsjZz
evnK/fWYsEH4O9QUHbu8lgM7cEH+UaHolrBCDF7pnhxSNdePe/dRuJRlM/o2iusLfBYiBDL8aZTs
fwTzFvOrA41P/CQlkUZLlU4pgFVY8+a1RKkh8WTYnQ5eAAFoSmO6IRQ3x4OR45GB0kPEegcxJdU5
iYcYHnNCkgptd2fasQY1/jiVHQA1L4kZiNGgd0z5y+g5kVLH8MDrOG6T9yOeHM3AYPZqEYZK3mlI
Gc0Jw0Oj28WELy4tlkMKMtSXc7t+5pUp2nEih6jm9YdhM5M3ePCiMfUZBXY1VAay7BJs8R3EGpsO
hx0VcWHUNFDjmq9GkYNaMKjp52+V0uSpLRMG99OwrRfgj+tbf4qr/yAFE2mdJQcv6yr5C3/xGQ/7
+pAasFOV3gV4C62AHcb/k172wTwcMlmyIr2+QdTWgcmSk+wEV9sC1fnMk5FHj9o5VgJMeQApaFKF
xawZCo1dzVRjscZKAffyNcTyZUePhRCtJ6D0zD+rCM0uRar9xcHSX9NyVNCkzeYZWemUn6zEdX2L
7jdz5jwL3G13jhArngOI38chQT2hcRxR8FUD/qpjknDPSgLxfmt/UbTfNrxgGHsopz+28UeJjZyJ
l0QSzq7vWH5lOibBXP+3MlyDESQ6LUUtbpCoyfzJ40QnCzdxAbUY/8B5ydhtv3Tmxn1fUVNlNiZ3
fjJ+GJb0ZT5UHoQktVLUiwIGtnTVobZuavAHB8cEmYQyUaUKdC/lgKL3k05NLRhemkaOx35D+Zcj
sE+kzZpYim7AuYWbGCFgwU/MrNzU1mHc/6/6NfsgVFLv9K6Rt+aDFfpHWnHH5W4BAx98eoTCxPzr
EsjX9i/6L3Ef/GG6pcAnItVBlWaeXMbCrux2A/HATVgIgbG6mmlsg6Cxh7YpyylCALwAAiPrylBv
GCn5TRBMRZL7B8cBHnKgHkIAPR+5JNe+kW/f3cgSoVnpmZRDY3DdKZd/ek2UmZ1NnLeWYWkNwJWv
5XfIRv3+Sxs3bQGoCGZ+ss9fu4kKVuFN9SSe8SSCBQPKhZcWRTPlQpx+ymZJJYRgb3qLJIxqF3Fk
2RI0Od7Gy3et1b/ke10hDvY6Z916YDRm2LXuFQSQRnpe6wdCg0WREjNAXAvB0E3Wo+IFeK9fuwZ0
1/doVPjaOL35DVy6foS1MOoOi3do7tPEMoay3O6y29k53FQcOQxRWKX8BlGLxRSgAe4Grkt6O4NB
cXWl0zWKvnzV7RXxXYdXfsieOFIYHBse7kSksvdztklKdBV8DWF59aXtg0BEQZ712Jni0vac30Q8
Gx0WaBTWK3TLu2ybtTTfukDdXzufN7xIu7eOIEeFGU0BG/q9TrkyX5hG7X2ezTyNY4ksHZUHOW7u
fsahVu7xTJnXFZapzpyB3etwUYZuAA3/G0yY/cWOZzI2bZqKbrUxkbt2M/pS03ABPkwOFpoEzeu1
Z4POv/W4H+iHPSShorNxgbYX2QjMm2dLNEo1HQDfY5j+6EldYXwwtbVgy52jBCKlh0VaQ4EVOPDR
oTKOZNcK+TyiPgJ0OpYkfqolhR6Rdy09QVT8aMs68LqtRRJftnd8xCqSiQ7zL4TLQzVrC1F5I9BX
RHSRDL/YI64jsnGYclwTt0dZlVp6AAXFD9D6SB1IYqfuuhDcMM2SnUjdxBjT2hOKoR4KngZK535Z
kXRRk6wnFsEfCnbEZtfiHdi4llVKE/XhOBTP31z5wRi375bqIQZee8GIrYbG+qR0xMkbdVma11jp
tnXgsuMGlo1oGNau+8+nYVwwf4k8RR6fUc1u+bijdVUc7xkeXOp5JYWrEytmR9B5a4fCQKxdFAAO
GiGoLzgGgOIR3vJTx3c4I4UuJMqCxC6DgfV6gE8W4QKVITzmmbz8nkpd3MdRvSdZXjixHiVyq86e
4MbLAeAFgj1FNcvt3tdF5ugOXkCsxCW0vakWerGCv2ymFCXrKYoF6MHF91K23MWEjZBRmfvpKLkI
XgpwdwL9/2e9A0gEP/gDkkSpmFY0+cQUvo1dZXW6AmA3md8stCwSHPrtDqSuOJdWXUSRcZWi9unw
GQI6USRtB9mNBDfulcobMW6JLteYcSf4S+j7ve6uCcOfy6RDt20tAiU0iwtZpAQL6orJTNohv9UW
OQNiO5S4OFy+MfduQIfd521hjnh/MathoH09ZVLTrBvTyVbLRh4lvC7taoF5T3Yn5dpCEfABRr1d
uYlupPHgtJcCaThFApQ6p7W6bBBdHd+d055hHCpjLuK58V04lpK3swdCz9bl7p4Sz79O6HxdLGJ/
MiT/9zSKGWjkE6pIvd1RUo1YEtmgepfs811x3BRM3D9ejzKfVfBCGLUr0KQdryxOSP5StRd8LEGn
DIzLBABq4QymOT9lH55guBef909K/v2FgBL4R1zO96r/PE+DuO6s5EAQd0zIYXOPF+/hTntpwdwZ
MOX749X29xJJgUXRfWJez8KdylmmKaQuSOytyyQ+vg/lqAHAfjlyXmHSxGOYmJLaXKxZSA/OeNHe
T6raWuEshVS7dkr/LZE8BQsYeHy8vbnjBpRzM4+i3omL6uGmLGh9++F//ClKTOJW1aRipcL6bSeK
UIfABZcYdt7oRT8vVnr3ZdMLK3EQzpuIyVbgyOBDW2mQR3OZ5yppdW8ftSa1yZKFenj8kqqkNwgC
GQi2Y8Y4+TM33PEyFQW0gyC0KXWEl86ZQd7bez0AEdtxTq+Q60Lyn0xs/1WkEggqENCgGs44uG5B
9aOL1dslsVAwYl9CF9YjQl48rhX/G/ag1OM18PlT97AeAG+I9Hv3+EH3myHQ3TLxYa9rw9DWmwof
yxSwiS5cmXXvHtxxfrYgKRX4kDhMaPymjAR5GUFZmV0RHmp9BMG4Zn+lb78a5ENQ1z3lWJ+69+fR
Elbctu4oS9olVACyEq+L/ib15QrgBU64q7PuBVwAxR99rt5w/3MXdxUxiYyewvJ1SGjFqIMJnSsw
fcZLdFfvPTIdB/T9x9jdnQlfFZAwpnkBWbYR10Rb6SyLK8hZ/mSm5pn0z8NftCI/x9KbJHXcGqGh
AVSWi34efQnDRER0uwJtu5ImmVNb77If1ZFXNLZitz41TjwcV1f33UtJB2ssZB7sP71dbIGUpGVc
O3/O4p3rq4HK9tOfasc+/1ewskAK0y3ZaUBN10tESN2Tbe8HDx9+2BPXDQvTjSTuIm2zriVRjLWm
EYzlQxsekPdsYb0pTO4T0qnviYCevz95Am5p0Wfmx9rMVB6GSDluYR+Qx0aF1OStBaYt2T0GVtQU
JR+rchhtGtz6DgXGbTFMUp9lf09vEP+kiD4logwClI4PaFnzFAiOIquEHYMWz55FJDcRvvJTGvTw
9IFSGXMTSYMr4wY5EFSY0KWojSXhI5JeshHpLthQVP9DQP2m7Du40fLYIEuM+Hn1+TyGmGy3Alwh
3uGpAp+OOFlZIwI4kRBgQPTIXc/LDU6b+TnxSvpFjjLZ3EbV0j/z8BH94PYzAkwQXi1z9Ydb/Dwp
vSiXpxxZocwkwJsbZMPOATwm5whgUNnKcNvTjyZ4MZ65/rfFvlW8wdHz1+FdbMUuTJm4lwadwABI
vN/LHDnW4VQ6hncUIny7UxU6MP4Aw0OpOS6nMAt8CBSnKpA+9u2nUHKwuClNJyN5AltuEYT7dfUv
xPFjwb8qylcKPHY/glBguZ6ahZy+kw2ccSeli/J0W3oKGPBXyxETQZAzoD6rMa+1HVavtfZo+ckM
/rCxEqgo6M14Hnp0fnFTClgt68L2RIMMwD7NC+VR9N9E2vMXIwLhMQ5UN9JQMM07TnPGz/QWB66h
n8w3WEDYQwrlRP4EwC5C0Ru2SWwz5ko7ZK9YISmSRlhSwUdqi99YXDBdfpOFZVGJUrvd6jz12ndk
awilK0CvUpXzG9JtQgD3rIpzGf1xyX2pWcd7d6E6of/B8u8WuFwuoz3qz7rNR9QhLBC1A5rqcAxD
Sa5oVhbEQsII9uf2rPNEXJvMy2SpREG1J4aTAacNmB9cPqhWkXCCUlz5g14HdQ+1TJ9I4+geJuQv
ZkhP60poy54FZQ1q1WEO+hpCj+3pYnfvrl0jfHXZ4BiWJSTZYDDW5blyvedPvI3rW3QjuslQJdcJ
yJeIs+MOs8zwZHG4Qb+/wQ6v5hByYGz7xCIFTRHK3I6bPWXAgjqHuznw3g4RKViXhdm9DqqryP0I
FPiVNnv5AeIRKUZDC6fbd0Ks0y/wjRZpPA3OQd7sA/eBRRBQrwSO1zsL0WA/HGyDr6+EeugB+lXY
A5a7v9GVdl2kSUI0Znqj8lyjaw9kb/zweDZ9SvJvbdyWTLnyPANHz/ydBi8A30AJHSWA3T5OLeaM
vCL8PVQGJ2BZ6QmNeqgKhJ7dmJToX4HIBPdCN8qBCotRvpNoIwjpysVDHvF11K1MvazUuSaTFQR7
+Ho9G3T9049y5LT96rfrFcfek/mmuf5n2niD9Awgia4fVjFkdZYgC1Nq8nr163e3i5cIqgsoGOnv
ixmXC0MtLxFvq0hzq+LPfuvJXe2PDmAuYvb6IdDXzHOWctjE8RvF5HR9B+c6+mdqTVDs4mYnI7Gz
Gr+JoniHvHF+5K4pfP1gL+AwUigBYlc6TiieXTj3AXXh/gDmaPTsF7yX2pGIi/siiVUc8wPr1Un8
0OZqlZ2TQdekQ4c1q6gc7obLD1NOi5ZM1Yi9PwaXROrg5XmWkh4O3M6jm+qzDJkEuReH6ZHlAnx2
6gddJaQG4xsPK6Unh5g63tSj4/FAhjDXX91+l0EcNu+OyXswFZF53qX1lCjs1iFeHKQ0TW23oCir
Xl9Me3Jwaw2dRk8xuX9ehWaOxLDPOY2lSX3TBR12b6mkyhK9hdt3IIFotpBbZzMqJd05smKOGPmw
cMxEndkLKSJ9PJc/2n1KMjxqFAFrnB+UENRpl4xZk6lLGTOocpEGMRMNK730f6a/7S3B5nYUPwUZ
Pj8zPPwvBIkxnzQQGx/5Cqi1yvD+lAr3W6BSTo6m3mH25q+m/pFu2uv4zSx16l0yT6EyxHlaF/Pm
wgIJqvZSKGLg+XVKHr+jFCG6JXwCyBDSciCekHyi4lv32KJDoU33B0l6tT8Vc2dsSuvfRzGJurqE
2YjRped/LXc8Y2t4ubYtwJF2zhbJmKAv4LyndRUUsYpdmKqg6rXc2ZMhFs11s6CurG0zv2V0E3ZE
yP8BzxzjtWM/WySlrFYE7gBamRaICve+jIpb3sNQxB4O94Dt+u/fhx7vm5AYBO2B/otqY6mH5Fi3
3XbSLSm5kcv9a+ytYBiHbrMO+clkE7D0QfZdF1tUpYX/2NFz1Q/ka1gE4vi7cVjoCfNm2ZFJtpxw
4aos8sbgHxX98z4eAT8Y+w42R1kUXyGhtvryq1QQ4tKvr7L9XtMKoSN/exaSo4X6rW11hNm4e/q2
WxJtQrxJHPdaKzRihj8RbXgjm2mICTSHwuWXFTeNcI142INBcjU9wtzw9PCVL9LHXFp3dRb+DRU+
kiODWzzzQcsK18AtTVNoj9zopWjxesy9xSWv2cfG2dZkKSz62Usm7YS121Q24W7oez27AeAkSxK2
tFzljMzBRusDyhQ8gXmDNmH7IPVgVeSyUTILbGHUxjxUxb+v7W+Zkw2FNz08g7X+MCwaiWu3y//L
vQYawCEixqhH+hYB3zGPimdGzzV95sEm5PVji0AA0qg3/Q+kAxnh9Mk1h5r/PCo9rg7CMhA2Seio
+dDHVMhfVuRkuFaCLaoCO9+3tHcYCUnexTJmnILnaM7JhsEKcowaCa9jvKJ6UBS8pxM0wCkapWMP
qUsUQqbkyX2KQZapggATsW9J5/LNvI1Ro0LZymePIwK6B+AmKK8P7lp9CuKdM5dLbAMjE7Ot9eFk
HnYI5MlhP/AaSDU2EURZr++cpwUaeLaMvEWAAToeSrClL0BzidkEZ0O4546gMz3+NqSTDq0s+6hG
p4wgfPy+OSX7Pot+zkn6fL+HeXFn+Of8nToRsHyklxYHflzNVQ2NTl7YNJnQOmV14MYF8keJzOZ9
ud3C5b6xbUXP0SwKUODDfyrzysk0rmF7LvnoaRoagjKSznODhiH7pyzIrXKNMOPxUeuHz0iJc6Sc
G1NuBUYV0/zHEDRAetEnHGd9m+0XZk900KnS5mF/h4609YCcAVcgqW0HlSzIcedoxw2263eRw1Pb
/PMwyGaF+js5nMq8b0t/39pA3HMgFXf+QPcR7CdbQd4q5B4/UMPH4LHQeXPfGj5QmXyMOBgVkKG5
3iBc2l6iGaUfD0UcFdbxeswwdfjEDha6i8wdbUOjs7Wj70dE0NTtgtJEtfRw0ovC+mymsX/ulKoH
podbRX1qoOmabyvKd07HQKUUQh/SjyL0ggTI2/EqtW0vp60Fqn1L+d1tpitKwHAratRdwJP/qee4
kd4/4Af+n9D3yRda/sYHGfEyz4KzoyAk+F8oOolzbFqcvFgapSgxhUhU9MJ6zd90aZwooYyDJnzH
d9LhM1NGyQ7cuxjAMZgfLQMnOCS+NWNfWdQ2w/sEFlmGb7iEwAgXd/2cKEJIOSk8XYmSQBTlOhmG
HwHNiMxFerjELtSouWP+yILYEkkvFiQ/uqFz8ecYIH/bEF8Wvj54qLQ3CEOEAFM6ztnupRSBx+lz
medBkzSZID2JPQoMtq61EmyfuWNhJdfSRfQShNZXluJiOTeLTplnTRV/Em7vzEUEvr1qFiEGUJj+
iBBsFkiyPop295UcOCttXAuURo5BZMtP81wlVVf5BQJSkrvNygGxUDhKX46nK2SmdxYCWHBd4/AL
s89dB+tlvCvZy/CtxRSM4w4W2f4JZ9DfB9VCMmZ/DOlBoMFSyYO0rynLT+sbIV54rslwCu4nSxhl
M7fhg0baB2vCq4jNs0Nts9qR9hdUp1Y6I8JT5J6GK5STBRmK+MC5PIYFSwRQGaV31kOOOp1plJRS
+I1JX+wWNLtNCQYKBPbtNN5T8u3EAHMYinIOvVhFpwNdFyrDXhTkXwiIhdf79l6a+NSJOoiflAKi
PGGfIldPbCVwM9ZbtVHwrgok6EF2HUq3XeX35dIfg8zze3f7vRPJUYwGHuJW4gGOavfPPom+6ZKa
bXrOYBgJHd8RAV0N8VhRh2gF0gH8GWgMbYlZkHIiDWelNdOORlaKncmSEUnBvy4KODIRi2H7RWdR
xvIlQsum9cTScVdVxrchq71Ns7ij5ILu6cLF7ELacMNPcJIue1+gpbJQ2s21PTlkL3+jubJK/Db1
kMoW3gHYOngpzzKmm+QzTJUz1r+rRiXVPGJjCu0uMAcTGOjGnVrr3XwHu/oo+8H6mUv+58/QUkiV
PeeYSnlz4/H8nKOg5T58oK8lovibak+50i5f40vmicYkcL1x5sEGIF7MZc4+33WH1Zx38/IwVcc5
MVOwAax39bxUfnfuCjTvK7210PWDBrizB1kcglpnpmfNsuU7iipK15EaELAFk1m7VjyT6h1sPeVr
JmfMDfGCUqk+/T+gxPaBrvuUqW3GKFbWEQ3csOkqLNcZtuZTmO0mnKlGPprAkpDqS6lRaqexuw7+
3skDqNoo+xmpjeu18BX6x0Ke6u9uPrcib+rz4IhlL5icfj71DtcvPtfqHyi5ZginwfsxJ1+yB9yc
6DxNxIxgNH8RWAM9/JMpBxPu+T6QhDZBsyLE21lV9XiQxqua012dvxvSZCKJWT5kDBDgq61QjQQl
gF6yWLNYgGgwsdbFJDU9AxS+kJwajEkm4iqf5639MxVz+PXYru8gtnoNn1oEiNqwgNMZ738x6U0O
AkzKgdG0rGyCa8LqfI7Uo5AEMxy4Mu2Xqw96xu8H/f12OzmIDFY+6H0HxWuBfdzOkLoJPGCFedNq
A9h48KewZtihhZYEAj8vi4sboQ+Z7nO/H86mLgjKRPYokz307I9EflZS0L2zjQJ1YygaqVgbP76k
qsjcTNxl1XDIdlkVwMh4pgrOqNNGwDtTiOFtNWJEAZ/MqNN6TUzlwobaXkj5dG45Uky3VfwG3DLb
RMlaFvzWQ8DnUwInSwnquqb0U7nHegYGuw1HrF6g+H0rkMuWE69f9RL/SoK93pnEbnFVv3LVSS0N
+/gdSLZ/NOYj+bCg1j8rXNEIUU8Sd1X2+9Hu0tNoKMJ2s0h2e4s14maYyf0wC7GirCGxt2owjh/2
QLFIX3C7oWDjNaub8drmlSfKR6T5JKOHy0tcuuAjbWbuiZ4me5rEJWSHGhVWhjU//Mvvy8gEA+nN
xNcq65cH9H42FAZnpwEt2IyT103vPx26YVa1DtE0/3yY2BKrXiaimsGXouHR8iwF2H3chjp6IUc4
WCeTTNmizrMyZtVEWLz34KF0+O5IDyI81xFyZ0XkRYQwLqHkNtEZI8F7qAprVg+cqGaGZTrvh1AI
d7YbMQ7QfJBum8xQUGWiyIZ0NlRPjzx1MMgYAJUUF0Ld0or/maT3X7WE3ggHnWHELLuCDuE5/G1z
lx6sJFYsMdovcmVaK4ACbeNMhDLOpNTxO18bQaIlfXUlFC8yOVz1xrmzNyVFYzaxd8oblcA3bejG
Hx5Pz+jUOQpIukE2tedPaOwD1B2j2hk28zJr9SYsnk7EoP26apfquzHVfXDJq/tsQ1zLBPRz36O3
2w3yN2GfPdWqpEGQHPwDrCzy2NQfVSx8qHh5IZOvsbNUKtY0tyWyKeGCBCGvUpUqEuo2eJrlTHHO
zscmsSimyRqyoHYCB7qAK91t5MWgJY/xd4A8FQCwNzCdBy4KQBTbvFb0qqQyFb9uXREYeqQeeoId
N/MbbwVZYIBDNMGrCy7Iuk9BcY3fqXrgUA7fDkZdTd2Kj3xWiPcUzEQZ78SdlrM0ap9ad548g4vZ
McKFkfB0BI0ZOtRHUGUAaxAqE/ntuaqpkM5oxnPfCFRDj9wz2xiD/g34YTziIWPioa9G4e3S9fpp
5UzkLU6919tnF7bbHuAchrLxJR17Wt7X3Ab7mGDZ8R/UTp0yzxj76B8dpoKYafToRXZvD6f80a4d
Jxcs++MkIrVF3zL5os0aUgKdadSIpXLs9BhyvqtLj6AlGuuIZvoiRy0WPhgAQMas/jt+Zh9dl630
QanPo/wkx5YHDC0hSSjCC909Tuggk2TQMrqj/c5Xl+Ecv3fU+3XStfKE2ojw1nHhB5V5KHyQcPcc
i+kZYqz3iYNn2lgjHgRdFOkCZszTB15GcpeLV7bAROv/2+gUGMAAyOoMT6TRaiQcC4yssPKzRXP8
A4FZCR3Dn52wnFBb/rcG242LjhxMY8jQ80E3mcybl7c5pbLJeIyKesSC8+OKhuT+7XEQRqhdZZfN
otm7sF4zcOrteBVIyLgvmkTTl1kP7KpMozSQa8tGLZjKAGOgiM1KM+rtQfvFk7tmrknjsIT21eLI
twlp30Sfe6LVsgAWCgr+aTuxVGjXGEdg4NupXR8m8YyosaPHmUOcz9M9WOCZylnjI9qLCqk4/Jnw
+naSCkjIEqCZ0o2CzkieEQbXwULfxXej8sdrt9sdUKHVsrbb5fQLmRuTlm2nTThzO0L4zI2PVRJy
SJuIHQjm17N7/QK14I8KqhNiNuKqCRXXOPn+lkB3fPfaiCVbHkIjIySPrd2hFIczsK28tIGpyJzg
0Bi1PkhuRoPj07MQt8bs96GLJCLtSZV174uzheT016m8daOcbfigqM/KhXHUHelGS0b0HI/qneQB
CCKf8i9aSCr3AJDCtSLEn2B9jfv8wh81BmhIn9yxy4AX1d8CxmSRyEq1nf1KgciKKiqUyhC0S1YP
aX1hEnoeT1Ze2st+B06WxGCmLN/yLfqIQnMIczs7ZsYutDzFsq0/8galR9gk5E1J/4cGU0V3+Vbt
13r2xGpf2iV7TbgoilMTnil5P8Mh5DddooTx+bQIkOgaSInBDHJ5EIzX2fMYoRFMoDUiyWpRYn2t
eeY/vczzXoxbKrxGDCk3CmLAVRRnPL/3KdnZCPXF16xmWm3Xhj5UMWpFACoXuLNGyBd3yexF/KXM
m7m6R24PZYEwe9tYoJ/+uKfg1bwnTZolXCOQkDrGwWfmmSEfAaS4oHUyAgWv3KwydAWvMHlZasrD
8BmACYPJrbtLuiWhFweB5g95Gq7W6em9Ma9LTC370UpNGe+ovxZykwkFPlEqNTpPtPJcT/6/0gcA
eYp5fhmvJFKeXE96fVaWmXRnQMYbHMnovHGTLugli0Rn5Bg1xOUDoBgNKQUwC8jQXncSUamrJLmX
M/GVJg+QWOPK9v5QOVYh8PQmZz4WEaYuK6vKyVFG4dKpNDudc6kA2GBJde7JmAuw9Qdz7CQG/+n6
9RFASeHTwcHop/237Q15o65kwK0YSA017XuAdzWKknCMQ4VRqt8N8/AfUjhcfRs1mpiElfzmqqjM
peNQecvwk3HEPI/X99mBKvOqXdQu6DWUH2JKjtEX2B6OpFg20bSh3KI/ctHjy9psABwChR2U+eEb
ycTz54DOZsTW6cQQlt9c+khDAw1TWZ2I3QSsVOkNc9opPkUV3UmsjRLj7NWSYNtJ6e7egNHWDfNE
2b/vjp2nHLCK8f/FdbvS3H4jsBZ8ralT9VkiMg6EkcR2UQzWW91TN4WzUwBc/H3aScn4YCaG6hZO
crMJrs5LDTEIVXdPhJ0AB9K7oULzAQJOTuPRU8RaEx2YRayabaRQRc5IxHhh+VYqwqjuk5xok/og
uc4BbthSoqLw6HrJk4ntbOlSKxSPiDak0mKgxA2bPeBBm4mfT0t6q8XXgVF4EClBSgLzEWuxA64j
5N7YeQQEFn7JrjJ6Je0w7y/jcp4H1XyyDH7+MOOQZp2UUDOnnd1rVtCp/D3BJooc1cxtCzcW8Bkx
JA887Xp0OS+xGhF8rtHeZZ4JKOiO5pYgL3Ifg+WqFvpuPXiIcTAqUapi4v5vsRe4t4TlHc07FpNP
NfLw0QpdEYLyxfmxF/FHuG7dgYMQPqeySdrFUyxJ5GWx89oDZgErqGnJlnvSBFnRsoXwOu9PcB2o
UxR1k1QJRDY6UN81uOOW/RXZNoU61YH7oTgbAa4Nig6J2cqu16eLsgGMUVVRF4nn5YXI3lwAE2DP
yla5NgH4kBRYe6IJ7exfZmuImOXHlfvMeHi7Uu2XMwBYdc6I4lmQ4yWTqP7WueYaQmJLZc2+dbbE
XiKhRwnzzuvFs3dwRJxbf3U6g/ZohhmrBM4YcL1/V3MT9bPirnJUJhgPAAiBeDLgqih18A3UVKHJ
bQAK9LSCqkr3duNGa2kOwxVdxbPZuOqKaexyxXinWwFKbDUIWhzgNoDPgq+zqx6gy3EQpSPEQgKQ
ZJ0mCZY/n4JnUVyZ1wtpjpMSYyciKwE8bfd9Qh/oB6ToKo7casCoDcvPb1/kVeiB9rYRSxY4j2cr
1Ly9kuesMeHkkLZdOs/hcZsDVqUyux1i9dTF2lz95aCGqbnmIBAeHoiV1Lb5wSvwfsI1KDZKlGam
PSLRwxPgM8ZHXtkDxNR4W7GPKweWLeK2Pl6q114iQViuBFvfFrOWu/h9neXz2mBglUWWZVAS95W7
dpb5uckhsqdNDLB0jg1/l/v40dRDYGDPa/6IE5bS6IwdOtw2EWcEQu8hSfS5mxh1SD0WD6W/4nX5
v/B8ESjiVyOe2K9vx+GKKKtdS5tq8icR2hUW5HtAJtnNhWVtiuwLyPl0+ZFZ5Ig7Z3mAFMox16gc
9ECm9qShBav00V314n3cTDD5DpHp2Jnx2dZ9csJs/u1qxIYX+SG4T0czvUtESwnyvSZ5zN6yCtu6
fu/1TBxPJQXNGCIJ1O4SgZyv4k0xVsk5K1lGc7fzWI63Cs3WLVJZJ5HA0yVoEDG0b1Ut8zjQSd1x
FSQYEQWxskB9s5YDBHS3o3zJwtD05eRWkS+VjkUQbJyq1/a/d8Q+Geyb7fOgD/EFb09eiiJc8p/R
x+YtloEhDm5+aFetOUeBKlNI7T21NC7wXj1buqVda9FrcsBl2c21FjMlEHoQrCT3qVwgxVWPQfMj
YnlfBOls+Fjih7d1JxWMev5iyAzlx2thy7O5QohXnD/O86rp4cOvqW4Uhbd1Djsy428l9LDpbVDq
ZQg2xaYYX14xvAUMnNW3GKIl8yr+b0fM1swX+v00MxfRWKYqHqRAwLDJJbRbfeNeiC7fiGzy0ixr
ljR/BdFWCb4t34JvgOth9G4Ax1Ry+AnmYcPgRDVXLITD46fgLONTK7QVnZxW3W2lIDEtRG1c7mOE
BZbbykUGNsoHp/IJQ+npxRb7G4E4f6fr64D5cB+75pCKae/hIOgwfb/AuQZVQiW2dgL+gfVtOL45
snjkiVxwLzguQbviE2rEhWLLwh3nEZVn/ttGpl62hEUWg7SUp55LPW83rCclj7lsGO/2Vhc7lWQh
rBiVIHyvEjabOrZ5w1DCGPX+/0ICPhsiwEQp3hYoE+Ycd5mkt2v8CIICfL3CUQ3lW5W1bAMT5fL/
HeED2fE2Yl9bI+J4MpyHVsUSJXLJJf7WH2YyWFvKx12+HDlkW+ONTNWPAMxSv/f9XmEHk/nYKPxz
rl/8dyPcb12iEA57+wKlDXavMx/Z5Y5+gA8V2IsMUMbVtOYNh/am+EwY/iM/RqQu7odapl2L7i3D
nely0Irw6E9mJipcW9DCv3+9OBkOw2UazbnQbvsA3LJ736/tnN3iPSAAI9KSh4xu/3AHwCGavg+q
jHr1MFuvjSYE/xLoJXL87E6/TY/NqtrPIdZRe1MJ8sgwpzaIQrVxsVpO6lY97UmLpd6fGerdicTl
0hmSl+XdFUjqwHWrYldEW+XLcgALOpdcYx8zIfCRXCKgermR6S/TCiNE6ij+yGsRdUbLzSI6SkAl
qFPxTt34MflgEJ/xCIo41FUDlRscStIs3iO5dRNv2lPPuj+VfmYII1YJpPj/xYIfnD50L/jtzQ7u
Bm1i/vD7ntudL4fJCWdIICKSTrCJA6Xzxkd0q6+8otUkqUIguyTvb3d8VBDzUTP0O0LrNtqWPdkS
3k08PUPIRucDIi2ojSAFMNtBwJQd8hxyJ+b9gd5CnW6lGV0KGgcXMlXB6LpEiQh/3W2i1bLG54K5
ii5A999UCOATqDzNdREaKbJm8v+L+42Ol8DfZyBu3vVMpuliiCAsg3tOUnoVXiARpwBCk5G9abb6
txeaRpe3s1SzB25m4rboGm+hjt7h9YCXao7PGr67w53S+Bx2YrAvl9r9kfQjx3aFFhKssTV/bn6k
IFd58HhrqFUIJlbbyI8UoVokQJV9lijPjLjumlRF8IVrpkXV2VYHHy1RL2bU5WAFu2EcJF41gX7S
IxrHxVfFcUSM1UTjnQzY6vsYyt/nIzAPWWsFZrnYKu7bJNMoELW1woHYzvw+hKMbsihvU7C+uzxG
uueIU2LtpTM4KY0Q+q8mZ8hxpomdl4hI1EQFRqRIik18cQRy+S3ZIrw+aQL4rI3JjRtItpHrGfAZ
lm4G4LG6E8Tyu1WU8PxQOPthRXONw7aTAVXijRjWowKjs271tFsnEPXUx7Ac4PU6mMUCkbyQCABk
TBciDYaQNzZynqQXDGusjjkEureSXr81PvUmg7KTqalTOhJ2Pbo0zZJCux3I04SxuMKwEwGdWxN+
IIHeVQEWfwOW9b0JIvMwuJBk+fn70OwrTwnWLu0zgKBsFC+eURR1wySLdGeiDY0sbkLAQ9mzDB92
gjYlXzYsnXVR4V7z66Koe4d6aK6ElSDGuHtbhNXOB9d6IPWEhA32q8HOYXjhZEXC/amYn2syRaQF
nbTc5ErXv63KsB8rW15jdD4ECMEYohOIqSLpJ/Ycl84vMo2fMgnrhsxygfIy9kr0Gz04FIoo+SPB
dx/L+eklY1UNtYKWbAPy8vDSkTwjEkP8CjSuWJM2V2pOAcwxUxgHy2C3W2qKQzEFHo1AjUR2IeRT
6sHoYuQSJat2q4YXXHhpSq+FGTh94gPaXCoDgGK5xuS5LU8I4kE9EB8tgq4TgFgbg40pNZD3NdHz
SPmHFoJtRnsgxoZkJdf/TSYXuzxvhuw+N/LWltn81JZ7kHQFcfj/K16PZ6viegiwKT990p93kFuF
UFXamchUzCHijHx7D+zlyS8Flcc+q49swa4hWtFGsgFd2sp9kGbETGOdGJb8+u84LMlvFhCjOLy3
XCr5P73fjnDz3+HDFTg2Uo1zvfdx9Ttvdd3ZrJ/hMsJa/IDs5A7KK2NvO4Dm68sI6TD/eGmpeRON
9NuRvHMCVfrUzBD/mVdhdFZk9V+nrLo4qandUqEV2oYB+N5qlrabvdj5dnDlmWP5+Ju/fJfeCkUt
0NnXZSynPmL+PP8VbipbhKLvArmkkyjLgc5u7bWeUg8/BeIVN5xGJNcjgAwY3PStyE4wh9xnbpmL
nBzJ3v6XO2Z2Z/4F/4TojrESzOjBw9N3fNNRt+k+Rdk8CHNigaU+sLBtjiWjdj0H2hp4gx+dseLe
mNLGdDUn5+hjmu0hjGkiYNkazxO+M779+Nco0Xr0ZHrDEcJa61yf+b+EhXmNRNTlkMjNYpOnQmIk
Thkrc/HvuOHU7PorVNvmG9AHd7z0HzAMIZlpqdpGQGohkaDwI54AYykqAZZxbaiy/Oqu5+jvJ0pB
KxPFrlYh/bOLIH5mg4aBuopqdmmA69I5oBohlPHGsvqYuEOrTKzW2oF0x06F3f4VE6o+2ph7vkx8
ozm/l5+rUI5ORG+MuZlZBjmOxT8hHspetMk6/523hxxtZB3LQi1UD6LPwE0R7ssqkDJtBsejpVS3
vTQNxRzT0vyzAaX0nTBQf+tdDMch27lAQhcBR6rQA2Ah8M1heTbHlKGsk4lgCQGA0U/lJDp1ijtX
MlrSXtHlckr2BcR50pOiU8Gtr8qEB3BpB3n1mGJ8kFetOUMiCSFgHFPHOiaAZL1LdObcoVtLe2NT
Dk5AEQ9BIL09RmzwUHZ7iz5j8m5hTdT8LF4wQbTy/ukClEpuUjx3sgIlIPjpiXDRL1XHe8zyBYKg
WZ0euJx9Ya47gAeD2DEGCCL69pVpeKp+vwKhVq28kvKr9mtM56wm08phm4Bgnw/G4jxcYo+QSFKd
nlwb/KEtqDbgWFvZx2Z0GVyfAx6jKgE6wkcAEL7OixsPWGBzdypXWDk1c0geSo2wpLpKbE5owREL
PIDGUmyOW775xhsGeRg95/0JiqeV+JrmvJ0b4MMCuHoBKQ2XR1teH/fkQa63oo2XS9AMt6djpx+U
B40RJ+LbzMwsvo2SzjDsuT+/fR+bafvd9PF27K5vkhTqB7DzYMkrlz54V9J3ONKpTA3nnxhgQNc7
DnzlyKhOT/isFeOsyg1SMuGkDLTOHqi80QlCGcy8CD4N6LCSAhjliOMRDmsqFyoLSo7Q8zhsM2e2
kc/OCnM22Bb7R0oR924BKFnIZysFNx2yADd4/KrpE4madJHV+OH0ejJ8Z6vS+EV6/mmwUQRTcuHc
4cUDuy2IFwsSGKnC2/8L6vAZ9lwG9PCiek8W0XeAq+KmkeZxXm7xbctiDVASRr5pzDnEPMrviUA8
lpeDfykhSfKZydQpZ8uPdhgaevktzNvFI/Reht8FMpGzPCMap5IRktlmHv5TVdxgOof47Gumvg7I
5+XN6jgndFIeUkkW2ys3IwEZJO5e5sK5pDKKL9vBjGvYx4UnaEmbaPOxA0F2dAvfelALoUurT6Jj
xLOmoawYbqN6LlqUkaiJ+mVi8SCDAPLjx8aBsahW/RlYqab1cXk1sQbX/4VqjBhPuftUkUzVrJrV
/qF1PXjDGXs/mLtt+8wHunJv6jMTmEOLQIDMFkm3u+w54IzDiyDgi9ibLvCxPlY3qh+t+8MBg+xw
Ja7rQ4Tpii2uL3+evvlwsWmBTlRWnks2im+VcAPdpnYzyFPVj2J7/MRVS9bC0FKUq98KcEI6qmn4
VlTAx7XUSerp6DPQTJFZCTWnCJznJP6RVZnVzZkTouL96mXiOJbKCcbL7pFhCJN6nvEsCKFXskIm
GNFmELH2f9Ki2BKtH5TG5JDKcaUpjljsG96oK4KXWMplAxdx1oCfZdIBqdOsOB3S99ijH7g+UYFv
RM0YuM7Cl/mOPCBAbk27bMpPplcDs+VgqsprLlnTU20sofJZE3thFDoW/0B3cAvhb41uEEpzP5dO
IjzDd7evSNVXEtdD+b4bc85DAeyZMeaysE2u0fWqI64fwSJMQ8C7KKFu5dN6m2FIZXkUSDj6v70T
Ge7Jh0bUb0M3gA4/zmNzVUXKyi8L+Pr6kWwE3rnzC8RPIikb4RfcpRaqre/OJpGEDPRMqFNfgOka
f3UhlR5g5Z8GjGmOEBB1z1HzkopaFsUfFUXfpeF7hYfzVprrFRtWC4P7jH2kvYkKQYr8V7TTzfVO
Aqb2uo4jeoz5hsj/+fhrEh+k7Wlyug6b/0F8tiFo33FgUaYH0SRBoj6Bwq/J7lw9Qv93eMssagXL
linmIyffjIH9xwDfn5UeLkuFvJsrt6om02J5APpSdMaorV/sX6KUQ2DN8ytUhPOHEkzVuWPfNFol
aj1z7cr5m6xKB8E5HKsrG/QOFamxYRRteGHS3oeITsLaVm8UpqT2TVx2H1bnUDDmJa/RuzDeNylY
5EIvNYSkFyGd37Hv8aXDb9siWf2XfBYqnALiaXpgC47Tbhr1/E9QPyFnigpeYkbJxwy3ywQ9TVCw
+Q2LKCp9jJm+lvCk4yr6tpoFcSvJ9ZexzOgIlM/VoXWblbC7YnH1VqQ8jZA+lceHO1X3HxL7W/vr
ynuJ3a8TanVtRMMvGDaNLy7TsHKzi2JpTz1wBhnT83ZCKbbjkfNBBVHQ1z9LckDqTs5eiUWMhocW
wb56IlsxwLhOosV6LXEmwhLfF7AcgsDxxQKvXe+IsuruW43ONvkX/C6Y+4mfZmsU8/Sb9BYjpdLY
dxpdkuCj6dXa3+bZ759tjiYE5LHPwiIqhEaL+1yPrPpU/JS+6gWgyt31mf3dz0ZWHTgl/IqvzcVk
7gv4ELYgApCAobhPG0INvzDZ7naKtpd5+yDPRF8AiMNXDcuN5NCwe19tjOBO9LRWYrwBn2I5So4+
WcmZl/y4oObimmZJCI9GotpetdAw6DUrsoa9vBAB+T6aQLE74bCSTJWtOo0Y2KY99CL3s1m28Bfu
qjJ1RCKUWfywckXgy/Qc4RW3AMVPwYx3Y73C+Tn61oKMNc2GV9Y+imAIXOtmUILdcMv/14yJhCFv
thzskuMK0SoJJuLLaL7+2gdJTxDAYungt2Du1YWbKBLxUV36byt5Vzo0c2xw7gghF/UF0kSvGGRd
hgSkid7BZaZaeSR0Mt73hO06AVqhtG8ovFHSYfJQK6N55U04KEqsXwqGAYcyJzftcsLIIpnFR+zo
dkILFk41yvclKnPWsOQ5xlJmcgVcgO8lJvT7Lh9bBNuTmYOfBy+dPIkqRpuugSfHpHnpvfCZIgdH
7f8NvcD+rIa+o4Ftci+6JsoUlxi1WLl4L59FiHD28ffVXvjp1efQozQb6j/DQv9jHkjcWiD8Jtz9
j7w5b2yPFVZirOW2fLnzI2qSRsKP+unLogkHlxEj+8D/50n4UFXm5uJ4qplDsD+JsCwtYCOhI1z+
Ao0gTaNOknCVY6dUZoUR+vUbc+Nf/8Hai6oM/P3ZXJxHMc70XbrvNiYwxMDhTGWVaQhkz9/PXE0i
mhvhmlFrjYd9IHkfsjo+1SzJsAWJPQYvsyYq7H23mwrGnIldAuf9nTe1QQwRR84anvqZVRagPUzS
leNrzPsri7uxfxKi3S7FPvSJrqQiXKQDrJp9eEw1OY2NTkWTjNIC90gzYVTNhudS92Sjd8f5+A1g
uNsW1QV2JB7wMAnspONN67LAjw2MRq2aWa6R0f7agC3Wez8yidnnkz/dM48zrE8Ojkr3J+AvwJr/
1lR904tOwdZMcgeTt6v3chfXycYjBUU7SFjeq5tG2bFln4vj/tuQvqcoYpolGPDMXsLYdoMA0Nv3
FlRozMMPlpotsxpxV9zBzU9Y9BphPwcH6voG1nh3RUEqj2PgZ43nssxNZg5mObfDs85QNe1nEcSB
2WXQiMphxWd8c0fpZhNDqvS8GPvv5zdJPqJTGJxec9ydd+f439Sav/rcJBnwLHG77nKq029mAA38
c3FZT/gemWlagDmUfeQkcrpd/xdLs5e8L1KTqGZjr9k5PXvVcD88UD3UShF9xjyR6VD6HeYd1Yvs
tmIYOXUNe4Xo4Lwku/tjeIfpVGxpiGRNfAxoegHMu9fXAJG4tVQot/XntBt7P/72IcdU1Tpc+B1Y
qo3nWP54QsjqE4LjSMWvjEB98/QT1VG0aHKKRgrH5yLQBTR1nyuvi29xOnbpSlixlzrgxBYxfJMY
fdI08lSOdeh9qgMblUWbFxZoRfDR2KcAuCwG0qRnfUZYo4uQ+RTxdap5GgDD8SyJqmZjN8suygtH
e5Dgla/pe8rwde/C8/i3g7zrC5xox3Z0h0MTVPEGogSea1tBn08X/LgVslyg/PfubmzmV6rGH7uC
95UiKjRtr/WKF3FlLjx5OE3UhAMWe7DotQ9UTZUWOJVPOk+i9fsAEDEMWw1IUOBsuGjtNG6Yxnsz
x9YFkoEcFO4QeNbXC62kYHFd9xccmcRZOy1HHg9rQEsH8fSyauGd4mttiMqeK/fsNytahsIexz0w
/o3kHjnEkxXUrakH7eRbj9RfItvMCu+wndU729S+LGL725YN/+xAPXLLoZb8rOCjQjlmps0iIu31
V9EQ5CI3+JFsenVv/OBC379JojpJ2ke4LkFm5bUgA+97kBA2YytL9DE3OsSbWa+0EevJQOcHg+NR
/J4TaSn1t58WPzRWcQrBiYPosstweH3BhES4dBNkXahOrGgiHK+HHfMeVi+JDZZK3b5vvlHl+RDe
dw8RilYz0OY6NZTUXwRwrhi4zBSygiKeYDa9RZdUIUElr7bd3PUAA4rvm3Lsgj2EeBONX9JVgd55
cJbUyrMqYlKP137JfDobeNIsku1S+OoQMydixR5BrS3n4nJloct/nlCDIYIiuy/bq2/Q3OeM8GS7
NM+0Ra5+TwAf5/5p/If/7OW6BWJuopAKTK+x89W5uIb6kR3c7FX6fkLBKccOiSc81HcSKjCCbYva
rwP1ZhCrVXuuuqEgvGNioyRuy1k6GImejcpiokXQnqwn15vA/jzHN4YkP8RLGRmQJas2EMKwmMOC
3jvAGpmIgFprNNLmsJMEqJ0eXp8YW1linDrDUF8+bphucCw+llw2jOOtzdbr0lgTy+GWODDE3GlC
j4NdQ9/zmAGDMTJ5UIisNPxJJusKkOmnc4XK0I8qj6ioqmEo3hxcfNhDP5El8D8yN/8gZzGt/X5v
VTJ0sfl7R0kk2k6fSpnUk2kzEEvdQieHhpTljVHrscgBrcZPa09M9NBQDfwGSLgAi3aW1Au3lXkw
QgnnYPuyPn3wkYeoV1BCs6wQvVIKI5HI24BFnScI/Z+FMlv8w32xShf7PQjERzNdqdffV/dkBjT9
GgpcSj93tLtyfDkcd44pHSFUESGO4gQ4RwDTHHKbnXR9nVtqheqPcJdB4u9TL4hZXRqEBMAGqEHE
IJdJ1eW41LDdbdD+x6wWdYv0njt/xq/ddyFBTWaDe9cwgmzkBFaTRpuIOBWa1DCFqt/sZQvM349F
EQDGbPA4iI/78PoSv2vEADTBrGl9aRYL64Es+4XZeogmezsvFoQmg5e3bBT8iptpRIDGCF5HnQvL
vavj2S4pRJn+3/gOeowHnv/v6DCVMK5lWMESb4o7iOl/uMM5Qt1svVIh7IEAaNS4KhRHLrv7+XZS
srDpRJCRaEAgiTgC1o1Vs/v5x7iDQLJh8BRg7s1g9rrEZyRsyjQ8JTH7dDOchw9YyFqnpTZF5Yb6
4WNZ3yNQnWTr2JkMaOLaKqjiWuO8gWcjk0cTb8e7X/hRLWXutKr6Wihk33pYfDO46fpsjlDzTuxJ
iogQ8qeM3060ZNAwfkXHuJCZP1HkEv3FqtyS3iObqqg1AY0PP1tmmhuHdNdLCqsGvaZsuJsIgAfp
jwjm3hI55Q+JaNVzIWSNhA4iFqzKRc3yQ983VWjkbLMbNUlrtmYey5segKn8mUm0VxD5Sx2JCTR5
16RY5wuemYfG06gL+pyEriI5fZv/09ycvheD4+U71Ed5/nHSX8IMzKyhCXrxRbDDp7qPAlcCFhSk
1FDnViDRu+WE9+Qz73yZEiICiww7g8/jeZQum1Y6jKFaF8mNLaDcPvBgesQcgjkXDKbWonDBgnD3
mA43hBEw/hEkOZobKvDKozrt22YuH/ZmdmleOEP/vyxzOutc2xd2eYh1cWvVQTUX5HXBMMkz64ki
oRErdrE7rqRJ5hFR2IYtGSoU2iFuHy8POJt6O+BSeIKdhJTVHvWSXg94d+SBnhlvHP6F+FfIgGeh
9r8qq1gk5D0V3aFGETLRd1HzignVYGwpHot4SI9anbviEh8PRnVRCI8eQPXjifYI6DIwGw9bNvRm
C4hDYXZTib+pgvSKI9hZqyXJw9YDRwIVthE76/1iLbUILaEk9oBHraKrOXL7DCjQuPGhV255PeaM
GYD4hRxueNweEJ3Y0rcVMMLTh+2t6O+CzgLaXDcaXisQTJdx+WcNy1xbct4EgGEU0RtaOkegNomD
x7PUrwjYGBsRvJpI8gf1paz18jbU2rk4WbIp0uPW1+w++KRI2zdxyCYzh624+vG1Il2B0JJ+fBoZ
pRA4+3UBsPCL9D9LA5EPoHyVTfYXairx1NfVUf2H49mquDgHyti0e+Y4pTTuLmvllpIyVwMxhiWS
Dq6Ier7N+b03xEAdp3DrEgfJnensv+FjwvH70/e2n+XDWCkD4tVIDSTkHbnC+JXlqC/Eil9XDeW3
7n4qpetgKHG65kmIj4yI6ndmuhh20VhOtzC/d4bKWSnUoeg3aeOFmDWuYRoQL2MEudxQ77LiGmfj
CKaC/QP+Uh4nRcfN354xhTBlRBxER6GYQC80wTGOxuTblutlq7j1UWPIdL93xPhl+VZIuuCahzBP
333gbDOO5m/gRiZ69/khSUJQ2kex9ERb+gM97KkBsGh3mttbGumyUeRjOAFalbEtoAqljjQ0per2
LjOnlbcBqJfmmyv66D/Pxbe6wtOzWqYCY6G6f6tOrd8kW4kuZLPmwWFc96/eyqys7mNn2CiRz6yt
C4sKXMAW5c4kSnB69sosODXH45iSBdE3C9XT3biR9aGx0rajSj2NNMSl84FP+vINE6t6aahhAGtG
W4FGPiKHsel+9OLffOkf1lVfDlvleRtLiPIQp9QPnLUmJ3RmNYYJeHGNR7OPF+M46PToDMoRRqpF
lX3PuIkzFZEmLhhd4julR0R5LNPbHJca2evZbRgXCk7APOIrtd/J7OLRO74A/SOome9fPbu1hqoF
VPhIue60EKxCr/8gjjTuUGfHumxDvjhRfkYAQDOMPjnPg+OGqbXcJKPtpdtCXvupt3oBovDPORZw
hBHKnhbYpU3Wy9KcLp+ECpQZATjQvlgsWOIvmYVpir8JLXEXr6UyAVJNfxUSuVGTgk/s4S+YP7pO
XhtTwn5/HDeSry0+zLe1tmvkE3CHmVw7JL9sw5TLvNNPZbUlGqZnDwtuSDioX3Pe5ZlUDz7bHo8Q
EDSiEycJfuR+MnVpzFfqsxzMz+DdnIXY5+arJYSFYv7TSDHYiT208B239rMp9BOkvCEXa9GVSnoR
Y5xPAsAXL0Yd/b0v9bofGfnFE6LyoUT9wwd1JR8MhCmvZrhcEYh1NyDMJ/v/KaNLBMpjiFAjwdfR
t+W7vlv84+TKikQ691/D6iYDpc8EjbRi8hMiBmN1+Ph7d7lG0qrwRIEtX9ReG0jINOl+rLVi7qcO
8Y82l8l5SIJiIg6qqAaZV0cusgosmzoYI7RdtIEWu7TR/fgrgchzie7mUkfjLH4KvBS1eAUgBVze
ot9Guoeb5ETx1MLemGau33Q8NbGI2XpgQZRtiEcoNCk9RRhB3xSlerOL0OnE+dw63LEu3o50qTkU
ZG80X2Jhn4k3QjdT+2UneMUFcYHJ9fuYHVwMPVgx7VSVwrbB3hZrFfcsKrYfsbQAmuUDqqn4NqZW
5QYslzrpLuWLZgbvBcfBLFiTiWDlkRwPqa/Jt91qDXvtaDR4Oc7dOph2j7Q+d3u+g/zlORphDjWO
CjS5PB13WbrxWL6oGg6ec0GicXbEXKSYegEaqk61YTpWNGx+elDN0hLtRfyFfcr+GtDHWD389u99
IKoG/dFbR5oUD6GAm67ldILdMey3RQDBa7+zsosjaAucZtWcXGGZ2XN7b1+s6jMACeze+mXVSKul
rB5sYvWrrKNOQPhUlVpDdCjCLsIBpKiG/otKQ3zRmhay5zc91a066T9PneYYpu3hxGFpFuHZFGI0
rIVG+KdTp4rK5w1zFR1yU2Rz3/3nowo2LG1XMHUURWI6dRFctKAdpiESiJMNMX8nZo3Cvk7LBg02
KSkqZqMPbtLez2dpXs3emUjoYjd4CsNQ0NxW90NOUz0Iz96rhwZlpzaB8sDTftDWes3+XG77tdhm
+wHeHfLIPeHEWTtCtfvifNdkJOcRhMXyqLnvwnL/JGaRlPz2tO7RLsV085tRjF8pTBRaBy1Ov3A0
fX9Yzge4lm17npjmpD+gaQ7uP1R4jfrcgdM/yMzod1XSJmkobI1xTi9W95WT2bxpS/nk2ilhmSfY
+eQq+K0v3SylTvFWZeshYQz7saVxmcuhhfGUtlicuVgSyH6lo289s6ooIJQuQhYxn1Rmr0GDjk7P
EUR7nWKGySJrAFnQqA3PA2dwCHnhzvZJkTf7K5RsaVrU5Sa8xwl47ATP9qQ4OV8CtDFlWThgZ2Pn
ytAl1PJ2RPUVe1EOfIMe1GFcynsZHKd9ubGHViUGC6QPT8ms6/OAgWwL1Lbe5LMpQR0Sz/cCVsW9
LM9ZdOgUL091ElrB+VuhqruFZ6BJuwsRXh/Kq3ecTwrXu8G5yQqsOfvq/k/7D/6/RRZh47EDSPzi
yeXhac9jwk0iEACLQb70+Ui6F38xLPMm/WFydfCjs8IyRDPvn8S0OS1z1c5/cfmiRiAsvZe6L5Zd
oOl4yPxk6c42LuznvnkBNf7V0DhrSynvTdu2NbU/FLTPMvcQYymPvpMZCV85iDMGltKW7Y4LiGA0
jzWaw8CZg+VUUR7/4fRisHPjcDoenX0YOsiQGpzG5UF8Kn7x1vcUSwYB5gU0jGEFp+zmWsjtGjRf
4Cllh51b1eI+pW5qX5bGEsRni/eEei/EMLH0M8hSO0eRscasP1784Nniu6x6LjoeRA93T1oB1527
ahkwAnsUzuCtStRmwMo+r6dayTiMYVSrjdB5vGF5HN4jcI14XagvHBe49MZ1n7sllnFWVymm7HHh
t+2OInUhBzQmI7GKUhFveU06MKBezssiEYC1S2CxdOVH13eeAlUPGlHg7nHrNbGebBlBeM30Oh/8
hBQDgem6P1MhX6QmH887Wsxw/JLcuSkjfh4nQY4932zIb++2c7z69tx6JxnF8FMdDl9mihrj14q/
ZA1enFE3ws8e2fGFAuffQpzXUOMPaRcCTxkPo1hPrwiR4lZO1w4XFGdIv6e7UPVpZf1xPG6ZX+Gp
HrdLMBeI8Kyw0h0s+5lRECYRSbVVTWNAQwJmvKA2UbyLyDP/U0oO9k+8hA00M7qMDG3TiFeWwASO
Pci2Auogk39YVLxtliB7O7+TcH0z+Di3Wj2tRYQypLvF4iVZvk3qodNJVR+AeBUAYDEN7kKOj60H
XU4qhidxYCicIf7xM1jEowVz9xPWV/PM6RepqK+9s8EpPG+1/rKFWs0KhSouBV+FJDlV8vhBSH3n
YTSrhKDujIx/S5jGsecScJ5UAV5N4AcD/AOtMyp0stpTtl7Ppc3tc96X3cg4/zIZLV1qbdgk4jxZ
Cx2I2PUPg449PyGQrT5/BjOzdDohgQr26GoHLgqY/2xjnq9tE+NMO8qUP7ervDIdcyn4cpoCfMu1
X3u3QtTJpvi2KFaCtJ1gU/yFIoqRCRPsSp7N1O2rpEPbmPDEreo5aFOhYgsUMixlRpBCPsq8sKg1
fqGKxLM75HdJFCJSSRq7Wo/J4I/JW5RsuVsFs2ItRAMjo6vfLgiUpzt4r4MABWp8I/IXOjczfR4Q
Uwf9eIRApsc27j1GzODYJQWdCanqu6TXXIMMCdD5MID79GltDD3H64qIUOvdxVf4OdZ7GGJrQ8Jc
xNtiZ6NyTVv6CrHW7kvF6eNb9QGVUCKn2JwED8qN/pcVkXV99RmSWvmgKqBxmvOvcZfz8abC6qSH
w3wXM9hIFE5YWC6g3PvI5Q7Y0MSO0dKnwbE87n1QnXrkIEaCRb2ib/CnLPeqBjr/ZTZohDz3WwgT
FlNfLoXF6/hFPwTz0W8/GPCR0sWnDPpiGwmShWLzliAWwPySsY9JzIsmG8bQouQ+aLs5aXO2MaiR
vKaIL6J60A+TSkFv4Av5jF229PdNuwAB9ptaw4eLHOkd762uapsg6MQtbPnRQiul4Z54yqvPmPM4
aFptBBGtK0y6+w6G82kaSjWJlKMCObHdxWI0JkE3N/jQrDcNoI+gMYoWwk6vVKFye+CrVzzGow2n
w8aqTS1+Fuagg23oQ5+3n2NCLVBdwhiW9JoTVWKhGovfz6oPZN4fHzDb7KMjBpESiY9gmGjJaq8P
aKB8Zv9bl2rFfb0tpPAedHw5i/iB3PRzQYlAuAg7yuubQ3s2MJSx4szxQpyRjspya1WIhr/ttZr+
cNByOkFEtdlOZG2I380E40cONUHcpQXTidjJ8xxYiGtyNfpV3LHK0tJZqL5r5Y0e4eSf1cl8UPUq
SpyRhnclWRyHe8AxxHoqxWqbRrx3GKTayVKnmG7ZeA89sINN7u4k+wPVuFc052hky8bOM9ErfqCo
ErtNfNMsBWZvRVsb50IVad90VDZVVHeaIvQV5kK+VT4bWKmWEsFN4L03aB3HWHqCDXeXhOj8GIje
3CKYx82NhLem8ZVCx4cAJn5PDWMADxDtcpKuh+Upvpyqx47YWTJG4wIMcTzksGPBnd/il+peRJxr
1YHoPDtdHBQ2+74BU+kD/hkfdtY+DwyYfvw5tJopVjnijcj56+/BumdwpLk5lqmSRfiWAWJe99ux
ZM+DBX3AOSQJyq9fOAGWzoCk1k4SlFZmcTl+h33hkhBBgR/beVFoO1Ah3hBr8BOGpFKRhvTAqUvN
xxijffwQjyGqYVtqdkmfU6uYTMZvSNFQOch5v0XwQC/wGI72LyOi+kyPo7RLnb5vm4tMRi+7FVq5
nBgQ9bJgfv6+HbOaP+PHwFDrL68g2Us3kKqP8o6cWnPSOp6/kY9+ESktE+Ecn4HAun3TlaRj//a9
0WKtz2396PBeb5k04IJDRS7Zm1+JU+//4fc23cblHM5W5VtSauUC8Am/cH5HZHgD5Vaxd1sr3Qo7
NhGTic2hbNYfaIuOoWu8IkNXG4it2KvpZn8lTvXToxkYQRGLv8ed1INl28eNWeHdirpgpxVVUO9q
Xk3H+cGKrffE7oZmhubHI3+Bg18NCCpgYt8IBZrkQau2IBlD9da35zASojckRBTabdyQGepEDGJE
RbVFjxqgRaETZqS1L3zEZZvCJyQgf600B3Hms5Zk0tJ3sJS1o4SnoJB70a8GuSNKH2pnl2su7LqR
tnA0FYBgrfqH8yZbBnA8GBqnac9Kr1/35NRBRrT0b1Ipfgp5vKa01vJ6ZSlDIClSyX7qopl2kWyA
tVOfoecIHoVQXdE+Fr+eSEdbcONXtNgUSBVHJ/D6/fdQaWTxQdqWdnFRkTaR7yGFLM/SW7Z0qYc+
m5a+J5LuibvLA6IhR5wJB9imgfVfZPLwikNSnt2DbFNi6cgMSyIqa3T6SmIKT9GXGI/8VDNuuipI
EQH+SWe8tiJP7EkujU2FRRsSA3hakUmP0+EDzDUy+eW4E2IehnML+53bb5ye4tt4txiAzw7AAeAC
kElRR3XOje6Z/LemfCu/Ock8/wYBts+0Wr4lu5lLpIT14m8vgzMKKgJ6vfBqZc1ynQP/+XngKkX/
gdtOuvoTuCU1/ApxvrGsdKo68lObTLml7i7b78NwXNVyqGJQm7U6+pJVXSfnyY1ri+ppL+TSNpuw
vIlpuqKQYtitCoz7fIyJPm/bex7V99E+oQVkwvMnmmxbqUR03NFYI+qwZf9aP4PehN9mIDLrTtPC
x8kG50JTX+oz8nhMItCEKEMiVmgnF8WjILbBWZt16jCmoiXYpJX0eB0GCHSTqkFpQ7sgzN/J4jE9
kBoaf6zVKPWmqa62P2fEL9aQn6qzN1fz3d68bOGFxg3FVh3Nj7USLuoUBDTczkIAI+9csTk89Xdu
mLAZkC1OwRTiw3r7Z84Jqh+VIKXH8Kn+YysX3L2AX53t5FmXcqcRRUIx+RLsmu95e68mTxNvH5sy
XNnXbHB7VOrFYWtwIA6Bscts6uOdbe/5zBYd/uNG+lsthumo8xBL4F5jeCW+XSvntztHTYFHyFm6
20KEQue1ObXHJseI5KGw9kDMF+bOUhN0bcLvb2OVDJw79FsYzK5IVbwLZ0Jy+zfIiMEOcVogPj3e
hM+Jq4iG3S+mb01UZVtOw3Khm4HlCiTUdIXDfWHHmHyHaOgljZJmZUUBRIIp3gjkAM2PY+jD1mUi
0kdxKQrgUryhSitBWukJwVHcB5fIpZ2dVwl+4qjlcQTX24nCMtGULWRgPulN5JYAfOE11fRmz9ue
tWXeFxMZwutm02RXhL/OBI5ypLciL0rKW/8NUGW/gKfo5Robku4cgiVCKAmLhUEEexSBXo3YUfj7
y2mCRW5BQrrHuCYMUBUgh2X/NiyMzqZUD/msFRAtUa58PXIoOtPrh1gTu6Jt0kJaX3DnNFi9rw1X
kMOu0dtpB9UJubPi4J12Oj0vsj0bv6YxoRRp4pjFpSSG3Lu9vWb+zcl8CcI5bZBJoRIgsqUZLCMN
1oJel2W1d9YUU9bqt+pEfoXCgLxrK4FWLt6ETP7WIU14jGLtPNqUC9+H9rglHi5vXpPgMWSA2EfU
e6K8P6Ro8C4W4xCHjxF3XfnUV5yhNzvGBGkCWrpP3coJvo+xb696Hd2RyLFWF0xaKeK9xHgIqdod
Xep6UjqIBLIi8q+4iXvZLew6zjN4HbTb3c2SgeCI+lgi6yROdGPW8rjh/f1uBwW2DvkSlj7c/Cwx
e2HJMsO8JyvIc/R2AkKvRAfGtryA8UcQFcuOj5OVi7TEqG5z34HM1dLLY01n/XeXvq12rutPzrAe
JqqMJhqqPw85zSug+cXvEigw6D1072ClMNPDd5HW3TjHnotmwro4d9I2KgE0FdSjyqMvL57ijQKt
PLTF/djmtaO/CsOvIhgmlhPfzoog+daSpv3ie0kotVoj3SuqhpS0w6HYVlpyWiaItEK0JlRqc+0f
4w9m2hgu33dXeXumg7GOLMAxW3TDKIuvxNNCrKk5zA9Wj9NPxjgA5UwbqkjG4p1lzv/GqwlEjw9N
xIaB9n6hghWCZmHYLNsuzjavmol69XQp6J7cQ+sayF0AV/V5VyWiBQbH2B5tfkxYKD53vPw2OZ9p
YMmbd+sDuAuRPwk1br8Pm87/GRq/dmmglGE47yzmqvDn3txyZwTWUfMwrFBz/yvZklC6uyffPuoY
8ZHzva1JsVv/RaK1wAmMGiDhu2M8QhNFAtt6D5leK8aTAfTWgv31UzGa+EHdOWlhybXnmFoQLpzs
44hKVM6PVoRzkCzXJceyYmPa9DhJg/6CPEVddyyFR2flUfvAV5WlZ0ribls4Oo+VC1wceZwSxOal
jL6CWxgHbTbqiOsFQeXcYb7Tagv4MV9aSLbeaL+ORhSuSRmpedoFae7dYE1virvtX7EipC/68DA1
Scqd4fH8YqgP4PcPfNiDPMgbGeawhB8DL4l7uDpL2HwlYSa50T681p80vWwQWZatfwpdA4mUM5gc
6h+cJuLdrjBY1kLpDUrUxFvGxciicV+/9vDUMHtEgVw/vEBS/J9GuhLmOCmzpRoIsXdmZqMy2H/C
17LGKLZf7YYvzJZ6uWADrflYgpOXRpkSLey7UtCA4yhL3+lyFClpr/2gkYLk+dslga46h/jbLapa
kctSPQGoiojhrbaOAb3CGHKPf5bLL+v+Gyoy0mquLS4MC9WrsZldld2M5kLsYHmQkymZQv9rzfSA
79H5cJtGpFM695kThBRN97PaosA9Ibc/euaXj7EXGLzin9P2huG75o0qS4dN1+nZJjT+zcska+wb
LqX2UGp5sbVjrl3gaHrUlJCXvoZSRq/lORyLSoKfsR/WO9eZxPgln2ka1mpD8ShP8Wc5FV/x5blK
MwRX0GXwHi5qRjS5YqRG5hdXUrirAkgTVJKCCoFFDM5hS+TyQIVeEREqSFz4CigXFjfLjQ605Zu+
gnEaUZCjzppwBAqzQ5lo7l5VgGL4g9sLtRmugRllGgCPp8yNeLLEq9zSQeSBLQDlYPyiqdy+nNDu
2Dj8Hmp5e5Di4ynr7KcSAEqrvxfFtbRxc3Psu8wmiTAQQmUW96OpXTww0C6Dz56kDYGv+rieNCm5
dT+e9BLUSrLM4gwjXV6vLXWZMLOiaK4zpTrctXWULfqLCH8Rlk+QRqDDxKzO6erI5HtO0Xq5A2DL
3Z1yklZ0O0LWnss+Y/NENqjK+9z12b397UGNHNaIww8S5Y/KEkmvJ+bnGdRJmE/EnXVnWLFZqcZu
hDGMqCpilKfIumxL3AJntXpTD2UXnszj6TlQyJUJcgL1ijWf3WeU9ogndimV69G+cZSPo7Go+bmb
QRdNU0xNE70Ryd32jHua+kA7BPNW3DGXgMeHrrn11UYpTRu0Psdfzdm7L9nkMW3SrIZwFiJIDgP7
Saph0E6GJNta+gJnbRzXZEb27XJxsW5Co8ijpinUmkxJvdnct/hoE76GgVJNZ5rN1vR1nqH/VUjd
h6NB1Yn28y31pfyi3TUdnCZQOLZfjfVYqh2Vz9DyfnhaKRDU8wwUa8qhpnq2lXZm4EfHHvNTuDji
3doc2R/KhjIEjkXkBvRVCnV/oPy961HTYyhF3obgZqLU+PTHQRHvjJqYQvzBYcL5XCci4HvAa6Q+
XUQjXgXp69gvgG1wtrJtEKdNQe/pCieX+qQ/aTQncIwSNbjUKl5L0db/WJd6EWibqtEwBmkFsiSN
GWUSJbfo0fNGaWVrluXjOpERy+q2Yb96HTbjWow5QJrNjzYAxxEpzY6dHdGbPVC0XXW3NohjawWY
onemZCsC0j5bXeWTE/jJpNt2r5+RWMAK77Esi5GBw2qaTS9zuvAO8Nfy+w9RMj7ifQ9k4kLauTFY
W6bGASI4PWQz6HFyIgd9NlNZzH8zxEj+ZPU8ev3nT42YrZ0eUt9Agy0x20eXhASpiOoPqlQWPgIY
Z6KwfuTBVLQr5zkyrqXztRQmAuZ/nMYw3LVCjHXe/k3BXrCXVhjzhtvi+VJPZopNyt2VdsEgPiaB
+xwWMMYMrvz9NK2vaeORL384vH6DW6mnoaHfmjg4XridNr7r5XY26pJooXfAAUL9FkEeKeTMRZbH
LBeGtR8ULpkpGw8ytfJHnYCbW8xP6zuhM/otsi4NOd3pMdCcn3hTXsAgOu76Qb8lp7Oqg71Jean9
lpyuGVSwFfceSY9YOVtXJF3QkT+5TiroLemnLdal3o8pJHfRnOrRq4S9O1xBp58OuS/lCRAWSTVJ
Lgdn2cWQq54cZMrofJwuCi4D1gyy5firY1ccsVKHq3LdHPxQh8mNKw0LGQY4dMhxo/B0M6yJBVK5
ETx4NRkhN5vuUTQhy22jRxNh7p2T1L9C3HkuoZ/P4CfD1hcER1tA23k3erhjFlp2BBuRnIn0zk15
BiOSkET6CEeXRS/f77OsNvUD4lg1Z9z+F5J/QF56Dod9Wp5jrp4o7TVlLV78B5EAAF/Qs1bn9Gd8
bh38kuuLCLSVKJkwngzAukcc/aMfF4Ekl4Kb6Z7KUOxPmgdRWc5tTIYWwWqeNTzeZPA4cnfMhrEP
cKM7Opkr+b94FkKc1W0zyM0HzKRKDHeoqf8lQHHOLxBU/f0yHd0PUd5m0AqVI+QHcMbfbT4GyPff
ZyRwTu2osIkI/pcE8MEmJcHvr/GWmyal0hsT9ezKHNVb7gZuibQPnIXKMWqgXFTkBy5Q87QAUhr2
bsUYzZ5egGwx8j/35uj7DHGPdoVLoM+ouno0w0OCr5CMMogLSUZMdWaW/jsqsL6/DpyVrfCv9pEl
nJ88d6wNau07T5AobcTBF447N1N8va1ve+mSFBJq1UGggoz+i+NP2r9LkSlOOu+BO3FjCDGwjM9e
jzQi7yMXDi5tQcYLIGhU1d4vA21q4WR/kYpMN0GUcAaM/GkuN4lZxVuP9NwzX6l2qDZYG4EX8eUk
VRKvYIZfnefWtO5GArBxHHGp2bAoblBVUYQmYm2KeEewNVH1Xzqp8QYq4/CPrVDdqrozkZ9ZjjZu
Yx73HsSuyxRoHR7KOImv0jJX7aAlL7hW0JUhHlMees0A5rdciMEzpUPWwIQDPRb1YtGehu1TJFnS
3Bquqc+uaYKeUUy0Ng9J7EV0UyM8xCtbf3BC+X7Mp08dhT+aqBzLhUGtKaJr9qfFJpcQke91QPE0
mMfd7EKXagtj+MRLfFNuBav0YFCSrSrj1fZKjD3Um1RfEyjhi5fbwEOx8uibyoHIM5upme820/vn
skVtcJ61CDjp99HfyBCMiSX/aGbkfVnk60Ms0yhpIWt67OLngegWNu+wV9DtdFKZZguD31OBVtS6
St4cd8byBptllWTasS+Qf5T/iaUIDK/L4aS5NQ5MQyUSFkrC2CRgppvEPqNzhx0lGR3A5PswKDQ2
Dx3sIsdMZAZkHYOn6AfIt7QLM/cpqgUCf1F5Dn+oFey1iyM1cZpIAm/EgUUEjWG87LE3jYDhoqKe
kjZa3n6eYecXJmbyB3+va3Bm/hLJVd3UMEpaDq1sL32NZvps9jK/aPiMrI3QxSKzPVozjoCO67KJ
mOxiUxUDPRHm6FC72p0urcKmCFU0ScLwnsboMIgInwJeuKt1m3//BvOTWjGrgsNHuBsu8brFhYTk
9tH4jhKYXrBHg1jchnbb6EqmX5lcbR9ygxOhf7O5XaAOfTC7Ra54vrk55/jHr4Z1L+S8OsbMACZ0
yt6Qi1XZr4Z9bi+3pt+O3xDgzrII/WwgfRRETZUNXMpNnBzBOCIYp1g1LIFpuR7hV7TSBZllUmKn
ToqNTJfHTSriwOgTdfVAg672rIUeOapZ4BM5bOsys6wtPEigAML+H3DMFA05eRox+whnz5PLrqYe
LxeN5UcPugYDuPwi27wZSPF3OQ807qw8gHPil96flb5O+P3V3b3foQucXK1dl+cbfBLiMkB0Aesf
m6OL23DJ2ChGYMHXTYu+frev1BHdy97MB/soVZlESr6Xjk20T1ZimjeUMvHToLWByUXmw1k0GVPL
CNW9THreTI0RWHUnwW/AP6zl8mfEX3N0uhCLikurGAGsd6qZDaojXUlQUycoILrPZ0/GVCIUT+v+
MMfRIabtHPPyK8KsCQmx6zM2cZgPZaH7LbyCae44L5voMSnSpvc0vx3SPMRaYturcyUznZQerFIg
egAeEbUBjg/p+oO9Vrbp1XIGzHNXlSq5ldLVIKujs+fG8qf5flc4uVP9VvtZLF+Qtwg8SMDQJN58
XilMA/h85yGmcYMW2QMDVEQgc65q3lFyxKqWHQVsy91wTCdd+E+zKQgjr2LE5ceWc/EcjRFGESIU
s4Q1VNa6CkmZGDRa+/bORS8CxuC10NY+PpYJGD9Jr2v2zDFSl+pOVQrFxXUAjzlKELijZR0H+Oen
FR6ASVIcMhq4lUWQmqJH6IgYHFLtmGUlayE7jUzzgSsq5/dL7ZSudEHES6ocSCSD10vQtke7fXF0
UQt0T2KEX1Buz3TR79vBpbzGc168hkw5JoDKO4bwT3/aNsIVndu1DTiCImGLnUVLFiq6xWM1FQot
UshvUPIP+l5L8E0n+Vc3CScL9Oowf20/aHAAMcTQPZS6VEt8+ZUTrLaCNyBhJaR1m2Z6S+4MLrXc
X+5oV8kLOzbD8UHehexKGWFsHoM6D2OjHip0/0ibt9FM9qyGUiiTt0VBAz3nAsHAjl8bNHvAVNG3
mfgCKqARMZBV8t09OT/AvbIOHDQQtslZFVlag2EQ9+DvcFS2sjeZtKlvJdM2Pd4JkPgPf8W8Xk+M
S1uUbDD6RWgUak0d+4nZjrybmIRZ+lZO4+rT6L9I5vwLcF7IsQXj+SUwZ54OFQf8JZAr1AyLtX4P
BYZ9Xwhv8N6g1gcllNdTt/EwJ6JFDppz4zbtuTOODv+ohz5dSkx34n245ZJw5Rs9B7dG9Eb5bnDW
ZduSHFOEyYm8kXTsbxRn9mL1M5K3lqTrgN1yw3bcPOfDpaQxpXRobo1sHKUOzk3yHPcKEDSui/8g
iS0nGh0SL2UcGXs64CaRnDgt9XkXtCyQeJF/mrKvFPTRXQBXeJTK5SQvPEIija8XNao8J58EmB43
RV1kzHq6HycFbsS2vBQihQ121pP/lnUEG8oWVNZ3Dj0HfmTW96Dg8g24wA1INvmb7rYsIqYMFHsr
meQNQaZRkGjYK6yTW2rgkJ6xolUFCXQGzWwpvNfoWlbuPCB1oUKf09BgyP5awK7tlYldckcHOQkK
4filBzlAiVcqKSZOVMujp5lqqlqXsEYv2ttDaTLjMAzS7hMqyllJ7Uy86RseHFSc+1RCsp2TCPTY
tFKTTxjrAOH3RVFtkpbs//XnugxtQr4n6GMvNmBCUmIK1CV7LTinRY46rSBxzR/gYqovF2xioXT5
vodivbSepSiSZd3cN1vbp393QOFqswPCIZIpre0sS8bfHMBVgz+XYaWecVQgukixyNe0gT4BzvZk
DOsgpe0adV8gynEJsprwS1pI82h45GvH2sf4yHnu+Aqa9DucBHxmesuuwWQcpQR1+tqpgq+s2K8e
Ub+TMHLldmoHLC5EgmEmgXysuB4FGkW7TWxR4MOa3ySwpJdS7OacVGpP3YLMKqUYh5zEIy7hSqXe
wD0cxnkmO8wI2MGeT3tMd4FW1jJAtBGLRIYgATA5kZV//0jujeB3uT5smJSMQkqQgMcRJcKh3O6n
5JMunGg7RBcAA2A6JnP4gdOWuJpe1IIC1zTUw4qHZl+xURQHWOIRQxW5bc3RgNgPij82DlV/nFno
tnG3JvQb/BAbKl2QFBJDJRXIrgaWJEilv2pgqzv5oNmRab2N4ZM0sdfUiEncQR/Q/2VPNfr8IINh
o+0xLhQPNms640ge6MyJzuV/mMeBxYiRJv+SGUTHZv3q3ZE3Lgt41Xh5qcQ3d5vovbmcUmeDXkVf
OoUCVzV7eONchShREw6Ef7eXrHocdKaet88Eb2o8hBrJqHzfwbbeyHFkqcIhZgmZknG3RAs7DA3+
fQkIlMHe3KBIDl6nchKTvys6T60IrkOIoHcusydsC1y9pvI/cST0IM8pv/VePJjlynDvhFyK6ncQ
US7UpFbAYDrdomebQ7ycVkO8fNbrxaozrgc/AfjU1Bq9wgNwvILWlwFjzePmMIzpyE+fJzJyaXQM
ZVYcXAWNHlfFcQclWU/HM5oX82I2ulvXvIdLCddWP0oG9+BViCI3/naJk9iy0M/n2XoPX0qW9za6
WVCJ+bppaDBgcO7M3ODjeljECnGkev/sYMqF6t7VIZOMgJExCazrmouYVMC61VI6cb4OqJIhcrdt
wrdedEVuMwixO19zA+U/on3+4X/d6ecKiX3BmXwwz0hDiQdM6bxN5ZpIguqzZ/uvyUt8c5DlTjzi
Stdx4q8Roh1IIy7xi7Waz6pm+K5nO4QOVnBQ/qT3v1vn85bHiSZ17bwp1mZGbDnpsmpnCyLcadMN
3sJy0KHLlTBtfEYEr1u/err3sbeZ6rw469Q5VULceKW+XFSS0oyPE9M+2eXBHBN99On7j/yKdgZe
d4it4gK/7njZe8atjPcd8emnseVu73igWD6ulBULoYp7ixVFzb9aiqnFCIxRZiy2qqJk8MIcDNBN
BxAKsnZ++OplhGZXaiDhDrB4ZG44hHMltZzUhhm0wNS7X2ETReyCyjBBWFpp38kE3o3ClxwUONCf
xob2EuYjlDUk0N40rwHLfZPBQECmIUOODkjGtXpndpIdXM6Sh86mba35uHR5HYqfzYK2va1xZ0pl
MjtRTKD469rG/UXQqbikCHxp1HF5j5pnhYyVIL/ZT0gkujbn8IzF4vD/LBc1Mwd/Akaa4H9RmPoz
kQKzCM1L41st8dbrw9CjsWudIjfIlNPDndqpzgTUtYLsx8OMKAXY8LGoLpN+QIY3O+ZDbxyXgTbI
8PHGN9jD91WEYnHcYGW7o95ymcU1IgcNoeinuUmykM232nYvPLJgcPJtcUo0F40yeqlgTvpRxHqs
QqP4eWSiW3EwpEpYtySatfHDLlO4SSmt4ORoNzDJnaMAVZb7ym7S++ufdbIAZb2EaObsEJhvMBbo
IyegpPogQuIm9+xpaXQI/+dm2YrLZvJ3OSIBS9jYnSFbQLB2xdrSikkjkRC1oQ0VEXurbRaxb8xn
RU8C442I22mses0aTz+S2bIfN20ybDXom+kkh0301gI7hbWuuQhecyMgSViJJeT2CU+BEQ9yfl0x
VcRxmkrmWEyRvL4SgpSQmMTn32S+quQVL3G9mHgTNpl/tRurInDnOfD4W/N+nY015OAOlh1mBz97
aWD8QcG7kmfQzBXNJXJIp1mlPYHMxgrqyWGnFRkYHAd12PDxwhofjb7jcq4xerfB/SKAwAd8MtBg
xpvLvhafSW4f73kcFo8IED89JBwO9YlJcQ3PZgUTXW/6Ljt8yFbRVGwFVJuie873E2O04XJZR5Se
ygiKBp8hV3v5Dvjb/gqRcyzyfYCsvBbYqWdXe+msK2rpgp5W9E9qYR3pGYuXxQUcfZoVC97s/FrU
1JVYcZyaqrvVCiYKKQQKTScEp9zUnOXekC++JU59x57TH3itS2UcCqwnvn2/uR2DoKwOwE2WwJa9
fs/Z4ZnDpvRzAobTHiPPwLOrvbNTZrfl0uk8TN1r/lHdKO8TsAKP/GjkWUtlB/BV4GxV6bJTUL+O
8oVVIYT6C7L8S4m6oB6TFBEvqzv9cv8IUKs5+O6pMr07kPF/6pw6ey9/dKErwteRgLoozuuz+eQ5
p3Y+rJm/9bpk58yooPOqmNSHT3NarNXQPmfGdPkL9JXeN5lYhNvzhY2FRTZmbH82y76k2eiBnDvY
T2IQe20SAw8zj9E9vxyJgTytAOVIIubkE1y4i+i5Z/Myc0tL0YlBwifkF31ikcxwgqw6ZxkbKHbO
04kToEistPGNFUF+ctzQv0mCyjNyaCg2x/FnTTk3fCj9dHaslU6/ZjF+DIk0WysIUGE3UuG4Fw02
Yqjho03gLZyIbWD3JohltQ01ppipZPEuCkoYsqSdM0RkyJBoVhfsk6e90csjrqLmMQ7jNu7dWpxz
61GxQyaWs1yPT9d2Sij5LhFLkhDpT+ZC9pz6rj3/LUAh1CMeFI50S1YAg66YLZe+Re0qBE8nMpvE
YwrQPeWWdpDnlOQ9BePf8jaS670uBxLcmOWXWwZFJoh5ycQiMeDpb+n8IOow4lYshRFvYEWygO4U
Jnx/SZpxx5BNnFPHmOrOcxNt9rsKEP42CAVj/YHjHqpd+zWpXP4OgaFBJuPUH2GPsB6ePZ4BMKQf
oTD8RHi5heGbVcaG3tyN0ySdu2LfpRCsGlxcluf4fLTOSdnv5UhPEqo+71BDCjfwjiPURXMbMu74
tTUCDxvCjsdikeV+0wD1hRAiayAU8fakoa0xOXesvQrLK7Vc572qXibxLcnIv4KW9HvsX3V6uXYJ
CK5RAc+WaxQtv+RX6dYWG0HVbTFmu9Pk5KSrlKLnYhDcz5jiIYe+JoyZYlYHH8ayXISHkWfYqWHO
bGAezaETMP+DsLAXUVdaC1mPdXJkdoTSKJLOFU2CgtNi+/puZPEYEp44hh+FOyIcuuVyztwVxQ/B
BauvR9bQirUjNLNXraU8nS+GScVRdkegXJOItlxfTn+wLeM99ZItJP97C8OcLJIPmuMTZmKwvNXH
EWVamU0IAKr9GV+6Nd0X6HHUfZzl5mxKaNlUrBkaiODuURqM6lQZzvAaARn+zZp1pcz16lncmfLZ
HwyE9uqbpecpEQPYjr6j6bN2ghPTJkgU0juZSVdAEz/EhVwoy8mo3+2XjWN0HkCSN6ht+OwGEYS4
cr60ApHVdOOaiOHxKunabUAeh9WugDdEx1Epzxn7tqUgYv2ikUwA2lKTLovw2g1XNG1t3HlKxfID
B2NczWfbOK6YkDxiPMCls95zoW6ZxxN3U6NorzzYBoLEDm+kHmD/anle2DdWrkq1/QwGjmoo3MoO
obDkxHjBOGrmy4Sj5en8u+xGD1VGxz8WOXKPI0OK2VWnWz13G5ZlNNqHjcCGrz6oZTziPTXWa3Ed
DfAlsUlyYfRdI226ooUIKbi3k7KxsLXRCMqE3ynLxy1IKMoITwmQB7TSTe+sRdvmGvlZJp/o794G
MCGn3FQLJNMfsHWCU3MeCVv+xu63PmVHUSpE988T8x4/JREWkfV5RS4UAqqVGc3/jOk+3UrngLLz
uvnvIxj/0I19FtnWrRUgac+4jkOiLigUlMGp98nJroCGMk+0Y1oIS8vqFxjqQTzvCHOBZm81Ysji
8h7pifwk9EjDJKIvGUUZ3ktILNxxCPYBo07dTQO11IHfLwy8HK9iZIUMCzZSnc59ejEA4MjrM/Dp
QBQJj3BO6/+4SeOHik0xu+Zhk2VIcY3yJrMwTmhCugMz5h4+hUWpXIDJXP6gqaPIxxyBKGlJJ5Gi
3JfQMangkJmGqiVY5u4wi/i6vUcT7AB5E1h/n6ofy/w+JpvyENOksXP+Bp9aEgQvrghaJtdmKQkW
ktnlQCGbcADV8UAeHEDxGGqG23Af/UueM7Bec7bjfSW469Nk+8FTPC4UOCaGUPACHKyoMf5Nc2qZ
t1jyRSTQxoyMuu1FdJwpqOl+9U5SVbxqvF9L0SonndvdY3aQPnORJ18tR7IonfwlGRQTsRuv0/wJ
fQ0kYuk4mpWd0HBO8mBclZxKRjI8+8z4zITvczl2rCnCDFVNzFSSBeTZuQOxn9DtwoJeOKpOp7Ul
B8pyXr2KsrGa9RXTWn+HVLtb3FQg66SIDBWIvBYYcXezjLsvJY7B1ND3X/HdoVnOAN0v5dm2fAf2
ERwj5sD1MMNAQ3hND41C8eXwxdwMLfKDPEkwNbJ65v84akEnBQ7G/oDtgcSLBL5Vg4MZrGdyFHhU
n9DKHPkrKgf2hFmaejat+GSe9OsBFqt5vHFfjiZNcr4clGJkp32coQzjr3JKVVOpIqmXTuOS0bOE
zKSTBJcbZMf9OIdQ39BZlMjqNccnlNxIXeHaMrGPonOb2eermSA1UqErfk9WfdL/BnPSQLiCA8t6
UwU0/jgqWBAl3LnQ8YEMdomAZxbkv4xr/LPA33Y1i3Ry+f5k4XxzNpvMGKCAgEz+V9b5KcPq+zhM
HtQbP3G2FNGoFiVPHreGULOVQRtC6JsUlIEpYhkDqvPRuH6ypNKe4lkFVi97h8olJs5BTJz0diMN
8rURuYjOXY9Hg8EVtqJ9Km7fcA+QdupMLG7oB8HvC1kffstVdkz+wzXD0GhtzRaXjesqfiP2dmv5
5fQ4FQ6MORzbakCX1px79K1h1eS39GQHGfYqotLw75BE5IEgqNatCFc2IPU5A/o+XoV2NuT7rRMa
MIIOyi7f+Vjl2Hg0d6WTO/n3nfF37Rs8Z1Cy601jb2G4Z3X0VxNF2I4sGAJNZWLkgAzBbWmTyYAT
OpoqSVefazMXzW4J6p+xapVVb5s3jri6YnOaavCkF36wjk3AASSZRW61xf0hG8Mc+W4A2nlm6b39
wqU7AeZn6SPBh0P9QNL9X+vevvbpxChx6GT/U1injWOWc3UKF1wW7CHqUx0r2qrUIgnnKp4m4Cn6
4WRH111/yMjxhwPeB60tRFfbfIqx2XZ/FTOyYoASEyZxh5KP0O9rv6flCumaUDq87AD+rJUD0z5z
MpAF75tdEG7Nupq4tRcLumqpcabjLhmNnLrMCDRnjBNt6P5Nd+k+CIZ25Wuk+VB9LhtwtA3YSTir
7ADxTrLjeVdQ/gIKTlZCCPOd6PQkWL8ovRP35bZL+0UhQTGNlmSWXfXvE9X28bCQpfqRNIQESw4X
YVnhmfgJf8FPulrTGQ3K19J0fMP1GaDDMU7oX4AzWInFf03Tbfw449WswddEbO7Y5p5JClzJWPJD
AEC02R4dnYvIP4voieauJeX/5P4W298QPHNs6O4OdUeK0evHADNh59+Fr3YiBS2UiZ9lEvYhUFqZ
JiPnnF7AKBez3UZrPDg5hI0Fy30qbAnq4660/vtz0Re3rg1947sTznqyIgwP1Ra/u/577yV3H5Xc
A5Sxe+jL1MZHwR7v3a1oI4rRbEacwWK5Khrrne0RnUA81VOPT6zJQIClTHyk4OL3Rj8rErJ/8uwW
pWmLdUL6AQUkZ8Tc+ZGIrpe3UgIT2BL3xGa1pzQeK0UjtuBuuX8Hr3M85fZz22W3prEdKXgta85f
mrbHdOjq9RLdvUFJtER9A17ZJVKrT25FS+Pj/aPf8KQ3khakta8cftRrP0JPTspOMwH5BoEQvDkD
2B2EtSTsRK4L1hDE45VC/vPInEYShBsisFz/D5n22hcTtomS45cXT1Y5dzFkFa9zxRkETtucZShR
SUNUMj/LO/aaJcZODcM9v+PTRGGsOli7T0w8fcsEeYZi2xV8sf1sPCTVk6KcypnyUtPfjchmKsBR
xskjThIM+vw9qj1X3fQAMqyRtt87ed7SSzivV0mNVegjNcGjnEDDmNGmVKbobYmDuaEqJMe8fgOD
AvOKjIHu/o6S14m20+p+HyfFgA1qkfYZyL3DYHP5kjS9XJu6c1pwHjT4TaO0sqFlM54VDTyViVAx
8Vwqng+aiGNnjb3T12zlWme+NLckcKvThbD0jlRGMmBqfrYJdmMmVhHd8dKfPHSPfJuYa4GtRAIQ
gG5wprieSeWtmc3R/lwFvrclg9H8t/Tf6qQtaMulXm1t4n9sltZHNICv6EvRngVGYYHmEP1x61kX
krWuMUnVN+c1fxxWH/LX5X007w8+XKufye0QKlUtbHJDzqfEPFIdbr1uit1sLgEo14GWvd1czCvo
gGxzlvV7OcLoi7BdvvYNaFpRWa7Bj/6vtn7oLkcz46MM9M/+Bk534oGAQr9DWJ3V/oUHY7aflI5C
UUkSEaiXGJzDZHDcu/9rXKV8/pTIWsqK8j9gQT9Ajo+2Ebs2F9I1jZ6c8XQx3s/Izg9TPSAxpZEs
CinuGxW57fsEjhv9W+0MmzLBj4/qhw2VzUA0QOZRrOXcDyfbG6BacQ0RtaVU5MzydsoiLUGRh3pe
mZgQorS+mh+ejcJAt7U1OMQuGqqRJ/jgQSOZnmzTPIgnpP5v0B+FEYDANisWGD2Ofz+e5xAxL03Z
eLIaTsSugswsnqi8PPaM7GJAbxvBMCfeY5zWNruxedHxl+Af7OL7r+6e9/MiS9ziUC7lJKf6zdny
t+EnPv3DjtC7zxGpDyIfo4KxoGltY+cH6Z81SgH1BSBARzs5B8P3rPh2imY+TzLAwg+vuRsGxC7J
HA8kJTtnBLDvuR8ets0bBsLo5hrV0JbZcqVF+vOpF9tuIruRXHYF+R35DSZeIAWhIrHifyEwpgX0
2SDtwxWMgtfyB0W/GHyWKOC3UNZuHIrPDl9v60DK+TY/pHfFjJlDz5zOIWsT6PcJLH1stYCFCt/D
+lF/Hf0uOPxFiJZBOd/HjnwNEKCMHRogLOA7oGqKllh7WIN+ARRXqr5FDWJMvW2Dm2HzOjYFlywp
et0nnE4FXVJWa9SQYCdxkp0abV9d6KXb5CWJSDaNHZnRttrrTnll2txkPdMeBI2NQU5AQGTlhcVp
ONOai21UGbrzMGOuQuhE9Gl/7l5S1E8CfjqwV5Quf0527jV0IMwXblp0pQ6f6rBBlglwpmXQQU2c
UGoDfHxyngYFqykPGodtdCmk6qmmAo0JZ/GuZL/kHrY+9gf6cPELZPsX1EeFET7yMFkxTOhy/Jp3
cGIMhF9ygRuob1h35WU1aW30Y3vJOdJNiFF5ElNKgTcLd8euZtkuX0ZZTcDQcbKny740ShUjqq+5
IY+MkqEjIPoikGTd3q81M9V4xsafolQeAy3uAFeTaqttqqQmLU7s5EEcsWvDG1waMvLsQwK18a0L
8Jhg6TZBsb7TY8T+i+dUae2U1nt+iaODvvCzQoQnkTHJPnacrs2kBxRN6uzcfsDaGiF3PFM8qCub
g3eaQsu2zJ8eE+AL6TANCaa4h6nD4P5tiJ3e/ojZZU3hsYJe9GJ9X0fn73gEjJRO0/PUsBMMBv8Q
T/22c9B4mkidBH2nMbn/YkmgA570GXPjKH4axo7jG5JjB1zrnipLxsccWjKlz05JIYPVbV5zRqdj
gdhcBZWwDvh7SoQY/A2QlrHFYa7q2Tpi2CnlougdhFescgCp+b+liDqBn1clVaATTX34PSBtIOZs
NGRligBNQCKC11BjAUJHzVyVWlK7G+pIoPFRp6GzarnGAcA0CDjspIiklkeryou4cmX8/EGwvGfp
XoEb7Bwa/QTUfK80DUQ7jnvnJms8ivjEwvohb80i0QV93pV2Xxig+r1rbtJP4FMMd1PTv2UUxu6Z
Ld+40uhanaIFlz2h/rH/vIj6TBjjlrkbx/K8u5i6BuPJGeiecVjbC4o+fvttaZ8xrq64BPfnd2Zh
NfIeLpXsG8Efp6kUanDgmPma73TdysS4lLtvzh9N2KExt1Q6qz+dAf0HSKB8vq/YGguLQMuOk+DN
hwrCabI5eX6ADywLi8/DRPPGFqgp9cuccX8The9XjV/3naoUv9uMRdaiGSmE599eW8dHjh5uGSkQ
LEZw8QFvZmo2gYL138zx7fWo7Eza7cjUBg28dFh/lkgdXLMhIxZT9F8K50H6Bq7QK7O5IDmLaNDo
gokgpHB9sLYf85MowrcSws8skTRR+dCPOx9KpUojYWVgvy8qfSNt8nECQqdeSY4u/cqi7khFq44H
ZQzyCDZe8Gsonu1yD5RxarVEvnpCa87+Q4f85xqy5NNV87djDDgdR0CGxOHV/RKLt3nXWAs1C/gS
dZ4WA2WVwN8gWZiQoIZHzK9z7uoO3A2gENpBJ17toMtF+dCjX84rHpT4wYuwhAURoGFsuW0ik+sh
EEE0QwwWr2M8TW7OmBk/AQZB3dlyH0knSsYrYWHTyPDtVyIli4tU2HqbTjYkOkrLytzK0QZRkb7e
Cf9DdFKnNpDyx/OViSZRDxutff0meyaSptvhM0CQ1PBLLdtkYIbJfBAB7eoob7xvyS8F9bONi/7/
nGpatvf8srw0Efqfqbv+FIY9NanzByHv7jwF1HvRy6YVmvhkljENwL2ABa56ycswojFRlXB+mnAT
ZmEf1GFUAKIpZmdD7gdL3+iiGZwHTHtNq6sX9y+prOkZp0/OpSN1LNUWw3rwbnBE4togh2vBUISm
ZW9tGXVgpWTTboI+TNZlcOjvGvh6rrCNG7hkD60iIpO7Js+QmWTkdthgHCwLqA1lneYAGBM/dPqP
O1FuCGqIx84RUBAy7fI0MdwMgEWM6euEygc+EmpMYRKsj2LeDEU9d/BGEwL1j9ewGuUpQYPvMOna
38w3DqmWXfk1Uqp1ioNAOQUO02FItXAeH/4NnOezRmBqKrfa/E4BJ5lUs0Dk0/hRbfA00Cq14K96
+G+EhXubrnd1VIWaYCrQKZ9n9wh81drfU/8LJ8JSGut52LfzPee58UQW6/+Mu/RRfpNXfjEsXNKd
y82i3orZxT2iLzzCb65IxISCZQtodeLBFZi9IouMx3bunuCjV6UKOjhTJrShb5GgfpWEBPB0SlSL
mlLgbCRHza7cZazglrP9ugh89yl4UICMzY7uQohcLJzoH6vtDdIf9mbJmZ6lqxyt/mqIwyc22inH
tG6xAzqubIfYyuWGm+jDPfu93nVzGq5JUFl/DUYdbIh2WTGYWGkJ25yHfC5I+OF5hZShj9/2Sb2h
eCQOht0pfqvQNBaKPj3Ln4FMnT0mpV7MLYWc/5iX7VKS2u3P7VvLsVAJLtzIWu2nvzuguUMFx4ho
W+rE/C4Dt3iU/UxXm5gJMphjxwyi2vx8+tUtiSKsYeQJKxcnZWiDJ5Ra32wqzwrqnSYGR08GJsMY
COtigvZTK2tfIw+7GyAvGO8BxWr1TVXkm235qr46XT8RP8TVDkIE33/H1IArrbSGi1d/7F/ORYw4
7Q02c1l1anouMsP4lHgmDhEJK64ht6blKhFPS9qmO6CiY+x84NOpXnCNfIiMNpyptKdkwyOlEdqV
7PZ8m/+0VcNtfdDS0Zk5AKoGQGGY7Srrtmz7wv6GOMkrle5P+4R3WgfMKWJD7rROUnQ8RFA0EQVN
vdAHia7UdU4cnY26LhF23ZGFuphSvo+L5Ih9Yzwd5mT4F4xCXMNgrqEUK9v8EWhPzLYyZQrz8fSK
h7iH78TM//4ds/8ouiwoAJ+fJy+0shU5RThit8IW4J5LTui42P4mP1kIu+c/nHVKmpjLnxNK1op/
Miu9pB46dWa+X/zTpFxArmpJk63BwuqkLi/mL6VcgdU0lBu03AjIMShOKk1ZBMunnBkNzn1Px1fk
FOVOh4CNPs4/lB/TcY9ntAgGaKLlofjZ0ERhGMoLVnkngJCDXXtlg1cUtase29PZFYd+ESh+6xpO
O8hNt2Fk2hSYl67JJsK5ANfkuCXBUVx6aI32jy5TsPTwjDqLMjk1jgDCPJnkoJsLHuX8v0ubF3eT
MoPiRXZoG6t08ODngQ0lctDzy7I5psEFhy6L5Dy+kmF4I/3VQRI1wLcw0GygufTWZ92OjnV2NiKM
3A5y/87UolqULmvKYQJ/BHiDAlf5+DNJK8BM+vlAbWdNYZG/IKVbzSxnSK+P7qteieHcwJnW7A3e
8kpqZo8dmE98SjUXavPNcBoTKMKyZWwxVPFekJCpgcV5E8Si0klfNetUKlvmbGIlUd0cdjHOFSs2
B5VQcCC53dD8VSY4deEfYVIybz2pKE31hcssPoAFmll2NWffHf6KpkvHwHZ2UpgCB6vgUu32gj+d
Jx7t0zhnXxZGsgU6iEK6sqkTRurVYnPSEJDHzZ0N0RFtuhMAsxSPDG36w0CeSHmtLf7EVLVeCqnC
9K7MO/q/ShuMhaSF52OoIL1ZyJLv27CIpM5/SOiY/7XjPFaYh4uQPENiln97XLgioQvMvoAUcqfh
65VeLukD/AqKU572Ihhv7wjALB/8xpAWJ6EMxClymuOWRPmCaXtWHrLVoBb60Z56pD52hxqFS5id
b2FZk7+jgSPjG53iiXb9pthA7UzfBJa52CKC0T8TE15KclRCJITIE151utbeLjIh83di+2nuOpQ1
Gaf706BbFXSmszxhEJPhb0+oSJgfUrFyPtukn3Vib7ng4aTWna6BPKx0cqY6CIfo/XFVgpfiFKuI
FSb1e32pBRFdEQjIcCeN58DCo/HqyK+OakjkbsxGF/f9v6ci5HJ8QlPJTmCWKXZktqJ/CgN7EP78
b4tOPX8V+pDgT3dZJ8Fz+w2vMiaeLODmw6uIZ+MXYUJ50f4scjGDWSsndSYfxf096rEqYazLxep2
tPgAqUIR75SFcJ5VS/E2/eNIdw3rT835ojYFBd3FCA9ysXqx6wjUtSg6ri4H91zRl+u2D/QpOpdp
LvKW4pqEpyMnZog+MYh86BLiKPo6Dgt8hziOb8s29KMk5US7/khQHsGH5eDpsuFJ8gByh/Db8qz7
za+3MYhTW3eF11scvdyWtKb7AzsANlMChzrxpnEMy6RgqbfgqZdGJwKW/KzOnExFrg5d7e7kF7xp
49FoHXyYSuFYKcB/0msY41J8XLOFeXjF8rvHfOHfT6OFz/jxCzx8TumSXRgKCz6cYG4Er4eOI8PE
DTV5alZZ6QiPipCHELH/nwKFZ/dvowkOhCR7HV+/3E3E/6+/+chLm42Mb1U+gaxHfYsp85G7x9CS
6QHW/ibR8L1U03g50ij0EvXzAWlY4usN1qNt/K6jmHdus9gQ5955YAqetMuKbbROx4eWNL/QP1Kv
mXExE2tTVZC2qi9slqzWEnjYxLwRQ/l3d3tv6UZtHea9fJPXCnPvE5iuJQDhZOndzym67jKkvWaG
BG1qVZRRQDAgCicyAKOPyUKJoFChLKLdYib7CcGiZI0kl+g/R47WpMiwkfi5bKMBEcADSd8OA+ka
Pq3JY78IzKXybRzuVH/gRc8lq1JbO6zH2awHQMko0gN+sObVW5bx4IK0QXGE68yB9BpCs6tcW5Qy
ONSSlMSId8wXBZHPc+/Je2KhME5LHumCmAfeian1EWAVgPZzg/8B6QH/d2TZkMXZYGdtXiIT+Pvm
nE+9khA/hv0Dpu3L+lcY+gbhjAR5gsw8VZaXl2QbD/Fq74VcVVLUTLxz/AfbRTWwjOJ+s86s+6sx
V4c2w848ht6gTWYNv/snyCTDYei4v52wIrzF3jCOXgqBfF24TtBdEIJhHaKrQssGUNRstGWxi6AA
2meGzou/Q+/w5om0EAgwpvtkuL6KZnRorDhLhKMdZt0PxRprLLfqCP2Ypv8weJpPuSba5Im+5+e+
6aiYNGZNOYYir+nkgj3Qvf30q7uTP647YHaJqRe7ZxEfV27QyEscV8t7ulunhfbmRjHg4jrlRcwr
lTxQ0XsrEtmpC8OEW6tCSdGcMfh0SIUDVu6N0Lo/LEhGHufKZpAkhGjqKfHtekjMgy4VTS4DZbi1
XWcRuwDHMOUmnvpHm8S3VDY20IQuuDSF1l033VGBe3UYGcDwxcGMnS0zKtVXbQO6edkEbe7qs0oA
6dhNG0KrXBpmiUOjka9NzcXBgWSMQvVb6L2CItpCH4a2MInOgav9crOk57YulP0ES0lZtjm0A9dv
bjSbiBmnsShw15bpKge+A2Fr25HlTlRAmANT6sXI3J9QpGyWZFYNhktP9BgCf6HWROULQAOjxjvq
pl9oMUmD0oRxo92fTA8ZPQjMFQ/u3/atAEa7p9bM409yE8WQicR2qTQo6YIfJnm2G8yu4soikdB1
em7W+JFDWbfjma70KfsRlXmFOppgCfrdGNiPXP1yBhW0E0Mb7n8+gd0xUfBrBaIL2ICyjtfs1dl7
XXBysUnP+nxqcvUCSKLY7RQb4KqiKhBEfLBk2lL27zctxUb3zAsCDSMr7+5Mr3ZX/NH1O/8ai9oA
gqhCYtDeqAb+KYABdA4SBOFuZ721/z60pw2iguMY/RRd/zlpwHhyJ5qY9H4udolv4qc7gu3pAYcF
8R1KtZKeMuU8MgpTH0uVoxv5C7IvGsYOKWwqRy4ja1BCOH5nP461CRW+/sxUv0MR4zi2hEQgJFuC
GQLEwLBqPTFhUMrWm6Sj/8bwyFUAJhzJNvJlgoFRiq2DXx6CFXO8fR8RnOaOVUy2tce2jezjJCtV
bIalUQzM+jdC933DR6NIGi+aG0FD9HdKU44SmLhQrxJTg6SoypKUQuek35yu6VWeTg3/RHD6qyzn
rIjikpPykg5Wmot80u42B/Sr39TLvSGquAloFJUySMi55mQRWlyM1hMEwrq6KfMKDKkveXA+ZW8Q
NMuxg9oCnCnKU9wqrusRVBFSPkBl4kr2PusPJmIigvmsTb199y/mcdcvhOeOtE5MRQtOe3HelJqH
dGusQUyXRdKIU+ZKqVARXa6Gh+OmkHpIMjE10MBdk7khEkmfwmD9Suedgvi4KBIt4ym94/0LfP5/
laSQFOc1wjAnzZfUnrMr0js3Z7io1++q+uFV36duTjX8Y/jpsWDmDJCb1yE+vPCBBoXjKKEjwvfT
JBoamKz/OhKXVlZlh3BvDTuEkC3o+lOIt8ZPkln2XqwpG1bl1NNPtazeZvLOgtbEerTdhDfKCUx0
4iLqKGl42k95VG8ciob1cZcnRusLhPYHF2A36d1mJZM77UGn3zX141RWrpa75SzNmVANXAE0bQiD
gn411wKg+sPlCt0VP9v1eGOLCFjYWMS0fQM2kxLZR0YA+Es0R0dzFHj5xXVOkcsiuoOzfQJie1G9
BCXM00VkGuH5lVo7VSA2ZZP9NLWASF6mbEc4CLmx+pko7b0u5Os0lbbN4zlJ1ReM8vC8iP5VeFZ4
z00Z4RV9QnpiOU42qw2gYKyczaWuT+gYdu2AYppJxYWPG5jcLQniWsmcpvR+e+CDzkwxsDKdU6cj
2wXRtcbWGXPMIvnMYmpipoennbKmZDaZ5782RjTSsNcxqscnBKVgVzuX25zj8ybP8vfDUQd/uihf
3Wbu2fL+BfEoKmhmKgetjIA3YZqRSBuNWrrdEBdLmPCyXTqJVwOgTL83Z3OuZeG9J3H2kGPZQC78
i5Q+4hbCwsrIddNLCpqYra0MTKSsVh702TFM5Lin4InD14i5QnzY9dEJ4/yNvKltPN6Yqe4+o74f
azt7UScFsOFtu13tRgiml4fMfxijeAUq52olR3BRTb+2gXfNzb1kPD2G+eOoMoVU/hMRJPAChkye
wh0/CFnUA5MhJcOPEiVXDeCX3B2r6zEUoOWK0nQTbeWrTlxCXjEJSMXhJUsn0AJ6oNf9NMPV6Yec
cglkJKfEC4oJHPnMuihosjjq3oY23LlVbVA+7Nmy8W1VqnUsbKbUZYFRHXgjKKoDrH+NNGhvIEFI
IrDcXyFQXOlzrV5OsHiHFs+UldvKo+WKbDRRnYlWFRL/oO4dPuxKyfshv6LwKj0blNyCHVOh/ITg
ZoGuRFfQ6xBvx24F7T0hUasHKumPnQfBVoKQLrHb5FTwd3YUEJx4DyvuqhYXtOWNtd6S8EcEmndB
qQ+wHBKHLidDEGXS7gdUyIXl/ybgeitlPJBVUdEuW8qDtNhNaAhYQZ5V2u2DLAV3RP68CJBDi3fF
eqhdFj2Arp7KEp8JGO9bmUbPpeo6iXIx6O+O0I//x9CJrTjioFkLI6yjQ+mbQ/IqhOmLomhx93j1
1+ivRlCV+HOzSbpRACpnluZhNJIhx9CHEQZ5bqczw8eYcSLxo6jd8Kn7egMSTN4DVshbi4q59pMR
9HpIBe4+AGSqoFlQhvqu3LXMAOizQ/HGmiqKnVrbWIlhuI3ocePBUW2LL8WUefA2R09Sc/aaqjC9
BaIw8dKY2kAqPe6PX5h6THlxjwE7JmkVmNkA+TIk4c7k5jFuOMsSBLyddyJ2X5cSh5ErMXx/cA7T
EblMYwvq0VGWoXOLlGjYSxeaCDyJegFHYM+15v1aoaTm2YD2wEobAGFxGBHYcgER0hM2yOa03PfB
y4QKQuonlvXpDRVzOv25yIri/GcienkiVL2Y8pRfZnOFNDfRue8pDlaDY4MhAadfX0yudoKU8i4A
eRJAKZSEWlfj3zgFKolrQVNCQHNy0dZ+KKa4wJotjCFXWHz1jweCWmddXqYZkkGhvhwVuSEdqENB
Yu7MDbtDvYe5A1HDFxSJDzs+cPNUNoPCDDJkDFykcUJqqwXJveobKTDCQCpk+74EWCqwpCLljnzb
IL/HGO0kXhozlnZz+2yaR9G5QXZsXC1GavBj0yE8HiLVr/3O711AfZ0tdiU+61nsZewxQnHGFbO9
BUIHLLDQbxaM8E8v4uVHgMJ15pyGHT0wI69LDYWO3cNU5SXV5pC4phF9nO0ZehFlRkgHErkDG4Cl
sc0N12ZSNslMh2fN4FQiUiMMng/E8WMhamUHxRbgQ4IYWLUUoIzJhiJ4NhM4ZOOXtAj4OA/rdWMk
2Ejz1Q4TaDxKi/y6DzIJ08dtnLJb+raDr0KMOBs9/970UC8tmPPLKEJuRDxWl83xBRcfMtAc9fy6
RkrcTloLAKWaHg+BGKGzoP/xN1WM2cdHbK1BJ865WThpKiayFFAHwYtCyRh6GVOQF3o1cjEbUlLy
0EsYI7qbJEzrNDuOrRKRF6VX7gHFBtWH/VopHAZd7hn6GcxY6r0KpaDRobYFqBlGt8ifqnzctD8G
PXnohB+SN56YbAtmBBqYDVadOPgLGHFeS9OaaO2/EMk6G7Z01WL3I3jnj/W9BWU/t8gPoLcnc5Me
8PuZvW3xdKvERxypbSZ4OK0Sx+NPhu42NPFduXQxPI//Kupn6YCHMToFg+RTJw/iq3pG6bdYq7Vb
iigAWFGtp3cRmwsbycfZBgiCRnbgbQ4OpC1A+dqDuTNHuoyb5zpUlymt0YV1iQ1BjCHTDBpvIo4D
MtaO6flUu1pr1JX7K5NOAKTwtv60/McbYc6b3AqiocRcfYwy5785gHCLOOnnD3j0vVUTF1hM5tX1
ukXOEWPFd490Iqocf0Lrb2BTucDvEDEpQ+gCHnF46taz1rQYmf8vtQDGUV9nnu0J3Z1Nxdaqe0Y4
2k/ILwZcrik+Saymou7wi2kIuQ9o8TQCAezsVWNogKYVulVTpqazgAL14CLIrbfg+H4kz4Tgvw/N
A32Wz3MTVG28WIb7MITVGh9KYCzktTvt2Z8enz3ZY+MyH4lb8QfA6UL0OcxNdb3HhMveWwqgCTGN
5wuO93JcNRGfGpjuch5F8lzD2iRVUDuKHnTCbpfPiNxh5pzGaHWeAM+W8YFTGR9yvnNLC6DWZNZg
Mxwk2z+eoshyMl9xuA/8c1uOHYloATEqWL2nG2ipCU3BnLvdYkZcUxhMnV4oMP6/w/WgGFXETqSa
vEj874Et7jPgRed5vZnvqYHCqyGQU5n3dC9tegj2ibsyoA3Pk82bY+iA7UZIEiwVj/ahMLQrCO05
riLeAc3t1DbkA3dCSDwQojB3Kt1HsgmRCwo6EiUDPG+ES9PLC0feV7AcTEs/WIsWVaiEYbuxpneB
cd00VJfXQkD2LJ7HB5O65+hYjOLAwZnLY0R2KsdSeShMjs3A6996Qb2NV40d+0ie8cge3sHlqMeh
nXQyNNCUG+nqK5/ITHhYTFk1ovuvg8L2D5oH9PkE5fI4ycbT6MESnxasdCHvdX6dzTy1ej65FbjR
ClOPRx8O1tgISUZyxaGE+QLh1/obWqFwk84RkyQMhU0hVK4ztBu33tI/4hzCEnqx7BQ91CC30zGC
Y8RMwlHSvnY7JOnjWGQHoeVTq7wCo2MX9I0XBZukY1fq2dDVetDLrT6mHUGFdJIs++bGr9Eh8AXt
WtZMLdtKbIsordrEeakzwD+pD7aDNkuyBbNR0LG9s7kgnVfxa6vQBexSzYUU5gIMBr88wpaxbwm+
qVpL5QS6+4VKUU/GYbGvAlD8tStEgrU1MWKl+LsY4HWo6dWz3JQnMsd2Mqn90Zc1MjEPvABCFSGq
2d51drf0fFQpI3a4a/SnIU18IfiA4ed0sGoBY8E6LlRezS1FkVQKpIfKvaHeF8YE/a2ZlX20IYKN
u77t7JUYd/hpvpQev86uwP32FLF07rp+vyqI3X68Qux3sqvg117dRIBtdxA/9wqMKR1J71TMkBOL
FZmpRyH7G2+oHu+xADXz9vKSoZgP2rZiIYmRm2b/+na/wwlbUvTVpsVK3thBrC2Jw/vDJTkqX1QO
UJ3zxRrjdzcWCmNqnlzmMG5v8OFdUMmA6fqIQjywewwOUAH71OquTEN8rzXpzr/3Ub4Nu1U8DH19
JReaxWjdfS+tvejRrblris7R8+nvJ9Sd+UoEYyYO6TeFeL7OE2B9K30ZPcsH4aYDsGKZ0OwyXN2V
r6qX4geDxXHbGV/p5beUV9qDKjJ95dJO15HYzAZttXEIdAB+eRsKOALPyhFM7Owa6KVuvDbu+LLm
34YIV9/a7SUfHgBn4WGPSLM9fC+yD8K2ZxeWqVwOGVGIgLCa3oK32lAHbXeGuDYrhCwoz+R4nslc
tf6u8BqT2toPVcyIGJu3D6Cqdeb8BLaLyvVFJ41WQJlW47RrCTjlhd2uI4+unsgILTfKcKLnc/vT
4R0X3Lz0Nz6JBy1LdIvHEfL3Y9neCJNusq1yr7GGZPWUHWXVcvzswlkb4GH/fOPQEy4WPL1+0VvX
X8ngYaG9u0A7itbNHJwWa0Vm7oNB+VtK8NiyDLZx07KZL23eqqTL55z6EnHhSg4M0E7/TE5M0kLl
GerV3dF6aAPbMEWftX1rOjU7Z4fx9z6qxSGr/PXWOvgCmQbFO+EtiQyP48jnik4Qci1EgvrqCKF/
EF2iEQr0AKC6k6KFW7ahkIlMHZMzfitfZpKtDGCthJxr8xS5RV+YTsFSz0OBcLD/Qq+Ixzl8uiXz
SsK3Ob2UKPzEICzlV08+xnEio2UtgkKxhLjKiIvWDNDFh3g3ysOj6aZQm1zaT3J1djwZ5JQGMZwc
aY/u6bih5C4Evt6YBQEBdodVntYLWADAZEFZ/NFyw/KfUV8zA+uxVrStW2roLky4Th5yGglerzFu
ZGKmihCJz2Q5CUowgBsw4zE4Pc3IKkvO/Me1h3lufAPRA446RTHrsDUsYHvv6qo9Ooi8fXtWdEsO
aCrJ+NFte5dDRPnkBi/3H1dTgHEMLzxWj5fMS7LOyKYenTMsdtKTldnsrm6AA3ec4aCYu7WIZwle
uXAqfOyiXyGwr7Cv819rCwcNqbbeMx4JOX1WrTSW9lT6iMvuxE6nKASFnoi4zkeRq6i9Vht3GOAN
9ReL1/B8eR3qMKr1YGQgCJPUXV6KVMJSVa1xoSL14lYhXaW4ngAV0jh2ASDlPq2OkiXTA3aa9DC2
HzQkbq/TXq8H0Cphl43f9VFJMOhmFvx6XVqC8HMQcO4OiY6LprXYC9IkcOyt6cNyi4rNu89J06eJ
VbkIgxnMek2g7Y/bCyfELpMBw+bJPjSyp8CGusflAlHl832pRlSYMqTfjo0Ww/CD0SaZ71neXF6U
H38fgsblMG/u93FaZAUg5HmaTN6qzRiM0MqbAimHrcPZYb8F24su3NbLUbRIQBDrBjtdg7XB56b3
rMandwoB2Isv977ueA689JavPk7ERrMNs4z9Bl4M4zWtBzFIjSTvwNewsnHnwfxkZ1KoP0wykq5M
0z2RBk0XpxSHD5ihkAM4QT5tJHc5exh5uGoOwLqtphJb8ZWQbo0SNCP2y9rDEVzGnY1qmcIXdZfB
uFGca44rJAND4tGA8Nghc9Rk3Yo3h9riMt7alC1prmZPJBySI5yzoFKAyYGpa3TqtiNEPq8sYTX5
RMS2UG3+C1+vL+/PzuWDZRQR1HePVkWMZ2gggrY6cIc3s7E7nksfxC5UVMlAgAzFV+erk6BKXNLj
n+0zhoJdekhgAU8trOGLMX5jO1cD52VDB1ozQ6Bbh3Mp35XbFonDpbCxf8+xVa0fkXwnPnR808i0
Sghk9c1xhaP3UVjb+8IHX79zqVRxYiLc2AOaGp4GEdiJm4HlFng0ijKdGyL2rhZAPJ1CGh6boVbV
G+Xdylbw8YO9xrEHuttJVwRnlIbiwjCy382GGT64w9MJKMkc4dnvNFi3SWN6IW8uccpyZzkCRJXl
bgzyCAckKfFdLCz1cPCJhO7GUuoNLzWk062tzekUiXcZwL5V8sfWWj9lyDMEvJf2o7+VgkicfDOv
nAYZtvFcCF1NE9bdzivovmI8OAZPx4HLYa0yR4X4rYb8gY2jUlVFruHcSe7vot1luZuEAEtOAVIy
CMgVxCamw8Pc6eXypgrDufuFwhHtKZPIp6lrdYtiQWLDK7rpj+NHFv+fNdXcIwp8kLbpemBjnyr8
QigjieoUMygDVeAkpkAd7dZgCeSJQrgn5ZU0oyALiIpRTRoyLhUAPwttxxOzuwMFZkv6tRGaZhhE
FeaH18n1fBPDpV56CERqQOJ0vntZfl1EPKZRqyggMco2wXQ26dEFNSDw3fKBDTNR8zPsQE2V+jhr
SLwRibQx3HqPYw4qA8wkNpjTqHiasvQHba6q+AyIBaffyta9SbSTUrMcHn/RDlLTYUfTaYVGtYlY
ovuuwjN8foQLMCgomdwkGMGt68kiL+5Y0nZmU7HGqumXtdrKWVU0MyPHlizxpHBobWdAttjGdc4L
JOOWWBvSKT45ZVi+ni09Y+U+dFN0rcmKDWJHbpLIMDO08GtXHWZAhgqDkELEFkr1ygXHZyU/tWeb
NjHR9rOLEIeEjTIshk5O9Nx/f/f32q0ggB9MD5B7EY6nQSv3zbuVDGAd5lJtnZrGRYnKyn4fpy6d
frvyGhPTPDB3kLTGJCNzsLbfIgpu1j8QQ1LkYzyeXgK2esOmkmjGvUPdVBgE3IrttvqwgvZL/x0e
WrWs4cLc9wWY8Q0GUXgYK5GTvCnHTlkHIhuOvpqE81odiB6OeX19J6p2KF8GYJmslN2VTqkIx+BL
PgX1uin2qllBHaSVy4JxanMsHc+Vvn9eX0SObiNCJTuFSojzFumz9CrJhcki9gzMhbiPtzbTu9Y7
O+X4YKqVPD4C6VzsteOxVpBhDmnpCG7fAy1DjFE0gZzLRlPc4c/e0dHz7yN/u/ymySW834pVqsEh
EnF7mfgRbdfMDa/hwdF3i/23pgIsW2+RJYZjC/Ess0k+97UcUl4eQmZsbLkSE5gEozuFiUjwz+EG
YCU6LK/M4XTZE1oB+Oib57YvhUNyAMUNlT9/g5RZr2Kal3apfDobtNPdRbdhX+Ya9olsW7mMyj6j
jaoLG8AKrBqMbJHSCeBP2inlc8HdrBCPBAP0TEo/lAI0pTuPeDxd7ZWIwSxdzdFc9nV8O6sNwtV7
2VzxuBT7jSoDzjQOt6gTdaBS36IZWtCBeB4O2Tol1UZON2XMkT+OB/vPGktOCudNdK0LCuwf6ha6
qvaSgW2ulTCy7BN8V6w/JRO+YO+c+1LhE/OJAUu/G1REMbNJFuhMvvqPxDUnan18spae6JX3Unvu
2GR4/Rt8wnK5917FH1JFrsyuapFSIP0eO4RN0NXisO//zL7Js/ADbhFqSAJtEKF+bhDZCR2Pdsln
CAebYGg3hC+Sz/2SXd+L3rd39sf6FA5fGOW3k2Okn8Lv7rpPjnLIjMGW1Q8fUiw5G+F4k1qavnlJ
yTA4Srajr49ulmdL2KYU236FHTtPxipYJoDtFeh3oPdPc9LfbHkRiZ8vungJPlzqyanPiHpTqF7K
W9d3LwDjWZ+kOZnLpOy7BcgDm1Gc8Sb5PIWKfkrI9snB8r8rfHOFEV8IECz+HwDgK59wfTFrIkuX
T+smTEzd1zhdSOhfK4Wwa0x0XInQlf1rsSByzMCsMVDnNQf2DWEtjtTRQ0U8qUpxbrK+0uBuCe61
5YXK13c6y6PDXqPaxAE3U/DkiJDpCYvcGJJVju5sZLKKBtG9JsbA5QVRLI+XBf82Q8uJ3gogrsDd
wGzgMvdCuJmw4zV4YaT3uetFyNmWdftnGXu1qHd+PWq1EjuuyPsWLb7qsF+w7tPgef7+/SxcCdG0
RjoZr51IzRRL2Tstro3I6dpe9QXWDdobMt9feSHKhzk55L504rLhytb+Nuxm7qgQsAY0iXBuvS7U
q0pFb2e1NeY4ZqsJTy+gnmokrKPPsaTg3FdFku9zWZ6qWt35YpaT0x6bdYx091Bl8+o44PtEvvTp
cjIyrBzwEF4lHc5x+/h4Kh2oh39vsezyVIjixo6DHLc0sLFOihKBo8FkSwZ0F6iNoMLvTh8cSnzS
dgh1hwjq2nlIrHf/7LJw9cS8rhCgBuJlyWjxjOTPi5typPJ3hK6x1D4s3oWXIADH/A2gjmZW+PVE
ktPxlZKBU70wDeGe96dMd8E/WYUFCmwQDB+LuLspyW6LV0pOn3L7k9t1TKjhPDOhUqrwqTdERI21
ZS4RpXFaV9k3yXJvQ2pg8GebEScxtPHTfdimoDrcDtowp4MZ7XTalcxB8jbiySp4vDeYNUTEFQUJ
wRqNqcwuDPpT24IV5qOgnxn6A2rzKrXpmYouX6yCUFf1P1a6mTwfKEG0VabyghgHApBaZtEE04LR
lrjEBmyUQBAAEZtGZnymqeYeABGpRJY55/1T518lG8OcVJDVOJ320e2p9EMlW6oK1Mz1jWRJWQYN
QIbPPSdapkJzve5ygALyGcH9ja2w3nba+a7Vc/5+aTHR/xIZ/GkhfJgeRY0OZLkdppEvPb++73Ex
el6iIAqirSFE21UVqi177ZrIOpj4TPRXvx16jkp4rRdGsgiSv5Jq5EGGEvHCNvm6IAwd5PI0cWf/
y9TDEwMQe6akw4k4FfcQP46yONpXk3YkUeR/mlFlGNOChzW0aHRIpdk5EjxwnRE4gcm8zW0bIueu
2A8ZArtPQxKjzU1ztel1dCRo3qzndpOdn0vYPUfr5mFWlgw0QIebROgUhYX8bx6nVax/a1RNZs8o
4VTEwgDApWb51Tht5rl42XQ1
`pragma protect end_protected

// 
